

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9585, n9587, n9588, n9589, n9590, n9591, n9592, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9607,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20037, n20038, n20039, n20040, n20041, n20042, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405,
         n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
         n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
         n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
         n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
         n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
         n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
         n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
         n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469,
         n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
         n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867;

  OAI21_X1 U11029 ( .B1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15301), .A(
        n15269), .ZN(n16026) );
  NOR2_X1 U11030 ( .A1(n17991), .A2(n16320), .ZN(n17633) );
  NOR2_X1 U11031 ( .A1(n14204), .A2(n14190), .ZN(n14192) );
  OAI21_X1 U11032 ( .B1(n15593), .B2(n15592), .A(n18483), .ZN(n17158) );
  NOR2_X1 U11033 ( .A1(n12227), .A2(n12229), .ZN(n19192) );
  INV_X1 U11034 ( .A(n17988), .ZN(n16646) );
  INV_X1 U11035 ( .A(n12735), .ZN(n12724) );
  NAND2_X1 U11036 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10438), .ZN(
        n12736) );
  INV_X1 U11037 ( .A(n10090), .ZN(n16839) );
  INV_X1 U11039 ( .A(n10962), .ZN(n16910) );
  INV_X1 U11040 ( .A(n16950), .ZN(n15510) );
  CLKBUF_X1 U11041 ( .A(n10239), .Z(n19057) );
  BUF_X1 U11042 ( .A(n11235), .Z(n13416) );
  NOR2_X1 U11043 ( .A1(n12509), .A2(n19045), .ZN(n12521) );
  CLKBUF_X2 U11044 ( .A(n10256), .Z(n10271) );
  NAND2_X1 U11045 ( .A1(n11052), .A2(n18590), .ZN(n10811) );
  NAND2_X2 U11046 ( .A1(n10097), .A2(n9707), .ZN(n11267) );
  INV_X2 U11047 ( .A(n20005), .ZN(n11270) );
  INV_X2 U11048 ( .A(n20032), .ZN(n12030) );
  INV_X1 U11049 ( .A(n11236), .ZN(n13383) );
  AND2_X1 U11050 ( .A1(n13432), .A2(n11148), .ZN(n11201) );
  AND2_X4 U11051 ( .A1(n11156), .A2(n13638), .ZN(n12130) );
  CLKBUF_X1 U11052 ( .A(n11240), .Z(n12111) );
  AND2_X1 U11053 ( .A1(n9781), .A2(n11155), .ZN(n11195) );
  AND2_X1 U11054 ( .A1(n13432), .A2(n11148), .ZN(n9672) );
  BUF_X2 U11055 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n19681) );
  NOR2_X2 U11056 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13433) );
  NAND2_X1 U11058 ( .A1(n13383), .A2(n20025), .ZN(n11936) );
  INV_X1 U11059 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10136) );
  INV_X1 U11060 ( .A(n15488), .ZN(n16908) );
  INV_X1 U11061 ( .A(n14002), .ZN(n14000) );
  NOR2_X1 U11062 ( .A1(n12227), .A2(n12234), .ZN(n13718) );
  NAND2_X1 U11064 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13978) );
  NAND2_X1 U11065 ( .A1(n9592), .A2(n20005), .ZN(n11295) );
  AND2_X1 U11066 ( .A1(n13418), .A2(n13438), .ZN(n19987) );
  BUF_X2 U11067 ( .A(n10325), .Z(n10403) );
  INV_X1 U11068 ( .A(n18865), .ZN(n9828) );
  NOR3_X2 U11069 ( .A1(n11045), .A2(n11070), .A3(n18434), .ZN(n13971) );
  CLKBUF_X2 U11070 ( .A(n13265), .Z(n14089) );
  INV_X1 U11071 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19732) );
  INV_X2 U11072 ( .A(n10264), .ZN(n13720) );
  AND2_X1 U11073 ( .A1(n12214), .A2(n12216), .ZN(n12601) );
  INV_X1 U11074 ( .A(n9732), .ZN(n16659) );
  INV_X1 U11075 ( .A(n17092), .ZN(n18024) );
  INV_X1 U11076 ( .A(n17549), .ZN(n17537) );
  INV_X1 U11077 ( .A(n17643), .ZN(n17614) );
  INV_X1 U11078 ( .A(n18631), .ZN(n17991) );
  INV_X1 U11079 ( .A(n15781), .ZN(n19934) );
  INV_X2 U11080 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18604) );
  INV_X2 U11081 ( .A(n11428), .ZN(n9650) );
  INV_X2 U11082 ( .A(n11428), .ZN(n9651) );
  AND2_X1 U11083 ( .A1(n14469), .A2(n9758), .ZN(n9585) );
  INV_X1 U11084 ( .A(n15785), .ZN(n14015) );
  AOI21_X2 U11085 ( .B1(n15004), .B2(n15003), .A(n15002), .ZN(n15230) );
  XNOR2_X2 U11086 ( .A(n11962), .B(n19957), .ZN(n19926) );
  NOR2_X1 U11087 ( .A1(n12227), .A2(n12228), .ZN(n12291) );
  AOI211_X2 U11088 ( .C1(n11037), .C2(n11029), .A(n11028), .B(n11027), .ZN(
        n11032) );
  XNOR2_X2 U11089 ( .A(n11956), .B(n19967), .ZN(n13526) );
  BUF_X8 U11091 ( .A(n16908), .Z(n9588) );
  AND2_X2 U11092 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10437) );
  INV_X4 U11093 ( .A(n13977), .ZN(n16929) );
  INV_X4 U11094 ( .A(n10447), .ZN(n12901) );
  NOR2_X2 U11095 ( .A1(n13544), .A2(n13543), .ZN(n13556) );
  BUF_X1 U11096 ( .A(n11091), .Z(n9589) );
  AND2_X4 U11097 ( .A1(n15425), .A2(n10299), .ZN(n12754) );
  NAND2_X2 U11098 ( .A1(n10054), .A2(n12396), .ZN(n15995) );
  NAND2_X2 U11099 ( .A1(n10238), .A2(n13720), .ZN(n10325) );
  NAND2_X1 U11100 ( .A1(n14406), .A2(n9590), .ZN(n14438) );
  NAND2_X2 U11101 ( .A1(n14214), .A2(n14216), .ZN(n14215) );
  CLKBUF_X1 U11102 ( .A(n14996), .Z(n14997) );
  NOR2_X1 U11103 ( .A1(n10939), .A2(n16191), .ZN(n11129) );
  NOR2_X2 U11104 ( .A1(n13844), .A2(n11564), .ZN(n13892) );
  AOI21_X1 U11105 ( .B1(n9681), .B2(n9634), .A(n9590), .ZN(n9631) );
  INV_X1 U11106 ( .A(n14479), .ZN(n9590) );
  NAND2_X1 U11107 ( .A1(n13827), .A2(n15397), .ZN(n13829) );
  NOR2_X1 U11108 ( .A1(n14896), .A2(n14897), .ZN(n14889) );
  NAND2_X1 U11109 ( .A1(n11962), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11963) );
  NAND2_X1 U11110 ( .A1(n11526), .A2(n11525), .ZN(n11993) );
  NAND2_X1 U11111 ( .A1(n13354), .A2(n13355), .ZN(n13356) );
  AND2_X1 U11112 ( .A1(n14192), .A2(n14177), .ZN(n14179) );
  NAND2_X1 U11113 ( .A1(n11437), .A2(n11436), .ZN(n11438) );
  AND2_X1 U11114 ( .A1(n13151), .A2(n12608), .ZN(n13219) );
  NAND2_X1 U11115 ( .A1(n12399), .A2(n12405), .ZN(n10786) );
  CLKBUF_X2 U11116 ( .A(n13633), .Z(n9664) );
  AND2_X1 U11117 ( .A1(n12364), .A2(n14852), .ZN(n12384) );
  NAND2_X1 U11118 ( .A1(n11416), .A2(n11372), .ZN(n13424) );
  NOR2_X1 U11119 ( .A1(n18586), .A2(n20825), .ZN(n16688) );
  AND2_X1 U11120 ( .A1(n10283), .A2(n10297), .ZN(n12209) );
  AND2_X1 U11121 ( .A1(n11405), .A2(n11403), .ZN(n11304) );
  NAND2_X1 U11122 ( .A1(n12213), .A2(n12212), .ZN(n12214) );
  OAI211_X1 U11123 ( .C1(n11360), .C2(n11153), .A(n11286), .B(n9639), .ZN(
        n11287) );
  AND2_X1 U11124 ( .A1(n9810), .A2(n9706), .ZN(n10412) );
  NAND2_X1 U11125 ( .A1(n10266), .A2(n9714), .ZN(n12437) );
  AND2_X1 U11126 ( .A1(n10792), .A2(n12521), .ZN(n10290) );
  CLKBUF_X2 U11127 ( .A(n10476), .Z(n10752) );
  NAND2_X1 U11128 ( .A1(n11235), .A2(n20032), .ZN(n11275) );
  NAND2_X1 U11129 ( .A1(n18017), .A2(n18009), .ZN(n18452) );
  NAND2_X1 U11130 ( .A1(n10767), .A2(n10264), .ZN(n10433) );
  CLKBUF_X2 U11131 ( .A(n10255), .Z(n10234) );
  NAND2_X2 U11133 ( .A1(n19742), .A2(n9597), .ZN(n10766) );
  AND2_X2 U11134 ( .A1(n10216), .A2(n10215), .ZN(n19742) );
  NAND2_X1 U11135 ( .A1(n10156), .A2(n10155), .ZN(n10239) );
  CLKBUF_X1 U11136 ( .A(n11293), .Z(n13186) );
  INV_X2 U11137 ( .A(n11930), .ZN(n9592) );
  OR2_X2 U11138 ( .A1(n11264), .A2(n11263), .ZN(n11930) );
  NAND2_X1 U11139 ( .A1(n10085), .A2(n10229), .ZN(n10056) );
  AND2_X1 U11140 ( .A1(n11163), .A2(n9699), .ZN(n11293) );
  CLKBUF_X2 U11141 ( .A(n11453), .Z(n11892) );
  BUF_X2 U11142 ( .A(n11195), .Z(n12137) );
  INV_X1 U11143 ( .A(n10858), .ZN(n10944) );
  AOI22_X1 U11144 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10152) );
  NOR2_X2 U11145 ( .A1(n10811), .A2(n10808), .ZN(n10867) );
  CLKBUF_X2 U11147 ( .A(n11310), .Z(n9665) );
  NAND4_X1 U11149 ( .A1(n10048), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        n11153), .A4(n15547), .ZN(n11428) );
  INV_X1 U11150 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18612) );
  NAND2_X1 U11151 ( .A1(n9600), .A2(n9821), .ZN(n14937) );
  OAI21_X1 U11152 ( .B1(n14035), .B2(n14034), .A(n14033), .ZN(n14038) );
  NAND2_X1 U11153 ( .A1(n13996), .A2(n13995), .ZN(n9600) );
  OAI21_X1 U11154 ( .B1(n13996), .B2(n13997), .A(n9601), .ZN(n14035) );
  AND2_X1 U11155 ( .A1(n12486), .A2(n12485), .ZN(n12487) );
  AND2_X1 U11156 ( .A1(n12582), .A2(n12581), .ZN(n12583) );
  AOI21_X1 U11157 ( .B1(n15085), .B2(n15410), .A(n9911), .ZN(n15089) );
  NAND2_X1 U11158 ( .A1(n14429), .A2(n14541), .ZN(n14019) );
  XNOR2_X1 U11159 ( .A(n9698), .B(n12157), .ZN(n14132) );
  NAND2_X1 U11160 ( .A1(n14428), .A2(n14438), .ZN(n14429) );
  NAND2_X1 U11161 ( .A1(n9826), .A2(n12406), .ZN(n10060) );
  INV_X1 U11162 ( .A(n14978), .ZN(n9826) );
  CLKBUF_X1 U11163 ( .A(n14187), .Z(n14188) );
  OR2_X1 U11164 ( .A1(n15341), .A2(n15312), .ZN(n15305) );
  NOR2_X1 U11165 ( .A1(n14947), .A2(n14948), .ZN(n12475) );
  NAND2_X2 U11166 ( .A1(n9623), .A2(n9622), .ZN(n14428) );
  NOR2_X1 U11167 ( .A1(n14947), .A2(n10034), .ZN(n14939) );
  NAND2_X1 U11168 ( .A1(n14969), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14947) );
  NAND2_X1 U11169 ( .A1(n14013), .A2(n14607), .ZN(n9622) );
  AND2_X1 U11170 ( .A1(n10013), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9623) );
  AOI21_X1 U11171 ( .B1(n15995), .B2(n15997), .A(n15996), .ZN(n14988) );
  OAI21_X2 U11172 ( .B1(n9762), .B2(n9766), .A(n12472), .ZN(n12971) );
  OR2_X1 U11173 ( .A1(n15024), .A2(n9617), .ZN(n16000) );
  NOR2_X1 U11174 ( .A1(n15024), .A2(n9616), .ZN(n14969) );
  OAI21_X1 U11175 ( .B1(n16060), .B2(n9765), .A(n9763), .ZN(n15024) );
  NAND2_X1 U11176 ( .A1(n14470), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14014) );
  NOR2_X1 U11177 ( .A1(n12099), .A2(n12098), .ZN(n12100) );
  NAND2_X1 U11178 ( .A1(n14820), .A2(n14819), .ZN(n14818) );
  NAND2_X1 U11179 ( .A1(n14285), .A2(n10028), .ZN(n14263) );
  AOI21_X1 U11180 ( .B1(n9915), .B2(n16104), .A(n9913), .ZN(n9912) );
  NAND2_X1 U11181 ( .A1(n11664), .A2(n11663), .ZN(n14289) );
  NAND2_X1 U11182 ( .A1(n9632), .A2(n9631), .ZN(n14470) );
  NAND2_X1 U11183 ( .A1(n9633), .A2(n15758), .ZN(n14490) );
  OR2_X1 U11184 ( .A1(n12096), .A2(n14026), .ZN(n15930) );
  NAND2_X1 U11185 ( .A1(n9783), .A2(n9782), .ZN(n9633) );
  XNOR2_X1 U11186 ( .A(n9693), .B(n10411), .ZN(n14792) );
  OAI21_X1 U11187 ( .B1(n12096), .B2(n12097), .A(n9693), .ZN(n15087) );
  NAND2_X1 U11188 ( .A1(n9819), .A2(n9621), .ZN(n14996) );
  NOR2_X1 U11189 ( .A1(n9615), .A2(n9614), .ZN(n9613) );
  AND2_X1 U11190 ( .A1(n11127), .A2(n9802), .ZN(n10939) );
  INV_X1 U11191 ( .A(n12466), .ZN(n9615) );
  NOR2_X1 U11192 ( .A1(n14812), .A2(n9991), .ZN(n12096) );
  NAND2_X1 U11193 ( .A1(n15377), .A2(n15376), .ZN(n15375) );
  AOI21_X1 U11194 ( .B1(n9766), .B2(n12472), .A(n9764), .ZN(n9763) );
  NAND2_X1 U11195 ( .A1(n9761), .A2(n12460), .ZN(n12465) );
  NAND3_X1 U11196 ( .A1(n9950), .A2(n9948), .A3(n9947), .ZN(n12775) );
  OR2_X1 U11197 ( .A1(n9657), .A2(n9953), .ZN(n9950) );
  INV_X1 U11198 ( .A(n9602), .ZN(n9601) );
  XNOR2_X1 U11199 ( .A(n12470), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16061) );
  INV_X1 U11200 ( .A(n14881), .ZN(n15105) );
  AND2_X1 U11201 ( .A1(n15070), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9614) );
  INV_X1 U11202 ( .A(n15758), .ZN(n9634) );
  NOR2_X1 U11203 ( .A1(n15070), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9612) );
  AND2_X1 U11204 ( .A1(n9778), .A2(n9636), .ZN(n9635) );
  NAND2_X1 U11205 ( .A1(n9594), .A2(n9711), .ZN(n14881) );
  OAI21_X1 U11206 ( .B1(n13995), .B2(n13997), .A(n14936), .ZN(n9602) );
  NAND2_X1 U11207 ( .A1(n10937), .A2(n10936), .ZN(n17291) );
  INV_X1 U11208 ( .A(n12469), .ZN(n12471) );
  AND2_X1 U11209 ( .A1(n9853), .A2(n15822), .ZN(n9852) );
  OR2_X1 U11210 ( .A1(n14761), .A2(n14751), .ZN(n14749) );
  OAI21_X1 U11211 ( .B1(n12459), .B2(n14000), .A(n18845), .ZN(n12303) );
  OR2_X1 U11212 ( .A1(n14890), .A2(n9928), .ZN(n9594) );
  NAND2_X1 U11213 ( .A1(n11997), .A2(n9637), .ZN(n9636) );
  OR2_X1 U11214 ( .A1(n12459), .A2(n15398), .ZN(n12460) );
  XNOR2_X1 U11215 ( .A(n12467), .B(n12461), .ZN(n12464) );
  AOI21_X1 U11216 ( .B1(n11981), .B2(n9775), .A(n9715), .ZN(n9774) );
  NAND2_X1 U11217 ( .A1(n12300), .A2(n12467), .ZN(n12459) );
  INV_X1 U11218 ( .A(n15793), .ZN(n9637) );
  NOR2_X1 U11219 ( .A1(n9702), .A2(n9779), .ZN(n9778) );
  OR2_X1 U11220 ( .A1(n13012), .A2(n13013), .ZN(n9711) );
  NAND2_X1 U11221 ( .A1(n14505), .A2(n12003), .ZN(n14497) );
  NOR2_X1 U11222 ( .A1(n13012), .A2(n9926), .ZN(n14867) );
  INV_X1 U11223 ( .A(n11997), .ZN(n9638) );
  AND2_X1 U11224 ( .A1(n10058), .A2(n10092), .ZN(n9611) );
  AND2_X1 U11225 ( .A1(n14498), .A2(n14496), .ZN(n15758) );
  NAND2_X1 U11226 ( .A1(n14889), .A2(n14888), .ZN(n13012) );
  NAND2_X1 U11227 ( .A1(n9607), .A2(n9609), .ZN(n12467) );
  AND2_X1 U11228 ( .A1(n15768), .A2(n15772), .ZN(n14498) );
  AND2_X1 U11229 ( .A1(n14518), .A2(n12010), .ZN(n14496) );
  AND2_X1 U11230 ( .A1(n12299), .A2(n12277), .ZN(n9607) );
  NAND2_X1 U11231 ( .A1(n19498), .A2(n19684), .ZN(n19424) );
  AND2_X1 U11232 ( .A1(n12323), .A2(n12322), .ZN(n12461) );
  OAI21_X1 U11233 ( .B1(n13573), .B2(n13574), .A(n12453), .ZN(n12456) );
  AND2_X1 U11234 ( .A1(n12298), .A2(n12297), .ZN(n12299) );
  XNOR2_X1 U11235 ( .A(n11993), .B(n11529), .ZN(n11982) );
  OR2_X1 U11236 ( .A1(n12320), .A2(n12319), .ZN(n12323) );
  NOR2_X1 U11237 ( .A1(n17329), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17328) );
  NOR2_X1 U11238 ( .A1(n17429), .A2(n17540), .ZN(n17372) );
  AND2_X1 U11239 ( .A1(n14762), .A2(n14763), .ZN(n14764) );
  AND2_X1 U11240 ( .A1(n14785), .A2(n14786), .ZN(n14762) );
  AOI21_X1 U11241 ( .B1(n11964), .B2(n11625), .A(n11498), .ZN(n13765) );
  OAI21_X1 U11242 ( .B1(n12244), .B2(n12243), .A(n12242), .ZN(n12274) );
  OAI21_X1 U11243 ( .B1(n12258), .B2(n12257), .A(n12256), .ZN(n12273) );
  INV_X1 U11244 ( .A(n17504), .ZN(n17476) );
  XNOR2_X1 U11245 ( .A(n11503), .B(n11501), .ZN(n11964) );
  AND2_X1 U11246 ( .A1(n15198), .A2(n14927), .ZN(n14785) );
  AND2_X1 U11247 ( .A1(n12980), .A2(n9739), .ZN(n15198) );
  OR2_X1 U11248 ( .A1(n12617), .A2(n9945), .ZN(n9942) );
  AND2_X1 U11249 ( .A1(n9704), .A2(n12236), .ZN(n12305) );
  AND2_X1 U11250 ( .A1(n12237), .A2(n12236), .ZN(n19313) );
  INV_X1 U11251 ( .A(n12232), .ZN(n12234) );
  INV_X1 U11252 ( .A(n11438), .ZN(n9591) );
  AND2_X1 U11253 ( .A1(n12237), .A2(n12232), .ZN(n19368) );
  AND2_X1 U11254 ( .A1(n10786), .A2(n10003), .ZN(n15953) );
  NAND2_X2 U11255 ( .A1(n19858), .A2(n11267), .ZN(n14322) );
  AND2_X1 U11256 ( .A1(n9704), .A2(n12233), .ZN(n12311) );
  NAND2_X1 U11257 ( .A1(n12589), .A2(n12588), .ZN(n12614) );
  NAND2_X1 U11258 ( .A1(n12208), .A2(n16115), .ZN(n12227) );
  AND2_X1 U11259 ( .A1(n12237), .A2(n12218), .ZN(n19343) );
  OR2_X1 U11260 ( .A1(n18872), .A2(n12601), .ZN(n12229) );
  AND2_X1 U11261 ( .A1(n18872), .A2(n13238), .ZN(n12232) );
  NOR2_X1 U11262 ( .A1(n15289), .A2(n10694), .ZN(n15270) );
  AND2_X1 U11263 ( .A1(n9817), .A2(n12350), .ZN(n9621) );
  NOR2_X1 U11264 ( .A1(n14636), .A2(n14635), .ZN(n14638) );
  AND2_X1 U11265 ( .A1(n10923), .A2(n9808), .ZN(n17478) );
  NAND2_X1 U11266 ( .A1(n9642), .A2(n9641), .ZN(n9644) );
  OR2_X1 U11267 ( .A1(n16115), .A2(n13332), .ZN(n12235) );
  NAND2_X1 U11268 ( .A1(n15313), .A2(n15314), .ZN(n15289) );
  AOI21_X1 U11269 ( .B1(n13394), .B2(n13393), .A(n19756), .ZN(n13418) );
  NAND2_X1 U11270 ( .A1(n9658), .A2(n12211), .ZN(n18872) );
  NAND2_X1 U11271 ( .A1(n12384), .A2(n14848), .ZN(n12399) );
  NAND2_X1 U11272 ( .A1(n12597), .A2(n12596), .ZN(n12611) );
  AND2_X1 U11273 ( .A1(n10021), .A2(n11318), .ZN(n11934) );
  AND2_X1 U11274 ( .A1(n15361), .A2(n9917), .ZN(n15313) );
  NAND2_X1 U11275 ( .A1(n10603), .A2(n10602), .ZN(n15361) );
  CLKBUF_X2 U11276 ( .A(n12593), .Z(n16115) );
  NOR2_X1 U11277 ( .A1(n12374), .A2(n10785), .ZN(n12364) );
  NAND4_X1 U11278 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(n16922), .A4(n13950), .ZN(n15535) );
  NAND2_X1 U11279 ( .A1(n9809), .A2(n12207), .ZN(n9995) );
  NOR2_X2 U11280 ( .A1(n17564), .A2(n10922), .ZN(n10924) );
  NOR2_X2 U11281 ( .A1(n19033), .A2(n19338), .ZN(n19034) );
  NAND2_X1 U11282 ( .A1(n12604), .A2(n12603), .ZN(n12605) );
  NAND2_X1 U11283 ( .A1(n11371), .A2(n11369), .ZN(n11367) );
  NAND2_X1 U11284 ( .A1(n12381), .A2(n9996), .ZN(n12374) );
  NAND2_X1 U11285 ( .A1(n15393), .A2(n10583), .ZN(n15387) );
  NOR2_X2 U11286 ( .A1(n9692), .A2(n12378), .ZN(n12381) );
  INV_X2 U11287 ( .A(n13752), .ZN(n18865) );
  OR2_X1 U11288 ( .A1(n9987), .A2(n9989), .ZN(n9986) );
  AND2_X2 U11289 ( .A1(n10306), .A2(n10305), .ZN(n12207) );
  NAND2_X1 U11290 ( .A1(n9603), .A2(n10297), .ZN(n9809) );
  AOI21_X1 U11291 ( .B1(n10917), .B2(n17580), .A(n11098), .ZN(n11101) );
  NAND2_X1 U11292 ( .A1(n12214), .A2(n10283), .ZN(n9603) );
  XNOR2_X1 U11293 ( .A(n11287), .B(n11360), .ZN(n11305) );
  NAND2_X1 U11294 ( .A1(n9605), .A2(n9604), .ZN(n10306) );
  OR2_X1 U11295 ( .A1(n12213), .A2(n12212), .ZN(n12216) );
  NAND2_X1 U11296 ( .A1(n11419), .A2(n11418), .ZN(n20153) );
  NOR2_X1 U11297 ( .A1(n10517), .A2(n9910), .ZN(n9909) );
  OR2_X1 U11298 ( .A1(n13277), .A2(n13276), .ZN(n9906) );
  NAND2_X1 U11299 ( .A1(n9640), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9639) );
  NAND3_X1 U11300 ( .A1(n10307), .A2(n10288), .A3(n10287), .ZN(n12213) );
  NOR2_X1 U11301 ( .A1(n19735), .A2(n10793), .ZN(n18876) );
  INV_X2 U11302 ( .A(n16998), .ZN(n16980) );
  NOR2_X1 U11303 ( .A1(n10499), .A2(n10498), .ZN(n10516) );
  AND2_X1 U11304 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n16984), .ZN(n16979) );
  NAND2_X1 U11305 ( .A1(n11360), .A2(n11284), .ZN(n9659) );
  NOR2_X1 U11306 ( .A1(n17602), .A2(n17601), .ZN(n17600) );
  NAND2_X1 U11307 ( .A1(n12336), .A2(n10234), .ZN(n12405) );
  AND4_X1 U11308 ( .A1(n10286), .A2(n10285), .A3(n16171), .A4(n10284), .ZN(
        n10287) );
  OAI21_X1 U11309 ( .B1(n11042), .B2(n13947), .A(n18420), .ZN(n11049) );
  NOR2_X1 U11310 ( .A1(n13391), .A2(n9630), .ZN(n13444) );
  NAND3_X1 U11311 ( .A1(n13413), .A2(n13415), .A3(n11273), .ZN(n11274) );
  INV_X1 U11312 ( .A(n10325), .ZN(n10406) );
  AND2_X1 U11313 ( .A1(n13212), .A2(n13211), .ZN(n13214) );
  NAND2_X1 U11314 ( .A1(n11280), .A2(n13389), .ZN(n11302) );
  AND2_X1 U11315 ( .A1(n12161), .A2(n12158), .ZN(n13413) );
  INV_X2 U11316 ( .A(n10405), .ZN(n10394) );
  NAND2_X1 U11317 ( .A1(n13245), .A2(n11272), .ZN(n11273) );
  INV_X1 U11318 ( .A(n9620), .ZN(n12560) );
  OAI21_X1 U11319 ( .B1(n13112), .B2(n10473), .A(n10472), .ZN(n13212) );
  NAND2_X1 U11320 ( .A1(n9628), .A2(n9626), .ZN(n13194) );
  NAND2_X1 U11321 ( .A1(n9628), .A2(n9627), .ZN(n12161) );
  NOR2_X1 U11322 ( .A1(n17622), .A2(n17621), .ZN(n17620) );
  AND2_X2 U11323 ( .A1(n10290), .A2(n12939), .ZN(n10291) );
  NOR2_X1 U11324 ( .A1(n13395), .A2(n11930), .ZN(n9627) );
  NAND2_X1 U11325 ( .A1(n10260), .A2(n12523), .ZN(n12545) );
  AND2_X1 U11326 ( .A1(n12260), .A2(n12259), .ZN(n12270) );
  INV_X1 U11327 ( .A(n11277), .ZN(n9628) );
  AND4_X1 U11328 ( .A1(n11299), .A2(n11298), .A3(n13403), .A4(n11297), .ZN(
        n11300) );
  INV_X1 U11329 ( .A(n12034), .ZN(n12052) );
  INV_X1 U11330 ( .A(n13395), .ZN(n9626) );
  NOR2_X1 U11331 ( .A1(n17133), .A2(n10916), .ZN(n10918) );
  NOR2_X1 U11332 ( .A1(n13425), .A2(n13379), .ZN(n13409) );
  NOR2_X1 U11333 ( .A1(n11271), .A2(n11270), .ZN(n13245) );
  NOR2_X1 U11334 ( .A1(n12266), .A2(n12265), .ZN(n12260) );
  NAND2_X1 U11335 ( .A1(n11421), .A2(n11420), .ZN(n12034) );
  NAND2_X1 U11336 ( .A1(n13270), .A2(n13269), .ZN(n9855) );
  NAND2_X1 U11337 ( .A1(n13189), .A2(n11270), .ZN(n13395) );
  OR2_X1 U11338 ( .A1(n11950), .A2(n11421), .ZN(n9641) );
  NAND3_X1 U11339 ( .A1(n9810), .A2(n9706), .A3(n13111), .ZN(n10278) );
  OR2_X1 U11340 ( .A1(n11421), .A2(n11994), .ZN(n11991) );
  NAND2_X1 U11341 ( .A1(n12437), .A2(n9596), .ZN(n12563) );
  OR2_X2 U11342 ( .A1(n10433), .A2(n10478), .ZN(n10755) );
  NOR2_X1 U11343 ( .A1(n10235), .A2(n10234), .ZN(n10236) );
  MUX2_X1 U11344 ( .A(n12427), .B(P2_EBX_REG_2__SCAN_IN), .S(n10768), .Z(
        n12266) );
  OR2_X1 U11345 ( .A1(n12443), .A2(n13720), .ZN(n13112) );
  NAND2_X1 U11346 ( .A1(n13416), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11421) );
  NOR2_X1 U11347 ( .A1(n11266), .A2(n11936), .ZN(n13191) );
  INV_X1 U11348 ( .A(n18003), .ZN(n11039) );
  INV_X1 U11349 ( .A(n11295), .ZN(n15572) );
  AND2_X1 U11350 ( .A1(n11281), .A2(n11267), .ZN(n11294) );
  AND2_X1 U11351 ( .A1(n10230), .A2(n10233), .ZN(n10266) );
  CLKBUF_X1 U11352 ( .A(n11289), .Z(n13593) );
  NAND2_X1 U11353 ( .A1(n13266), .A2(n14089), .ZN(n14107) );
  AND2_X2 U11354 ( .A1(n10601), .A2(n10600), .ZN(n14002) );
  INV_X1 U11355 ( .A(n17006), .ZN(n18009) );
  CLKBUF_X1 U11356 ( .A(n10258), .Z(n10259) );
  NAND2_X1 U11357 ( .A1(n10865), .A2(n10864), .ZN(n17150) );
  AND2_X2 U11358 ( .A1(n9597), .A2(n19732), .ZN(n9595) );
  INV_X1 U11359 ( .A(n11265), .ZN(n11235) );
  INV_X1 U11360 ( .A(n10255), .ZN(n10767) );
  AND2_X1 U11361 ( .A1(n12515), .A2(n9597), .ZN(n9596) );
  OR2_X1 U11362 ( .A1(n10494), .A2(n10493), .ZN(n12442) );
  OR2_X1 U11364 ( .A1(n10511), .A2(n10510), .ZN(n10765) );
  NAND2_X1 U11365 ( .A1(n10192), .A2(n10191), .ZN(n19045) );
  NAND2_X1 U11366 ( .A1(n10098), .A2(n11193), .ZN(n11265) );
  AND2_X1 U11367 ( .A1(n11293), .A2(n20032), .ZN(n11290) );
  NAND2_X2 U11368 ( .A1(n10057), .A2(n10056), .ZN(n12515) );
  NAND2_X1 U11369 ( .A1(n10168), .A2(n10167), .ZN(n10256) );
  NAND2_X1 U11370 ( .A1(n10144), .A2(n10143), .ZN(n10258) );
  NAND2_X1 U11371 ( .A1(n10088), .A2(n10087), .ZN(n10215) );
  NAND2_X1 U11372 ( .A1(n9705), .A2(n10073), .ZN(n10057) );
  NAND3_X2 U11373 ( .A1(n11252), .A2(n11251), .A3(n10095), .ZN(n20005) );
  NAND4_X2 U11374 ( .A1(n11183), .A2(n11181), .A3(n11182), .A4(n11180), .ZN(
        n20032) );
  AND4_X1 U11375 ( .A1(n11192), .A2(n11191), .A3(n11190), .A4(n11189), .ZN(
        n11193) );
  AND4_X1 U11376 ( .A1(n11244), .A2(n11243), .A3(n11242), .A4(n11241), .ZN(
        n11252) );
  AND4_X1 U11377 ( .A1(n11162), .A2(n11161), .A3(n11160), .A4(n11159), .ZN(
        n9699) );
  AND4_X1 U11378 ( .A1(n11152), .A2(n11151), .A3(n11150), .A4(n11149), .ZN(
        n11163) );
  AND4_X1 U11379 ( .A1(n11179), .A2(n11178), .A3(n11177), .A4(n11176), .ZN(
        n11180) );
  AND4_X1 U11380 ( .A1(n11171), .A2(n11170), .A3(n11169), .A4(n11168), .ZN(
        n11182) );
  AND4_X1 U11381 ( .A1(n11175), .A2(n11174), .A3(n11173), .A4(n11172), .ZN(
        n11181) );
  AND4_X1 U11382 ( .A1(n11167), .A2(n11166), .A3(n11165), .A4(n11164), .ZN(
        n11183) );
  AND2_X2 U11383 ( .A1(n10223), .A2(n10136), .ZN(n12747) );
  AND3_X1 U11384 ( .A1(n10209), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10208), .ZN(n10210) );
  INV_X2 U11385 ( .A(n10944), .ZN(n16953) );
  INV_X2 U11386 ( .A(n9665), .ZN(n12135) );
  INV_X2 U11387 ( .A(n16307), .ZN(U215) );
  NOR2_X2 U11388 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n9656), .ZN(
        n11453) );
  BUF_X4 U11389 ( .A(n10890), .Z(n16951) );
  NAND2_X1 U11390 ( .A1(n9790), .A2(n9789), .ZN(n10962) );
  BUF_X2 U11391 ( .A(n11253), .Z(n12112) );
  INV_X2 U11392 ( .A(n9666), .ZN(n9667) );
  BUF_X2 U11393 ( .A(n11194), .Z(n12129) );
  OR2_X1 U11394 ( .A1(n10044), .A2(n9617), .ZN(n9616) );
  CLKBUF_X3 U11395 ( .A(n11194), .Z(n12106) );
  OR2_X1 U11396 ( .A1(n16692), .A2(n10807), .ZN(n9695) );
  NOR2_X1 U11397 ( .A1(n10811), .A2(n10810), .ZN(n10853) );
  OR2_X1 U11398 ( .A1(n10811), .A2(n16693), .ZN(n10090) );
  INV_X1 U11399 ( .A(n10447), .ZN(n12777) );
  INV_X2 U11400 ( .A(n16309), .ZN(n16311) );
  INV_X4 U11401 ( .A(n9694), .ZN(n16945) );
  OR2_X1 U11402 ( .A1(n13978), .A2(n10808), .ZN(n13977) );
  AND2_X2 U11403 ( .A1(n10435), .A2(n10299), .ZN(n10226) );
  CLKBUF_X3 U11404 ( .A(n11240), .Z(n12136) );
  AND2_X2 U11405 ( .A1(n12892), .A2(n10136), .ZN(n10522) );
  AND2_X4 U11406 ( .A1(n11155), .A2(n13430), .ZN(n11200) );
  AND2_X1 U11407 ( .A1(n11155), .A2(n13456), .ZN(n11253) );
  AND2_X1 U11408 ( .A1(n9781), .A2(n13637), .ZN(n11194) );
  OR2_X1 U11409 ( .A1(n10811), .A2(n16692), .ZN(n10809) );
  NOR2_X1 U11410 ( .A1(n9619), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15425) );
  AND2_X1 U11411 ( .A1(n9599), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10129) );
  AND3_X1 U11412 ( .A1(n12014), .A2(n12013), .A3(n14603), .ZN(n9758) );
  AND2_X2 U11413 ( .A1(n13637), .A2(n13430), .ZN(n11458) );
  NOR2_X1 U11414 ( .A1(n9645), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11156) );
  NAND2_X1 U11415 ( .A1(n10436), .A2(n10299), .ZN(n10447) );
  NOR2_X1 U11416 ( .A1(n19681), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12755) );
  NAND2_X1 U11417 ( .A1(n13456), .A2(n13638), .ZN(n11310) );
  AND2_X2 U11418 ( .A1(n13456), .A2(n13637), .ZN(n11336) );
  NOR2_X1 U11419 ( .A1(n15547), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11158) );
  AND2_X1 U11420 ( .A1(n13431), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11155) );
  AND2_X1 U11421 ( .A1(n13433), .A2(n11154), .ZN(n11240) );
  AND2_X2 U11422 ( .A1(n13456), .A2(n13637), .ZN(n9673) );
  NAND2_X1 U11423 ( .A1(n18604), .A2(n18612), .ZN(n16692) );
  AND2_X2 U11425 ( .A1(n15435), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12892) );
  NAND2_X2 U11426 ( .A1(n11052), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9791) );
  OR2_X1 U11427 ( .A1(n16693), .A2(n13978), .ZN(n9694) );
  NAND2_X1 U11428 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16693) );
  AND2_X1 U11429 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15435) );
  INV_X1 U11430 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15415) );
  INV_X1 U11431 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9599) );
  INV_X1 U11432 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9619) );
  INV_X1 U11433 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9598) );
  AND2_X1 U11434 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11154) );
  AND2_X1 U11435 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13638) );
  NOR2_X1 U11436 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11148) );
  INV_X1 U11437 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18457) );
  INV_X1 U11438 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11153) );
  NOR2_X2 U11439 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13637) );
  INV_X1 U11440 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9645) );
  INV_X2 U11441 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15547) );
  INV_X1 U11442 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10048) );
  NOR2_X2 U11443 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13456) );
  INV_X4 U11444 ( .A(n9597), .ZN(n10264) );
  NOR2_X1 U11445 ( .A1(n19742), .A2(n9597), .ZN(n13137) );
  NAND2_X2 U11446 ( .A1(n10205), .A2(n10204), .ZN(n9597) );
  INV_X1 U11447 ( .A(n9906), .ZN(n13278) );
  NAND3_X1 U11448 ( .A1(n9906), .A2(n9908), .A3(n9909), .ZN(n15393) );
  AND2_X2 U11449 ( .A1(n9598), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10435) );
  NOR2_X1 U11450 ( .A1(n19741), .A2(n9599), .ZN(n9933) );
  INV_X1 U11451 ( .A(n10303), .ZN(n9604) );
  INV_X1 U11452 ( .A(n10304), .ZN(n9605) );
  INV_X1 U11453 ( .A(n12455), .ZN(n9609) );
  OAI21_X1 U11454 ( .B1(n12455), .B2(n12454), .A(n9610), .ZN(n12300) );
  INV_X1 U11457 ( .A(n12299), .ZN(n9610) );
  NAND2_X1 U11458 ( .A1(n10060), .A2(n9611), .ZN(n13992) );
  AOI21_X2 U11459 ( .B1(n15379), .B2(n9613), .A(n9612), .ZN(n16060) );
  NAND2_X1 U11460 ( .A1(n15380), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15379) );
  INV_X1 U11461 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n9617) );
  NAND2_X1 U11462 ( .A1(n13829), .A2(n12458), .ZN(n13914) );
  NAND3_X1 U11463 ( .A1(n13829), .A2(n9618), .A3(n12458), .ZN(n9761) );
  INV_X1 U11464 ( .A(n13915), .ZN(n9618) );
  NAND3_X1 U11465 ( .A1(n10218), .A2(n10217), .A3(n12540), .ZN(n12551) );
  NAND4_X1 U11466 ( .A1(n10218), .A2(n10217), .A3(n12540), .A4(n12521), .ZN(
        n9620) );
  NAND2_X2 U11467 ( .A1(n15375), .A2(n9682), .ZN(n9819) );
  INV_X1 U11468 ( .A(n12456), .ZN(n9654) );
  NAND2_X1 U11469 ( .A1(n9585), .A2(n14014), .ZN(n14406) );
  NAND2_X2 U11470 ( .A1(n14014), .A2(n14469), .ZN(n14013) );
  NAND2_X1 U11471 ( .A1(n14014), .A2(n14479), .ZN(n10013) );
  NAND3_X1 U11472 ( .A1(n9625), .A2(n11963), .A3(n9624), .ZN(n15807) );
  NAND2_X1 U11473 ( .A1(n10015), .A2(n19926), .ZN(n9624) );
  INV_X1 U11474 ( .A(n9777), .ZN(n10015) );
  NAND3_X1 U11475 ( .A1(n10014), .A2(n19926), .A3(n13526), .ZN(n9625) );
  NAND2_X1 U11476 ( .A1(n9777), .A2(n10016), .ZN(n10014) );
  NAND2_X1 U11477 ( .A1(n15807), .A2(n15806), .ZN(n15805) );
  NOR2_X1 U11478 ( .A1(n13194), .A2(n9592), .ZN(n13987) );
  NOR2_X1 U11479 ( .A1(n9629), .A2(n13194), .ZN(n13179) );
  INV_X1 U11480 ( .A(n13377), .ZN(n9629) );
  INV_X1 U11481 ( .A(n13194), .ZN(n9630) );
  NAND3_X1 U11482 ( .A1(n9783), .A2(n9782), .A3(n9681), .ZN(n9632) );
  OAI21_X2 U11483 ( .B1(n9850), .B2(n9638), .A(n9635), .ZN(n14527) );
  NAND2_X1 U11484 ( .A1(n13878), .A2(n11997), .ZN(n9780) );
  NAND2_X1 U11485 ( .A1(n9850), .A2(n15793), .ZN(n13878) );
  NAND3_X1 U11486 ( .A1(n12007), .A2(n12000), .A3(n14527), .ZN(n12008) );
  INV_X1 U11487 ( .A(n11284), .ZN(n9640) );
  NAND2_X2 U11488 ( .A1(n11274), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11360) );
  NAND3_X1 U11489 ( .A1(n11416), .A2(n11372), .A3(n20578), .ZN(n9642) );
  NAND2_X2 U11491 ( .A1(n11390), .A2(n11391), .ZN(n11439) );
  XNOR2_X2 U11492 ( .A(n9644), .B(n11389), .ZN(n11390) );
  NOR2_X1 U11493 ( .A1(n13914), .A2(n13915), .ZN(n9646) );
  AND2_X1 U11494 ( .A1(n19742), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13111) );
  NAND2_X4 U11495 ( .A1(n11993), .A2(n11992), .ZN(n15785) );
  INV_X2 U11496 ( .A(n11271), .ZN(n13378) );
  AND2_X1 U11497 ( .A1(n9932), .A2(n10280), .ZN(n9647) );
  XNOR2_X1 U11498 ( .A(n12456), .B(n12457), .ZN(n13827) );
  NOR2_X2 U11499 ( .A1(n10924), .A2(n17881), .ZN(n17845) );
  OAI211_X1 U11500 ( .C1(n10394), .C2(n10772), .A(n10313), .B(n10312), .ZN(
        n10314) );
  CLKBUF_X1 U11501 ( .A(n15796), .Z(n9648) );
  OAI211_X1 U11502 ( .C1(n13526), .C2(n10015), .A(n19926), .B(n10014), .ZN(
        n9649) );
  NAND2_X1 U11503 ( .A1(n9788), .A2(n9787), .ZN(n11503) );
  NAND2_X1 U11504 ( .A1(n14438), .A2(n14428), .ZN(n9652) );
  AND2_X2 U11505 ( .A1(n11157), .A2(n13430), .ZN(n9670) );
  CLKBUF_X1 U11506 ( .A(n11311), .Z(n11757) );
  NAND2_X1 U11507 ( .A1(n15379), .A2(n12466), .ZN(n9653) );
  NAND2_X1 U11508 ( .A1(n12496), .A2(n10766), .ZN(n12540) );
  NAND2_X1 U11509 ( .A1(n12276), .A2(n12275), .ZN(n12455) );
  AND2_X1 U11510 ( .A1(n10256), .A2(n10239), .ZN(n10233) );
  CLKBUF_X1 U11511 ( .A(n15805), .Z(n9655) );
  NAND2_X1 U11512 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n11156), .ZN(
        n9656) );
  NAND2_X2 U11513 ( .A1(n13359), .A2(n12620), .ZN(n13701) );
  NAND2_X2 U11514 ( .A1(n9940), .A2(n9939), .ZN(n13359) );
  OR2_X1 U11515 ( .A1(n16000), .A2(n10045), .ZN(n14976) );
  AND2_X2 U11516 ( .A1(n14846), .A2(n14847), .ZN(n9657) );
  INV_X1 U11517 ( .A(n9657), .ZN(n14841) );
  NAND2_X1 U11518 ( .A1(n12209), .A2(n12214), .ZN(n9658) );
  AOI21_X2 U11519 ( .B1(n11048), .B2(n13964), .A(n11047), .ZN(n18432) );
  NOR2_X2 U11520 ( .A1(n17991), .A2(n17781), .ZN(n17789) );
  NAND2_X1 U11521 ( .A1(n11109), .A2(n17547), .ZN(n17843) );
  NOR2_X2 U11522 ( .A1(n17647), .A2(n16208), .ZN(n17552) );
  NAND2_X1 U11523 ( .A1(n9936), .A2(n9934), .ZN(n12890) );
  OR2_X1 U11524 ( .A1(n12580), .A2(n16073), .ZN(n12486) );
  OR2_X1 U11525 ( .A1(n12467), .A2(n12468), .ZN(n12469) );
  INV_X1 U11526 ( .A(n14290), .ZN(n9660) );
  NOR2_X4 U11527 ( .A1(n14215), .A2(n9661), .ZN(n14285) );
  NAND2_X1 U11528 ( .A1(n11663), .A2(n9660), .ZN(n9661) );
  INV_X1 U11529 ( .A(n10028), .ZN(n9662) );
  AND2_X2 U11530 ( .A1(n9663), .A2(n14285), .ZN(n14256) );
  NOR2_X1 U11531 ( .A1(n14264), .A2(n9662), .ZN(n9663) );
  NOR2_X2 U11532 ( .A1(n17169), .A2(n17024), .ZN(n17016) );
  NOR3_X2 U11533 ( .A1(n17181), .A2(n17083), .A3(n17048), .ZN(n17044) );
  NAND2_X1 U11534 ( .A1(n9995), .A2(n10306), .ZN(n10315) );
  OAI21_X1 U11535 ( .B1(n13656), .B2(n12022), .A(n11933), .ZN(n13354) );
  NAND2_X2 U11536 ( .A1(n10268), .A2(n10255), .ZN(n10263) );
  NAND2_X2 U11537 ( .A1(n11367), .A2(n11366), .ZN(n11416) );
  OR2_X2 U11538 ( .A1(n15305), .A2(n15254), .ZN(n15269) );
  AOI21_X1 U11539 ( .B1(n9659), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11361), .ZN(n11370) );
  OR2_X1 U11540 ( .A1(n11360), .A2(n11359), .ZN(n11369) );
  OAI21_X2 U11541 ( .B1(n14988), .B2(n14989), .A(n12404), .ZN(n14978) );
  NAND2_X1 U11542 ( .A1(n13356), .A2(n11949), .ZN(n11956) );
  AND2_X2 U11543 ( .A1(n13785), .A2(n13927), .ZN(n13868) );
  NOR2_X2 U11544 ( .A1(n13701), .A2(n12621), .ZN(n13785) );
  NOR2_X1 U11545 ( .A1(n14019), .A2(n14419), .ZN(n14408) );
  XNOR2_X2 U11546 ( .A(n10318), .B(n10316), .ZN(n12206) );
  OAI21_X2 U11547 ( .B1(n18433), .B2(n11049), .A(n18432), .ZN(n18438) );
  NOR2_X1 U11548 ( .A1(n11153), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9781) );
  AND2_X1 U11549 ( .A1(n11265), .A2(n11267), .ZN(n11206) );
  XNOR2_X1 U11550 ( .A(n11416), .B(n20153), .ZN(n13633) );
  XNOR2_X2 U11551 ( .A(n10315), .B(n12206), .ZN(n13332) );
  OAI21_X2 U11552 ( .B1(n14418), .B2(n9725), .A(n10009), .ZN(n10012) );
  AND2_X2 U11553 ( .A1(n13892), .A2(n10029), .ZN(n14214) );
  AND2_X1 U11554 ( .A1(n11157), .A2(n13430), .ZN(n9669) );
  AND2_X1 U11555 ( .A1(n11157), .A2(n13430), .ZN(n11320) );
  AND2_X1 U11556 ( .A1(n13432), .A2(n11148), .ZN(n9671) );
  AND4_X4 U11557 ( .A1(n15547), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A4(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11258) );
  AND2_X1 U11558 ( .A1(n10291), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9674) );
  AND2_X1 U11559 ( .A1(n10291), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9675) );
  AND2_X4 U11560 ( .A1(n10291), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10405) );
  AND2_X2 U11561 ( .A1(n12901), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10527) );
  NAND2_X1 U11562 ( .A1(n13330), .A2(n13331), .ZN(n9946) );
  NOR2_X1 U11563 ( .A1(n16138), .A2(n10264), .ZN(n13131) );
  OAI21_X1 U11564 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n11052), .A(
        n11055), .ZN(n11056) );
  OR2_X1 U11565 ( .A1(n11054), .A2(n11053), .ZN(n11055) );
  OR2_X1 U11566 ( .A1(n11421), .A2(n11986), .ZN(n11353) );
  AND2_X1 U11567 ( .A1(n12755), .A2(n10436), .ZN(n12748) );
  INV_X1 U11568 ( .A(n10269), .ZN(n9810) );
  NOR2_X1 U11569 ( .A1(n16368), .A2(n9884), .ZN(n9883) );
  NAND2_X1 U11570 ( .A1(n18000), .A2(n17092), .ZN(n11045) );
  NAND2_X1 U11571 ( .A1(n10043), .A2(n11926), .ZN(n10042) );
  INV_X1 U11572 ( .A(n14176), .ZN(n10043) );
  NAND2_X1 U11573 ( .A1(n9590), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9853) );
  INV_X1 U11574 ( .A(n11447), .ZN(n11711) );
  INV_X1 U11575 ( .A(n11471), .ZN(n12150) );
  NAND2_X1 U11576 ( .A1(n11957), .A2(n13187), .ZN(n11961) );
  AND2_X1 U11577 ( .A1(n11278), .A2(n13401), .ZN(n11301) );
  NAND3_X1 U11578 ( .A1(n11265), .A2(n20005), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12053) );
  NAND2_X1 U11579 ( .A1(n11270), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11420) );
  NOR2_X1 U11580 ( .A1(n9999), .A2(n10782), .ZN(n9998) );
  AND2_X1 U11581 ( .A1(n12336), .A2(n12334), .ZN(n12337) );
  AND2_X1 U11582 ( .A1(n12324), .A2(n10776), .ZN(n12336) );
  NOR2_X1 U11583 ( .A1(n12325), .A2(n12330), .ZN(n10776) );
  NOR2_X1 U11584 ( .A1(n9981), .A2(n9980), .ZN(n9979) );
  INV_X1 U11585 ( .A(n13887), .ZN(n9980) );
  OR2_X1 U11586 ( .A1(n13990), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10092) );
  OAI21_X1 U11587 ( .B1(n10270), .B2(n19057), .A(n10271), .ZN(n10272) );
  AOI21_X1 U11588 ( .B1(n10915), .B2(n9966), .A(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n9962) );
  INV_X1 U11589 ( .A(n11711), .ZN(n12155) );
  NAND2_X1 U11590 ( .A1(n15796), .A2(n15794), .ZN(n9850) );
  XNOR2_X1 U11591 ( .A(n12420), .B(n13998), .ZN(n15922) );
  AND2_X1 U11592 ( .A1(n15953), .A2(n10389), .ZN(n12413) );
  CLKBUF_X1 U11593 ( .A(n10759), .Z(n10760) );
  INV_X1 U11594 ( .A(n12613), .ZN(n9945) );
  NOR2_X1 U11595 ( .A1(n12616), .A2(n12615), .ZN(n13301) );
  AND2_X1 U11596 ( .A1(n14889), .A2(n9924), .ZN(n14869) );
  NOR2_X1 U11597 ( .A1(n9926), .A2(n9925), .ZN(n9924) );
  NAND2_X1 U11598 ( .A1(n14866), .A2(n14888), .ZN(n9925) );
  NAND2_X1 U11599 ( .A1(n14869), .A2(n12081), .ZN(n12085) );
  INV_X1 U11600 ( .A(n13560), .ZN(n9910) );
  NAND2_X1 U11601 ( .A1(n12535), .A2(n19598), .ZN(n12578) );
  AND2_X1 U11602 ( .A1(n19741), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12600) );
  XNOR2_X1 U11603 ( .A(n12605), .B(n12606), .ZN(n13149) );
  OR2_X1 U11604 ( .A1(n12614), .A2(n12591), .ZN(n12592) );
  AND2_X1 U11605 ( .A1(n12510), .A2(n12508), .ZN(n16138) );
  NAND2_X1 U11606 ( .A1(n16402), .A2(n9732), .ZN(n9887) );
  NAND2_X1 U11607 ( .A1(n9732), .A2(n17359), .ZN(n9902) );
  NAND2_X1 U11608 ( .A1(n16450), .A2(n9732), .ZN(n9901) );
  NAND2_X1 U11609 ( .A1(n15539), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11127) );
  NAND2_X1 U11610 ( .A1(n11100), .A2(n10918), .ZN(n16215) );
  NAND2_X1 U11611 ( .A1(n15088), .A2(n16105), .ZN(n9916) );
  INV_X1 U11612 ( .A(n16097), .ZN(n15410) );
  NAND2_X1 U11613 ( .A1(n10291), .A2(n9733), .ZN(n10249) );
  INV_X1 U11614 ( .A(n11478), .ZN(n9849) );
  NAND2_X1 U11615 ( .A1(n12066), .A2(n11235), .ZN(n13389) );
  OR2_X1 U11616 ( .A1(n11330), .A2(n11329), .ZN(n11986) );
  NAND2_X1 U11617 ( .A1(n11232), .A2(n11231), .ZN(n11234) );
  NAND2_X1 U11618 ( .A1(n13383), .A2(n20032), .ZN(n11232) );
  NAND2_X1 U11619 ( .A1(n11293), .A2(n11265), .ZN(n11233) );
  AND2_X1 U11620 ( .A1(n10274), .A2(n12538), .ZN(n10275) );
  NAND2_X1 U11621 ( .A1(n10129), .A2(n15415), .ZN(n10135) );
  INV_X1 U11622 ( .A(n12277), .ZN(n12454) );
  NAND2_X1 U11623 ( .A1(n10289), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10307) );
  NAND2_X1 U11624 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19720), .ZN(
        n12261) );
  NOR2_X1 U11625 ( .A1(n17143), .A2(n10909), .ZN(n10913) );
  NAND2_X1 U11626 ( .A1(n10905), .A2(n17150), .ZN(n10909) );
  NAND2_X1 U11627 ( .A1(n11270), .A2(n9592), .ZN(n11289) );
  AND2_X1 U11628 ( .A1(n10027), .A2(n10026), .ZN(n10025) );
  INV_X1 U11629 ( .A(n14462), .ZN(n10026) );
  AND2_X1 U11630 ( .A1(n14250), .A2(n14257), .ZN(n10027) );
  OR2_X1 U11631 ( .A1(n15785), .A2(n12009), .ZN(n14518) );
  INV_X1 U11632 ( .A(n13893), .ZN(n14307) );
  INV_X1 U11633 ( .A(n14259), .ZN(n9871) );
  AND2_X1 U11634 ( .A1(n9864), .A2(n9717), .ZN(n9863) );
  OR2_X1 U11635 ( .A1(n11342), .A2(n11341), .ZN(n11941) );
  NAND2_X1 U11636 ( .A1(n13188), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11284) );
  INV_X1 U11637 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20407) );
  INV_X1 U11638 ( .A(n20052), .ZN(n20160) );
  NAND2_X1 U11639 ( .A1(n11930), .A2(n20032), .ZN(n12022) );
  NAND2_X1 U11640 ( .A1(n10421), .A2(n10420), .ZN(n12503) );
  NOR2_X1 U11641 ( .A1(n10006), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10005) );
  INV_X1 U11642 ( .A(n10007), .ZN(n10006) );
  NOR2_X1 U11643 ( .A1(n9997), .A2(n12371), .ZN(n9996) );
  INV_X1 U11644 ( .A(n9998), .ZN(n9997) );
  AND2_X1 U11645 ( .A1(n10777), .A2(n12341), .ZN(n10002) );
  NAND2_X1 U11646 ( .A1(n12405), .A2(n10778), .ZN(n12349) );
  INV_X1 U11647 ( .A(n10766), .ZN(n10792) );
  NAND2_X1 U11648 ( .A1(n12825), .A2(n12827), .ZN(n12828) );
  INV_X1 U11649 ( .A(n12748), .ZN(n12713) );
  INV_X1 U11650 ( .A(n14859), .ZN(n9955) );
  AND2_X1 U11651 ( .A1(n12981), .A2(n15231), .ZN(n9923) );
  NOR2_X1 U11652 ( .A1(n9919), .A2(n10621), .ZN(n9918) );
  INV_X1 U11653 ( .A(n15360), .ZN(n9919) );
  NAND2_X1 U11654 ( .A1(n10239), .A2(n10767), .ZN(n10257) );
  AND2_X1 U11655 ( .A1(n10234), .A2(n19732), .ZN(n10469) );
  NOR2_X1 U11656 ( .A1(n12397), .A2(n10050), .ZN(n10049) );
  INV_X1 U11657 ( .A(n10051), .ZN(n10050) );
  NOR2_X1 U11658 ( .A1(n18685), .A2(n9832), .ZN(n9831) );
  INV_X1 U11659 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9832) );
  OR2_X1 U11660 ( .A1(n9844), .A2(n16018), .ZN(n9843) );
  NAND2_X1 U11661 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n9844) );
  NOR2_X1 U11662 ( .A1(n13675), .A2(n9985), .ZN(n9984) );
  INV_X1 U11663 ( .A(n13534), .ZN(n9985) );
  INV_X1 U11664 ( .A(n10278), .ZN(n10238) );
  XNOR2_X1 U11665 ( .A(n12087), .B(n12086), .ZN(n14001) );
  NOR2_X1 U11666 ( .A1(n14957), .A2(n10059), .ZN(n10058) );
  NAND2_X1 U11667 ( .A1(n14965), .A2(n9685), .ZN(n10059) );
  AND2_X1 U11668 ( .A1(n9923), .A2(n9922), .ZN(n9921) );
  INV_X1 U11669 ( .A(n13872), .ZN(n9922) );
  NAND2_X1 U11670 ( .A1(n9982), .A2(n10358), .ZN(n9981) );
  INV_X1 U11671 ( .A(n12985), .ZN(n9982) );
  NOR2_X1 U11672 ( .A1(n10599), .A2(n10598), .ZN(n10600) );
  AND3_X1 U11673 ( .A1(n10587), .A2(n10586), .A3(n10585), .ZN(n10601) );
  INV_X1 U11674 ( .A(n16061), .ZN(n9766) );
  AND2_X1 U11675 ( .A1(n10469), .A2(n10264), .ZN(n10726) );
  AOI21_X1 U11676 ( .B1(n16944), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A(n9772), .ZN(n9771) );
  INV_X1 U11677 ( .A(n10999), .ZN(n9772) );
  NOR2_X1 U11678 ( .A1(n13978), .A2(n16692), .ZN(n10889) );
  NOR2_X1 U11679 ( .A1(n9905), .A2(n9690), .ZN(n9903) );
  AND2_X1 U11680 ( .A1(n15540), .A2(n16193), .ZN(n11125) );
  AND2_X1 U11681 ( .A1(n11059), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11061) );
  OAI21_X1 U11682 ( .B1(n10920), .B2(n16208), .A(n17546), .ZN(n10921) );
  NOR2_X1 U11683 ( .A1(n9962), .A2(n9963), .ZN(n9961) );
  INV_X1 U11684 ( .A(n10899), .ZN(n10900) );
  NAND2_X1 U11685 ( .A1(n20678), .A2(n13588), .ZN(n13848) );
  OR2_X1 U11686 ( .A1(n15580), .A2(n12160), .ZN(n12170) );
  NOR2_X1 U11687 ( .A1(n15744), .A2(n13379), .ZN(n13312) );
  NAND2_X1 U11688 ( .A1(n14058), .A2(n10041), .ZN(n10040) );
  INV_X1 U11689 ( .A(n10041), .ZN(n10039) );
  OAI21_X1 U11690 ( .B1(n11471), .B2(n14433), .A(n11904), .ZN(n14176) );
  AND2_X1 U11691 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n11769), .ZN(
        n11770) );
  INV_X1 U11692 ( .A(n11768), .ZN(n11769) );
  NAND2_X1 U11693 ( .A1(n11770), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11814) );
  AND2_X1 U11694 ( .A1(n11734), .A2(n9742), .ZN(n10028) );
  INV_X1 U11695 ( .A(n14273), .ZN(n11734) );
  NAND2_X1 U11696 ( .A1(n12008), .A2(n14479), .ZN(n9782) );
  NOR2_X1 U11697 ( .A1(n10031), .A2(n10030), .ZN(n10029) );
  NAND2_X1 U11698 ( .A1(n10032), .A2(n9730), .ZN(n10031) );
  INV_X1 U11699 ( .A(n13894), .ZN(n10030) );
  NAND2_X1 U11700 ( .A1(n13892), .A2(n13894), .ZN(n13893) );
  INV_X1 U11701 ( .A(n13765), .ZN(n11499) );
  AOI21_X1 U11702 ( .B1(n11974), .B2(n11625), .A(n11521), .ZN(n13791) );
  INV_X1 U11703 ( .A(n13266), .ZN(n14129) );
  NOR2_X1 U11704 ( .A1(n14419), .A2(n14410), .ZN(n10011) );
  NOR2_X1 U11705 ( .A1(n14406), .A2(n14584), .ZN(n14016) );
  NAND2_X1 U11706 ( .A1(n14497), .A2(n14498), .ZN(n12006) );
  NOR2_X1 U11707 ( .A1(n11356), .A2(n11355), .ZN(n11357) );
  INV_X1 U11708 ( .A(n11439), .ZN(n9788) );
  NAND2_X1 U11709 ( .A1(n9664), .A2(n20578), .ZN(n11437) );
  AND2_X1 U11710 ( .A1(n20006), .A2(n20657), .ZN(n20011) );
  INV_X1 U11711 ( .A(n20152), .ZN(n20405) );
  AND2_X1 U11712 ( .A1(n20160), .A2(n20338), .ZN(n20474) );
  NOR2_X1 U11713 ( .A1(n13656), .A2(n9591), .ZN(n20465) );
  NOR2_X1 U11714 ( .A1(n12053), .A2(n12022), .ZN(n12056) );
  AOI221_X1 U11715 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n12023), 
        .C1(n11469), .C2(n12023), .A(n12021), .ZN(n12167) );
  NOR2_X1 U11716 ( .A1(n15580), .A2(n15585), .ZN(n15570) );
  OR2_X1 U11717 ( .A1(n15931), .A2(n18865), .ZN(n9840) );
  INV_X1 U11718 ( .A(n12423), .ZN(n10790) );
  AND2_X1 U11719 ( .A1(n12409), .A2(n12408), .ZN(n15945) );
  NOR2_X1 U11720 ( .A1(n15965), .A2(n18865), .ZN(n15958) );
  OR2_X1 U11721 ( .A1(n15958), .A2(n15959), .ZN(n9829) );
  AND2_X1 U11722 ( .A1(n12340), .A2(n12339), .ZN(n18798) );
  INV_X1 U11723 ( .A(n10239), .ZN(n10268) );
  AND2_X1 U11724 ( .A1(n12619), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13700) );
  NAND2_X1 U11725 ( .A1(n12775), .A2(n10080), .ZN(n14824) );
  XNOR2_X1 U11726 ( .A(n10101), .B(n10100), .ZN(n14051) );
  NAND2_X1 U11727 ( .A1(n10102), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10101) );
  NAND2_X1 U11728 ( .A1(n10111), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10110) );
  NOR2_X2 U11729 ( .A1(n14856), .A2(n14855), .ZN(n14857) );
  NOR2_X2 U11730 ( .A1(n13729), .A2(n13730), .ZN(n13731) );
  INV_X1 U11731 ( .A(n12097), .ZN(n9990) );
  INV_X1 U11732 ( .A(n14935), .ZN(n14032) );
  NAND2_X1 U11733 ( .A1(n10038), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10034) );
  NAND2_X1 U11734 ( .A1(n12475), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14940) );
  NAND2_X1 U11735 ( .A1(n13994), .A2(n20693), .ZN(n13995) );
  NAND2_X1 U11736 ( .A1(n9823), .A2(n9820), .ZN(n12418) );
  NAND2_X1 U11737 ( .A1(n9822), .A2(n9821), .ZN(n9820) );
  NAND2_X1 U11738 ( .A1(n9826), .A2(n9824), .ZN(n9823) );
  INV_X1 U11739 ( .A(n10058), .ZN(n9822) );
  INV_X1 U11740 ( .A(n15367), .ZN(n15366) );
  AND2_X1 U11741 ( .A1(n9709), .A2(n15325), .ZN(n9817) );
  AND2_X1 U11742 ( .A1(n13565), .A2(n15394), .ZN(n9908) );
  NAND2_X1 U11743 ( .A1(n13571), .A2(n13830), .ZN(n9816) );
  OR2_X1 U11744 ( .A1(n13571), .A2(n13830), .ZN(n9815) );
  AOI21_X1 U11745 ( .B1(n18872), .B2(n12600), .A(n12599), .ZN(n13148) );
  XNOR2_X1 U11746 ( .A(n12611), .B(n12609), .ZN(n13220) );
  AND2_X1 U11747 ( .A1(n19304), .A2(n19303), .ZN(n19278) );
  NOR2_X1 U11748 ( .A1(n19304), .A2(n19303), .ZN(n19498) );
  INV_X1 U11749 ( .A(n19544), .ZN(n19338) );
  NAND2_X1 U11750 ( .A1(n11046), .A2(n11040), .ZN(n11072) );
  NOR2_X1 U11751 ( .A1(n13969), .A2(n17224), .ZN(n18420) );
  INV_X1 U11752 ( .A(n12191), .ZN(n18428) );
  INV_X1 U11753 ( .A(n17293), .ZN(n9892) );
  NOR2_X1 U11754 ( .A1(n16402), .A2(n17306), .ZN(n16401) );
  AND2_X1 U11755 ( .A1(n9901), .A2(n9737), .ZN(n16430) );
  INV_X1 U11756 ( .A(n17348), .ZN(n9900) );
  OR2_X1 U11757 ( .A1(n16452), .A2(n16453), .ZN(n16450) );
  INV_X1 U11758 ( .A(n10809), .ZN(n16943) );
  NAND2_X1 U11759 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10859) );
  INV_X1 U11760 ( .A(n16693), .ZN(n9789) );
  NAND2_X1 U11761 ( .A1(n9882), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9876) );
  OR2_X1 U11762 ( .A1(n16350), .A2(n9880), .ZN(n9879) );
  NAND2_X1 U11763 ( .A1(n16350), .A2(n9878), .ZN(n9877) );
  NAND2_X1 U11764 ( .A1(n17276), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16340) );
  NOR2_X1 U11765 ( .A1(n16340), .A2(n16390), .ZN(n16350) );
  NOR2_X1 U11766 ( .A1(n17485), .A2(n17436), .ZN(n17433) );
  NOR2_X1 U11767 ( .A1(n17291), .A2(n10938), .ZN(n15540) );
  OR2_X1 U11768 ( .A1(n17431), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10938) );
  OR2_X1 U11769 ( .A1(n10934), .A2(n10084), .ZN(n10935) );
  OAI211_X1 U11770 ( .C1(n17314), .C2(n17678), .A(n17313), .B(n9744), .ZN(
        n17302) );
  NAND2_X1 U11771 ( .A1(n9795), .A2(n17666), .ZN(n9796) );
  INV_X1 U11772 ( .A(n17302), .ZN(n9795) );
  OR2_X1 U11773 ( .A1(n17431), .A2(n17328), .ZN(n17313) );
  NOR3_X1 U11774 ( .A1(n17328), .A2(n17350), .A3(n17702), .ZN(n17314) );
  OR2_X1 U11775 ( .A1(n17845), .A2(n17546), .ZN(n9808) );
  NOR2_X2 U11776 ( .A1(n11022), .A2(n11021), .ZN(n18631) );
  INV_X1 U11777 ( .A(n9961), .ZN(n9801) );
  INV_X1 U11778 ( .A(n17570), .ZN(n9799) );
  NAND2_X1 U11779 ( .A1(n9962), .A2(n17585), .ZN(n9960) );
  NOR2_X1 U11780 ( .A1(n10915), .A2(n9966), .ZN(n9963) );
  NAND2_X1 U11781 ( .A1(n13965), .A2(n13964), .ZN(n18419) );
  OR3_X1 U11782 ( .A1(n15580), .A2(n19756), .A3(n15560), .ZN(n19944) );
  INV_X1 U11783 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20665) );
  NOR2_X1 U11784 ( .A1(n16173), .A2(n13030), .ZN(n13031) );
  OR2_X1 U11785 ( .A1(n16142), .A2(n18657), .ZN(n19735) );
  AND2_X1 U11786 ( .A1(n9840), .A2(n9839), .ZN(n15925) );
  OAI21_X1 U11787 ( .B1(n9840), .B2(n9839), .A(n18882), .ZN(n9838) );
  OR2_X1 U11788 ( .A1(n14869), .A2(n14868), .ZN(n15092) );
  OR2_X1 U11789 ( .A1(n13043), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n18871) );
  INV_X1 U11790 ( .A(n18874), .ZN(n18901) );
  NAND2_X1 U11791 ( .A1(n9941), .A2(n9946), .ZN(n9944) );
  INV_X1 U11792 ( .A(n9942), .ZN(n9941) );
  INV_X1 U11793 ( .A(n19706), .ZN(n19026) );
  XNOR2_X1 U11794 ( .A(n12085), .B(n10758), .ZN(n18905) );
  OR2_X1 U11795 ( .A1(n13128), .A2(n12940), .ZN(n12941) );
  INV_X1 U11796 ( .A(n18953), .ZN(n18963) );
  AND2_X1 U11797 ( .A1(n13110), .A2(n19744), .ZN(n18990) );
  AND2_X1 U11798 ( .A1(n16059), .A2(n19702), .ZN(n16067) );
  AND2_X1 U11799 ( .A1(n16059), .A2(n13115), .ZN(n16052) );
  INV_X1 U11800 ( .A(n16052), .ZN(n19025) );
  NAND2_X1 U11801 ( .A1(n12441), .A2(n13720), .ZN(n16072) );
  INV_X1 U11802 ( .A(n16067), .ZN(n19020) );
  NAND2_X1 U11803 ( .A1(n18905), .A2(n15410), .ZN(n14045) );
  INV_X1 U11804 ( .A(n15087), .ZN(n9915) );
  NAND2_X1 U11805 ( .A1(n15086), .A2(n9914), .ZN(n9913) );
  INV_X1 U11806 ( .A(n15084), .ZN(n9914) );
  AND2_X1 U11807 ( .A1(n12084), .A2(n12085), .ZN(n15085) );
  AND2_X1 U11808 ( .A1(n12579), .A2(n19723), .ZN(n16105) );
  OR2_X1 U11809 ( .A1(n12578), .A2(n12564), .ZN(n16097) );
  OR2_X1 U11810 ( .A1(n12578), .A2(n19724), .ZN(n15405) );
  INV_X1 U11811 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19710) );
  NAND2_X1 U11812 ( .A1(n12601), .A2(n12600), .ZN(n12604) );
  AND2_X1 U11813 ( .A1(n19278), .A2(n19476), .ZN(n19247) );
  INV_X1 U11814 ( .A(n17223), .ZN(n17164) );
  NAND2_X1 U11815 ( .A1(n18473), .A2(n18483), .ZN(n16320) );
  INV_X1 U11816 ( .A(n16361), .ZN(n9873) );
  XNOR2_X1 U11817 ( .A(n16359), .B(n9875), .ZN(n9874) );
  INV_X1 U11818 ( .A(n16360), .ZN(n9875) );
  INV_X1 U11819 ( .A(n16696), .ZN(n20820) );
  NOR2_X1 U11820 ( .A1(n10827), .A2(n10826), .ZN(n17133) );
  NOR2_X1 U11821 ( .A1(n17158), .A2(n18024), .ZN(n17149) );
  OR2_X1 U11822 ( .A1(n9969), .A2(n16189), .ZN(n9968) );
  NOR2_X1 U11823 ( .A1(n17845), .A2(n10925), .ZN(n17551) );
  NOR2_X1 U11824 ( .A1(n9712), .A2(n11129), .ZN(n16190) );
  AOI22_X1 U11825 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10175) );
  INV_X1 U11826 ( .A(n12036), .ZN(n12032) );
  AOI22_X1 U11827 ( .A1(n12029), .A2(n12028), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20407), .ZN(n12025) );
  AND2_X1 U11828 ( .A1(n11438), .A2(n11478), .ZN(n9787) );
  OR2_X1 U11829 ( .A1(n11464), .A2(n11463), .ZN(n11965) );
  OAI21_X1 U11830 ( .B1(n11275), .B2(n11231), .A(n11294), .ZN(n11282) );
  NOR2_X1 U11831 ( .A1(n12025), .A2(n12026), .ZN(n12024) );
  AOI21_X1 U11832 ( .B1(n10429), .B2(n10427), .A(n10418), .ZN(n10426) );
  NAND2_X1 U11833 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12893) );
  AOI22_X1 U11834 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12278), .B1(
        n12305), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12241) );
  AND2_X1 U11835 ( .A1(n12514), .A2(n10271), .ZN(n10260) );
  NAND2_X1 U11836 ( .A1(n9704), .A2(n12218), .ZN(n12312) );
  AND4_X1 U11837 ( .A1(n10133), .A2(n10132), .A3(n10131), .A4(n10130), .ZN(
        n10134) );
  AND3_X1 U11838 ( .A1(n10138), .A2(n10137), .A3(n10136), .ZN(n10142) );
  AOI21_X1 U11839 ( .B1(n10226), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n10139), .ZN(n10141) );
  NAND2_X1 U11840 ( .A1(n18590), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10807) );
  NAND2_X1 U11841 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18612), .ZN(
        n10810) );
  AOI21_X1 U11842 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18457), .A(
        n11051), .ZN(n11053) );
  NAND3_X1 U11843 ( .A1(n11301), .A2(n11283), .A3(n11302), .ZN(n13188) );
  NOR2_X1 U11844 ( .A1(n14153), .A2(n10042), .ZN(n10041) );
  AND2_X1 U11845 ( .A1(n11642), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11646) );
  OR2_X1 U11846 ( .A1(n9722), .A2(n11601), .ZN(n10032) );
  NAND2_X1 U11847 ( .A1(n9591), .A2(n11478), .ZN(n9846) );
  NOR2_X1 U11848 ( .A1(n14160), .A2(n9858), .ZN(n9857) );
  INV_X1 U11849 ( .A(n14163), .ZN(n9858) );
  INV_X1 U11850 ( .A(n14220), .ZN(n9868) );
  OR2_X1 U11851 ( .A1(n15785), .A2(n14737), .ZN(n12010) );
  AND2_X1 U11852 ( .A1(n14318), .A2(n14312), .ZN(n9869) );
  NOR2_X1 U11853 ( .A1(n14324), .A2(n14323), .ZN(n14319) );
  AND2_X1 U11854 ( .A1(n13555), .A2(n9865), .ZN(n9864) );
  INV_X1 U11855 ( .A(n15899), .ZN(n9865) );
  INV_X1 U11856 ( .A(n14101), .ZN(n14113) );
  NAND2_X1 U11857 ( .A1(n10017), .A2(n10018), .ZN(n11946) );
  AOI21_X1 U11858 ( .B1(n10020), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11939), 
        .ZN(n10018) );
  NAND2_X1 U11860 ( .A1(n11348), .A2(n11347), .ZN(n11411) );
  OR2_X1 U11861 ( .A1(n11386), .A2(n11385), .ZN(n11387) );
  INV_X1 U11862 ( .A(n11387), .ZN(n11950) );
  AND3_X1 U11863 ( .A1(n11353), .A2(n11352), .A3(n11351), .ZN(n11354) );
  OR2_X1 U11864 ( .A1(n11435), .A2(n11434), .ZN(n11966) );
  AOI21_X1 U11865 ( .B1(n11275), .B2(n11236), .A(n13236), .ZN(n11237) );
  AND2_X1 U11866 ( .A1(n10048), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11157) );
  INV_X1 U11867 ( .A(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11246) );
  INV_X1 U11868 ( .A(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11245) );
  INV_X1 U11869 ( .A(n12053), .ZN(n12057) );
  NAND2_X1 U11870 ( .A1(n13191), .A2(n11267), .ZN(n11271) );
  OR2_X1 U11871 ( .A1(n13649), .A2(n13648), .ZN(n15565) );
  NOR2_X1 U11872 ( .A1(n10008), .A2(n12402), .ZN(n10007) );
  NAND2_X1 U11873 ( .A1(n12337), .A2(n10002), .ZN(n12346) );
  AND2_X1 U11874 ( .A1(n12337), .A2(n10777), .ZN(n12342) );
  NAND2_X1 U11875 ( .A1(n12270), .A2(n12269), .ZN(n12302) );
  NAND2_X1 U11876 ( .A1(n10300), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10288) );
  CLKBUF_X1 U11877 ( .A(n12754), .Z(n12929) );
  NAND2_X1 U11878 ( .A1(n12847), .A2(n9935), .ZN(n9934) );
  OR2_X1 U11879 ( .A1(n14815), .A2(n9746), .ZN(n9936) );
  INV_X1 U11880 ( .A(n12871), .ZN(n9935) );
  AND2_X1 U11881 ( .A1(n9931), .A2(n9930), .ZN(n9929) );
  INV_X1 U11882 ( .A(n14908), .ZN(n9930) );
  AND2_X1 U11883 ( .A1(n14752), .A2(n12999), .ZN(n9931) );
  AND3_X1 U11884 ( .A1(n10268), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13720), 
        .ZN(n12869) );
  INV_X1 U11885 ( .A(n13869), .ZN(n9956) );
  NOR2_X1 U11886 ( .A1(n16058), .A2(n9834), .ZN(n9833) );
  INV_X1 U11887 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n9834) );
  NAND2_X1 U11888 ( .A1(n9992), .A2(n12477), .ZN(n9991) );
  NOR2_X1 U11889 ( .A1(n9994), .A2(n13009), .ZN(n9992) );
  INV_X1 U11890 ( .A(n14024), .ZN(n9994) );
  NAND2_X1 U11891 ( .A1(n9928), .A2(n9927), .ZN(n9926) );
  INV_X1 U11892 ( .A(n12562), .ZN(n9927) );
  NOR2_X1 U11893 ( .A1(n15096), .A2(n20693), .ZN(n10038) );
  NOR2_X1 U11894 ( .A1(n13997), .A2(n9825), .ZN(n9824) );
  INV_X1 U11895 ( .A(n12406), .ZN(n9825) );
  OR2_X1 U11896 ( .A1(n10046), .A2(n12557), .ZN(n10045) );
  NAND2_X1 U11897 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10046) );
  AND2_X1 U11898 ( .A1(n14764), .A2(n14752), .ZN(n14754) );
  NOR2_X1 U11899 ( .A1(n10052), .A2(n15285), .ZN(n10051) );
  INV_X1 U11900 ( .A(n15265), .ZN(n10052) );
  OR2_X1 U11901 ( .A1(n10548), .A2(n10547), .ZN(n12277) );
  NAND2_X1 U11902 ( .A1(n10324), .A2(n9988), .ZN(n9987) );
  INV_X1 U11903 ( .A(n13325), .ZN(n9988) );
  AOI21_X1 U11904 ( .B1(n10300), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10314), .ZN(n10316) );
  OR2_X1 U11905 ( .A1(n10325), .A2(n10536), .ZN(n10313) );
  OR2_X1 U11906 ( .A1(n10533), .A2(n10532), .ZN(n12254) );
  CLKBUF_X1 U11907 ( .A(n12521), .Z(n12541) );
  NAND2_X1 U11908 ( .A1(n10198), .A2(n10136), .ZN(n10205) );
  NAND2_X1 U11909 ( .A1(n10203), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10204) );
  INV_X1 U11910 ( .A(n12229), .ZN(n12236) );
  AOI22_X1 U11911 ( .A1(n12812), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10224) );
  AND2_X1 U11912 ( .A1(n10228), .A2(n10227), .ZN(n10229) );
  NAND3_X1 U11913 ( .A1(n19688), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19544), 
        .ZN(n13716) );
  AND2_X1 U11914 ( .A1(n12503), .A2(n10431), .ZN(n16131) );
  NOR2_X1 U11915 ( .A1(n17995), .A2(n11025), .ZN(n11030) );
  OR2_X1 U11916 ( .A1(n16693), .A2(n10807), .ZN(n15509) );
  NOR2_X1 U11917 ( .A1(n10808), .A2(n10807), .ZN(n10852) );
  NOR3_X1 U11918 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18604), .A3(
        n13978), .ZN(n10842) );
  NOR2_X1 U11919 ( .A1(n11044), .A2(n11073), .ZN(n13969) );
  AND2_X1 U11920 ( .A1(n9881), .A2(n9880), .ZN(n9878) );
  NAND2_X1 U11921 ( .A1(n17349), .A2(n17377), .ZN(n17378) );
  INV_X1 U11922 ( .A(n16318), .ZN(n11073) );
  NAND2_X1 U11923 ( .A1(n9697), .A2(n9961), .ZN(n9797) );
  NAND2_X1 U11924 ( .A1(n17600), .A2(n9697), .ZN(n9798) );
  OR2_X1 U11925 ( .A1(n18024), .A2(n15590), .ZN(n11042) );
  NOR2_X1 U11926 ( .A1(n10950), .A2(n10949), .ZN(n11037) );
  NAND2_X1 U11927 ( .A1(n17880), .A2(n11069), .ZN(n16213) );
  AND2_X1 U11928 ( .A1(n11685), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11698) );
  NAND2_X1 U11929 ( .A1(n13271), .A2(n13266), .ZN(n9854) );
  OR2_X1 U11930 ( .A1(n13349), .A2(n13348), .ZN(n13544) );
  INV_X1 U11931 ( .A(n20001), .ZN(n20002) );
  AND2_X1 U11932 ( .A1(n14412), .A2(n12150), .ZN(n12151) );
  OR2_X1 U11933 ( .A1(n12104), .A2(n12103), .ZN(n13589) );
  AND2_X1 U11934 ( .A1(n11883), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11884) );
  AOI21_X1 U11935 ( .B1(n12150), .B2(n14444), .A(n11881), .ZN(n14189) );
  AND2_X1 U11936 ( .A1(n11842), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11843) );
  NAND2_X1 U11937 ( .A1(n11843), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11882) );
  AND2_X1 U11938 ( .A1(n10025), .A2(n11840), .ZN(n10024) );
  NOR2_X1 U11939 ( .A1(n11814), .A2(n15617), .ZN(n11815) );
  NAND2_X1 U11940 ( .A1(n11815), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11841) );
  AND2_X1 U11941 ( .A1(n15620), .A2(n12150), .ZN(n11787) );
  AND2_X1 U11942 ( .A1(n11772), .A2(n11771), .ZN(n14257) );
  NOR2_X1 U11943 ( .A1(n11730), .A2(n11729), .ZN(n11731) );
  NAND2_X1 U11944 ( .A1(n11731), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11768) );
  NAND2_X1 U11945 ( .A1(n11698), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11730) );
  AND2_X1 U11946 ( .A1(n11646), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11665) );
  INV_X1 U11947 ( .A(n14298), .ZN(n11663) );
  NOR2_X1 U11948 ( .A1(n11628), .A2(n15709), .ZN(n11642) );
  INV_X1 U11949 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15709) );
  NAND2_X1 U11950 ( .A1(n11584), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11628) );
  NAND2_X1 U11951 ( .A1(n11550), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11565) );
  INV_X1 U11952 ( .A(n13909), .ZN(n11564) );
  CLKBUF_X1 U11953 ( .A(n13794), .Z(n13795) );
  AND2_X1 U11954 ( .A1(n11518), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11530) );
  INV_X1 U11955 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11494) );
  NOR2_X1 U11956 ( .A1(n11495), .A2(n11494), .ZN(n11518) );
  NAND2_X1 U11957 ( .A1(n11473), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11495) );
  CLKBUF_X1 U11958 ( .A(n13546), .Z(n13547) );
  NAND2_X1 U11959 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11443) );
  OR2_X1 U11960 ( .A1(n14246), .A2(n14202), .ZN(n14204) );
  NAND2_X1 U11961 ( .A1(n14638), .A2(n14244), .ZN(n14246) );
  NAND2_X1 U11962 ( .A1(n14269), .A2(n9745), .ZN(n14636) );
  INV_X1 U11963 ( .A(n14252), .ZN(n9870) );
  OAI21_X1 U11964 ( .B1(n14490), .B2(n9773), .A(n9590), .ZN(n14469) );
  NAND2_X1 U11965 ( .A1(n14269), .A2(n9741), .ZN(n14261) );
  NAND2_X1 U11966 ( .A1(n14269), .A2(n14266), .ZN(n14265) );
  OR2_X1 U11967 ( .A1(n14284), .A2(n14277), .ZN(n14279) );
  NOR2_X1 U11968 ( .A1(n14279), .A2(n14268), .ZN(n14269) );
  NAND2_X1 U11969 ( .A1(n14294), .A2(n14282), .ZN(n14284) );
  AND2_X1 U11970 ( .A1(n14302), .A2(n14292), .ZN(n14294) );
  OR2_X1 U11971 ( .A1(n15785), .A2(n15837), .ZN(n15772) );
  OR2_X1 U11972 ( .A1(n15785), .A2(n12004), .ZN(n15768) );
  AND2_X1 U11973 ( .A1(n14319), .A2(n9866), .ZN(n14302) );
  AND2_X1 U11974 ( .A1(n9727), .A2(n9867), .ZN(n9866) );
  INV_X1 U11975 ( .A(n14299), .ZN(n9867) );
  NAND2_X1 U11976 ( .A1(n14319), .A2(n9727), .ZN(n14300) );
  NOR2_X1 U11977 ( .A1(n14520), .A2(n9786), .ZN(n14505) );
  OR2_X1 U11978 ( .A1(n12001), .A2(n14519), .ZN(n9786) );
  INV_X1 U11979 ( .A(n14520), .ZN(n9785) );
  INV_X1 U11980 ( .A(n12001), .ZN(n9784) );
  NAND2_X1 U11981 ( .A1(n14319), .A2(n9869), .ZN(n14314) );
  INV_X1 U11982 ( .A(n19987), .ZN(n14736) );
  INV_X1 U11983 ( .A(n11998), .ZN(n9779) );
  AND2_X1 U11984 ( .A1(n13902), .A2(n13901), .ZN(n13907) );
  OR2_X1 U11985 ( .A1(n15860), .A2(n13907), .ZN(n14324) );
  OR2_X1 U11986 ( .A1(n15858), .A2(n15857), .ZN(n15860) );
  INV_X1 U11987 ( .A(n11981), .ZN(n9776) );
  INV_X1 U11988 ( .A(n11973), .ZN(n9775) );
  AND2_X1 U11989 ( .A1(n13807), .A2(n13806), .ZN(n13808) );
  NAND2_X1 U11990 ( .A1(n13556), .A2(n9864), .ZN(n15896) );
  NAND2_X1 U11991 ( .A1(n13556), .A2(n13555), .ZN(n15898) );
  INV_X1 U11992 ( .A(n13525), .ZN(n10016) );
  NAND2_X1 U11993 ( .A1(n13526), .A2(n13525), .ZN(n13528) );
  AND2_X1 U11994 ( .A1(n15869), .A2(n14736), .ZN(n14557) );
  AND2_X1 U11995 ( .A1(n14536), .A2(n19990), .ZN(n14534) );
  NAND2_X1 U11996 ( .A1(n11288), .A2(n11345), .ZN(n11405) );
  OR3_X1 U11997 ( .A1(n13450), .A2(n13449), .A3(n13448), .ZN(n13646) );
  NOR2_X1 U11998 ( .A1(n13656), .A2(n11438), .ZN(n20249) );
  INV_X1 U11999 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20406) );
  AND2_X1 U12000 ( .A1(n13657), .A2(n20658), .ZN(n20248) );
  AOI21_X1 U12001 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20665), .A(n20052), 
        .ZN(n20523) );
  AND2_X1 U12002 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20160), .ZN(n20042) );
  OAI221_X2 U12003 ( .B1(n15915), .B2(n20649), .C1(n15920), .C2(n20649), .A(
        n20578), .ZN(n20052) );
  AND2_X1 U12004 ( .A1(n10774), .A2(n10771), .ZN(n12502) );
  INV_X1 U12005 ( .A(n15926), .ZN(n9839) );
  NOR2_X1 U12006 ( .A1(n10004), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10003) );
  INV_X1 U12007 ( .A(n10005), .ZN(n10004) );
  NAND2_X1 U12008 ( .A1(n10786), .A2(n10005), .ZN(n15968) );
  OR2_X1 U12009 ( .A1(n12994), .A2(n14993), .ZN(n9827) );
  NAND2_X1 U12010 ( .A1(n12381), .A2(n9998), .ZN(n12372) );
  AND2_X1 U12011 ( .A1(n10002), .A2(n10001), .ZN(n10000) );
  NAND2_X1 U12012 ( .A1(n12349), .A2(n12355), .ZN(n12359) );
  XNOR2_X1 U12013 ( .A(n12302), .B(n12301), .ZN(n18845) );
  CLKBUF_X1 U12014 ( .A(n10792), .Z(n12536) );
  INV_X1 U12015 ( .A(n10755), .ZN(n10756) );
  NOR2_X1 U12016 ( .A1(n14805), .A2(n14804), .ZN(n14803) );
  XNOR2_X1 U12017 ( .A(n12825), .B(n12826), .ZN(n14820) );
  NAND2_X1 U12018 ( .A1(n14764), .A2(n9931), .ZN(n14907) );
  NOR2_X1 U12019 ( .A1(n9949), .A2(n14837), .ZN(n9948) );
  INV_X1 U12020 ( .A(n9952), .ZN(n9949) );
  NAND2_X1 U12021 ( .A1(n9687), .A2(n14850), .ZN(n9954) );
  NAND2_X1 U12022 ( .A1(n12980), .A2(n9921), .ZN(n15196) );
  NAND2_X1 U12023 ( .A1(n12980), .A2(n9923), .ZN(n15233) );
  CLKBUF_X1 U12024 ( .A(n13869), .Z(n13870) );
  AND2_X1 U12025 ( .A1(n12980), .A2(n12981), .ZN(n15232) );
  AND2_X1 U12026 ( .A1(n9726), .A2(n15331), .ZN(n9917) );
  NOR2_X1 U12027 ( .A1(n10270), .A2(n10256), .ZN(n10240) );
  OAI21_X1 U12028 ( .B1(n10755), .B2(n18674), .A(n10475), .ZN(n13211) );
  INV_X1 U12029 ( .A(n13052), .ZN(n13717) );
  NAND2_X1 U12030 ( .A1(n9845), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10105) );
  NOR2_X1 U12031 ( .A1(n10105), .A2(n14941), .ZN(n10102) );
  NAND2_X1 U12032 ( .A1(n10107), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10109) );
  OR2_X1 U12033 ( .A1(n14749), .A2(n12997), .ZN(n14832) );
  NOR2_X2 U12034 ( .A1(n14832), .A2(n14833), .ZN(n14831) );
  AND2_X1 U12035 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n10099), .ZN(
        n10111) );
  AND2_X1 U12036 ( .A1(n12395), .A2(n15029), .ZN(n12396) );
  NAND2_X1 U12037 ( .A1(n14758), .A2(n14759), .ZN(n14761) );
  AND2_X1 U12038 ( .A1(n9686), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9830) );
  NAND2_X1 U12039 ( .A1(n10115), .A2(n9686), .ZN(n10128) );
  NAND2_X1 U12040 ( .A1(n9979), .A2(n9978), .ZN(n9977) );
  INV_X1 U12041 ( .A(n13938), .ZN(n9978) );
  NAND2_X1 U12042 ( .A1(n9976), .A2(n9979), .ZN(n13937) );
  INV_X1 U12043 ( .A(n13699), .ZN(n9976) );
  NAND2_X1 U12044 ( .A1(n9842), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9841) );
  INV_X1 U12045 ( .A(n9843), .ZN(n9842) );
  NAND2_X1 U12046 ( .A1(n10118), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10127) );
  INV_X1 U12047 ( .A(n13780), .ZN(n9983) );
  NAND2_X1 U12048 ( .A1(n13535), .A2(n9703), .ZN(n13779) );
  NAND2_X1 U12049 ( .A1(n10121), .A2(n9679), .ZN(n10126) );
  NAND2_X1 U12050 ( .A1(n13535), .A2(n13534), .ZN(n13674) );
  NAND2_X1 U12051 ( .A1(n10121), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10125) );
  INV_X1 U12052 ( .A(n15074), .ZN(n10062) );
  INV_X1 U12053 ( .A(n15072), .ZN(n10061) );
  INV_X1 U12054 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15076) );
  NOR2_X1 U12055 ( .A1(n13921), .A2(n9836), .ZN(n9835) );
  NAND2_X1 U12056 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9836) );
  NOR2_X1 U12057 ( .A1(n10122), .A2(n20796), .ZN(n10124) );
  NAND2_X1 U12058 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10122) );
  INV_X1 U12059 ( .A(n10300), .ZN(n10311) );
  INV_X1 U12060 ( .A(n10038), .ZN(n10037) );
  NAND2_X1 U12061 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10036) );
  INV_X1 U12062 ( .A(n14979), .ZN(n14036) );
  INV_X1 U12063 ( .A(n15922), .ZN(n13999) );
  NAND2_X1 U12064 ( .A1(n15922), .A2(n9754), .ZN(n14935) );
  NAND2_X1 U12065 ( .A1(n14940), .A2(n9759), .ZN(n12580) );
  NAND2_X1 U12066 ( .A1(n9760), .A2(n20693), .ZN(n9759) );
  NOR2_X1 U12067 ( .A1(n13007), .A2(n14002), .ZN(n13990) );
  OAI21_X1 U12068 ( .B1(n12411), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12412), .ZN(n14957) );
  OR2_X1 U12069 ( .A1(n10045), .A2(n15116), .ZN(n10044) );
  INV_X1 U12070 ( .A(n12472), .ZN(n9765) );
  INV_X1 U12071 ( .A(n15164), .ZN(n9764) );
  INV_X1 U12072 ( .A(n15195), .ZN(n9920) );
  NOR2_X1 U12073 ( .A1(n13699), .A2(n9981), .ZN(n13930) );
  NAND2_X1 U12074 ( .A1(n15361), .A2(n9726), .ZN(n15352) );
  INV_X1 U12075 ( .A(n10063), .ZN(n9818) );
  AND2_X1 U12076 ( .A1(n12569), .A2(n13576), .ZN(n15316) );
  INV_X1 U12077 ( .A(n16060), .ZN(n9762) );
  AND2_X1 U12078 ( .A1(n10064), .A2(n16063), .ZN(n10063) );
  OR2_X1 U12079 ( .A1(n16064), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10064) );
  AND2_X1 U12080 ( .A1(n16064), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10065) );
  AND2_X1 U12081 ( .A1(n18823), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15072) );
  OAI21_X1 U12082 ( .B1(n12465), .B2(n12463), .A(n12462), .ZN(n15380) );
  INV_X1 U12083 ( .A(n12460), .ZN(n13917) );
  AND2_X1 U12084 ( .A1(n10258), .A2(n10255), .ZN(n10230) );
  INV_X1 U12085 ( .A(n19368), .ZN(n19372) );
  NAND2_X1 U12086 ( .A1(n10185), .A2(n10136), .ZN(n10192) );
  NAND2_X1 U12087 ( .A1(n10190), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10191) );
  NAND2_X1 U12088 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19544), .ZN(n19049) );
  NOR2_X2 U12089 ( .A1(n13715), .A2(n13716), .ZN(n19062) );
  INV_X1 U12090 ( .A(n19540), .ZN(n19497) );
  OR2_X1 U12091 ( .A1(n19304), .A2(n19716), .ZN(n19475) );
  INV_X1 U12092 ( .A(n19049), .ZN(n19067) );
  AND2_X1 U12093 ( .A1(n13133), .A2(n13132), .ZN(n16129) );
  INV_X1 U12094 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19733) );
  NAND2_X1 U12095 ( .A1(n16646), .A2(n17991), .ZN(n11044) );
  NOR2_X1 U12096 ( .A1(n11011), .A2(n11010), .ZN(n11050) );
  INV_X1 U12097 ( .A(n11030), .ZN(n11041) );
  INV_X1 U12098 ( .A(n18645), .ZN(n18634) );
  AND2_X1 U12099 ( .A1(n16379), .A2(n9732), .ZN(n16366) );
  NOR2_X1 U12100 ( .A1(n16366), .A2(n16367), .ZN(n16365) );
  NAND2_X1 U12101 ( .A1(n9891), .A2(n9732), .ZN(n9888) );
  OR2_X1 U12103 ( .A1(n16381), .A2(n16382), .ZN(n16379) );
  INV_X1 U12104 ( .A(n16340), .ZN(n16341) );
  AND2_X1 U12105 ( .A1(n16422), .A2(n9732), .ZN(n16409) );
  OR2_X1 U12106 ( .A1(n16424), .A2(n17331), .ZN(n16422) );
  NOR2_X1 U12107 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16512), .ZN(n16496) );
  NOR2_X1 U12108 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16562), .ZN(n16543) );
  NOR2_X1 U12109 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16638), .ZN(n16624) );
  INV_X1 U12110 ( .A(n17604), .ZN(n16642) );
  NOR2_X1 U12111 ( .A1(n10997), .A2(n9770), .ZN(n9769) );
  NAND2_X1 U12112 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17123), .ZN(n17119) );
  AOI22_X1 U12113 ( .A1(n10877), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10841) );
  NAND2_X1 U12114 ( .A1(n10853), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10838) );
  NOR2_X1 U12115 ( .A1(n18490), .A2(n18424), .ZN(n17223) );
  NAND2_X1 U12116 ( .A1(n16350), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16349) );
  NOR2_X1 U12117 ( .A1(n17305), .A2(n17304), .ZN(n17276) );
  NOR2_X1 U12118 ( .A1(n17788), .A2(n17649), .ZN(n17274) );
  AND2_X1 U12119 ( .A1(n17408), .A2(n9688), .ZN(n17330) );
  NAND2_X1 U12120 ( .A1(n17408), .A2(n9903), .ZN(n17339) );
  INV_X1 U12121 ( .A(n17486), .ZN(n17407) );
  NOR2_X1 U12122 ( .A1(n17422), .A2(n17421), .ZN(n17408) );
  NAND2_X1 U12123 ( .A1(n9895), .A2(n9898), .ZN(n17485) );
  NOR2_X1 U12124 ( .A1(n9896), .A2(n16501), .ZN(n9895) );
  NAND2_X1 U12125 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n9734), .ZN(
        n9896) );
  NOR2_X1 U12126 ( .A1(n17587), .A2(n9894), .ZN(n9899) );
  INV_X1 U12127 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9894) );
  AND2_X1 U12128 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17604) );
  XNOR2_X1 U12129 ( .A(n10905), .B(n10903), .ZN(n17635) );
  INV_X1 U12130 ( .A(n11125), .ZN(n9802) );
  NOR2_X1 U12131 ( .A1(n17290), .A2(n10070), .ZN(n15539) );
  NAND2_X1 U12132 ( .A1(n17349), .A2(n10932), .ZN(n17329) );
  NAND2_X1 U12133 ( .A1(n17430), .A2(n11083), .ZN(n10931) );
  NAND2_X1 U12134 ( .A1(n17378), .A2(n9792), .ZN(n17350) );
  AND2_X1 U12135 ( .A1(n17364), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9792) );
  NAND2_X1 U12136 ( .A1(n17430), .A2(n17759), .ZN(n17377) );
  OAI21_X1 U12137 ( .B1(n17468), .B2(n17796), .A(n17546), .ZN(n10929) );
  AOI211_X1 U12138 ( .C1(n17468), .C2(n17546), .A(n9958), .B(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9957) );
  NOR2_X1 U12139 ( .A1(n17431), .A2(n9959), .ZN(n9958) );
  INV_X1 U12140 ( .A(n17796), .ZN(n9959) );
  NOR2_X1 U12141 ( .A1(n17820), .A2(n17429), .ZN(n17790) );
  AND2_X1 U12142 ( .A1(n10924), .A2(n9971), .ZN(n17505) );
  NOR2_X1 U12143 ( .A1(n9972), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9971) );
  INV_X1 U12144 ( .A(n9973), .ZN(n9972) );
  NOR2_X1 U12145 ( .A1(n9974), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9973) );
  INV_X1 U12146 ( .A(n9975), .ZN(n9974) );
  INV_X1 U12147 ( .A(n17789), .ZN(n18426) );
  NOR2_X1 U12148 ( .A1(n17431), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9975) );
  INV_X1 U12149 ( .A(n17845), .ZN(n17820) );
  NAND3_X1 U12150 ( .A1(n10887), .A2(n10886), .A3(n10885), .ZN(n16208) );
  OAI21_X1 U12151 ( .B1(n11066), .B2(n11065), .A(n11064), .ZN(n16317) );
  OAI211_X1 U12152 ( .C1(n17620), .C2(n9806), .A(n9804), .B(n9803), .ZN(n17612) );
  NAND2_X1 U12153 ( .A1(n17620), .A2(n9805), .ZN(n9803) );
  NOR2_X1 U12154 ( .A1(n17612), .A2(n17926), .ZN(n17611) );
  INV_X1 U12155 ( .A(n18438), .ZN(n18451) );
  NAND2_X1 U12156 ( .A1(n18634), .A2(n13971), .ZN(n18427) );
  NOR2_X1 U12157 ( .A1(n11036), .A2(n11047), .ZN(n13965) );
  AOI21_X1 U12158 ( .B1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B2(n10877), .A(
        n10900), .ZN(n10901) );
  NOR2_X1 U12159 ( .A1(n10898), .A2(n10897), .ZN(n10902) );
  NAND2_X1 U12160 ( .A1(n17642), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17641) );
  NAND3_X1 U12161 ( .A1(n10960), .A2(n10959), .A3(n10958), .ZN(n17988) );
  INV_X1 U12162 ( .A(n11050), .ZN(n17995) );
  NOR2_X2 U12163 ( .A1(n10991), .A2(n10990), .ZN(n18017) );
  NAND2_X1 U12164 ( .A1(n18486), .A2(n17986), .ZN(n18178) );
  OAI22_X1 U12165 ( .A1(n18421), .A2(n16213), .B1(n12191), .B2(n18426), .ZN(
        n18473) );
  INV_X1 U12166 ( .A(n13717), .ZN(n13715) );
  INV_X1 U12167 ( .A(n13451), .ZN(n19756) );
  NOR2_X1 U12168 ( .A1(n19820), .A2(n14217), .ZN(n15730) );
  AND3_X1 U12169 ( .A1(n13603), .A2(n13600), .A3(n13598), .ZN(n19815) );
  INV_X1 U12170 ( .A(n19816), .ZN(n19828) );
  AND2_X1 U12171 ( .A1(n13848), .A2(n13611), .ZN(n19816) );
  AND2_X1 U12172 ( .A1(n13848), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19832) );
  OR2_X1 U12173 ( .A1(n13604), .A2(n13602), .ZN(n19833) );
  AND2_X2 U12174 ( .A1(n13230), .A2(n13451), .ZN(n19858) );
  AND2_X1 U12175 ( .A1(n13312), .A2(n20002), .ZN(n15747) );
  INV_X1 U12176 ( .A(n14404), .ZN(n15748) );
  OR2_X1 U12177 ( .A1(n13450), .A2(n12173), .ZN(n12174) );
  INV_X1 U12178 ( .A(n15744), .ZN(n14401) );
  AND2_X1 U12179 ( .A1(n13248), .A2(n13247), .ZN(n19867) );
  AND2_X1 U12180 ( .A1(n13451), .A2(n15570), .ZN(n13247) );
  INV_X2 U12181 ( .A(n13468), .ZN(n19922) );
  OR2_X1 U12182 ( .A1(n11927), .A2(n11926), .ZN(n11928) );
  INV_X1 U12183 ( .A(n19938), .ZN(n19925) );
  CLKBUF_X1 U12184 ( .A(n13341), .Z(n13342) );
  AND2_X1 U12185 ( .A1(n19938), .A2(n12071), .ZN(n15781) );
  INV_X1 U12186 ( .A(n19944), .ZN(n19930) );
  XNOR2_X1 U12187 ( .A(n9859), .B(n14131), .ZN(n14563) );
  NAND2_X1 U12188 ( .A1(n14179), .A2(n9691), .ZN(n9860) );
  XNOR2_X1 U12189 ( .A(n10012), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14565) );
  NAND2_X1 U12190 ( .A1(n9780), .A2(n11998), .ZN(n13943) );
  NAND2_X1 U12191 ( .A1(n9655), .A2(n11973), .ZN(n15802) );
  NAND2_X1 U12192 ( .A1(n13272), .A2(n13266), .ZN(n13343) );
  XNOR2_X1 U12193 ( .A(n9855), .B(n13271), .ZN(n13272) );
  AND2_X1 U12194 ( .A1(n13418), .A2(n13417), .ZN(n19973) );
  AND2_X1 U12195 ( .A1(n13418), .A2(n13412), .ZN(n19993) );
  NAND2_X1 U12196 ( .A1(n9788), .A2(n11438), .ZN(n11477) );
  AOI21_X1 U12197 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20578), .A(n15907), 
        .ZN(n15906) );
  OAI211_X1 U12198 ( .C1(n20014), .C2(n20581), .A(n20335), .B(n20009), .ZN(
        n20047) );
  OAI22_X1 U12199 ( .A1(n20016), .A2(n20015), .B1(n20338), .B2(n20155), .ZN(
        n20046) );
  INV_X1 U12200 ( .A(n20067), .ZN(n20074) );
  OR2_X1 U12201 ( .A1(n20118), .A2(n20326), .ZN(n20151) );
  OAI221_X1 U12202 ( .B1(n20176), .B2(n20412), .C1(n20176), .C2(n20161), .A(
        n20474), .ZN(n20179) );
  INV_X1 U12203 ( .A(n20241), .ZN(n20202) );
  OAI211_X1 U12204 ( .C1(n20293), .C2(n20412), .A(n20335), .B(n20278), .ZN(
        n20296) );
  INV_X1 U12205 ( .A(n20271), .ZN(n20295) );
  INV_X1 U12206 ( .A(n20404), .ZN(n20391) );
  OAI211_X1 U12207 ( .C1(n20431), .C2(n20412), .A(n20474), .B(n20411), .ZN(
        n20433) );
  AND2_X1 U12208 ( .A1(n20465), .A2(n20405), .ZN(n20460) );
  OAI211_X1 U12209 ( .C1(n20505), .C2(n20475), .A(n20474), .B(n20473), .ZN(
        n20509) );
  AND2_X1 U12210 ( .A1(n11930), .A2(n20042), .ZN(n20530) );
  AND2_X1 U12211 ( .A1(n11236), .A2(n20042), .ZN(n20536) );
  AND2_X1 U12212 ( .A1(n11265), .A2(n20042), .ZN(n20548) );
  AND2_X1 U12213 ( .A1(n20032), .A2(n20042), .ZN(n20554) );
  AND2_X1 U12214 ( .A1(n11231), .A2(n20042), .ZN(n20560) );
  NOR2_X1 U12215 ( .A1(n20665), .A2(n20516), .ZN(n20566) );
  AND2_X1 U12216 ( .A1(n20465), .A2(n20248), .ZN(n20571) );
  AND2_X1 U12217 ( .A1(n11267), .A2(n20042), .ZN(n20567) );
  AND2_X2 U12218 ( .A1(n12065), .A2(n12064), .ZN(n15580) );
  INV_X1 U12219 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20577) );
  AOI21_X1 U12220 ( .B1(n18905), .B2(n18877), .A(n10798), .ZN(n10799) );
  NOR2_X1 U12221 ( .A1(n15087), .A2(n18871), .ZN(n12098) );
  NAND2_X1 U12222 ( .A1(n12095), .A2(n12094), .ZN(n12099) );
  NAND2_X1 U12223 ( .A1(n15085), .A2(n18877), .ZN(n12095) );
  NOR2_X1 U12224 ( .A1(n15943), .A2(n15944), .ZN(n15942) );
  AND2_X1 U12225 ( .A1(n9829), .A2(n9828), .ZN(n15943) );
  INV_X1 U12226 ( .A(n9829), .ZN(n15957) );
  AND2_X1 U12227 ( .A1(n9827), .A2(n9828), .ZN(n15966) );
  NOR2_X1 U12228 ( .A1(n14747), .A2(n18865), .ZN(n12994) );
  INV_X1 U12229 ( .A(n9827), .ZN(n12993) );
  AND2_X1 U12230 ( .A1(n14744), .A2(n16004), .ZN(n14747) );
  NAND2_X1 U12231 ( .A1(n12381), .A2(n12380), .ZN(n12376) );
  NAND2_X1 U12232 ( .A1(n12090), .A2(n12089), .ZN(n18889) );
  NOR2_X1 U12233 ( .A1(n12605), .A2(n13120), .ZN(n19303) );
  OR2_X1 U12234 ( .A1(n10725), .A2(n10724), .ZN(n13702) );
  OR2_X1 U12235 ( .A1(n10708), .A2(n10707), .ZN(n13727) );
  NAND2_X1 U12236 ( .A1(n9942), .A2(n9943), .ZN(n9939) );
  AND2_X1 U12237 ( .A1(n13301), .A2(n9750), .ZN(n9943) );
  INV_X1 U12238 ( .A(n14854), .ZN(n14860) );
  INV_X1 U12239 ( .A(n18968), .ZN(n18945) );
  NOR2_X1 U12240 ( .A1(n18945), .A2(n18964), .ZN(n18951) );
  NAND2_X1 U12241 ( .A1(n9946), .A2(n12613), .ZN(n13305) );
  INV_X1 U12242 ( .A(n18937), .ZN(n18972) );
  INV_X2 U12243 ( .A(n18978), .ZN(n19007) );
  INV_X1 U12244 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16058) );
  NAND2_X1 U12245 ( .A1(n18659), .A2(n12478), .ZN(n16059) );
  INV_X1 U12246 ( .A(n16072), .ZN(n19013) );
  AND2_X1 U12247 ( .A1(n15349), .A2(n12556), .ZN(n16086) );
  NOR2_X1 U12248 ( .A1(n16099), .A2(n12567), .ZN(n15349) );
  NOR2_X1 U12249 ( .A1(n13278), .A2(n9907), .ZN(n15395) );
  NAND2_X1 U12250 ( .A1(n9909), .A2(n13565), .ZN(n9907) );
  AOI21_X1 U12251 ( .B1(n9815), .B2(n9813), .A(n9743), .ZN(n9812) );
  INV_X1 U12252 ( .A(n9815), .ZN(n9814) );
  INV_X1 U12253 ( .A(n9816), .ZN(n9813) );
  NAND2_X1 U12254 ( .A1(n13570), .A2(n9816), .ZN(n9811) );
  NOR2_X1 U12255 ( .A1(n13278), .A2(n10517), .ZN(n13561) );
  INV_X1 U12256 ( .A(n12601), .ZN(n13238) );
  AND2_X1 U12257 ( .A1(n15213), .A2(n13281), .ZN(n15367) );
  INV_X1 U12258 ( .A(n15405), .ZN(n16102) );
  INV_X1 U12259 ( .A(n19303), .ZN(n19716) );
  INV_X1 U12260 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19700) );
  OR2_X1 U12261 ( .A1(n13149), .A2(n13148), .ZN(n13150) );
  OR2_X1 U12262 ( .A1(n13220), .A2(n13219), .ZN(n13221) );
  NAND2_X1 U12263 ( .A1(n13708), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19678) );
  INV_X1 U12264 ( .A(n16138), .ZN(n13708) );
  INV_X1 U12265 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13139) );
  OR2_X1 U12266 ( .A1(n19136), .A2(n19338), .ZN(n19154) );
  INV_X1 U12267 ( .A(n19196), .ZN(n19214) );
  AND2_X1 U12268 ( .A1(n19278), .A2(n19684), .ZN(n19213) );
  NAND2_X1 U12269 ( .A1(n13714), .A2(n13713), .ZN(n19264) );
  OR2_X1 U12270 ( .A1(n19274), .A2(n19273), .ZN(n19300) );
  INV_X1 U12271 ( .A(n19361), .ZN(n19362) );
  NOR2_X2 U12272 ( .A1(n19475), .A2(n19337), .ZN(n19392) );
  INV_X1 U12273 ( .A(n19424), .ZN(n19416) );
  INV_X1 U12274 ( .A(n19556), .ZN(n19438) );
  INV_X1 U12275 ( .A(n19562), .ZN(n19442) );
  INV_X1 U12276 ( .A(n19568), .ZN(n19446) );
  INV_X1 U12277 ( .A(n19574), .ZN(n19450) );
  INV_X1 U12278 ( .A(n19586), .ZN(n19456) );
  OAI22_X1 U12279 ( .A1(n19066), .A2(n19065), .B1(n19064), .B2(n19063), .ZN(
        n19462) );
  INV_X1 U12280 ( .A(n19533), .ZN(n19521) );
  INV_X1 U12281 ( .A(n19580), .ZN(n19520) );
  OAI21_X1 U12282 ( .B1(n19508), .B2(n19507), .A(n19506), .ZN(n19529) );
  INV_X1 U12283 ( .A(n19596), .ZN(n19528) );
  AND2_X1 U12284 ( .A1(n13720), .A2(n19067), .ZN(n19551) );
  AND2_X1 U12285 ( .A1(n10234), .A2(n19067), .ZN(n19575) );
  OAI22_X1 U12286 ( .A1(n14375), .A2(n19065), .B1(n19056), .B2(n19063), .ZN(
        n19583) );
  AND2_X1 U12287 ( .A1(n19057), .A2(n19067), .ZN(n19581) );
  NOR2_X2 U12288 ( .A1(n19475), .A2(n19540), .ZN(n19592) );
  INV_X1 U12289 ( .A(n19462), .ZN(n19597) );
  INV_X1 U12290 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n19601) );
  AND2_X1 U12291 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10432), .ZN(n19598) );
  AND2_X1 U12292 ( .A1(n16176), .A2(n16175), .ZN(n19608) );
  AND3_X1 U12293 ( .A1(n20805), .A2(n19662), .A3(n19618), .ZN(n19744) );
  NOR2_X1 U12294 ( .A1(n11036), .A2(n11050), .ZN(n16318) );
  NOR2_X1 U12295 ( .A1(n11041), .A2(n11072), .ZN(n17224) );
  NOR2_X1 U12296 ( .A1(n16401), .A2(n16659), .ZN(n16389) );
  NAND2_X1 U12297 ( .A1(n9901), .A2(n9902), .ZN(n16431) );
  AND2_X1 U12298 ( .A1(n16450), .A2(n9732), .ZN(n16445) );
  NOR2_X1 U12299 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n20822), .ZN(n20821) );
  NAND2_X1 U12300 ( .A1(n16337), .A2(n18474), .ZN(n16691) );
  NOR2_X1 U12301 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16572), .ZN(n16571) );
  INV_X1 U12302 ( .A(n16691), .ZN(n20827) );
  NAND2_X1 U12303 ( .A1(n16336), .A2(n17963), .ZN(n16703) );
  INV_X1 U12304 ( .A(n20834), .ZN(n16700) );
  NOR2_X1 U12305 ( .A1(n16836), .A2(n16851), .ZN(n16821) );
  NAND2_X1 U12306 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n16867), .ZN(n16851) );
  NOR2_X2 U12307 ( .A1(n13949), .A2(n15535), .ZN(n16880) );
  NAND2_X1 U12308 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17028), .ZN(n17024) );
  NOR2_X1 U12309 ( .A1(n17173), .A2(n17033), .ZN(n17028) );
  INV_X1 U12310 ( .A(n17038), .ZN(n17034) );
  NAND2_X1 U12311 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17034), .ZN(n17033) );
  NOR2_X1 U12312 ( .A1(n17092), .A2(n17043), .ZN(n17039) );
  AND2_X1 U12313 ( .A1(n17050), .A2(n17077), .ZN(n17072) );
  NAND2_X1 U12314 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17087), .ZN(n17083) );
  INV_X1 U12315 ( .A(n17075), .ZN(n17082) );
  NOR2_X1 U12316 ( .A1(n17119), .A2(n17093), .ZN(n17095) );
  NOR2_X1 U12317 ( .A1(n10817), .A2(n10816), .ZN(n17130) );
  NOR2_X1 U12318 ( .A1(n10837), .A2(n10836), .ZN(n17143) );
  INV_X1 U12319 ( .A(n10851), .ZN(n10865) );
  INV_X1 U12320 ( .A(n17147), .ZN(n17156) );
  NOR2_X1 U12321 ( .A1(n17164), .A2(n17163), .ZN(n17216) );
  CLKBUF_X1 U12322 ( .A(n17263), .Z(n17266) );
  NOR2_X1 U12323 ( .A1(n17266), .A2(n18631), .ZN(n17267) );
  NOR3_X1 U12324 ( .A1(n17649), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n16185), .ZN(n9767) );
  NAND2_X1 U12325 ( .A1(n17408), .A2(n17396), .ZN(n17386) );
  NAND3_X1 U12326 ( .A1(n17433), .A2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17422) );
  INV_X1 U12327 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17421) );
  INV_X1 U12328 ( .A(n17372), .ZN(n17444) );
  AND3_X1 U12329 ( .A1(n9898), .A2(n9897), .A3(n9899), .ZN(n17461) );
  INV_X1 U12330 ( .A(n16501), .ZN(n9897) );
  NAND2_X1 U12331 ( .A1(n9898), .A2(n9899), .ZN(n17561) );
  NOR2_X1 U12332 ( .A1(n17588), .A2(n17587), .ZN(n17572) );
  NOR2_X1 U12333 ( .A1(n17614), .A2(n17541), .ZN(n17640) );
  INV_X1 U12334 ( .A(n17647), .ZN(n17636) );
  OAI21_X1 U12335 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18625), .A(n16320), 
        .ZN(n17643) );
  OR2_X1 U12336 ( .A1(n16320), .A2(n18631), .ZN(n17647) );
  NAND2_X1 U12337 ( .A1(n9796), .A2(n9793), .ZN(n10937) );
  INV_X1 U12338 ( .A(n10935), .ZN(n9793) );
  NAND2_X1 U12339 ( .A1(n9796), .A2(n9794), .ZN(n17290) );
  NOR2_X1 U12340 ( .A1(n10935), .A2(n10936), .ZN(n9794) );
  INV_X1 U12341 ( .A(n9796), .ZN(n17301) );
  INV_X1 U12342 ( .A(n17781), .ZN(n17880) );
  INV_X1 U12343 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18646) );
  NAND2_X1 U12344 ( .A1(n18451), .A2(n17831), .ZN(n17781) );
  NOR2_X1 U12345 ( .A1(n9808), .A2(n10925), .ZN(n17545) );
  NAND2_X1 U12346 ( .A1(n9800), .A2(n9960), .ZN(n17571) );
  AND2_X1 U12347 ( .A1(n9800), .A2(n9697), .ZN(n17569) );
  NAND2_X1 U12348 ( .A1(n9965), .A2(n9801), .ZN(n9800) );
  NAND2_X1 U12349 ( .A1(n9965), .A2(n9963), .ZN(n17584) );
  OR2_X1 U12350 ( .A1(n13965), .A2(n11049), .ZN(n18437) );
  NOR2_X1 U12351 ( .A1(n17965), .A2(n17961), .ZN(n17954) );
  INV_X1 U12352 ( .A(n18437), .ZN(n18453) );
  INV_X1 U12353 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18463) );
  INV_X1 U12354 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18467) );
  INV_X1 U12355 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18605) );
  INV_X1 U12356 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18486) );
  INV_X1 U12357 ( .A(n18490), .ZN(n18483) );
  INV_X1 U12358 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18586) );
  AND2_X1 U12360 ( .A1(n12185), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20001)
         );
  NOR2_X1 U12362 ( .A1(n15925), .A2(n9838), .ZN(n15927) );
  AND2_X1 U12363 ( .A1(n12959), .A2(n12958), .ZN(n12960) );
  OAI21_X1 U12364 ( .B1(n14792), .B2(n19020), .A(n14053), .ZN(n14054) );
  OAI211_X1 U12365 ( .C1(n14792), .C2(n15404), .A(n14046), .B(n14045), .ZN(
        n14047) );
  NOR2_X1 U12366 ( .A1(n14044), .A2(n10068), .ZN(n14046) );
  NAND2_X1 U12367 ( .A1(n9916), .A2(n9912), .ZN(n9911) );
  AOI21_X1 U12368 ( .B1(n15102), .B2(n16105), .A(n15101), .ZN(n15103) );
  AOI21_X1 U12369 ( .B1(n9874), .B2(n18487), .A(n9872), .ZN(n16364) );
  NAND2_X1 U12370 ( .A1(n9873), .A2(n9729), .ZN(n9872) );
  AOI21_X1 U12371 ( .B1(n12203), .B2(n17633), .A(n12202), .ZN(n12204) );
  NAND2_X1 U12372 ( .A1(n12201), .A2(n12200), .ZN(n12202) );
  NOR2_X1 U12373 ( .A1(n9968), .A2(n9710), .ZN(n9967) );
  NOR2_X1 U12374 ( .A1(n11145), .A2(n11144), .ZN(n11146) );
  OAI211_X1 U12375 ( .C1(n11121), .C2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11120), .B(n11119), .ZN(n11122) );
  NOR2_X2 U12376 ( .A1(n10810), .A2(n9791), .ZN(n10858) );
  NAND2_X1 U12377 ( .A1(n14307), .A2(n9722), .ZN(n14308) );
  AND2_X1 U12378 ( .A1(n10060), .A2(n9685), .ZN(n9676) );
  NAND3_X1 U12379 ( .A1(n9879), .A2(n9877), .A3(n9876), .ZN(n9732) );
  OAI21_X2 U12380 ( .B1(n11391), .B2(n11390), .A(n11439), .ZN(n13656) );
  INV_X1 U12381 ( .A(n9651), .ZN(n11911) );
  INV_X1 U12382 ( .A(n10853), .ZN(n11016) );
  OR2_X1 U12383 ( .A1(n10127), .A2(n9841), .ZN(n9677) );
  NAND2_X1 U12384 ( .A1(n9956), .A2(n12666), .ZN(n13934) );
  NAND2_X1 U12385 ( .A1(n14285), .A2(n9742), .ZN(n14271) );
  NAND2_X1 U12386 ( .A1(n9676), .A2(n14965), .ZN(n14955) );
  NAND2_X1 U12387 ( .A1(n11930), .A2(n20025), .ZN(n13265) );
  INV_X1 U12388 ( .A(n10122), .ZN(n9837) );
  AND4_X1 U12389 ( .A1(n9837), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9678) );
  AND2_X1 U12390 ( .A1(n12357), .A2(n15300), .ZN(n15285) );
  AND2_X1 U12391 ( .A1(n9833), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9679) );
  NAND2_X1 U12392 ( .A1(n14527), .A2(n12000), .ZN(n14495) );
  AND3_X1 U12393 ( .A1(n9798), .A2(n9797), .A3(n9720), .ZN(n9680) );
  OR2_X1 U12394 ( .A1(n16000), .A2(n10046), .ZN(n14975) );
  AND2_X1 U12395 ( .A1(n14489), .A2(n9757), .ZN(n9681) );
  AND2_X1 U12396 ( .A1(n9819), .A2(n9709), .ZN(n15326) );
  AND2_X1 U12397 ( .A1(n10053), .A2(n10055), .ZN(n15264) );
  NAND2_X1 U12398 ( .A1(n10062), .A2(n10061), .ZN(n16062) );
  AND2_X1 U12399 ( .A1(n12328), .A2(n9731), .ZN(n9682) );
  INV_X1 U12400 ( .A(n10915), .ZN(n9964) );
  AND2_X1 U12401 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n10914), .ZN(
        n10915) );
  XNOR2_X1 U12402 ( .A(n11356), .B(n11354), .ZN(n11398) );
  NOR2_X1 U12403 ( .A1(n10022), .A2(n9592), .ZN(n10020) );
  AND2_X1 U12404 ( .A1(n9679), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9683) );
  NAND2_X1 U12405 ( .A1(n10115), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10114) );
  OR2_X1 U12406 ( .A1(n10127), .A2(n9844), .ZN(n9684) );
  NAND2_X1 U12407 ( .A1(n14036), .A2(n12557), .ZN(n9685) );
  OR2_X1 U12408 ( .A1(n13308), .A2(n13307), .ZN(n13306) );
  AND2_X1 U12409 ( .A1(n9831), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9686) );
  AND2_X1 U12410 ( .A1(n12666), .A2(n9955), .ZN(n9687) );
  AND2_X1 U12411 ( .A1(n9903), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9688) );
  AND2_X1 U12412 ( .A1(n11397), .A2(n11415), .ZN(n9689) );
  NAND2_X1 U12413 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n9690) );
  AND2_X1 U12414 ( .A1(n9857), .A2(n14127), .ZN(n9691) );
  INV_X1 U12415 ( .A(n17588), .ZN(n9898) );
  OR2_X1 U12416 ( .A1(n12359), .A2(n12358), .ZN(n9692) );
  NOR2_X1 U12417 ( .A1(n10810), .A2(n10807), .ZN(n10888) );
  NAND2_X1 U12418 ( .A1(n14490), .A2(n14489), .ZN(n14475) );
  OR3_X1 U12419 ( .A1(n14812), .A2(n9990), .A3(n9991), .ZN(n9693) );
  AND2_X1 U12420 ( .A1(n10927), .A2(n10926), .ZN(n9696) );
  AND2_X1 U12421 ( .A1(n9960), .A2(n9799), .ZN(n9697) );
  OR2_X1 U12422 ( .A1(n14175), .A2(n10040), .ZN(n9698) );
  NAND2_X1 U12423 ( .A1(n10053), .A2(n10051), .ZN(n12966) );
  NOR2_X1 U12424 ( .A1(n10120), .A2(n15076), .ZN(n10121) );
  AND2_X1 U12425 ( .A1(n10121), .A2(n9833), .ZN(n10119) );
  AND2_X1 U12426 ( .A1(n10786), .A2(n10007), .ZN(n9700) );
  AND2_X1 U12427 ( .A1(n9657), .A2(n12732), .ZN(n9701) );
  NOR2_X1 U12428 ( .A1(n14479), .A2(n11999), .ZN(n9702) );
  AND2_X1 U12429 ( .A1(n9984), .A2(n13736), .ZN(n9703) );
  AND2_X1 U12430 ( .A1(n14285), .A2(n14286), .ZN(n14275) );
  AND2_X1 U12431 ( .A1(n13332), .A2(n16115), .ZN(n9704) );
  AND2_X1 U12432 ( .A1(n14256), .A2(n14257), .ZN(n14249) );
  NAND2_X1 U12433 ( .A1(n14256), .A2(n10027), .ZN(n14248) );
  AND3_X1 U12434 ( .A1(n10220), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10219), .ZN(n9705) );
  AND4_X1 U12435 ( .A1(n10268), .A2(n10258), .A3(n10256), .A4(n12515), .ZN(
        n9706) );
  AND2_X1 U12436 ( .A1(n9704), .A2(n12232), .ZN(n12281) );
  NOR2_X1 U12437 ( .A1(n11236), .A2(n20025), .ZN(n11279) );
  NAND2_X1 U12438 ( .A1(n9819), .A2(n10063), .ZN(n15342) );
  AND4_X1 U12439 ( .A1(n11199), .A2(n11196), .A3(n11197), .A4(n11198), .ZN(
        n9707) );
  NOR3_X1 U12440 ( .A1(n14003), .A2(n14002), .A3(n14006), .ZN(n9708) );
  NOR2_X1 U12441 ( .A1(n15343), .A2(n9818), .ZN(n9709) );
  AND2_X1 U12442 ( .A1(n17372), .A2(n9767), .ZN(n9710) );
  NAND2_X1 U12443 ( .A1(n10276), .A2(n10275), .ZN(n10289) );
  AND2_X1 U12444 ( .A1(n10939), .A2(n16191), .ZN(n9712) );
  OR2_X1 U12445 ( .A1(n10278), .A2(n13720), .ZN(n9713) );
  INV_X1 U12446 ( .A(n10258), .ZN(n10270) );
  INV_X1 U12447 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13431) );
  AND2_X1 U12448 ( .A1(n12515), .A2(n19045), .ZN(n9714) );
  NOR2_X1 U12449 ( .A1(n12302), .A2(n12301), .ZN(n12324) );
  INV_X2 U12450 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10299) );
  NAND2_X1 U12451 ( .A1(n9819), .A2(n9817), .ZN(n15306) );
  AND2_X1 U12452 ( .A1(n15800), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9715) );
  OR2_X1 U12453 ( .A1(n14175), .A2(n10042), .ZN(n12126) );
  NOR2_X1 U12454 ( .A1(n16000), .A2(n16001), .ZN(n14987) );
  NAND2_X1 U12455 ( .A1(n14831), .A2(n14821), .ZN(n14809) );
  AND2_X1 U12456 ( .A1(n12846), .A2(n10066), .ZN(n12847) );
  NAND2_X1 U12457 ( .A1(n14825), .A2(n10091), .ZN(n12825) );
  NAND2_X1 U12458 ( .A1(n14256), .A2(n10025), .ZN(n9716) );
  INV_X1 U12459 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20796) );
  INV_X1 U12460 ( .A(n19742), .ZN(n19027) );
  AND2_X1 U12461 ( .A1(n12592), .A2(n13300), .ZN(n13330) );
  INV_X1 U12462 ( .A(n12233), .ZN(n12226) );
  AND2_X1 U12463 ( .A1(n15889), .A2(n13808), .ZN(n9717) );
  AND2_X1 U12464 ( .A1(n9703), .A2(n9983), .ZN(n9718) );
  AND2_X1 U12465 ( .A1(n9938), .A2(n9937), .ZN(n9719) );
  NAND2_X1 U12466 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n10919), .ZN(
        n9720) );
  INV_X1 U12467 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13921) );
  OR2_X1 U12468 ( .A1(n12076), .A2(n12075), .ZN(P1_U2971) );
  NAND2_X1 U12469 ( .A1(n20050), .A2(n11371), .ZN(n13459) );
  NAND2_X1 U12470 ( .A1(n11586), .A2(n11585), .ZN(n9722) );
  NOR2_X1 U12471 ( .A1(n15272), .A2(n10730), .ZN(n12980) );
  AND2_X1 U12472 ( .A1(n9956), .A2(n9687), .ZN(n9723) );
  NOR2_X1 U12473 ( .A1(n9677), .A2(n18709), .ZN(n10115) );
  INV_X1 U12474 ( .A(n11282), .ZN(n12066) );
  NOR2_X1 U12475 ( .A1(n10127), .A2(n16032), .ZN(n10117) );
  NOR2_X1 U12476 ( .A1(n10127), .A2(n9843), .ZN(n10116) );
  AND2_X1 U12477 ( .A1(n10121), .A2(n9683), .ZN(n10118) );
  AND2_X1 U12478 ( .A1(n10115), .A2(n9831), .ZN(n9724) );
  OR2_X1 U12479 ( .A1(n14420), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9725) );
  OAI21_X1 U12480 ( .B1(n13570), .B2(n9814), .A(n9812), .ZN(n13839) );
  NAND2_X1 U12481 ( .A1(n15375), .A2(n12328), .ZN(n15074) );
  AND2_X1 U12482 ( .A1(n9918), .A2(n15351), .ZN(n9726) );
  AND2_X1 U12483 ( .A1(n9869), .A2(n9868), .ZN(n9727) );
  OR2_X1 U12484 ( .A1(n13699), .A2(n12985), .ZN(n9728) );
  OR2_X1 U12485 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16353), .ZN(n9729) );
  INV_X1 U12486 ( .A(n13997), .ZN(n9821) );
  AND2_X1 U12487 ( .A1(n14309), .A2(n14317), .ZN(n9730) );
  NOR2_X1 U12488 ( .A1(n15072), .A2(n10065), .ZN(n9731) );
  NOR2_X1 U12489 ( .A1(n13699), .A2(n9977), .ZN(n10364) );
  AND2_X1 U12491 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n9733) );
  AND2_X1 U12492 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n9734) );
  INV_X1 U12493 ( .A(n9905), .ZN(n9904) );
  NAND2_X1 U12494 ( .A1(n17396), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9905) );
  AND2_X1 U12495 ( .A1(n9811), .A2(n9815), .ZN(n9735) );
  AND2_X1 U12496 ( .A1(n14857), .A2(n14776), .ZN(n14758) );
  AND2_X1 U12497 ( .A1(n9785), .A2(n9784), .ZN(n9736) );
  AND2_X1 U12498 ( .A1(n9902), .A2(n9900), .ZN(n9737) );
  AND2_X1 U12499 ( .A1(n9696), .A2(n10929), .ZN(n9738) );
  AND2_X1 U12500 ( .A1(n9921), .A2(n9920), .ZN(n9739) );
  AND2_X1 U12501 ( .A1(n9887), .A2(n9890), .ZN(n9740) );
  INV_X1 U12502 ( .A(n15285), .ZN(n10055) );
  INV_X1 U12503 ( .A(n9768), .ZN(n17831) );
  OR2_X1 U12504 ( .A1(n18437), .A2(n18449), .ZN(n9768) );
  NAND2_X1 U12505 ( .A1(n9944), .A2(n13301), .ZN(n13303) );
  OAI22_X1 U12506 ( .A1(n14051), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19741), 
        .B2(n10409), .ZN(n13752) );
  INV_X1 U12507 ( .A(n12801), .ZN(n9953) );
  NAND2_X1 U12508 ( .A1(n15361), .A2(n15360), .ZN(n15362) );
  NAND2_X1 U12509 ( .A1(n9906), .A2(n9909), .ZN(n13562) );
  NAND2_X1 U12510 ( .A1(n13769), .A2(n13770), .ZN(n13729) );
  NAND2_X1 U12511 ( .A1(n20114), .A2(n11303), .ZN(n20050) );
  OR2_X1 U12512 ( .A1(n12578), .A2(n12561), .ZN(n15404) );
  INV_X1 U12513 ( .A(n15404), .ZN(n16104) );
  AND2_X1 U12514 ( .A1(n10115), .A2(n9830), .ZN(n10112) );
  INV_X1 U12515 ( .A(n12380), .ZN(n9999) );
  NOR2_X1 U12516 ( .A1(n13308), .A2(n9986), .ZN(n13360) );
  AND2_X1 U12517 ( .A1(n14266), .A2(n9871), .ZN(n9741) );
  AND2_X1 U12518 ( .A1(n13535), .A2(n9718), .ZN(n13769) );
  AND2_X1 U12519 ( .A1(n15361), .A2(n9918), .ZN(n15350) );
  AND2_X1 U12520 ( .A1(n14319), .A2(n14318), .ZN(n14311) );
  AND2_X1 U12521 ( .A1(n14286), .A2(n14276), .ZN(n9742) );
  NAND2_X1 U12522 ( .A1(n10023), .A2(n13760), .ZN(n13570) );
  XOR2_X1 U12523 ( .A(n18862), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n9743) );
  INV_X1 U12524 ( .A(n17600), .ZN(n9965) );
  INV_X1 U12525 ( .A(n12398), .ZN(n10008) );
  OR2_X1 U12526 ( .A1(n17546), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9744) );
  NAND2_X1 U12527 ( .A1(n10924), .A2(n9973), .ZN(n17518) );
  INV_X1 U12528 ( .A(n11305), .ZN(n20114) );
  OAI211_X1 U12529 ( .C1(n10273), .C2(n10272), .A(n13135), .B(n19027), .ZN(
        n12538) );
  INV_X1 U12530 ( .A(n9845), .ZN(n10106) );
  NOR2_X1 U12531 ( .A1(n10109), .A2(n14949), .ZN(n9845) );
  INV_X2 U12532 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20578) );
  NOR2_X1 U12533 ( .A1(n10110), .A2(n14970), .ZN(n10107) );
  AND2_X1 U12534 ( .A1(n9741), .A2(n9870), .ZN(n9745) );
  AND2_X1 U12535 ( .A1(n10241), .A2(n10240), .ZN(n12939) );
  INV_X1 U12536 ( .A(n9891), .ZN(n9890) );
  OAI21_X1 U12537 ( .B1(n16659), .B2(n9893), .A(n9892), .ZN(n9891) );
  INV_X1 U12538 ( .A(n17276), .ZN(n12194) );
  INV_X1 U12539 ( .A(n9882), .ZN(n9881) );
  NAND2_X1 U12540 ( .A1(n9883), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9882) );
  OR2_X1 U12541 ( .A1(n12871), .A2(n14814), .ZN(n9746) );
  INV_X1 U12542 ( .A(n13307), .ZN(n10324) );
  NOR2_X1 U12543 ( .A1(n13308), .A2(n9987), .ZN(n9747) );
  AND2_X1 U12544 ( .A1(n10924), .A2(n9975), .ZN(n9748) );
  NOR2_X1 U12545 ( .A1(n16445), .A2(n17359), .ZN(n9749) );
  AND2_X1 U12546 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9750) );
  AND2_X1 U12547 ( .A1(n9965), .A2(n9964), .ZN(n9751) );
  AND2_X1 U12548 ( .A1(n13535), .A2(n9984), .ZN(n9752) );
  INV_X1 U12549 ( .A(n17306), .ZN(n9893) );
  AND2_X1 U12550 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13432) );
  AND2_X1 U12551 ( .A1(n16350), .A2(n9883), .ZN(n9753) );
  NAND2_X1 U12552 ( .A1(n10231), .A2(n10266), .ZN(n13135) );
  AND2_X1 U12553 ( .A1(n14000), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9754) );
  OR2_X1 U12554 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9755) );
  INV_X1 U12555 ( .A(n13013), .ZN(n9928) );
  INV_X1 U12556 ( .A(n9862), .ZN(n13853) );
  NAND2_X1 U12557 ( .A1(n13556), .A2(n9863), .ZN(n9862) );
  INV_X1 U12558 ( .A(n19942), .ZN(n20003) );
  AND2_X1 U12559 ( .A1(n11929), .A2(n20657), .ZN(n19942) );
  NAND2_X1 U12560 ( .A1(n17604), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17588) );
  AND2_X1 U12561 ( .A1(n17408), .A2(n9904), .ZN(n9756) );
  AND2_X1 U12562 ( .A1(n12011), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9757) );
  INV_X1 U12563 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n9880) );
  INV_X1 U12564 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n10001) );
  INV_X1 U12565 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9884) );
  AOI21_X1 U12566 ( .B1(n12079), .B2(n12078), .A(n19606), .ZN(n12080) );
  AOI22_X2 U12567 ( .A1(DATAI_23_), .A2(n20041), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n20040), .ZN(n20512) );
  AOI22_X2 U12568 ( .A1(DATAI_18_), .A2(n20041), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n20040), .ZN(n20488) );
  INV_X1 U12569 ( .A(n12475), .ZN(n9760) );
  NAND2_X1 U12570 ( .A1(n10253), .A2(n10252), .ZN(n10281) );
  NAND3_X1 U12571 ( .A1(n9647), .A2(n10253), .A3(n10252), .ZN(n10297) );
  NAND2_X1 U12572 ( .A1(n9932), .A2(n10280), .ZN(n10282) );
  OAI21_X1 U12573 ( .B1(n9761), .B2(n13917), .A(n13916), .ZN(n15412) );
  INV_X2 U12574 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18590) );
  NAND4_X2 U12575 ( .A1(n10996), .A2(n9769), .A3(n10994), .A4(n10995), .ZN(
        n17092) );
  NAND3_X1 U12576 ( .A1(n9771), .A2(n10993), .A3(n10998), .ZN(n9770) );
  NAND3_X1 U12577 ( .A1(n10078), .A2(n12012), .A3(n14476), .ZN(n9773) );
  OAI21_X2 U12578 ( .B1(n15805), .B2(n9776), .A(n9774), .ZN(n15796) );
  NAND2_X1 U12579 ( .A1(n11956), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9777) );
  NAND2_X1 U12580 ( .A1(n13528), .A2(n9777), .ZN(n19927) );
  NAND2_X1 U12581 ( .A1(n14018), .A2(n14019), .ZN(n14418) );
  AND2_X2 U12582 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13430) );
  NAND2_X1 U12583 ( .A1(n9851), .A2(n9852), .ZN(n9783) );
  INV_X1 U12584 ( .A(n9791), .ZN(n9790) );
  NOR2_X1 U12585 ( .A1(n16692), .A2(n9791), .ZN(n10877) );
  NAND2_X1 U12586 ( .A1(n17425), .A2(n17546), .ZN(n17349) );
  NOR2_X1 U12587 ( .A1(n17620), .A2(n10908), .ZN(n10911) );
  NAND2_X1 U12588 ( .A1(n9805), .A2(n10908), .ZN(n9804) );
  INV_X1 U12589 ( .A(n10910), .ZN(n9805) );
  NAND2_X1 U12590 ( .A1(n10910), .A2(n9807), .ZN(n9806) );
  INV_X1 U12591 ( .A(n10908), .ZN(n9807) );
  NAND2_X1 U12592 ( .A1(n17478), .A2(n17755), .ZN(n10928) );
  INV_X1 U12593 ( .A(n13332), .ZN(n12208) );
  AND2_X1 U12594 ( .A1(n13332), .A2(n13222), .ZN(n12237) );
  NAND2_X1 U12595 ( .A1(n13332), .A2(n12600), .ZN(n12589) );
  XNOR2_X1 U12596 ( .A(n9809), .B(n12207), .ZN(n12593) );
  NAND3_X1 U12597 ( .A1(n9837), .A2(n9835), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10120) );
  NAND3_X1 U12598 ( .A1(n9837), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10123) );
  NOR2_X1 U12599 ( .A1(n15932), .A2(n15933), .ZN(n15931) );
  OAI211_X1 U12600 ( .C1(n9848), .C2(n11439), .A(n9847), .B(n9846), .ZN(n11957) );
  NAND2_X1 U12601 ( .A1(n11439), .A2(n11478), .ZN(n9847) );
  NAND2_X1 U12602 ( .A1(n11438), .A2(n9849), .ZN(n9848) );
  NAND4_X1 U12603 ( .A1(n12007), .A2(n14527), .A3(n12000), .A4(n9590), .ZN(
        n9851) );
  NAND3_X1 U12604 ( .A1(n20050), .A2(n11371), .A3(n20578), .ZN(n10021) );
  NAND2_X1 U12605 ( .A1(n9855), .A2(n9854), .ZN(n13349) );
  NAND2_X1 U12606 ( .A1(n14179), .A2(n9857), .ZN(n9861) );
  NAND2_X1 U12607 ( .A1(n9861), .A2(n14128), .ZN(n9856) );
  NAND2_X1 U12608 ( .A1(n9856), .A2(n9860), .ZN(n9859) );
  NAND2_X1 U12609 ( .A1(n14179), .A2(n14163), .ZN(n14117) );
  INV_X1 U12610 ( .A(n9861), .ZN(n14159) );
  NAND3_X1 U12611 ( .A1(n13556), .A2(n9863), .A3(n13852), .ZN(n15858) );
  NOR2_X1 U12612 ( .A1(n16365), .A2(n16659), .ZN(n16359) );
  INV_X1 U12613 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n9885) );
  NAND2_X1 U12614 ( .A1(n9886), .A2(n9888), .ZN(n16381) );
  NAND2_X1 U12615 ( .A1(n16402), .A2(n9732), .ZN(n9886) );
  NAND2_X1 U12616 ( .A1(n14764), .A2(n9929), .ZN(n14896) );
  NAND2_X1 U12617 ( .A1(n10289), .A2(n9933), .ZN(n9932) );
  INV_X1 U12618 ( .A(n12847), .ZN(n9937) );
  OR2_X2 U12619 ( .A1(n14815), .A2(n14814), .ZN(n9938) );
  INV_X1 U12620 ( .A(n9938), .ZN(n14813) );
  XNOR2_X1 U12621 ( .A(n12846), .B(n10066), .ZN(n14815) );
  NAND3_X1 U12622 ( .A1(n13330), .A2(n9943), .A3(n13331), .ZN(n9940) );
  NAND2_X1 U12623 ( .A1(n9657), .A2(n9951), .ZN(n9947) );
  NAND3_X1 U12624 ( .A1(n9950), .A2(n9952), .A3(n9947), .ZN(n14838) );
  NOR2_X1 U12625 ( .A1(n12801), .A2(n14842), .ZN(n9951) );
  NAND2_X1 U12626 ( .A1(n12801), .A2(n14842), .ZN(n9952) );
  INV_X1 U12627 ( .A(n12775), .ZN(n14836) );
  NOR2_X2 U12628 ( .A1(n13869), .A2(n9954), .ZN(n14846) );
  NAND2_X1 U12629 ( .A1(n9696), .A2(n9957), .ZN(n17425) );
  INV_X1 U12630 ( .A(n17585), .ZN(n9966) );
  NAND2_X1 U12631 ( .A1(n9970), .A2(n9967), .ZN(P3_U2800) );
  AOI21_X1 U12632 ( .B1(n16192), .B2(n16206), .A(n16191), .ZN(n9969) );
  NAND2_X1 U12633 ( .A1(n16190), .A2(n17537), .ZN(n9970) );
  NAND2_X1 U12634 ( .A1(n10924), .A2(n17881), .ZN(n10923) );
  INV_X2 U12635 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11052) );
  INV_X1 U12636 ( .A(n13366), .ZN(n9989) );
  NOR3_X1 U12637 ( .A1(n14812), .A2(n13009), .A3(n9993), .ZN(n14025) );
  NOR2_X1 U12638 ( .A1(n14812), .A2(n13009), .ZN(n13008) );
  INV_X1 U12639 ( .A(n12477), .ZN(n9993) );
  NAND2_X1 U12640 ( .A1(n10767), .A2(n19045), .ZN(n10269) );
  NAND2_X1 U12641 ( .A1(n12337), .A2(n10000), .ZN(n10778) );
  INV_X1 U12642 ( .A(n10778), .ZN(n12354) );
  NAND2_X1 U12643 ( .A1(n10786), .A2(n12398), .ZN(n12401) );
  INV_X1 U12644 ( .A(n14019), .ZN(n10010) );
  NAND2_X1 U12645 ( .A1(n10010), .A2(n10011), .ZN(n10009) );
  NAND2_X1 U12646 ( .A1(n13459), .A2(n10020), .ZN(n10017) );
  INV_X1 U12647 ( .A(n11318), .ZN(n10022) );
  OR2_X1 U12648 ( .A1(n13573), .A2(n14000), .ZN(n10023) );
  XNOR2_X1 U12649 ( .A(n12273), .B(n12274), .ZN(n13573) );
  NAND2_X1 U12650 ( .A1(n14256), .A2(n10024), .ZN(n14200) );
  INV_X1 U12651 ( .A(n14947), .ZN(n10033) );
  NAND2_X1 U12652 ( .A1(n10033), .A2(n10035), .ZN(n14039) );
  NOR2_X1 U12653 ( .A1(n10037), .A2(n10036), .ZN(n10035) );
  NOR2_X1 U12654 ( .A1(n14175), .A2(n10039), .ZN(n14152) );
  NOR2_X1 U12655 ( .A1(n14175), .A2(n14176), .ZN(n11927) );
  NAND3_X1 U12656 ( .A1(n10047), .A2(n13529), .A3(n13530), .ZN(n13546) );
  INV_X1 U12657 ( .A(n13549), .ZN(n10047) );
  AOI21_X1 U12658 ( .B1(n11957), .B2(n11625), .A(n11476), .ZN(n13549) );
  INV_X1 U12659 ( .A(n13546), .ZN(n11500) );
  NAND2_X1 U12660 ( .A1(n13529), .A2(n13530), .ZN(n13548) );
  NAND2_X1 U12661 ( .A1(n13657), .A2(n11625), .ZN(n11402) );
  XNOR2_X1 U12662 ( .A(n11934), .B(n11398), .ZN(n13657) );
  NAND2_X1 U12663 ( .A1(n14996), .A2(n14998), .ZN(n10053) );
  NAND2_X1 U12664 ( .A1(n10053), .A2(n10049), .ZN(n10054) );
  AND2_X1 U12665 ( .A1(n20025), .A2(n20042), .ZN(n20542) );
  OAI21_X1 U12666 ( .B1(n13656), .B2(n11660), .A(n11396), .ZN(n11397) );
  NAND2_X1 U12667 ( .A1(n13264), .A2(n13263), .ZN(n13340) );
  NAND2_X1 U12668 ( .A1(n11234), .A2(n11233), .ZN(n11238) );
  INV_X1 U12669 ( .A(n11526), .ZN(n11517) );
  AND2_X1 U12670 ( .A1(n12231), .A2(n12230), .ZN(n12240) );
  AOI22_X1 U12671 ( .A1(n10226), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12892), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10227) );
  AOI22_X1 U12672 ( .A1(n10226), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12892), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10219) );
  AOI22_X1 U12673 ( .A1(n10226), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12892), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10177) );
  AOI22_X1 U12674 ( .A1(n10226), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12892), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10153) );
  NAND2_X1 U12675 ( .A1(n10257), .A2(n10263), .ZN(n12517) );
  AOI21_X1 U12676 ( .B1(n14132), .B2(n19942), .A(n14022), .ZN(n14023) );
  NAND2_X1 U12677 ( .A1(n14132), .A2(n12175), .ZN(n12190) );
  AOI22_X1 U12678 ( .A1(n10226), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10132) );
  NAND2_X1 U12679 ( .A1(n19858), .A2(n13236), .ZN(n14329) );
  AND2_X1 U12680 ( .A1(n12845), .A2(n12869), .ZN(n10066) );
  INV_X1 U12681 ( .A(n10889), .ZN(n15488) );
  INV_X1 U12682 ( .A(n10842), .ZN(n16950) );
  OR2_X1 U12684 ( .A1(n15744), .A2(n13311), .ZN(n14404) );
  OR2_X1 U12685 ( .A1(n15930), .A2(n15404), .ZN(n10067) );
  AND3_X1 U12686 ( .A1(n15082), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16078), .ZN(n10068) );
  NOR2_X1 U12687 ( .A1(n14785), .A2(n14928), .ZN(n10069) );
  OR2_X1 U12688 ( .A1(n17546), .A2(n20801), .ZN(n10070) );
  AND4_X1 U12689 ( .A1(n10894), .A2(n10893), .A3(n10892), .A4(n10891), .ZN(
        n10071) );
  BUF_X4 U12690 ( .A(n10867), .Z(n15523) );
  BUF_X4 U12691 ( .A(n10852), .Z(n16944) );
  OR2_X1 U12692 ( .A1(n10089), .A2(n13670), .ZN(n10072) );
  AND2_X1 U12693 ( .A1(n10222), .A2(n10221), .ZN(n10073) );
  AND2_X1 U12694 ( .A1(n13917), .A2(n12468), .ZN(n10074) );
  AND4_X1 U12695 ( .A1(n12287), .A2(n12286), .A3(n12285), .A4(n12284), .ZN(
        n10075) );
  OR2_X1 U12696 ( .A1(n14130), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10076) );
  AND4_X1 U12697 ( .A1(n11223), .A2(n11222), .A3(n11221), .A4(n11220), .ZN(
        n10077) );
  AND2_X1 U12698 ( .A1(n14662), .A2(n15820), .ZN(n10078) );
  AND2_X1 U12699 ( .A1(n12265), .A2(n12262), .ZN(n10079) );
  NAND2_X1 U12700 ( .A1(n9701), .A2(n9953), .ZN(n10080) );
  INV_X1 U12701 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10936) );
  INV_X1 U12702 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12013) );
  INV_X1 U12703 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10906) );
  OR3_X1 U12704 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17363), .ZN(n10081) );
  AND2_X1 U12705 ( .A1(n10207), .A2(n10206), .ZN(n10082) );
  OR2_X1 U12706 ( .A1(n14130), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10083) );
  AND2_X1 U12707 ( .A1(n17431), .A2(n17653), .ZN(n10084) );
  AND3_X1 U12708 ( .A1(n10225), .A2(n10136), .A3(n10224), .ZN(n10085) );
  AND2_X1 U12709 ( .A1(n18909), .A2(n18921), .ZN(n10086) );
  AND3_X1 U12710 ( .A1(n10214), .A2(n10136), .A3(n10213), .ZN(n10087) );
  AND2_X1 U12711 ( .A1(n10212), .A2(n10211), .ZN(n10088) );
  INV_X2 U12712 ( .A(n17431), .ZN(n17546) );
  INV_X1 U12713 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19780) );
  OR2_X1 U12714 ( .A1(n11421), .A2(n11350), .ZN(n11318) );
  OR2_X1 U12715 ( .A1(n12618), .A2(n13738), .ZN(n10089) );
  INV_X2 U12716 ( .A(n10090), .ZN(n16962) );
  NOR2_X1 U12717 ( .A1(n17644), .A2(n17614), .ZN(n17342) );
  OR3_X1 U12718 ( .A1(n12801), .A2(n12800), .A3(n14830), .ZN(n10091) );
  AND2_X1 U12719 ( .A1(n15327), .A2(n15324), .ZN(n10093) );
  NAND2_X1 U12720 ( .A1(n12237), .A2(n12233), .ZN(n12306) );
  AND4_X1 U12721 ( .A1(n12295), .A2(n12294), .A3(n12293), .A4(n12292), .ZN(
        n10094) );
  AND3_X1 U12722 ( .A1(n11250), .A2(n11249), .A3(n11248), .ZN(n10095) );
  AND4_X1 U12723 ( .A1(n11230), .A2(n11229), .A3(n11228), .A4(n11227), .ZN(
        n10096) );
  AND4_X1 U12724 ( .A1(n11205), .A2(n11204), .A3(n11203), .A4(n11202), .ZN(
        n10097) );
  AND3_X1 U12725 ( .A1(n11188), .A2(n11187), .A3(n11186), .ZN(n10098) );
  NAND2_X1 U12726 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10248) );
  AOI22_X1 U12727 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n12030), .B1(n12034), 
        .B2(n11930), .ZN(n12045) );
  INV_X1 U12728 ( .A(n11293), .ZN(n11231) );
  INV_X1 U12729 ( .A(n11935), .ZN(n11350) );
  AND3_X1 U12730 ( .A1(n10270), .A2(n10268), .A3(n10271), .ZN(n10193) );
  NOR2_X1 U12731 ( .A1(n10325), .A2(n10247), .ZN(n10251) );
  AOI22_X1 U12732 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19368), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12249) );
  AND2_X1 U12733 ( .A1(n10193), .A2(n10269), .ZN(n10218) );
  AND2_X1 U12734 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10139) );
  AOI22_X1 U12735 ( .A1(n10226), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12892), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10171) );
  NAND2_X1 U12736 ( .A1(n12020), .A2(n12019), .ZN(n12029) );
  INV_X1 U12737 ( .A(n15757), .ZN(n12007) );
  OR2_X1 U12738 ( .A1(n11491), .A2(n11490), .ZN(n11976) );
  OR2_X1 U12739 ( .A1(n11317), .A2(n11316), .ZN(n11935) );
  INV_X1 U12740 ( .A(n12172), .ZN(n11268) );
  INV_X1 U12741 ( .A(n12228), .ZN(n12218) );
  INV_X1 U12742 ( .A(n12161), .ZN(n12168) );
  INV_X1 U12743 ( .A(n14242), .ZN(n11840) );
  INV_X1 U12744 ( .A(n13791), .ZN(n11522) );
  OR2_X1 U12745 ( .A1(n11516), .A2(n11515), .ZN(n11984) );
  INV_X1 U12746 ( .A(n11275), .ZN(n13189) );
  NAND2_X1 U12747 ( .A1(n10417), .A2(n10416), .ZN(n10429) );
  INV_X1 U12748 ( .A(n12826), .ZN(n12827) );
  NOR2_X1 U12749 ( .A1(n10581), .A2(n10580), .ZN(n12321) );
  NAND3_X1 U12750 ( .A1(n10142), .A2(n10141), .A3(n10140), .ZN(n10143) );
  NOR2_X1 U12751 ( .A1(n11077), .A2(n11058), .ZN(n11051) );
  OR2_X1 U12752 ( .A1(n12102), .A2(n14165), .ZN(n12104) );
  NOR2_X1 U12753 ( .A1(n11267), .A2(n20581), .ZN(n11447) );
  AOI21_X1 U12754 ( .B1(n20406), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12024), .ZN(n12023) );
  INV_X1 U12755 ( .A(n13646), .ZN(n15553) );
  NAND2_X1 U12756 ( .A1(n10790), .A2(n12421), .ZN(n12420) );
  NAND2_X1 U12757 ( .A1(n10310), .A2(n10309), .ZN(n10318) );
  AND2_X1 U12758 ( .A1(n13702), .A2(n13700), .ZN(n12620) );
  INV_X1 U12759 ( .A(n12869), .ZN(n12616) );
  INV_X1 U12760 ( .A(n12926), .ZN(n12915) );
  INV_X1 U12761 ( .A(n14827), .ZN(n12798) );
  NOR2_X1 U12762 ( .A1(n10565), .A2(n10564), .ZN(n12296) );
  INV_X1 U12763 ( .A(n12461), .ZN(n12468) );
  NAND2_X1 U12764 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18272), .ZN(
        n11058) );
  NOR2_X1 U12765 ( .A1(n17557), .A2(n17558), .ZN(n11104) );
  NAND2_X1 U12766 ( .A1(n17431), .A2(n17786), .ZN(n10926) );
  INV_X1 U12767 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n20770) );
  INV_X1 U12768 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10917) );
  INV_X1 U12769 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16949) );
  INV_X1 U12770 ( .A(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n20846) );
  AND2_X1 U12771 ( .A1(n11665), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11685) );
  NAND2_X1 U12772 ( .A1(n12170), .A2(n12169), .ZN(n13450) );
  AOI21_X1 U12773 ( .B1(n12153), .B2(n12152), .A(n12151), .ZN(n14058) );
  NAND2_X1 U12774 ( .A1(n13983), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12123) );
  AND2_X1 U12775 ( .A1(n20581), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12154) );
  INV_X1 U12776 ( .A(n11660), .ZN(n11625) );
  INV_X1 U12777 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20327) );
  INV_X1 U12778 ( .A(n10797), .ZN(n10798) );
  NAND2_X1 U12779 ( .A1(n9719), .A2(n12871), .ZN(n12872) );
  AND2_X1 U12780 ( .A1(n12521), .A2(n13137), .ZN(n12938) );
  NOR2_X1 U12781 ( .A1(n15936), .A2(n14002), .ZN(n13993) );
  AND2_X1 U12782 ( .A1(n16086), .A2(n12572), .ZN(n12574) );
  AND2_X1 U12783 ( .A1(n12382), .A2(n12973), .ZN(n15002) );
  OR2_X1 U12784 ( .A1(n18753), .A2(n14002), .ZN(n12390) );
  BUF_X1 U12785 ( .A(n12280), .Z(n19133) );
  AOI22_X1 U12786 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n18457), .B2(n18604), .ZN(
        n11077) );
  NAND2_X1 U12787 ( .A1(n11035), .A2(n11034), .ZN(n13947) );
  INV_X2 U12788 ( .A(n11016), .ZN(n16926) );
  INV_X1 U12789 ( .A(n17130), .ZN(n11100) );
  INV_X1 U12790 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10903) );
  INV_X1 U12791 ( .A(n18427), .ZN(n18449) );
  NAND2_X1 U12792 ( .A1(n11884), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12102) );
  AND2_X1 U12793 ( .A1(n14205), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14194) );
  INV_X1 U12794 ( .A(n19806), .ZN(n15659) );
  AND2_X1 U12795 ( .A1(n20005), .A2(n13597), .ZN(n13603) );
  NAND2_X1 U12796 ( .A1(n13604), .A2(n13603), .ZN(n19820) );
  NAND2_X1 U12797 ( .A1(n13551), .A2(n14089), .ZN(n14130) );
  OR2_X1 U12798 ( .A1(n15744), .A2(n13313), .ZN(n14389) );
  OR2_X1 U12799 ( .A1(n13987), .A2(n13246), .ZN(n13248) );
  INV_X1 U12800 ( .A(n14058), .ZN(n14059) );
  OAI21_X1 U12801 ( .B1(n11471), .B2(n14452), .A(n11862), .ZN(n14201) );
  NAND2_X1 U12802 ( .A1(n13186), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11660) );
  NOR2_X1 U12803 ( .A1(n11565), .A2(n19780), .ZN(n11583) );
  NAND2_X1 U12804 ( .A1(n19944), .A2(n12068), .ZN(n19938) );
  AND2_X1 U12805 ( .A1(n19990), .A2(n14704), .ZN(n15869) );
  INV_X1 U12806 ( .A(n20548), .ZN(n20355) );
  AND2_X1 U12807 ( .A1(n20160), .A2(n20466), .ZN(n20335) );
  NAND2_X1 U12808 ( .A1(n11477), .A2(n11440), .ZN(n20004) );
  INV_X1 U12809 ( .A(n13929), .ZN(n10358) );
  AND2_X1 U12810 ( .A1(n10656), .A2(n10655), .ZN(n13738) );
  INV_X1 U12811 ( .A(n14825), .ZN(n14826) );
  NAND2_X1 U12812 ( .A1(n18953), .A2(n12954), .ZN(n14930) );
  OAI21_X1 U12813 ( .B1(n12952), .B2(n12951), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13052) );
  INV_X1 U12814 ( .A(n19011), .ZN(n18831) );
  INV_X1 U12815 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14006) );
  INV_X1 U12816 ( .A(n12574), .ZN(n15131) );
  OR2_X1 U12817 ( .A1(n12578), .A2(n12550), .ZN(n15213) );
  NOR2_X1 U12818 ( .A1(n19678), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13710) );
  OR2_X1 U12819 ( .A1(n19081), .A2(n19076), .ZN(n19122) );
  INV_X1 U12820 ( .A(n19305), .ZN(n19337) );
  OR2_X1 U12821 ( .A1(n19696), .A2(n19026), .ZN(n19540) );
  INV_X1 U12822 ( .A(n11049), .ZN(n13964) );
  NOR2_X1 U12823 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16487), .ZN(n16477) );
  NOR2_X1 U12824 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16536), .ZN(n16520) );
  NOR2_X1 U12825 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16609), .ZN(n16584) );
  NOR2_X1 U12826 ( .A1(n10863), .A2(n10862), .ZN(n10864) );
  OR3_X2 U12827 ( .A1(n10849), .A2(n10848), .A3(n10847), .ZN(n10905) );
  NOR2_X1 U12828 ( .A1(n17712), .A2(n17336), .ZN(n17690) );
  OR2_X1 U12829 ( .A1(n11118), .A2(n16191), .ZN(n11120) );
  NOR2_X1 U12830 ( .A1(n17678), .A2(n17324), .ZN(n17323) );
  INV_X1 U12831 ( .A(n17816), .ZN(n17885) );
  NAND2_X1 U12832 ( .A1(n11103), .A2(n17573), .ZN(n17558) );
  NOR2_X1 U12833 ( .A1(n11084), .A2(n15595), .ZN(n11092) );
  AOI211_X1 U12834 ( .C1(n16929), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n10957), .B(n10956), .ZN(n10958) );
  INV_X1 U12835 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18478) );
  OR3_X1 U12836 ( .A1(n15580), .A2(n19756), .A3(n13180), .ZN(n20678) );
  AND2_X1 U12837 ( .A1(n13848), .A2(n13591), .ZN(n19811) );
  INV_X1 U12838 ( .A(n19833), .ZN(n19818) );
  NAND2_X1 U12839 ( .A1(n13848), .A2(n19820), .ZN(n19806) );
  INV_X1 U12840 ( .A(n14329), .ZN(n19853) );
  AND2_X1 U12841 ( .A1(n15577), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13451) );
  NAND2_X1 U12842 ( .A1(n12174), .A2(n13451), .ZN(n15744) );
  INV_X1 U12843 ( .A(n13469), .ZN(n19921) );
  OR2_X1 U12844 ( .A1(n20678), .A2(n13335), .ZN(n19916) );
  AND2_X1 U12845 ( .A1(n11583), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11584) );
  AND2_X1 U12846 ( .A1(n11530), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11550) );
  AND2_X1 U12847 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11442), .ZN(
        n11473) );
  INV_X1 U12848 ( .A(n14557), .ZN(n15874) );
  NOR2_X1 U12849 ( .A1(n15869), .A2(n14534), .ZN(n19969) );
  NOR2_X1 U12850 ( .A1(n20412), .A2(n15580), .ZN(n20649) );
  NOR2_X1 U12851 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15908) );
  OR2_X1 U12852 ( .A1(n13657), .A2(n20658), .ZN(n20152) );
  OAI22_X1 U12853 ( .A1(n20084), .A2(n20083), .B1(n20338), .B2(n20212), .ZN(
        n20107) );
  NAND2_X1 U12854 ( .A1(n20004), .A2(n13656), .ZN(n20118) );
  INV_X1 U12855 ( .A(n20156), .ZN(n20178) );
  NOR2_X1 U12856 ( .A1(n20665), .A2(n20243), .ZN(n20265) );
  INV_X1 U12857 ( .A(n20369), .ZN(n20330) );
  OR2_X1 U12858 ( .A1(n13657), .A2(n20078), .ZN(n20305) );
  OAI22_X1 U12859 ( .A1(n20340), .A2(n20339), .B1(n20338), .B2(n20467), .ZN(
        n20371) );
  OAI22_X1 U12860 ( .A1(n20416), .A2(n20415), .B1(n20466), .B2(n20414), .ZN(
        n20432) );
  OR2_X1 U12861 ( .A1(n20004), .A2(n13658), .ZN(n20380) );
  INV_X1 U12862 ( .A(n20476), .ZN(n20508) );
  AND2_X1 U12863 ( .A1(n20577), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15577) );
  INV_X1 U12864 ( .A(n20627), .ZN(n20639) );
  OAI21_X1 U12865 ( .B1(n14792), .B2(n18871), .A(n10799), .ZN(n10800) );
  INV_X1 U12866 ( .A(n18890), .ZN(n18849) );
  AND2_X1 U12867 ( .A1(n19735), .A2(n10764), .ZN(n18890) );
  INV_X1 U12868 ( .A(n19606), .ZN(n18882) );
  NOR2_X1 U12869 ( .A1(n14025), .A2(n14024), .ZN(n14026) );
  NAND2_X1 U12870 ( .A1(n13121), .A2(n19598), .ZN(n13122) );
  INV_X1 U12871 ( .A(n18954), .ZN(n18964) );
  INV_X1 U12872 ( .A(n19737), .ZN(n19008) );
  INV_X1 U12873 ( .A(n13108), .ZN(n13104) );
  INV_X1 U12874 ( .A(n16059), .ZN(n19012) );
  NAND2_X1 U12875 ( .A1(n10067), .A2(n15100), .ZN(n15101) );
  AND2_X1 U12876 ( .A1(n13279), .A2(n9906), .ZN(n13816) );
  OR2_X1 U12877 ( .A1(n13710), .A2(n13709), .ZN(n19544) );
  NAND2_X1 U12878 ( .A1(n13151), .A2(n13150), .ZN(n19706) );
  OAI21_X1 U12879 ( .B1(n19037), .B2(n19036), .A(n19035), .ZN(n19070) );
  NOR2_X1 U12880 ( .A1(n19337), .A2(n19187), .ZN(n19124) );
  INV_X1 U12881 ( .A(n19130), .ZN(n19153) );
  INV_X1 U12882 ( .A(n19684), .ZN(n19403) );
  INV_X1 U12883 ( .A(n19246), .ZN(n19236) );
  NAND2_X1 U12884 ( .A1(n19304), .A2(n19716), .ZN(n19187) );
  INV_X1 U12885 ( .A(n19336), .ZN(n19328) );
  AND2_X1 U12886 ( .A1(n19696), .A2(n19026), .ZN(n19305) );
  OAI21_X1 U12887 ( .B1(n19375), .B2(n19390), .A(n19544), .ZN(n19393) );
  AND2_X1 U12888 ( .A1(n19696), .A2(n19706), .ZN(n19684) );
  INV_X1 U12889 ( .A(n19550), .ZN(n19499) );
  NOR2_X1 U12890 ( .A1(n19696), .A2(n19706), .ZN(n19476) );
  NOR2_X2 U12891 ( .A1(n13717), .A2(n13716), .ZN(n19061) );
  INV_X1 U12892 ( .A(n15589), .ZN(n19725) );
  INV_X1 U12893 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20805) );
  NOR2_X1 U12894 ( .A1(n18643), .A2(n16646), .ZN(n16337) );
  NOR2_X1 U12895 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16437), .ZN(n16421) );
  NOR2_X1 U12896 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16457), .ZN(n16444) );
  INV_X1 U12897 ( .A(n16703), .ZN(n20825) );
  INV_X1 U12898 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16668) );
  NAND2_X1 U12899 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n16821), .ZN(n16783) );
  NAND2_X1 U12900 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n16880), .ZN(n16879) );
  NAND2_X1 U12901 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16971), .ZN(n16966) );
  AOI21_X1 U12902 ( .B1(n18428), .B2(n13971), .A(n13948), .ZN(n15591) );
  NOR2_X1 U12903 ( .A1(n10981), .A2(n10980), .ZN(n17006) );
  INV_X1 U12904 ( .A(n17149), .ZN(n17142) );
  INV_X1 U12905 ( .A(n17274), .ZN(n17658) );
  INV_X1 U12906 ( .A(n17790), .ZN(n17712) );
  NAND2_X1 U12907 ( .A1(n17755), .A2(n17843), .ZN(n17788) );
  OR2_X1 U12908 ( .A1(n18178), .A2(n18324), .ZN(n18006) );
  NOR2_X1 U12909 ( .A1(n11135), .A2(n17969), .ZN(n11145) );
  INV_X1 U12910 ( .A(n17482), .ZN(n17830) );
  INV_X1 U12911 ( .A(n17891), .ZN(n17872) );
  NOR2_X1 U12912 ( .A1(n17596), .A2(n17595), .ZN(n17594) );
  INV_X1 U12913 ( .A(n17952), .ZN(n17961) );
  INV_X1 U12914 ( .A(n18249), .ZN(n18242) );
  INV_X1 U12915 ( .A(n18317), .ZN(n18319) );
  INV_X1 U12916 ( .A(n18006), .ZN(n18364) );
  INV_X1 U12917 ( .A(U212), .ZN(n16272) );
  INV_X1 U12918 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20468) );
  INV_X1 U12919 ( .A(n19832), .ZN(n19791) );
  INV_X1 U12920 ( .A(n19815), .ZN(n19835) );
  INV_X1 U12921 ( .A(n19811), .ZN(n19795) );
  OR2_X1 U12922 ( .A1(n12072), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n19823) );
  INV_X1 U12923 ( .A(n14563), .ZN(n14231) );
  NAND2_X1 U12924 ( .A1(n13312), .A2(n20001), .ZN(n15751) );
  INV_X1 U12925 ( .A(n13541), .ZN(n13690) );
  INV_X1 U12926 ( .A(n14397), .ZN(n14403) );
  INV_X1 U12927 ( .A(n19867), .ZN(n19886) );
  INV_X1 U12928 ( .A(n19916), .ZN(n13469) );
  INV_X1 U12929 ( .A(n19993), .ZN(n19953) );
  OR2_X1 U12930 ( .A1(n14733), .A2(n14729), .ZN(n15894) );
  INV_X1 U12931 ( .A(n19973), .ZN(n19998) );
  INV_X1 U12932 ( .A(n19999), .ZN(n20664) );
  OR2_X1 U12933 ( .A1(n20118), .A2(n20152), .ZN(n20067) );
  OR2_X1 U12934 ( .A1(n20118), .A2(n20305), .ZN(n20111) );
  OR2_X1 U12935 ( .A1(n20118), .A2(n20375), .ZN(n20156) );
  NAND2_X1 U12936 ( .A1(n20249), .A2(n20405), .ZN(n20206) );
  NAND2_X1 U12937 ( .A1(n20249), .A2(n20437), .ZN(n20241) );
  NAND2_X1 U12938 ( .A1(n20249), .A2(n20464), .ZN(n20264) );
  NAND2_X1 U12939 ( .A1(n20272), .A2(n20405), .ZN(n20325) );
  OR2_X1 U12940 ( .A1(n20380), .A2(n20305), .ZN(n20369) );
  OR2_X1 U12941 ( .A1(n20380), .A2(n20326), .ZN(n20404) );
  OR2_X1 U12942 ( .A1(n20380), .A2(n20375), .ZN(n20436) );
  NAND2_X1 U12943 ( .A1(n20465), .A2(n20437), .ZN(n20476) );
  NAND2_X1 U12944 ( .A1(n20465), .A2(n20464), .ZN(n20575) );
  INV_X2 U12945 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20581) );
  INV_X1 U12946 ( .A(n20648), .ZN(n20583) );
  INV_X1 U12947 ( .A(n20598), .ZN(n20673) );
  NAND2_X1 U12948 ( .A1(n12440), .A2(n12439), .ZN(n18659) );
  INV_X1 U12949 ( .A(n10800), .ZN(n10801) );
  INV_X1 U12950 ( .A(n18876), .ZN(n18888) );
  INV_X1 U12951 ( .A(n18889), .ZN(n18857) );
  INV_X1 U12952 ( .A(n18877), .ZN(n18893) );
  XNOR2_X1 U12953 ( .A(n13330), .B(n13331), .ZN(n19304) );
  INV_X1 U12954 ( .A(n13122), .ZN(n14796) );
  NAND2_X1 U12955 ( .A1(n13218), .A2(n13221), .ZN(n19696) );
  AND2_X1 U12956 ( .A1(n12941), .A2(n19598), .ZN(n18953) );
  NAND2_X1 U12957 ( .A1(n18953), .A2(n12942), .ZN(n18968) );
  OR2_X1 U12958 ( .A1(n18990), .A2(n19008), .ZN(n18978) );
  INV_X1 U12959 ( .A(n18990), .ZN(n19010) );
  NAND2_X1 U12960 ( .A1(n13031), .A2(n10264), .ZN(n13108) );
  INV_X1 U12961 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16046) );
  INV_X1 U12962 ( .A(n19015), .ZN(n16073) );
  INV_X1 U12963 ( .A(n16105), .ZN(n15413) );
  INV_X1 U12964 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19720) );
  INV_X1 U12965 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16155) );
  INV_X1 U12966 ( .A(n19124), .ZN(n19103) );
  NAND2_X1 U12967 ( .A1(n19305), .A2(n19278), .ZN(n19130) );
  OR2_X1 U12968 ( .A1(n19187), .A2(n19403), .ZN(n19186) );
  OR2_X1 U12969 ( .A1(n19187), .A2(n19218), .ZN(n19246) );
  INV_X1 U12970 ( .A(n19247), .ZN(n19267) );
  INV_X1 U12971 ( .A(n19300), .ZN(n19293) );
  NAND2_X1 U12972 ( .A1(n19278), .A2(n19497), .ZN(n19336) );
  NAND2_X1 U12973 ( .A1(n19498), .A2(n19305), .ZN(n19361) );
  INV_X1 U12974 ( .A(n19463), .ZN(n19429) );
  INV_X1 U12975 ( .A(n19583), .ZN(n19459) );
  NAND2_X1 U12976 ( .A1(n19498), .A2(n19476), .ZN(n19496) );
  NAND2_X1 U12977 ( .A1(n19477), .A2(n19476), .ZN(n19533) );
  NAND2_X1 U12978 ( .A1(n19498), .A2(n19497), .ZN(n19596) );
  INV_X1 U12979 ( .A(n19673), .ZN(n19609) );
  AOI21_X1 U12980 ( .B1(n18420), .B2(n18419), .A(n17164), .ZN(n18651) );
  INV_X1 U12981 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17587) );
  INV_X1 U12982 ( .A(n16688), .ZN(n20832) );
  NOR2_X1 U12983 ( .A1(n16754), .A2(n16707), .ZN(n16758) );
  NOR2_X1 U12984 ( .A1(n16854), .A2(n16879), .ZN(n16867) );
  NOR2_X2 U12985 ( .A1(n16997), .A2(n18024), .ZN(n16998) );
  AND2_X1 U12986 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17115), .ZN(n17118) );
  INV_X1 U12987 ( .A(n16208), .ZN(n17126) );
  INV_X1 U12988 ( .A(n17155), .ZN(n17144) );
  OR2_X1 U12989 ( .A1(n18628), .A2(n17216), .ZN(n17218) );
  NAND2_X1 U12990 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17640), .ZN(n17504) );
  AOI22_X1 U12991 ( .A1(n17843), .A2(n17633), .B1(n17552), .B2(n17845), .ZN(
        n17540) );
  INV_X1 U12992 ( .A(n17633), .ZN(n17648) );
  INV_X1 U12993 ( .A(n17954), .ZN(n17925) );
  INV_X1 U12994 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18272) );
  INV_X1 U12995 ( .A(n18583), .ZN(n18495) );
  INV_X1 U12996 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18509) );
  CLKBUF_X1 U12997 ( .A(n18565), .Z(n18571) );
  INV_X1 U12998 ( .A(n16270), .ZN(n16275) );
  NAND2_X1 U12999 ( .A1(n12190), .A2(n12189), .ZN(P1_U2873) );
  OAI21_X1 U13000 ( .B1(n12077), .B2(n12101), .A(n12100), .ZN(P2_U2825) );
  INV_X1 U13001 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16032) );
  INV_X1 U13002 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16018) );
  INV_X1 U13003 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18709) );
  INV_X1 U13004 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18685) );
  INV_X1 U13005 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15019) );
  NAND2_X1 U13006 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n10112), .ZN(
        n10113) );
  INV_X1 U13007 ( .A(n10113), .ZN(n10099) );
  INV_X1 U13008 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14970) );
  INV_X1 U13009 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14949) );
  INV_X1 U13010 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10103) );
  INV_X1 U13011 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14941) );
  XNOR2_X1 U13012 ( .A(n10102), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14008) );
  INV_X1 U13013 ( .A(n14008), .ZN(n12078) );
  INV_X1 U13014 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10100) );
  INV_X2 U13015 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19741) );
  INV_X1 U13016 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10409) );
  AOI21_X1 U13017 ( .B1(n14941), .B2(n10105), .A(n10102), .ZN(n15926) );
  NAND2_X1 U13018 ( .A1(n10106), .A2(n10103), .ZN(n10104) );
  NAND2_X1 U13019 ( .A1(n10105), .A2(n10104), .ZN(n12482) );
  INV_X1 U13020 ( .A(n12482), .ZN(n15933) );
  AOI21_X1 U13021 ( .B1(n14949), .B2(n10109), .A(n9845), .ZN(n14951) );
  OR2_X1 U13022 ( .A1(n10107), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10108) );
  NAND2_X1 U13023 ( .A1(n10109), .A2(n10108), .ZN(n14960) );
  INV_X1 U13024 ( .A(n14960), .ZN(n15944) );
  AOI21_X1 U13025 ( .B1(n14970), .B2(n10110), .A(n10107), .ZN(n15959) );
  OAI21_X1 U13026 ( .B1(n10111), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n10110), .ZN(n14982) );
  INV_X1 U13027 ( .A(n14982), .ZN(n15967) );
  INV_X1 U13028 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14990) );
  AOI21_X1 U13029 ( .B1(n14990), .B2(n10113), .A(n10111), .ZN(n14993) );
  OAI21_X1 U13030 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n10112), .A(
        n10113), .ZN(n16004) );
  AOI21_X1 U13031 ( .B1(n15019), .B2(n10128), .A(n10112), .ZN(n15023) );
  AOI21_X1 U13032 ( .B1(n18685), .B2(n10114), .A(n9724), .ZN(n18684) );
  AOI21_X1 U13033 ( .B1(n18709), .B2(n9677), .A(n10115), .ZN(n18707) );
  AOI21_X1 U13034 ( .B1(n16018), .B2(n9684), .A(n10116), .ZN(n18729) );
  AOI21_X1 U13035 ( .B1(n16032), .B2(n10127), .A(n10117), .ZN(n18756) );
  AOI21_X1 U13036 ( .B1(n16046), .B2(n10126), .A(n10118), .ZN(n18780) );
  AOI21_X1 U13037 ( .B1(n16058), .B2(n10125), .A(n10119), .ZN(n18804) );
  AOI21_X1 U13038 ( .B1(n15076), .B2(n10120), .A(n10121), .ZN(n18821) );
  AOI21_X1 U13039 ( .B1(n13921), .B2(n10123), .A(n9678), .ZN(n18843) );
  AOI21_X1 U13040 ( .B1(n20796), .B2(n10122), .A(n10124), .ZN(n13755) );
  INV_X1 U13041 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13020) );
  INV_X1 U13042 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20759) );
  AOI22_X1 U13043 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13020), .B1(n20759), 
        .B2(n19741), .ZN(n18898) );
  INV_X1 U13044 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13025) );
  AOI22_X1 U13045 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13025), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19741), .ZN(n15422) );
  NOR2_X1 U13046 ( .A1(n18898), .A2(n15422), .ZN(n15421) );
  OAI21_X1 U13047 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n10122), .ZN(n13813) );
  NAND2_X1 U13048 ( .A1(n15421), .A2(n13813), .ZN(n13753) );
  NOR2_X1 U13049 ( .A1(n13755), .A2(n13753), .ZN(n18864) );
  OAI21_X1 U13050 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n10124), .A(
        n10123), .ZN(n19024) );
  NAND2_X1 U13051 ( .A1(n18864), .A2(n19024), .ZN(n18842) );
  NOR2_X1 U13052 ( .A1(n18843), .A2(n18842), .ZN(n18835) );
  OAI21_X1 U13053 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9678), .A(
        n10120), .ZN(n18836) );
  NAND2_X1 U13054 ( .A1(n18835), .A2(n18836), .ZN(n18820) );
  NOR2_X1 U13055 ( .A1(n18821), .A2(n18820), .ZN(n18812) );
  OAI21_X1 U13056 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n10121), .A(
        n10125), .ZN(n18813) );
  NAND2_X1 U13057 ( .A1(n18812), .A2(n18813), .ZN(n18802) );
  NOR2_X1 U13058 ( .A1(n18804), .A2(n18802), .ZN(n18786) );
  OAI21_X1 U13059 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n10119), .A(
        n10126), .ZN(n18788) );
  NAND2_X1 U13060 ( .A1(n18786), .A2(n18788), .ZN(n18781) );
  NOR2_X1 U13061 ( .A1(n18780), .A2(n18781), .ZN(n18779) );
  OAI21_X1 U13062 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n10118), .A(
        n10127), .ZN(n18766) );
  NAND2_X1 U13063 ( .A1(n18779), .A2(n18766), .ZN(n18755) );
  NOR2_X1 U13064 ( .A1(n18756), .A2(n18755), .ZN(n18746) );
  OAI21_X1 U13065 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n10117), .A(
        n9684), .ZN(n18747) );
  NAND2_X1 U13066 ( .A1(n18746), .A2(n18747), .ZN(n18728) );
  NOR2_X1 U13067 ( .A1(n18729), .A2(n18728), .ZN(n18721) );
  OAI21_X1 U13068 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n10116), .A(
        n9677), .ZN(n18722) );
  NAND2_X1 U13069 ( .A1(n18721), .A2(n18722), .ZN(n18705) );
  NOR2_X1 U13070 ( .A1(n18707), .A2(n18705), .ZN(n18694) );
  OAI21_X1 U13071 ( .B1(n10115), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n10114), .ZN(n18695) );
  NAND2_X1 U13072 ( .A1(n18694), .A2(n18695), .ZN(n18682) );
  NOR2_X1 U13073 ( .A1(n18684), .A2(n18682), .ZN(n14784) );
  OAI21_X1 U13074 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n9724), .A(
        n10128), .ZN(n15034) );
  NAND2_X1 U13075 ( .A1(n14784), .A2(n15034), .ZN(n14771) );
  OAI21_X1 U13076 ( .B1(n15023), .B2(n14771), .A(n13752), .ZN(n14744) );
  NOR2_X1 U13077 ( .A1(n15967), .A2(n15966), .ZN(n15965) );
  NOR2_X1 U13078 ( .A1(n18865), .A2(n15942), .ZN(n13006) );
  NOR2_X1 U13079 ( .A1(n14951), .A2(n13006), .ZN(n13005) );
  NOR2_X1 U13080 ( .A1(n18865), .A2(n13005), .ZN(n15932) );
  NOR2_X1 U13081 ( .A1(n18865), .A2(n15925), .ZN(n12079) );
  NOR2_X1 U13082 ( .A1(n12078), .A2(n12079), .ZN(n12077) );
  INV_X1 U13083 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19682) );
  NAND4_X1 U13084 ( .A1(n19741), .A2(n19733), .A3(n19682), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19606) );
  NOR2_X1 U13085 ( .A1(n18865), .A2(n19606), .ZN(n18899) );
  NAND2_X1 U13086 ( .A1(n12077), .A2(n18899), .ZN(n10802) );
  AND2_X4 U13087 ( .A1(n10435), .A2(n19681), .ZN(n12776) );
  AOI22_X1 U13088 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12892), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10133) );
  AND2_X4 U13089 ( .A1(n15435), .A2(n15415), .ZN(n10442) );
  AND2_X4 U13090 ( .A1(n10437), .A2(n10299), .ZN(n10434) );
  AOI22_X1 U13091 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10131) );
  INV_X2 U13092 ( .A(n10135), .ZN(n12812) );
  AOI22_X1 U13093 ( .A1(n12812), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12777), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10130) );
  NAND2_X1 U13094 ( .A1(n10134), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10144) );
  AOI22_X1 U13095 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10138) );
  INV_X2 U13096 ( .A(n10135), .ZN(n10223) );
  AOI22_X1 U13097 ( .A1(n12812), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10137) );
  AOI22_X1 U13098 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12892), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10140) );
  AOI22_X1 U13099 ( .A1(n10226), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12892), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U13100 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10147) );
  AOI22_X1 U13101 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U13102 ( .A1(n12812), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12777), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10145) );
  NAND4_X1 U13103 ( .A1(n10148), .A2(n10147), .A3(n10146), .A4(n10145), .ZN(
        n10149) );
  NAND2_X1 U13104 ( .A1(n10149), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10156) );
  AOI22_X1 U13105 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10151) );
  AOI22_X1 U13106 ( .A1(n12812), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12777), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10150) );
  NAND4_X1 U13107 ( .A1(n10153), .A2(n10152), .A3(n10151), .A4(n10150), .ZN(
        n10154) );
  NAND2_X1 U13108 ( .A1(n10154), .A2(n10136), .ZN(n10155) );
  AOI22_X1 U13109 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10226), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10160) );
  AOI22_X1 U13110 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10159) );
  AOI22_X1 U13111 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12812), .B1(
        n12777), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10158) );
  AOI22_X1 U13112 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12892), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10157) );
  NAND4_X1 U13113 ( .A1(n10160), .A2(n10159), .A3(n10158), .A4(n10157), .ZN(
        n10161) );
  NAND2_X1 U13114 ( .A1(n10161), .A2(n10136), .ZN(n10168) );
  AOI22_X1 U13115 ( .A1(n10226), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12892), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10165) );
  AOI22_X1 U13116 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U13117 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U13118 ( .A1(n12812), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12777), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10162) );
  NAND4_X1 U13119 ( .A1(n10165), .A2(n10164), .A3(n10163), .A4(n10162), .ZN(
        n10166) );
  NAND2_X1 U13120 ( .A1(n10166), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10167) );
  AOI22_X1 U13121 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U13122 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10170) );
  AOI22_X1 U13123 ( .A1(n12812), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10169) );
  NAND4_X1 U13124 ( .A1(n10172), .A2(n10171), .A3(n10170), .A4(n10169), .ZN(
        n10173) );
  NAND2_X1 U13125 ( .A1(n10173), .A2(n10136), .ZN(n10180) );
  AOI22_X1 U13126 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U13127 ( .A1(n12812), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10174) );
  NAND4_X1 U13128 ( .A1(n10177), .A2(n10176), .A3(n10175), .A4(n10174), .ZN(
        n10178) );
  NAND2_X1 U13129 ( .A1(n10178), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10179) );
  NAND2_X2 U13130 ( .A1(n10180), .A2(n10179), .ZN(n10255) );
  AOI22_X1 U13131 ( .A1(n10226), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U13132 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12892), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10183) );
  AOI22_X1 U13133 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10182) );
  AOI22_X1 U13134 ( .A1(n10223), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10181) );
  NAND4_X1 U13135 ( .A1(n10184), .A2(n10183), .A3(n10182), .A4(n10181), .ZN(
        n10185) );
  AOI22_X1 U13136 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10226), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10189) );
  AOI22_X1 U13137 ( .A1(n12892), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10188) );
  AOI22_X1 U13138 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U13139 ( .A1(n10223), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10186) );
  NAND4_X1 U13140 ( .A1(n10189), .A2(n10188), .A3(n10187), .A4(n10186), .ZN(
        n10190) );
  AOI22_X1 U13141 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10226), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10197) );
  AOI22_X1 U13142 ( .A1(n12812), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12777), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U13143 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10195) );
  AOI22_X1 U13144 ( .A1(n12892), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10194) );
  NAND4_X1 U13145 ( .A1(n10197), .A2(n10196), .A3(n10195), .A4(n10194), .ZN(
        n10198) );
  AOI22_X1 U13146 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10202) );
  AOI22_X1 U13147 ( .A1(n10226), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12892), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10201) );
  AOI22_X1 U13148 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10200) );
  AOI22_X1 U13149 ( .A1(n12812), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10199) );
  NAND4_X1 U13150 ( .A1(n10202), .A2(n10201), .A3(n10200), .A4(n10199), .ZN(
        n10203) );
  INV_X1 U13151 ( .A(n19045), .ZN(n12546) );
  NAND2_X1 U13152 ( .A1(n10433), .A2(n12546), .ZN(n10217) );
  AOI22_X1 U13153 ( .A1(n10226), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12892), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10207) );
  AOI22_X1 U13154 ( .A1(n12812), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12777), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10206) );
  AOI22_X1 U13155 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10209) );
  AOI22_X1 U13156 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10208) );
  NAND2_X1 U13157 ( .A1(n10082), .A2(n10210), .ZN(n10216) );
  AOI22_X1 U13158 ( .A1(n10226), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12892), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10212) );
  AOI22_X1 U13159 ( .A1(n12812), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12777), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10211) );
  AOI22_X1 U13160 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10214) );
  AOI22_X1 U13161 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10213) );
  INV_X1 U13162 ( .A(n13137), .ZN(n12496) );
  AOI22_X1 U13163 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10220) );
  AOI22_X1 U13164 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10222) );
  AOI22_X1 U13165 ( .A1(n12812), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12777), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10221) );
  AOI22_X1 U13166 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10225) );
  AOI22_X1 U13167 ( .A1(n12754), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10228) );
  NAND2_X1 U13168 ( .A1(n12560), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10294) );
  NOR2_X1 U13169 ( .A1(n12515), .A2(n19045), .ZN(n10231) );
  INV_X1 U13170 ( .A(n13135), .ZN(n10232) );
  NAND2_X1 U13171 ( .A1(n10232), .A2(n19027), .ZN(n10759) );
  INV_X1 U13172 ( .A(n10233), .ZN(n10235) );
  NAND2_X1 U13173 ( .A1(n12938), .A2(n10236), .ZN(n10237) );
  NAND2_X1 U13174 ( .A1(n10759), .A2(n10237), .ZN(n12559) );
  NAND2_X1 U13175 ( .A1(n12559), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10279) );
  NAND3_X2 U13176 ( .A1(n10294), .A2(n10279), .A3(n9713), .ZN(n10300) );
  INV_X4 U13177 ( .A(n10311), .ZN(n10404) );
  NAND2_X1 U13178 ( .A1(n10404), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10246) );
  INV_X1 U13179 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n10729) );
  INV_X1 U13180 ( .A(n10257), .ZN(n10241) );
  NAND2_X1 U13181 ( .A1(n10405), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10243) );
  NAND2_X1 U13182 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10242) );
  OAI211_X1 U13183 ( .C1(n10729), .C2(n10403), .A(n10243), .B(n10242), .ZN(
        n10244) );
  INV_X1 U13184 ( .A(n10244), .ZN(n10245) );
  NAND2_X1 U13185 ( .A1(n10246), .A2(n10245), .ZN(n13697) );
  INV_X1 U13186 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10247) );
  NAND2_X1 U13187 ( .A1(n10249), .A2(n10248), .ZN(n10250) );
  NOR2_X1 U13188 ( .A1(n10251), .A2(n10250), .ZN(n10253) );
  NAND2_X1 U13189 ( .A1(n10300), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10252) );
  INV_X1 U13190 ( .A(n12939), .ZN(n10254) );
  NAND2_X1 U13191 ( .A1(n10254), .A2(n12546), .ZN(n10262) );
  NAND2_X1 U13192 ( .A1(n10263), .A2(n10270), .ZN(n12514) );
  NAND2_X1 U13193 ( .A1(n12517), .A2(n10259), .ZN(n12523) );
  NAND2_X1 U13194 ( .A1(n12545), .A2(n19045), .ZN(n10261) );
  NAND3_X1 U13195 ( .A1(n10262), .A2(n10261), .A3(n19742), .ZN(n10265) );
  NAND2_X1 U13196 ( .A1(n10263), .A2(n10264), .ZN(n12539) );
  NAND2_X1 U13197 ( .A1(n10265), .A2(n12539), .ZN(n10276) );
  INV_X1 U13198 ( .A(n10412), .ZN(n10267) );
  NAND3_X1 U13199 ( .A1(n12563), .A2(n19742), .A3(n10267), .ZN(n10274) );
  OAI211_X1 U13200 ( .C1(n10268), .C2(n10767), .A(n10269), .B(n12515), .ZN(
        n10273) );
  NOR2_X1 U13201 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19734) );
  NAND2_X1 U13202 ( .A1(n19734), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10277) );
  AND3_X1 U13203 ( .A1(n10279), .A2(n10278), .A3(n10277), .ZN(n10280) );
  NAND2_X1 U13204 ( .A1(n10281), .A2(n10282), .ZN(n10283) );
  NAND2_X1 U13205 ( .A1(n10406), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10286) );
  NAND2_X1 U13206 ( .A1(n9674), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10285) );
  INV_X1 U13207 ( .A(n19734), .ZN(n16171) );
  NAND2_X1 U13208 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10284) );
  INV_X1 U13209 ( .A(n10291), .ZN(n15438) );
  AOI21_X1 U13210 ( .B1(n15438), .B2(n15415), .A(n19741), .ZN(n10292) );
  OAI21_X1 U13211 ( .B1(n10289), .B2(n10290), .A(n10292), .ZN(n10296) );
  NAND2_X1 U13212 ( .A1(n19734), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10293) );
  AND2_X1 U13213 ( .A1(n10294), .A2(n10293), .ZN(n10295) );
  NAND2_X1 U13214 ( .A1(n10296), .A2(n10295), .ZN(n12212) );
  AOI21_X1 U13215 ( .B1(n19741), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10298) );
  OAI21_X2 U13216 ( .B1(n10307), .B2(n10299), .A(n10298), .ZN(n10303) );
  INV_X1 U13217 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n13818) );
  NAND2_X1 U13218 ( .A1(n10300), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10302) );
  AOI22_X1 U13219 ( .A1(n9675), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10301) );
  OAI211_X1 U13220 ( .C1(n10403), .C2(n13818), .A(n10302), .B(n10301), .ZN(
        n10304) );
  NAND2_X1 U13221 ( .A1(n10303), .A2(n10304), .ZN(n10305) );
  INV_X1 U13222 ( .A(n10307), .ZN(n10308) );
  NAND2_X1 U13223 ( .A1(n10308), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10310) );
  NAND2_X1 U13224 ( .A1(n19734), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10309) );
  INV_X1 U13225 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10772) );
  INV_X1 U13226 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n10536) );
  NAND2_X1 U13227 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10312) );
  NAND2_X1 U13228 ( .A1(n10315), .A2(n12206), .ZN(n10320) );
  INV_X1 U13229 ( .A(n10316), .ZN(n10317) );
  OR2_X1 U13230 ( .A1(n10318), .A2(n10317), .ZN(n10319) );
  NAND2_X1 U13231 ( .A1(n10320), .A2(n10319), .ZN(n13308) );
  INV_X1 U13232 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n10551) );
  NAND2_X1 U13233 ( .A1(n10405), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n10322) );
  NAND2_X1 U13234 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10321) );
  OAI211_X1 U13235 ( .C1(n10551), .C2(n10403), .A(n10322), .B(n10321), .ZN(
        n10323) );
  AOI21_X1 U13236 ( .B1(n10404), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n10323), .ZN(n13307) );
  INV_X1 U13237 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n10328) );
  NAND2_X1 U13238 ( .A1(n10405), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n10327) );
  NAND2_X1 U13239 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10326) );
  OAI211_X1 U13240 ( .C1(n10328), .C2(n10403), .A(n10327), .B(n10326), .ZN(
        n10329) );
  AOI21_X1 U13241 ( .B1(n10404), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n10329), .ZN(n13325) );
  INV_X1 U13242 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n10332) );
  NAND2_X1 U13243 ( .A1(n10404), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10331) );
  AOI22_X1 U13244 ( .A1(n10405), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10330) );
  OAI211_X1 U13245 ( .C1(n10403), .C2(n10332), .A(n10331), .B(n10330), .ZN(
        n13366) );
  INV_X1 U13246 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n10335) );
  NAND2_X1 U13247 ( .A1(n10404), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10334) );
  AOI22_X1 U13248 ( .A1(n10405), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10333) );
  OAI211_X1 U13249 ( .C1(n10403), .C2(n10335), .A(n10334), .B(n10333), .ZN(
        n13361) );
  AND2_X2 U13250 ( .A1(n13360), .A2(n13361), .ZN(n13535) );
  INV_X1 U13251 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16091) );
  AOI22_X1 U13252 ( .A1(n10405), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10337) );
  NAND2_X1 U13253 ( .A1(n10406), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10336) );
  OAI211_X1 U13254 ( .C1(n10311), .C2(n16091), .A(n10337), .B(n10336), .ZN(
        n13534) );
  INV_X1 U13255 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n10638) );
  NAND2_X1 U13256 ( .A1(n10405), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10339) );
  NAND2_X1 U13257 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10338) );
  OAI211_X1 U13258 ( .C1(n10638), .C2(n10403), .A(n10339), .B(n10338), .ZN(
        n10340) );
  AOI21_X1 U13259 ( .B1(n10404), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n10340), .ZN(n13675) );
  INV_X1 U13260 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n10659) );
  NAND2_X1 U13261 ( .A1(n10404), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10342) );
  AOI22_X1 U13262 ( .A1(n10405), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10341) );
  OAI211_X1 U13263 ( .C1(n10403), .C2(n10659), .A(n10342), .B(n10341), .ZN(
        n13736) );
  INV_X1 U13264 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n10676) );
  NAND2_X1 U13265 ( .A1(n10405), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10344) );
  NAND2_X1 U13266 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10343) );
  OAI211_X1 U13267 ( .C1(n10676), .C2(n10403), .A(n10344), .B(n10343), .ZN(
        n10345) );
  AOI21_X1 U13268 ( .B1(n10404), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n10345), .ZN(n13780) );
  INV_X1 U13269 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n10693) );
  NAND2_X1 U13270 ( .A1(n10404), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10347) );
  AOI22_X1 U13271 ( .A1(n10405), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n10346) );
  OAI211_X1 U13272 ( .C1(n10325), .C2(n10693), .A(n10347), .B(n10346), .ZN(
        n13770) );
  INV_X1 U13273 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n10711) );
  NAND2_X1 U13274 ( .A1(n10405), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10349) );
  NAND2_X1 U13275 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10348) );
  OAI211_X1 U13276 ( .C1(n10711), .C2(n10403), .A(n10349), .B(n10348), .ZN(
        n10350) );
  AOI21_X1 U13277 ( .B1(n10404), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n10350), .ZN(n13730) );
  NAND2_X1 U13278 ( .A1(n13697), .A2(n13731), .ZN(n13699) );
  INV_X1 U13279 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10353) );
  INV_X1 U13280 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n10456) );
  OR2_X1 U13281 ( .A1(n10403), .A2(n10456), .ZN(n10352) );
  NAND2_X1 U13282 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10351) );
  OAI211_X1 U13283 ( .C1(n10394), .C2(n10353), .A(n10352), .B(n10351), .ZN(
        n10354) );
  AOI21_X1 U13284 ( .B1(n10404), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n10354), .ZN(n12985) );
  INV_X1 U13285 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n10781) );
  INV_X1 U13286 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n10732) );
  OR2_X1 U13287 ( .A1(n10403), .A2(n10732), .ZN(n10356) );
  NAND2_X1 U13288 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10355) );
  OAI211_X1 U13289 ( .C1(n10394), .C2(n10781), .A(n10356), .B(n10355), .ZN(
        n10357) );
  AOI21_X1 U13290 ( .B1(n10404), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10357), .ZN(n13929) );
  INV_X1 U13291 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19641) );
  NAND2_X1 U13292 ( .A1(n10404), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10360) );
  AOI22_X1 U13293 ( .A1(n10405), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n10359) );
  OAI211_X1 U13294 ( .C1(n10403), .C2(n19641), .A(n10360), .B(n10359), .ZN(
        n13887) );
  INV_X1 U13295 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n13941) );
  INV_X1 U13296 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19643) );
  OR2_X1 U13297 ( .A1(n10325), .A2(n19643), .ZN(n10362) );
  NAND2_X1 U13298 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10361) );
  OAI211_X1 U13299 ( .C1(n10394), .C2(n13941), .A(n10362), .B(n10361), .ZN(
        n10363) );
  AOI21_X1 U13300 ( .B1(n10404), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n10363), .ZN(n13938) );
  INV_X1 U13301 ( .A(n10364), .ZN(n14856) );
  INV_X1 U13302 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n10367) );
  INV_X1 U13303 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19645) );
  OR2_X1 U13304 ( .A1(n10403), .A2(n19645), .ZN(n10366) );
  NAND2_X1 U13305 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10365) );
  OAI211_X1 U13306 ( .C1(n10394), .C2(n10367), .A(n10366), .B(n10365), .ZN(
        n10368) );
  AOI21_X1 U13307 ( .B1(n10404), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n10368), .ZN(n14855) );
  INV_X1 U13308 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19647) );
  NAND2_X1 U13309 ( .A1(n10404), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10370) );
  AOI22_X1 U13310 ( .A1(n10405), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n10369) );
  OAI211_X1 U13311 ( .C1(n10403), .C2(n19647), .A(n10370), .B(n10369), .ZN(
        n14776) );
  INV_X1 U13312 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19649) );
  NAND2_X1 U13313 ( .A1(n10404), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10372) );
  AOI22_X1 U13314 ( .A1(n10405), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n10371) );
  OAI211_X1 U13315 ( .C1(n10403), .C2(n19649), .A(n10372), .B(n10371), .ZN(
        n14759) );
  INV_X1 U13316 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n10375) );
  INV_X1 U13317 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n10741) );
  OR2_X1 U13318 ( .A1(n10403), .A2(n10741), .ZN(n10374) );
  NAND2_X1 U13319 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10373) );
  OAI211_X1 U13320 ( .C1(n10394), .C2(n10375), .A(n10374), .B(n10373), .ZN(
        n10376) );
  AOI21_X1 U13321 ( .B1(n10404), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n10376), .ZN(n14751) );
  INV_X1 U13322 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10787) );
  INV_X1 U13323 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n10377) );
  OR2_X1 U13324 ( .A1(n10403), .A2(n10377), .ZN(n10379) );
  NAND2_X1 U13325 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10378) );
  OAI211_X1 U13326 ( .C1(n10394), .C2(n10787), .A(n10379), .B(n10378), .ZN(
        n10380) );
  AOI21_X1 U13327 ( .B1(n10404), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n10380), .ZN(n12997) );
  INV_X1 U13328 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n14834) );
  INV_X1 U13329 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n10381) );
  OR2_X1 U13330 ( .A1(n10403), .A2(n10381), .ZN(n10383) );
  NAND2_X1 U13331 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10382) );
  OAI211_X1 U13332 ( .C1(n10394), .C2(n14834), .A(n10383), .B(n10382), .ZN(
        n10384) );
  AOI21_X1 U13333 ( .B1(n10404), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n10384), .ZN(n14833) );
  INV_X1 U13334 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19654) );
  NAND2_X1 U13335 ( .A1(n10404), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10386) );
  AOI22_X1 U13336 ( .A1(n10405), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n10385) );
  OAI211_X1 U13337 ( .C1(n10403), .C2(n19654), .A(n10386), .B(n10385), .ZN(
        n14821) );
  INV_X1 U13338 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n10389) );
  INV_X1 U13339 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n14958) );
  OR2_X1 U13340 ( .A1(n10403), .A2(n14958), .ZN(n10388) );
  NAND2_X1 U13341 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10387) );
  OAI211_X1 U13342 ( .C1(n10394), .C2(n10389), .A(n10388), .B(n10387), .ZN(
        n10390) );
  AOI21_X1 U13343 ( .B1(n10404), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n10390), .ZN(n14810) );
  OR2_X2 U13344 ( .A1(n14809), .A2(n14810), .ZN(n14812) );
  INV_X1 U13345 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n10393) );
  INV_X1 U13346 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19658) );
  OR2_X1 U13347 ( .A1(n10403), .A2(n19658), .ZN(n10392) );
  NAND2_X1 U13348 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10391) );
  OAI211_X1 U13349 ( .C1(n10394), .C2(n10393), .A(n10392), .B(n10391), .ZN(
        n10395) );
  AOI21_X1 U13350 ( .B1(n10404), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10395), .ZN(n13009) );
  INV_X1 U13351 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n10398) );
  NAND2_X1 U13352 ( .A1(n10404), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10397) );
  AOI22_X1 U13353 ( .A1(n10405), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n10396) );
  OAI211_X1 U13354 ( .C1(n10403), .C2(n10398), .A(n10397), .B(n10396), .ZN(
        n12477) );
  INV_X1 U13355 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19659) );
  NAND2_X1 U13356 ( .A1(n10404), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10400) );
  AOI22_X1 U13357 ( .A1(n10405), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10399) );
  OAI211_X1 U13358 ( .C1(n10403), .C2(n19659), .A(n10400), .B(n10399), .ZN(
        n14024) );
  INV_X1 U13359 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n14007) );
  NAND2_X1 U13360 ( .A1(n10404), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10402) );
  AOI22_X1 U13361 ( .A1(n10405), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n10401) );
  OAI211_X1 U13362 ( .C1(n10403), .C2(n14007), .A(n10402), .B(n10401), .ZN(
        n12097) );
  AOI22_X1 U13363 ( .A1(n10405), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n10408) );
  NAND2_X1 U13364 ( .A1(n10406), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n10407) );
  OAI211_X1 U13365 ( .C1(n10311), .C2(n10409), .A(n10408), .B(n10407), .ZN(
        n10410) );
  INV_X1 U13366 ( .A(n10410), .ZN(n10411) );
  NAND2_X1 U13367 ( .A1(n10412), .A2(n19742), .ZN(n16173) );
  MUX2_X1 U13368 ( .A(n19710), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12489) );
  INV_X1 U13369 ( .A(n12261), .ZN(n10413) );
  NAND2_X1 U13370 ( .A1(n12489), .A2(n10413), .ZN(n10415) );
  NAND2_X1 U13371 ( .A1(n19710), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10414) );
  NAND2_X1 U13372 ( .A1(n10415), .A2(n10414), .ZN(n10424) );
  XNOR2_X1 U13373 ( .A(n19681), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10422) );
  NAND2_X1 U13374 ( .A1(n10424), .A2(n10422), .ZN(n10417) );
  NAND2_X1 U13375 ( .A1(n19700), .A2(n19681), .ZN(n10416) );
  XNOR2_X1 U13376 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10427) );
  NOR2_X1 U13377 ( .A1(n10136), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10418) );
  NAND2_X1 U13378 ( .A1(n16155), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10419) );
  NAND2_X1 U13379 ( .A1(n10426), .A2(n10419), .ZN(n10421) );
  NAND2_X1 U13380 ( .A1(n13139), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n10420) );
  XNOR2_X1 U13381 ( .A(n12489), .B(n12261), .ZN(n12491) );
  INV_X1 U13382 ( .A(n10422), .ZN(n10423) );
  XNOR2_X1 U13383 ( .A(n10424), .B(n10423), .ZN(n12497) );
  NOR2_X1 U13384 ( .A1(n16155), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10425) );
  NAND2_X1 U13385 ( .A1(n10426), .A2(n10425), .ZN(n10774) );
  INV_X1 U13386 ( .A(n10427), .ZN(n10428) );
  XNOR2_X1 U13387 ( .A(n10429), .B(n10428), .ZN(n10771) );
  NAND2_X1 U13388 ( .A1(n12497), .A2(n12502), .ZN(n12431) );
  INV_X1 U13389 ( .A(n12431), .ZN(n10430) );
  NAND2_X1 U13390 ( .A1(n12491), .A2(n10430), .ZN(n10431) );
  NAND2_X1 U13391 ( .A1(n19601), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10762) );
  INV_X1 U13392 ( .A(n10762), .ZN(n10432) );
  NAND2_X1 U13393 ( .A1(n16131), .A2(n19598), .ZN(n13030) );
  NAND2_X1 U13394 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19740) );
  NAND2_X1 U13395 ( .A1(n13031), .A2(n19740), .ZN(n13037) );
  OR2_X1 U13396 ( .A1(n13037), .A2(n10264), .ZN(n13043) );
  NAND2_X1 U13397 ( .A1(n10271), .A2(n19732), .ZN(n10478) );
  NOR2_X1 U13398 ( .A1(n10271), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10476) );
  AOI22_X1 U13399 ( .A1(n10752), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10455) );
  AND2_X2 U13400 ( .A1(n12776), .A2(n10136), .ZN(n12741) );
  AND2_X2 U13401 ( .A1(n10442), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10518) );
  AOI22_X1 U13402 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10446) );
  AND2_X2 U13403 ( .A1(n12754), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10457) );
  AND2_X2 U13404 ( .A1(n10434), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12697) );
  AOI22_X1 U13405 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10445) );
  INV_X1 U13406 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12924) );
  NAND2_X1 U13407 ( .A1(n10435), .A2(n12755), .ZN(n10592) );
  NOR2_X1 U13408 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10436) );
  INV_X1 U13409 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12737) );
  OAI22_X1 U13410 ( .A1(n12924), .A2(n10592), .B1(n12713), .B2(n12737), .ZN(
        n10441) );
  NAND2_X2 U13411 ( .A1(n10437), .A2(n12755), .ZN(n12734) );
  INV_X1 U13412 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12925) );
  INV_X1 U13413 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10439) );
  NAND3_X1 U13414 ( .A1(n19681), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12433) );
  INV_X1 U13415 ( .A(n12433), .ZN(n10438) );
  OAI22_X1 U13416 ( .A1(n12734), .A2(n12925), .B1(n10439), .B2(n12736), .ZN(
        n10440) );
  NOR2_X1 U13417 ( .A1(n10441), .A2(n10440), .ZN(n10444) );
  AND2_X2 U13418 ( .A1(n10442), .A2(n10136), .ZN(n12746) );
  AOI22_X1 U13419 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n12746), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10443) );
  NAND4_X1 U13420 ( .A1(n10446), .A2(n10445), .A3(n10444), .A4(n10443), .ZN(
        n10453) );
  INV_X1 U13421 ( .A(n10223), .ZN(n12923) );
  AND2_X2 U13422 ( .A1(n10223), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12723) );
  AOI22_X1 U13423 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12747), .B1(
        n12723), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10451) );
  NAND2_X1 U13424 ( .A1(n15425), .A2(n12755), .ZN(n12735) );
  AOI22_X1 U13425 ( .A1(n10527), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10450) );
  AND2_X2 U13426 ( .A1(n10226), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12725) );
  NAND2_X1 U13427 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10449) );
  AND2_X2 U13428 ( .A1(n12776), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12432) );
  NAND2_X1 U13429 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10448) );
  NAND4_X1 U13430 ( .A1(n10451), .A2(n10450), .A3(n10449), .A4(n10448), .ZN(
        n10452) );
  NOR2_X1 U13431 ( .A1(n10453), .A2(n10452), .ZN(n12621) );
  INV_X1 U13432 ( .A(n12621), .ZN(n13787) );
  NAND2_X1 U13433 ( .A1(n10726), .A2(n13787), .ZN(n10454) );
  OAI211_X1 U13434 ( .C1(n10755), .C2(n10456), .A(n10455), .B(n10454), .ZN(
        n12981) );
  AOI22_X1 U13435 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10461) );
  AOI22_X1 U13436 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10460) );
  AOI22_X1 U13437 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10527), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10459) );
  AOI22_X1 U13438 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12746), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10458) );
  NAND4_X1 U13439 ( .A1(n10461), .A2(n10460), .A3(n10459), .A4(n10458), .ZN(
        n10468) );
  INV_X1 U13440 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12628) );
  INV_X1 U13441 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12627) );
  OAI22_X1 U13442 ( .A1(n10592), .A2(n12628), .B1(n12734), .B2(n12627), .ZN(
        n10462) );
  INV_X1 U13443 ( .A(n10462), .ZN(n10466) );
  AOI22_X1 U13444 ( .A1(n12724), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10465) );
  AOI22_X1 U13445 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10464) );
  INV_X1 U13446 ( .A(n12736), .ZN(n10644) );
  AOI22_X1 U13447 ( .A1(n12747), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10644), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10463) );
  NAND4_X1 U13448 ( .A1(n10466), .A2(n10465), .A3(n10464), .A4(n10463), .ZN(
        n10467) );
  NOR2_X1 U13449 ( .A1(n10468), .A2(n10467), .ZN(n12443) );
  INV_X1 U13450 ( .A(n10469), .ZN(n10473) );
  INV_X1 U13451 ( .A(n10263), .ZN(n12942) );
  NAND2_X1 U13452 ( .A1(n12942), .A2(n9595), .ZN(n10513) );
  NOR2_X1 U13453 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19732), .ZN(
        n19717) );
  INV_X1 U13454 ( .A(n19717), .ZN(n10470) );
  NAND2_X1 U13455 ( .A1(n10478), .A2(n10470), .ZN(n10471) );
  AND2_X1 U13456 ( .A1(n10513), .A2(n10471), .ZN(n10472) );
  INV_X1 U13457 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18674) );
  INV_X1 U13458 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13039) );
  NAND2_X1 U13459 ( .A1(n19732), .A2(n13039), .ZN(n10474) );
  AOI22_X1 U13460 ( .A1(n10478), .A2(n10474), .B1(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13720), .ZN(n10475) );
  AOI22_X1 U13461 ( .A1(n10476), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10477) );
  OAI21_X1 U13462 ( .B1(n10755), .B2(n10247), .A(n10477), .ZN(n10497) );
  XNOR2_X1 U13463 ( .A(n13214), .B(n10497), .ZN(n13024) );
  INV_X1 U13464 ( .A(n10478), .ZN(n10480) );
  AND2_X1 U13465 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10479) );
  AOI21_X1 U13466 ( .B1(n10480), .B2(n10263), .A(n10479), .ZN(n10496) );
  AOI22_X1 U13467 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13468 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10487) );
  INV_X1 U13469 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12638) );
  NAND2_X1 U13470 ( .A1(n12748), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10481) );
  OAI21_X1 U13471 ( .B1(n10592), .B2(n12638), .A(n10481), .ZN(n10484) );
  INV_X1 U13472 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12637) );
  INV_X1 U13473 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10482) );
  OAI22_X1 U13474 ( .A1(n12734), .A2(n12637), .B1(n10482), .B2(n12736), .ZN(
        n10483) );
  NOR2_X1 U13475 ( .A1(n10484), .A2(n10483), .ZN(n10486) );
  AOI22_X1 U13476 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12746), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10485) );
  NAND4_X1 U13477 ( .A1(n10488), .A2(n10487), .A3(n10486), .A4(n10485), .ZN(
        n10494) );
  AOI22_X1 U13478 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12747), .B1(
        n12723), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13479 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n10527), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10491) );
  NAND2_X1 U13480 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10490) );
  NAND2_X1 U13481 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10489) );
  NAND4_X1 U13482 ( .A1(n10492), .A2(n10491), .A3(n10490), .A4(n10489), .ZN(
        n10493) );
  NAND2_X1 U13483 ( .A1(n10726), .A2(n12442), .ZN(n10495) );
  NAND2_X1 U13484 ( .A1(n10496), .A2(n10495), .ZN(n13023) );
  NOR2_X1 U13485 ( .A1(n13024), .A2(n13023), .ZN(n10499) );
  NOR2_X1 U13486 ( .A1(n13214), .A2(n10497), .ZN(n10498) );
  AOI22_X1 U13487 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12741), .B1(
        n12432), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10506) );
  INV_X1 U13488 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12806) );
  INV_X1 U13489 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12651) );
  OAI22_X1 U13490 ( .A1(n12806), .A2(n12735), .B1(n12734), .B2(n12651), .ZN(
        n10502) );
  INV_X1 U13491 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12652) );
  INV_X1 U13492 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10500) );
  OAI22_X1 U13493 ( .A1(n10592), .A2(n12652), .B1(n10500), .B2(n12736), .ZN(
        n10501) );
  NOR2_X1 U13494 ( .A1(n10502), .A2(n10501), .ZN(n10505) );
  AOI22_X1 U13495 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10504) );
  AOI22_X1 U13496 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12746), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10503) );
  NAND4_X1 U13497 ( .A1(n10506), .A2(n10505), .A3(n10504), .A4(n10503), .ZN(
        n10511) );
  AOI22_X1 U13498 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U13499 ( .A1(n10527), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10508) );
  AOI22_X1 U13500 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12747), .B1(
        n12723), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10507) );
  NAND3_X1 U13501 ( .A1(n10509), .A2(n10508), .A3(n10507), .ZN(n10510) );
  NAND2_X1 U13502 ( .A1(n10726), .A2(n10765), .ZN(n10512) );
  OAI211_X1 U13503 ( .C1(n19732), .C2(n19700), .A(n10513), .B(n10512), .ZN(
        n10515) );
  XNOR2_X1 U13504 ( .A(n10516), .B(n10515), .ZN(n13277) );
  INV_X1 U13505 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12553) );
  AOI22_X1 U13506 ( .A1(n10752), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10514) );
  OAI21_X1 U13507 ( .B1(n10755), .B2(n13818), .A(n10514), .ZN(n13276) );
  NOR2_X1 U13508 ( .A1(n10516), .A2(n10515), .ZN(n10517) );
  AOI22_X1 U13509 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U13510 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10525) );
  INV_X1 U13511 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12668) );
  NAND2_X1 U13512 ( .A1(n12748), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10519) );
  OAI21_X1 U13513 ( .B1(n12668), .B2(n10592), .A(n10519), .ZN(n10521) );
  INV_X1 U13514 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12667) );
  INV_X1 U13515 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12590) );
  OAI22_X1 U13516 ( .A1(n12734), .A2(n12667), .B1(n12736), .B2(n12590), .ZN(
        n10520) );
  NOR2_X1 U13517 ( .A1(n10521), .A2(n10520), .ZN(n10524) );
  AOI22_X1 U13518 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12746), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10523) );
  NAND4_X1 U13519 ( .A1(n10526), .A2(n10525), .A3(n10524), .A4(n10523), .ZN(
        n10533) );
  AOI22_X1 U13520 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10531) );
  AOI22_X1 U13521 ( .A1(n10527), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10530) );
  NAND2_X1 U13522 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10529) );
  NAND2_X1 U13523 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10528) );
  NAND4_X1 U13524 ( .A1(n10531), .A2(n10530), .A3(n10529), .A4(n10528), .ZN(
        n10532) );
  AOI22_X1 U13525 ( .A1(n10726), .A2(n12254), .B1(n10752), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13526 ( .A1(n9595), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n10534) );
  OAI211_X1 U13527 ( .C1(n10536), .C2(n10755), .A(n10535), .B(n10534), .ZN(
        n13560) );
  AOI22_X1 U13528 ( .A1(n10752), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10550) );
  AOI22_X1 U13529 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10542) );
  AOI22_X1 U13530 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U13531 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10540) );
  INV_X1 U13532 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12852) );
  INV_X1 U13533 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12682) );
  OAI22_X1 U13534 ( .A1(n12735), .A2(n12852), .B1(n12734), .B2(n12682), .ZN(
        n10538) );
  INV_X1 U13535 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12683) );
  INV_X1 U13536 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12615) );
  OAI22_X1 U13537 ( .A1(n10592), .A2(n12683), .B1(n12736), .B2(n12615), .ZN(
        n10537) );
  NOR2_X1 U13538 ( .A1(n10538), .A2(n10537), .ZN(n10539) );
  NAND4_X1 U13539 ( .A1(n10542), .A2(n10541), .A3(n10540), .A4(n10539), .ZN(
        n10548) );
  AOI22_X1 U13540 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10527), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10546) );
  AOI22_X1 U13541 ( .A1(n12747), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10545) );
  NAND2_X1 U13542 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10544) );
  NAND2_X1 U13543 ( .A1(n12746), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10543) );
  NAND4_X1 U13544 ( .A1(n10546), .A2(n10545), .A3(n10544), .A4(n10543), .ZN(
        n10547) );
  NAND2_X1 U13545 ( .A1(n10726), .A2(n12277), .ZN(n10549) );
  OAI211_X1 U13546 ( .C1(n10755), .C2(n10551), .A(n10550), .B(n10549), .ZN(
        n13565) );
  AOI22_X1 U13547 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10559) );
  AOI22_X1 U13548 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10558) );
  INV_X1 U13549 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12699) );
  NAND2_X1 U13550 ( .A1(n12748), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10552) );
  OAI21_X1 U13551 ( .B1(n12699), .B2(n10592), .A(n10552), .ZN(n10555) );
  INV_X1 U13552 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12698) );
  INV_X1 U13553 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10553) );
  OAI22_X1 U13554 ( .A1(n12734), .A2(n12698), .B1(n10553), .B2(n12736), .ZN(
        n10554) );
  NOR2_X1 U13555 ( .A1(n10555), .A2(n10554), .ZN(n10557) );
  AOI22_X1 U13556 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12746), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10556) );
  NAND4_X1 U13557 ( .A1(n10559), .A2(n10558), .A3(n10557), .A4(n10556), .ZN(
        n10565) );
  AOI22_X1 U13558 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10563) );
  AOI22_X1 U13559 ( .A1(n10527), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10562) );
  NAND2_X1 U13560 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10561) );
  NAND2_X1 U13561 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10560) );
  NAND4_X1 U13562 ( .A1(n10563), .A2(n10562), .A3(n10561), .A4(n10560), .ZN(
        n10564) );
  INV_X1 U13563 ( .A(n12296), .ZN(n10566) );
  AOI22_X1 U13564 ( .A1(n10756), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n10726), 
        .B2(n10566), .ZN(n10568) );
  AOI22_X1 U13565 ( .A1(n10752), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10567) );
  NAND2_X1 U13566 ( .A1(n10568), .A2(n10567), .ZN(n15394) );
  AOI22_X1 U13567 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12741), .B1(
        n12432), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10576) );
  INV_X1 U13568 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12715) );
  NAND2_X1 U13569 ( .A1(n12748), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10569) );
  OAI21_X1 U13570 ( .B1(n10592), .B2(n12715), .A(n10569), .ZN(n10572) );
  INV_X1 U13571 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12714) );
  INV_X1 U13572 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10570) );
  OAI22_X1 U13573 ( .A1(n12734), .A2(n12714), .B1(n10570), .B2(n12736), .ZN(
        n10571) );
  NOR2_X1 U13574 ( .A1(n10572), .A2(n10571), .ZN(n10575) );
  AOI22_X1 U13575 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10574) );
  AOI22_X1 U13576 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10518), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10573) );
  NAND4_X1 U13577 ( .A1(n10576), .A2(n10575), .A3(n10574), .A4(n10573), .ZN(
        n10581) );
  AOI22_X1 U13578 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12746), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10579) );
  AOI22_X1 U13579 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10527), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10578) );
  AOI22_X1 U13580 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12747), .B1(
        n12723), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10577) );
  NAND3_X1 U13581 ( .A1(n10579), .A2(n10578), .A3(n10577), .ZN(n10580) );
  INV_X1 U13582 ( .A(n12321), .ZN(n10582) );
  NAND2_X1 U13583 ( .A1(n10726), .A2(n10582), .ZN(n10583) );
  AOI22_X1 U13584 ( .A1(n10752), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10584) );
  OAI21_X1 U13585 ( .B1(n10755), .B2(n10332), .A(n10584), .ZN(n15385) );
  NAND2_X1 U13586 ( .A1(n15387), .A2(n15385), .ZN(n10603) );
  AOI22_X1 U13587 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12746), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10587) );
  AOI22_X1 U13588 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n10527), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10586) );
  AOI22_X1 U13589 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12747), .B1(
        n12723), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10585) );
  NAND2_X1 U13590 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10591) );
  NAND2_X1 U13591 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10590) );
  NAND2_X1 U13592 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10589) );
  NAND2_X1 U13593 ( .A1(n10518), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10588) );
  NAND4_X1 U13594 ( .A1(n10591), .A2(n10590), .A3(n10589), .A4(n10588), .ZN(
        n10599) );
  NAND2_X1 U13595 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10597) );
  INV_X1 U13596 ( .A(n10592), .ZN(n10645) );
  AOI22_X1 U13597 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10596) );
  INV_X1 U13598 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12738) );
  INV_X1 U13599 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12922) );
  OAI22_X1 U13600 ( .A1(n12734), .A2(n12738), .B1(n12922), .B2(n12736), .ZN(
        n10593) );
  INV_X1 U13601 ( .A(n10593), .ZN(n10595) );
  NAND2_X1 U13602 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10594) );
  NAND4_X1 U13603 ( .A1(n10597), .A2(n10596), .A3(n10595), .A4(n10594), .ZN(
        n10598) );
  NAND2_X1 U13604 ( .A1(n10726), .A2(n14000), .ZN(n10602) );
  AOI22_X1 U13605 ( .A1(n10752), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10604) );
  OAI21_X1 U13606 ( .B1(n10755), .B2(n10335), .A(n10604), .ZN(n15360) );
  INV_X1 U13607 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U13608 ( .A1(n10752), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13609 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10611) );
  AOI22_X1 U13610 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10610) );
  AOI22_X1 U13611 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10609) );
  INV_X1 U13612 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12759) );
  OAI22_X1 U13613 ( .A1(n12735), .A2(n12627), .B1(n12734), .B2(n12759), .ZN(
        n10607) );
  INV_X1 U13614 ( .A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12626) );
  INV_X1 U13615 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10605) );
  OAI22_X1 U13616 ( .A1(n10592), .A2(n12626), .B1(n12736), .B2(n10605), .ZN(
        n10606) );
  NOR2_X1 U13617 ( .A1(n10607), .A2(n10606), .ZN(n10608) );
  NAND4_X1 U13618 ( .A1(n10611), .A2(n10610), .A3(n10609), .A4(n10608), .ZN(
        n10617) );
  AOI22_X1 U13619 ( .A1(n12747), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10527), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U13620 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10614) );
  NAND2_X1 U13621 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10613) );
  NAND2_X1 U13622 ( .A1(n12746), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10612) );
  NAND4_X1 U13623 ( .A1(n10615), .A2(n10614), .A3(n10613), .A4(n10612), .ZN(
        n10616) );
  NOR2_X1 U13624 ( .A1(n10617), .A2(n10616), .ZN(n13536) );
  INV_X1 U13625 ( .A(n13536), .ZN(n13538) );
  NAND2_X1 U13626 ( .A1(n10726), .A2(n13538), .ZN(n10618) );
  OAI211_X1 U13627 ( .C1(n10755), .C2(n10620), .A(n10619), .B(n10618), .ZN(
        n16094) );
  INV_X1 U13628 ( .A(n16094), .ZN(n10621) );
  AOI22_X1 U13629 ( .A1(n10752), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10637) );
  AOI22_X1 U13630 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10629) );
  AOI22_X1 U13631 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10628) );
  INV_X1 U13632 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12779) );
  OAI22_X1 U13633 ( .A1(n12779), .A2(n10592), .B1(n12713), .B2(n12638), .ZN(
        n10625) );
  INV_X1 U13634 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10623) );
  INV_X1 U13635 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10622) );
  OAI22_X1 U13636 ( .A1(n12734), .A2(n10623), .B1(n10622), .B2(n12736), .ZN(
        n10624) );
  NOR2_X1 U13637 ( .A1(n10625), .A2(n10624), .ZN(n10627) );
  AOI22_X1 U13638 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n10522), .B1(
        n12746), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10626) );
  NAND4_X1 U13639 ( .A1(n10629), .A2(n10628), .A3(n10627), .A4(n10626), .ZN(
        n10635) );
  AOI22_X1 U13640 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12747), .B1(
        n12723), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10633) );
  AOI22_X1 U13641 ( .A1(n10527), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10632) );
  NAND2_X1 U13642 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10631) );
  NAND2_X1 U13643 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10630) );
  NAND4_X1 U13644 ( .A1(n10633), .A2(n10632), .A3(n10631), .A4(n10630), .ZN(
        n10634) );
  NOR2_X1 U13645 ( .A1(n10635), .A2(n10634), .ZN(n13670) );
  INV_X1 U13646 ( .A(n13670), .ZN(n13672) );
  NAND2_X1 U13647 ( .A1(n10726), .A2(n13672), .ZN(n10636) );
  OAI211_X1 U13648 ( .C1(n10755), .C2(n10638), .A(n10637), .B(n10636), .ZN(
        n15351) );
  AOI22_X1 U13649 ( .A1(n10752), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10658) );
  NAND2_X1 U13650 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10642) );
  NAND2_X1 U13651 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10641) );
  NAND2_X1 U13652 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10640) );
  NAND2_X1 U13653 ( .A1(n10518), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10639) );
  NAND4_X1 U13654 ( .A1(n10642), .A2(n10641), .A3(n10640), .A4(n10639), .ZN(
        n10651) );
  NAND2_X1 U13655 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10649) );
  INV_X1 U13656 ( .A(n12734), .ZN(n10643) );
  AOI22_X1 U13657 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12724), .B1(
        n10643), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10648) );
  AOI22_X1 U13658 ( .A1(n10645), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n10644), .ZN(n10647) );
  NAND2_X1 U13659 ( .A1(n12697), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10646) );
  NAND4_X1 U13660 ( .A1(n10649), .A2(n10648), .A3(n10647), .A4(n10646), .ZN(
        n10650) );
  NOR2_X1 U13661 ( .A1(n10651), .A2(n10650), .ZN(n10656) );
  AOI22_X1 U13662 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n10522), .B1(
        n12746), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10654) );
  AOI22_X1 U13663 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12747), .B1(
        n12723), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U13664 ( .A1(n10527), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10652) );
  AND3_X1 U13665 ( .A1(n10654), .A2(n10653), .A3(n10652), .ZN(n10655) );
  INV_X1 U13666 ( .A(n13738), .ZN(n13741) );
  NAND2_X1 U13667 ( .A1(n10726), .A2(n13741), .ZN(n10657) );
  OAI211_X1 U13668 ( .C1(n10755), .C2(n10659), .A(n10658), .B(n10657), .ZN(
        n15331) );
  AOI22_X1 U13669 ( .A1(n10752), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10675) );
  AOI22_X1 U13670 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U13671 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10666) );
  INV_X1 U13672 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12830) );
  OAI22_X1 U13673 ( .A1(n10592), .A2(n12830), .B1(n12713), .B2(n12668), .ZN(
        n10663) );
  INV_X1 U13674 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10661) );
  INV_X1 U13675 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10660) );
  OAI22_X1 U13676 ( .A1(n12734), .A2(n10661), .B1(n12736), .B2(n10660), .ZN(
        n10662) );
  NOR2_X1 U13677 ( .A1(n10663), .A2(n10662), .ZN(n10665) );
  AOI22_X1 U13678 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12746), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10664) );
  NAND4_X1 U13679 ( .A1(n10667), .A2(n10666), .A3(n10665), .A4(n10664), .ZN(
        n10673) );
  AOI22_X1 U13680 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U13681 ( .A1(n10527), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10670) );
  NAND2_X1 U13682 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10669) );
  NAND2_X1 U13683 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10668) );
  NAND4_X1 U13684 ( .A1(n10671), .A2(n10670), .A3(n10669), .A4(n10668), .ZN(
        n10672) );
  OR2_X1 U13685 ( .A1(n10673), .A2(n10672), .ZN(n13777) );
  NAND2_X1 U13686 ( .A1(n10726), .A2(n13777), .ZN(n10674) );
  OAI211_X1 U13687 ( .C1(n10755), .C2(n10676), .A(n10675), .B(n10674), .ZN(
        n15314) );
  AOI22_X1 U13688 ( .A1(n10752), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U13689 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10684) );
  AOI22_X1 U13690 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10683) );
  OAI22_X1 U13691 ( .A1(n10592), .A2(n12852), .B1(n12713), .B2(n12683), .ZN(
        n10680) );
  INV_X1 U13692 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10678) );
  INV_X1 U13693 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10677) );
  OAI22_X1 U13694 ( .A1(n12734), .A2(n10678), .B1(n12736), .B2(n10677), .ZN(
        n10679) );
  NOR2_X1 U13695 ( .A1(n10680), .A2(n10679), .ZN(n10682) );
  AOI22_X1 U13696 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12746), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10681) );
  NAND4_X1 U13697 ( .A1(n10684), .A2(n10683), .A3(n10682), .A4(n10681), .ZN(
        n10690) );
  AOI22_X1 U13698 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U13699 ( .A1(n10527), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10687) );
  NAND2_X1 U13700 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10686) );
  NAND2_X1 U13701 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10685) );
  NAND4_X1 U13702 ( .A1(n10688), .A2(n10687), .A3(n10686), .A4(n10685), .ZN(
        n10689) );
  OR2_X1 U13703 ( .A1(n10690), .A2(n10689), .ZN(n13768) );
  NAND2_X1 U13704 ( .A1(n10726), .A2(n13768), .ZN(n10691) );
  OAI211_X1 U13705 ( .C1(n10755), .C2(n10693), .A(n10692), .B(n10691), .ZN(
        n15291) );
  INV_X1 U13706 ( .A(n15291), .ZN(n10694) );
  AOI22_X1 U13707 ( .A1(n10752), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10710) );
  AOI22_X1 U13708 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10702) );
  AOI22_X1 U13709 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10701) );
  INV_X1 U13710 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12875) );
  OAI22_X1 U13711 ( .A1(n10592), .A2(n12875), .B1(n12713), .B2(n12699), .ZN(
        n10698) );
  INV_X1 U13712 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10696) );
  INV_X1 U13713 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10695) );
  OAI22_X1 U13714 ( .A1(n12734), .A2(n10696), .B1(n12736), .B2(n10695), .ZN(
        n10697) );
  NOR2_X1 U13715 ( .A1(n10698), .A2(n10697), .ZN(n10700) );
  AOI22_X1 U13716 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12746), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10699) );
  NAND4_X1 U13717 ( .A1(n10702), .A2(n10701), .A3(n10700), .A4(n10699), .ZN(
        n10708) );
  AOI22_X1 U13718 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10706) );
  AOI22_X1 U13719 ( .A1(n10527), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10705) );
  NAND2_X1 U13720 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10704) );
  NAND2_X1 U13721 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10703) );
  NAND4_X1 U13722 ( .A1(n10706), .A2(n10705), .A3(n10704), .A4(n10703), .ZN(
        n10707) );
  NAND2_X1 U13723 ( .A1(n10726), .A2(n13727), .ZN(n10709) );
  OAI211_X1 U13724 ( .C1(n10755), .C2(n10711), .A(n10710), .B(n10709), .ZN(
        n15271) );
  NAND2_X1 U13725 ( .A1(n15270), .A2(n15271), .ZN(n15272) );
  AOI22_X1 U13726 ( .A1(n10752), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10728) );
  AOI22_X1 U13727 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10719) );
  AOI22_X1 U13728 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10718) );
  INV_X1 U13729 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12903) );
  OAI22_X1 U13730 ( .A1(n12903), .A2(n10592), .B1(n12713), .B2(n12715), .ZN(
        n10715) );
  INV_X1 U13731 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10713) );
  INV_X1 U13732 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10712) );
  OAI22_X1 U13733 ( .A1(n12734), .A2(n10713), .B1(n10712), .B2(n12736), .ZN(
        n10714) );
  NOR2_X1 U13734 ( .A1(n10715), .A2(n10714), .ZN(n10717) );
  AOI22_X1 U13735 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10518), .B1(
        n12746), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10716) );
  NAND4_X1 U13736 ( .A1(n10719), .A2(n10718), .A3(n10717), .A4(n10716), .ZN(
        n10725) );
  AOI22_X1 U13737 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12747), .B1(
        n10527), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10723) );
  AOI22_X1 U13738 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10722) );
  NAND2_X1 U13739 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10721) );
  NAND2_X1 U13740 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10720) );
  NAND4_X1 U13741 ( .A1(n10723), .A2(n10722), .A3(n10721), .A4(n10720), .ZN(
        n10724) );
  NAND2_X1 U13742 ( .A1(n10726), .A2(n13702), .ZN(n10727) );
  OAI211_X1 U13743 ( .C1(n10755), .C2(n10729), .A(n10728), .B(n10727), .ZN(
        n15250) );
  INV_X1 U13744 ( .A(n15250), .ZN(n10730) );
  AOI22_X1 U13745 ( .A1(n10752), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10731) );
  OAI21_X1 U13746 ( .B1(n10755), .B2(n10732), .A(n10731), .ZN(n15231) );
  NAND2_X1 U13747 ( .A1(n10756), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U13748 ( .A1(n10752), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10733) );
  AND2_X1 U13749 ( .A1(n10734), .A2(n10733), .ZN(n13872) );
  NAND2_X1 U13750 ( .A1(n10756), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n10736) );
  AOI22_X1 U13751 ( .A1(n10752), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10735) );
  AND2_X1 U13752 ( .A1(n10736), .A2(n10735), .ZN(n15195) );
  AOI22_X1 U13753 ( .A1(n10752), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10737) );
  OAI21_X1 U13754 ( .B1(n10755), .B2(n19645), .A(n10737), .ZN(n14927) );
  AOI22_X1 U13755 ( .A1(n10752), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10738) );
  OAI21_X1 U13756 ( .B1(n10755), .B2(n19647), .A(n10738), .ZN(n14786) );
  AOI22_X1 U13757 ( .A1(n10752), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10739) );
  OAI21_X1 U13758 ( .B1(n10755), .B2(n19649), .A(n10739), .ZN(n14763) );
  AOI22_X1 U13759 ( .A1(n10752), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10740) );
  OAI21_X1 U13760 ( .B1(n10755), .B2(n10741), .A(n10740), .ZN(n14752) );
  AOI22_X1 U13761 ( .A1(n10752), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10742) );
  OAI21_X1 U13762 ( .B1(n10755), .B2(n10377), .A(n10742), .ZN(n12999) );
  NAND2_X1 U13763 ( .A1(n10756), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U13764 ( .A1(n10752), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10743) );
  AND2_X1 U13765 ( .A1(n10744), .A2(n10743), .ZN(n14908) );
  NAND2_X1 U13766 ( .A1(n10756), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n10746) );
  AOI22_X1 U13767 ( .A1(n10752), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10745) );
  AND2_X1 U13768 ( .A1(n10746), .A2(n10745), .ZN(n14897) );
  AOI22_X1 U13769 ( .A1(n10752), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10747) );
  OAI21_X1 U13770 ( .B1(n10755), .B2(n14958), .A(n10747), .ZN(n14888) );
  NAND2_X1 U13771 ( .A1(n10756), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U13772 ( .A1(n10752), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10748) );
  AND2_X1 U13773 ( .A1(n10749), .A2(n10748), .ZN(n13013) );
  NAND2_X1 U13774 ( .A1(n10756), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n10751) );
  AOI22_X1 U13775 ( .A1(n10752), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10750) );
  AND2_X1 U13776 ( .A1(n10751), .A2(n10750), .ZN(n12562) );
  AOI22_X1 U13777 ( .A1(n10752), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10753) );
  OAI21_X1 U13778 ( .B1(n10755), .B2(n19659), .A(n10753), .ZN(n14866) );
  AOI22_X1 U13779 ( .A1(n10752), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n9595), .B2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10754) );
  OAI21_X1 U13780 ( .B1(n10755), .B2(n14007), .A(n10754), .ZN(n12081) );
  AOI222_X1 U13781 ( .A1(n10756), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n10752), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n9595), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10757) );
  INV_X1 U13782 ( .A(n10757), .ZN(n10758) );
  NAND2_X1 U13783 ( .A1(n10760), .A2(n16173), .ZN(n16133) );
  NAND2_X1 U13784 ( .A1(n16133), .A2(n16131), .ZN(n16142) );
  INV_X1 U13785 ( .A(n19598), .ZN(n18657) );
  NAND2_X1 U13786 ( .A1(n20805), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19753) );
  INV_X2 U13787 ( .A(n19753), .ZN(n19752) );
  NAND2_X2 U13788 ( .A1(n19752), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19662) );
  NOR2_X1 U13789 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n18656) );
  INV_X1 U13790 ( .A(n18656), .ZN(n19618) );
  NAND2_X1 U13791 ( .A1(n19740), .A2(n19744), .ZN(n16139) );
  NOR2_X1 U13792 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n16139), .ZN(n16170) );
  NAND3_X1 U13793 ( .A1(n19742), .A2(n10264), .A3(n16170), .ZN(n10761) );
  NOR2_X2 U13794 ( .A1(n19735), .A2(n10761), .ZN(n18877) );
  NOR2_X2 U13795 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19688) );
  AND2_X2 U13796 ( .A1(n19734), .A2(n19688), .ZN(n19011) );
  NOR3_X1 U13797 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10762), .A3(n19732), 
        .ZN(n16167) );
  OR2_X1 U13798 ( .A1(n19011), .A2(n16167), .ZN(n10763) );
  NOR2_X1 U13799 ( .A1(n18882), .A2(n10763), .ZN(n10764) );
  NAND2_X1 U13800 ( .A1(n18849), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18874) );
  INV_X1 U13801 ( .A(n10765), .ZN(n12449) );
  INV_X1 U13802 ( .A(n12497), .ZN(n12495) );
  MUX2_X1 U13803 ( .A(n12449), .B(n12495), .S(n10766), .Z(n12427) );
  BUF_X1 U13804 ( .A(n10767), .Z(n10768) );
  INV_X1 U13805 ( .A(n12442), .ZN(n10770) );
  INV_X1 U13806 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13123) );
  INV_X1 U13807 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n20734) );
  NAND2_X1 U13808 ( .A1(n13123), .A2(n20734), .ZN(n10769) );
  MUX2_X1 U13809 ( .A(n10770), .B(n10769), .S(n10768), .Z(n12265) );
  MUX2_X1 U13810 ( .A(n12254), .B(n10771), .S(n10766), .Z(n10773) );
  MUX2_X1 U13811 ( .A(n10773), .B(n10772), .S(n10768), .Z(n12259) );
  MUX2_X1 U13812 ( .A(n12277), .B(n10774), .S(n10766), .Z(n10775) );
  INV_X1 U13813 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n18856) );
  MUX2_X1 U13814 ( .A(n10775), .B(n18856), .S(n10768), .Z(n12269) );
  MUX2_X1 U13815 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n12296), .S(n10234), .Z(
        n12301) );
  MUX2_X1 U13816 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n12321), .S(n10234), .Z(
        n12325) );
  MUX2_X1 U13817 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n14002), .S(n10234), .Z(
        n12330) );
  NAND2_X1 U13818 ( .A1(n10768), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12334) );
  INV_X1 U13819 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10777) );
  INV_X1 U13820 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n12341) );
  NAND2_X1 U13821 ( .A1(n10768), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12355) );
  INV_X1 U13822 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10779) );
  NOR2_X1 U13823 ( .A1(n10234), .A2(n10779), .ZN(n12358) );
  INV_X1 U13824 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n10780) );
  NOR2_X1 U13825 ( .A1(n10234), .A2(n10780), .ZN(n12378) );
  NAND2_X1 U13826 ( .A1(n10768), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12380) );
  NOR2_X1 U13827 ( .A1(n10234), .A2(n10781), .ZN(n10782) );
  INV_X1 U13828 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10783) );
  NOR2_X1 U13829 ( .A1(n10234), .A2(n10783), .ZN(n12371) );
  NOR2_X1 U13830 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(P2_EBX_REG_19__SCAN_IN), 
        .ZN(n10784) );
  NOR2_X1 U13831 ( .A1(n10234), .A2(n10784), .ZN(n10785) );
  INV_X1 U13832 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n14852) );
  INV_X1 U13833 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n14848) );
  NAND2_X1 U13834 ( .A1(n10768), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12398) );
  NOR2_X1 U13835 ( .A1(n10234), .A2(n10787), .ZN(n12402) );
  INV_X1 U13836 ( .A(n12405), .ZN(n10788) );
  NOR2_X1 U13837 ( .A1(n12413), .A2(n10788), .ZN(n12409) );
  INV_X1 U13838 ( .A(n12409), .ZN(n10789) );
  NAND2_X1 U13839 ( .A1(n10768), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12414) );
  NAND2_X1 U13840 ( .A1(n10789), .A2(n12414), .ZN(n12423) );
  NAND2_X1 U13841 ( .A1(n10768), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12421) );
  INV_X1 U13842 ( .A(n12420), .ZN(n10791) );
  NAND2_X1 U13843 ( .A1(n10768), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13998) );
  NAND2_X1 U13844 ( .A1(n10791), .A2(n13998), .ZN(n12087) );
  NAND2_X1 U13845 ( .A1(n10768), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12086) );
  INV_X1 U13846 ( .A(n12086), .ZN(n10794) );
  NAND2_X1 U13847 ( .A1(n19682), .A2(n19740), .ZN(n12088) );
  NAND3_X1 U13848 ( .A1(n12536), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n12088), 
        .ZN(n10793) );
  NOR3_X1 U13849 ( .A1(n12087), .A2(n10794), .A3(n18888), .ZN(n10796) );
  INV_X1 U13850 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n14795) );
  OR2_X1 U13851 ( .A1(n13108), .A2(n16170), .ZN(n12090) );
  INV_X1 U13852 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19664) );
  OAI22_X1 U13853 ( .A1(n14795), .A2(n12090), .B1(n19664), .B2(n18849), .ZN(
        n10795) );
  AOI211_X1 U13854 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n18901), .A(
        n10796), .B(n10795), .ZN(n10797) );
  NAND2_X1 U13855 ( .A1(n10802), .A2(n10801), .ZN(P2_U2824) );
  AOI22_X1 U13856 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U13857 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10890), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10805) );
  INV_X2 U13858 ( .A(n10962), .ZN(n16947) );
  AOI22_X1 U13859 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10804) );
  AOI22_X1 U13860 ( .A1(n16883), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15510), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10803) );
  NAND4_X1 U13861 ( .A1(n10806), .A2(n10805), .A3(n10804), .A4(n10803), .ZN(
        n10817) );
  INV_X2 U13862 ( .A(n13977), .ZN(n16946) );
  AOI22_X1 U13863 ( .A1(n16946), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16952), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10815) );
  AOI22_X1 U13865 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U13866 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10813) );
  INV_X2 U13867 ( .A(n11016), .ZN(n16872) );
  AOI22_X1 U13868 ( .A1(n16839), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10812) );
  NAND4_X1 U13869 ( .A1(n10815), .A2(n10814), .A3(n10813), .A4(n10812), .ZN(
        n10816) );
  AOI22_X1 U13870 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10890), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U13871 ( .A1(n16946), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10820) );
  INV_X4 U13872 ( .A(n15509), .ZN(n16955) );
  INV_X2 U13873 ( .A(n10809), .ZN(n15525) );
  AOI22_X1 U13874 ( .A1(n16955), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10819) );
  AOI22_X1 U13875 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15510), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10818) );
  NAND4_X1 U13876 ( .A1(n10821), .A2(n10820), .A3(n10819), .A4(n10818), .ZN(
        n10827) );
  AOI22_X1 U13877 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10825) );
  AOI22_X1 U13878 ( .A1(n16839), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16952), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10824) );
  INV_X2 U13879 ( .A(n9695), .ZN(n16954) );
  AOI22_X1 U13880 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U13881 ( .A1(n16883), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10822) );
  NAND4_X1 U13882 ( .A1(n10825), .A2(n10824), .A3(n10823), .A4(n10822), .ZN(
        n10826) );
  AOI22_X1 U13883 ( .A1(n16839), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16844), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10831) );
  AOI22_X1 U13884 ( .A1(n16883), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10830) );
  AOI22_X1 U13885 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10829) );
  AOI22_X1 U13886 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15510), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10828) );
  NAND4_X1 U13887 ( .A1(n10831), .A2(n10830), .A3(n10829), .A4(n10828), .ZN(
        n10837) );
  AOI22_X1 U13888 ( .A1(n16946), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10835) );
  AOI22_X1 U13889 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10834) );
  AOI22_X1 U13890 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10833) );
  AOI22_X1 U13891 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10832) );
  NAND4_X1 U13892 ( .A1(n10835), .A2(n10834), .A3(n10833), .A4(n10832), .ZN(
        n10836) );
  AOI22_X1 U13893 ( .A1(n16946), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10890), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U13894 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16844), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10839) );
  NAND3_X1 U13895 ( .A1(n10840), .A2(n10839), .A3(n10838), .ZN(n10849) );
  INV_X1 U13896 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n16993) );
  OAI21_X1 U13897 ( .B1(n9694), .B2(n16993), .A(n10841), .ZN(n10848) );
  AOI22_X1 U13898 ( .A1(n16839), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10858), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U13899 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10867), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U13900 ( .A1(n10852), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10842), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10844) );
  AOI22_X1 U13901 ( .A1(n10889), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10843) );
  NAND4_X1 U13902 ( .A1(n10846), .A2(n10845), .A3(n10844), .A4(n10843), .ZN(
        n10847) );
  INV_X1 U13903 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n20848) );
  AOI22_X1 U13904 ( .A1(n16955), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10850) );
  OAI21_X1 U13905 ( .B1(n10962), .B2(n20848), .A(n10850), .ZN(n10851) );
  AOI22_X1 U13906 ( .A1(n10877), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10889), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U13907 ( .A1(n16927), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10890), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10856) );
  AOI22_X1 U13908 ( .A1(n10853), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10852), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U13909 ( .A1(n15510), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10867), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10854) );
  NAND4_X1 U13910 ( .A1(n10857), .A2(n10856), .A3(n10855), .A4(n10854), .ZN(
        n10863) );
  AOI22_X1 U13911 ( .A1(n16839), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10861) );
  AOI22_X1 U13912 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10860) );
  NAND3_X1 U13913 ( .A1(n10861), .A2(n10860), .A3(n10859), .ZN(n10862) );
  AOI22_X1 U13914 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10876) );
  AOI22_X1 U13915 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10875) );
  AOI22_X1 U13916 ( .A1(n16928), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10866) );
  OAI21_X1 U13917 ( .B1(n10944), .B2(n20846), .A(n10866), .ZN(n10873) );
  AOI22_X1 U13918 ( .A1(n15523), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U13919 ( .A1(n16946), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10870) );
  INV_X2 U13920 ( .A(n9695), .ZN(n16927) );
  AOI22_X1 U13921 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U13922 ( .A1(n16839), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10868) );
  NAND4_X1 U13923 ( .A1(n10871), .A2(n10870), .A3(n10869), .A4(n10868), .ZN(
        n10872) );
  AOI211_X1 U13924 ( .C1(n16911), .C2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n10873), .B(n10872), .ZN(n10874) );
  NAND3_X1 U13925 ( .A1(n10876), .A2(n10875), .A3(n10874), .ZN(n17137) );
  NAND2_X1 U13926 ( .A1(n10913), .A2(n17137), .ZN(n10916) );
  AOI22_X1 U13927 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10887) );
  AOI22_X1 U13928 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n16844), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10886) );
  AOI22_X1 U13929 ( .A1(n16946), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16952), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10878) );
  OAI21_X1 U13930 ( .B1(n11016), .B2(n20770), .A(n10878), .ZN(n10884) );
  AOI22_X1 U13931 ( .A1(n16883), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10882) );
  AOI22_X1 U13932 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10881) );
  AOI22_X1 U13933 ( .A1(n16955), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10880) );
  AOI22_X1 U13934 ( .A1(n16928), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10879) );
  NAND4_X1 U13935 ( .A1(n10882), .A2(n10881), .A3(n10880), .A4(n10879), .ZN(
        n10883) );
  AOI211_X1 U13936 ( .C1(n16962), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n10884), .B(n10883), .ZN(n10885) );
  NOR2_X4 U13937 ( .A1(n16215), .A2(n17126), .ZN(n17431) );
  INV_X1 U13938 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17678) );
  INV_X1 U13939 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17926) );
  NOR2_X1 U13940 ( .A1(n10905), .A2(n10903), .ZN(n10904) );
  AOI22_X1 U13941 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10894) );
  AOI22_X1 U13942 ( .A1(n16839), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10893) );
  AOI22_X1 U13943 ( .A1(n10853), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10889), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10892) );
  AOI22_X1 U13944 ( .A1(n16946), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10890), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10891) );
  AOI22_X1 U13945 ( .A1(n16953), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15510), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10895) );
  OAI21_X1 U13946 ( .B1(n9694), .B2(n16949), .A(n10895), .ZN(n10898) );
  AOI22_X1 U13947 ( .A1(n10852), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10867), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10896) );
  INV_X1 U13948 ( .A(n10896), .ZN(n10897) );
  AOI22_X1 U13949 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10899) );
  NAND3_X1 U13950 ( .A1(n10071), .A2(n10902), .A3(n10901), .ZN(n17642) );
  NOR2_X1 U13951 ( .A1(n17641), .A2(n17635), .ZN(n17634) );
  NOR2_X1 U13952 ( .A1(n10904), .A2(n17634), .ZN(n17622) );
  XNOR2_X1 U13953 ( .A(n10905), .B(n17150), .ZN(n10907) );
  XNOR2_X1 U13954 ( .A(n10907), .B(n10906), .ZN(n17621) );
  NOR2_X1 U13955 ( .A1(n10906), .A2(n10907), .ZN(n10908) );
  XNOR2_X1 U13956 ( .A(n10909), .B(n17143), .ZN(n10910) );
  NOR2_X1 U13957 ( .A1(n10911), .A2(n10910), .ZN(n10912) );
  NOR2_X1 U13958 ( .A1(n17611), .A2(n10912), .ZN(n17602) );
  INV_X1 U13959 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17917) );
  XOR2_X1 U13960 ( .A(n10913), .B(n17137), .Z(n10914) );
  XOR2_X1 U13961 ( .A(n17917), .B(n10914), .Z(n17601) );
  XNOR2_X1 U13962 ( .A(n10916), .B(n17133), .ZN(n17585) );
  INV_X1 U13963 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17902) );
  XNOR2_X1 U13964 ( .A(n10918), .B(n17130), .ZN(n10919) );
  XOR2_X1 U13965 ( .A(n17902), .B(n10919), .Z(n17570) );
  INV_X1 U13966 ( .A(n16215), .ZN(n10920) );
  XNOR2_X1 U13967 ( .A(n9680), .B(n10921), .ZN(n17565) );
  INV_X1 U13968 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17894) );
  NOR2_X1 U13969 ( .A1(n17565), .A2(n17894), .ZN(n17564) );
  NOR2_X1 U13970 ( .A1(n9680), .A2(n10921), .ZN(n10922) );
  INV_X1 U13971 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17881) );
  INV_X1 U13972 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17859) );
  INV_X1 U13973 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17851) );
  NAND2_X1 U13974 ( .A1(n17505), .A2(n17851), .ZN(n17477) );
  NOR2_X1 U13975 ( .A1(n17477), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17450) );
  INV_X1 U13976 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17842) );
  NAND2_X1 U13977 ( .A1(n17450), .A2(n17842), .ZN(n17468) );
  INV_X1 U13978 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17811) );
  INV_X1 U13979 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17804) );
  NAND2_X1 U13980 ( .A1(n17811), .A2(n17804), .ZN(n17796) );
  INV_X1 U13981 ( .A(n10923), .ZN(n10925) );
  NAND2_X1 U13982 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17507) );
  NOR2_X1 U13983 ( .A1(n17507), .A2(n17851), .ZN(n17825) );
  NAND2_X1 U13984 ( .A1(n17825), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17806) );
  INV_X1 U13985 ( .A(n17806), .ZN(n17481) );
  INV_X1 U13986 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17483) );
  NOR2_X1 U13987 ( .A1(n17483), .A2(n17811), .ZN(n17459) );
  NAND2_X1 U13988 ( .A1(n17481), .A2(n17459), .ZN(n17778) );
  NOR2_X1 U13989 ( .A1(n17778), .A2(n17804), .ZN(n17755) );
  NAND2_X1 U13990 ( .A1(n10928), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10927) );
  INV_X1 U13991 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17786) );
  INV_X1 U13992 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17769) );
  NAND2_X1 U13993 ( .A1(n10929), .A2(n10928), .ZN(n17430) );
  NOR2_X1 U13994 ( .A1(n17786), .A2(n17769), .ZN(n17759) );
  NAND2_X1 U13995 ( .A1(n17759), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17715) );
  INV_X1 U13996 ( .A(n17715), .ZN(n17730) );
  NAND2_X1 U13997 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17719) );
  INV_X1 U13998 ( .A(n17719), .ZN(n17732) );
  NAND3_X1 U13999 ( .A1(n17730), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n17732), .ZN(n17717) );
  INV_X1 U14000 ( .A(n17717), .ZN(n17651) );
  NAND2_X1 U14001 ( .A1(n17651), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17672) );
  INV_X1 U14002 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17702) );
  NOR2_X1 U14003 ( .A1(n17672), .A2(n17702), .ZN(n11083) );
  NOR2_X1 U14004 ( .A1(n17431), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17414) );
  INV_X1 U14005 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17401) );
  NAND2_X1 U14006 ( .A1(n17414), .A2(n17401), .ZN(n10930) );
  NOR2_X1 U14007 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n10930), .ZN(
        n17379) );
  INV_X1 U14008 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17718) );
  NAND2_X1 U14009 ( .A1(n17379), .A2(n17718), .ZN(n17363) );
  NAND2_X1 U14010 ( .A1(n10931), .A2(n10081), .ZN(n10932) );
  INV_X1 U14011 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17406) );
  NAND2_X1 U14012 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17732), .ZN(
        n10933) );
  NOR2_X1 U14013 ( .A1(n17406), .A2(n10933), .ZN(n17364) );
  NOR2_X1 U14014 ( .A1(n17314), .A2(n17546), .ZN(n10934) );
  NAND2_X1 U14015 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17653) );
  INV_X1 U14016 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16193) );
  INV_X1 U14017 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n20801) );
  INV_X1 U14018 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16191) );
  AOI22_X1 U14019 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U14020 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U14021 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U14022 ( .A1(n16928), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10940) );
  NAND4_X1 U14023 ( .A1(n10943), .A2(n10942), .A3(n10941), .A4(n10940), .ZN(
        n10950) );
  AOI22_X1 U14024 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10948) );
  AOI22_X1 U14025 ( .A1(n16844), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10947) );
  INV_X2 U14026 ( .A(n10944), .ZN(n16883) );
  AOI22_X1 U14027 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16883), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10946) );
  AOI22_X1 U14028 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16952), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10945) );
  NAND4_X1 U14029 ( .A1(n10948), .A2(n10947), .A3(n10946), .A4(n10945), .ZN(
        n10949) );
  AOI22_X1 U14030 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U14031 ( .A1(n10890), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U14032 ( .A1(n16927), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10951) );
  OAI21_X1 U14033 ( .B1(n10809), .B2(n16949), .A(n10951), .ZN(n10957) );
  AOI22_X1 U14034 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10955) );
  AOI22_X1 U14035 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10954) );
  AOI22_X1 U14036 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16883), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10953) );
  AOI22_X1 U14037 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10952) );
  NAND4_X1 U14038 ( .A1(n10955), .A2(n10954), .A3(n10953), .A4(n10952), .ZN(
        n10956) );
  AOI22_X1 U14039 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16952), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10971) );
  AOI22_X1 U14040 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U14041 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10961) );
  OAI21_X1 U14042 ( .B1(n10962), .B2(n20846), .A(n10961), .ZN(n10968) );
  AOI22_X1 U14043 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10966) );
  AOI22_X1 U14044 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10965) );
  AOI22_X1 U14045 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10964) );
  INV_X2 U14046 ( .A(n16950), .ZN(n16928) );
  AOI22_X1 U14047 ( .A1(n9587), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10963) );
  NAND4_X1 U14048 ( .A1(n10966), .A2(n10965), .A3(n10964), .A4(n10963), .ZN(
        n10967) );
  AOI211_X1 U14049 ( .C1(n16926), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n10968), .B(n10967), .ZN(n10969) );
  NAND3_X1 U14050 ( .A1(n10971), .A2(n10970), .A3(n10969), .ZN(n18003) );
  NOR2_X1 U14051 ( .A1(n17988), .A2(n18003), .ZN(n11000) );
  AOI22_X1 U14052 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10975) );
  AOI22_X1 U14053 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10974) );
  AOI22_X1 U14054 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10973) );
  AOI22_X1 U14055 ( .A1(n16844), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10972) );
  NAND4_X1 U14056 ( .A1(n10975), .A2(n10974), .A3(n10973), .A4(n10972), .ZN(
        n10981) );
  AOI22_X1 U14057 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10979) );
  AOI22_X1 U14058 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10978) );
  AOI22_X1 U14059 ( .A1(n16955), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10977) );
  AOI22_X1 U14060 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10976) );
  NAND4_X1 U14061 ( .A1(n10979), .A2(n10978), .A3(n10977), .A4(n10976), .ZN(
        n10980) );
  AOI22_X1 U14062 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10985) );
  AOI22_X1 U14063 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10984) );
  AOI22_X1 U14064 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10983) );
  AOI22_X1 U14065 ( .A1(n16928), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10982) );
  NAND4_X1 U14066 ( .A1(n10985), .A2(n10984), .A3(n10983), .A4(n10982), .ZN(
        n10991) );
  AOI22_X1 U14067 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10989) );
  AOI22_X1 U14068 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10988) );
  AOI22_X1 U14069 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10987) );
  AOI22_X1 U14070 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10986) );
  NAND4_X1 U14071 ( .A1(n10989), .A2(n10988), .A3(n10987), .A4(n10986), .ZN(
        n10990) );
  NOR2_X1 U14072 ( .A1(n17006), .A2(n18017), .ZN(n11001) );
  AOI22_X1 U14073 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10999) );
  AOI22_X1 U14074 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n16955), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n16910), .ZN(n10998) );
  AOI22_X1 U14075 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10992) );
  OAI21_X1 U14076 ( .B1(n10090), .B2(n20770), .A(n10992), .ZN(n10997) );
  AOI22_X1 U14077 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n15525), .ZN(n10996) );
  AOI22_X1 U14078 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n16927), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n16951), .ZN(n10995) );
  AOI22_X1 U14079 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16911), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U14080 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n16928), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n16883), .ZN(n10993) );
  NAND4_X1 U14081 ( .A1(n11037), .A2(n11000), .A3(n11001), .A4(n17092), .ZN(
        n11036) );
  INV_X1 U14082 ( .A(n11001), .ZN(n11024) );
  AOI22_X1 U14083 ( .A1(n16872), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U14084 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11004) );
  AOI22_X1 U14085 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11003) );
  AOI22_X1 U14086 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11002) );
  NAND4_X1 U14087 ( .A1(n11005), .A2(n11004), .A3(n11003), .A4(n11002), .ZN(
        n11011) );
  AOI22_X1 U14088 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16883), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11009) );
  AOI22_X1 U14089 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11008) );
  AOI22_X1 U14090 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11007) );
  AOI22_X1 U14091 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11006) );
  NAND4_X1 U14092 ( .A1(n11009), .A2(n11008), .A3(n11007), .A4(n11006), .ZN(
        n11010) );
  AOI22_X1 U14093 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11015) );
  AOI22_X1 U14094 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11014) );
  AOI22_X1 U14095 ( .A1(n16883), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11013) );
  AOI22_X1 U14096 ( .A1(n16928), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11012) );
  NAND4_X1 U14097 ( .A1(n11015), .A2(n11014), .A3(n11013), .A4(n11012), .ZN(
        n11022) );
  AOI22_X1 U14098 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11020) );
  AOI22_X1 U14099 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11019) );
  AOI22_X1 U14100 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11018) );
  AOI22_X1 U14101 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11017) );
  NAND4_X1 U14102 ( .A1(n11020), .A2(n11019), .A3(n11018), .A4(n11017), .ZN(
        n11021) );
  NAND2_X1 U14103 ( .A1(n11050), .A2(n11044), .ZN(n11074) );
  AOI21_X1 U14104 ( .B1(n17092), .B2(n11024), .A(n11039), .ZN(n11023) );
  AOI21_X1 U14105 ( .B1(n11024), .B2(n11074), .A(n11023), .ZN(n11033) );
  NAND2_X1 U14106 ( .A1(n18631), .A2(n16646), .ZN(n15590) );
  AND2_X1 U14107 ( .A1(n11044), .A2(n11042), .ZN(n11029) );
  NAND2_X1 U14108 ( .A1(n11039), .A2(n18017), .ZN(n11025) );
  NOR2_X1 U14109 ( .A1(n17006), .A2(n11025), .ZN(n11028) );
  NAND2_X1 U14110 ( .A1(n11050), .A2(n18009), .ZN(n11070) );
  NAND2_X1 U14111 ( .A1(n18631), .A2(n17988), .ZN(n11043) );
  AOI21_X1 U14112 ( .B1(n17092), .B2(n18452), .A(n11043), .ZN(n11071) );
  AOI21_X1 U14113 ( .B1(n11070), .B2(n11041), .A(n11071), .ZN(n11026) );
  NOR2_X1 U14114 ( .A1(n11026), .A2(n11037), .ZN(n11027) );
  NOR2_X1 U14115 ( .A1(n18017), .A2(n11070), .ZN(n11078) );
  OAI21_X1 U14116 ( .B1(n11030), .B2(n11078), .A(n16646), .ZN(n11031) );
  NAND3_X1 U14117 ( .A1(n11033), .A2(n11032), .A3(n11031), .ZN(n11047) );
  NOR2_X1 U14118 ( .A1(n18017), .A2(n18009), .ZN(n11035) );
  NAND2_X1 U14119 ( .A1(n11050), .A2(n11037), .ZN(n18433) );
  INV_X1 U14120 ( .A(n18433), .ZN(n11034) );
  INV_X1 U14121 ( .A(n11037), .ZN(n18000) );
  INV_X1 U14122 ( .A(n11045), .ZN(n11046) );
  OAI211_X1 U14123 ( .C1(n18009), .C2(n18017), .A(n11039), .B(n18452), .ZN(
        n11038) );
  OAI22_X1 U14124 ( .A1(n11039), .A2(n18452), .B1(n16646), .B2(n11038), .ZN(
        n11040) );
  NAND2_X1 U14125 ( .A1(n11044), .A2(n11043), .ZN(n18645) );
  NAND2_X1 U14126 ( .A1(n18017), .A2(n18003), .ZN(n18434) );
  NOR2_X1 U14127 ( .A1(n18631), .A2(n11046), .ZN(n11048) );
  XNOR2_X1 U14128 ( .A(n17991), .B(n11050), .ZN(n11069) );
  INV_X1 U14129 ( .A(n16213), .ZN(n18422) );
  AOI22_X1 U14130 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18463), .B2(n11052), .ZN(
        n11054) );
  XNOR2_X1 U14131 ( .A(n11053), .B(n11054), .ZN(n11067) );
  OAI22_X1 U14132 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18467), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11056), .ZN(n11060) );
  NOR2_X1 U14133 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18467), .ZN(
        n11057) );
  NAND2_X1 U14134 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11056), .ZN(
        n11059) );
  AOI22_X1 U14135 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11060), .B1(
        n11057), .B2(n11059), .ZN(n11063) );
  OAI211_X1 U14136 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18272), .A(
        n11063), .B(n11058), .ZN(n11076) );
  XOR2_X1 U14137 ( .A(n11077), .B(n11058), .Z(n11066) );
  OAI22_X1 U14138 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18478), .B1(
        n11061), .B2(n11060), .ZN(n11065) );
  INV_X1 U14139 ( .A(n11067), .ZN(n11062) );
  AOI21_X1 U14140 ( .B1(n11063), .B2(n11062), .A(n11065), .ZN(n11075) );
  INV_X1 U14141 ( .A(n11075), .ZN(n11064) );
  OAI21_X1 U14142 ( .B1(n11067), .B2(n11076), .A(n16317), .ZN(n18421) );
  NOR4_X1 U14143 ( .A1(n18631), .A2(n18017), .A3(n18421), .A4(n17995), .ZN(
        n11082) );
  NAND2_X1 U14144 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18509), .ZN(n18641) );
  INV_X2 U14145 ( .A(n18641), .ZN(n18640) );
  NAND2_X1 U14146 ( .A1(n18640), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18575) );
  NOR2_X1 U14147 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18496) );
  INV_X1 U14148 ( .A(n18496), .ZN(n11068) );
  NAND3_X1 U14149 ( .A1(n18509), .A2(n18568), .A3(n11068), .ZN(n18629) );
  INV_X1 U14150 ( .A(n18629), .ZN(n13968) );
  NAND2_X1 U14151 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18632) );
  OAI21_X1 U14152 ( .B1(n13968), .B2(n11069), .A(n18632), .ZN(n16316) );
  NAND2_X1 U14153 ( .A1(n16317), .A2(n11070), .ZN(n11080) );
  AOI221_X1 U14154 ( .B1(n11074), .B2(n11073), .C1(n11072), .C2(n11073), .A(
        n11071), .ZN(n13973) );
  OAI21_X1 U14155 ( .B1(n11077), .B2(n11076), .A(n11075), .ZN(n12191) );
  OAI21_X1 U14156 ( .B1(n11078), .B2(n18003), .A(n18428), .ZN(n11079) );
  OAI211_X1 U14157 ( .C1(n16316), .C2(n11080), .A(n13973), .B(n11079), .ZN(
        n11081) );
  NOR2_X1 U14158 ( .A1(n18646), .A2(n18486), .ZN(n18626) );
  NAND2_X1 U14159 ( .A1(n18605), .A2(n18626), .ZN(n18490) );
  OAI21_X2 U14160 ( .B1(n11082), .B2(n11081), .A(n18483), .ZN(n17952) );
  NAND3_X1 U14161 ( .A1(n16208), .A2(n18422), .A3(n17961), .ZN(n17891) );
  NAND2_X1 U14162 ( .A1(n16190), .A2(n17872), .ZN(n11124) );
  INV_X1 U14163 ( .A(n17755), .ZN(n17429) );
  INV_X1 U14164 ( .A(n11083), .ZN(n17336) );
  NAND2_X1 U14165 ( .A1(n17690), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17324) );
  NAND2_X1 U14166 ( .A1(n17323), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17273) );
  NAND2_X1 U14167 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11110) );
  NOR2_X1 U14168 ( .A1(n17273), .A2(n11110), .ZN(n16210) );
  INV_X1 U14169 ( .A(n16210), .ZN(n16194) );
  NAND2_X1 U14170 ( .A1(n18422), .A2(n17961), .ZN(n17967) );
  NOR2_X1 U14171 ( .A1(n16208), .A2(n17967), .ZN(n17816) );
  NAND2_X1 U14172 ( .A1(n17789), .A2(n17961), .ZN(n17969) );
  INV_X1 U14173 ( .A(n17969), .ZN(n17951) );
  INV_X1 U14174 ( .A(n10905), .ZN(n11084) );
  INV_X1 U14175 ( .A(n17642), .ZN(n15595) );
  NOR2_X1 U14176 ( .A1(n11092), .A2(n17150), .ZN(n11087) );
  NOR2_X1 U14177 ( .A1(n17143), .A2(n11087), .ZN(n11095) );
  NAND2_X1 U14178 ( .A1(n11095), .A2(n17137), .ZN(n11086) );
  NOR2_X1 U14179 ( .A1(n17133), .A2(n11086), .ZN(n11099) );
  NAND2_X1 U14180 ( .A1(n11099), .A2(n11100), .ZN(n11085) );
  NOR2_X1 U14181 ( .A1(n17126), .A2(n11085), .ZN(n11108) );
  XOR2_X1 U14182 ( .A(n17126), .B(n11085), .Z(n17557) );
  XOR2_X1 U14183 ( .A(n17133), .B(n11086), .Z(n17582) );
  XOR2_X1 U14184 ( .A(n17143), .B(n11087), .Z(n11088) );
  NAND2_X1 U14185 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11088), .ZN(
        n11094) );
  XOR2_X1 U14186 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n11088), .Z(
        n17610) );
  AOI21_X1 U14187 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10905), .A(
        n17642), .ZN(n11090) );
  INV_X1 U14188 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17960) );
  NOR2_X1 U14189 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n10905), .ZN(
        n11089) );
  AOI221_X1 U14190 ( .B1(n17642), .B2(n10905), .C1(n11090), .C2(n17960), .A(
        n11089), .ZN(n11091) );
  NAND2_X1 U14191 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n9589), .ZN(
        n11093) );
  XOR2_X1 U14192 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n9589), .Z(n17625) );
  XNOR2_X1 U14193 ( .A(n17150), .B(n11092), .ZN(n17624) );
  NAND2_X1 U14194 ( .A1(n17625), .A2(n17624), .ZN(n17623) );
  NAND2_X1 U14195 ( .A1(n11093), .A2(n17623), .ZN(n17609) );
  NAND2_X1 U14196 ( .A1(n17610), .A2(n17609), .ZN(n17608) );
  NAND2_X1 U14197 ( .A1(n11094), .A2(n17608), .ZN(n11096) );
  NOR2_X1 U14198 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11096), .ZN(
        n11097) );
  XOR2_X1 U14199 ( .A(n17137), .B(n11095), .Z(n17596) );
  XOR2_X1 U14200 ( .A(n17917), .B(n11096), .Z(n17595) );
  NOR2_X2 U14201 ( .A1(n11097), .A2(n17594), .ZN(n17581) );
  NAND2_X1 U14202 ( .A1(n17582), .A2(n17581), .ZN(n17580) );
  NOR2_X1 U14203 ( .A1(n17582), .A2(n17581), .ZN(n11098) );
  XOR2_X1 U14204 ( .A(n11100), .B(n11099), .Z(n11102) );
  NAND2_X1 U14205 ( .A1(n11101), .A2(n11102), .ZN(n11103) );
  XOR2_X1 U14206 ( .A(n11102), .B(n11101), .Z(n17574) );
  NAND2_X1 U14207 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17574), .ZN(
        n17573) );
  NOR2_X2 U14208 ( .A1(n11104), .A2(n17894), .ZN(n11105) );
  NAND2_X1 U14209 ( .A1(n11108), .A2(n11105), .ZN(n11109) );
  INV_X1 U14210 ( .A(n11105), .ZN(n11107) );
  NAND2_X1 U14211 ( .A1(n17557), .A2(n17558), .ZN(n17556) );
  NAND2_X1 U14212 ( .A1(n11108), .A2(n11107), .ZN(n11106) );
  OAI211_X1 U14213 ( .C1(n11108), .C2(n11107), .A(n17556), .B(n11106), .ZN(
        n17548) );
  NAND2_X1 U14214 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17548), .ZN(
        n17547) );
  INV_X1 U14215 ( .A(n17672), .ZN(n17271) );
  INV_X1 U14216 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17666) );
  NAND2_X1 U14217 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17679) );
  INV_X1 U14218 ( .A(n17679), .ZN(n17673) );
  NAND2_X1 U14219 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17673), .ZN(
        n17667) );
  NOR2_X1 U14220 ( .A1(n17666), .A2(n17667), .ZN(n11112) );
  NAND2_X1 U14221 ( .A1(n17271), .A2(n11112), .ZN(n17649) );
  NOR2_X1 U14222 ( .A1(n11110), .A2(n17658), .ZN(n16209) );
  NAND3_X1 U14223 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17795) );
  NOR3_X1 U14224 ( .A1(n17917), .A2(n17926), .A3(n10917), .ZN(n17753) );
  AOI21_X1 U14225 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17915) );
  INV_X1 U14226 ( .A(n17915), .ZN(n17936) );
  NAND2_X1 U14227 ( .A1(n17753), .A2(n17936), .ZN(n17878) );
  NOR2_X1 U14228 ( .A1(n17795), .A2(n17878), .ZN(n17776) );
  NAND2_X1 U14229 ( .A1(n17755), .A2(n17776), .ZN(n17757) );
  AOI21_X1 U14230 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18438), .A(
        n18437), .ZN(n17937) );
  NAND2_X1 U14231 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17914) );
  INV_X1 U14232 ( .A(n17914), .ZN(n11111) );
  NAND2_X1 U14233 ( .A1(n11111), .A2(n17753), .ZN(n17877) );
  NOR2_X1 U14234 ( .A1(n17877), .A2(n17795), .ZN(n17777) );
  NAND2_X1 U14235 ( .A1(n17755), .A2(n17777), .ZN(n17711) );
  OAI22_X1 U14236 ( .A1(n18427), .A2(n17757), .B1(n17937), .B2(n17711), .ZN(
        n16218) );
  NAND2_X1 U14237 ( .A1(n17271), .A2(n16218), .ZN(n17677) );
  NAND2_X1 U14238 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n11112), .ZN(
        n17272) );
  NOR4_X1 U14239 ( .A1(n20801), .A2(n17952), .A3(n17677), .A4(n17272), .ZN(
        n11140) );
  AOI21_X1 U14240 ( .B1(n17951), .B2(n16209), .A(n11140), .ZN(n11113) );
  OAI21_X1 U14241 ( .B1(n16194), .B2(n17885), .A(n11113), .ZN(n15542) );
  NAND2_X1 U14242 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15542), .ZN(
        n11121) );
  NOR2_X1 U14243 ( .A1(n17880), .A2(n17952), .ZN(n17955) );
  NAND3_X1 U14244 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16185) );
  NOR2_X1 U14245 ( .A1(n17273), .A2(n16185), .ZN(n16184) );
  OAI21_X1 U14246 ( .B1(n16185), .B2(n17658), .A(n17951), .ZN(n11117) );
  NAND2_X1 U14247 ( .A1(n18605), .A2(n18586), .ZN(n18593) );
  NOR3_X1 U14248 ( .A1(n18593), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(
        P3_STATE2_REG_0__SCAN_IN), .ZN(n11114) );
  INV_X2 U14249 ( .A(n11114), .ZN(n17963) );
  INV_X2 U14250 ( .A(n17963), .ZN(n17965) );
  OAI21_X1 U14251 ( .B1(n17649), .B2(n17757), .A(n18449), .ZN(n17654) );
  NAND2_X1 U14252 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17777), .ZN(
        n17866) );
  NOR2_X1 U14253 ( .A1(n17429), .A2(n17866), .ZN(n17780) );
  NAND2_X1 U14254 ( .A1(n17271), .A2(n17780), .ZN(n17650) );
  OAI21_X1 U14255 ( .B1(n17272), .B2(n17650), .A(n18438), .ZN(n11116) );
  OAI21_X1 U14256 ( .B1(n17649), .B2(n17711), .A(n18437), .ZN(n11115) );
  NAND4_X1 U14257 ( .A1(n17925), .A2(n17654), .A3(n11116), .A4(n11115), .ZN(
        n16212) );
  NAND2_X1 U14258 ( .A1(n17963), .A2(n16212), .ZN(n11138) );
  OAI211_X1 U14259 ( .C1(n16184), .C2(n17885), .A(n11117), .B(n11138), .ZN(
        n15538) );
  AOI21_X1 U14260 ( .B1(n17955), .B2(n16185), .A(n15538), .ZN(n11118) );
  NAND2_X1 U14261 ( .A1(n17965), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n11119) );
  INV_X1 U14262 ( .A(n11122), .ZN(n11123) );
  NAND2_X1 U14263 ( .A1(n11124), .A2(n11123), .ZN(P3_U2832) );
  NOR2_X1 U14264 ( .A1(n17431), .A2(n11125), .ZN(n11130) );
  INV_X1 U14265 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18591) );
  AND2_X1 U14266 ( .A1(n18591), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11126) );
  NOR2_X1 U14267 ( .A1(n11130), .A2(n11126), .ZN(n11128) );
  AOI22_X1 U14268 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16191), .B1(
        n11128), .B2(n11127), .ZN(n11133) );
  AOI22_X1 U14269 ( .A1(n17431), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n18591), .B2(n17546), .ZN(n11132) );
  OAI21_X1 U14270 ( .B1(n11130), .B2(n11129), .A(n11132), .ZN(n11131) );
  OAI21_X1 U14271 ( .B1(n11133), .B2(n11132), .A(n11131), .ZN(n12192) );
  NAND2_X1 U14272 ( .A1(n12192), .A2(n17872), .ZN(n11147) );
  OR3_X1 U14273 ( .A1(n16185), .A2(n17658), .A3(n16191), .ZN(n11134) );
  XOR2_X1 U14274 ( .A(n11134), .B(n18591), .Z(n12203) );
  INV_X1 U14275 ( .A(n12203), .ZN(n11135) );
  NOR3_X1 U14276 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16193), .A3(
        n16191), .ZN(n11141) );
  NAND2_X1 U14277 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16184), .ZN(
        n11136) );
  AOI22_X1 U14278 ( .A1(n16210), .A2(n11141), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n11136), .ZN(n12193) );
  OR2_X1 U14279 ( .A1(n12193), .A2(n17885), .ZN(n11143) );
  INV_X1 U14280 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18572) );
  NOR2_X1 U14281 ( .A1(n17963), .A2(n18572), .ZN(n12199) );
  OAI21_X1 U14282 ( .B1(n16191), .B2(n16185), .A(n17955), .ZN(n11137) );
  AOI21_X1 U14283 ( .B1(n11138), .B2(n11137), .A(n18591), .ZN(n11139) );
  AOI211_X1 U14284 ( .C1(n11141), .C2(n11140), .A(n12199), .B(n11139), .ZN(
        n11142) );
  NAND2_X1 U14285 ( .A1(n11143), .A2(n11142), .ZN(n11144) );
  NAND2_X1 U14286 ( .A1(n11147), .A2(n11146), .ZN(P3_U2831) );
  AOI22_X1 U14287 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9650), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11152) );
  AOI22_X1 U14288 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11151) );
  AOI22_X1 U14289 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9671), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11150) );
  AND2_X2 U14290 ( .A1(n13430), .A2(n13638), .ZN(n11311) );
  AOI22_X1 U14291 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11311), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11149) );
  AOI22_X1 U14292 ( .A1(n11195), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11162) );
  AOI22_X1 U14293 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12130), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11161) );
  AOI22_X1 U14294 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11458), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11160) );
  AND2_X4 U14295 ( .A1(n13433), .A2(n11158), .ZN(n11373) );
  AOI22_X1 U14296 ( .A1(n11453), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11159) );
  NAND2_X1 U14297 ( .A1(n11195), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11167) );
  NAND2_X1 U14298 ( .A1(n11453), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11166) );
  NAND2_X1 U14299 ( .A1(n11373), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11165) );
  NAND2_X1 U14300 ( .A1(n12111), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11164) );
  NAND2_X1 U14301 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11171) );
  NAND2_X1 U14302 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11170) );
  NAND2_X1 U14303 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11169) );
  NAND2_X1 U14304 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11168) );
  NAND2_X1 U14305 ( .A1(n9651), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11175) );
  NAND2_X1 U14306 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11174) );
  NAND2_X1 U14307 ( .A1(n11336), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11173) );
  NAND2_X1 U14308 ( .A1(n11258), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11172) );
  NAND2_X1 U14309 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11179) );
  NAND2_X1 U14310 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11178) );
  NAND2_X1 U14311 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11177) );
  NAND2_X1 U14312 ( .A1(n11311), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11176) );
  AOI22_X1 U14313 ( .A1(n9651), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11188) );
  AOI22_X1 U14314 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9671), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11187) );
  AOI22_X1 U14315 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11311), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11185) );
  AOI22_X1 U14316 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11458), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11184) );
  AND2_X1 U14317 ( .A1(n11185), .A2(n11184), .ZN(n11186) );
  AOI22_X1 U14318 ( .A1(n11453), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11192) );
  AOI22_X1 U14319 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11191) );
  AOI22_X1 U14320 ( .A1(n11195), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11190) );
  AOI22_X1 U14321 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11189) );
  AOI22_X1 U14322 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11194), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11199) );
  AOI22_X1 U14323 ( .A1(n11453), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11198) );
  AOI22_X1 U14324 ( .A1(n11195), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11197) );
  AOI22_X1 U14325 ( .A1(n11336), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11196) );
  AOI22_X1 U14326 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11458), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11205) );
  AOI22_X1 U14327 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12135), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11204) );
  AOI22_X1 U14328 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11203) );
  AOI22_X1 U14329 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11311), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11202) );
  NAND2_X1 U14330 ( .A1(n11290), .A2(n11206), .ZN(n11280) );
  AOI22_X1 U14331 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11210) );
  AOI22_X1 U14332 ( .A1(n11195), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11209) );
  AOI22_X1 U14333 ( .A1(n11453), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11208) );
  AOI22_X1 U14334 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11207) );
  NAND4_X1 U14335 ( .A1(n11210), .A2(n11209), .A3(n11208), .A4(n11207), .ZN(
        n11219) );
  INV_X1 U14336 ( .A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11212) );
  INV_X1 U14337 ( .A(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11211) );
  OAI22_X1 U14338 ( .A1(n11428), .A2(n11212), .B1(n9666), .B2(n11211), .ZN(
        n11213) );
  INV_X1 U14339 ( .A(n11213), .ZN(n11217) );
  AOI22_X1 U14340 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11458), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11216) );
  AOI22_X1 U14341 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11201), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11215) );
  AOI22_X1 U14342 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11311), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11214) );
  NAND4_X1 U14343 ( .A1(n11217), .A2(n11216), .A3(n11215), .A4(n11214), .ZN(
        n11218) );
  OR2_X2 U14344 ( .A1(n11219), .A2(n11218), .ZN(n20025) );
  NAND2_X1 U14345 ( .A1(n11280), .A2(n20025), .ZN(n11239) );
  AOI22_X1 U14346 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11223) );
  AOI22_X1 U14347 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11222) );
  AOI22_X1 U14348 ( .A1(n11453), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11221) );
  AOI22_X1 U14349 ( .A1(n11195), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11220) );
  AOI22_X1 U14350 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11230) );
  AOI22_X1 U14351 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11458), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11229) );
  INV_X1 U14352 ( .A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11225) );
  INV_X1 U14353 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11224) );
  OAI22_X1 U14354 ( .A1(n11428), .A2(n11225), .B1(n9665), .B2(n11224), .ZN(
        n11226) );
  INV_X1 U14355 ( .A(n11226), .ZN(n11228) );
  AOI22_X1 U14356 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11311), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11227) );
  NAND2_X1 U14357 ( .A1(n10077), .A2(n10096), .ZN(n11236) );
  INV_X1 U14358 ( .A(n11267), .ZN(n13236) );
  NAND3_X1 U14359 ( .A1(n11239), .A2(n11238), .A3(n11237), .ZN(n11277) );
  AOI22_X1 U14360 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11244) );
  AOI22_X1 U14361 ( .A1(n11453), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11243) );
  AOI22_X1 U14362 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11242) );
  AOI22_X1 U14363 ( .A1(n11195), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11241) );
  OAI22_X1 U14364 ( .A1(n11428), .A2(n11246), .B1(n9665), .B2(n11245), .ZN(
        n11247) );
  INV_X1 U14365 ( .A(n11247), .ZN(n11251) );
  AOI22_X1 U14366 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11311), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11250) );
  AOI22_X1 U14367 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11458), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11249) );
  AOI22_X1 U14368 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11201), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11248) );
  AOI22_X1 U14369 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11257) );
  AOI22_X1 U14370 ( .A1(n12135), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11256) );
  AOI22_X1 U14371 ( .A1(n11453), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11255) );
  AOI22_X1 U14372 ( .A1(n11195), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11254) );
  NAND4_X1 U14373 ( .A1(n11257), .A2(n11256), .A3(n11255), .A4(n11254), .ZN(
        n11264) );
  AOI22_X1 U14374 ( .A1(n9651), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11201), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11262) );
  AOI22_X1 U14375 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11458), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11261) );
  AOI22_X1 U14376 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11260) );
  AOI22_X1 U14377 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11311), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11259) );
  NAND4_X1 U14378 ( .A1(n11262), .A2(n11261), .A3(n11260), .A4(n11259), .ZN(
        n11263) );
  NAND3_X1 U14379 ( .A1(n12030), .A2(n11293), .A3(n11235), .ZN(n11266) );
  AND2_X2 U14380 ( .A1(n11930), .A2(n20005), .ZN(n13266) );
  NAND2_X1 U14381 ( .A1(n13378), .A2(n13266), .ZN(n12158) );
  INV_X1 U14382 ( .A(n11289), .ZN(n11269) );
  NAND2_X1 U14383 ( .A1(n11279), .A2(n12030), .ZN(n12172) );
  NAND2_X1 U14384 ( .A1(n11269), .A2(n11268), .ZN(n13425) );
  NAND2_X1 U14385 ( .A1(n11231), .A2(n11267), .ZN(n13379) );
  INV_X1 U14386 ( .A(n13409), .ZN(n13415) );
  NAND2_X1 U14387 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20589) );
  OAI21_X1 U14388 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(n20589), .ZN(n13184) );
  INV_X1 U14389 ( .A(n13184), .ZN(n11272) );
  OAI22_X1 U14390 ( .A1(n13416), .A2(n11295), .B1(n11275), .B2(n13265), .ZN(
        n11276) );
  MUX2_X1 U14391 ( .A(n11930), .B(n11236), .S(n20005), .Z(n13396) );
  NOR2_X1 U14392 ( .A1(n11276), .A2(n13396), .ZN(n11278) );
  NAND2_X1 U14393 ( .A1(n11277), .A2(n11270), .ZN(n13401) );
  INV_X1 U14394 ( .A(n11279), .ZN(n11283) );
  NAND2_X1 U14395 ( .A1(n12030), .A2(n11231), .ZN(n11281) );
  NAND2_X1 U14396 ( .A1(n15908), .A2(n20578), .ZN(n12072) );
  NAND2_X1 U14397 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11363) );
  OAI21_X1 U14398 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11363), .ZN(n20332) );
  OR2_X1 U14399 ( .A1(n15577), .A2(n20327), .ZN(n11358) );
  OAI21_X1 U14400 ( .B1(n12072), .B2(n20332), .A(n11358), .ZN(n11285) );
  INV_X1 U14401 ( .A(n11285), .ZN(n11286) );
  NAND2_X1 U14402 ( .A1(n9659), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11288) );
  MUX2_X1 U14403 ( .A(n15577), .B(n12072), .S(n20665), .Z(n11345) );
  AND2_X1 U14404 ( .A1(n13593), .A2(n14089), .ZN(n13177) );
  INV_X1 U14405 ( .A(n11290), .ZN(n11291) );
  NAND2_X1 U14406 ( .A1(n11291), .A2(n20025), .ZN(n11292) );
  NAND2_X1 U14407 ( .A1(n13177), .A2(n11292), .ZN(n11299) );
  INV_X1 U14408 ( .A(n15908), .ZN(n20651) );
  NOR2_X1 U14409 ( .A1(n20651), .A2(n20578), .ZN(n11298) );
  NAND2_X1 U14410 ( .A1(n11279), .A2(n13186), .ZN(n13403) );
  INV_X1 U14411 ( .A(n11294), .ZN(n11296) );
  NAND2_X1 U14412 ( .A1(n11296), .A2(n15572), .ZN(n11297) );
  OAI211_X1 U14413 ( .C1(n9592), .C2(n11302), .A(n11301), .B(n11300), .ZN(
        n11403) );
  INV_X1 U14414 ( .A(n11304), .ZN(n11303) );
  AOI22_X1 U14416 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11309) );
  AOI22_X1 U14417 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11308) );
  AOI22_X1 U14418 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11307) );
  AOI22_X1 U14419 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11306) );
  NAND4_X1 U14420 ( .A1(n11309), .A2(n11308), .A3(n11307), .A4(n11306), .ZN(
        n11317) );
  AOI22_X1 U14421 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11315) );
  AOI22_X1 U14422 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11314) );
  AOI22_X1 U14423 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11313) );
  AOI22_X1 U14424 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11312) );
  NAND4_X1 U14425 ( .A1(n11315), .A2(n11314), .A3(n11313), .A4(n11312), .ZN(
        n11316) );
  INV_X1 U14426 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U14427 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U14428 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11323) );
  AOI22_X1 U14429 ( .A1(n11319), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11201), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11322) );
  INV_X1 U14430 ( .A(n11320), .ZN(n11331) );
  AOI22_X1 U14431 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11321) );
  NAND4_X1 U14432 ( .A1(n11324), .A2(n11323), .A3(n11322), .A4(n11321), .ZN(
        n11330) );
  AOI22_X1 U14433 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11328) );
  AOI22_X1 U14434 ( .A1(n11195), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11327) );
  AOI22_X1 U14435 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14436 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11325) );
  NAND4_X1 U14437 ( .A1(n11328), .A2(n11327), .A3(n11326), .A4(n11325), .ZN(
        n11329) );
  AOI21_X1 U14438 ( .B1(n13416), .B2(n11986), .A(n20578), .ZN(n11344) );
  AOI22_X1 U14439 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11335) );
  AOI22_X1 U14440 ( .A1(n9651), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11334) );
  AOI22_X1 U14441 ( .A1(n11319), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9671), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14442 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11311), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11332) );
  NAND4_X1 U14443 ( .A1(n11335), .A2(n11334), .A3(n11333), .A4(n11332), .ZN(
        n11342) );
  AOI22_X1 U14444 ( .A1(n12135), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11340) );
  AOI22_X1 U14445 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11339) );
  AOI22_X1 U14446 ( .A1(n11195), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11338) );
  AOI22_X1 U14447 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11337) );
  NAND4_X1 U14448 ( .A1(n11340), .A2(n11339), .A3(n11338), .A4(n11337), .ZN(
        n11341) );
  NAND2_X1 U14449 ( .A1(n11270), .A2(n11941), .ZN(n11343) );
  OAI211_X1 U14450 ( .C1(n12053), .C2(n11673), .A(n11344), .B(n11343), .ZN(
        n11412) );
  NAND2_X1 U14451 ( .A1(n11345), .A2(n20578), .ZN(n11348) );
  INV_X1 U14452 ( .A(n11986), .ZN(n11994) );
  INV_X1 U14453 ( .A(n11941), .ZN(n11346) );
  MUX2_X1 U14454 ( .A(n11353), .B(n11991), .S(n11346), .Z(n11347) );
  NAND2_X1 U14455 ( .A1(n11412), .A2(n11411), .ZN(n11349) );
  NAND2_X1 U14456 ( .A1(n11349), .A2(n11991), .ZN(n11356) );
  OR2_X1 U14457 ( .A1(n11420), .A2(n11350), .ZN(n11352) );
  NAND2_X1 U14458 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11351) );
  INV_X1 U14459 ( .A(n11354), .ZN(n11355) );
  AND2_X1 U14461 ( .A1(n11358), .A2(n11153), .ZN(n11359) );
  NOR2_X1 U14462 ( .A1(n15577), .A2(n20407), .ZN(n11361) );
  INV_X1 U14463 ( .A(n12072), .ZN(n11365) );
  INV_X1 U14464 ( .A(n11363), .ZN(n11362) );
  NAND2_X1 U14465 ( .A1(n11362), .A2(n20407), .ZN(n20376) );
  NAND2_X1 U14466 ( .A1(n11363), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11364) );
  NAND2_X1 U14467 ( .A1(n20376), .A2(n11364), .ZN(n20012) );
  NAND2_X1 U14468 ( .A1(n11365), .A2(n20012), .ZN(n11368) );
  NAND2_X1 U14469 ( .A1(n11370), .A2(n11368), .ZN(n11366) );
  NAND4_X1 U14470 ( .A1(n11371), .A2(n11370), .A3(n11369), .A4(n11368), .ZN(
        n11372) );
  AOI22_X1 U14471 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11377) );
  AOI22_X1 U14472 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11376) );
  AOI22_X1 U14473 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11375) );
  AOI22_X1 U14474 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11374) );
  NAND4_X1 U14475 ( .A1(n11377), .A2(n11376), .A3(n11375), .A4(n11374), .ZN(
        n11386) );
  INV_X1 U14476 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11379) );
  INV_X1 U14477 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11378) );
  OAI22_X1 U14478 ( .A1(n11911), .A2(n11379), .B1(n9666), .B2(n11378), .ZN(
        n11380) );
  INV_X1 U14479 ( .A(n11380), .ZN(n11384) );
  AOI22_X1 U14480 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14481 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11201), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11382) );
  AOI22_X1 U14482 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11381) );
  NAND4_X1 U14483 ( .A1(n11384), .A2(n11383), .A3(n11382), .A4(n11381), .ZN(
        n11385) );
  INV_X1 U14484 ( .A(n11420), .ZN(n11388) );
  AOI22_X1 U14485 ( .A1(n11388), .A2(n11387), .B1(n12057), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11389) );
  INV_X1 U14486 ( .A(n13379), .ZN(n11392) );
  NAND2_X1 U14487 ( .A1(n11392), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11470) );
  NAND2_X1 U14488 ( .A1(n20581), .A2(n20468), .ZN(n11471) );
  XNOR2_X1 U14489 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13612) );
  AOI21_X1 U14490 ( .B1(n12150), .B2(n13612), .A(n12154), .ZN(n11394) );
  NAND2_X1 U14491 ( .A1(n11447), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11393) );
  OAI211_X1 U14492 ( .C1(n11470), .C2(n13431), .A(n11394), .B(n11393), .ZN(
        n11395) );
  INV_X1 U14493 ( .A(n11395), .ZN(n11396) );
  NAND2_X1 U14494 ( .A1(n12154), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11415) );
  AOI22_X1 U14495 ( .A1(n11447), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20581), .ZN(n11400) );
  INV_X1 U14496 ( .A(n11470), .ZN(n11406) );
  NAND2_X1 U14497 ( .A1(n11406), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11399) );
  AND2_X1 U14498 ( .A1(n11400), .A2(n11399), .ZN(n11401) );
  NAND2_X1 U14499 ( .A1(n11402), .A2(n11401), .ZN(n13264) );
  INV_X1 U14500 ( .A(n11403), .ZN(n11404) );
  XNOR2_X1 U14501 ( .A(n11405), .B(n11404), .ZN(n20660) );
  NAND2_X1 U14502 ( .A1(n20660), .A2(n11625), .ZN(n11410) );
  AOI22_X1 U14503 ( .A1(n11447), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20581), .ZN(n11408) );
  NAND2_X1 U14504 ( .A1(n11406), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11407) );
  AND2_X1 U14505 ( .A1(n11408), .A2(n11407), .ZN(n11409) );
  NAND2_X1 U14506 ( .A1(n11410), .A2(n11409), .ZN(n13226) );
  XNOR2_X1 U14507 ( .A(n11412), .B(n11411), .ZN(n20078) );
  AOI21_X1 U14508 ( .B1(n20078), .B2(n13186), .A(n20581), .ZN(n13225) );
  NAND2_X1 U14509 ( .A1(n13226), .A2(n13225), .ZN(n13224) );
  OR2_X1 U14510 ( .A1(n13226), .A2(n11471), .ZN(n11413) );
  NAND2_X1 U14511 ( .A1(n13224), .A2(n11413), .ZN(n13263) );
  INV_X1 U14512 ( .A(n13340), .ZN(n11414) );
  NAND2_X1 U14513 ( .A1(n9689), .A2(n11414), .ZN(n13341) );
  NAND2_X1 U14514 ( .A1(n13341), .A2(n11415), .ZN(n13529) );
  NAND2_X1 U14515 ( .A1(n9659), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11419) );
  NAND3_X1 U14516 ( .A1(n20406), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20243) );
  NOR3_X1 U14517 ( .A1(n20406), .A2(n20407), .A3(n20327), .ZN(n20525) );
  INV_X1 U14518 ( .A(n20525), .ZN(n20516) );
  INV_X1 U14519 ( .A(n20566), .ZN(n20514) );
  OAI21_X1 U14520 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20265), .A(
        n20514), .ZN(n20273) );
  OAI22_X1 U14521 ( .A1(n12072), .A2(n20273), .B1(n15577), .B2(n20406), .ZN(
        n11417) );
  INV_X1 U14522 ( .A(n11417), .ZN(n11418) );
  AOI22_X1 U14523 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U14524 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U14525 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14526 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11422) );
  NAND4_X1 U14527 ( .A1(n11425), .A2(n11424), .A3(n11423), .A4(n11422), .ZN(
        n11435) );
  INV_X1 U14528 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11427) );
  INV_X1 U14529 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11426) );
  OAI22_X1 U14530 ( .A1(n11428), .A2(n11427), .B1(n9665), .B2(n11426), .ZN(
        n11429) );
  INV_X1 U14531 ( .A(n11429), .ZN(n11433) );
  AOI22_X1 U14532 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11432) );
  AOI22_X1 U14533 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U14534 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11430) );
  NAND4_X1 U14535 ( .A1(n11433), .A2(n11432), .A3(n11431), .A4(n11430), .ZN(
        n11434) );
  AOI22_X1 U14536 ( .A1(n12034), .A2(n11966), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n12057), .ZN(n11436) );
  NAND2_X1 U14537 ( .A1(n11439), .A2(n9591), .ZN(n11440) );
  INV_X1 U14538 ( .A(n20004), .ZN(n11441) );
  NAND2_X1 U14539 ( .A1(n11441), .A2(n11625), .ZN(n11452) );
  INV_X1 U14540 ( .A(n11443), .ZN(n11442) );
  INV_X1 U14541 ( .A(n11473), .ZN(n11446) );
  INV_X1 U14542 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11444) );
  NAND2_X1 U14543 ( .A1(n11444), .A2(n11443), .ZN(n11445) );
  NAND2_X1 U14544 ( .A1(n11446), .A2(n11445), .ZN(n13687) );
  AOI22_X1 U14545 ( .A1(n13687), .A2(n12150), .B1(n12154), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11449) );
  NAND2_X1 U14546 ( .A1(n12155), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11448) );
  OAI211_X1 U14547 ( .C1(n11470), .C2(n10048), .A(n11449), .B(n11448), .ZN(
        n11450) );
  INV_X1 U14548 ( .A(n11450), .ZN(n11451) );
  NAND2_X1 U14549 ( .A1(n11452), .A2(n11451), .ZN(n13530) );
  AOI22_X1 U14550 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12130), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11457) );
  AOI22_X1 U14551 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11456) );
  AOI22_X1 U14552 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11455) );
  AOI22_X1 U14553 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11336), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11454) );
  NAND4_X1 U14554 ( .A1(n11457), .A2(n11456), .A3(n11455), .A4(n11454), .ZN(
        n11464) );
  AOI22_X1 U14555 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12135), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U14556 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9671), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11461) );
  AOI22_X1 U14557 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12112), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14558 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11459) );
  NAND4_X1 U14559 ( .A1(n11462), .A2(n11461), .A3(n11460), .A4(n11459), .ZN(
        n11463) );
  NAND2_X1 U14560 ( .A1(n12034), .A2(n11965), .ZN(n11466) );
  NAND2_X1 U14561 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11465) );
  NAND2_X1 U14562 ( .A1(n11466), .A2(n11465), .ZN(n11478) );
  INV_X1 U14563 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n11469) );
  NAND2_X1 U14564 ( .A1(n20581), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11468) );
  NAND2_X1 U14565 ( .A1(n12155), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11467) );
  OAI211_X1 U14566 ( .C1(n11470), .C2(n11469), .A(n11468), .B(n11467), .ZN(
        n11472) );
  NAND2_X1 U14567 ( .A1(n11472), .A2(n11471), .ZN(n11475) );
  OAI21_X1 U14568 ( .B1(n11473), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11495), .ZN(n19933) );
  NAND2_X1 U14569 ( .A1(n19933), .A2(n12150), .ZN(n11474) );
  NAND2_X1 U14570 ( .A1(n11475), .A2(n11474), .ZN(n11476) );
  AOI22_X1 U14571 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U14572 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U14573 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14574 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11479) );
  NAND4_X1 U14575 ( .A1(n11482), .A2(n11481), .A3(n11480), .A4(n11479), .ZN(
        n11491) );
  INV_X1 U14576 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11484) );
  INV_X1 U14577 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11483) );
  OAI22_X1 U14578 ( .A1(n11911), .A2(n11484), .B1(n9666), .B2(n11483), .ZN(
        n11485) );
  INV_X1 U14579 ( .A(n11485), .ZN(n11489) );
  AOI22_X1 U14580 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11488) );
  AOI22_X1 U14581 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11201), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11487) );
  INV_X1 U14582 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U14583 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11486) );
  NAND4_X1 U14584 ( .A1(n11489), .A2(n11488), .A3(n11487), .A4(n11486), .ZN(
        n11490) );
  NAND2_X1 U14585 ( .A1(n12034), .A2(n11976), .ZN(n11493) );
  NAND2_X1 U14586 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11492) );
  NAND2_X1 U14587 ( .A1(n11493), .A2(n11492), .ZN(n11501) );
  INV_X1 U14588 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13766) );
  AND2_X1 U14589 ( .A1(n11495), .A2(n11494), .ZN(n11496) );
  OR2_X1 U14590 ( .A1(n11496), .A2(n11518), .ZN(n19814) );
  AOI22_X1 U14591 ( .A1(n19814), .A2(n12150), .B1(n12154), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11497) );
  OAI21_X1 U14592 ( .B1(n11711), .B2(n13766), .A(n11497), .ZN(n11498) );
  NAND2_X1 U14593 ( .A1(n11500), .A2(n11499), .ZN(n13764) );
  INV_X1 U14594 ( .A(n13764), .ZN(n11523) );
  INV_X1 U14595 ( .A(n11501), .ZN(n11502) );
  NOR2_X2 U14596 ( .A1(n11503), .A2(n11502), .ZN(n11526) );
  AOI22_X1 U14597 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U14598 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11506) );
  AOI22_X1 U14599 ( .A1(n11336), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U14600 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11504) );
  NAND4_X1 U14601 ( .A1(n11507), .A2(n11506), .A3(n11505), .A4(n11504), .ZN(
        n11516) );
  INV_X1 U14602 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11509) );
  INV_X1 U14603 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11508) );
  OAI22_X1 U14604 ( .A1(n11911), .A2(n11509), .B1(n9665), .B2(n11508), .ZN(
        n11510) );
  INV_X1 U14605 ( .A(n11510), .ZN(n11514) );
  AOI22_X1 U14606 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U14607 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14608 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11511) );
  NAND4_X1 U14609 ( .A1(n11514), .A2(n11513), .A3(n11512), .A4(n11511), .ZN(
        n11515) );
  AOI22_X1 U14610 ( .A1(n12034), .A2(n11984), .B1(n12057), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11524) );
  NAND2_X1 U14611 ( .A1(n11517), .A2(n11524), .ZN(n11974) );
  INV_X1 U14612 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n19874) );
  NOR2_X1 U14613 ( .A1(n11518), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11519) );
  OR2_X1 U14614 ( .A1(n11530), .A2(n11519), .ZN(n19804) );
  AOI22_X1 U14615 ( .A1(n19804), .A2(n12150), .B1(n12154), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11520) );
  OAI21_X1 U14616 ( .B1(n11711), .B2(n19874), .A(n11520), .ZN(n11521) );
  NAND2_X1 U14617 ( .A1(n11523), .A2(n11522), .ZN(n13793) );
  INV_X1 U14618 ( .A(n11524), .ZN(n11525) );
  NAND2_X1 U14619 ( .A1(n12034), .A2(n11986), .ZN(n11528) );
  NAND2_X1 U14620 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11527) );
  NAND2_X1 U14621 ( .A1(n11528), .A2(n11527), .ZN(n11529) );
  INV_X1 U14622 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11533) );
  NOR2_X1 U14623 ( .A1(n11530), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11531) );
  OR2_X1 U14624 ( .A1(n11550), .A2(n11531), .ZN(n19803) );
  AOI22_X1 U14625 ( .A1(n19803), .A2(n12150), .B1(n12154), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11532) );
  OAI21_X1 U14626 ( .B1(n11711), .B2(n11533), .A(n11532), .ZN(n11534) );
  AOI21_X1 U14627 ( .B1(n11982), .B2(n11625), .A(n11534), .ZN(n13796) );
  AOI22_X1 U14629 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14630 ( .A1(n9651), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11537) );
  AOI22_X1 U14631 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14632 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11535) );
  NAND4_X1 U14633 ( .A1(n11538), .A2(n11537), .A3(n11536), .A4(n11535), .ZN(
        n11544) );
  AOI22_X1 U14634 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11542) );
  AOI22_X1 U14635 ( .A1(n12135), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11541) );
  AOI22_X1 U14636 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11201), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11540) );
  AOI22_X1 U14637 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11539) );
  NAND4_X1 U14638 ( .A1(n11542), .A2(n11541), .A3(n11540), .A4(n11539), .ZN(
        n11543) );
  OAI21_X1 U14639 ( .B1(n11544), .B2(n11543), .A(n11625), .ZN(n11549) );
  NAND2_X1 U14640 ( .A1(n12155), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11548) );
  INV_X1 U14641 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11545) );
  XNOR2_X1 U14642 ( .A(n11550), .B(n11545), .ZN(n13881) );
  OR2_X1 U14643 ( .A1(n13881), .A2(n11471), .ZN(n11547) );
  NAND2_X1 U14644 ( .A1(n12154), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11546) );
  NAND4_X1 U14645 ( .A1(n11549), .A2(n11548), .A3(n11547), .A4(n11546), .ZN(
        n13843) );
  NAND2_X1 U14646 ( .A1(n13794), .A2(n13843), .ZN(n13844) );
  XOR2_X1 U14647 ( .A(n19780), .B(n11565), .Z(n19779) );
  AOI22_X1 U14648 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U14649 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U14650 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11552) );
  AOI22_X1 U14651 ( .A1(n11336), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11551) );
  NAND4_X1 U14652 ( .A1(n11554), .A2(n11553), .A3(n11552), .A4(n11551), .ZN(
        n11560) );
  AOI22_X1 U14653 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U14654 ( .A1(n9651), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U14655 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11201), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U14656 ( .A1(n9669), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11555) );
  NAND4_X1 U14657 ( .A1(n11558), .A2(n11557), .A3(n11556), .A4(n11555), .ZN(
        n11559) );
  OR2_X1 U14658 ( .A1(n11560), .A2(n11559), .ZN(n11561) );
  AOI22_X1 U14659 ( .A1(n11625), .A2(n11561), .B1(n12154), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11563) );
  NAND2_X1 U14660 ( .A1(n12155), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11562) );
  OAI211_X1 U14661 ( .C1(n19779), .C2(n11471), .A(n11563), .B(n11562), .ZN(
        n13909) );
  INV_X1 U14662 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11566) );
  XNOR2_X1 U14663 ( .A(n11583), .B(n11566), .ZN(n15729) );
  OR2_X1 U14664 ( .A1(n15729), .A2(n11471), .ZN(n11582) );
  AOI22_X1 U14665 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14666 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U14667 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U14668 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11567) );
  NAND4_X1 U14669 ( .A1(n11570), .A2(n11569), .A3(n11568), .A4(n11567), .ZN(
        n11576) );
  AOI22_X1 U14670 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11574) );
  AOI22_X1 U14671 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U14672 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11572) );
  AOI22_X1 U14673 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11571) );
  NAND4_X1 U14674 ( .A1(n11574), .A2(n11573), .A3(n11572), .A4(n11571), .ZN(
        n11575) );
  NOR2_X1 U14675 ( .A1(n11576), .A2(n11575), .ZN(n11579) );
  NAND2_X1 U14676 ( .A1(n12155), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11578) );
  NAND2_X1 U14677 ( .A1(n12154), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11577) );
  OAI211_X1 U14678 ( .C1(n11660), .C2(n11579), .A(n11578), .B(n11577), .ZN(
        n11580) );
  INV_X1 U14679 ( .A(n11580), .ZN(n11581) );
  NAND2_X1 U14680 ( .A1(n11582), .A2(n11581), .ZN(n13894) );
  NAND2_X1 U14681 ( .A1(n12155), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n11586) );
  OAI21_X1 U14682 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11584), .A(
        n11628), .ZN(n15792) );
  AOI22_X1 U14683 ( .A1(n12150), .A2(n15792), .B1(n12154), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11585) );
  AOI22_X1 U14684 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11590) );
  AOI22_X1 U14685 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U14686 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U14687 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11587) );
  NAND4_X1 U14688 ( .A1(n11590), .A2(n11589), .A3(n11588), .A4(n11587), .ZN(
        n11599) );
  INV_X1 U14689 ( .A(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11592) );
  INV_X1 U14690 ( .A(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11591) );
  OAI22_X1 U14691 ( .A1(n11911), .A2(n11592), .B1(n9666), .B2(n11591), .ZN(
        n11593) );
  INV_X1 U14692 ( .A(n11593), .ZN(n11597) );
  AOI22_X1 U14693 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U14694 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9671), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U14695 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11594) );
  NAND4_X1 U14696 ( .A1(n11597), .A2(n11596), .A3(n11595), .A4(n11594), .ZN(
        n11598) );
  OR2_X1 U14697 ( .A1(n11599), .A2(n11598), .ZN(n11600) );
  NAND2_X1 U14698 ( .A1(n11625), .A2(n11600), .ZN(n14328) );
  INV_X1 U14699 ( .A(n14328), .ZN(n11601) );
  XOR2_X1 U14700 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11642), .Z(
        n15698) );
  AOI22_X1 U14701 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14702 ( .A1(n12135), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14703 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U14704 ( .A1(n11373), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11602) );
  NAND4_X1 U14705 ( .A1(n11605), .A2(n11604), .A3(n11603), .A4(n11602), .ZN(
        n11613) );
  INV_X1 U14706 ( .A(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11606) );
  INV_X1 U14707 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11754) );
  OAI22_X1 U14708 ( .A1(n11911), .A2(n11606), .B1(n11908), .B2(n11754), .ZN(
        n11607) );
  INV_X1 U14709 ( .A(n11607), .ZN(n11611) );
  AOI22_X1 U14710 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U14711 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9671), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U14712 ( .A1(n9670), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11608) );
  NAND4_X1 U14713 ( .A1(n11611), .A2(n11610), .A3(n11609), .A4(n11608), .ZN(
        n11612) );
  OR2_X1 U14714 ( .A1(n11613), .A2(n11612), .ZN(n11614) );
  AOI22_X1 U14715 ( .A1(n11625), .A2(n11614), .B1(n12154), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11616) );
  NAND2_X1 U14716 ( .A1(n12155), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11615) );
  OAI211_X1 U14717 ( .C1(n15698), .C2(n11471), .A(n11616), .B(n11615), .ZN(
        n14309) );
  INV_X1 U14718 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14399) );
  AOI22_X1 U14719 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11620) );
  AOI22_X1 U14720 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U14721 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14722 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11319), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11617) );
  NAND4_X1 U14723 ( .A1(n11620), .A2(n11619), .A3(n11618), .A4(n11617), .ZN(
        n11627) );
  AOI22_X1 U14724 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12135), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14725 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_8__4__SCAN_IN), .B2(n9672), .ZN(n11623) );
  AOI22_X1 U14726 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12112), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14727 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11621) );
  NAND4_X1 U14728 ( .A1(n11624), .A2(n11623), .A3(n11622), .A4(n11621), .ZN(
        n11626) );
  OAI21_X1 U14729 ( .B1(n11627), .B2(n11626), .A(n11625), .ZN(n11631) );
  XOR2_X1 U14730 ( .A(n15709), .B(n11628), .Z(n15780) );
  INV_X1 U14731 ( .A(n15780), .ZN(n11629) );
  AOI22_X1 U14732 ( .A1(n12150), .A2(n11629), .B1(n12154), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11630) );
  OAI211_X1 U14733 ( .C1(n11711), .C2(n14399), .A(n11631), .B(n11630), .ZN(
        n14317) );
  AOI22_X1 U14734 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U14735 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U14736 ( .A1(n11373), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11633) );
  AOI22_X1 U14737 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11632) );
  NAND4_X1 U14738 ( .A1(n11635), .A2(n11634), .A3(n11633), .A4(n11632), .ZN(
        n11641) );
  AOI22_X1 U14739 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11639) );
  AOI22_X1 U14740 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11638) );
  AOI22_X1 U14741 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9671), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11637) );
  AOI22_X1 U14742 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11636) );
  NAND4_X1 U14743 ( .A1(n11639), .A2(n11638), .A3(n11637), .A4(n11636), .ZN(
        n11640) );
  NOR2_X1 U14744 ( .A1(n11641), .A2(n11640), .ZN(n11645) );
  XNOR2_X1 U14745 ( .A(n11646), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14511) );
  NAND2_X1 U14746 ( .A1(n14511), .A2(n12150), .ZN(n11644) );
  AOI22_X1 U14747 ( .A1(n12155), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n12154), 
        .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11643) );
  OAI211_X1 U14748 ( .C1(n11645), .C2(n11660), .A(n11644), .B(n11643), .ZN(
        n14216) );
  INV_X1 U14749 ( .A(n14215), .ZN(n11664) );
  XOR2_X1 U14750 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n11665), .Z(
        n15775) );
  INV_X1 U14751 ( .A(n15775), .ZN(n11662) );
  AOI22_X1 U14752 ( .A1(n12135), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11650) );
  AOI22_X1 U14753 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U14754 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U14755 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11647) );
  NAND4_X1 U14756 ( .A1(n11650), .A2(n11649), .A3(n11648), .A4(n11647), .ZN(
        n11656) );
  AOI22_X1 U14757 ( .A1(n9651), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11654) );
  AOI22_X1 U14758 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14759 ( .A1(n11319), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11201), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14760 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11651) );
  NAND4_X1 U14761 ( .A1(n11654), .A2(n11653), .A3(n11652), .A4(n11651), .ZN(
        n11655) );
  NOR2_X1 U14762 ( .A1(n11656), .A2(n11655), .ZN(n11659) );
  NAND2_X1 U14763 ( .A1(n12155), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11658) );
  NAND2_X1 U14764 ( .A1(n12154), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11657) );
  OAI211_X1 U14765 ( .C1(n11660), .C2(n11659), .A(n11658), .B(n11657), .ZN(
        n11661) );
  AOI21_X1 U14766 ( .B1(n11662), .B2(n12150), .A(n11661), .ZN(n14298) );
  INV_X1 U14767 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15681) );
  XNOR2_X1 U14768 ( .A(n11685), .B(n15681), .ZN(n15678) );
  NAND2_X1 U14769 ( .A1(n15678), .A2(n12150), .ZN(n11684) );
  AOI22_X1 U14770 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11669) );
  AOI22_X1 U14771 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11458), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U14772 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11667) );
  AOI22_X1 U14773 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11666) );
  NAND4_X1 U14774 ( .A1(n11669), .A2(n11668), .A3(n11667), .A4(n11666), .ZN(
        n11680) );
  NAND2_X1 U14775 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11671) );
  NAND2_X1 U14776 ( .A1(n11757), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11670) );
  AND3_X1 U14777 ( .A1(n11671), .A2(n11471), .A3(n11670), .ZN(n11678) );
  INV_X1 U14778 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11672) );
  OAI22_X1 U14779 ( .A1(n11908), .A2(n11673), .B1(n9666), .B2(n11672), .ZN(
        n11674) );
  INV_X1 U14780 ( .A(n11674), .ZN(n11677) );
  AOI22_X1 U14781 ( .A1(n12129), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14782 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11201), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11675) );
  NAND4_X1 U14783 ( .A1(n11678), .A2(n11677), .A3(n11676), .A4(n11675), .ZN(
        n11679) );
  INV_X1 U14784 ( .A(n11280), .ZN(n13983) );
  NAND2_X1 U14785 ( .A1(n12123), .A2(n11471), .ZN(n11786) );
  OAI21_X1 U14786 ( .B1(n11680), .B2(n11679), .A(n11786), .ZN(n11682) );
  AOI22_X1 U14787 ( .A1(n12155), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20581), .ZN(n11681) );
  NAND2_X1 U14788 ( .A1(n11682), .A2(n11681), .ZN(n11683) );
  NAND2_X1 U14789 ( .A1(n11684), .A2(n11683), .ZN(n14290) );
  XOR2_X1 U14790 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11698), .Z(
        n15762) );
  AOI22_X1 U14791 ( .A1(n12155), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n12154), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U14792 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U14793 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U14794 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14795 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11686) );
  NAND4_X1 U14796 ( .A1(n11689), .A2(n11688), .A3(n11687), .A4(n11686), .ZN(
        n11695) );
  AOI22_X1 U14797 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14798 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11458), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14799 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9671), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14800 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11690) );
  NAND4_X1 U14801 ( .A1(n11693), .A2(n11692), .A3(n11691), .A4(n11690), .ZN(
        n11694) );
  INV_X1 U14802 ( .A(n12123), .ZN(n12146) );
  OAI21_X1 U14803 ( .B1(n11695), .B2(n11694), .A(n12146), .ZN(n11696) );
  OAI211_X1 U14804 ( .C1(n15762), .C2(n11471), .A(n11697), .B(n11696), .ZN(
        n14286) );
  XNOR2_X1 U14805 ( .A(n11730), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15663) );
  AOI22_X1 U14806 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11704) );
  AOI22_X1 U14807 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11703) );
  AOI22_X1 U14808 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11702) );
  NAND2_X1 U14809 ( .A1(n11373), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11700) );
  NAND2_X1 U14810 ( .A1(n11311), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11699) );
  AND3_X1 U14811 ( .A1(n11700), .A2(n11471), .A3(n11699), .ZN(n11701) );
  NAND4_X1 U14812 ( .A1(n11704), .A2(n11703), .A3(n11702), .A4(n11701), .ZN(
        n11710) );
  AOI22_X1 U14813 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U14814 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11707) );
  AOI22_X1 U14815 ( .A1(n9651), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11706) );
  AOI22_X1 U14816 ( .A1(n12111), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11705) );
  NAND4_X1 U14817 ( .A1(n11708), .A2(n11707), .A3(n11706), .A4(n11705), .ZN(
        n11709) );
  OR2_X1 U14818 ( .A1(n11710), .A2(n11709), .ZN(n11713) );
  INV_X1 U14819 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14380) );
  INV_X1 U14820 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11729) );
  OAI22_X1 U14821 ( .A1(n11711), .A2(n14380), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n11729), .ZN(n11712) );
  AOI21_X1 U14822 ( .B1(n11786), .B2(n11713), .A(n11712), .ZN(n11714) );
  AOI21_X1 U14823 ( .B1(n15663), .B2(n12150), .A(n11714), .ZN(n14276) );
  AOI22_X1 U14824 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11718) );
  AOI22_X1 U14825 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11717) );
  AOI22_X1 U14826 ( .A1(n9651), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(n9671), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U14827 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11715) );
  NAND4_X1 U14828 ( .A1(n11718), .A2(n11717), .A3(n11716), .A4(n11715), .ZN(
        n11724) );
  AOI22_X1 U14829 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11722) );
  AOI22_X1 U14830 ( .A1(n11336), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11721) );
  AOI22_X1 U14831 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11458), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U14832 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11719) );
  NAND4_X1 U14833 ( .A1(n11722), .A2(n11721), .A3(n11720), .A4(n11719), .ZN(
        n11723) );
  NOR2_X1 U14834 ( .A1(n11724), .A2(n11723), .ZN(n11728) );
  OAI21_X1 U14835 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20468), .A(
        n20581), .ZN(n11725) );
  INV_X1 U14836 ( .A(n11725), .ZN(n11726) );
  AOI21_X1 U14837 ( .B1(n12155), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11726), .ZN(
        n11727) );
  OAI21_X1 U14838 ( .B1(n12123), .B2(n11728), .A(n11727), .ZN(n11733) );
  OAI21_X1 U14839 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n11731), .A(
        n11768), .ZN(n15756) );
  OR2_X1 U14840 ( .A1(n11471), .A2(n15756), .ZN(n11732) );
  NAND2_X1 U14841 ( .A1(n11733), .A2(n11732), .ZN(n14273) );
  AOI22_X1 U14842 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U14843 ( .A1(n12135), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U14844 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11200), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U14845 ( .A1(n11373), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11735) );
  NAND4_X1 U14846 ( .A1(n11738), .A2(n11737), .A3(n11736), .A4(n11735), .ZN(
        n11744) );
  AOI22_X1 U14847 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11742) );
  AOI22_X1 U14848 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11458), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U14849 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_9__4__SCAN_IN), .B2(n9671), .ZN(n11740) );
  AOI22_X1 U14850 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11311), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11739) );
  NAND4_X1 U14851 ( .A1(n11742), .A2(n11741), .A3(n11740), .A4(n11739), .ZN(
        n11743) );
  NOR2_X1 U14852 ( .A1(n11744), .A2(n11743), .ZN(n11747) );
  INV_X1 U14853 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15649) );
  AOI21_X1 U14854 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15649), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11745) );
  AOI21_X1 U14855 ( .B1(n12155), .B2(P1_EAX_REG_20__SCAN_IN), .A(n11745), .ZN(
        n11746) );
  OAI21_X1 U14856 ( .B1(n12123), .B2(n11747), .A(n11746), .ZN(n11749) );
  XNOR2_X1 U14857 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n11768), .ZN(
        n15640) );
  NAND2_X1 U14858 ( .A1(n12150), .A2(n15640), .ZN(n11748) );
  NAND2_X1 U14859 ( .A1(n11749), .A2(n11748), .ZN(n14264) );
  AOI22_X1 U14860 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11753) );
  AOI22_X1 U14861 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U14862 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12111), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U14863 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11750) );
  NAND4_X1 U14864 ( .A1(n11753), .A2(n11752), .A3(n11751), .A4(n11750), .ZN(
        n11763) );
  INV_X1 U14865 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11755) );
  OAI22_X1 U14866 ( .A1(n11911), .A2(n11755), .B1(n9665), .B2(n11754), .ZN(
        n11756) );
  INV_X1 U14867 ( .A(n11756), .ZN(n11761) );
  AOI22_X1 U14868 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U14869 ( .A1(n11458), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9671), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11759) );
  AOI22_X1 U14870 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11758) );
  NAND4_X1 U14871 ( .A1(n11761), .A2(n11760), .A3(n11759), .A4(n11758), .ZN(
        n11762) );
  NOR2_X1 U14872 ( .A1(n11763), .A2(n11762), .ZN(n11767) );
  NAND2_X1 U14873 ( .A1(n20581), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11764) );
  NAND2_X1 U14874 ( .A1(n11471), .A2(n11764), .ZN(n11765) );
  AOI21_X1 U14875 ( .B1(n12155), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11765), .ZN(
        n11766) );
  OAI21_X1 U14876 ( .B1(n12123), .B2(n11767), .A(n11766), .ZN(n11772) );
  OAI21_X1 U14877 ( .B1(n11770), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n11814), .ZN(n15627) );
  OR2_X1 U14878 ( .A1(n15627), .A2(n11471), .ZN(n11771) );
  AOI22_X1 U14879 ( .A1(n9651), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11320), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11778) );
  NAND2_X1 U14880 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11774) );
  NAND2_X1 U14881 ( .A1(n11311), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11773) );
  AND3_X1 U14882 ( .A1(n11774), .A2(n11471), .A3(n11773), .ZN(n11777) );
  AOI22_X1 U14883 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U14884 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11775) );
  NAND4_X1 U14885 ( .A1(n11778), .A2(n11777), .A3(n11776), .A4(n11775), .ZN(
        n11784) );
  AOI22_X1 U14886 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U14887 ( .A1(n11373), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U14888 ( .A1(n12135), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11458), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U14889 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11779) );
  NAND4_X1 U14890 ( .A1(n11782), .A2(n11781), .A3(n11780), .A4(n11779), .ZN(
        n11783) );
  OR2_X1 U14891 ( .A1(n11784), .A2(n11783), .ZN(n11785) );
  NAND2_X1 U14892 ( .A1(n11786), .A2(n11785), .ZN(n11789) );
  AOI22_X1 U14893 ( .A1(n12155), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20581), .ZN(n11788) );
  XNOR2_X1 U14894 ( .A(n11814), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15620) );
  AOI21_X1 U14895 ( .B1(n11789), .B2(n11788), .A(n11787), .ZN(n14250) );
  AOI22_X1 U14896 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U14897 ( .A1(n9673), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U14898 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(n9671), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U14899 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11790) );
  NAND4_X1 U14900 ( .A1(n11793), .A2(n11792), .A3(n11791), .A4(n11790), .ZN(
        n11799) );
  AOI22_X1 U14901 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U14902 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11796) );
  AOI22_X1 U14903 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11795) );
  AOI22_X1 U14904 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11794) );
  NAND4_X1 U14905 ( .A1(n11797), .A2(n11796), .A3(n11795), .A4(n11794), .ZN(
        n11798) );
  NOR2_X1 U14906 ( .A1(n11799), .A2(n11798), .ZN(n11819) );
  AOI22_X1 U14907 ( .A1(n12135), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11803) );
  AOI22_X1 U14908 ( .A1(n9651), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11201), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U14909 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U14910 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11800) );
  NAND4_X1 U14911 ( .A1(n11803), .A2(n11802), .A3(n11801), .A4(n11800), .ZN(
        n11809) );
  AOI22_X1 U14912 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11807) );
  AOI22_X1 U14913 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11806) );
  AOI22_X1 U14914 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11805) );
  AOI22_X1 U14915 ( .A1(n12111), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11804) );
  NAND4_X1 U14916 ( .A1(n11807), .A2(n11806), .A3(n11805), .A4(n11804), .ZN(
        n11808) );
  NOR2_X1 U14917 ( .A1(n11809), .A2(n11808), .ZN(n11820) );
  XNOR2_X1 U14918 ( .A(n11819), .B(n11820), .ZN(n11813) );
  NAND2_X1 U14919 ( .A1(n20581), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11810) );
  NAND2_X1 U14920 ( .A1(n11471), .A2(n11810), .ZN(n11811) );
  AOI21_X1 U14921 ( .B1(n12155), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11811), .ZN(
        n11812) );
  OAI21_X1 U14922 ( .B1(n11813), .B2(n12123), .A(n11812), .ZN(n11818) );
  INV_X1 U14923 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15617) );
  OR2_X1 U14924 ( .A1(n11815), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11816) );
  AND2_X1 U14925 ( .A1(n11841), .A2(n11816), .ZN(n15607) );
  NAND2_X1 U14926 ( .A1(n15607), .A2(n12150), .ZN(n11817) );
  NAND2_X1 U14927 ( .A1(n11818), .A2(n11817), .ZN(n14462) );
  NOR2_X1 U14928 ( .A1(n11820), .A2(n11819), .ZN(n11858) );
  AOI22_X1 U14929 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U14930 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11823) );
  AOI22_X1 U14931 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11822) );
  AOI22_X1 U14932 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11821) );
  NAND4_X1 U14933 ( .A1(n11824), .A2(n11823), .A3(n11822), .A4(n11821), .ZN(
        n11833) );
  INV_X1 U14934 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11826) );
  INV_X1 U14935 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11825) );
  OAI22_X1 U14936 ( .A1(n11911), .A2(n11826), .B1(n9665), .B2(n11825), .ZN(
        n11827) );
  INV_X1 U14937 ( .A(n11827), .ZN(n11831) );
  AOI22_X1 U14938 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11830) );
  AOI22_X1 U14939 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11201), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U14940 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11828) );
  NAND4_X1 U14941 ( .A1(n11831), .A2(n11830), .A3(n11829), .A4(n11828), .ZN(
        n11832) );
  OR2_X1 U14942 ( .A1(n11833), .A2(n11832), .ZN(n11857) );
  XNOR2_X1 U14943 ( .A(n11858), .B(n11857), .ZN(n11837) );
  NAND2_X1 U14944 ( .A1(n20581), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11834) );
  NAND2_X1 U14945 ( .A1(n11471), .A2(n11834), .ZN(n11835) );
  AOI21_X1 U14946 ( .B1(n12155), .B2(P1_EAX_REG_24__SCAN_IN), .A(n11835), .ZN(
        n11836) );
  OAI21_X1 U14947 ( .B1(n11837), .B2(n12123), .A(n11836), .ZN(n11839) );
  XNOR2_X1 U14948 ( .A(n11841), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15601) );
  NAND2_X1 U14949 ( .A1(n15601), .A2(n12150), .ZN(n11838) );
  NAND2_X1 U14950 ( .A1(n11839), .A2(n11838), .ZN(n14242) );
  INV_X1 U14951 ( .A(n11841), .ZN(n11842) );
  INV_X1 U14952 ( .A(n11843), .ZN(n11845) );
  INV_X1 U14953 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11844) );
  NAND2_X1 U14954 ( .A1(n11845), .A2(n11844), .ZN(n11846) );
  NAND2_X1 U14955 ( .A1(n11882), .A2(n11846), .ZN(n14452) );
  AOI22_X1 U14956 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12112), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U14957 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(n9672), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U14958 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U14959 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11847) );
  NAND4_X1 U14960 ( .A1(n11850), .A2(n11849), .A3(n11848), .A4(n11847), .ZN(
        n11856) );
  AOI22_X1 U14961 ( .A1(n12135), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11854) );
  AOI22_X1 U14962 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11853) );
  AOI22_X1 U14963 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11852) );
  AOI22_X1 U14964 ( .A1(n12111), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11851) );
  NAND4_X1 U14965 ( .A1(n11854), .A2(n11853), .A3(n11852), .A4(n11851), .ZN(
        n11855) );
  NOR2_X1 U14966 ( .A1(n11856), .A2(n11855), .ZN(n11864) );
  NAND2_X1 U14967 ( .A1(n11858), .A2(n11857), .ZN(n11863) );
  XNOR2_X1 U14968 ( .A(n11864), .B(n11863), .ZN(n11861) );
  AOI21_X1 U14969 ( .B1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20581), .A(
        n12150), .ZN(n11860) );
  NAND2_X1 U14970 ( .A1(n12155), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n11859) );
  OAI211_X1 U14971 ( .C1(n11861), .C2(n12123), .A(n11860), .B(n11859), .ZN(
        n11862) );
  NOR2_X2 U14972 ( .A1(n14200), .A2(n14201), .ZN(n14187) );
  XNOR2_X1 U14973 ( .A(n11882), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14444) );
  INV_X1 U14974 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14440) );
  AOI21_X1 U14975 ( .B1(n14440), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11880) );
  NOR2_X1 U14976 ( .A1(n11864), .A2(n11863), .ZN(n11900) );
  AOI22_X1 U14977 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11868) );
  AOI22_X1 U14978 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U14979 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11866) );
  AOI22_X1 U14980 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11865) );
  NAND4_X1 U14981 ( .A1(n11868), .A2(n11867), .A3(n11866), .A4(n11865), .ZN(
        n11877) );
  INV_X1 U14982 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11870) );
  INV_X1 U14983 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11869) );
  OAI22_X1 U14984 ( .A1(n11911), .A2(n11870), .B1(n9666), .B2(n11869), .ZN(
        n11871) );
  INV_X1 U14985 ( .A(n11871), .ZN(n11875) );
  AOI22_X1 U14986 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U14987 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11873) );
  AOI22_X1 U14988 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11757), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11872) );
  NAND4_X1 U14989 ( .A1(n11875), .A2(n11874), .A3(n11873), .A4(n11872), .ZN(
        n11876) );
  OR2_X1 U14990 ( .A1(n11877), .A2(n11876), .ZN(n11899) );
  XNOR2_X1 U14991 ( .A(n11900), .B(n11899), .ZN(n11878) );
  NOR2_X1 U14992 ( .A1(n11878), .A2(n12123), .ZN(n11879) );
  AOI211_X1 U14993 ( .C1(n12155), .C2(P1_EAX_REG_26__SCAN_IN), .A(n11880), .B(
        n11879), .ZN(n11881) );
  NAND2_X1 U14994 ( .A1(n14187), .A2(n14189), .ZN(n14175) );
  INV_X1 U14995 ( .A(n11882), .ZN(n11883) );
  INV_X1 U14996 ( .A(n11884), .ZN(n11886) );
  INV_X1 U14997 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11885) );
  NAND2_X1 U14998 ( .A1(n11886), .A2(n11885), .ZN(n11887) );
  NAND2_X1 U14999 ( .A1(n12102), .A2(n11887), .ZN(n14433) );
  AOI22_X1 U15000 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U15001 ( .A1(n9651), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        P1_INSTQUEUE_REG_10__4__SCAN_IN), .B2(n11201), .ZN(n11890) );
  AOI22_X1 U15002 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11889) );
  AOI22_X1 U15003 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11311), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11888) );
  NAND4_X1 U15004 ( .A1(n11891), .A2(n11890), .A3(n11889), .A4(n11888), .ZN(
        n11898) );
  AOI22_X1 U15005 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n9667), .B1(
        n12106), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11896) );
  AOI22_X1 U15006 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U15007 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11458), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U15008 ( .A1(n12111), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11893) );
  NAND4_X1 U15009 ( .A1(n11896), .A2(n11895), .A3(n11894), .A4(n11893), .ZN(
        n11897) );
  NOR2_X1 U15010 ( .A1(n11898), .A2(n11897), .ZN(n11906) );
  NAND2_X1 U15011 ( .A1(n11900), .A2(n11899), .ZN(n11905) );
  XNOR2_X1 U15012 ( .A(n11906), .B(n11905), .ZN(n11903) );
  AOI21_X1 U15013 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20581), .A(
        n12150), .ZN(n11902) );
  NAND2_X1 U15014 ( .A1(n12155), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n11901) );
  OAI211_X1 U15015 ( .C1(n11903), .C2(n12123), .A(n11902), .B(n11901), .ZN(
        n11904) );
  XNOR2_X1 U15016 ( .A(n12102), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14172) );
  INV_X1 U15017 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14165) );
  OAI21_X1 U15018 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14165), .A(n11471), 
        .ZN(n11924) );
  NOR2_X1 U15019 ( .A1(n11906), .A2(n11905), .ZN(n12120) );
  INV_X1 U15020 ( .A(n12130), .ZN(n11908) );
  INV_X1 U15021 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11907) );
  NOR2_X1 U15022 ( .A1(n11908), .A2(n11907), .ZN(n11913) );
  INV_X1 U15023 ( .A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11910) );
  OAI22_X1 U15024 ( .A1(n11911), .A2(n11910), .B1(n9665), .B2(n11909), .ZN(
        n11912) );
  AOI211_X1 U15025 ( .C1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .C2(n11458), .A(
        n11913), .B(n11912), .ZN(n11921) );
  AOI22_X1 U15026 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11917) );
  AOI22_X1 U15027 ( .A1(n11200), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9673), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11916) );
  AOI22_X1 U15028 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U15029 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11914) );
  AND4_X1 U15030 ( .A1(n11917), .A2(n11916), .A3(n11915), .A4(n11914), .ZN(
        n11920) );
  AOI22_X1 U15031 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11919) );
  AOI22_X1 U15032 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11311), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11918) );
  NAND4_X1 U15033 ( .A1(n11921), .A2(n11920), .A3(n11919), .A4(n11918), .ZN(
        n12119) );
  XNOR2_X1 U15034 ( .A(n12120), .B(n12119), .ZN(n11922) );
  NOR2_X1 U15035 ( .A1(n11922), .A2(n12123), .ZN(n11923) );
  AOI211_X1 U15036 ( .C1(n12155), .C2(P1_EAX_REG_28__SCAN_IN), .A(n11924), .B(
        n11923), .ZN(n11925) );
  AOI21_X1 U15037 ( .B1(n12150), .B2(n14172), .A(n11925), .ZN(n11926) );
  NAND2_X1 U15038 ( .A1(n11928), .A2(n12126), .ZN(n14235) );
  NAND3_X1 U15039 ( .A1(n20578), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15912) );
  INV_X1 U15040 ( .A(n15912), .ZN(n11929) );
  NOR2_X2 U15041 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20657) );
  NOR2_X1 U15042 ( .A1(n14235), .A2(n20003), .ZN(n12076) );
  NAND2_X1 U15043 ( .A1(n11941), .A2(n11935), .ZN(n11951) );
  XNOR2_X1 U15044 ( .A(n11951), .B(n11950), .ZN(n11932) );
  NAND2_X1 U15045 ( .A1(n11270), .A2(n20025), .ZN(n11940) );
  INV_X1 U15046 ( .A(n11940), .ZN(n11931) );
  AOI21_X1 U15047 ( .B1(n11932), .B2(n15572), .A(n11931), .ZN(n11933) );
  XNOR2_X1 U15048 ( .A(n11941), .B(n11935), .ZN(n11938) );
  INV_X1 U15049 ( .A(n11936), .ZN(n11937) );
  OAI211_X1 U15050 ( .C1(n11938), .C2(n11295), .A(n11937), .B(n20032), .ZN(
        n11939) );
  OR2_X1 U15051 ( .A1(n20078), .A2(n12022), .ZN(n11944) );
  OAI21_X1 U15052 ( .B1(n11295), .B2(n11941), .A(n11940), .ZN(n11942) );
  INV_X1 U15053 ( .A(n11942), .ZN(n11943) );
  NAND2_X1 U15054 ( .A1(n11944), .A2(n11943), .ZN(n19936) );
  NAND2_X1 U15055 ( .A1(n19936), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n19935) );
  XNOR2_X1 U15056 ( .A(n11946), .B(n19935), .ZN(n13296) );
  NAND2_X1 U15057 ( .A1(n13296), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13297) );
  INV_X1 U15058 ( .A(n19935), .ZN(n11945) );
  NAND2_X1 U15059 ( .A1(n11946), .A2(n11945), .ZN(n11947) );
  NAND2_X1 U15060 ( .A1(n13297), .A2(n11947), .ZN(n11948) );
  INV_X1 U15061 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19984) );
  XNOR2_X1 U15062 ( .A(n11948), .B(n19984), .ZN(n13355) );
  NAND2_X1 U15063 ( .A1(n11948), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11949) );
  INV_X1 U15064 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19967) );
  OR2_X1 U15065 ( .A1(n20004), .A2(n12022), .ZN(n11955) );
  NAND2_X1 U15066 ( .A1(n11951), .A2(n11950), .ZN(n11968) );
  INV_X1 U15067 ( .A(n11966), .ZN(n11952) );
  XNOR2_X1 U15068 ( .A(n11968), .B(n11952), .ZN(n11953) );
  NAND2_X1 U15069 ( .A1(n11953), .A2(n15572), .ZN(n11954) );
  NAND2_X1 U15070 ( .A1(n11955), .A2(n11954), .ZN(n13525) );
  INV_X1 U15071 ( .A(n12022), .ZN(n13187) );
  NAND2_X1 U15072 ( .A1(n11968), .A2(n11966), .ZN(n11958) );
  XNOR2_X1 U15073 ( .A(n11958), .B(n11965), .ZN(n11959) );
  NAND2_X1 U15074 ( .A1(n11959), .A2(n15572), .ZN(n11960) );
  NAND2_X1 U15075 ( .A1(n11961), .A2(n11960), .ZN(n11962) );
  INV_X1 U15076 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19957) );
  NAND2_X1 U15077 ( .A1(n11964), .A2(n13187), .ZN(n11971) );
  AND2_X1 U15078 ( .A1(n11966), .A2(n11965), .ZN(n11967) );
  NAND2_X1 U15079 ( .A1(n11968), .A2(n11967), .ZN(n11975) );
  XNOR2_X1 U15080 ( .A(n11975), .B(n11976), .ZN(n11969) );
  NAND2_X1 U15081 ( .A1(n11969), .A2(n15572), .ZN(n11970) );
  NAND2_X1 U15082 ( .A1(n11971), .A2(n11970), .ZN(n11972) );
  INV_X1 U15083 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15868) );
  XNOR2_X1 U15084 ( .A(n11972), .B(n15868), .ZN(n15806) );
  NAND2_X1 U15085 ( .A1(n11972), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11973) );
  NAND3_X1 U15086 ( .A1(n11993), .A2(n13187), .A3(n11974), .ZN(n11980) );
  INV_X1 U15087 ( .A(n11975), .ZN(n11977) );
  NAND2_X1 U15088 ( .A1(n11977), .A2(n11976), .ZN(n11983) );
  XNOR2_X1 U15089 ( .A(n11983), .B(n11984), .ZN(n11978) );
  NAND2_X1 U15090 ( .A1(n11978), .A2(n15572), .ZN(n11979) );
  NAND2_X1 U15091 ( .A1(n11980), .A2(n11979), .ZN(n15800) );
  OR2_X1 U15092 ( .A1(n15800), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11981) );
  NAND2_X1 U15093 ( .A1(n11982), .A2(n13187), .ZN(n11989) );
  INV_X1 U15094 ( .A(n11983), .ZN(n11985) );
  NAND2_X1 U15095 ( .A1(n11985), .A2(n11984), .ZN(n11995) );
  XNOR2_X1 U15096 ( .A(n11995), .B(n11986), .ZN(n11987) );
  NAND2_X1 U15097 ( .A1(n11987), .A2(n15572), .ZN(n11988) );
  NAND2_X1 U15098 ( .A1(n11989), .A2(n11988), .ZN(n11990) );
  OR2_X1 U15099 ( .A1(n11990), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15794) );
  NAND2_X1 U15100 ( .A1(n11990), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15793) );
  NOR2_X1 U15101 ( .A1(n11991), .A2(n12022), .ZN(n11992) );
  OR3_X1 U15102 ( .A1(n11995), .A2(n11994), .A3(n11295), .ZN(n11996) );
  NAND2_X1 U15103 ( .A1(n15785), .A2(n11996), .ZN(n13879) );
  OR2_X1 U15104 ( .A1(n13879), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11997) );
  NAND2_X1 U15105 ( .A1(n13879), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11998) );
  INV_X4 U15106 ( .A(n14015), .ZN(n14479) );
  INV_X1 U15107 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11999) );
  NAND2_X1 U15108 ( .A1(n15785), .A2(n11999), .ZN(n12000) );
  INV_X1 U15109 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14727) );
  OR2_X1 U15110 ( .A1(n15785), .A2(n14727), .ZN(n14506) );
  NAND2_X1 U15111 ( .A1(n15785), .A2(n14727), .ZN(n14517) );
  NAND2_X1 U15112 ( .A1(n14506), .A2(n14517), .ZN(n14520) );
  AND2_X1 U15113 ( .A1(n15785), .A2(n14737), .ZN(n12001) );
  NAND2_X1 U15114 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12002) );
  AND2_X1 U15115 ( .A1(n15785), .A2(n12002), .ZN(n14519) );
  INV_X1 U15116 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14068) );
  NAND2_X1 U15117 ( .A1(n14479), .A2(n14068), .ZN(n12003) );
  NOR2_X1 U15118 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12004) );
  XNOR2_X1 U15119 ( .A(n14479), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14501) );
  NAND2_X1 U15120 ( .A1(n14479), .A2(n15837), .ZN(n15771) );
  AND2_X1 U15121 ( .A1(n14501), .A2(n15771), .ZN(n12005) );
  NAND2_X1 U15122 ( .A1(n12006), .A2(n12005), .ZN(n15757) );
  INV_X1 U15123 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14694) );
  INV_X1 U15124 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15822) );
  NOR2_X1 U15125 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12009) );
  XNOR2_X1 U15126 ( .A(n14479), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14489) );
  NAND2_X1 U15127 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14546) );
  INV_X1 U15128 ( .A(n14546), .ZN(n12011) );
  INV_X1 U15129 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12012) );
  INV_X1 U15130 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14662) );
  INV_X1 U15131 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15820) );
  INV_X1 U15132 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12014) );
  AND2_X1 U15133 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14604) );
  NAND2_X1 U15134 ( .A1(n14604), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14607) );
  NAND2_X1 U15135 ( .A1(n14479), .A2(n14607), .ZN(n14437) );
  NAND3_X1 U15136 ( .A1(n14013), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n14437), .ZN(n12015) );
  OAI21_X1 U15137 ( .B1(n14406), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12015), .ZN(n12017) );
  INV_X1 U15138 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14430) );
  MUX2_X1 U15139 ( .A(n14430), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n15785), .Z(n12016) );
  NAND2_X1 U15140 ( .A1(n12017), .A2(n12016), .ZN(n12018) );
  INV_X1 U15141 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14589) );
  XNOR2_X1 U15142 ( .A(n12018), .B(n14589), .ZN(n14594) );
  XNOR2_X1 U15143 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12033) );
  NAND2_X1 U15144 ( .A1(n20665), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12036) );
  NAND2_X1 U15145 ( .A1(n12033), .A2(n12032), .ZN(n12020) );
  NAND2_X1 U15146 ( .A1(n20327), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12019) );
  XNOR2_X1 U15147 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12028) );
  XNOR2_X1 U15148 ( .A(n10048), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12026) );
  INV_X1 U15149 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20000) );
  NOR2_X1 U15150 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20000), .ZN(
        n12021) );
  NAND2_X1 U15151 ( .A1(n12167), .A2(n12056), .ZN(n12065) );
  NAND2_X1 U15152 ( .A1(n12167), .A2(n12034), .ZN(n12063) );
  NAND3_X1 U15153 ( .A1(n11469), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n12023), .ZN(n12165) );
  INV_X1 U15154 ( .A(n12056), .ZN(n12060) );
  AOI21_X1 U15155 ( .B1(n12026), .B2(n12025), .A(n12024), .ZN(n12027) );
  INV_X1 U15156 ( .A(n12027), .ZN(n12164) );
  XNOR2_X1 U15157 ( .A(n12029), .B(n12028), .ZN(n12162) );
  NAND2_X1 U15158 ( .A1(n12030), .A2(n20005), .ZN(n12031) );
  NAND2_X1 U15159 ( .A1(n12031), .A2(n9592), .ZN(n12051) );
  XNOR2_X1 U15160 ( .A(n12033), .B(n12032), .ZN(n12163) );
  INV_X1 U15161 ( .A(n12045), .ZN(n12035) );
  NOR2_X1 U15162 ( .A1(n12163), .A2(n12035), .ZN(n12041) );
  OAI21_X1 U15163 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20665), .A(
        n12036), .ZN(n12037) );
  NOR2_X1 U15164 ( .A1(n12052), .A2(n12037), .ZN(n12040) );
  INV_X1 U15165 ( .A(n12037), .ZN(n12038) );
  OAI211_X1 U15166 ( .C1(n11270), .C2(n11275), .A(n12038), .B(n12051), .ZN(
        n12039) );
  OAI21_X1 U15167 ( .B1(n12056), .B2(n12040), .A(n12039), .ZN(n12042) );
  AND2_X1 U15168 ( .A1(n12041), .A2(n12042), .ZN(n12050) );
  INV_X1 U15169 ( .A(n12163), .ZN(n12044) );
  NOR2_X1 U15170 ( .A1(n12045), .A2(n12042), .ZN(n12043) );
  AOI211_X1 U15171 ( .C1(n12045), .C2(n11930), .A(n12044), .B(n12043), .ZN(
        n12049) );
  INV_X1 U15172 ( .A(n12051), .ZN(n12047) );
  NOR2_X1 U15173 ( .A1(n12052), .A2(n12162), .ZN(n12046) );
  AOI211_X1 U15174 ( .C1(n12057), .C2(n12162), .A(n12047), .B(n12046), .ZN(
        n12048) );
  OAI33_X1 U15175 ( .A1(n12162), .A2(n12052), .A3(n12051), .B1(n12050), .B2(
        n12049), .B3(n12048), .ZN(n12055) );
  NAND2_X1 U15176 ( .A1(n12053), .A2(n12164), .ZN(n12054) );
  AOI22_X1 U15177 ( .A1(n12056), .A2(n12164), .B1(n12055), .B2(n12054), .ZN(
        n12059) );
  NOR2_X1 U15178 ( .A1(n12057), .A2(n12165), .ZN(n12058) );
  OAI22_X1 U15179 ( .A1(n12165), .A2(n12060), .B1(n12059), .B2(n12058), .ZN(
        n12061) );
  AOI21_X1 U15180 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20578), .A(
        n12061), .ZN(n12062) );
  NAND2_X1 U15181 ( .A1(n12063), .A2(n12062), .ZN(n12064) );
  AOI21_X1 U15182 ( .B1(n11280), .B2(n11270), .A(n11936), .ZN(n12067) );
  NAND2_X1 U15183 ( .A1(n12067), .A2(n12066), .ZN(n13386) );
  OR2_X1 U15184 ( .A1(n13386), .A2(n11275), .ZN(n15560) );
  INV_X1 U15185 ( .A(n20657), .ZN(n20515) );
  NAND2_X1 U15186 ( .A1(n20515), .A2(n12072), .ZN(n20676) );
  NAND2_X1 U15187 ( .A1(n20676), .A2(n20578), .ZN(n12068) );
  NAND2_X1 U15188 ( .A1(n20578), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12070) );
  NAND2_X1 U15189 ( .A1(n20468), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12069) );
  AND2_X1 U15190 ( .A1(n12070), .A2(n12069), .ZN(n19939) );
  INV_X1 U15191 ( .A(n19939), .ZN(n12071) );
  INV_X2 U15192 ( .A(n19823), .ZN(n19950) );
  NAND2_X1 U15193 ( .A1(n19950), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14587) );
  OAI21_X1 U15194 ( .B1(n19938), .B2(n14165), .A(n14587), .ZN(n12073) );
  AOI21_X1 U15195 ( .B1(n15781), .B2(n14172), .A(n12073), .ZN(n12074) );
  OAI21_X1 U15196 ( .B1(n14594), .B2(n19944), .A(n12074), .ZN(n12075) );
  INV_X1 U15197 ( .A(n12080), .ZN(n12101) );
  INV_X1 U15198 ( .A(n14869), .ZN(n12083) );
  INV_X1 U15199 ( .A(n12081), .ZN(n12082) );
  NAND2_X1 U15200 ( .A1(n12083), .A2(n12082), .ZN(n12084) );
  INV_X1 U15201 ( .A(n14001), .ZN(n14003) );
  NAND3_X1 U15202 ( .A1(n14795), .A2(n13031), .A3(n12088), .ZN(n12089) );
  NAND2_X1 U15203 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n18889), .ZN(n12092) );
  AOI22_X1 U15204 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18901), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n18890), .ZN(n12091) );
  OAI211_X1 U15205 ( .C1(n14003), .C2(n18888), .A(n12092), .B(n12091), .ZN(
        n12093) );
  INV_X1 U15206 ( .A(n12093), .ZN(n12094) );
  INV_X1 U15207 ( .A(n12104), .ZN(n12105) );
  INV_X1 U15208 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12103) );
  OAI21_X1 U15209 ( .B1(n12105), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n13589), .ZN(n14424) );
  AOI22_X1 U15210 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12110) );
  AOI22_X1 U15211 ( .A1(n9667), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n9673), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U15212 ( .A1(n12106), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11201), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15213 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11311), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12107) );
  NAND4_X1 U15214 ( .A1(n12110), .A2(n12109), .A3(n12108), .A4(n12107), .ZN(
        n12118) );
  AOI22_X1 U15215 ( .A1(n9651), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12130), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12116) );
  AOI22_X1 U15216 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U15217 ( .A1(n12111), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12114) );
  AOI22_X1 U15218 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11319), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12113) );
  NAND4_X1 U15219 ( .A1(n12116), .A2(n12115), .A3(n12114), .A4(n12113), .ZN(
        n12117) );
  NOR2_X1 U15220 ( .A1(n12118), .A2(n12117), .ZN(n12128) );
  NAND2_X1 U15221 ( .A1(n12120), .A2(n12119), .ZN(n12127) );
  XNOR2_X1 U15222 ( .A(n12128), .B(n12127), .ZN(n12124) );
  AOI21_X1 U15223 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20581), .A(
        n12150), .ZN(n12122) );
  NAND2_X1 U15224 ( .A1(n12155), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12121) );
  OAI211_X1 U15225 ( .C1(n12124), .C2(n12123), .A(n12122), .B(n12121), .ZN(
        n12125) );
  OAI21_X1 U15226 ( .B1(n11471), .B2(n14424), .A(n12125), .ZN(n14153) );
  NOR2_X1 U15227 ( .A1(n12128), .A2(n12127), .ZN(n12145) );
  AOI22_X1 U15228 ( .A1(n12130), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12129), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U15229 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9672), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15230 ( .A1(n11319), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11258), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12132) );
  AOI22_X1 U15231 ( .A1(n11320), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11311), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12131) );
  NAND4_X1 U15232 ( .A1(n12134), .A2(n12133), .A3(n12132), .A4(n12131), .ZN(
        n12143) );
  AOI22_X1 U15233 ( .A1(n12112), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11200), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U15234 ( .A1(n12135), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11336), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12140) );
  AOI22_X1 U15235 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11373), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U15236 ( .A1(n12137), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12136), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12138) );
  NAND4_X1 U15237 ( .A1(n12141), .A2(n12140), .A3(n12139), .A4(n12138), .ZN(
        n12142) );
  NOR2_X1 U15238 ( .A1(n12143), .A2(n12142), .ZN(n12144) );
  XNOR2_X1 U15239 ( .A(n12145), .B(n12144), .ZN(n12147) );
  NAND2_X1 U15240 ( .A1(n12147), .A2(n12146), .ZN(n12153) );
  NAND2_X1 U15241 ( .A1(n20581), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12148) );
  NAND2_X1 U15242 ( .A1(n11471), .A2(n12148), .ZN(n12149) );
  AOI21_X1 U15243 ( .B1(n12155), .B2(P1_EAX_REG_30__SCAN_IN), .A(n12149), .ZN(
        n12152) );
  XNOR2_X1 U15244 ( .A(n13589), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14412) );
  AOI22_X1 U15245 ( .A1(n12155), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12154), .ZN(n12156) );
  INV_X1 U15246 ( .A(n12156), .ZN(n12157) );
  NAND2_X1 U15247 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20677) );
  INV_X1 U15248 ( .A(n20677), .ZN(n20585) );
  OR2_X1 U15249 ( .A1(n13386), .A2(n13593), .ZN(n13436) );
  OAI21_X1 U15250 ( .B1(n12158), .B2(n20585), .A(n13436), .ZN(n12159) );
  INV_X1 U15251 ( .A(n12159), .ZN(n12160) );
  NOR3_X1 U15252 ( .A1(n12164), .A2(n12163), .A3(n12162), .ZN(n12166) );
  OAI21_X1 U15253 ( .B1(n12167), .B2(n12166), .A(n12165), .ZN(n13377) );
  NAND3_X1 U15254 ( .A1(n12168), .A2(n13377), .A3(n20677), .ZN(n12169) );
  NAND3_X1 U15255 ( .A1(n13416), .A2(n13236), .A3(n11231), .ZN(n12171) );
  OR2_X1 U15256 ( .A1(n12172), .A2(n12171), .ZN(n13227) );
  NOR2_X1 U15257 ( .A1(n13227), .A2(n13593), .ZN(n12173) );
  AND2_X1 U15258 ( .A1(n14401), .A2(n13236), .ZN(n12175) );
  NOR4_X1 U15259 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n12179) );
  NOR4_X1 U15260 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_ADDRESS_REG_19__SCAN_IN), .A3(P1_ADDRESS_REG_18__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n12178) );
  NOR4_X1 U15261 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n12177) );
  NOR4_X1 U15262 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n12176) );
  AND4_X1 U15263 ( .A1(n12179), .A2(n12178), .A3(n12177), .A4(n12176), .ZN(
        n12184) );
  NOR4_X1 U15264 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_2__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12182) );
  NOR4_X1 U15265 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(
        P1_ADDRESS_REG_23__SCAN_IN), .A3(P1_ADDRESS_REG_22__SCAN_IN), .A4(
        P1_ADDRESS_REG_21__SCAN_IN), .ZN(n12181) );
  NOR4_X1 U15266 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P1_ADDRESS_REG_27__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_25__SCAN_IN), .ZN(n12180) );
  INV_X1 U15267 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20604) );
  AND4_X1 U15268 ( .A1(n12182), .A2(n12181), .A3(n12180), .A4(n20604), .ZN(
        n12183) );
  NAND2_X1 U15269 ( .A1(n12184), .A2(n12183), .ZN(n12185) );
  AOI22_X1 U15270 ( .A1(n15747), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15744), .ZN(n12186) );
  INV_X1 U15271 ( .A(n12186), .ZN(n12188) );
  INV_X1 U15272 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19066) );
  NOR2_X1 U15273 ( .A1(n15751), .A2(n19066), .ZN(n12187) );
  NOR2_X1 U15274 ( .A1(n12188), .A2(n12187), .ZN(n12189) );
  NAND2_X1 U15275 ( .A1(n16208), .A2(n17636), .ZN(n17549) );
  NAND2_X1 U15276 ( .A1(n12192), .A2(n17537), .ZN(n12205) );
  INV_X1 U15277 ( .A(n17552), .ZN(n17454) );
  OR2_X1 U15278 ( .A1(n12193), .A2(n17454), .ZN(n12201) );
  INV_X1 U15279 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17639) );
  NAND4_X1 U15280 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16501) );
  NAND2_X1 U15281 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17487) );
  INV_X1 U15282 ( .A(n17487), .ZN(n17462) );
  NAND2_X1 U15283 ( .A1(n17462), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17436) );
  INV_X1 U15284 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n20831) );
  INV_X1 U15285 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17341) );
  NAND3_X1 U15286 ( .A1(n17330), .A2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17305) );
  INV_X1 U15287 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17304) );
  INV_X1 U15288 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16390) );
  INV_X1 U15289 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16368) );
  OAI21_X1 U15290 ( .B1(n18605), .B2(n18646), .A(n18586), .ZN(n18625) );
  INV_X1 U15291 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18630) );
  NOR2_X1 U15292 ( .A1(n18605), .A2(n18630), .ZN(n17541) );
  NOR2_X1 U15293 ( .A1(n12194), .A2(n16390), .ZN(n17275) );
  NAND2_X1 U15294 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17275), .ZN(
        n16198) );
  NOR2_X1 U15295 ( .A1(n16368), .A2(n16198), .ZN(n12195) );
  NAND2_X1 U15296 ( .A1(n18486), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17644) );
  NAND2_X1 U15297 ( .A1(n18478), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18599) );
  OAI221_X1 U15298 ( .B1(n18646), .B2(P3_STATE2_REG_1__SCAN_IN), .C1(
        P3_STATE2_REG_2__SCAN_IN), .C2(n18605), .A(n18599), .ZN(n17986) );
  NAND3_X1 U15299 ( .A1(n18646), .A2(n18586), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18324) );
  AOI21_X1 U15300 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17342), .A(
        n18364), .ZN(n17486) );
  NAND2_X1 U15301 ( .A1(n12195), .A2(n17407), .ZN(n16188) );
  XNOR2_X1 U15302 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12197) );
  INV_X1 U15303 ( .A(n17342), .ZN(n17384) );
  NOR2_X1 U15304 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17384), .ZN(
        n16195) );
  INV_X1 U15305 ( .A(n16349), .ZN(n12196) );
  OR2_X1 U15306 ( .A1(n18006), .A2(n12195), .ZN(n16199) );
  OAI211_X1 U15307 ( .C1(n12196), .C2(n17644), .A(n17643), .B(n16199), .ZN(
        n16202) );
  NOR2_X1 U15308 ( .A1(n16195), .A2(n16202), .ZN(n16187) );
  OAI22_X1 U15309 ( .A1(n16188), .A2(n12197), .B1(n16187), .B2(n9880), .ZN(
        n12198) );
  AOI211_X1 U15310 ( .C1(n9732), .C2(n17476), .A(n12199), .B(n12198), .ZN(
        n12200) );
  NAND2_X1 U15311 ( .A1(n12205), .A2(n12204), .ZN(P3_U2799) );
  INV_X1 U15312 ( .A(n12209), .ZN(n12215) );
  INV_X1 U15313 ( .A(n12214), .ZN(n12210) );
  NAND2_X1 U15314 ( .A1(n12215), .A2(n12210), .ZN(n12211) );
  NAND2_X1 U15315 ( .A1(n12215), .A2(n12601), .ZN(n12228) );
  AOI22_X1 U15316 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n13718), .B1(
        n12291), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12225) );
  INV_X1 U15317 ( .A(n12593), .ZN(n13222) );
  AOI22_X1 U15318 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19192), .B1(
        n19343), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12224) );
  INV_X1 U15319 ( .A(n12216), .ZN(n12217) );
  NOR2_X1 U15320 ( .A1(n9658), .A2(n12217), .ZN(n12233) );
  NOR2_X2 U15321 ( .A1(n12235), .A2(n12226), .ZN(n12279) );
  AOI22_X1 U15322 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12279), .B1(
        n19368), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12223) );
  INV_X1 U15323 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12219) );
  OAI21_X1 U15324 ( .B1(n12312), .B2(n12219), .A(n13720), .ZN(n12221) );
  INV_X1 U15325 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12786) );
  NOR2_X1 U15326 ( .A1(n12306), .A2(n12786), .ZN(n12220) );
  NOR2_X1 U15327 ( .A1(n12221), .A2(n12220), .ZN(n12222) );
  NAND4_X1 U15328 ( .A1(n12225), .A2(n12224), .A3(n12223), .A4(n12222), .ZN(
        n12244) );
  NOR2_X1 U15329 ( .A1(n12227), .A2(n12226), .ZN(n12278) );
  NOR2_X2 U15330 ( .A1(n12235), .A2(n12228), .ZN(n12289) );
  NAND2_X1 U15331 ( .A1(n12289), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12231) );
  NOR2_X2 U15332 ( .A1(n12235), .A2(n12229), .ZN(n12290) );
  NAND2_X1 U15333 ( .A1(n12290), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12230) );
  AOI22_X1 U15334 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n12281), .B1(
        n12311), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12239) );
  NOR2_X1 U15335 ( .A1(n12235), .A2(n12234), .ZN(n12280) );
  AOI22_X1 U15336 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12280), .B1(
        n19313), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12238) );
  NAND4_X1 U15337 ( .A1(n12241), .A2(n12240), .A3(n12239), .A4(n12238), .ZN(
        n12243) );
  INV_X1 U15338 ( .A(n13112), .ZN(n12444) );
  NAND2_X1 U15339 ( .A1(n12444), .A2(n12442), .ZN(n12448) );
  NAND2_X1 U15340 ( .A1(n12448), .A2(n12449), .ZN(n12242) );
  INV_X1 U15341 ( .A(n12306), .ZN(n12245) );
  AOI22_X1 U15342 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n13718), .B1(
        n12305), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15343 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12279), .B1(
        n19343), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15344 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19192), .B1(
        n12291), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12246) );
  NAND4_X1 U15345 ( .A1(n12249), .A2(n12248), .A3(n12247), .A4(n12246), .ZN(
        n12258) );
  AOI22_X1 U15346 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12278), .B1(
        n12290), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12253) );
  INV_X1 U15347 ( .A(n12312), .ZN(n12288) );
  AOI22_X1 U15348 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n12311), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15349 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12280), .B1(
        n12281), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U15350 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12289), .B1(
        n19313), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12250) );
  NAND4_X1 U15351 ( .A1(n12253), .A2(n12252), .A3(n12251), .A4(n12250), .ZN(
        n12257) );
  INV_X1 U15352 ( .A(n12254), .ZN(n12255) );
  NAND2_X1 U15353 ( .A1(n10264), .A2(n12255), .ZN(n12256) );
  XNOR2_X1 U15354 ( .A(n12260), .B(n12259), .ZN(n13760) );
  OAI21_X1 U15355 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19720), .A(
        n12261), .ZN(n12490) );
  MUX2_X1 U15356 ( .A(n12490), .B(n12443), .S(n12536), .Z(n12429) );
  MUX2_X1 U15357 ( .A(n12429), .B(n13123), .S(n10768), .Z(n18887) );
  NOR2_X1 U15358 ( .A1(n18887), .A2(n13020), .ZN(n12263) );
  NAND3_X1 U15359 ( .A1(n10768), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n12262) );
  NAND2_X1 U15360 ( .A1(n12263), .A2(n10079), .ZN(n12264) );
  XOR2_X1 U15361 ( .A(n12263), .B(n10079), .Z(n13019) );
  NAND2_X1 U15362 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13019), .ZN(
        n13018) );
  NAND2_X1 U15363 ( .A1(n12264), .A2(n13018), .ZN(n12268) );
  XNOR2_X1 U15364 ( .A(n12266), .B(n12265), .ZN(n13822) );
  XOR2_X1 U15365 ( .A(n12553), .B(n12268), .Z(n13201) );
  NOR2_X1 U15366 ( .A1(n13822), .A2(n13201), .ZN(n12267) );
  AOI21_X1 U15367 ( .B1(n12268), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n12267), .ZN(n13571) );
  INV_X1 U15368 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13830) );
  XNOR2_X1 U15369 ( .A(n12270), .B(n12269), .ZN(n18862) );
  INV_X1 U15370 ( .A(n18862), .ZN(n12271) );
  NAND2_X1 U15371 ( .A1(n12271), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12272) );
  NAND2_X1 U15372 ( .A1(n13839), .A2(n12272), .ZN(n13920) );
  INV_X1 U15373 ( .A(n12273), .ZN(n12276) );
  INV_X1 U15374 ( .A(n12274), .ZN(n12275) );
  AOI22_X1 U15375 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n13718), .B1(
        n12278), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12287) );
  AOI22_X1 U15376 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19192), .B1(
        n12279), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U15377 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19133), .B1(
        n12281), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12285) );
  INV_X1 U15378 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12282) );
  INV_X1 U15379 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12882) );
  OAI22_X1 U15380 ( .A1(n12282), .A2(n19372), .B1(n12306), .B2(n12882), .ZN(
        n12283) );
  INV_X1 U15381 ( .A(n12283), .ZN(n12284) );
  AOI22_X1 U15382 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n12311), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12295) );
  AOI22_X1 U15383 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n12289), .B1(
        n19313), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12294) );
  AOI22_X1 U15384 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n12290), .B1(
        n12305), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15385 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n12291), .B1(
        n19343), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12292) );
  NAND2_X1 U15386 ( .A1(n10075), .A2(n10094), .ZN(n12298) );
  NAND2_X1 U15387 ( .A1(n12296), .A2(n10264), .ZN(n12297) );
  INV_X1 U15388 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15398) );
  XNOR2_X1 U15389 ( .A(n12303), .B(n15398), .ZN(n13918) );
  NAND2_X1 U15390 ( .A1(n13920), .A2(n13918), .ZN(n13919) );
  NAND2_X1 U15391 ( .A1(n12303), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12304) );
  NAND2_X1 U15392 ( .A1(n13919), .A2(n12304), .ZN(n15377) );
  AOI22_X1 U15393 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19192), .B1(
        n12291), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12310) );
  AOI22_X1 U15394 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n13718), .B1(
        n12305), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U15395 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12279), .B1(
        n19343), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12308) );
  AOI22_X1 U15396 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19368), .B1(
        n12245), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12307) );
  NAND4_X1 U15397 ( .A1(n12310), .A2(n12309), .A3(n12308), .A4(n12307), .ZN(
        n12320) );
  AOI22_X1 U15398 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12278), .B1(
        n12290), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12318) );
  AOI22_X1 U15399 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19133), .B1(
        n12281), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U15400 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12289), .B1(
        n19313), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12316) );
  INV_X1 U15401 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12313) );
  INV_X1 U15402 ( .A(n12311), .ZN(n19535) );
  INV_X1 U15403 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12895) );
  OAI22_X1 U15404 ( .A1(n12313), .A2(n19535), .B1(n12312), .B2(n12895), .ZN(
        n12314) );
  INV_X1 U15405 ( .A(n12314), .ZN(n12315) );
  NAND4_X1 U15406 ( .A1(n12318), .A2(n12317), .A3(n12316), .A4(n12315), .ZN(
        n12319) );
  NAND2_X1 U15407 ( .A1(n12321), .A2(n10264), .ZN(n12322) );
  NAND2_X1 U15408 ( .A1(n12464), .A2(n14002), .ZN(n12326) );
  INV_X1 U15409 ( .A(n12325), .ZN(n12329) );
  XNOR2_X1 U15410 ( .A(n12324), .B(n12329), .ZN(n18830) );
  NAND2_X1 U15411 ( .A1(n12326), .A2(n18830), .ZN(n12327) );
  INV_X1 U15412 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15383) );
  XNOR2_X1 U15413 ( .A(n12327), .B(n15383), .ZN(n15376) );
  NAND2_X1 U15414 ( .A1(n12327), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12328) );
  NAND2_X1 U15415 ( .A1(n12324), .A2(n12329), .ZN(n12332) );
  INV_X1 U15416 ( .A(n12330), .ZN(n12331) );
  XNOR2_X1 U15417 ( .A(n12332), .B(n12331), .ZN(n18823) );
  INV_X1 U15418 ( .A(n18823), .ZN(n12333) );
  INV_X1 U15419 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15069) );
  NAND2_X1 U15420 ( .A1(n12333), .A2(n15069), .ZN(n16063) );
  INV_X1 U15421 ( .A(n12334), .ZN(n12335) );
  XNOR2_X1 U15422 ( .A(n12336), .B(n12335), .ZN(n18809) );
  AND2_X1 U15423 ( .A1(n18809), .A2(n14000), .ZN(n16064) );
  INV_X1 U15424 ( .A(n12342), .ZN(n12340) );
  NAND2_X1 U15425 ( .A1(n10768), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12338) );
  MUX2_X1 U15426 ( .A(n12338), .B(n10768), .S(n12337), .Z(n12339) );
  AOI21_X1 U15427 ( .B1(n18798), .B2(n14000), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15343) );
  NOR2_X1 U15428 ( .A1(n12342), .A2(n12341), .ZN(n12343) );
  NAND2_X1 U15429 ( .A1(n10768), .A2(n12343), .ZN(n12344) );
  AND2_X1 U15430 ( .A1(n12405), .A2(n12344), .ZN(n12345) );
  NAND2_X1 U15431 ( .A1(n12346), .A2(n12345), .ZN(n18790) );
  OR2_X1 U15432 ( .A1(n18790), .A2(n14002), .ZN(n12353) );
  INV_X1 U15433 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15333) );
  NAND2_X1 U15434 ( .A1(n12353), .A2(n15333), .ZN(n15325) );
  NAND2_X1 U15435 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n12346), .ZN(n12347) );
  NOR2_X1 U15436 ( .A1(n10234), .A2(n12347), .ZN(n12348) );
  NOR2_X1 U15437 ( .A1(n12349), .A2(n12348), .ZN(n18775) );
  AOI21_X1 U15438 ( .B1(n18775), .B2(n14000), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15309) );
  INV_X1 U15439 ( .A(n15309), .ZN(n12350) );
  INV_X1 U15440 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n20698) );
  NOR2_X1 U15441 ( .A1(n14002), .A2(n20698), .ZN(n12351) );
  NAND2_X1 U15442 ( .A1(n18775), .A2(n12351), .ZN(n15307) );
  INV_X1 U15443 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15348) );
  NOR2_X1 U15444 ( .A1(n14002), .A2(n15348), .ZN(n12352) );
  NAND2_X1 U15445 ( .A1(n18798), .A2(n12352), .ZN(n15327) );
  OR2_X1 U15446 ( .A1(n15333), .A2(n12353), .ZN(n15324) );
  AND2_X1 U15447 ( .A1(n15307), .A2(n10093), .ZN(n15283) );
  OR2_X1 U15448 ( .A1(n12355), .A2(n12354), .ZN(n12356) );
  NAND2_X1 U15449 ( .A1(n12359), .A2(n12356), .ZN(n18764) );
  INV_X1 U15450 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15300) );
  OR3_X1 U15451 ( .A1(n18764), .A2(n14002), .A3(n15300), .ZN(n15284) );
  AND2_X1 U15452 ( .A1(n15283), .A2(n15284), .ZN(n14998) );
  OR2_X1 U15453 ( .A1(n18764), .A2(n14002), .ZN(n12357) );
  NAND2_X1 U15454 ( .A1(n12359), .A2(n12358), .ZN(n12360) );
  NAND2_X1 U15455 ( .A1(n9692), .A2(n12360), .ZN(n18753) );
  INV_X1 U15456 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15274) );
  NAND2_X1 U15457 ( .A1(n12390), .A2(n15274), .ZN(n15265) );
  NAND2_X1 U15458 ( .A1(n10768), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12361) );
  MUX2_X1 U15459 ( .A(n12361), .B(n10768), .S(n12364), .Z(n12363) );
  INV_X1 U15460 ( .A(n12384), .ZN(n12362) );
  NAND2_X1 U15461 ( .A1(n12363), .A2(n12362), .ZN(n12393) );
  INV_X1 U15462 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15172) );
  OAI21_X1 U15463 ( .B1(n12393), .B2(n14002), .A(n15172), .ZN(n15030) );
  INV_X1 U15464 ( .A(n12364), .ZN(n12367) );
  INV_X1 U15465 ( .A(n12374), .ZN(n12365) );
  NAND2_X1 U15466 ( .A1(n12365), .A2(n13941), .ZN(n12369) );
  NAND3_X1 U15467 ( .A1(n12369), .A2(P2_EBX_REG_19__SCAN_IN), .A3(n10768), 
        .ZN(n12366) );
  NAND2_X1 U15468 ( .A1(n12367), .A2(n12366), .ZN(n18686) );
  OR2_X1 U15469 ( .A1(n18686), .A2(n14002), .ZN(n12386) );
  INV_X1 U15470 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15189) );
  NAND2_X1 U15471 ( .A1(n12386), .A2(n15189), .ZN(n15039) );
  NAND2_X1 U15472 ( .A1(n12374), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12368) );
  MUX2_X1 U15473 ( .A(n12368), .B(n12374), .S(n10234), .Z(n12370) );
  NAND2_X1 U15474 ( .A1(n12370), .A2(n12369), .ZN(n18698) );
  INV_X1 U15475 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15205) );
  OAI21_X1 U15476 ( .B1(n18698), .B2(n14002), .A(n15205), .ZN(n15041) );
  AND2_X1 U15477 ( .A1(n15039), .A2(n15041), .ZN(n15027) );
  AND2_X1 U15478 ( .A1(n15030), .A2(n15027), .ZN(n15013) );
  NAND2_X1 U15479 ( .A1(n12372), .A2(n12371), .ZN(n12373) );
  AND2_X1 U15480 ( .A1(n12374), .A2(n12373), .ZN(n18708) );
  AOI21_X1 U15481 ( .B1(n18708), .B2(n14000), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15010) );
  NAND3_X1 U15482 ( .A1(n12376), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n10768), 
        .ZN(n12375) );
  OAI211_X1 U15483 ( .C1(n12376), .C2(P2_EBX_REG_16__SCAN_IN), .A(n12375), .B(
        n12405), .ZN(n18719) );
  INV_X1 U15484 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n20838) );
  OAI21_X1 U15485 ( .B1(n18719), .B2(n14002), .A(n20838), .ZN(n12377) );
  OR3_X1 U15486 ( .A1(n18719), .A2(n14002), .A3(n20838), .ZN(n15005) );
  NAND2_X1 U15487 ( .A1(n12377), .A2(n15005), .ZN(n15229) );
  INV_X1 U15488 ( .A(n12378), .ZN(n12379) );
  XNOR2_X1 U15489 ( .A(n9692), .B(n12379), .ZN(n18740) );
  AOI21_X1 U15490 ( .B1(n18740), .B2(n14000), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14999) );
  XNOR2_X1 U15491 ( .A(n12381), .B(n9999), .ZN(n18731) );
  NAND2_X1 U15492 ( .A1(n18731), .A2(n14000), .ZN(n12382) );
  INV_X1 U15493 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12973) );
  NOR4_X1 U15494 ( .A1(n15010), .A2(n15229), .A3(n14999), .A4(n15002), .ZN(
        n12385) );
  NAND2_X1 U15495 ( .A1(n10768), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12383) );
  OAI211_X1 U15496 ( .C1(n12384), .C2(n12383), .A(n12405), .B(n12399), .ZN(
        n14770) );
  OAI21_X1 U15497 ( .B1(n14770), .B2(n14002), .A(n9617), .ZN(n15015) );
  NAND3_X1 U15498 ( .A1(n15013), .A2(n12385), .A3(n15015), .ZN(n12397) );
  NOR3_X1 U15499 ( .A1(n14770), .A2(n14002), .A3(n9617), .ZN(n15014) );
  NOR3_X1 U15500 ( .A1(n18698), .A2(n14002), .A3(n15205), .ZN(n15050) );
  NOR2_X1 U15501 ( .A1(n12386), .A2(n15189), .ZN(n15011) );
  NOR2_X1 U15502 ( .A1(n14002), .A2(n12973), .ZN(n12387) );
  AND2_X1 U15503 ( .A1(n18731), .A2(n12387), .ZN(n12968) );
  INV_X1 U15504 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15244) );
  NOR2_X1 U15505 ( .A1(n14002), .A2(n15244), .ZN(n12388) );
  AND2_X1 U15506 ( .A1(n18740), .A2(n12388), .ZN(n12967) );
  NOR2_X1 U15507 ( .A1(n12968), .A2(n12967), .ZN(n15003) );
  INV_X1 U15508 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15221) );
  NOR2_X1 U15509 ( .A1(n14002), .A2(n15221), .ZN(n12389) );
  NAND2_X1 U15510 ( .A1(n18708), .A2(n12389), .ZN(n15008) );
  INV_X1 U15511 ( .A(n12390), .ZN(n12391) );
  NAND2_X1 U15512 ( .A1(n12391), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15266) );
  NAND4_X1 U15513 ( .A1(n15003), .A2(n15008), .A3(n15005), .A4(n15266), .ZN(
        n12392) );
  NOR4_X1 U15514 ( .A1(n15014), .A2(n15050), .A3(n15011), .A4(n12392), .ZN(
        n12395) );
  INV_X1 U15515 ( .A(n12393), .ZN(n14788) );
  NOR2_X1 U15516 ( .A1(n14002), .A2(n15172), .ZN(n12394) );
  NAND2_X1 U15517 ( .A1(n14788), .A2(n12394), .ZN(n15029) );
  NAND2_X1 U15518 ( .A1(n12399), .A2(n10008), .ZN(n12400) );
  NAND2_X1 U15519 ( .A1(n12401), .A2(n12400), .ZN(n14757) );
  INV_X1 U15520 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16001) );
  OAI21_X1 U15521 ( .B1(n14757), .B2(n14002), .A(n16001), .ZN(n15997) );
  NOR3_X1 U15522 ( .A1(n14757), .A2(n14002), .A3(n16001), .ZN(n15996) );
  AOI21_X1 U15523 ( .B1(n12402), .B2(n12401), .A(n9700), .ZN(n12995) );
  NAND2_X1 U15524 ( .A1(n12995), .A2(n14000), .ZN(n12403) );
  XOR2_X1 U15525 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n12403), .Z(
        n14989) );
  NAND3_X1 U15526 ( .A1(n12995), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n14000), .ZN(n12404) );
  AND2_X1 U15527 ( .A1(n12405), .A2(n14000), .ZN(n14979) );
  NAND2_X1 U15528 ( .A1(n14979), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12406) );
  INV_X1 U15529 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12557) );
  INV_X1 U15530 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15116) );
  NAND2_X1 U15531 ( .A1(n14036), .A2(n15116), .ZN(n14965) );
  NAND2_X1 U15532 ( .A1(n10768), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12407) );
  OR2_X1 U15533 ( .A1(n15953), .A2(n12407), .ZN(n12408) );
  INV_X1 U15534 ( .A(n15945), .ZN(n12410) );
  NOR2_X1 U15535 ( .A1(n12410), .A2(n14002), .ZN(n12411) );
  NAND3_X1 U15536 ( .A1(n15945), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14000), .ZN(n12412) );
  OR2_X1 U15537 ( .A1(n14036), .A2(n15116), .ZN(n14966) );
  NAND2_X1 U15538 ( .A1(n12412), .A2(n14966), .ZN(n13997) );
  INV_X1 U15539 ( .A(n12413), .ZN(n12416) );
  INV_X1 U15540 ( .A(n12414), .ZN(n12415) );
  NAND2_X1 U15541 ( .A1(n12416), .A2(n12415), .ZN(n12417) );
  NAND2_X1 U15542 ( .A1(n12423), .A2(n12417), .ZN(n13007) );
  XNOR2_X1 U15543 ( .A(n12418), .B(n13990), .ZN(n14946) );
  INV_X1 U15544 ( .A(n12418), .ZN(n12419) );
  AOI22_X1 U15545 ( .A1(n14946), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n13990), .B2(n12419), .ZN(n12426) );
  INV_X1 U15546 ( .A(n12421), .ZN(n12422) );
  NAND2_X1 U15547 ( .A1(n12423), .A2(n12422), .ZN(n12424) );
  NAND2_X1 U15548 ( .A1(n12420), .A2(n12424), .ZN(n15936) );
  INV_X1 U15549 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n20693) );
  XNOR2_X1 U15550 ( .A(n13993), .B(n20693), .ZN(n12425) );
  XNOR2_X1 U15551 ( .A(n12426), .B(n12425), .ZN(n12537) );
  INV_X1 U15552 ( .A(n12489), .ZN(n12428) );
  OAI21_X1 U15553 ( .B1(n12429), .B2(n12428), .A(n12427), .ZN(n12430) );
  INV_X1 U15554 ( .A(n12503), .ZN(n12507) );
  AOI21_X1 U15555 ( .B1(n12430), .B2(n12502), .A(n12507), .ZN(n19727) );
  OAI21_X1 U15556 ( .B1(n12490), .B2(n12431), .A(n16131), .ZN(n12436) );
  INV_X1 U15557 ( .A(n12432), .ZN(n12435) );
  NAND2_X1 U15558 ( .A1(n13139), .A2(n12433), .ZN(n13136) );
  INV_X1 U15559 ( .A(n13136), .ZN(n12434) );
  AOI21_X1 U15560 ( .B1(n12435), .B2(n12434), .A(P2_FLUSH_REG_SCAN_IN), .ZN(
        n19714) );
  MUX2_X1 U15561 ( .A(n12436), .B(n19714), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n15589) );
  MUX2_X1 U15562 ( .A(n19727), .B(n19725), .S(n13720), .Z(n12440) );
  NAND2_X1 U15563 ( .A1(n19742), .A2(n19598), .ZN(n12438) );
  NOR2_X1 U15564 ( .A1(n12437), .A2(n12438), .ZN(n12439) );
  INV_X1 U15565 ( .A(n18659), .ZN(n12441) );
  NAND2_X1 U15566 ( .A1(n12537), .A2(n19013), .ZN(n12488) );
  XNOR2_X1 U15567 ( .A(n12443), .B(n12442), .ZN(n12446) );
  NOR2_X1 U15568 ( .A1(n12444), .A2(n13020), .ZN(n12445) );
  NAND2_X1 U15569 ( .A1(n12446), .A2(n12445), .ZN(n12447) );
  XOR2_X1 U15570 ( .A(n12446), .B(n12445), .Z(n13022) );
  NAND2_X1 U15571 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13022), .ZN(
        n13021) );
  NAND2_X1 U15572 ( .A1(n12447), .A2(n13021), .ZN(n12450) );
  XNOR2_X1 U15573 ( .A(n12553), .B(n12450), .ZN(n13204) );
  XNOR2_X1 U15574 ( .A(n12449), .B(n12448), .ZN(n13203) );
  NAND2_X1 U15575 ( .A1(n13204), .A2(n13203), .ZN(n13202) );
  NAND2_X1 U15576 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12450), .ZN(
        n12451) );
  NAND2_X1 U15577 ( .A1(n13202), .A2(n12451), .ZN(n12452) );
  XNOR2_X1 U15578 ( .A(n12452), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13574) );
  NAND2_X1 U15579 ( .A1(n12452), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12453) );
  XNOR2_X1 U15580 ( .A(n12455), .B(n12454), .ZN(n12457) );
  INV_X1 U15581 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15397) );
  NAND2_X1 U15582 ( .A1(n9654), .A2(n12457), .ZN(n12458) );
  AND2_X1 U15583 ( .A1(n12459), .A2(n15398), .ZN(n13915) );
  INV_X1 U15584 ( .A(n12464), .ZN(n12463) );
  AOI21_X1 U15585 ( .B1(n9646), .B2(n12463), .A(n10074), .ZN(n12462) );
  NAND2_X1 U15586 ( .A1(n12465), .A2(n12464), .ZN(n12466) );
  XNOR2_X1 U15587 ( .A(n12469), .B(n14000), .ZN(n15070) );
  NAND2_X1 U15588 ( .A1(n12471), .A2(n14000), .ZN(n12470) );
  NAND3_X1 U15589 ( .A1(n12471), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n14000), .ZN(n12472) );
  AND2_X1 U15590 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15242) );
  NAND2_X1 U15591 ( .A1(n15242), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12978) );
  NAND3_X1 U15592 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12974) );
  NOR2_X1 U15593 ( .A1(n12978), .A2(n12974), .ZN(n12972) );
  NOR3_X1 U15594 ( .A1(n20838), .A2(n12973), .A3(n15221), .ZN(n15054) );
  NAND2_X1 U15595 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15054), .ZN(
        n15171) );
  INV_X1 U15596 ( .A(n15171), .ZN(n12473) );
  AND2_X1 U15597 ( .A1(n12972), .A2(n12473), .ZN(n15173) );
  AND2_X1 U15598 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12474) );
  AND2_X1 U15599 ( .A1(n15173), .A2(n12474), .ZN(n15164) );
  INV_X1 U15600 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14948) );
  NOR2_X2 U15601 ( .A1(n18659), .A2(n13720), .ZN(n19015) );
  INV_X1 U15602 ( .A(n14025), .ZN(n12476) );
  OAI21_X1 U15603 ( .B1(n13008), .B2(n12477), .A(n12476), .ZN(n15941) );
  INV_X1 U15604 ( .A(n15941), .ZN(n12484) );
  NAND2_X1 U15605 ( .A1(n19601), .A2(n19732), .ZN(n19685) );
  INV_X1 U15606 ( .A(n19685), .ZN(n19600) );
  OR2_X1 U15607 ( .A1(n19688), .A2(n19600), .ZN(n19712) );
  NAND2_X1 U15608 ( .A1(n19712), .A2(n19741), .ZN(n12478) );
  AND2_X1 U15609 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19702) );
  INV_X1 U15610 ( .A(n12600), .ZN(n12480) );
  NAND2_X1 U15611 ( .A1(n19682), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12479) );
  NAND2_X1 U15612 ( .A1(n12480), .A2(n12479), .ZN(n13115) );
  INV_X1 U15613 ( .A(n19011), .ZN(n18847) );
  NAND2_X1 U15614 ( .A1(n19011), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12566) );
  NAND2_X1 U15615 ( .A1(n19012), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12481) );
  OAI211_X1 U15616 ( .C1(n19025), .C2(n12482), .A(n12566), .B(n12481), .ZN(
        n12483) );
  AOI21_X1 U15617 ( .B1(n12484), .B2(n16067), .A(n12483), .ZN(n12485) );
  NAND2_X1 U15618 ( .A1(n12487), .A2(n12488), .ZN(P2_U2986) );
  OAI21_X1 U15619 ( .B1(n12490), .B2(n12428), .A(n12536), .ZN(n12494) );
  INV_X1 U15620 ( .A(n12490), .ZN(n12492) );
  OAI211_X1 U15621 ( .C1(n13720), .C2(n12492), .A(n19027), .B(n12491), .ZN(
        n12493) );
  OAI211_X1 U15622 ( .C1(n12496), .C2(n12495), .A(n12494), .B(n12493), .ZN(
        n12501) );
  INV_X1 U15623 ( .A(n13111), .ZN(n19743) );
  NAND2_X1 U15624 ( .A1(n19743), .A2(n13720), .ZN(n12498) );
  MUX2_X1 U15625 ( .A(n12498), .B(n10766), .S(n12497), .Z(n12500) );
  INV_X1 U15626 ( .A(n12502), .ZN(n12499) );
  AOI21_X1 U15627 ( .B1(n12501), .B2(n12500), .A(n12499), .ZN(n12505) );
  NOR2_X1 U15628 ( .A1(n12502), .A2(n12536), .ZN(n12504) );
  OAI21_X1 U15629 ( .B1(n12505), .B2(n12504), .A(n12503), .ZN(n12506) );
  MUX2_X1 U15630 ( .A(n12506), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19741), .Z(n12510) );
  NAND2_X1 U15631 ( .A1(n12507), .A2(n13111), .ZN(n12508) );
  INV_X1 U15632 ( .A(n16139), .ZN(n13129) );
  NAND3_X1 U15633 ( .A1(n13131), .A2(n12509), .A3(n13129), .ZN(n12534) );
  INV_X1 U15634 ( .A(n13131), .ZN(n12512) );
  AOI21_X1 U15635 ( .B1(n12510), .B2(n19027), .A(n10259), .ZN(n12511) );
  NAND2_X1 U15636 ( .A1(n12512), .A2(n12511), .ZN(n12533) );
  NOR2_X1 U15637 ( .A1(n19027), .A2(n13720), .ZN(n12518) );
  INV_X1 U15638 ( .A(n12518), .ZN(n12513) );
  NOR2_X1 U15639 ( .A1(n12437), .A2(n12513), .ZN(n19723) );
  NAND2_X1 U15640 ( .A1(n12514), .A2(n12515), .ZN(n12516) );
  NAND2_X1 U15641 ( .A1(n10760), .A2(n12516), .ZN(n12527) );
  INV_X1 U15642 ( .A(n10271), .ZN(n12943) );
  OR2_X1 U15643 ( .A1(n12517), .A2(n12943), .ZN(n12519) );
  NAND2_X1 U15644 ( .A1(n12519), .A2(n12518), .ZN(n12547) );
  NAND3_X1 U15645 ( .A1(n10412), .A2(n16131), .A3(n13129), .ZN(n12525) );
  OAI21_X1 U15646 ( .B1(n10259), .B2(n13720), .A(n19027), .ZN(n12520) );
  NAND2_X1 U15647 ( .A1(n12520), .A2(n10271), .ZN(n12522) );
  AOI21_X1 U15648 ( .B1(n12522), .B2(n12515), .A(n12541), .ZN(n12524) );
  AND4_X1 U15649 ( .A1(n12547), .A2(n12525), .A3(n12524), .A4(n12523), .ZN(
        n12526) );
  AND2_X1 U15650 ( .A1(n12527), .A2(n12526), .ZN(n13125) );
  MUX2_X1 U15651 ( .A(n10412), .B(n12509), .S(n10264), .Z(n12528) );
  NAND3_X1 U15652 ( .A1(n12528), .A2(n16131), .A3(n19740), .ZN(n12530) );
  INV_X1 U15653 ( .A(n12437), .ZN(n16157) );
  NAND3_X1 U15654 ( .A1(n16157), .A2(n13720), .A3(n19725), .ZN(n12529) );
  NAND3_X1 U15655 ( .A1(n13125), .A2(n12530), .A3(n12529), .ZN(n12531) );
  AOI21_X1 U15656 ( .B1(n19727), .B2(n19723), .A(n12531), .ZN(n12532) );
  NAND3_X1 U15657 ( .A1(n12534), .A2(n12533), .A3(n12532), .ZN(n12535) );
  NAND2_X1 U15658 ( .A1(n16157), .A2(n12536), .ZN(n19724) );
  NAND2_X1 U15659 ( .A1(n12537), .A2(n16102), .ZN(n12584) );
  NAND3_X1 U15660 ( .A1(n10254), .A2(n12541), .A3(n12539), .ZN(n12544) );
  INV_X1 U15661 ( .A(n12540), .ZN(n13034) );
  OR2_X1 U15662 ( .A1(n10270), .A2(n12541), .ZN(n12542) );
  AOI22_X1 U15663 ( .A1(n13034), .A2(n12542), .B1(n19742), .B2(n12509), .ZN(
        n12543) );
  NAND3_X1 U15664 ( .A1(n12538), .A2(n12544), .A3(n12543), .ZN(n12549) );
  NAND2_X1 U15665 ( .A1(n12545), .A2(n13720), .ZN(n15414) );
  AOI21_X1 U15666 ( .B1(n15414), .B2(n12547), .A(n12546), .ZN(n12548) );
  OR2_X1 U15667 ( .A1(n12549), .A2(n12548), .ZN(n16114) );
  NOR2_X1 U15668 ( .A1(n16114), .A2(n10291), .ZN(n12550) );
  NAND3_X1 U15669 ( .A1(n10264), .A2(n12515), .A3(n10234), .ZN(n12552) );
  OR2_X1 U15670 ( .A1(n12551), .A2(n12552), .ZN(n15434) );
  OR2_X1 U15671 ( .A1(n12578), .A2(n15434), .ZN(n13281) );
  NAND2_X1 U15672 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13287) );
  OR2_X1 U15673 ( .A1(n12553), .A2(n13287), .ZN(n12554) );
  NAND2_X1 U15674 ( .A1(n15434), .A2(n12554), .ZN(n12555) );
  NAND2_X1 U15675 ( .A1(n15366), .A2(n12555), .ZN(n16099) );
  INV_X1 U15676 ( .A(n13287), .ZN(n13290) );
  NOR2_X1 U15677 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13290), .ZN(
        n13834) );
  NOR2_X1 U15678 ( .A1(n15398), .A2(n15397), .ZN(n15396) );
  NAND2_X1 U15679 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15396), .ZN(
        n15365) );
  NOR4_X1 U15680 ( .A1(n13834), .A2(n15383), .A3(n15069), .A4(n15365), .ZN(
        n16092) );
  NAND2_X1 U15681 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n16092), .ZN(
        n12567) );
  AND2_X1 U15682 ( .A1(n15164), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12556) );
  INV_X1 U15683 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15153) );
  NOR3_X1 U15684 ( .A1(n12557), .A2(n15153), .A3(n16001), .ZN(n12572) );
  NAND2_X1 U15685 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12573) );
  OR2_X1 U15686 ( .A1(n15131), .A2(n12573), .ZN(n12575) );
  NOR2_X1 U15687 ( .A1(n12575), .A2(n14948), .ZN(n15094) );
  INV_X1 U15688 ( .A(n16173), .ZN(n12558) );
  OR2_X1 U15689 ( .A1(n12559), .A2(n12558), .ZN(n16145) );
  AOI21_X1 U15690 ( .B1(n16145), .B2(n10264), .A(n12560), .ZN(n12561) );
  AOI21_X1 U15691 ( .B1(n12562), .B2(n9711), .A(n14867), .ZN(n15939) );
  NOR2_X1 U15692 ( .A1(n12563), .A2(n12551), .ZN(n16130) );
  AOI21_X1 U15693 ( .B1(n13720), .B2(n16133), .A(n16130), .ZN(n12564) );
  NAND2_X1 U15694 ( .A1(n15939), .A2(n15410), .ZN(n12565) );
  OAI211_X1 U15695 ( .C1(n15941), .C2(n15404), .A(n12566), .B(n12565), .ZN(
        n12577) );
  NAND2_X1 U15696 ( .A1(n15366), .A2(n12567), .ZN(n12569) );
  AND2_X1 U15697 ( .A1(n12578), .A2(n18831), .ZN(n12571) );
  AOI21_X1 U15698 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n13290), .A(
        n15213), .ZN(n12568) );
  NOR2_X1 U15699 ( .A1(n12571), .A2(n12568), .ZN(n13576) );
  INV_X1 U15700 ( .A(n15316), .ZN(n15347) );
  NAND2_X1 U15701 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15164), .ZN(
        n12570) );
  NOR2_X1 U15702 ( .A1(n15347), .A2(n12570), .ZN(n16081) );
  INV_X1 U15703 ( .A(n12571), .ZN(n13288) );
  AND2_X1 U15704 ( .A1(n15367), .A2(n13288), .ZN(n15315) );
  AOI21_X1 U15705 ( .B1(n16081), .B2(n12572), .A(n15315), .ZN(n15141) );
  AOI21_X1 U15706 ( .B1(n12574), .B2(n12573), .A(n15141), .ZN(n14042) );
  INV_X1 U15707 ( .A(n14042), .ZN(n15123) );
  NOR2_X1 U15708 ( .A1(n12575), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15110) );
  NOR2_X1 U15709 ( .A1(n15123), .A2(n15110), .ZN(n15097) );
  NOR2_X1 U15710 ( .A1(n15097), .A2(n20693), .ZN(n12576) );
  AOI211_X1 U15711 ( .C1(n15094), .C2(n20693), .A(n12577), .B(n12576), .ZN(
        n12582) );
  INV_X1 U15712 ( .A(n12578), .ZN(n12579) );
  OR2_X1 U15713 ( .A1(n12580), .A2(n15413), .ZN(n12581) );
  NAND2_X1 U15714 ( .A1(n12584), .A2(n12583), .ZN(P2_U3018) );
  NAND2_X1 U15715 ( .A1(n19057), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12585) );
  NAND2_X1 U15716 ( .A1(n12585), .A2(n19732), .ZN(n12602) );
  NOR2_X1 U15717 ( .A1(n19700), .A2(n19710), .ZN(n19536) );
  NAND2_X1 U15718 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19536), .ZN(
        n12594) );
  INV_X1 U15719 ( .A(n12594), .ZN(n12586) );
  NAND2_X1 U15720 ( .A1(n12586), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19534) );
  INV_X1 U15721 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19693) );
  NAND2_X1 U15722 ( .A1(n19693), .A2(n12594), .ZN(n12587) );
  AND3_X1 U15723 ( .A1(n19534), .A2(n19688), .A3(n12587), .ZN(n19425) );
  AOI21_X1 U15724 ( .B1(n12602), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19425), .ZN(n12588) );
  NOR2_X1 U15725 ( .A1(n12616), .A2(n12590), .ZN(n12591) );
  NAND2_X1 U15726 ( .A1(n12614), .A2(n12591), .ZN(n13300) );
  NAND2_X1 U15727 ( .A1(n12593), .A2(n12600), .ZN(n12597) );
  NAND2_X1 U15728 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19397) );
  NAND2_X1 U15729 ( .A1(n19397), .A2(n19700), .ZN(n12595) );
  AND2_X1 U15730 ( .A1(n12595), .A2(n12594), .ZN(n19188) );
  AOI22_X1 U15731 ( .A1(n12602), .A2(n19681), .B1(n19688), .B2(n19188), .ZN(
        n12596) );
  NAND2_X1 U15732 ( .A1(n12869), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12609) );
  NAND2_X1 U15733 ( .A1(n12602), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12598) );
  NAND2_X1 U15734 ( .A1(n19710), .A2(n19720), .ZN(n19306) );
  AND2_X1 U15735 ( .A1(n19397), .A2(n19306), .ZN(n19189) );
  NAND2_X1 U15736 ( .A1(n19189), .A2(n19688), .ZN(n19370) );
  NAND2_X1 U15737 ( .A1(n12598), .A2(n19370), .ZN(n12599) );
  AOI22_X1 U15738 ( .A1(n12602), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19688), .B2(n19720), .ZN(n12603) );
  NAND2_X1 U15739 ( .A1(n12869), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12606) );
  NAND2_X1 U15740 ( .A1(n13148), .A2(n13149), .ZN(n13151) );
  INV_X1 U15741 ( .A(n12605), .ZN(n12607) );
  NAND2_X1 U15742 ( .A1(n12607), .A2(n12606), .ZN(n12608) );
  NAND2_X1 U15743 ( .A1(n13220), .A2(n13219), .ZN(n13218) );
  INV_X1 U15744 ( .A(n12609), .ZN(n12610) );
  NAND2_X1 U15745 ( .A1(n12611), .A2(n12610), .ZN(n12612) );
  NAND2_X2 U15746 ( .A1(n13218), .A2(n12612), .ZN(n13331) );
  NAND2_X1 U15747 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19057), .ZN(
        n12613) );
  AND2_X1 U15748 ( .A1(n12614), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12617) );
  NAND2_X1 U15749 ( .A1(n13768), .A2(n13777), .ZN(n12618) );
  NOR2_X1 U15750 ( .A1(n10072), .A2(n13536), .ZN(n13724) );
  AND2_X1 U15751 ( .A1(n13727), .A2(n13724), .ZN(n12619) );
  AOI22_X1 U15752 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12625) );
  AOI22_X1 U15753 ( .A1(n10527), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12624) );
  NAND2_X1 U15754 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12623) );
  NAND2_X1 U15755 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12622) );
  NAND4_X1 U15756 ( .A1(n12625), .A2(n12624), .A3(n12623), .A4(n12622), .ZN(
        n12636) );
  AOI22_X1 U15757 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12634) );
  AOI22_X1 U15758 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12633) );
  OAI22_X1 U15759 ( .A1(n10592), .A2(n12627), .B1(n12713), .B2(n12626), .ZN(
        n12630) );
  INV_X1 U15760 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n19250) );
  OAI22_X1 U15761 ( .A1(n12734), .A2(n19250), .B1(n12736), .B2(n12628), .ZN(
        n12629) );
  NOR2_X1 U15762 ( .A1(n12630), .A2(n12629), .ZN(n12632) );
  AOI22_X1 U15763 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12746), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12631) );
  NAND4_X1 U15764 ( .A1(n12634), .A2(n12633), .A3(n12632), .A4(n12631), .ZN(
        n12635) );
  OR2_X1 U15765 ( .A1(n12636), .A2(n12635), .ZN(n13927) );
  AOI22_X1 U15766 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12644) );
  AOI22_X1 U15767 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12643) );
  OAI22_X1 U15768 ( .A1(n12637), .A2(n10592), .B1(n12713), .B2(n12779), .ZN(
        n12640) );
  INV_X1 U15769 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13723) );
  OAI22_X1 U15770 ( .A1(n12734), .A2(n13723), .B1(n12638), .B2(n12736), .ZN(
        n12639) );
  NOR2_X1 U15771 ( .A1(n12640), .A2(n12639), .ZN(n12642) );
  AOI22_X1 U15772 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12746), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12641) );
  NAND4_X1 U15773 ( .A1(n12644), .A2(n12643), .A3(n12642), .A4(n12641), .ZN(
        n12650) );
  AOI22_X1 U15774 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12747), .B1(
        n12723), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12648) );
  AOI22_X1 U15775 ( .A1(n10527), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12647) );
  NAND2_X1 U15776 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12646) );
  NAND2_X1 U15777 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12645) );
  NAND4_X1 U15778 ( .A1(n12648), .A2(n12647), .A3(n12646), .A4(n12645), .ZN(
        n12649) );
  OR2_X1 U15779 ( .A1(n12650), .A2(n12649), .ZN(n13871) );
  NAND2_X1 U15780 ( .A1(n13868), .A2(n13871), .ZN(n13869) );
  AOI22_X1 U15781 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12659) );
  AOI22_X1 U15782 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12658) );
  OAI22_X1 U15783 ( .A1(n12651), .A2(n10592), .B1(n12713), .B2(n12806), .ZN(
        n12655) );
  INV_X1 U15784 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12653) );
  OAI22_X1 U15785 ( .A1(n12734), .A2(n12653), .B1(n12652), .B2(n12736), .ZN(
        n12654) );
  NOR2_X1 U15786 ( .A1(n12655), .A2(n12654), .ZN(n12657) );
  AOI22_X1 U15787 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n12746), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12656) );
  NAND4_X1 U15788 ( .A1(n12659), .A2(n12658), .A3(n12657), .A4(n12656), .ZN(
        n12665) );
  AOI22_X1 U15789 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12747), .B1(
        n12723), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U15790 ( .A1(n10527), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12662) );
  NAND2_X1 U15791 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n12661) );
  NAND2_X1 U15792 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12660) );
  NAND4_X1 U15793 ( .A1(n12663), .A2(n12662), .A3(n12661), .A4(n12660), .ZN(
        n12664) );
  NOR2_X1 U15794 ( .A1(n12665), .A2(n12664), .ZN(n13936) );
  INV_X1 U15795 ( .A(n13936), .ZN(n12666) );
  AOI22_X1 U15796 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12675) );
  AOI22_X1 U15797 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12674) );
  OAI22_X1 U15798 ( .A1(n10592), .A2(n12667), .B1(n12713), .B2(n12830), .ZN(
        n12671) );
  INV_X1 U15799 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12669) );
  OAI22_X1 U15800 ( .A1(n12734), .A2(n12669), .B1(n12736), .B2(n12668), .ZN(
        n12670) );
  NOR2_X1 U15801 ( .A1(n12671), .A2(n12670), .ZN(n12673) );
  AOI22_X1 U15802 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12746), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12672) );
  NAND4_X1 U15803 ( .A1(n12675), .A2(n12674), .A3(n12673), .A4(n12672), .ZN(
        n12681) );
  AOI22_X1 U15804 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12679) );
  AOI22_X1 U15805 ( .A1(n10527), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12678) );
  NAND2_X1 U15806 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12677) );
  NAND2_X1 U15807 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12676) );
  NAND4_X1 U15808 ( .A1(n12679), .A2(n12678), .A3(n12677), .A4(n12676), .ZN(
        n12680) );
  NOR2_X1 U15809 ( .A1(n12681), .A2(n12680), .ZN(n14859) );
  AOI22_X1 U15810 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12690) );
  AOI22_X1 U15811 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12689) );
  OAI22_X1 U15812 ( .A1(n10592), .A2(n12682), .B1(n12713), .B2(n12852), .ZN(
        n12686) );
  INV_X1 U15813 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12684) );
  OAI22_X1 U15814 ( .A1(n12734), .A2(n12684), .B1(n12736), .B2(n12683), .ZN(
        n12685) );
  NOR2_X1 U15815 ( .A1(n12686), .A2(n12685), .ZN(n12688) );
  AOI22_X1 U15816 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12746), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12687) );
  NAND4_X1 U15817 ( .A1(n12690), .A2(n12689), .A3(n12688), .A4(n12687), .ZN(
        n12696) );
  AOI22_X1 U15818 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12694) );
  AOI22_X1 U15819 ( .A1(n10527), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12693) );
  NAND2_X1 U15820 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12692) );
  NAND2_X1 U15821 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12691) );
  NAND4_X1 U15822 ( .A1(n12694), .A2(n12693), .A3(n12692), .A4(n12691), .ZN(
        n12695) );
  OR2_X1 U15823 ( .A1(n12696), .A2(n12695), .ZN(n14850) );
  AOI22_X1 U15824 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12706) );
  AOI22_X1 U15825 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12705) );
  OAI22_X1 U15826 ( .A1(n10592), .A2(n12698), .B1(n12713), .B2(n12875), .ZN(
        n12702) );
  INV_X1 U15827 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12700) );
  OAI22_X1 U15828 ( .A1(n12734), .A2(n12700), .B1(n12736), .B2(n12699), .ZN(
        n12701) );
  NOR2_X1 U15829 ( .A1(n12702), .A2(n12701), .ZN(n12704) );
  AOI22_X1 U15830 ( .A1(n10522), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12746), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12703) );
  NAND4_X1 U15831 ( .A1(n12706), .A2(n12705), .A3(n12704), .A4(n12703), .ZN(
        n12712) );
  AOI22_X1 U15832 ( .A1(n12723), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12747), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12710) );
  AOI22_X1 U15833 ( .A1(n10527), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12709) );
  NAND2_X1 U15834 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12708) );
  NAND2_X1 U15835 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12707) );
  NAND4_X1 U15836 ( .A1(n12710), .A2(n12709), .A3(n12708), .A4(n12707), .ZN(
        n12711) );
  OR2_X1 U15837 ( .A1(n12712), .A2(n12711), .ZN(n14847) );
  AOI22_X1 U15838 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12722) );
  AOI22_X1 U15839 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12721) );
  OAI22_X1 U15840 ( .A1(n12714), .A2(n10592), .B1(n12713), .B2(n12903), .ZN(
        n12718) );
  INV_X1 U15841 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12716) );
  OAI22_X1 U15842 ( .A1(n12734), .A2(n12716), .B1(n12715), .B2(n12736), .ZN(
        n12717) );
  NOR2_X1 U15843 ( .A1(n12718), .A2(n12717), .ZN(n12720) );
  AOI22_X1 U15844 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12746), .B1(
        n10522), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12719) );
  NAND4_X1 U15845 ( .A1(n12722), .A2(n12721), .A3(n12720), .A4(n12719), .ZN(
        n12731) );
  AOI22_X1 U15846 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12747), .B1(
        n12723), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U15847 ( .A1(n10527), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12724), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12728) );
  NAND2_X1 U15848 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12727) );
  NAND2_X1 U15849 ( .A1(n12432), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12726) );
  NAND4_X1 U15850 ( .A1(n12729), .A2(n12728), .A3(n12727), .A4(n12726), .ZN(
        n12730) );
  NOR2_X1 U15851 ( .A1(n12731), .A2(n12730), .ZN(n14842) );
  INV_X1 U15852 ( .A(n14842), .ZN(n12732) );
  AOI22_X1 U15853 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12432), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12745) );
  INV_X1 U15854 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12733) );
  OAI22_X1 U15855 ( .A1(n12925), .A2(n12735), .B1(n12734), .B2(n12733), .ZN(
        n12740) );
  OAI22_X1 U15856 ( .A1(n10592), .A2(n12738), .B1(n12737), .B2(n12736), .ZN(
        n12739) );
  NOR2_X1 U15857 ( .A1(n12740), .A2(n12739), .ZN(n12744) );
  AOI22_X1 U15858 ( .A1(n10457), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12697), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12743) );
  AOI22_X1 U15859 ( .A1(n12741), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10518), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12742) );
  NAND4_X1 U15860 ( .A1(n12745), .A2(n12744), .A3(n12743), .A4(n12742), .ZN(
        n12753) );
  AOI22_X1 U15861 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n10522), .B1(
        n12746), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U15862 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12747), .B1(
        n12723), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12750) );
  AOI22_X1 U15863 ( .A1(n10527), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12748), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12749) );
  NAND3_X1 U15864 ( .A1(n12751), .A2(n12750), .A3(n12749), .ZN(n12752) );
  NOR2_X1 U15865 ( .A1(n12753), .A2(n12752), .ZN(n12794) );
  AOI22_X1 U15866 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12764) );
  AOI22_X1 U15867 ( .A1(n10434), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10223), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12763) );
  AOI22_X1 U15868 ( .A1(n12892), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12762) );
  INV_X1 U15869 ( .A(n10226), .ZN(n12926) );
  INV_X1 U15870 ( .A(n12755), .ZN(n12757) );
  NAND2_X1 U15871 ( .A1(n19681), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12756) );
  NAND2_X1 U15872 ( .A1(n12757), .A2(n12756), .ZN(n12921) );
  NAND2_X1 U15873 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12758) );
  OAI211_X1 U15874 ( .C1(n12926), .C2(n12759), .A(n12921), .B(n12758), .ZN(
        n12760) );
  INV_X1 U15875 ( .A(n12760), .ZN(n12761) );
  NAND4_X1 U15876 ( .A1(n12764), .A2(n12763), .A3(n12762), .A4(n12761), .ZN(
        n12773) );
  AOI22_X1 U15877 ( .A1(n12915), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12771) );
  AOI22_X1 U15878 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12770) );
  AOI22_X1 U15879 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10223), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12769) );
  INV_X1 U15880 ( .A(n12892), .ZN(n16121) );
  INV_X1 U15881 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12766) );
  INV_X1 U15882 ( .A(n12921), .ZN(n12894) );
  NAND2_X1 U15883 ( .A1(n12901), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12765) );
  OAI211_X1 U15884 ( .C1(n16121), .C2(n12766), .A(n12894), .B(n12765), .ZN(
        n12767) );
  INV_X1 U15885 ( .A(n12767), .ZN(n12768) );
  NAND4_X1 U15886 ( .A1(n12771), .A2(n12770), .A3(n12769), .A4(n12768), .ZN(
        n12772) );
  NAND2_X1 U15887 ( .A1(n12773), .A2(n12772), .ZN(n12800) );
  NOR2_X1 U15888 ( .A1(n10264), .A2(n12800), .ZN(n12774) );
  XOR2_X1 U15889 ( .A(n12794), .B(n12774), .Z(n12801) );
  INV_X1 U15890 ( .A(n12800), .ZN(n12795) );
  NAND2_X1 U15891 ( .A1(n10264), .A2(n12795), .ZN(n14837) );
  AOI22_X1 U15892 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12784) );
  AOI22_X1 U15893 ( .A1(n12915), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12783) );
  AOI22_X1 U15894 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12782) );
  NAND2_X1 U15895 ( .A1(n10223), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12778) );
  OAI211_X1 U15896 ( .C1(n16121), .C2(n12779), .A(n12778), .B(n12921), .ZN(
        n12780) );
  INV_X1 U15897 ( .A(n12780), .ZN(n12781) );
  NAND4_X1 U15898 ( .A1(n12784), .A2(n12783), .A3(n12782), .A4(n12781), .ZN(
        n12793) );
  AOI22_X1 U15899 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12791) );
  AOI22_X1 U15900 ( .A1(n12915), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12790) );
  AOI22_X1 U15901 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12789) );
  NAND2_X1 U15902 ( .A1(n10223), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12785) );
  OAI211_X1 U15903 ( .C1(n16121), .C2(n12786), .A(n12785), .B(n12894), .ZN(
        n12787) );
  INV_X1 U15904 ( .A(n12787), .ZN(n12788) );
  NAND4_X1 U15905 ( .A1(n12791), .A2(n12790), .A3(n12789), .A4(n12788), .ZN(
        n12792) );
  NAND2_X1 U15906 ( .A1(n12793), .A2(n12792), .ZN(n12799) );
  INV_X1 U15907 ( .A(n12794), .ZN(n12796) );
  NAND2_X1 U15908 ( .A1(n12796), .A2(n12795), .ZN(n12802) );
  XOR2_X1 U15909 ( .A(n12799), .B(n12802), .Z(n12797) );
  NAND2_X1 U15910 ( .A1(n12797), .A2(n12869), .ZN(n14827) );
  NAND2_X1 U15911 ( .A1(n14824), .A2(n12798), .ZN(n14825) );
  INV_X1 U15912 ( .A(n12799), .ZN(n12803) );
  NAND2_X1 U15913 ( .A1(n10264), .A2(n12803), .ZN(n14830) );
  INV_X1 U15914 ( .A(n12802), .ZN(n12804) );
  AND2_X1 U15915 ( .A1(n12804), .A2(n12803), .ZN(n12822) );
  AOI22_X1 U15916 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12811) );
  AOI22_X1 U15917 ( .A1(n12915), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12810) );
  AOI22_X1 U15918 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12809) );
  NAND2_X1 U15919 ( .A1(n10223), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12805) );
  OAI211_X1 U15920 ( .C1(n16121), .C2(n12806), .A(n12805), .B(n12921), .ZN(
        n12807) );
  INV_X1 U15921 ( .A(n12807), .ZN(n12808) );
  NAND4_X1 U15922 ( .A1(n12811), .A2(n12810), .A3(n12809), .A4(n12808), .ZN(
        n12821) );
  AOI22_X1 U15923 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12819) );
  AOI22_X1 U15924 ( .A1(n12915), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12818) );
  AOI22_X1 U15925 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12817) );
  INV_X1 U15926 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12814) );
  NAND2_X1 U15927 ( .A1(n10223), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12813) );
  OAI211_X1 U15928 ( .C1(n16121), .C2(n12814), .A(n12813), .B(n12894), .ZN(
        n12815) );
  INV_X1 U15929 ( .A(n12815), .ZN(n12816) );
  NAND4_X1 U15930 ( .A1(n12819), .A2(n12818), .A3(n12817), .A4(n12816), .ZN(
        n12820) );
  AND2_X1 U15931 ( .A1(n12821), .A2(n12820), .ZN(n12823) );
  NAND2_X1 U15932 ( .A1(n12822), .A2(n12823), .ZN(n12848) );
  OAI211_X1 U15933 ( .C1(n12822), .C2(n12823), .A(n12869), .B(n12848), .ZN(
        n12826) );
  INV_X1 U15934 ( .A(n12823), .ZN(n12824) );
  NOR2_X1 U15935 ( .A1(n13720), .A2(n12824), .ZN(n14819) );
  NAND2_X1 U15936 ( .A1(n14818), .A2(n12828), .ZN(n12846) );
  AOI22_X1 U15937 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12835) );
  AOI22_X1 U15938 ( .A1(n12915), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12834) );
  AOI22_X1 U15939 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12833) );
  NAND2_X1 U15940 ( .A1(n10223), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12829) );
  OAI211_X1 U15941 ( .C1(n16121), .C2(n12830), .A(n12829), .B(n12921), .ZN(
        n12831) );
  INV_X1 U15942 ( .A(n12831), .ZN(n12832) );
  NAND4_X1 U15943 ( .A1(n12835), .A2(n12834), .A3(n12833), .A4(n12832), .ZN(
        n12844) );
  AOI22_X1 U15944 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12842) );
  AOI22_X1 U15945 ( .A1(n12915), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12841) );
  AOI22_X1 U15946 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12840) );
  INV_X1 U15947 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12837) );
  NAND2_X1 U15948 ( .A1(n10223), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12836) );
  OAI211_X1 U15949 ( .C1(n16121), .C2(n12837), .A(n12836), .B(n12894), .ZN(
        n12838) );
  INV_X1 U15950 ( .A(n12838), .ZN(n12839) );
  NAND4_X1 U15951 ( .A1(n12842), .A2(n12841), .A3(n12840), .A4(n12839), .ZN(
        n12843) );
  AND2_X1 U15952 ( .A1(n12844), .A2(n12843), .ZN(n12849) );
  XNOR2_X1 U15953 ( .A(n12848), .B(n12849), .ZN(n12845) );
  NAND2_X1 U15954 ( .A1(n10264), .A2(n12849), .ZN(n14814) );
  INV_X1 U15955 ( .A(n12848), .ZN(n12850) );
  NAND2_X1 U15956 ( .A1(n12850), .A2(n12849), .ZN(n12868) );
  INV_X1 U15957 ( .A(n12868), .ZN(n12870) );
  AOI22_X1 U15958 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12857) );
  AOI22_X1 U15959 ( .A1(n12915), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12856) );
  AOI22_X1 U15960 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12855) );
  NAND2_X1 U15961 ( .A1(n10223), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12851) );
  OAI211_X1 U15962 ( .C1(n16121), .C2(n12852), .A(n12851), .B(n12921), .ZN(
        n12853) );
  INV_X1 U15963 ( .A(n12853), .ZN(n12854) );
  NAND4_X1 U15964 ( .A1(n12857), .A2(n12856), .A3(n12855), .A4(n12854), .ZN(
        n12866) );
  AOI22_X1 U15965 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12864) );
  AOI22_X1 U15966 ( .A1(n12915), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12863) );
  AOI22_X1 U15967 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12862) );
  INV_X1 U15968 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12859) );
  NAND2_X1 U15969 ( .A1(n10223), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12858) );
  OAI211_X1 U15970 ( .C1(n16121), .C2(n12859), .A(n12858), .B(n12894), .ZN(
        n12860) );
  INV_X1 U15971 ( .A(n12860), .ZN(n12861) );
  NAND4_X1 U15972 ( .A1(n12864), .A2(n12863), .A3(n12862), .A4(n12861), .ZN(
        n12865) );
  NAND2_X1 U15973 ( .A1(n12866), .A2(n12865), .ZN(n12867) );
  INV_X1 U15974 ( .A(n12867), .ZN(n12873) );
  OR2_X1 U15975 ( .A1(n12868), .A2(n12867), .ZN(n14797) );
  OAI211_X1 U15976 ( .C1(n12870), .C2(n12873), .A(n14797), .B(n12869), .ZN(
        n12871) );
  INV_X1 U15977 ( .A(n12890), .ZN(n14798) );
  NAND2_X1 U15978 ( .A1(n14798), .A2(n12872), .ZN(n14805) );
  NAND2_X1 U15979 ( .A1(n10264), .A2(n12873), .ZN(n14804) );
  AOI22_X1 U15980 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12880) );
  AOI22_X1 U15981 ( .A1(n12915), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12879) );
  AOI22_X1 U15982 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12878) );
  NAND2_X1 U15983 ( .A1(n10223), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12874) );
  OAI211_X1 U15984 ( .C1(n16121), .C2(n12875), .A(n12874), .B(n12921), .ZN(
        n12876) );
  INV_X1 U15985 ( .A(n12876), .ZN(n12877) );
  NAND4_X1 U15986 ( .A1(n12880), .A2(n12879), .A3(n12878), .A4(n12877), .ZN(
        n12889) );
  AOI22_X1 U15987 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12887) );
  AOI22_X1 U15988 ( .A1(n12915), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12886) );
  AOI22_X1 U15989 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12885) );
  NAND2_X1 U15990 ( .A1(n10223), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12881) );
  OAI211_X1 U15991 ( .C1(n16121), .C2(n12882), .A(n12881), .B(n12894), .ZN(
        n12883) );
  INV_X1 U15992 ( .A(n12883), .ZN(n12884) );
  NAND4_X1 U15993 ( .A1(n12887), .A2(n12886), .A3(n12885), .A4(n12884), .ZN(
        n12888) );
  AND2_X1 U15994 ( .A1(n12889), .A2(n12888), .ZN(n14799) );
  OAI21_X1 U15995 ( .B1(n14803), .B2(n12890), .A(n14799), .ZN(n14029) );
  NAND2_X1 U15996 ( .A1(n13720), .A2(n14799), .ZN(n12891) );
  NOR2_X1 U15997 ( .A1(n14797), .A2(n12891), .ZN(n12912) );
  AOI22_X1 U15998 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12900) );
  AOI22_X1 U15999 ( .A1(n10434), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10223), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12899) );
  AOI22_X1 U16000 ( .A1(n12892), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12898) );
  OAI211_X1 U16001 ( .C1(n12926), .C2(n12895), .A(n12894), .B(n12893), .ZN(
        n12896) );
  INV_X1 U16002 ( .A(n12896), .ZN(n12897) );
  NAND4_X1 U16003 ( .A1(n12900), .A2(n12899), .A3(n12898), .A4(n12897), .ZN(
        n12910) );
  AOI22_X1 U16004 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12908) );
  AOI22_X1 U16005 ( .A1(n12915), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12907) );
  AOI22_X1 U16006 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12906) );
  NAND2_X1 U16007 ( .A1(n10223), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12902) );
  OAI211_X1 U16008 ( .C1(n16121), .C2(n12903), .A(n12902), .B(n12921), .ZN(
        n12904) );
  INV_X1 U16009 ( .A(n12904), .ZN(n12905) );
  NAND4_X1 U16010 ( .A1(n12908), .A2(n12907), .A3(n12906), .A4(n12905), .ZN(
        n12909) );
  AND2_X1 U16011 ( .A1(n12910), .A2(n12909), .ZN(n12911) );
  NAND2_X1 U16012 ( .A1(n12912), .A2(n12911), .ZN(n12913) );
  OAI21_X1 U16013 ( .B1(n12912), .B2(n12911), .A(n12913), .ZN(n14028) );
  NOR2_X1 U16014 ( .A1(n14029), .A2(n14028), .ZN(n14027) );
  INV_X1 U16015 ( .A(n12913), .ZN(n12914) );
  NOR2_X1 U16016 ( .A1(n14027), .A2(n12914), .ZN(n12937) );
  AOI22_X1 U16017 ( .A1(n12915), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12917) );
  AOI22_X1 U16018 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10223), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12916) );
  NAND2_X1 U16019 ( .A1(n12917), .A2(n12916), .ZN(n12935) );
  INV_X1 U16020 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12920) );
  AOI22_X1 U16021 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12919) );
  AOI21_X1 U16022 ( .B1(n12901), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n12921), .ZN(n12918) );
  OAI211_X1 U16023 ( .C1(n16121), .C2(n12920), .A(n12919), .B(n12918), .ZN(
        n12934) );
  OAI21_X1 U16024 ( .B1(n12923), .B2(n12922), .A(n12921), .ZN(n12928) );
  OAI22_X1 U16025 ( .A1(n12926), .A2(n12925), .B1(n16121), .B2(n12924), .ZN(
        n12927) );
  AOI211_X1 U16026 ( .C1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .C2(n10442), .A(
        n12928), .B(n12927), .ZN(n12932) );
  AOI22_X1 U16027 ( .A1(n10434), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12901), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12931) );
  AOI22_X1 U16028 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12929), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12930) );
  NAND3_X1 U16029 ( .A1(n12932), .A2(n12931), .A3(n12930), .ZN(n12933) );
  OAI21_X1 U16030 ( .B1(n12935), .B2(n12934), .A(n12933), .ZN(n12936) );
  XNOR2_X1 U16031 ( .A(n12937), .B(n12936), .ZN(n14126) );
  NAND2_X1 U16032 ( .A1(n12540), .A2(n19740), .ZN(n16140) );
  OAI22_X1 U16033 ( .A1(n16138), .A2(n15434), .B1(n16142), .B2(n16140), .ZN(
        n13128) );
  AND2_X1 U16034 ( .A1(n12939), .A2(n12938), .ZN(n12940) );
  NAND2_X1 U16035 ( .A1(n18953), .A2(n12943), .ZN(n18954) );
  AOI22_X1 U16036 ( .A1(n15085), .A2(n18964), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n18963), .ZN(n12959) );
  NAND2_X1 U16037 ( .A1(n18953), .A2(n10233), .ZN(n13210) );
  NOR4_X1 U16038 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12947) );
  NOR4_X1 U16039 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12946) );
  NOR4_X1 U16040 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12945) );
  NOR4_X1 U16041 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12944) );
  NAND4_X1 U16042 ( .A1(n12947), .A2(n12946), .A3(n12945), .A4(n12944), .ZN(
        n12952) );
  NOR4_X1 U16043 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_27__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n12950) );
  NOR4_X1 U16044 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12949) );
  NOR4_X1 U16045 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12948) );
  INV_X1 U16046 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19627) );
  NAND4_X1 U16047 ( .A1(n12950), .A2(n12949), .A3(n12948), .A4(n19627), .ZN(
        n12951) );
  NOR2_X2 U16048 ( .A1(n13210), .A2(n13717), .ZN(n18910) );
  NOR2_X2 U16049 ( .A1(n13210), .A2(n13715), .ZN(n18911) );
  AOI22_X1 U16050 ( .A1(n18910), .A2(BUF2_REG_30__SCAN_IN), .B1(n18911), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n12953) );
  INV_X1 U16051 ( .A(n12953), .ZN(n12957) );
  AND2_X1 U16052 ( .A1(n10768), .A2(n10271), .ZN(n12954) );
  INV_X1 U16053 ( .A(n14930), .ZN(n18909) );
  NAND2_X1 U16054 ( .A1(n13052), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12956) );
  INV_X1 U16055 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14330) );
  OR2_X1 U16056 ( .A1(n13715), .A2(n14330), .ZN(n12955) );
  NAND2_X1 U16057 ( .A1(n12956), .A2(n12955), .ZN(n18921) );
  NOR2_X1 U16058 ( .A1(n12957), .A2(n10086), .ZN(n12958) );
  OAI21_X1 U16059 ( .B1(n14126), .B2(n18968), .A(n12960), .ZN(P2_U2889) );
  NOR2_X1 U16060 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12962) );
  NOR4_X1 U16061 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12961) );
  NAND4_X1 U16062 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12962), .A4(n12961), .ZN(n12965) );
  NOR2_X1 U16063 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12965), .ZN(n16299)
         );
  INV_X1 U16064 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20674) );
  NOR3_X1 U16065 ( .A1(P1_BE_N_REG_3__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20674), .ZN(n12964) );
  NOR4_X1 U16066 ( .A1(P1_BE_N_REG_1__SCAN_IN), .A2(P1_BE_N_REG_2__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12963) );
  NAND4_X1 U16067 ( .A1(n20001), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12964), .A4(
        n12963), .ZN(U214) );
  NOR2_X1 U16068 ( .A1(n13715), .A2(n12965), .ZN(n16226) );
  NAND2_X1 U16069 ( .A1(n16226), .A2(U214), .ZN(U212) );
  NAND2_X1 U16070 ( .A1(n12966), .A2(n15266), .ZN(n15246) );
  OR2_X1 U16071 ( .A1(n14999), .A2(n12967), .ZN(n15245) );
  NOR2_X1 U16072 ( .A1(n15246), .A2(n15245), .ZN(n15248) );
  NOR2_X1 U16073 ( .A1(n15248), .A2(n14999), .ZN(n12970) );
  NOR2_X1 U16074 ( .A1(n15002), .A2(n12968), .ZN(n12969) );
  XNOR2_X1 U16075 ( .A(n12970), .B(n12969), .ZN(n16014) );
  NOR2_X1 U16076 ( .A1(n16014), .A2(n15405), .ZN(n12992) );
  NAND2_X1 U16077 ( .A1(n12971), .A2(n12972), .ZN(n15243) );
  XNOR2_X1 U16078 ( .A(n15243), .B(n12973), .ZN(n16013) );
  NOR2_X1 U16079 ( .A1(n16013), .A2(n15413), .ZN(n12991) );
  INV_X1 U16080 ( .A(n12974), .ZN(n12977) );
  NAND2_X1 U16081 ( .A1(n15316), .A2(n12977), .ZN(n12975) );
  INV_X1 U16082 ( .A(n15315), .ZN(n16078) );
  NAND2_X1 U16083 ( .A1(n12975), .A2(n16078), .ZN(n15296) );
  NAND2_X1 U16084 ( .A1(n15366), .A2(n12978), .ZN(n12976) );
  NAND2_X1 U16085 ( .A1(n15296), .A2(n12976), .ZN(n15215) );
  AND2_X1 U16086 ( .A1(n15215), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12990) );
  AND2_X1 U16087 ( .A1(n15349), .A2(n12977), .ZN(n15275) );
  INV_X1 U16088 ( .A(n12978), .ZN(n12979) );
  NAND2_X1 U16089 ( .A1(n15275), .A2(n12979), .ZN(n15219) );
  NOR2_X1 U16090 ( .A1(n12981), .A2(n12980), .ZN(n12982) );
  OR2_X1 U16091 ( .A1(n15232), .A2(n12982), .ZN(n18920) );
  INV_X1 U16092 ( .A(n18920), .ZN(n12984) );
  NOR2_X1 U16093 ( .A1(n10456), .A2(n18847), .ZN(n12983) );
  AOI21_X1 U16094 ( .B1(n15410), .B2(n12984), .A(n12983), .ZN(n12988) );
  NAND2_X1 U16095 ( .A1(n13699), .A2(n12985), .ZN(n12986) );
  AND2_X1 U16096 ( .A1(n9728), .A2(n12986), .ZN(n18733) );
  NAND2_X1 U16097 ( .A1(n16104), .A2(n18733), .ZN(n12987) );
  OAI211_X1 U16098 ( .C1(n15219), .C2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n12988), .B(n12987), .ZN(n12989) );
  OR4_X1 U16099 ( .A1(n12992), .A2(n12991), .A3(n12990), .A4(n12989), .ZN(
        P2_U3031) );
  AOI211_X1 U16100 ( .C1(n14993), .C2(n12994), .A(n12993), .B(n19606), .ZN(
        n13004) );
  OAI22_X1 U16101 ( .A1(n14990), .A2(n18874), .B1(n10377), .B2(n18849), .ZN(
        n13003) );
  INV_X1 U16102 ( .A(n12995), .ZN(n12996) );
  OAI22_X1 U16103 ( .A1(n12996), .A2(n18888), .B1(n10787), .B2(n18857), .ZN(
        n13002) );
  NAND2_X1 U16104 ( .A1(n14749), .A2(n12997), .ZN(n12998) );
  NAND2_X1 U16105 ( .A1(n14832), .A2(n12998), .ZN(n15146) );
  OR2_X1 U16106 ( .A1(n14754), .A2(n12999), .ZN(n13000) );
  NAND2_X1 U16107 ( .A1(n14907), .A2(n13000), .ZN(n15150) );
  OAI22_X1 U16108 ( .A1(n15146), .A2(n18871), .B1(n15150), .B2(n18893), .ZN(
        n13001) );
  OR4_X1 U16109 ( .A1(n13004), .A2(n13003), .A3(n13002), .A4(n13001), .ZN(
        P2_U2832) );
  AOI211_X1 U16110 ( .C1(n14951), .C2(n13006), .A(n13005), .B(n19606), .ZN(
        n13017) );
  OAI22_X1 U16111 ( .A1(n14949), .A2(n18874), .B1(n19658), .B2(n18849), .ZN(
        n13016) );
  OAI22_X1 U16112 ( .A1(n13007), .A2(n18888), .B1(n18857), .B2(n10393), .ZN(
        n13015) );
  INV_X1 U16113 ( .A(n13008), .ZN(n13011) );
  NAND2_X1 U16114 ( .A1(n14812), .A2(n13009), .ZN(n13010) );
  NAND2_X1 U16115 ( .A1(n13011), .A2(n13010), .ZN(n15108) );
  INV_X1 U16116 ( .A(n13012), .ZN(n14890) );
  OAI22_X1 U16117 ( .A1(n15108), .A2(n18871), .B1(n14881), .B2(n18893), .ZN(
        n13014) );
  OR4_X1 U16118 ( .A1(n13017), .A2(n13016), .A3(n13015), .A4(n13014), .ZN(
        P2_U2828) );
  OAI21_X1 U16119 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13019), .A(
        n13018), .ZN(n13140) );
  NAND2_X1 U16120 ( .A1(n19011), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13141) );
  OAI21_X1 U16121 ( .B1(n13140), .B2(n15405), .A(n13141), .ZN(n13029) );
  AOI211_X1 U16122 ( .C1(n13025), .C2(n13020), .A(n13290), .B(n15367), .ZN(
        n13028) );
  OAI21_X1 U16123 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13022), .A(
        n13021), .ZN(n13142) );
  INV_X1 U16124 ( .A(n18872), .ZN(n13143) );
  OAI22_X1 U16125 ( .A1(n15413), .A2(n13142), .B1(n13143), .B2(n15404), .ZN(
        n13027) );
  XNOR2_X1 U16126 ( .A(n13024), .B(n13023), .ZN(n19708) );
  INV_X1 U16127 ( .A(n19708), .ZN(n13317) );
  OAI22_X1 U16128 ( .A1(n13288), .A2(n13025), .B1(n16097), .B2(n13317), .ZN(
        n13026) );
  OR4_X1 U16129 ( .A1(n13029), .A2(n13028), .A3(n13027), .A4(n13026), .ZN(
        P2_U3045) );
  NOR2_X1 U16130 ( .A1(n10760), .A2(n13030), .ZN(n18897) );
  INV_X1 U16131 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13033) );
  INV_X1 U16132 ( .A(n13031), .ZN(n13032) );
  NAND2_X1 U16133 ( .A1(n19688), .A2(n19601), .ZN(n13035) );
  OAI211_X1 U16134 ( .C1(n18897), .C2(n13033), .A(n13032), .B(n13035), .ZN(
        P2_U2814) );
  INV_X1 U16135 ( .A(n19735), .ZN(n18653) );
  NOR2_X1 U16136 ( .A1(n18653), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n13036)
         );
  AOI22_X1 U16137 ( .A1(n13036), .A2(n13035), .B1(n13034), .B2(n18653), .ZN(
        P2_U3612) );
  INV_X1 U16138 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13038) );
  NAND2_X1 U16139 ( .A1(n13108), .A2(n13037), .ZN(n13046) );
  INV_X1 U16140 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13155) );
  OAI22_X1 U16141 ( .A1(n13715), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13717), .ZN(n19033) );
  OAI222_X1 U16142 ( .A1(n13038), .A2(n13046), .B1(n13108), .B2(n13155), .C1(
        n13043), .C2(n19033), .ZN(P2_U2952) );
  INV_X1 U16143 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n13040) );
  OAI222_X1 U16144 ( .A1(n13040), .A2(n13046), .B1(n13043), .B2(n19033), .C1(
        n13108), .C2(n13039), .ZN(P2_U2967) );
  INV_X1 U16145 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13042) );
  AOI22_X1 U16146 ( .A1(n13717), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13715), .ZN(n18919) );
  INV_X1 U16147 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13041) );
  OAI222_X1 U16148 ( .A1(n13042), .A2(n13046), .B1(n13043), .B2(n18919), .C1(
        n13041), .C2(n13108), .ZN(P2_U2982) );
  INV_X1 U16149 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n18985) );
  INV_X1 U16150 ( .A(n13043), .ZN(n13092) );
  NAND2_X1 U16151 ( .A1(n13052), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13045) );
  INV_X1 U16152 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16254) );
  OR2_X1 U16153 ( .A1(n13715), .A2(n16254), .ZN(n13044) );
  NAND2_X1 U16154 ( .A1(n13045), .A2(n13044), .ZN(n18926) );
  NAND2_X1 U16155 ( .A1(n13092), .A2(n18926), .ZN(n13057) );
  INV_X2 U16156 ( .A(n13046), .ZN(n13105) );
  NAND2_X1 U16157 ( .A1(n13105), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13047) );
  OAI211_X1 U16158 ( .C1(n18985), .C2(n13108), .A(n13057), .B(n13047), .ZN(
        P2_U2979) );
  INV_X1 U16159 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n18981) );
  NAND2_X1 U16160 ( .A1(n13092), .A2(n18921), .ZN(n13059) );
  NAND2_X1 U16161 ( .A1(n13105), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13048) );
  OAI211_X1 U16162 ( .C1(n18981), .C2(n13108), .A(n13059), .B(n13048), .ZN(
        P2_U2981) );
  INV_X1 U16163 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13169) );
  NAND2_X1 U16164 ( .A1(n13052), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13050) );
  INV_X1 U16165 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16260) );
  OR2_X1 U16166 ( .A1(n13715), .A2(n16260), .ZN(n13049) );
  NAND2_X1 U16167 ( .A1(n13050), .A2(n13049), .ZN(n18938) );
  NAND2_X1 U16168 ( .A1(n13092), .A2(n18938), .ZN(n13063) );
  NAND2_X1 U16169 ( .A1(n13105), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13051) );
  OAI211_X1 U16170 ( .C1(n13169), .C2(n13108), .A(n13063), .B(n13051), .ZN(
        P2_U2960) );
  INV_X1 U16171 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13159) );
  NAND2_X1 U16172 ( .A1(n13052), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13054) );
  INV_X1 U16173 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16257) );
  OR2_X1 U16174 ( .A1(n13715), .A2(n16257), .ZN(n13053) );
  NAND2_X1 U16175 ( .A1(n13054), .A2(n13053), .ZN(n18931) );
  NAND2_X1 U16176 ( .A1(n13092), .A2(n18931), .ZN(n13061) );
  NAND2_X1 U16177 ( .A1(n13105), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13055) );
  OAI211_X1 U16178 ( .C1(n13159), .C2(n13108), .A(n13061), .B(n13055), .ZN(
        P2_U2962) );
  INV_X1 U16179 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13171) );
  NAND2_X1 U16180 ( .A1(n13105), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13056) );
  OAI211_X1 U16181 ( .C1(n13171), .C2(n13108), .A(n13057), .B(n13056), .ZN(
        P2_U2964) );
  INV_X1 U16182 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13173) );
  NAND2_X1 U16183 ( .A1(n13105), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13058) );
  OAI211_X1 U16184 ( .C1(n13173), .C2(n13108), .A(n13059), .B(n13058), .ZN(
        P2_U2966) );
  INV_X1 U16185 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n18989) );
  NAND2_X1 U16186 ( .A1(n13105), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13060) );
  OAI211_X1 U16187 ( .C1(n18989), .C2(n13108), .A(n13061), .B(n13060), .ZN(
        P2_U2977) );
  INV_X1 U16188 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n18993) );
  NAND2_X1 U16189 ( .A1(n13105), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13062) );
  OAI211_X1 U16190 ( .C1(n18993), .C2(n13108), .A(n13063), .B(n13062), .ZN(
        P2_U2975) );
  AOI22_X1 U16191 ( .A1(n13105), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n13104), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13065) );
  AOI22_X1 U16192 ( .A1(n13717), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13715), .ZN(n18973) );
  INV_X1 U16193 ( .A(n18973), .ZN(n13064) );
  NAND2_X1 U16194 ( .A1(n13092), .A2(n13064), .ZN(n13074) );
  NAND2_X1 U16195 ( .A1(n13065), .A2(n13074), .ZN(P2_U2953) );
  AOI22_X1 U16196 ( .A1(n13105), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n13104), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13066) );
  OAI22_X1 U16197 ( .A1(n13715), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13717), .ZN(n19042) );
  INV_X1 U16198 ( .A(n19042), .ZN(n15990) );
  NAND2_X1 U16199 ( .A1(n13092), .A2(n15990), .ZN(n13098) );
  NAND2_X1 U16200 ( .A1(n13066), .A2(n13098), .ZN(P2_U2969) );
  AOI22_X1 U16201 ( .A1(n13105), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n13104), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n13068) );
  AOI22_X1 U16202 ( .A1(n13717), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13715), .ZN(n19046) );
  INV_X1 U16203 ( .A(n19046), .ZN(n13067) );
  NAND2_X1 U16204 ( .A1(n13092), .A2(n13067), .ZN(n13080) );
  NAND2_X1 U16205 ( .A1(n13068), .A2(n13080), .ZN(P2_U2970) );
  AOI22_X1 U16206 ( .A1(n13105), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n13104), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13069) );
  OAI22_X1 U16207 ( .A1(n13715), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13717), .ZN(n19050) );
  INV_X1 U16208 ( .A(n19050), .ZN(n15982) );
  NAND2_X1 U16209 ( .A1(n13092), .A2(n15982), .ZN(n13094) );
  NAND2_X1 U16210 ( .A1(n13069), .A2(n13094), .ZN(P2_U2971) );
  AOI22_X1 U16211 ( .A1(n13105), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n13104), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13071) );
  AOI22_X1 U16212 ( .A1(n13717), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13715), .ZN(n19053) );
  INV_X1 U16213 ( .A(n19053), .ZN(n13070) );
  NAND2_X1 U16214 ( .A1(n13092), .A2(n13070), .ZN(n13076) );
  NAND2_X1 U16215 ( .A1(n13071), .A2(n13076), .ZN(P2_U2972) );
  AOI22_X1 U16216 ( .A1(n13105), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n13104), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13073) );
  AOI22_X1 U16217 ( .A1(n13717), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13715), .ZN(n19069) );
  INV_X1 U16218 ( .A(n19069), .ZN(n13072) );
  NAND2_X1 U16219 ( .A1(n13092), .A2(n13072), .ZN(n13078) );
  NAND2_X1 U16220 ( .A1(n13073), .A2(n13078), .ZN(P2_U2974) );
  AOI22_X1 U16221 ( .A1(n13105), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n13104), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13075) );
  NAND2_X1 U16222 ( .A1(n13075), .A2(n13074), .ZN(P2_U2968) );
  AOI22_X1 U16223 ( .A1(n13105), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n13104), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13077) );
  NAND2_X1 U16224 ( .A1(n13077), .A2(n13076), .ZN(P2_U2957) );
  AOI22_X1 U16225 ( .A1(n13105), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n13104), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13079) );
  NAND2_X1 U16226 ( .A1(n13079), .A2(n13078), .ZN(P2_U2959) );
  AOI22_X1 U16227 ( .A1(n13105), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n13104), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13081) );
  NAND2_X1 U16228 ( .A1(n13081), .A2(n13080), .ZN(P2_U2955) );
  AOI22_X1 U16229 ( .A1(n13105), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n13104), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13082) );
  OAI22_X1 U16230 ( .A1(n13715), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13717), .ZN(n19058) );
  INV_X1 U16231 ( .A(n19058), .ZN(n15976) );
  NAND2_X1 U16232 ( .A1(n13092), .A2(n15976), .ZN(n13106) );
  NAND2_X1 U16233 ( .A1(n13082), .A2(n13106), .ZN(P2_U2973) );
  AOI22_X1 U16234 ( .A1(n13105), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n13104), .ZN(n13085) );
  INV_X1 U16235 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n14350) );
  NOR2_X1 U16236 ( .A1(n13715), .A2(n14350), .ZN(n13083) );
  AOI21_X1 U16237 ( .B1(n13715), .B2(BUF2_REG_11__SCAN_IN), .A(n13083), .ZN(
        n18929) );
  INV_X1 U16238 ( .A(n18929), .ZN(n13084) );
  NAND2_X1 U16239 ( .A1(n13092), .A2(n13084), .ZN(n13096) );
  NAND2_X1 U16240 ( .A1(n13085), .A2(n13096), .ZN(P2_U2963) );
  AOI22_X1 U16241 ( .A1(n13105), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n13104), .ZN(n13088) );
  INV_X1 U16242 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13911) );
  NOR2_X1 U16243 ( .A1(n13715), .A2(n13911), .ZN(n13086) );
  AOI21_X1 U16244 ( .B1(n13715), .B2(BUF2_REG_9__SCAN_IN), .A(n13086), .ZN(
        n18934) );
  INV_X1 U16245 ( .A(n18934), .ZN(n13087) );
  NAND2_X1 U16246 ( .A1(n13092), .A2(n13087), .ZN(n13100) );
  NAND2_X1 U16247 ( .A1(n13088), .A2(n13100), .ZN(P2_U2961) );
  AOI22_X1 U16248 ( .A1(n13105), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n13104), .ZN(n13093) );
  INV_X1 U16249 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n13089) );
  NOR2_X1 U16250 ( .A1(n13717), .A2(n13089), .ZN(n13090) );
  AOI21_X1 U16251 ( .B1(BUF1_REG_13__SCAN_IN), .B2(n13717), .A(n13090), .ZN(
        n18924) );
  INV_X1 U16252 ( .A(n18924), .ZN(n13091) );
  NAND2_X1 U16253 ( .A1(n13092), .A2(n13091), .ZN(n13102) );
  NAND2_X1 U16254 ( .A1(n13093), .A2(n13102), .ZN(P2_U2980) );
  AOI22_X1 U16255 ( .A1(n13105), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n13104), .ZN(n13095) );
  NAND2_X1 U16256 ( .A1(n13095), .A2(n13094), .ZN(P2_U2956) );
  AOI22_X1 U16257 ( .A1(n13105), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n13104), .ZN(n13097) );
  NAND2_X1 U16258 ( .A1(n13097), .A2(n13096), .ZN(P2_U2978) );
  AOI22_X1 U16259 ( .A1(n13105), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n13104), .ZN(n13099) );
  NAND2_X1 U16260 ( .A1(n13099), .A2(n13098), .ZN(P2_U2954) );
  AOI22_X1 U16261 ( .A1(n13105), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n13104), .ZN(n13101) );
  NAND2_X1 U16262 ( .A1(n13101), .A2(n13100), .ZN(P2_U2976) );
  AOI22_X1 U16263 ( .A1(n13105), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n13104), .ZN(n13103) );
  NAND2_X1 U16264 ( .A1(n13103), .A2(n13102), .ZN(P2_U2965) );
  AOI22_X1 U16265 ( .A1(n13105), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n13104), .ZN(n13107) );
  NAND2_X1 U16266 ( .A1(n13107), .A2(n13106), .ZN(P2_U2958) );
  INV_X1 U16267 ( .A(n10760), .ZN(n13130) );
  NAND3_X1 U16268 ( .A1(n13131), .A2(n13130), .A3(n19598), .ZN(n13109) );
  NAND2_X1 U16269 ( .A1(n13109), .A2(n13108), .ZN(n13110) );
  NAND2_X1 U16270 ( .A1(n18990), .A2(n13111), .ZN(n18975) );
  INV_X1 U16271 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13874) );
  NAND2_X1 U16272 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n19713) );
  NOR2_X1 U16273 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19713), .ZN(n13167) );
  INV_X1 U16274 ( .A(n13167), .ZN(n19737) );
  INV_X1 U16275 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n16246) );
  INV_X1 U16276 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n20775) );
  OAI222_X1 U16277 ( .A1(n18975), .A2(n13874), .B1(n18978), .B2(n16246), .C1(
        n19737), .C2(n20775), .ZN(P2_U2934) );
  XNOR2_X1 U16278 ( .A(n18887), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13242) );
  NAND2_X1 U16279 ( .A1(n19011), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13237) );
  INV_X1 U16280 ( .A(n13237), .ZN(n13114) );
  XNOR2_X1 U16281 ( .A(n13112), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13239) );
  NOR2_X1 U16282 ( .A1(n16073), .A2(n13239), .ZN(n13113) );
  AOI211_X1 U16283 ( .C1(n13242), .C2(n19013), .A(n13114), .B(n13113), .ZN(
        n13117) );
  OAI21_X1 U16284 ( .B1(n19012), .B2(n13115), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13116) );
  OAI211_X1 U16285 ( .C1(n19020), .C2(n13238), .A(n13117), .B(n13116), .ZN(
        P2_U3014) );
  NAND2_X1 U16286 ( .A1(n13179), .A2(n13451), .ZN(n13587) );
  INV_X1 U16287 ( .A(n13245), .ZN(n13180) );
  NAND2_X1 U16288 ( .A1(n20657), .A2(n20577), .ZN(n19759) );
  NAND2_X1 U16289 ( .A1(n20678), .A2(n19759), .ZN(n13174) );
  AOI21_X1 U16290 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(n13587), .A(n13174), 
        .ZN(n13118) );
  INV_X1 U16291 ( .A(n13118), .ZN(P1_U2801) );
  NAND2_X1 U16292 ( .A1(n13720), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13119) );
  AND4_X1 U16293 ( .A1(n13119), .A2(n10268), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19732), .ZN(n13120) );
  NAND2_X1 U16294 ( .A1(n16138), .A2(n16130), .ZN(n13126) );
  NAND2_X1 U16295 ( .A1(n13126), .A2(n15438), .ZN(n13121) );
  NAND2_X1 U16296 ( .A1(n14796), .A2(n10271), .ZN(n14854) );
  MUX2_X1 U16297 ( .A(n13238), .B(n13123), .S(n14861), .Z(n13124) );
  OAI21_X1 U16298 ( .B1(n19716), .B2(n14854), .A(n13124), .ZN(P2_U2887) );
  NAND2_X1 U16299 ( .A1(n13126), .A2(n13125), .ZN(n13127) );
  NOR2_X1 U16300 ( .A1(n13128), .A2(n13127), .ZN(n13133) );
  NAND3_X1 U16301 ( .A1(n13131), .A2(n13130), .A3(n13129), .ZN(n13132) );
  NOR2_X1 U16302 ( .A1(n19741), .A2(n19713), .ZN(n16182) );
  AOI22_X1 U16303 ( .A1(n19741), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n16182), 
        .B2(P2_FLUSH_REG_SCAN_IN), .ZN(n13134) );
  OAI21_X1 U16304 ( .B1(n16129), .B2(n18657), .A(n13134), .ZN(n19679) );
  INV_X1 U16305 ( .A(n19679), .ZN(n15431) );
  NAND2_X1 U16306 ( .A1(n13137), .A2(n13136), .ZN(n16160) );
  OR4_X1 U16307 ( .A1(n15431), .A2(n19685), .A3(n13135), .A4(n16160), .ZN(
        n13138) );
  OAI21_X1 U16308 ( .B1(n13139), .B2(n19679), .A(n13138), .ZN(P2_U3595) );
  INV_X1 U16309 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18873) );
  OAI22_X1 U16310 ( .A1(n13140), .A2(n16072), .B1(n18873), .B2(n16059), .ZN(
        n13146) );
  OAI21_X1 U16311 ( .B1(n16073), .B2(n13142), .A(n13141), .ZN(n13145) );
  OAI22_X1 U16312 ( .A1(n13143), .A2(n19020), .B1(n19025), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13144) );
  OR3_X1 U16313 ( .A1(n13146), .A2(n13145), .A3(n13144), .ZN(P2_U3013) );
  INV_X1 U16314 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14870) );
  AOI22_X1 U16315 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n19007), .B1(n19008), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13147) );
  OAI21_X1 U16316 ( .B1(n14870), .B2(n18975), .A(n13147), .ZN(P2_U2922) );
  NOR2_X1 U16317 ( .A1(n14796), .A2(n20734), .ZN(n13152) );
  AOI21_X1 U16318 ( .B1(n18872), .B2(n14796), .A(n13152), .ZN(n13153) );
  OAI21_X1 U16319 ( .B1(n19026), .B2(n14854), .A(n13153), .ZN(P2_U2886) );
  AOI22_X1 U16320 ( .A1(n13167), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13154) );
  OAI21_X1 U16321 ( .B1(n13155), .B2(n18975), .A(n13154), .ZN(P2_U2935) );
  INV_X1 U16322 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14929) );
  AOI22_X1 U16323 ( .A1(n13167), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13156) );
  OAI21_X1 U16324 ( .B1(n14929), .B2(n18975), .A(n13156), .ZN(P2_U2932) );
  INV_X1 U16325 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n14914) );
  AOI22_X1 U16326 ( .A1(n13167), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13157) );
  OAI21_X1 U16327 ( .B1(n14914), .B2(n18975), .A(n13157), .ZN(P2_U2928) );
  AOI22_X1 U16328 ( .A1(n13167), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13158) );
  OAI21_X1 U16329 ( .B1(n13159), .B2(n18975), .A(n13158), .ZN(P2_U2925) );
  INV_X1 U16330 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13161) );
  AOI22_X1 U16331 ( .A1(n13167), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13160) );
  OAI21_X1 U16332 ( .B1(n13161), .B2(n18975), .A(n13160), .ZN(P2_U2931) );
  INV_X1 U16333 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14920) );
  AOI22_X1 U16334 ( .A1(n13167), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13162) );
  OAI21_X1 U16335 ( .B1(n14920), .B2(n18975), .A(n13162), .ZN(P2_U2930) );
  INV_X1 U16336 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13164) );
  AOI22_X1 U16337 ( .A1(n13167), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13163) );
  OAI21_X1 U16338 ( .B1(n13164), .B2(n18975), .A(n13163), .ZN(P2_U2929) );
  INV_X1 U16339 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14900) );
  AOI22_X1 U16340 ( .A1(n13167), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13165) );
  OAI21_X1 U16341 ( .B1(n14900), .B2(n18975), .A(n13165), .ZN(P2_U2926) );
  INV_X1 U16342 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14882) );
  AOI22_X1 U16343 ( .A1(n13167), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13166) );
  OAI21_X1 U16344 ( .B1(n14882), .B2(n18975), .A(n13166), .ZN(P2_U2924) );
  AOI22_X1 U16345 ( .A1(n13167), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13168) );
  OAI21_X1 U16346 ( .B1(n13169), .B2(n18975), .A(n13168), .ZN(P2_U2927) );
  AOI22_X1 U16347 ( .A1(n19008), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13170) );
  OAI21_X1 U16348 ( .B1(n13171), .B2(n18975), .A(n13170), .ZN(P2_U2923) );
  AOI22_X1 U16349 ( .A1(n19008), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13172) );
  OAI21_X1 U16350 ( .B1(n13173), .B2(n18975), .A(n13172), .ZN(P2_U2921) );
  OR2_X1 U16351 ( .A1(n13174), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n13175) );
  INV_X1 U16352 ( .A(n13587), .ZN(n20675) );
  NOR2_X1 U16353 ( .A1(n13175), .A2(n20675), .ZN(n13178) );
  INV_X1 U16354 ( .A(n13175), .ZN(n13176) );
  NAND2_X1 U16355 ( .A1(n20678), .A2(n13587), .ZN(n13597) );
  OAI22_X1 U16356 ( .A1(n13178), .A2(n13177), .B1(n13176), .B2(n13597), .ZN(
        P1_U3487) );
  NAND2_X1 U16357 ( .A1(n15580), .A2(n13593), .ZN(n13183) );
  INV_X1 U16358 ( .A(n13179), .ZN(n13181) );
  NAND2_X1 U16359 ( .A1(n13181), .A2(n13180), .ZN(n13182) );
  NAND2_X1 U16360 ( .A1(n13183), .A2(n13182), .ZN(n19757) );
  OR2_X1 U16361 ( .A1(n13184), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n15585) );
  NAND3_X1 U16362 ( .A1(n14129), .A2(n13593), .A3(n15585), .ZN(n13185) );
  AND2_X1 U16363 ( .A1(n13185), .A2(n20677), .ZN(n20681) );
  OR2_X1 U16364 ( .A1(n19757), .A2(n20681), .ZN(n15562) );
  NAND2_X1 U16365 ( .A1(n15562), .A2(n13451), .ZN(n19763) );
  INV_X1 U16366 ( .A(n19763), .ZN(n13200) );
  INV_X1 U16367 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13199) );
  NAND2_X1 U16368 ( .A1(n13187), .A2(n13186), .ZN(n13387) );
  NOR2_X1 U16369 ( .A1(n13188), .A2(n13387), .ZN(n13438) );
  NOR2_X1 U16370 ( .A1(n11269), .A2(n13189), .ZN(n13190) );
  OR2_X1 U16371 ( .A1(n13386), .A2(n13190), .ZN(n13414) );
  NAND2_X1 U16372 ( .A1(n13191), .A2(n20005), .ZN(n13192) );
  NAND2_X1 U16373 ( .A1(n13414), .A2(n13192), .ZN(n13193) );
  MUX2_X1 U16374 ( .A(n13438), .B(n13193), .S(n15580), .Z(n13196) );
  NOR2_X1 U16375 ( .A1(n13377), .A2(n13194), .ZN(n13195) );
  OR2_X1 U16376 ( .A1(n13196), .A2(n13195), .ZN(n13197) );
  NAND2_X1 U16377 ( .A1(n13197), .A2(n11267), .ZN(n15561) );
  OR2_X1 U16378 ( .A1(n15561), .A2(n19763), .ZN(n13198) );
  OAI21_X1 U16379 ( .B1(n13200), .B2(n13199), .A(n13198), .ZN(P1_U3484) );
  INV_X1 U16380 ( .A(n13813), .ZN(n13208) );
  XNOR2_X1 U16381 ( .A(n13822), .B(n13201), .ZN(n13282) );
  OAI22_X1 U16382 ( .A1(n16072), .A2(n13282), .B1(n13818), .B2(n18847), .ZN(
        n13207) );
  OAI21_X1 U16383 ( .B1(n13204), .B2(n13203), .A(n13202), .ZN(n13280) );
  INV_X1 U16384 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13205) );
  OAI22_X1 U16385 ( .A1(n13280), .A2(n16073), .B1(n13205), .B2(n16059), .ZN(
        n13206) );
  AOI211_X1 U16386 ( .C1(n16052), .C2(n13208), .A(n13207), .B(n13206), .ZN(
        n13209) );
  OAI21_X1 U16387 ( .B1(n13222), .B2(n19020), .A(n13209), .ZN(P2_U3012) );
  NAND2_X1 U16388 ( .A1(n14930), .A2(n13210), .ZN(n18937) );
  NOR2_X1 U16389 ( .A1(n13212), .A2(n13211), .ZN(n13213) );
  OR2_X1 U16390 ( .A1(n13214), .A2(n13213), .ZN(n18892) );
  NOR2_X1 U16391 ( .A1(n18954), .A2(n18892), .ZN(n13216) );
  NOR2_X1 U16392 ( .A1(n19716), .A2(n18892), .ZN(n18967) );
  AOI211_X1 U16393 ( .C1(n19716), .C2(n18892), .A(n18968), .B(n18967), .ZN(
        n13215) );
  AOI211_X1 U16394 ( .C1(P2_EAX_REG_0__SCAN_IN), .C2(n18963), .A(n13216), .B(
        n13215), .ZN(n13217) );
  OAI21_X1 U16395 ( .B1(n18972), .B2(n19033), .A(n13217), .ZN(P2_U2919) );
  INV_X1 U16396 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13817) );
  MUX2_X1 U16397 ( .A(n13222), .B(n13817), .S(n13122), .Z(n13223) );
  OAI21_X1 U16398 ( .B1(n19696), .B2(n14854), .A(n13223), .ZN(P2_U2885) );
  OAI21_X1 U16399 ( .B1(n13226), .B2(n13225), .A(n13224), .ZN(n19937) );
  NAND2_X1 U16400 ( .A1(n15580), .A2(n13438), .ZN(n13443) );
  INV_X1 U16401 ( .A(n13227), .ZN(n13228) );
  NAND2_X1 U16402 ( .A1(n13228), .A2(n13266), .ZN(n13229) );
  NAND2_X1 U16403 ( .A1(n13443), .A2(n13229), .ZN(n13230) );
  INV_X1 U16404 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13691) );
  INV_X1 U16405 ( .A(n20025), .ZN(n13231) );
  NAND2_X1 U16406 ( .A1(n13231), .A2(n20005), .ZN(n13551) );
  INV_X1 U16407 ( .A(n13551), .ZN(n13232) );
  OR2_X1 U16408 ( .A1(n14130), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13235) );
  NAND2_X1 U16409 ( .A1(n13551), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13234) );
  NAND2_X1 U16410 ( .A1(n14089), .A2(n13691), .ZN(n13233) );
  NAND2_X1 U16411 ( .A1(n13234), .A2(n13233), .ZN(n13271) );
  NAND2_X1 U16412 ( .A1(n13235), .A2(n13271), .ZN(n19986) );
  OAI222_X1 U16413 ( .A1(n19937), .A2(n14322), .B1(n13691), .B2(n19858), .C1(
        n19986), .C2(n14329), .ZN(P1_U2872) );
  OAI21_X1 U16414 ( .B1(n15404), .B2(n13238), .A(n13237), .ZN(n13241) );
  OAI22_X1 U16415 ( .A1(n15413), .A2(n13239), .B1(n16097), .B2(n18892), .ZN(
        n13240) );
  AOI211_X1 U16416 ( .C1(n16102), .C2(n13242), .A(n13241), .B(n13240), .ZN(
        n13244) );
  MUX2_X1 U16417 ( .A(n15367), .B(n13288), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13243) );
  NAND2_X1 U16418 ( .A1(n13244), .A2(n13243), .ZN(P2_U3046) );
  INV_X1 U16419 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13250) );
  NAND2_X1 U16420 ( .A1(n13245), .A2(n9592), .ZN(n13411) );
  INV_X1 U16421 ( .A(n13411), .ZN(n13246) );
  NAND2_X1 U16422 ( .A1(n19867), .A2(n20005), .ZN(n13523) );
  NAND2_X1 U16423 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15920) );
  INV_X1 U16424 ( .A(n15920), .ZN(n15918) );
  NAND2_X1 U16425 ( .A1(n20578), .A2(n15918), .ZN(n19869) );
  INV_X2 U16426 ( .A(n19869), .ZN(n19884) );
  NOR2_X4 U16427 ( .A1(n19867), .A2(n19884), .ZN(n19871) );
  AOI22_X1 U16428 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13249) );
  OAI21_X1 U16429 ( .B1(n13250), .B2(n13523), .A(n13249), .ZN(P1_U2911) );
  INV_X1 U16430 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13252) );
  AOI22_X1 U16431 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13251) );
  OAI21_X1 U16432 ( .B1(n13252), .B2(n13523), .A(n13251), .ZN(P1_U2906) );
  INV_X1 U16433 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13254) );
  AOI22_X1 U16434 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13253) );
  OAI21_X1 U16435 ( .B1(n13254), .B2(n13523), .A(n13253), .ZN(P1_U2908) );
  INV_X1 U16436 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13256) );
  AOI22_X1 U16437 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13255) );
  OAI21_X1 U16438 ( .B1(n13256), .B2(n13523), .A(n13255), .ZN(P1_U2909) );
  INV_X1 U16439 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13258) );
  AOI22_X1 U16440 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13257) );
  OAI21_X1 U16441 ( .B1(n13258), .B2(n13523), .A(n13257), .ZN(P1_U2910) );
  INV_X1 U16442 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13260) );
  AOI22_X1 U16443 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13259) );
  OAI21_X1 U16444 ( .B1(n13260), .B2(n13523), .A(n13259), .ZN(P1_U2907) );
  INV_X1 U16445 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13262) );
  AOI22_X1 U16446 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13261) );
  OAI21_X1 U16447 ( .B1(n13262), .B2(n13523), .A(n13261), .ZN(P1_U2912) );
  OAI21_X1 U16448 ( .B1(n13264), .B2(n13263), .A(n13340), .ZN(n13631) );
  INV_X1 U16449 ( .A(n13265), .ZN(n14128) );
  AND2_X2 U16450 ( .A1(n14128), .A2(n13266), .ZN(n14101) );
  INV_X1 U16451 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13620) );
  NAND2_X1 U16452 ( .A1(n14101), .A2(n13620), .ZN(n13270) );
  INV_X1 U16453 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19972) );
  NAND2_X1 U16454 ( .A1(n13551), .A2(n19972), .ZN(n13268) );
  NAND2_X1 U16455 ( .A1(n13266), .A2(n13620), .ZN(n13267) );
  NAND3_X1 U16456 ( .A1(n13268), .A2(n14089), .A3(n13267), .ZN(n13269) );
  OR2_X1 U16457 ( .A1(n13272), .A2(n13266), .ZN(n13273) );
  AND2_X1 U16458 ( .A1(n13273), .A2(n13343), .ZN(n13619) );
  OAI22_X1 U16459 ( .A1(n14329), .A2(n13619), .B1(n13620), .B2(n19858), .ZN(
        n13274) );
  INV_X1 U16460 ( .A(n13274), .ZN(n13275) );
  OAI21_X1 U16461 ( .B1(n13631), .B2(n14322), .A(n13275), .ZN(P1_U2871) );
  NAND2_X1 U16462 ( .A1(n13277), .A2(n13276), .ZN(n13279) );
  OAI22_X1 U16463 ( .A1(n15413), .A2(n13280), .B1(n13818), .B2(n18847), .ZN(
        n13284) );
  INV_X1 U16464 ( .A(n13281), .ZN(n15211) );
  NAND2_X1 U16465 ( .A1(n15211), .A2(n13834), .ZN(n13575) );
  OAI21_X1 U16466 ( .B1(n13282), .B2(n15405), .A(n13575), .ZN(n13283) );
  NOR2_X1 U16467 ( .A1(n13284), .A2(n13283), .ZN(n13286) );
  NAND2_X1 U16468 ( .A1(n16115), .A2(n16104), .ZN(n13285) );
  OAI211_X1 U16469 ( .C1(n13816), .C2(n16097), .A(n13286), .B(n13285), .ZN(
        n13294) );
  NOR2_X1 U16470 ( .A1(n15213), .A2(n13287), .ZN(n13292) );
  NAND2_X1 U16471 ( .A1(n15211), .A2(n13290), .ZN(n13289) );
  OAI211_X1 U16472 ( .C1(n13290), .C2(n15213), .A(n13289), .B(n13288), .ZN(
        n13291) );
  MUX2_X1 U16473 ( .A(n13292), .B(n13291), .S(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n13293) );
  OR2_X1 U16474 ( .A1(n13294), .A2(n13293), .ZN(P2_U3044) );
  INV_X1 U16475 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13626) );
  NAND2_X1 U16476 ( .A1(n19950), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n13420) );
  OAI21_X1 U16477 ( .B1(n19938), .B2(n13626), .A(n13420), .ZN(n13295) );
  AOI21_X1 U16478 ( .B1(n15781), .B2(n13626), .A(n13295), .ZN(n13299) );
  OR2_X1 U16479 ( .A1(n13296), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13419) );
  NAND3_X1 U16480 ( .A1(n13419), .A2(n13297), .A3(n19930), .ZN(n13298) );
  OAI211_X1 U16481 ( .C1(n13631), .C2(n20003), .A(n13299), .B(n13298), .ZN(
        P1_U2998) );
  INV_X1 U16482 ( .A(n13301), .ZN(n13302) );
  NAND2_X1 U16483 ( .A1(n13300), .A2(n13302), .ZN(n13304) );
  OAI21_X1 U16484 ( .B1(n13305), .B2(n13304), .A(n13303), .ZN(n18855) );
  NAND2_X1 U16485 ( .A1(n13308), .A2(n13307), .ZN(n13309) );
  NAND2_X1 U16486 ( .A1(n13306), .A2(n13309), .ZN(n19019) );
  MUX2_X1 U16487 ( .A(n19019), .B(n18856), .S(n13122), .Z(n13310) );
  OAI21_X1 U16488 ( .B1(n18855), .B2(n14854), .A(n13310), .ZN(P2_U2883) );
  NAND2_X1 U16489 ( .A1(n12030), .A2(n11267), .ZN(n13313) );
  NAND2_X1 U16490 ( .A1(n13313), .A2(n13379), .ZN(n13311) );
  INV_X1 U16491 ( .A(n13312), .ZN(n13314) );
  NAND2_X1 U16492 ( .A1(n13314), .A2(n14389), .ZN(n14397) );
  NAND2_X1 U16493 ( .A1(n20002), .A2(DATAI_0_), .ZN(n13316) );
  NAND2_X1 U16494 ( .A1(n20001), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13315) );
  AND2_X1 U16495 ( .A1(n13316), .A2(n13315), .ZN(n20010) );
  INV_X1 U16496 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19887) );
  OAI222_X1 U16497 ( .A1(n14404), .A2(n19937), .B1(n14403), .B2(n20010), .C1(
        n14401), .C2(n19887), .ZN(P1_U2904) );
  XNOR2_X1 U16498 ( .A(n19696), .B(n13816), .ZN(n13321) );
  NAND2_X1 U16499 ( .A1(n19026), .A2(n13317), .ZN(n13318) );
  OAI21_X1 U16500 ( .B1(n19026), .B2(n13317), .A(n13318), .ZN(n18966) );
  NOR2_X1 U16501 ( .A1(n18966), .A2(n18967), .ZN(n18965) );
  INV_X1 U16502 ( .A(n13318), .ZN(n13319) );
  NOR2_X1 U16503 ( .A1(n18965), .A2(n13319), .ZN(n13320) );
  NOR2_X1 U16504 ( .A1(n13320), .A2(n13321), .ZN(n13559) );
  AOI21_X1 U16505 ( .B1(n13321), .B2(n13320), .A(n13559), .ZN(n13324) );
  AOI22_X1 U16506 ( .A1(n18937), .A2(n15990), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n18963), .ZN(n13323) );
  INV_X1 U16507 ( .A(n13816), .ZN(n19698) );
  NAND2_X1 U16508 ( .A1(n19698), .A2(n18964), .ZN(n13322) );
  OAI211_X1 U16509 ( .C1(n13324), .C2(n18968), .A(n13323), .B(n13322), .ZN(
        P2_U2917) );
  XOR2_X1 U16510 ( .A(n13303), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13329)
         );
  AND2_X1 U16511 ( .A1(n13306), .A2(n13325), .ZN(n13326) );
  OR2_X1 U16512 ( .A1(n13326), .A2(n9747), .ZN(n18850) );
  INV_X1 U16513 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13327) );
  MUX2_X1 U16514 ( .A(n18850), .B(n13327), .S(n14861), .Z(n13328) );
  OAI21_X1 U16515 ( .B1(n13329), .B2(n14854), .A(n13328), .ZN(P2_U2882) );
  INV_X1 U16516 ( .A(n19304), .ZN(n19690) );
  INV_X1 U16517 ( .A(n12208), .ZN(n15433) );
  MUX2_X1 U16518 ( .A(P2_EBX_REG_3__SCAN_IN), .B(n15433), .S(n14796), .Z(
        n13333) );
  AOI21_X1 U16519 ( .B1(n19690), .B2(n14860), .A(n13333), .ZN(n13334) );
  INV_X1 U16520 ( .A(n13334), .ZN(P2_U2884) );
  AND2_X1 U16521 ( .A1(n11295), .A2(n20585), .ZN(n13335) );
  OR2_X1 U16522 ( .A1(n19916), .A2(n11930), .ZN(n13468) );
  INV_X1 U16523 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13339) );
  NOR2_X2 U16524 ( .A1(n19916), .A2(n9592), .ZN(n19906) );
  INV_X1 U16525 ( .A(n19906), .ZN(n13338) );
  NOR2_X1 U16526 ( .A1(n20002), .A2(n20706), .ZN(n13336) );
  AOI21_X1 U16527 ( .B1(DATAI_15_), .B2(n20002), .A(n13336), .ZN(n14394) );
  INV_X1 U16528 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13337) );
  OAI222_X1 U16529 ( .A1(n13468), .A2(n13339), .B1(n13338), .B2(n14394), .C1(
        n13337), .C2(n13469), .ZN(P1_U2967) );
  OAI21_X1 U16530 ( .B1(n9689), .B2(n11414), .A(n13342), .ZN(n13618) );
  INV_X1 U16531 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13606) );
  NAND2_X1 U16532 ( .A1(n14101), .A2(n13606), .ZN(n13347) );
  NAND2_X1 U16533 ( .A1(n13551), .A2(n19984), .ZN(n13345) );
  NAND2_X1 U16534 ( .A1(n13266), .A2(n13606), .ZN(n13344) );
  NAND3_X1 U16535 ( .A1(n13345), .A2(n14089), .A3(n13344), .ZN(n13346) );
  AND2_X1 U16536 ( .A1(n13347), .A2(n13346), .ZN(n13348) );
  NAND2_X1 U16537 ( .A1(n13349), .A2(n13348), .ZN(n13350) );
  NAND2_X1 U16538 ( .A1(n13544), .A2(n13350), .ZN(n13596) );
  OAI22_X1 U16539 ( .A1(n14329), .A2(n13596), .B1(n13606), .B2(n19858), .ZN(
        n13351) );
  INV_X1 U16540 ( .A(n13351), .ZN(n13352) );
  OAI21_X1 U16541 ( .B1(n13618), .B2(n14322), .A(n13352), .ZN(P1_U2870) );
  INV_X1 U16542 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13609) );
  NOR2_X1 U16543 ( .A1(n19823), .A2(n13609), .ZN(n19975) );
  NOR2_X1 U16544 ( .A1(n19934), .A2(n13612), .ZN(n13353) );
  AOI211_X1 U16545 ( .C1(n19925), .C2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n19975), .B(n13353), .ZN(n13358) );
  OR2_X1 U16546 ( .A1(n13355), .A2(n13354), .ZN(n19974) );
  NAND3_X1 U16547 ( .A1(n19974), .A2(n13356), .A3(n19930), .ZN(n13357) );
  OAI211_X1 U16548 ( .C1(n13618), .C2(n20003), .A(n13358), .B(n13357), .ZN(
        P1_U2997) );
  XNOR2_X1 U16549 ( .A(n13359), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13365) );
  NOR2_X1 U16550 ( .A1(n13360), .A2(n13361), .ZN(n13362) );
  OR2_X1 U16551 ( .A1(n13535), .A2(n13362), .ZN(n18825) );
  INV_X1 U16552 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13363) );
  MUX2_X1 U16553 ( .A(n18825), .B(n13363), .S(n14861), .Z(n13364) );
  OAI21_X1 U16554 ( .B1(n13365), .B2(n14854), .A(n13364), .ZN(P2_U2880) );
  NOR2_X1 U16555 ( .A1(n9747), .A2(n13366), .ZN(n13367) );
  OR2_X1 U16556 ( .A1(n13360), .A2(n13367), .ZN(n18841) );
  NOR2_X1 U16557 ( .A1(n13303), .A2(n10553), .ZN(n13369) );
  INV_X1 U16558 ( .A(n13359), .ZN(n13368) );
  OAI211_X1 U16559 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13369), .A(
        n13368), .B(n14860), .ZN(n13371) );
  NAND2_X1 U16560 ( .A1(n13122), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13370) );
  OAI211_X1 U16561 ( .C1(n18841), .C2(n14861), .A(n13371), .B(n13370), .ZN(
        P2_U2881) );
  NAND2_X1 U16562 ( .A1(n20002), .A2(DATAI_1_), .ZN(n13373) );
  NAND2_X1 U16563 ( .A1(n20001), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13372) );
  AND2_X1 U16564 ( .A1(n13373), .A2(n13372), .ZN(n20019) );
  INV_X1 U16565 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19883) );
  OAI222_X1 U16566 ( .A1(n14404), .A2(n13631), .B1(n14403), .B2(n20019), .C1(
        n14401), .C2(n19883), .ZN(P1_U2903) );
  NAND2_X1 U16567 ( .A1(n20002), .A2(DATAI_2_), .ZN(n13375) );
  NAND2_X1 U16568 ( .A1(n20001), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13374) );
  AND2_X1 U16569 ( .A1(n13375), .A2(n13374), .ZN(n20022) );
  INV_X1 U16570 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19881) );
  OAI222_X1 U16571 ( .A1(n14404), .A2(n13618), .B1(n20022), .B2(n14403), .C1(
        n14401), .C2(n19881), .ZN(P1_U2902) );
  AOI21_X1 U16572 ( .B1(n11930), .B2(n15585), .A(n20585), .ZN(n13376) );
  NAND2_X1 U16573 ( .A1(n13377), .A2(n13376), .ZN(n13385) );
  NAND2_X1 U16574 ( .A1(n9592), .A2(n15585), .ZN(n13599) );
  AND2_X1 U16575 ( .A1(n13599), .A2(n20677), .ZN(n13381) );
  NAND2_X1 U16576 ( .A1(n13379), .A2(n20005), .ZN(n13380) );
  AOI21_X1 U16577 ( .B1(n13378), .B2(n13381), .A(n13380), .ZN(n13382) );
  OR2_X1 U16578 ( .A1(n15580), .A2(n13382), .ZN(n13384) );
  MUX2_X1 U16579 ( .A(n13385), .B(n13384), .S(n13383), .Z(n13394) );
  INV_X1 U16580 ( .A(n13387), .ZN(n13392) );
  INV_X1 U16581 ( .A(n13386), .ZN(n13390) );
  AND2_X1 U16582 ( .A1(n13387), .A2(n20005), .ZN(n13388) );
  NAND2_X1 U16583 ( .A1(n13389), .A2(n13388), .ZN(n13400) );
  AND2_X1 U16584 ( .A1(n13390), .A2(n13400), .ZN(n13391) );
  AOI21_X1 U16585 ( .B1(n15580), .B2(n13392), .A(n13444), .ZN(n13393) );
  NAND2_X1 U16586 ( .A1(n13418), .A2(n13987), .ZN(n19990) );
  NAND2_X1 U16587 ( .A1(n13396), .A2(n13395), .ZN(n13398) );
  NAND2_X1 U16588 ( .A1(n14130), .A2(n11936), .ZN(n13397) );
  OAI211_X1 U16589 ( .C1(n12066), .C2(n14089), .A(n13398), .B(n13397), .ZN(
        n13399) );
  INV_X1 U16590 ( .A(n13399), .ZN(n13402) );
  AND3_X1 U16591 ( .A1(n13402), .A2(n13401), .A3(n13400), .ZN(n13428) );
  NAND2_X1 U16592 ( .A1(n13428), .A2(n13403), .ZN(n13404) );
  NAND2_X1 U16593 ( .A1(n13418), .A2(n13404), .ZN(n14704) );
  INV_X1 U16594 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14536) );
  NOR2_X1 U16595 ( .A1(n14557), .A2(n14534), .ZN(n13408) );
  OR2_X1 U16596 ( .A1(n14704), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13406) );
  OR2_X1 U16597 ( .A1(n13418), .A2(n19950), .ZN(n13405) );
  NAND2_X1 U16598 ( .A1(n13406), .A2(n13405), .ZN(n19970) );
  AOI21_X1 U16599 ( .B1(n19987), .B2(n14536), .A(n19970), .ZN(n19991) );
  INV_X1 U16600 ( .A(n19991), .ZN(n13407) );
  MUX2_X1 U16601 ( .A(n13408), .B(n13407), .S(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n13423) );
  NAND2_X1 U16602 ( .A1(n13409), .A2(n13416), .ZN(n13410) );
  NAND2_X1 U16603 ( .A1(n13411), .A2(n13410), .ZN(n13412) );
  OAI211_X1 U16604 ( .C1(n13416), .C2(n13415), .A(n13413), .B(n13414), .ZN(
        n13417) );
  NAND3_X1 U16605 ( .A1(n13419), .A2(n19973), .A3(n13297), .ZN(n13421) );
  OAI211_X1 U16606 ( .C1(n13619), .C2(n19953), .A(n13421), .B(n13420), .ZN(
        n13422) );
  OR2_X1 U16607 ( .A1(n13423), .A2(n13422), .ZN(P1_U3030) );
  INV_X1 U16608 ( .A(n13425), .ZN(n13426) );
  NOR2_X1 U16609 ( .A1(n13378), .A2(n13426), .ZN(n13427) );
  AND2_X1 U16610 ( .A1(n13428), .A2(n13427), .ZN(n13429) );
  AND2_X1 U16611 ( .A1(n13429), .A2(n12161), .ZN(n13636) );
  XNOR2_X1 U16612 ( .A(n13430), .B(n13431), .ZN(n13442) );
  AND2_X1 U16613 ( .A1(n11279), .A2(n13442), .ZN(n13435) );
  NOR2_X1 U16614 ( .A1(n13433), .A2(n13432), .ZN(n13434) );
  AOI22_X1 U16615 ( .A1(n13636), .A2(n13435), .B1(n13987), .B2(n13434), .ZN(
        n13441) );
  INV_X1 U16616 ( .A(n13436), .ZN(n13437) );
  OR2_X1 U16617 ( .A1(n13438), .A2(n13437), .ZN(n13641) );
  INV_X1 U16618 ( .A(n13442), .ZN(n13439) );
  NAND2_X1 U16619 ( .A1(n13641), .A2(n13439), .ZN(n13440) );
  OAI211_X1 U16620 ( .C1(n13424), .C2(n13636), .A(n13441), .B(n13440), .ZN(
        n13632) );
  INV_X1 U16621 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14540) );
  AOI22_X1 U16622 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n19972), .B2(n14540), .ZN(
        n13463) );
  NOR2_X1 U16623 ( .A1(n20577), .A2(n14536), .ZN(n13462) );
  INV_X1 U16624 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20412) );
  AOI222_X1 U16625 ( .A1(n13632), .A2(n15908), .B1(n13463), .B2(n13462), .C1(
        n20649), .C2(n13442), .ZN(n13455) );
  INV_X1 U16626 ( .A(n13443), .ZN(n13449) );
  INV_X1 U16627 ( .A(n13444), .ZN(n13447) );
  OAI211_X1 U16628 ( .C1(n13987), .C2(n13378), .A(n15570), .B(n20677), .ZN(
        n13446) );
  NAND3_X1 U16629 ( .A1(n11270), .A2(n13383), .A3(n11930), .ZN(n13445) );
  NAND3_X1 U16630 ( .A1(n13447), .A2(n13446), .A3(n13445), .ZN(n13448) );
  NAND2_X1 U16631 ( .A1(n13646), .A2(n13451), .ZN(n13453) );
  NOR2_X1 U16632 ( .A1(n20578), .A2(n15920), .ZN(n13654) );
  NAND2_X1 U16633 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13654), .ZN(n13452) );
  NAND2_X1 U16634 ( .A1(n13453), .A2(n13452), .ZN(n15907) );
  NAND2_X1 U16635 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n15906), .ZN(
        n13454) );
  OAI21_X1 U16636 ( .B1(n13455), .B2(n15906), .A(n13454), .ZN(P1_U3472) );
  INV_X1 U16637 ( .A(n13456), .ZN(n13458) );
  INV_X1 U16638 ( .A(n13430), .ZN(n13457) );
  NAND2_X1 U16639 ( .A1(n13458), .A2(n13457), .ZN(n13460) );
  INV_X1 U16640 ( .A(n13460), .ZN(n13465) );
  INV_X1 U16641 ( .A(n13459), .ZN(n20470) );
  INV_X1 U16642 ( .A(n13636), .ZN(n13984) );
  INV_X1 U16643 ( .A(n13987), .ZN(n15546) );
  OAI22_X1 U16644 ( .A1(n15546), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n13460), .B2(n11280), .ZN(n13461) );
  AOI21_X1 U16645 ( .B1(n20470), .B2(n13984), .A(n13461), .ZN(n15548) );
  INV_X1 U16646 ( .A(n13462), .ZN(n13986) );
  OAI22_X1 U16647 ( .A1(n15548), .A2(n20651), .B1(n13986), .B2(n13463), .ZN(
        n13464) );
  AOI21_X1 U16648 ( .B1(n20649), .B2(n13465), .A(n13464), .ZN(n13467) );
  NAND2_X1 U16649 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n15906), .ZN(
        n13466) );
  OAI21_X1 U16650 ( .B1(n13467), .B2(n15906), .A(n13466), .ZN(P1_U3473) );
  AOI22_X1 U16651 ( .A1(n19922), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n19921), .ZN(n13471) );
  INV_X1 U16652 ( .A(n20010), .ZN(n13470) );
  NAND2_X1 U16653 ( .A1(n19906), .A2(n13470), .ZN(n13488) );
  NAND2_X1 U16654 ( .A1(n13471), .A2(n13488), .ZN(P1_U2937) );
  AOI22_X1 U16655 ( .A1(n19922), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n19921), .ZN(n13473) );
  INV_X1 U16656 ( .A(n20019), .ZN(n13472) );
  NAND2_X1 U16657 ( .A1(n19906), .A2(n13472), .ZN(n13505) );
  NAND2_X1 U16658 ( .A1(n13473), .A2(n13505), .ZN(P1_U2953) );
  AOI22_X1 U16659 ( .A1(n19922), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n19921), .ZN(n13476) );
  NAND2_X1 U16660 ( .A1(n20002), .A2(DATAI_4_), .ZN(n13475) );
  NAND2_X1 U16661 ( .A1(n20001), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13474) );
  AND2_X1 U16662 ( .A1(n13475), .A2(n13474), .ZN(n20029) );
  INV_X1 U16663 ( .A(n20029), .ZN(n15740) );
  NAND2_X1 U16664 ( .A1(n19906), .A2(n15740), .ZN(n13483) );
  NAND2_X1 U16665 ( .A1(n13476), .A2(n13483), .ZN(P1_U2956) );
  AOI22_X1 U16666 ( .A1(n19922), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n19921), .ZN(n13478) );
  INV_X1 U16667 ( .A(n20022), .ZN(n13477) );
  NAND2_X1 U16668 ( .A1(n19906), .A2(n13477), .ZN(n13501) );
  NAND2_X1 U16669 ( .A1(n13478), .A2(n13501), .ZN(P1_U2939) );
  AOI22_X1 U16670 ( .A1(n19922), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n19921), .ZN(n13482) );
  NAND2_X1 U16671 ( .A1(n20002), .A2(DATAI_5_), .ZN(n13480) );
  NAND2_X1 U16672 ( .A1(n20001), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13479) );
  AND2_X1 U16673 ( .A1(n13480), .A2(n13479), .ZN(n20033) );
  INV_X1 U16674 ( .A(n20033), .ZN(n13481) );
  NAND2_X1 U16675 ( .A1(n19906), .A2(n13481), .ZN(n13507) );
  NAND2_X1 U16676 ( .A1(n13482), .A2(n13507), .ZN(P1_U2957) );
  AOI22_X1 U16677 ( .A1(n19922), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n19921), .ZN(n13484) );
  NAND2_X1 U16678 ( .A1(n13484), .A2(n13483), .ZN(P1_U2941) );
  AOI22_X1 U16679 ( .A1(n19922), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n19921), .ZN(n13487) );
  NAND2_X1 U16680 ( .A1(n20002), .A2(DATAI_7_), .ZN(n13486) );
  NAND2_X1 U16681 ( .A1(n20001), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13485) );
  AND2_X1 U16682 ( .A1(n13486), .A2(n13485), .ZN(n20045) );
  INV_X1 U16683 ( .A(n20045), .ZN(n15736) );
  NAND2_X1 U16684 ( .A1(n19906), .A2(n15736), .ZN(n13490) );
  NAND2_X1 U16685 ( .A1(n13487), .A2(n13490), .ZN(P1_U2959) );
  AOI22_X1 U16686 ( .A1(n19922), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n19921), .ZN(n13489) );
  NAND2_X1 U16687 ( .A1(n13489), .A2(n13488), .ZN(P1_U2952) );
  AOI22_X1 U16688 ( .A1(n19922), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n19921), .ZN(n13491) );
  NAND2_X1 U16689 ( .A1(n13491), .A2(n13490), .ZN(P1_U2944) );
  AOI22_X1 U16690 ( .A1(n19922), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n19921), .ZN(n13495) );
  NAND2_X1 U16691 ( .A1(n20002), .A2(DATAI_6_), .ZN(n13493) );
  NAND2_X1 U16692 ( .A1(n20001), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13492) );
  AND2_X1 U16693 ( .A1(n13493), .A2(n13492), .ZN(n20037) );
  INV_X1 U16694 ( .A(n20037), .ZN(n13494) );
  NAND2_X1 U16695 ( .A1(n19906), .A2(n13494), .ZN(n13496) );
  NAND2_X1 U16696 ( .A1(n13495), .A2(n13496), .ZN(P1_U2958) );
  AOI22_X1 U16697 ( .A1(n19922), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n19921), .ZN(n13497) );
  NAND2_X1 U16698 ( .A1(n13497), .A2(n13496), .ZN(P1_U2943) );
  AOI22_X1 U16699 ( .A1(n19922), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n19921), .ZN(n13500) );
  NAND2_X1 U16700 ( .A1(n20002), .A2(DATAI_3_), .ZN(n13499) );
  NAND2_X1 U16701 ( .A1(n20001), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13498) );
  AND2_X1 U16702 ( .A1(n13499), .A2(n13498), .ZN(n20026) );
  INV_X1 U16703 ( .A(n20026), .ZN(n15745) );
  NAND2_X1 U16704 ( .A1(n19906), .A2(n15745), .ZN(n13503) );
  NAND2_X1 U16705 ( .A1(n13500), .A2(n13503), .ZN(P1_U2955) );
  AOI22_X1 U16706 ( .A1(n19922), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n19921), .ZN(n13502) );
  NAND2_X1 U16707 ( .A1(n13502), .A2(n13501), .ZN(P1_U2954) );
  AOI22_X1 U16708 ( .A1(n19922), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n19921), .ZN(n13504) );
  NAND2_X1 U16709 ( .A1(n13504), .A2(n13503), .ZN(P1_U2940) );
  AOI22_X1 U16710 ( .A1(n19922), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n19921), .ZN(n13506) );
  NAND2_X1 U16711 ( .A1(n13506), .A2(n13505), .ZN(P1_U2938) );
  AOI22_X1 U16712 ( .A1(n19922), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n19921), .ZN(n13508) );
  NAND2_X1 U16713 ( .A1(n13508), .A2(n13507), .ZN(P1_U2942) );
  INV_X1 U16714 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13510) );
  AOI22_X1 U16715 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13509) );
  OAI21_X1 U16716 ( .B1(n13510), .B2(n13523), .A(n13509), .ZN(P1_U2913) );
  INV_X1 U16717 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13512) );
  AOI22_X1 U16718 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13511) );
  OAI21_X1 U16719 ( .B1(n13512), .B2(n13523), .A(n13511), .ZN(P1_U2916) );
  INV_X1 U16720 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13514) );
  AOI22_X1 U16721 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13513) );
  OAI21_X1 U16722 ( .B1(n13514), .B2(n13523), .A(n13513), .ZN(P1_U2917) );
  INV_X1 U16723 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13516) );
  AOI22_X1 U16724 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13515) );
  OAI21_X1 U16725 ( .B1(n13516), .B2(n13523), .A(n13515), .ZN(P1_U2915) );
  INV_X1 U16726 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13518) );
  AOI22_X1 U16727 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13517) );
  OAI21_X1 U16728 ( .B1(n13518), .B2(n13523), .A(n13517), .ZN(P1_U2919) );
  INV_X1 U16729 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13520) );
  AOI22_X1 U16730 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13519) );
  OAI21_X1 U16731 ( .B1(n13520), .B2(n13523), .A(n13519), .ZN(P1_U2914) );
  AOI22_X1 U16732 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13521) );
  OAI21_X1 U16733 ( .B1(n14380), .B2(n13523), .A(n13521), .ZN(P1_U2918) );
  INV_X1 U16734 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13524) );
  AOI22_X1 U16735 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13522) );
  OAI21_X1 U16736 ( .B1(n13524), .B2(n13523), .A(n13522), .ZN(P1_U2920) );
  OR2_X1 U16737 ( .A1(n13526), .A2(n13525), .ZN(n13527) );
  NAND2_X1 U16738 ( .A1(n13528), .A2(n13527), .ZN(n19962) );
  XOR2_X1 U16739 ( .A(n13529), .B(n13530), .Z(n13541) );
  NAND2_X1 U16740 ( .A1(n19950), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n19959) );
  NAND2_X1 U16741 ( .A1(n19925), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13531) );
  OAI211_X1 U16742 ( .C1(n19934), .C2(n13687), .A(n19959), .B(n13531), .ZN(
        n13532) );
  AOI21_X1 U16743 ( .B1(n13541), .B2(n19942), .A(n13532), .ZN(n13533) );
  OAI21_X1 U16744 ( .B1(n19944), .B2(n19962), .A(n13533), .ZN(P1_U2996) );
  OAI21_X1 U16745 ( .B1(n13535), .B2(n13534), .A(n13674), .ZN(n18819) );
  NAND2_X1 U16746 ( .A1(n13359), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13537) );
  INV_X1 U16747 ( .A(n13537), .ZN(n13725) );
  OR2_X1 U16748 ( .A1(n13537), .A2(n13536), .ZN(n13671) );
  OAI211_X1 U16749 ( .C1(n13725), .C2(n13538), .A(n14860), .B(n13671), .ZN(
        n13540) );
  INV_X1 U16750 ( .A(n14796), .ZN(n14861) );
  NAND2_X1 U16751 ( .A1(n14861), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13539) );
  OAI211_X1 U16752 ( .C1(n18819), .C2(n13122), .A(n13540), .B(n13539), .ZN(
        P2_U2879) );
  INV_X1 U16753 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19879) );
  OAI222_X1 U16754 ( .A1(n14404), .A2(n13690), .B1(n14403), .B2(n20026), .C1(
        n14401), .C2(n19879), .ZN(P1_U2901) );
  MUX2_X1 U16755 ( .A(n14107), .B(n14089), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13542) );
  OAI21_X1 U16756 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14130), .A(
        n13542), .ZN(n13543) );
  AND2_X1 U16757 ( .A1(n13544), .A2(n13543), .ZN(n13545) );
  OR2_X1 U16758 ( .A1(n13545), .A2(n13556), .ZN(n19958) );
  INV_X1 U16759 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n20690) );
  OAI222_X1 U16760 ( .A1(n19958), .A2(n14329), .B1(n19858), .B2(n20690), .C1(
        n13690), .C2(n14322), .ZN(P1_U2869) );
  NAND2_X1 U16761 ( .A1(n13548), .A2(n13549), .ZN(n13550) );
  AND2_X1 U16762 ( .A1(n13547), .A2(n13550), .ZN(n19929) );
  INV_X1 U16763 ( .A(n19929), .ZN(n13558) );
  INV_X1 U16764 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n19834) );
  MUX2_X1 U16765 ( .A(n14113), .B(n13551), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n13554) );
  NAND2_X1 U16766 ( .A1(n14129), .A2(n13232), .ZN(n14097) );
  NAND2_X1 U16767 ( .A1(n14129), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13552) );
  AND2_X1 U16768 ( .A1(n14097), .A2(n13552), .ZN(n13553) );
  NAND2_X1 U16769 ( .A1(n13554), .A2(n13553), .ZN(n13555) );
  OR2_X1 U16770 ( .A1(n13556), .A2(n13555), .ZN(n13557) );
  NAND2_X1 U16771 ( .A1(n15898), .A2(n13557), .ZN(n19952) );
  OAI222_X1 U16772 ( .A1(n13558), .A2(n14322), .B1(n19858), .B2(n19834), .C1(
        n19952), .C2(n14329), .ZN(P1_U2868) );
  INV_X1 U16773 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19877) );
  OAI222_X1 U16774 ( .A1(n14404), .A2(n13558), .B1(n14403), .B2(n20029), .C1(
        n14401), .C2(n19877), .ZN(P1_U2900) );
  AOI21_X1 U16775 ( .B1(n13816), .B2(n19696), .A(n13559), .ZN(n18958) );
  OR2_X1 U16776 ( .A1(n13561), .A2(n13560), .ZN(n13563) );
  NAND2_X1 U16777 ( .A1(n13563), .A2(n13562), .ZN(n18955) );
  XNOR2_X1 U16778 ( .A(n19304), .B(n18955), .ZN(n18959) );
  NOR2_X1 U16779 ( .A1(n18958), .A2(n18959), .ZN(n18957) );
  INV_X1 U16780 ( .A(n18955), .ZN(n19689) );
  NOR2_X1 U16781 ( .A1(n19690), .A2(n19689), .ZN(n13566) );
  INV_X1 U16782 ( .A(n13562), .ZN(n13564) );
  XNOR2_X1 U16783 ( .A(n13565), .B(n13564), .ZN(n13831) );
  OAI21_X1 U16784 ( .B1(n18957), .B2(n13566), .A(n13831), .ZN(n18947) );
  XOR2_X1 U16785 ( .A(n18855), .B(n18947), .Z(n13569) );
  INV_X1 U16786 ( .A(n13831), .ZN(n18859) );
  AOI22_X1 U16787 ( .A1(n18964), .A2(n18859), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n18963), .ZN(n13568) );
  NAND2_X1 U16788 ( .A1(n18937), .A2(n15982), .ZN(n13567) );
  OAI211_X1 U16789 ( .C1(n13569), .C2(n18968), .A(n13568), .B(n13567), .ZN(
        P2_U2915) );
  XNOR2_X1 U16790 ( .A(n13571), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13572) );
  XNOR2_X1 U16791 ( .A(n13570), .B(n13572), .ZN(n13751) );
  XNOR2_X1 U16792 ( .A(n13573), .B(n13574), .ZN(n13747) );
  INV_X1 U16793 ( .A(n13747), .ZN(n13582) );
  NAND2_X1 U16794 ( .A1(n19011), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n13745) );
  INV_X1 U16795 ( .A(n13745), .ZN(n13579) );
  NOR2_X1 U16796 ( .A1(n13834), .A2(n16099), .ZN(n13577) );
  NAND2_X1 U16797 ( .A1(n13576), .A2(n13575), .ZN(n15364) );
  MUX2_X1 U16798 ( .A(n13577), .B(n15364), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n13578) );
  AOI211_X1 U16799 ( .C1(n15433), .C2(n16104), .A(n13579), .B(n13578), .ZN(
        n13580) );
  OAI21_X1 U16800 ( .B1(n18955), .B2(n16097), .A(n13580), .ZN(n13581) );
  AOI21_X1 U16801 ( .B1(n13582), .B2(n16105), .A(n13581), .ZN(n13583) );
  OAI21_X1 U16802 ( .B1(n13751), .B2(n15405), .A(n13583), .ZN(P2_U3043) );
  NAND2_X1 U16803 ( .A1(n20581), .A2(n20577), .ZN(n15915) );
  INV_X1 U16804 ( .A(n15915), .ZN(n20680) );
  NAND2_X1 U16805 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20680), .ZN(n15914) );
  NAND2_X1 U16806 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20578), .ZN(n13584) );
  OAI22_X1 U16807 ( .A1(n20578), .A2(n15914), .B1(n13584), .B2(n11471), .ZN(
        n13585) );
  NOR2_X1 U16808 ( .A1(n13585), .A2(n19950), .ZN(n13586) );
  AND2_X1 U16809 ( .A1(n13587), .A2(n13586), .ZN(n13588) );
  INV_X1 U16810 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14414) );
  NOR2_X1 U16811 ( .A1(n13589), .A2(n14414), .ZN(n13590) );
  XNOR2_X1 U16812 ( .A(n13590), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14021) );
  NOR2_X1 U16813 ( .A1(n14021), .A2(n20577), .ZN(n13591) );
  INV_X1 U16814 ( .A(n13597), .ZN(n13592) );
  NOR2_X1 U16815 ( .A1(n13593), .A2(n13592), .ZN(n13594) );
  OR2_X1 U16816 ( .A1(n19811), .A2(n13594), .ZN(n19837) );
  INV_X1 U16817 ( .A(n19837), .ZN(n13696) );
  AND2_X1 U16818 ( .A1(n11930), .A2(n13597), .ZN(n13595) );
  AND2_X1 U16819 ( .A1(n13595), .A2(n11270), .ZN(n13681) );
  INV_X1 U16820 ( .A(n13681), .ZN(n19829) );
  INV_X1 U16821 ( .A(n13596), .ZN(n19976) );
  AND2_X1 U16822 ( .A1(n11930), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13600) );
  NAND2_X1 U16823 ( .A1(n20677), .A2(n20468), .ZN(n13598) );
  INV_X1 U16824 ( .A(n13598), .ZN(n15571) );
  AND2_X1 U16825 ( .A1(n13599), .A2(n15571), .ZN(n13604) );
  INV_X1 U16826 ( .A(n13600), .ZN(n13601) );
  NAND2_X1 U16827 ( .A1(n13601), .A2(n13603), .ZN(n13602) );
  NAND2_X1 U16828 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n13680) );
  OAI21_X1 U16829 ( .B1(P1_REIP_REG_2__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .A(n13680), .ZN(n13605) );
  OAI22_X1 U16830 ( .A1(n13606), .A2(n19833), .B1(n19820), .B2(n13605), .ZN(
        n13607) );
  AOI21_X1 U16831 ( .B1(n19976), .B2(n19815), .A(n13607), .ZN(n13608) );
  OAI21_X1 U16832 ( .B1(n13848), .B2(n13609), .A(n13608), .ZN(n13610) );
  AOI21_X1 U16833 ( .B1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19832), .A(
        n13610), .ZN(n13615) );
  AND2_X1 U16834 ( .A1(n14021), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13611) );
  INV_X1 U16835 ( .A(n13612), .ZN(n13613) );
  NAND2_X1 U16836 ( .A1(n19816), .A2(n13613), .ZN(n13614) );
  OAI211_X1 U16837 ( .C1(n13424), .C2(n19829), .A(n13615), .B(n13614), .ZN(
        n13616) );
  INV_X1 U16838 ( .A(n13616), .ZN(n13617) );
  OAI21_X1 U16839 ( .B1(n13618), .B2(n13696), .A(n13617), .ZN(P1_U2838) );
  INV_X1 U16840 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13624) );
  INV_X1 U16841 ( .A(n13619), .ZN(n13622) );
  OAI22_X1 U16842 ( .A1(n13620), .A2(n19833), .B1(n19820), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n13621) );
  AOI21_X1 U16843 ( .B1(n13622), .B2(n19815), .A(n13621), .ZN(n13623) );
  OAI21_X1 U16844 ( .B1(n13848), .B2(n13624), .A(n13623), .ZN(n13625) );
  AOI21_X1 U16845 ( .B1(n19816), .B2(n13626), .A(n13625), .ZN(n13628) );
  NAND2_X1 U16846 ( .A1(n19832), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13627) );
  OAI211_X1 U16847 ( .C1(n13459), .C2(n19829), .A(n13628), .B(n13627), .ZN(
        n13629) );
  INV_X1 U16848 ( .A(n13629), .ZN(n13630) );
  OAI21_X1 U16849 ( .B1(n13631), .B2(n13696), .A(n13630), .ZN(P1_U2839) );
  NOR2_X1 U16850 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20577), .ZN(n13653) );
  MUX2_X1 U16851 ( .A(n13632), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15553), .Z(n15555) );
  AOI22_X1 U16852 ( .A1(n13653), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15555), .B2(n20577), .ZN(n13649) );
  XNOR2_X1 U16853 ( .A(n13432), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13644) );
  NAND2_X1 U16854 ( .A1(n13430), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13634) );
  NAND2_X1 U16855 ( .A1(n13634), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13635) );
  NAND2_X1 U16856 ( .A1(n11331), .A2(n13635), .ZN(n20650) );
  NAND3_X1 U16857 ( .A1(n13636), .A2(n11279), .A3(n20650), .ZN(n13643) );
  MUX2_X1 U16858 ( .A(n13637), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n13430), .Z(n13639) );
  NOR2_X1 U16859 ( .A1(n13639), .A2(n13638), .ZN(n13640) );
  NAND2_X1 U16860 ( .A1(n13641), .A2(n13640), .ZN(n13642) );
  OAI211_X1 U16861 ( .C1(n15546), .C2(n13644), .A(n13643), .B(n13642), .ZN(
        n13645) );
  AOI21_X1 U16862 ( .B1(n9664), .B2(n13984), .A(n13645), .ZN(n20652) );
  MUX2_X1 U16863 ( .A(n10048), .B(n20652), .S(n13646), .Z(n15556) );
  INV_X1 U16864 ( .A(n15556), .ZN(n13647) );
  AOI22_X1 U16865 ( .A1(n13647), .A2(n20577), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13653), .ZN(n13648) );
  INV_X1 U16866 ( .A(n20153), .ZN(n20410) );
  NOR2_X1 U16867 ( .A1(n11416), .A2(n20410), .ZN(n13650) );
  XOR2_X1 U16868 ( .A(n11469), .B(n13650), .Z(n19830) );
  NOR2_X1 U16869 ( .A1(n19830), .A2(n12161), .ZN(n15909) );
  OAI21_X1 U16870 ( .B1(n15909), .B2(n15553), .A(n20577), .ZN(n13651) );
  AOI21_X1 U16871 ( .B1(n15553), .B2(n11469), .A(n13651), .ZN(n13652) );
  AOI21_X1 U16872 ( .B1(n13653), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13652), .ZN(n15567) );
  OAI21_X1 U16873 ( .B1(n15565), .B2(n13456), .A(n15567), .ZN(n15575) );
  OAI21_X1 U16874 ( .B1(n15575), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13654), .ZN(
        n13655) );
  NAND2_X1 U16875 ( .A1(n13655), .A2(n20052), .ZN(n19999) );
  OR2_X1 U16876 ( .A1(n13657), .A2(n20468), .ZN(n20302) );
  NAND2_X1 U16877 ( .A1(n13657), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20521) );
  OAI22_X1 U16878 ( .A1(n20465), .A2(n20302), .B1(n20249), .B2(n20521), .ZN(
        n13659) );
  INV_X1 U16879 ( .A(n13656), .ZN(n13658) );
  NAND2_X1 U16880 ( .A1(n13659), .A2(n20380), .ZN(n13661) );
  AOI21_X1 U16881 ( .B1(n20004), .B2(n20468), .A(n20515), .ZN(n13660) );
  NAND2_X1 U16882 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20412), .ZN(n20659) );
  AOI22_X1 U16883 ( .A1(n13661), .A2(n13660), .B1(n20659), .B2(n9664), .ZN(
        n13663) );
  NAND2_X1 U16884 ( .A1(n20664), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13662) );
  OAI21_X1 U16885 ( .B1(n20664), .B2(n13663), .A(n13662), .ZN(P1_U3475) );
  NOR2_X1 U16886 ( .A1(n13657), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20441) );
  NOR2_X1 U16887 ( .A1(n20441), .A2(n20515), .ZN(n13664) );
  AOI22_X1 U16888 ( .A1(n13664), .A2(n20521), .B1(n20470), .B2(n20659), .ZN(
        n13666) );
  NAND2_X1 U16889 ( .A1(n20664), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13665) );
  OAI21_X1 U16890 ( .B1(n20664), .B2(n13666), .A(n13665), .ZN(P1_U3477) );
  XOR2_X1 U16891 ( .A(n20521), .B(n13656), .Z(n13667) );
  INV_X1 U16892 ( .A(n13424), .ZN(n20007) );
  AOI22_X1 U16893 ( .A1(n13667), .A2(n20657), .B1(n20007), .B2(n20659), .ZN(
        n13669) );
  NAND2_X1 U16894 ( .A1(n20664), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13668) );
  OAI21_X1 U16895 ( .B1(n20664), .B2(n13669), .A(n13668), .ZN(P1_U3476) );
  INV_X1 U16896 ( .A(n13671), .ZN(n13673) );
  OR2_X1 U16897 ( .A1(n13671), .A2(n13670), .ZN(n13739) );
  OAI211_X1 U16898 ( .C1(n13673), .C2(n13672), .A(n14860), .B(n13739), .ZN(
        n13679) );
  NAND2_X1 U16899 ( .A1(n13675), .A2(n13674), .ZN(n13677) );
  INV_X1 U16900 ( .A(n9752), .ZN(n13676) );
  AND2_X1 U16901 ( .A1(n13677), .A2(n13676), .ZN(n18806) );
  NAND2_X1 U16902 ( .A1(n18806), .A2(n14796), .ZN(n13678) );
  OAI211_X1 U16903 ( .C1(n14796), .C2(n10777), .A(n13679), .B(n13678), .ZN(
        P2_U2878) );
  NOR2_X1 U16904 ( .A1(n19820), .A2(n13680), .ZN(n19827) );
  INV_X1 U16905 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20602) );
  NAND2_X1 U16906 ( .A1(n9664), .A2(n13681), .ZN(n13686) );
  OAI221_X1 U16907 ( .B1(n19820), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n19820), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n13848), .ZN(n13682) );
  AOI22_X1 U16908 ( .A1(n19818), .A2(P1_EBX_REG_3__SCAN_IN), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n13682), .ZN(n13683) );
  OAI21_X1 U16909 ( .B1(n19958), .B2(n19835), .A(n13683), .ZN(n13684) );
  AOI21_X1 U16910 ( .B1(n19832), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13684), .ZN(n13685) );
  OAI211_X1 U16911 ( .C1(n19828), .C2(n13687), .A(n13686), .B(n13685), .ZN(
        n13688) );
  AOI21_X1 U16912 ( .B1(n19827), .B2(n20602), .A(n13688), .ZN(n13689) );
  OAI21_X1 U16913 ( .B1(n13690), .B2(n13696), .A(n13689), .ZN(P1_U2837) );
  OAI22_X1 U16914 ( .A1(n19986), .A2(n19835), .B1(n19833), .B2(n13691), .ZN(
        n13694) );
  INV_X1 U16915 ( .A(n20660), .ZN(n20115) );
  OAI21_X1 U16916 ( .B1(n19832), .B2(n19816), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13692) );
  OAI21_X1 U16917 ( .B1(n20115), .B2(n19829), .A(n13692), .ZN(n13693) );
  AOI211_X1 U16918 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(n19806), .A(n13694), .B(
        n13693), .ZN(n13695) );
  OAI21_X1 U16919 ( .B1(n13696), .B2(n19937), .A(n13695), .ZN(P1_U2840) );
  OR2_X1 U16920 ( .A1(n13697), .A2(n13731), .ZN(n13698) );
  NAND2_X1 U16921 ( .A1(n13699), .A2(n13698), .ZN(n18751) );
  NAND2_X1 U16922 ( .A1(n13359), .A2(n13700), .ZN(n13726) );
  INV_X1 U16923 ( .A(n13726), .ZN(n13703) );
  OAI211_X1 U16924 ( .C1(n13703), .C2(n13702), .A(n14860), .B(n13701), .ZN(
        n13705) );
  NAND2_X1 U16925 ( .A1(n14861), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13704) );
  OAI211_X1 U16926 ( .C1(n18751), .C2(n14861), .A(n13705), .B(n13704), .ZN(
        P2_U2873) );
  NOR2_X2 U16927 ( .A1(n19540), .A2(n19187), .ZN(n19299) );
  OAI21_X1 U16928 ( .B1(n19247), .B2(n19299), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13707) );
  NAND2_X1 U16929 ( .A1(n19693), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19217) );
  INV_X1 U16930 ( .A(n19217), .ZN(n19270) );
  NAND2_X1 U16931 ( .A1(n19189), .A2(n19270), .ZN(n13706) );
  NAND2_X1 U16932 ( .A1(n13707), .A2(n13706), .ZN(n13714) );
  OAI21_X1 U16933 ( .B1(n13718), .B2(n19733), .A(n19732), .ZN(n13712) );
  INV_X1 U16934 ( .A(n19536), .ZN(n19542) );
  NOR3_X2 U16935 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19542), .ZN(n19262) );
  INV_X1 U16936 ( .A(n19262), .ZN(n13711) );
  AOI21_X1 U16937 ( .B1(n19601), .B2(n19733), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19739) );
  AND2_X1 U16938 ( .A1(n19739), .A2(n19713), .ZN(n13709) );
  AOI21_X1 U16939 ( .B1(n13712), .B2(n13711), .A(n19338), .ZN(n13713) );
  INV_X1 U16940 ( .A(n19264), .ZN(n19251) );
  AOI22_X1 U16941 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19062), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19061), .ZN(n19556) );
  AOI22_X1 U16942 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19062), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19061), .ZN(n19441) );
  INV_X1 U16943 ( .A(n19441), .ZN(n19553) );
  AOI22_X1 U16944 ( .A1(n19247), .A2(n19438), .B1(n19299), .B2(n19553), .ZN(
        n13722) );
  OAI21_X1 U16945 ( .B1(n13718), .B2(n19262), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13719) );
  OAI21_X1 U16946 ( .B1(n19217), .B2(n19370), .A(n13719), .ZN(n19263) );
  NOR2_X2 U16947 ( .A1(n18973), .A2(n19338), .ZN(n19552) );
  AOI22_X1 U16948 ( .A1(n19263), .A2(n19552), .B1(n19551), .B2(n19262), .ZN(
        n13721) );
  OAI211_X1 U16949 ( .C1(n19251), .C2(n13723), .A(n13722), .B(n13721), .ZN(
        P2_U3097) );
  AND2_X1 U16950 ( .A1(n13725), .A2(n13724), .ZN(n13728) );
  OAI211_X1 U16951 ( .C1(n13728), .C2(n13727), .A(n13726), .B(n14860), .ZN(
        n13735) );
  NAND2_X1 U16952 ( .A1(n13730), .A2(n13729), .ZN(n13733) );
  INV_X1 U16953 ( .A(n13731), .ZN(n13732) );
  AND2_X1 U16954 ( .A1(n13733), .A2(n13732), .ZN(n16029) );
  NAND2_X1 U16955 ( .A1(n16029), .A2(n14796), .ZN(n13734) );
  OAI211_X1 U16956 ( .C1(n14796), .C2(n10779), .A(n13735), .B(n13734), .ZN(
        P2_U2874) );
  OR2_X1 U16957 ( .A1(n13736), .A2(n9752), .ZN(n13737) );
  NAND2_X1 U16958 ( .A1(n13737), .A2(n13779), .ZN(n18793) );
  INV_X1 U16959 ( .A(n13739), .ZN(n13742) );
  NOR2_X1 U16960 ( .A1(n13739), .A2(n13738), .ZN(n13778) );
  INV_X1 U16961 ( .A(n13778), .ZN(n13740) );
  OAI211_X1 U16962 ( .C1(n13742), .C2(n13741), .A(n13740), .B(n14860), .ZN(
        n13744) );
  NAND2_X1 U16963 ( .A1(n14861), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n13743) );
  OAI211_X1 U16964 ( .C1(n18793), .C2(n13122), .A(n13744), .B(n13743), .ZN(
        P2_U2877) );
  NAND2_X1 U16965 ( .A1(n16052), .A2(n13755), .ZN(n13746) );
  OAI211_X1 U16966 ( .C1(n20796), .C2(n16059), .A(n13746), .B(n13745), .ZN(
        n13749) );
  NOR2_X1 U16967 ( .A1(n13747), .A2(n16073), .ZN(n13748) );
  AOI211_X1 U16968 ( .C1(n16067), .C2(n15433), .A(n13749), .B(n13748), .ZN(
        n13750) );
  OAI21_X1 U16969 ( .B1(n16072), .B2(n13751), .A(n13750), .ZN(P2_U3011) );
  INV_X1 U16970 ( .A(n18897), .ZN(n13826) );
  NAND2_X1 U16971 ( .A1(n9828), .A2(n13753), .ZN(n13754) );
  XNOR2_X1 U16972 ( .A(n13755), .B(n13754), .ZN(n13756) );
  NAND2_X1 U16973 ( .A1(n13756), .A2(n18882), .ZN(n13763) );
  INV_X1 U16974 ( .A(n18871), .ZN(n18896) );
  OAI22_X1 U16975 ( .A1(n20796), .A2(n18874), .B1(n18893), .B2(n18955), .ZN(
        n13758) );
  NOR2_X1 U16976 ( .A1(n18849), .A2(n10536), .ZN(n13757) );
  AOI211_X1 U16977 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n18889), .A(n13758), .B(
        n13757), .ZN(n13759) );
  OAI21_X1 U16978 ( .B1(n13760), .B2(n18888), .A(n13759), .ZN(n13761) );
  AOI21_X1 U16979 ( .B1(n15433), .B2(n18896), .A(n13761), .ZN(n13762) );
  OAI211_X1 U16980 ( .C1(n19304), .C2(n13826), .A(n13763), .B(n13762), .ZN(
        P2_U2852) );
  AOI21_X1 U16981 ( .B1(n13765), .B2(n13547), .A(n11523), .ZN(n19855) );
  INV_X1 U16982 ( .A(n19855), .ZN(n13767) );
  OAI222_X1 U16983 ( .A1(n13767), .A2(n14404), .B1(n20033), .B2(n14403), .C1(
        n13766), .C2(n14401), .ZN(P1_U2899) );
  AND2_X1 U16984 ( .A1(n13778), .A2(n13777), .ZN(n13775) );
  XNOR2_X1 U16985 ( .A(n13775), .B(n13768), .ZN(n13774) );
  OR2_X1 U16986 ( .A1(n13770), .A2(n13769), .ZN(n13771) );
  NAND2_X1 U16987 ( .A1(n13771), .A2(n13729), .ZN(n18772) );
  INV_X1 U16988 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n13772) );
  MUX2_X1 U16989 ( .A(n18772), .B(n13772), .S(n14861), .Z(n13773) );
  OAI21_X1 U16990 ( .B1(n13774), .B2(n14854), .A(n13773), .ZN(P2_U2875) );
  INV_X1 U16991 ( .A(n13775), .ZN(n13776) );
  OAI211_X1 U16992 ( .C1(n13778), .C2(n13777), .A(n13776), .B(n14860), .ZN(
        n13784) );
  NAND2_X1 U16993 ( .A1(n13780), .A2(n13779), .ZN(n13782) );
  INV_X1 U16994 ( .A(n13769), .ZN(n13781) );
  AND2_X1 U16995 ( .A1(n13782), .A2(n13781), .ZN(n18773) );
  NAND2_X1 U16996 ( .A1(n18773), .A2(n14796), .ZN(n13783) );
  OAI211_X1 U16997 ( .C1(n14796), .C2(n10001), .A(n13784), .B(n13783), .ZN(
        P2_U2876) );
  INV_X1 U16998 ( .A(n13701), .ZN(n13788) );
  INV_X1 U16999 ( .A(n13785), .ZN(n13786) );
  OAI211_X1 U17000 ( .C1(n13788), .C2(n13787), .A(n13786), .B(n14860), .ZN(
        n13790) );
  NAND2_X1 U17001 ( .A1(n18733), .A2(n14796), .ZN(n13789) );
  OAI211_X1 U17002 ( .C1(n14796), .C2(n10353), .A(n13790), .B(n13789), .ZN(
        P2_U2872) );
  XOR2_X1 U17003 ( .A(n13764), .B(n13791), .Z(n19849) );
  INV_X1 U17004 ( .A(n19849), .ZN(n13792) );
  OAI222_X1 U17005 ( .A1(n14404), .A2(n13792), .B1(n19874), .B2(n14401), .C1(
        n14403), .C2(n20037), .ZN(P1_U2898) );
  AOI21_X1 U17006 ( .B1(n13796), .B2(n13793), .A(n13795), .ZN(n15797) );
  INV_X1 U17007 ( .A(n15797), .ZN(n19796) );
  INV_X1 U17008 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n19857) );
  NAND2_X1 U17009 ( .A1(n13266), .A2(n19857), .ZN(n13798) );
  NAND2_X1 U17010 ( .A1(n14089), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13797) );
  NAND3_X1 U17011 ( .A1(n13798), .A2(n13551), .A3(n13797), .ZN(n13799) );
  OAI21_X1 U17012 ( .B1(n14107), .B2(P1_EBX_REG_5__SCAN_IN), .A(n13799), .ZN(
        n15899) );
  MUX2_X1 U17013 ( .A(n14113), .B(n13551), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n13802) );
  NAND2_X1 U17014 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14129), .ZN(
        n13800) );
  AND2_X1 U17015 ( .A1(n14097), .A2(n13800), .ZN(n13801) );
  NAND2_X1 U17016 ( .A1(n13802), .A2(n13801), .ZN(n15889) );
  INV_X1 U17017 ( .A(n14107), .ZN(n13803) );
  INV_X1 U17018 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n19789) );
  NAND2_X1 U17019 ( .A1(n13803), .A2(n19789), .ZN(n13807) );
  NAND2_X1 U17020 ( .A1(n13266), .A2(n19789), .ZN(n13805) );
  NAND2_X1 U17021 ( .A1(n14089), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13804) );
  NAND3_X1 U17022 ( .A1(n13805), .A2(n13551), .A3(n13804), .ZN(n13806) );
  INV_X1 U17023 ( .A(n15889), .ZN(n13810) );
  INV_X1 U17024 ( .A(n13808), .ZN(n13809) );
  OAI21_X1 U17025 ( .B1(n15896), .B2(n13810), .A(n13809), .ZN(n13811) );
  AND2_X1 U17026 ( .A1(n9862), .A2(n13811), .ZN(n19800) );
  INV_X1 U17027 ( .A(n19858), .ZN(n14303) );
  AOI22_X1 U17028 ( .A1(n19800), .A2(n19853), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n14303), .ZN(n13812) );
  OAI21_X1 U17029 ( .B1(n19796), .B2(n14322), .A(n13812), .ZN(P1_U2865) );
  NOR2_X1 U17030 ( .A1(n18865), .A2(n15421), .ZN(n13814) );
  XNOR2_X1 U17031 ( .A(n13814), .B(n13813), .ZN(n13815) );
  NAND2_X1 U17032 ( .A1(n13815), .A2(n18882), .ZN(n13825) );
  OAI22_X1 U17033 ( .A1(n18857), .A2(n13817), .B1(n13816), .B2(n18893), .ZN(
        n13820) );
  NOR2_X1 U17034 ( .A1(n18849), .A2(n13818), .ZN(n13819) );
  AOI211_X1 U17035 ( .C1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .C2(n18901), .A(
        n13820), .B(n13819), .ZN(n13821) );
  OAI21_X1 U17036 ( .B1(n13822), .B2(n18888), .A(n13821), .ZN(n13823) );
  AOI21_X1 U17037 ( .B1(n16115), .B2(n18896), .A(n13823), .ZN(n13824) );
  OAI211_X1 U17038 ( .C1(n13826), .C2(n19696), .A(n13825), .B(n13824), .ZN(
        P2_U2853) );
  OAI222_X1 U17039 ( .A1(n19796), .A2(n14404), .B1(n14401), .B2(n11533), .C1(
        n14403), .C2(n20045), .ZN(P1_U2897) );
  OR2_X1 U17040 ( .A1(n13827), .A2(n15397), .ZN(n13828) );
  NAND2_X1 U17041 ( .A1(n13829), .A2(n13828), .ZN(n19016) );
  AOI21_X1 U17042 ( .B1(n15366), .B2(n13830), .A(n15364), .ZN(n15399) );
  INV_X1 U17043 ( .A(n15399), .ZN(n13833) );
  OAI22_X1 U17044 ( .A1(n16097), .A2(n13831), .B1(n10551), .B2(n18847), .ZN(
        n13832) );
  AOI21_X1 U17045 ( .B1(n13833), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13832), .ZN(n13838) );
  INV_X1 U17046 ( .A(n13834), .ZN(n13835) );
  NAND2_X1 U17047 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13835), .ZN(
        n13836) );
  NOR2_X1 U17048 ( .A1(n16099), .A2(n13836), .ZN(n15402) );
  NAND2_X1 U17049 ( .A1(n15402), .A2(n15397), .ZN(n13837) );
  OAI211_X1 U17050 ( .C1(n19019), .C2(n15404), .A(n13838), .B(n13837), .ZN(
        n13841) );
  NAND2_X1 U17051 ( .A1(n9735), .A2(n9743), .ZN(n19014) );
  AND3_X1 U17052 ( .A1(n13839), .A2(n16102), .A3(n19014), .ZN(n13840) );
  AOI211_X1 U17053 ( .C1(n16105), .C2(n19016), .A(n13841), .B(n13840), .ZN(
        n13842) );
  INV_X1 U17054 ( .A(n13842), .ZN(P2_U3042) );
  INV_X1 U17055 ( .A(n13843), .ZN(n13847) );
  INV_X1 U17056 ( .A(n13795), .ZN(n13846) );
  INV_X1 U17057 ( .A(n13844), .ZN(n13845) );
  AOI21_X1 U17058 ( .B1(n13847), .B2(n13846), .A(n13845), .ZN(n13885) );
  INV_X1 U17059 ( .A(n13885), .ZN(n13867) );
  INV_X1 U17060 ( .A(n13848), .ZN(n19792) );
  INV_X1 U17061 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n19794) );
  NAND4_X1 U17062 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n19819)
         );
  NAND2_X1 U17063 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19793) );
  NOR3_X1 U17064 ( .A1(n19794), .A2(n19819), .A3(n19793), .ZN(n13858) );
  NAND2_X1 U17065 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n13858), .ZN(n14217) );
  NOR2_X1 U17066 ( .A1(n19792), .A2(n14217), .ZN(n14218) );
  OR2_X1 U17067 ( .A1(n14218), .A2(n15659), .ZN(n19783) );
  INV_X1 U17068 ( .A(n19783), .ZN(n13857) );
  MUX2_X1 U17069 ( .A(n14113), .B(n13551), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n13851) );
  NAND2_X1 U17070 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n14129), .ZN(
        n13849) );
  AND2_X1 U17071 ( .A1(n14097), .A2(n13849), .ZN(n13850) );
  NAND2_X1 U17072 ( .A1(n13851), .A2(n13850), .ZN(n13852) );
  OR2_X1 U17073 ( .A1(n13853), .A2(n13852), .ZN(n13854) );
  NAND2_X1 U17074 ( .A1(n15858), .A2(n13854), .ZN(n15877) );
  AOI22_X1 U17075 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19832), .B1(
        n13881), .B2(n19816), .ZN(n13855) );
  OAI211_X1 U17076 ( .C1(n19835), .C2(n15877), .A(n13855), .B(n19823), .ZN(
        n13856) );
  AOI21_X1 U17077 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n13857), .A(n13856), .ZN(
        n13864) );
  INV_X1 U17078 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13861) );
  INV_X1 U17079 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n13859) );
  NAND2_X1 U17080 ( .A1(n13859), .A2(n13858), .ZN(n13860) );
  OAI22_X1 U17081 ( .A1(n13861), .A2(n19833), .B1(n19820), .B2(n13860), .ZN(
        n13862) );
  INV_X1 U17082 ( .A(n13862), .ZN(n13863) );
  OAI211_X1 U17083 ( .C1(n13867), .C2(n19795), .A(n13864), .B(n13863), .ZN(
        P1_U2832) );
  INV_X1 U17084 ( .A(DATAI_8_), .ZN(n13865) );
  MUX2_X1 U17085 ( .A(n13865), .B(n16260), .S(n20001), .Z(n19888) );
  INV_X1 U17086 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13866) );
  OAI222_X1 U17087 ( .A1(n13867), .A2(n14404), .B1(n19888), .B2(n14403), .C1(
        n13866), .C2(n14401), .ZN(P1_U2896) );
  OAI222_X1 U17088 ( .A1(n13867), .A2(n14322), .B1(n19858), .B2(n13861), .C1(
        n15877), .C2(n14329), .ZN(P1_U2864) );
  OAI21_X1 U17089 ( .B1(n13868), .B2(n13871), .A(n13870), .ZN(n13891) );
  NAND2_X1 U17090 ( .A1(n15233), .A2(n13872), .ZN(n13873) );
  AND2_X1 U17091 ( .A1(n15196), .A2(n13873), .ZN(n18714) );
  OAI22_X1 U17092 ( .A1(n14930), .A2(n18973), .B1(n18953), .B2(n13874), .ZN(
        n13875) );
  AOI21_X1 U17093 ( .B1(n18964), .B2(n18714), .A(n13875), .ZN(n13877) );
  AOI22_X1 U17094 ( .A1(n18910), .A2(BUF2_REG_17__SCAN_IN), .B1(n18911), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n13876) );
  OAI211_X1 U17095 ( .C1(n13891), .C2(n18968), .A(n13877), .B(n13876), .ZN(
        P2_U2902) );
  XOR2_X1 U17096 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n13879), .Z(
        n13880) );
  XNOR2_X1 U17097 ( .A(n13878), .B(n13880), .ZN(n15876) );
  INV_X1 U17098 ( .A(n13881), .ZN(n13883) );
  AOI22_X1 U17099 ( .A1(n19925), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19950), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13882) );
  OAI21_X1 U17100 ( .B1(n19934), .B2(n13883), .A(n13882), .ZN(n13884) );
  AOI21_X1 U17101 ( .B1(n13885), .B2(n19942), .A(n13884), .ZN(n13886) );
  OAI21_X1 U17102 ( .B1(n15876), .B2(n19944), .A(n13886), .ZN(P1_U2991) );
  NAND2_X1 U17103 ( .A1(n14861), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n13890) );
  OR2_X1 U17104 ( .A1(n13930), .A2(n13887), .ZN(n13888) );
  AND2_X1 U17105 ( .A1(n13937), .A2(n13888), .ZN(n18713) );
  NAND2_X1 U17106 ( .A1(n18713), .A2(n14796), .ZN(n13889) );
  OAI211_X1 U17107 ( .C1(n13891), .C2(n14854), .A(n13890), .B(n13889), .ZN(
        P2_U2870) );
  OAI21_X1 U17108 ( .B1(n13892), .B2(n13894), .A(n13893), .ZN(n15726) );
  INV_X1 U17109 ( .A(DATAI_10_), .ZN(n13896) );
  NAND2_X1 U17110 ( .A1(n20001), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13895) );
  OAI21_X1 U17111 ( .B1(n20001), .B2(n13896), .A(n13895), .ZN(n19894) );
  AOI22_X1 U17112 ( .A1(n14397), .A2(n19894), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15744), .ZN(n13897) );
  OAI21_X1 U17113 ( .B1(n15726), .B2(n14404), .A(n13897), .ZN(P1_U2894) );
  INV_X1 U17114 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15724) );
  NAND2_X1 U17115 ( .A1(n14101), .A2(n15724), .ZN(n13902) );
  INV_X1 U17116 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13898) );
  NAND2_X1 U17117 ( .A1(n13551), .A2(n13898), .ZN(n13900) );
  NAND2_X1 U17118 ( .A1(n13266), .A2(n15724), .ZN(n13899) );
  NAND3_X1 U17119 ( .A1(n13900), .A2(n14089), .A3(n13899), .ZN(n13901) );
  INV_X1 U17120 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n19847) );
  NAND2_X1 U17121 ( .A1(n13266), .A2(n19847), .ZN(n13904) );
  NAND2_X1 U17122 ( .A1(n14089), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13903) );
  NAND3_X1 U17123 ( .A1(n13904), .A2(n13551), .A3(n13903), .ZN(n13905) );
  OAI21_X1 U17124 ( .B1(n14107), .B2(P1_EBX_REG_9__SCAN_IN), .A(n13905), .ZN(
        n15857) );
  INV_X1 U17125 ( .A(n14324), .ZN(n13906) );
  AOI21_X1 U17126 ( .B1(n13907), .B2(n15860), .A(n13906), .ZN(n15849) );
  AOI22_X1 U17127 ( .A1(n15849), .A2(n19853), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14303), .ZN(n13908) );
  OAI21_X1 U17128 ( .B1(n15726), .B2(n14322), .A(n13908), .ZN(P1_U2862) );
  NOR2_X1 U17129 ( .A1(n13845), .A2(n13909), .ZN(n13910) );
  OR2_X1 U17130 ( .A1(n13892), .A2(n13910), .ZN(n19844) );
  INV_X1 U17131 ( .A(DATAI_9_), .ZN(n13912) );
  MUX2_X1 U17132 ( .A(n13912), .B(n13911), .S(n20001), .Z(n19891) );
  INV_X1 U17133 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n13913) );
  OAI222_X1 U17134 ( .A1(n19844), .A2(n14404), .B1(n19891), .B2(n14403), .C1(
        n13913), .C2(n14401), .ZN(P1_U2895) );
  OAI21_X1 U17135 ( .B1(n13917), .B2(n13915), .A(n13914), .ZN(n13916) );
  OAI21_X1 U17136 ( .B1(n13918), .B2(n13920), .A(n13919), .ZN(n15406) );
  NOR2_X1 U17137 ( .A1(n15406), .A2(n16072), .ZN(n13925) );
  NOR2_X1 U17138 ( .A1(n18850), .A2(n19020), .ZN(n13924) );
  OAI22_X1 U17139 ( .A1(n16059), .A2(n13921), .B1(n10328), .B2(n18847), .ZN(
        n13923) );
  AND2_X1 U17140 ( .A1(n16052), .A2(n18843), .ZN(n13922) );
  NOR4_X1 U17141 ( .A1(n13925), .A2(n13924), .A3(n13923), .A4(n13922), .ZN(
        n13926) );
  OAI21_X1 U17142 ( .B1(n16073), .B2(n15412), .A(n13926), .ZN(P2_U3009) );
  NOR2_X1 U17143 ( .A1(n13785), .A2(n13927), .ZN(n13928) );
  OR2_X1 U17144 ( .A1(n13868), .A2(n13928), .ZN(n18914) );
  AND2_X1 U17145 ( .A1(n9728), .A2(n13929), .ZN(n13931) );
  OR2_X1 U17146 ( .A1(n13931), .A2(n13930), .ZN(n18727) );
  NOR2_X1 U17147 ( .A1(n18727), .A2(n13122), .ZN(n13932) );
  AOI21_X1 U17148 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n13122), .A(n13932), .ZN(
        n13933) );
  OAI21_X1 U17149 ( .B1(n18914), .B2(n14854), .A(n13933), .ZN(P2_U2871) );
  INV_X1 U17150 ( .A(n13934), .ZN(n13935) );
  AOI21_X1 U17151 ( .B1(n13936), .B2(n13870), .A(n13935), .ZN(n15991) );
  NAND2_X1 U17152 ( .A1(n15991), .A2(n14860), .ZN(n13940) );
  AOI21_X1 U17153 ( .B1(n13938), .B2(n13937), .A(n10364), .ZN(n18701) );
  NAND2_X1 U17154 ( .A1(n18701), .A2(n14796), .ZN(n13939) );
  OAI211_X1 U17155 ( .C1(n14796), .C2(n13941), .A(n13940), .B(n13939), .ZN(
        P2_U2869) );
  MUX2_X1 U17156 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n11999), .S(
        n15785), .Z(n13942) );
  XNOR2_X1 U17157 ( .A(n13943), .B(n13942), .ZN(n15864) );
  NAND2_X1 U17158 ( .A1(n15864), .A2(n19930), .ZN(n13946) );
  NAND2_X1 U17159 ( .A1(n19950), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n15861) );
  OAI21_X1 U17160 ( .B1(n19938), .B2(n19780), .A(n15861), .ZN(n13944) );
  AOI21_X1 U17161 ( .B1(n15781), .B2(n19779), .A(n13944), .ZN(n13945) );
  OAI211_X1 U17162 ( .C1(n20003), .C2(n19844), .A(n13946), .B(n13945), .ZN(
        P1_U2990) );
  INV_X1 U17163 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n13949) );
  INV_X1 U17164 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16587) );
  INV_X1 U17165 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n16610) );
  INV_X1 U17166 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n16975) );
  INV_X1 U17167 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n16671) );
  NOR3_X1 U17168 ( .A1(n17092), .A2(n18003), .A3(n13947), .ZN(n13948) );
  NOR4_X4 U17169 ( .A1(n18631), .A2(n16646), .A3(n15591), .A4(n18490), .ZN(
        n16994) );
  NAND3_X1 U17170 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(n16994), .ZN(n16987) );
  NOR2_X2 U17171 ( .A1(n16671), .A2(n16987), .ZN(n16984) );
  AND2_X2 U17172 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16979), .ZN(n16983) );
  NAND2_X2 U17173 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n16983), .ZN(n16972) );
  NOR3_X4 U17174 ( .A1(n16610), .A2(n16975), .A3(n16972), .ZN(n16971) );
  NOR2_X4 U17175 ( .A1(n16587), .A2(n16966), .ZN(n16922) );
  INV_X1 U17176 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16563) );
  INV_X1 U17177 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n16921) );
  NOR2_X1 U17178 ( .A1(n16563), .A2(n16921), .ZN(n13950) );
  INV_X1 U17179 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n16550) );
  NAND3_X1 U17180 ( .A1(n18024), .A2(n16922), .A3(n13950), .ZN(n16882) );
  NOR2_X1 U17181 ( .A1(n16550), .A2(n16882), .ZN(n16895) );
  AOI21_X1 U17182 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n16895), .A(
        P3_EBX_REG_14__SCAN_IN), .ZN(n13951) );
  NOR2_X1 U17183 ( .A1(n16880), .A2(n13951), .ZN(n13963) );
  AOI22_X1 U17184 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13955) );
  AOI22_X1 U17185 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13954) );
  AOI22_X1 U17186 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13953) );
  AOI22_X1 U17187 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13952) );
  NAND4_X1 U17188 ( .A1(n13955), .A2(n13954), .A3(n13953), .A4(n13952), .ZN(
        n13961) );
  AOI22_X1 U17189 ( .A1(n16883), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13959) );
  AOI22_X1 U17190 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13958) );
  AOI22_X1 U17191 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13957) );
  AOI22_X1 U17192 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13956) );
  NAND4_X1 U17193 ( .A1(n13959), .A2(n13958), .A3(n13957), .A4(n13956), .ZN(
        n13960) );
  NOR2_X1 U17194 ( .A1(n13961), .A2(n13960), .ZN(n17098) );
  INV_X1 U17195 ( .A(n17098), .ZN(n13962) );
  INV_X1 U17196 ( .A(n16994), .ZN(n16997) );
  MUX2_X1 U17197 ( .A(n13963), .B(n13962), .S(n16998), .Z(P3_U2689) );
  INV_X1 U17198 ( .A(n18419), .ZN(n13967) );
  OAI21_X1 U17199 ( .B1(n13978), .B2(n18604), .A(n18478), .ZN(n13966) );
  NAND2_X1 U17200 ( .A1(n13967), .A2(n13966), .ZN(n18430) );
  NOR2_X1 U17201 ( .A1(n18593), .A2(n18430), .ZN(n13976) );
  INV_X1 U17202 ( .A(n17224), .ZN(n13970) );
  NOR2_X1 U17203 ( .A1(n17991), .A2(n13970), .ZN(n18475) );
  OAI21_X1 U17204 ( .B1(n13969), .B2(n18475), .A(n13968), .ZN(n17163) );
  NAND2_X1 U17205 ( .A1(n16317), .A2(n18632), .ZN(n13974) );
  AOI221_X2 U17206 ( .B1(n18631), .B2(n18419), .C1(n13970), .C2(n18419), .A(
        n13974), .ZN(n15593) );
  AOI21_X1 U17207 ( .B1(n18428), .B2(n13971), .A(n15593), .ZN(n13972) );
  OAI211_X1 U17208 ( .C1(n17163), .C2(n13974), .A(n13973), .B(n13972), .ZN(
        n18450) );
  NOR2_X1 U17209 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18586), .ZN(n17987) );
  INV_X1 U17210 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n17972) );
  NAND2_X1 U17211 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18626), .ZN(n18584) );
  NOR2_X1 U17212 ( .A1(n17972), .A2(n18584), .ZN(n13975) );
  AOI211_X1 U17213 ( .C1(n18483), .C2(n18450), .A(n17987), .B(n13975), .ZN(
        n18613) );
  MUX2_X1 U17214 ( .A(n13976), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18613), .Z(P3_U3284) );
  OAI211_X1 U17215 ( .C1(n13978), .C2(n18604), .A(n13977), .B(n18478), .ZN(
        n17971) );
  NOR2_X1 U17216 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n17971), .ZN(n13979) );
  OAI21_X1 U17217 ( .B1(n13979), .B2(n18584), .A(n18178), .ZN(n17982) );
  INV_X1 U17218 ( .A(n17982), .ZN(n13980) );
  NOR2_X1 U17219 ( .A1(n18625), .A2(n17541), .ZN(n17975) );
  AOI21_X1 U17220 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n17975), .ZN(n17976) );
  NOR2_X1 U17221 ( .A1(n13980), .A2(n17976), .ZN(n13982) );
  INV_X1 U17222 ( .A(n18324), .ZN(n17977) );
  NOR2_X1 U17223 ( .A1(n18586), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18028) );
  OR2_X1 U17224 ( .A1(n18028), .A2(n13980), .ZN(n17974) );
  OR2_X1 U17225 ( .A1(n17977), .A2(n17974), .ZN(n13981) );
  MUX2_X1 U17226 ( .A(n13982), .B(n13981), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  AOI22_X1 U17227 ( .A1(n20660), .A2(n13984), .B1(n13983), .B2(n15547), .ZN(
        n15545) );
  OAI21_X1 U17228 ( .B1(n15545), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20577), 
        .ZN(n13985) );
  AOI22_X1 U17229 ( .A1(n20649), .A2(n15547), .B1(n13986), .B2(n13985), .ZN(
        n13989) );
  AOI21_X1 U17230 ( .B1(n13987), .B2(n15908), .A(n15906), .ZN(n13988) );
  OAI22_X1 U17231 ( .A1(n13989), .A2(n15906), .B1(n13988), .B2(n15547), .ZN(
        P1_U3474) );
  OAI21_X1 U17232 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n13993), .ZN(n13991) );
  NAND2_X1 U17233 ( .A1(n13992), .A2(n13991), .ZN(n13996) );
  INV_X1 U17234 ( .A(n13993), .ZN(n13994) );
  INV_X1 U17235 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15096) );
  OAI21_X1 U17236 ( .B1(n13999), .B2(n14002), .A(n15096), .ZN(n14936) );
  NAND2_X1 U17237 ( .A1(n14035), .A2(n14935), .ZN(n14005) );
  AOI21_X1 U17238 ( .B1(n14001), .B2(n14000), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14034) );
  NOR2_X1 U17239 ( .A1(n14034), .A2(n9708), .ZN(n14004) );
  XNOR2_X1 U17240 ( .A(n14005), .B(n14004), .ZN(n15090) );
  XNOR2_X1 U17241 ( .A(n14939), .B(n14006), .ZN(n15088) );
  NOR2_X1 U17242 ( .A1(n18847), .A2(n14007), .ZN(n15084) );
  NOR2_X1 U17243 ( .A1(n19025), .A2(n14008), .ZN(n14009) );
  AOI211_X1 U17244 ( .C1(n19012), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15084), .B(n14009), .ZN(n14010) );
  OAI21_X1 U17245 ( .B1(n15087), .B2(n19020), .A(n14010), .ZN(n14011) );
  AOI21_X1 U17246 ( .B1(n15088), .B2(n19015), .A(n14011), .ZN(n14012) );
  OAI21_X1 U17247 ( .B1(n15090), .B2(n16072), .A(n14012), .ZN(P2_U2984) );
  INV_X1 U17248 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14608) );
  AND2_X1 U17249 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14541) );
  NAND2_X1 U17250 ( .A1(n14430), .A2(n14589), .ZN(n14584) );
  NAND2_X1 U17251 ( .A1(n14016), .A2(n14428), .ZN(n14017) );
  NAND2_X1 U17252 ( .A1(n14017), .A2(n9590), .ZN(n14018) );
  OR2_X1 U17253 ( .A1(n15785), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14420) );
  NAND2_X1 U17254 ( .A1(n14479), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14419) );
  NAND2_X1 U17255 ( .A1(n19950), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14560) );
  NAND2_X1 U17256 ( .A1(n19925), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14020) );
  OAI211_X1 U17257 ( .C1(n19934), .C2(n14021), .A(n14560), .B(n14020), .ZN(
        n14022) );
  OAI21_X1 U17258 ( .B1(n14565), .B2(n19944), .A(n14023), .ZN(P1_U2968) );
  INV_X1 U17259 ( .A(n14027), .ZN(n14865) );
  NAND2_X1 U17260 ( .A1(n14029), .A2(n14028), .ZN(n14864) );
  NAND3_X1 U17261 ( .A1(n14865), .A2(n14860), .A3(n14864), .ZN(n14031) );
  NAND2_X1 U17262 ( .A1(n13122), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14030) );
  OAI211_X1 U17263 ( .C1(n14861), .C2(n15930), .A(n14031), .B(n14030), .ZN(
        P2_U2858) );
  NOR2_X1 U17264 ( .A1(n9708), .A2(n14032), .ZN(n14033) );
  XNOR2_X1 U17265 ( .A(n14036), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14037) );
  XNOR2_X1 U17266 ( .A(n14038), .B(n14037), .ZN(n14057) );
  XNOR2_X1 U17267 ( .A(n14039), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14055) );
  NAND3_X1 U17268 ( .A1(n15094), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15081) );
  NOR3_X1 U17269 ( .A1(n15081), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14006), .ZN(n14041) );
  NAND2_X1 U17270 ( .A1(n19011), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14050) );
  INV_X1 U17271 ( .A(n14050), .ZN(n14040) );
  OR2_X1 U17272 ( .A1(n14041), .A2(n14040), .ZN(n14044) );
  NOR3_X1 U17273 ( .A1(n15096), .A2(n20693), .A3(n14948), .ZN(n14043) );
  OAI211_X1 U17274 ( .C1(n15367), .C2(n14043), .A(n14042), .B(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15082) );
  AOI21_X1 U17275 ( .B1(n14055), .B2(n16105), .A(n14047), .ZN(n14048) );
  OAI21_X1 U17276 ( .B1(n14057), .B2(n15405), .A(n14048), .ZN(P2_U3015) );
  NAND2_X1 U17277 ( .A1(n19012), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14049) );
  OAI211_X1 U17278 ( .C1(n19025), .C2(n14051), .A(n14050), .B(n14049), .ZN(
        n14052) );
  INV_X1 U17279 ( .A(n14052), .ZN(n14053) );
  AOI21_X1 U17280 ( .B1(n14055), .B2(n19015), .A(n14054), .ZN(n14056) );
  OAI21_X1 U17281 ( .B1(n14057), .B2(n16072), .A(n14056), .ZN(P2_U2983) );
  XNOR2_X1 U17282 ( .A(n14152), .B(n14059), .ZN(n14416) );
  INV_X1 U17283 ( .A(n14416), .ZN(n14123) );
  INV_X1 U17284 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14122) );
  MUX2_X1 U17285 ( .A(n14107), .B(n14089), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n14062) );
  INV_X1 U17286 ( .A(n14130), .ZN(n14060) );
  INV_X1 U17287 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14535) );
  NAND2_X1 U17288 ( .A1(n14060), .A2(n14535), .ZN(n14061) );
  NAND2_X1 U17289 ( .A1(n14062), .A2(n14061), .ZN(n14323) );
  MUX2_X1 U17290 ( .A(n14113), .B(n13551), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n14065) );
  NAND2_X1 U17291 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14129), .ZN(
        n14063) );
  AND2_X1 U17292 ( .A1(n14097), .A2(n14063), .ZN(n14064) );
  NAND2_X1 U17293 ( .A1(n14065), .A2(n14064), .ZN(n14318) );
  MUX2_X1 U17294 ( .A(n14107), .B(n14089), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n14066) );
  OAI21_X1 U17295 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n14130), .A(
        n14066), .ZN(n14067) );
  INV_X1 U17296 ( .A(n14067), .ZN(n14312) );
  INV_X1 U17297 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n20836) );
  NAND2_X1 U17298 ( .A1(n14101), .A2(n20836), .ZN(n14072) );
  NAND2_X1 U17299 ( .A1(n13551), .A2(n14068), .ZN(n14070) );
  NAND2_X1 U17300 ( .A1(n13266), .A2(n20836), .ZN(n14069) );
  NAND3_X1 U17301 ( .A1(n14070), .A2(n14089), .A3(n14069), .ZN(n14071) );
  AND2_X1 U17302 ( .A1(n14072), .A2(n14071), .ZN(n14220) );
  MUX2_X1 U17303 ( .A(n14107), .B(n14089), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n14073) );
  NAND2_X1 U17304 ( .A1(n14073), .A2(n10076), .ZN(n14299) );
  NAND2_X1 U17305 ( .A1(n13551), .A2(n14694), .ZN(n14075) );
  INV_X1 U17306 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n20755) );
  NAND2_X1 U17307 ( .A1(n13266), .A2(n20755), .ZN(n14074) );
  NAND3_X1 U17308 ( .A1(n14075), .A2(n14089), .A3(n14074), .ZN(n14076) );
  OAI21_X1 U17309 ( .B1(n14113), .B2(P1_EBX_REG_16__SCAN_IN), .A(n14076), .ZN(
        n14292) );
  MUX2_X1 U17310 ( .A(n14107), .B(n14089), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n14077) );
  OAI21_X1 U17311 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n14130), .A(
        n14077), .ZN(n14078) );
  INV_X1 U17312 ( .A(n14078), .ZN(n14282) );
  INV_X1 U17313 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n20798) );
  NAND2_X1 U17314 ( .A1(n14101), .A2(n20798), .ZN(n14082) );
  NAND2_X1 U17315 ( .A1(n13551), .A2(n15820), .ZN(n14080) );
  NAND2_X1 U17316 ( .A1(n13266), .A2(n20798), .ZN(n14079) );
  NAND3_X1 U17317 ( .A1(n14080), .A2(n14089), .A3(n14079), .ZN(n14081) );
  AND2_X1 U17318 ( .A1(n14082), .A2(n14081), .ZN(n14277) );
  MUX2_X1 U17319 ( .A(n14107), .B(n14089), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n14083) );
  NAND2_X1 U17320 ( .A1(n14083), .A2(n10083), .ZN(n14268) );
  MUX2_X1 U17321 ( .A(n14113), .B(n13551), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n14086) );
  NAND2_X1 U17322 ( .A1(n14129), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14084) );
  AND2_X1 U17323 ( .A1(n14097), .A2(n14084), .ZN(n14085) );
  NAND2_X1 U17324 ( .A1(n14086), .A2(n14085), .ZN(n14266) );
  MUX2_X1 U17325 ( .A(n14107), .B(n14089), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n14087) );
  OAI21_X1 U17326 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n14130), .A(
        n14087), .ZN(n14259) );
  INV_X1 U17327 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15616) );
  NAND2_X1 U17328 ( .A1(n14101), .A2(n15616), .ZN(n14092) );
  INV_X1 U17329 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14657) );
  NAND2_X1 U17330 ( .A1(n13551), .A2(n14657), .ZN(n14090) );
  NAND2_X1 U17331 ( .A1(n13266), .A2(n15616), .ZN(n14088) );
  NAND3_X1 U17332 ( .A1(n14090), .A2(n14089), .A3(n14088), .ZN(n14091) );
  AND2_X1 U17333 ( .A1(n14092), .A2(n14091), .ZN(n14252) );
  INV_X1 U17334 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n20738) );
  NAND2_X1 U17335 ( .A1(n13266), .A2(n20738), .ZN(n14094) );
  NAND2_X1 U17336 ( .A1(n14089), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14093) );
  NAND3_X1 U17337 ( .A1(n14094), .A2(n13551), .A3(n14093), .ZN(n14095) );
  OAI21_X1 U17338 ( .B1(n14107), .B2(P1_EBX_REG_23__SCAN_IN), .A(n14095), .ZN(
        n14635) );
  MUX2_X1 U17339 ( .A(n14113), .B(n13551), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n14099) );
  NAND2_X1 U17340 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n14129), .ZN(
        n14096) );
  AND2_X1 U17341 ( .A1(n14097), .A2(n14096), .ZN(n14098) );
  NAND2_X1 U17342 ( .A1(n14099), .A2(n14098), .ZN(n14244) );
  MUX2_X1 U17343 ( .A(n14107), .B(n14089), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n14100) );
  OAI21_X1 U17344 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n14130), .A(
        n14100), .ZN(n14202) );
  INV_X1 U17345 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14102) );
  NAND2_X1 U17346 ( .A1(n14101), .A2(n14102), .ZN(n14106) );
  NAND2_X1 U17347 ( .A1(n13551), .A2(n14608), .ZN(n14104) );
  NAND2_X1 U17348 ( .A1(n13266), .A2(n14102), .ZN(n14103) );
  NAND3_X1 U17349 ( .A1(n14104), .A2(n14089), .A3(n14103), .ZN(n14105) );
  AND2_X1 U17350 ( .A1(n14106), .A2(n14105), .ZN(n14190) );
  MUX2_X1 U17351 ( .A(n14107), .B(n14089), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n14108) );
  OAI21_X1 U17352 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14130), .A(
        n14108), .ZN(n14109) );
  INV_X1 U17353 ( .A(n14109), .ZN(n14177) );
  NAND2_X1 U17354 ( .A1(n13551), .A2(n14589), .ZN(n14111) );
  INV_X1 U17355 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14234) );
  NAND2_X1 U17356 ( .A1(n13266), .A2(n14234), .ZN(n14110) );
  NAND3_X1 U17357 ( .A1(n14111), .A2(n14089), .A3(n14110), .ZN(n14112) );
  OAI21_X1 U17358 ( .B1(n14113), .B2(P1_EBX_REG_28__SCAN_IN), .A(n14112), .ZN(
        n14163) );
  INV_X1 U17359 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14114) );
  NAND2_X1 U17360 ( .A1(n13266), .A2(n14114), .ZN(n14116) );
  OR2_X1 U17361 ( .A1(n14130), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14115) );
  NAND2_X1 U17362 ( .A1(n14115), .A2(n14116), .ZN(n14118) );
  MUX2_X1 U17363 ( .A(n14116), .B(n14118), .S(n14089), .Z(n14160) );
  OAI22_X1 U17364 ( .A1(n14159), .A2(n14089), .B1(n14118), .B2(n14117), .ZN(
        n14121) );
  NAND2_X1 U17365 ( .A1(n14130), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n14120) );
  NAND2_X1 U17366 ( .A1(n14129), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14119) );
  NAND2_X1 U17367 ( .A1(n14120), .A2(n14119), .ZN(n14127) );
  XNOR2_X1 U17368 ( .A(n14121), .B(n14127), .ZN(n14571) );
  OAI222_X1 U17369 ( .A1(n14322), .A2(n14123), .B1(n14122), .B2(n19858), .C1(
        n14571), .C2(n14329), .ZN(P1_U2842) );
  NOR2_X1 U17370 ( .A1(n15087), .A2(n13122), .ZN(n14124) );
  AOI21_X1 U17371 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n14861), .A(n14124), .ZN(
        n14125) );
  OAI21_X1 U17372 ( .B1(n14126), .B2(n14854), .A(n14125), .ZN(P2_U2857) );
  AOI22_X1 U17373 ( .A1(n14130), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n14129), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14131) );
  NAND2_X1 U17374 ( .A1(n14132), .A2(n19811), .ZN(n14143) );
  NAND2_X1 U17375 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14139) );
  INV_X1 U17376 ( .A(n14139), .ZN(n14136) );
  INV_X1 U17377 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20619) );
  INV_X1 U17378 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n14219) );
  INV_X1 U17379 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20615) );
  NAND4_X1 U17380 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(P1_REIP_REG_11__SCAN_IN), .ZN(n15697) );
  OR3_X1 U17381 ( .A1(n14219), .A2(n20615), .A3(n15697), .ZN(n15671) );
  INV_X1 U17382 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20620) );
  INV_X1 U17383 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n15831) );
  NOR4_X1 U17384 ( .A1(n20619), .A2(n15671), .A3(n20620), .A4(n15831), .ZN(
        n15658) );
  INV_X1 U17385 ( .A(n15658), .ZN(n14133) );
  NAND2_X1 U17386 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n15650) );
  NOR3_X1 U17387 ( .A1(n14217), .A2(n14133), .A3(n15650), .ZN(n15613) );
  INV_X1 U17388 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20628) );
  NAND2_X1 U17389 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15621) );
  NOR2_X1 U17390 ( .A1(n20628), .A2(n15621), .ZN(n15609) );
  NAND3_X1 U17391 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n15613), .A3(n15609), 
        .ZN(n15596) );
  NOR2_X1 U17392 ( .A1(n19792), .A2(n15596), .ZN(n15602) );
  AND2_X1 U17393 ( .A1(n15602), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14205) );
  NAND2_X1 U17394 ( .A1(n14194), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14180) );
  NAND2_X1 U17395 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14134) );
  NOR2_X1 U17396 ( .A1(n14180), .A2(n14134), .ZN(n14138) );
  INV_X1 U17397 ( .A(n14138), .ZN(n14135) );
  NAND2_X1 U17398 ( .A1(n14135), .A2(n19806), .ZN(n14167) );
  OAI21_X1 U17399 ( .B1(n15659), .B2(n14136), .A(n14167), .ZN(n14148) );
  INV_X1 U17400 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14137) );
  INV_X1 U17401 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14230) );
  OAI22_X1 U17402 ( .A1(n19791), .A2(n14137), .B1(n14230), .B2(n19833), .ZN(
        n14141) );
  INV_X1 U17403 ( .A(n19820), .ZN(n15615) );
  NAND2_X1 U17404 ( .A1(n14138), .A2(n15615), .ZN(n14155) );
  NOR3_X1 U17405 ( .A1(n14155), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14139), 
        .ZN(n14140) );
  AOI211_X1 U17406 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14148), .A(n14141), 
        .B(n14140), .ZN(n14142) );
  OAI211_X1 U17407 ( .C1(n14231), .C2(n19835), .A(n14143), .B(n14142), .ZN(
        P1_U2809) );
  NAND2_X1 U17408 ( .A1(n14416), .A2(n19811), .ZN(n14151) );
  INV_X1 U17409 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14422) );
  INV_X1 U17410 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14144) );
  OAI21_X1 U17411 ( .B1(n14155), .B2(n14422), .A(n14144), .ZN(n14149) );
  INV_X1 U17412 ( .A(n14412), .ZN(n14146) );
  AOI22_X1 U17413 ( .A1(n19832), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n19818), .ZN(n14145) );
  OAI21_X1 U17414 ( .B1(n19828), .B2(n14146), .A(n14145), .ZN(n14147) );
  AOI21_X1 U17415 ( .B1(n14149), .B2(n14148), .A(n14147), .ZN(n14150) );
  OAI211_X1 U17416 ( .C1(n19835), .C2(n14571), .A(n14151), .B(n14150), .ZN(
        P1_U2810) );
  AOI21_X1 U17417 ( .B1(n14153), .B2(n12126), .A(n14152), .ZN(n14426) );
  INV_X1 U17418 ( .A(n14426), .ZN(n14233) );
  INV_X1 U17419 ( .A(n14167), .ZN(n14158) );
  AOI22_X1 U17420 ( .A1(n19832), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        n19818), .B2(P1_EBX_REG_29__SCAN_IN), .ZN(n14154) );
  OAI21_X1 U17421 ( .B1(n19828), .B2(n14424), .A(n14154), .ZN(n14157) );
  NOR2_X1 U17422 ( .A1(n14155), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14156) );
  AOI211_X1 U17423 ( .C1(n14158), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14157), 
        .B(n14156), .ZN(n14162) );
  AOI21_X1 U17424 ( .B1(n14160), .B2(n14117), .A(n14159), .ZN(n14579) );
  NAND2_X1 U17425 ( .A1(n14579), .A2(n19815), .ZN(n14161) );
  OAI211_X1 U17426 ( .C1(n14233), .C2(n19795), .A(n14162), .B(n14161), .ZN(
        P1_U2811) );
  OR2_X1 U17427 ( .A1(n14179), .A2(n14163), .ZN(n14164) );
  NAND2_X1 U17428 ( .A1(n14117), .A2(n14164), .ZN(n14583) );
  INV_X1 U17429 ( .A(n14235), .ZN(n14343) );
  NAND2_X1 U17430 ( .A1(n14343), .A2(n19811), .ZN(n14174) );
  OAI22_X1 U17431 ( .A1(n19791), .A2(n14165), .B1(n19833), .B2(n14234), .ZN(
        n14171) );
  INV_X1 U17432 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14169) );
  INV_X1 U17433 ( .A(n14180), .ZN(n14166) );
  NAND2_X1 U17434 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n14166), .ZN(n14168) );
  AOI21_X1 U17435 ( .B1(n14169), .B2(n14168), .A(n14167), .ZN(n14170) );
  AOI211_X1 U17436 ( .C1(n19816), .C2(n14172), .A(n14171), .B(n14170), .ZN(
        n14173) );
  OAI211_X1 U17437 ( .C1(n19835), .C2(n14583), .A(n14174), .B(n14173), .ZN(
        P1_U2812) );
  AOI21_X1 U17438 ( .B1(n14176), .B2(n14175), .A(n11927), .ZN(n14435) );
  INV_X1 U17439 ( .A(n14435), .ZN(n14238) );
  NOR2_X1 U17440 ( .A1(n14192), .A2(n14177), .ZN(n14178) );
  OR2_X1 U17441 ( .A1(n14179), .A2(n14178), .ZN(n14236) );
  INV_X1 U17442 ( .A(n14236), .ZN(n14600) );
  NOR3_X1 U17443 ( .A1(n14180), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n19820), 
        .ZN(n14185) );
  NAND3_X1 U17444 ( .A1(n14180), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n19806), 
        .ZN(n14183) );
  INV_X1 U17445 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14237) );
  NOR2_X1 U17446 ( .A1(n19833), .A2(n14237), .ZN(n14181) );
  AOI21_X1 U17447 ( .B1(n19832), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14181), .ZN(n14182) );
  OAI211_X1 U17448 ( .C1(n19828), .C2(n14433), .A(n14183), .B(n14182), .ZN(
        n14184) );
  AOI211_X1 U17449 ( .C1(n14600), .C2(n19815), .A(n14185), .B(n14184), .ZN(
        n14186) );
  OAI21_X1 U17450 ( .B1(n14238), .B2(n19795), .A(n14186), .ZN(P1_U2813) );
  OAI21_X1 U17451 ( .B1(n14188), .B2(n14189), .A(n14175), .ZN(n14441) );
  AND2_X1 U17452 ( .A1(n14204), .A2(n14190), .ZN(n14191) );
  NOR2_X1 U17453 ( .A1(n14192), .A2(n14191), .ZN(n14614) );
  NOR2_X1 U17454 ( .A1(n14194), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14193) );
  AOI211_X1 U17455 ( .C1(n14194), .C2(P1_REIP_REG_26__SCAN_IN), .A(n15659), 
        .B(n14193), .ZN(n14198) );
  INV_X1 U17456 ( .A(n14444), .ZN(n14196) );
  AOI22_X1 U17457 ( .A1(n19832), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n19818), .B2(P1_EBX_REG_26__SCAN_IN), .ZN(n14195) );
  OAI21_X1 U17458 ( .B1(n19828), .B2(n14196), .A(n14195), .ZN(n14197) );
  AOI211_X1 U17459 ( .C1(n14614), .C2(n19815), .A(n14198), .B(n14197), .ZN(
        n14199) );
  OAI21_X1 U17460 ( .B1(n14441), .B2(n19795), .A(n14199), .ZN(P1_U2814) );
  AOI21_X1 U17461 ( .B1(n14201), .B2(n14200), .A(n14188), .ZN(n14454) );
  INV_X1 U17462 ( .A(n14454), .ZN(n14241) );
  NAND2_X1 U17463 ( .A1(n14246), .A2(n14202), .ZN(n14203) );
  NAND2_X1 U17464 ( .A1(n14204), .A2(n14203), .ZN(n14622) );
  INV_X1 U17465 ( .A(n14622), .ZN(n14212) );
  INV_X1 U17466 ( .A(n14205), .ZN(n14206) );
  NOR3_X1 U17467 ( .A1(n14206), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n19820), 
        .ZN(n14211) );
  NAND3_X1 U17468 ( .A1(n14206), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n19806), 
        .ZN(n14209) );
  INV_X1 U17469 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14240) );
  NOR2_X1 U17470 ( .A1(n19833), .A2(n14240), .ZN(n14207) );
  AOI21_X1 U17471 ( .B1(n19832), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14207), .ZN(n14208) );
  OAI211_X1 U17472 ( .C1(n19828), .C2(n14452), .A(n14209), .B(n14208), .ZN(
        n14210) );
  AOI211_X1 U17473 ( .C1(n14212), .C2(n19815), .A(n14211), .B(n14210), .ZN(
        n14213) );
  OAI21_X1 U17474 ( .B1(n14241), .B2(n19795), .A(n14213), .ZN(P1_U2815) );
  OAI21_X1 U17475 ( .B1(n14214), .B2(n14216), .A(n14215), .ZN(n14516) );
  INV_X1 U17476 ( .A(n14516), .ZN(n14228) );
  NAND2_X1 U17477 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n15716) );
  INV_X1 U17478 ( .A(n15730), .ZN(n19781) );
  NOR2_X1 U17479 ( .A1(n15716), .A2(n19781), .ZN(n15721) );
  NAND3_X1 U17480 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(n15721), .ZN(n15707) );
  INV_X1 U17481 ( .A(n14218), .ZN(n15715) );
  OAI21_X1 U17482 ( .B1(n15671), .B2(n15715), .A(n19806), .ZN(n15696) );
  AOI221_X1 U17483 ( .B1(n20615), .B2(n14219), .C1(n15707), .C2(n14219), .A(
        n15696), .ZN(n14227) );
  NAND2_X1 U17484 ( .A1(n14314), .A2(n14220), .ZN(n14221) );
  NAND2_X1 U17485 ( .A1(n14300), .A2(n14221), .ZN(n14710) );
  OAI21_X1 U17486 ( .B1(n19833), .B2(n20836), .A(n19823), .ZN(n14222) );
  AOI21_X1 U17487 ( .B1(n19832), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n14222), .ZN(n14225) );
  INV_X1 U17488 ( .A(n14511), .ZN(n14223) );
  NAND2_X1 U17489 ( .A1(n19816), .A2(n14223), .ZN(n14224) );
  OAI211_X1 U17490 ( .C1(n14710), .C2(n19835), .A(n14225), .B(n14224), .ZN(
        n14226) );
  AOI211_X1 U17491 ( .C1(n14228), .C2(n19811), .A(n14227), .B(n14226), .ZN(
        n14229) );
  INV_X1 U17492 ( .A(n14229), .ZN(P1_U2826) );
  OAI22_X1 U17493 ( .A1(n14231), .A2(n14329), .B1(n19858), .B2(n14230), .ZN(
        P1_U2841) );
  AOI22_X1 U17494 ( .A1(n14579), .A2(n19853), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14303), .ZN(n14232) );
  OAI21_X1 U17495 ( .B1(n14233), .B2(n14322), .A(n14232), .ZN(P1_U2843) );
  OAI222_X1 U17496 ( .A1(n14322), .A2(n14235), .B1(n14234), .B2(n19858), .C1(
        n14583), .C2(n14329), .ZN(P1_U2844) );
  OAI222_X1 U17497 ( .A1(n14322), .A2(n14238), .B1(n14237), .B2(n19858), .C1(
        n14236), .C2(n14329), .ZN(P1_U2845) );
  AOI22_X1 U17498 ( .A1(n14614), .A2(n19853), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n14303), .ZN(n14239) );
  OAI21_X1 U17499 ( .B1(n14441), .B2(n14322), .A(n14239), .ZN(P1_U2846) );
  OAI222_X1 U17500 ( .A1(n14322), .A2(n14241), .B1(n14240), .B2(n19858), .C1(
        n14622), .C2(n14329), .ZN(P1_U2847) );
  NAND2_X1 U17501 ( .A1(n9716), .A2(n14242), .ZN(n14243) );
  AND2_X1 U17502 ( .A1(n14200), .A2(n14243), .ZN(n15603) );
  INV_X1 U17503 ( .A(n15603), .ZN(n14247) );
  INV_X1 U17504 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n15597) );
  OR2_X1 U17505 ( .A1(n14638), .A2(n14244), .ZN(n14245) );
  NAND2_X1 U17506 ( .A1(n14246), .A2(n14245), .ZN(n15606) );
  OAI222_X1 U17507 ( .A1(n14322), .A2(n14247), .B1(n19858), .B2(n15597), .C1(
        n15606), .C2(n14329), .ZN(P1_U2848) );
  OR2_X1 U17508 ( .A1(n14249), .A2(n14250), .ZN(n14251) );
  AND2_X1 U17509 ( .A1(n14248), .A2(n14251), .ZN(n15623) );
  INV_X1 U17510 ( .A(n14322), .ZN(n19854) );
  NAND2_X1 U17511 ( .A1(n14261), .A2(n14252), .ZN(n14253) );
  NAND2_X1 U17512 ( .A1(n14636), .A2(n14253), .ZN(n15626) );
  OAI22_X1 U17513 ( .A1(n15626), .A2(n14329), .B1(n15616), .B2(n19858), .ZN(
        n14254) );
  AOI21_X1 U17514 ( .B1(n15623), .B2(n19854), .A(n14254), .ZN(n14255) );
  INV_X1 U17515 ( .A(n14255), .ZN(P1_U2850) );
  NOR2_X1 U17516 ( .A1(n14256), .A2(n14257), .ZN(n14258) );
  NOR2_X1 U17517 ( .A1(n14258), .A2(n14249), .ZN(n15637) );
  INV_X1 U17518 ( .A(n15637), .ZN(n14379) );
  NAND2_X1 U17519 ( .A1(n14265), .A2(n14259), .ZN(n14260) );
  AND2_X1 U17520 ( .A1(n14261), .A2(n14260), .ZN(n15636) );
  AOI22_X1 U17521 ( .A1(n15636), .A2(n19853), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n14303), .ZN(n14262) );
  OAI21_X1 U17522 ( .B1(n14379), .B2(n14322), .A(n14262), .ZN(P1_U2851) );
  XNOR2_X1 U17523 ( .A(n14263), .B(n14264), .ZN(n15641) );
  INV_X1 U17524 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14267) );
  OAI21_X1 U17525 ( .B1(n14269), .B2(n14266), .A(n14265), .ZN(n15645) );
  OAI222_X1 U17526 ( .A1(n15641), .A2(n14322), .B1(n14267), .B2(n19858), .C1(
        n15645), .C2(n14329), .ZN(P1_U2852) );
  AND2_X1 U17527 ( .A1(n14279), .A2(n14268), .ZN(n14270) );
  OR2_X1 U17528 ( .A1(n14270), .A2(n14269), .ZN(n15662) );
  INV_X1 U17529 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15651) );
  INV_X1 U17530 ( .A(n14263), .ZN(n14272) );
  AOI21_X1 U17531 ( .B1(n14273), .B2(n14271), .A(n14272), .ZN(n15752) );
  INV_X1 U17532 ( .A(n15752), .ZN(n14274) );
  OAI222_X1 U17533 ( .A1(n15662), .A2(n14329), .B1(n15651), .B2(n19858), .C1(
        n14274), .C2(n14322), .ZN(P1_U2853) );
  OAI21_X1 U17534 ( .B1(n14275), .B2(n14276), .A(n14271), .ZN(n14384) );
  INV_X1 U17535 ( .A(n14384), .ZN(n15667) );
  NAND2_X1 U17536 ( .A1(n14284), .A2(n14277), .ZN(n14278) );
  NAND2_X1 U17537 ( .A1(n14279), .A2(n14278), .ZN(n15813) );
  OAI22_X1 U17538 ( .A1(n15813), .A2(n14329), .B1(n20798), .B2(n19858), .ZN(
        n14280) );
  AOI21_X1 U17539 ( .B1(n15667), .B2(n19854), .A(n14280), .ZN(n14281) );
  INV_X1 U17540 ( .A(n14281), .ZN(P1_U2854) );
  OR2_X1 U17541 ( .A1(n14294), .A2(n14282), .ZN(n14283) );
  NAND2_X1 U17542 ( .A1(n14284), .A2(n14283), .ZN(n15824) );
  INV_X1 U17543 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14288) );
  NOR2_X1 U17544 ( .A1(n14285), .A2(n14286), .ZN(n14287) );
  OR2_X1 U17545 ( .A1(n14275), .A2(n14287), .ZN(n15764) );
  OAI222_X1 U17546 ( .A1(n15824), .A2(n14329), .B1(n14288), .B2(n19858), .C1(
        n15764), .C2(n14322), .ZN(P1_U2855) );
  AND2_X1 U17547 ( .A1(n14289), .A2(n14290), .ZN(n14291) );
  NOR2_X1 U17548 ( .A1(n14285), .A2(n14291), .ZN(n15684) );
  NOR2_X1 U17549 ( .A1(n14302), .A2(n14292), .ZN(n14293) );
  OR2_X1 U17550 ( .A1(n14294), .A2(n14293), .ZN(n15688) );
  OAI22_X1 U17551 ( .A1(n15688), .A2(n14329), .B1(n20755), .B2(n19858), .ZN(
        n14295) );
  AOI21_X1 U17552 ( .B1(n15684), .B2(n19854), .A(n14295), .ZN(n14296) );
  INV_X1 U17553 ( .A(n14296), .ZN(P1_U2856) );
  INV_X1 U17554 ( .A(n14289), .ZN(n14297) );
  AOI21_X1 U17555 ( .B1(n14298), .B2(n14215), .A(n14297), .ZN(n15776) );
  INV_X1 U17556 ( .A(n15776), .ZN(n14395) );
  AND2_X1 U17557 ( .A1(n14300), .A2(n14299), .ZN(n14301) );
  NOR2_X1 U17558 ( .A1(n14302), .A2(n14301), .ZN(n15835) );
  AOI22_X1 U17559 ( .A1(n15835), .A2(n19853), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n14303), .ZN(n14304) );
  OAI21_X1 U17560 ( .B1(n14395), .B2(n14322), .A(n14304), .ZN(P1_U2857) );
  OAI22_X1 U17561 ( .A1(n14710), .A2(n14329), .B1(n20836), .B2(n19858), .ZN(
        n14305) );
  INV_X1 U17562 ( .A(n14305), .ZN(n14306) );
  OAI21_X1 U17563 ( .B1(n14516), .B2(n14322), .A(n14306), .ZN(P1_U2858) );
  OAI21_X1 U17564 ( .B1(n14307), .B2(n9722), .A(n14308), .ZN(n14327) );
  OAI21_X1 U17565 ( .B1(n14327), .B2(n14328), .A(n14308), .ZN(n14316) );
  AOI21_X1 U17566 ( .B1(n14316), .B2(n14317), .A(n14309), .ZN(n14310) );
  OR2_X1 U17567 ( .A1(n14310), .A2(n14214), .ZN(n15702) );
  INV_X1 U17568 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15701) );
  OR2_X1 U17569 ( .A1(n14311), .A2(n14312), .ZN(n14313) );
  AND2_X1 U17570 ( .A1(n14314), .A2(n14313), .ZN(n15705) );
  INV_X1 U17571 ( .A(n15705), .ZN(n14315) );
  OAI222_X1 U17572 ( .A1(n15702), .A2(n14322), .B1(n15701), .B2(n19858), .C1(
        n14315), .C2(n14329), .ZN(P1_U2859) );
  XOR2_X1 U17573 ( .A(n14317), .B(n14316), .Z(n15779) );
  INV_X1 U17574 ( .A(n15779), .ZN(n14400) );
  INV_X1 U17575 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n20835) );
  INV_X1 U17576 ( .A(n14318), .ZN(n14320) );
  INV_X1 U17577 ( .A(n14319), .ZN(n14326) );
  AOI21_X1 U17578 ( .B1(n14320), .B2(n14326), .A(n14311), .ZN(n15708) );
  INV_X1 U17579 ( .A(n15708), .ZN(n14321) );
  OAI222_X1 U17580 ( .A1(n14400), .A2(n14322), .B1(n19858), .B2(n20835), .C1(
        n14321), .C2(n14329), .ZN(P1_U2860) );
  NAND2_X1 U17581 ( .A1(n14324), .A2(n14323), .ZN(n14325) );
  NAND2_X1 U17582 ( .A1(n14326), .A2(n14325), .ZN(n15840) );
  INV_X1 U17583 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15717) );
  XOR2_X1 U17584 ( .A(n14328), .B(n14327), .Z(n15789) );
  INV_X1 U17585 ( .A(n15789), .ZN(n14405) );
  OAI222_X1 U17586 ( .A1(n15840), .A2(n14329), .B1(n15717), .B2(n19858), .C1(
        n14405), .C2(n14322), .ZN(P1_U2861) );
  NAND2_X1 U17587 ( .A1(n14416), .A2(n15748), .ZN(n14335) );
  INV_X1 U17588 ( .A(DATAI_14_), .ZN(n14331) );
  MUX2_X1 U17589 ( .A(n14331), .B(n14330), .S(n20001), .Z(n19904) );
  NAND2_X1 U17590 ( .A1(n15744), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n14332) );
  OAI21_X1 U17591 ( .B1(n14389), .B2(n19904), .A(n14332), .ZN(n14333) );
  AOI21_X1 U17592 ( .B1(n15747), .B2(DATAI_30_), .A(n14333), .ZN(n14334) );
  OAI211_X1 U17593 ( .C1(n15751), .C2(n16228), .A(n14335), .B(n14334), .ZN(
        P1_U2874) );
  INV_X1 U17594 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n14340) );
  NAND2_X1 U17595 ( .A1(n15747), .A2(DATAI_29_), .ZN(n14339) );
  INV_X1 U17596 ( .A(n14389), .ZN(n15746) );
  INV_X1 U17597 ( .A(DATAI_13_), .ZN(n14337) );
  NAND2_X1 U17598 ( .A1(n20001), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14336) );
  OAI21_X1 U17599 ( .B1(n20001), .B2(n14337), .A(n14336), .ZN(n19902) );
  AOI22_X1 U17600 ( .A1(n15746), .A2(n19902), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n15744), .ZN(n14338) );
  OAI211_X1 U17601 ( .C1(n15751), .C2(n14340), .A(n14339), .B(n14338), .ZN(
        n14341) );
  AOI21_X1 U17602 ( .B1(n14426), .B2(n15748), .A(n14341), .ZN(n14342) );
  INV_X1 U17603 ( .A(n14342), .ZN(P1_U2875) );
  INV_X1 U17604 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n14349) );
  NAND2_X1 U17605 ( .A1(n14343), .A2(n15748), .ZN(n14348) );
  INV_X1 U17606 ( .A(DATAI_12_), .ZN(n14344) );
  MUX2_X1 U17607 ( .A(n14344), .B(n16254), .S(n20001), .Z(n19899) );
  NAND2_X1 U17608 ( .A1(n15744), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n14345) );
  OAI21_X1 U17609 ( .B1(n14389), .B2(n19899), .A(n14345), .ZN(n14346) );
  AOI21_X1 U17610 ( .B1(n15747), .B2(DATAI_28_), .A(n14346), .ZN(n14347) );
  OAI211_X1 U17611 ( .C1(n15751), .C2(n14349), .A(n14348), .B(n14347), .ZN(
        P1_U2876) );
  INV_X1 U17612 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n14356) );
  NAND2_X1 U17613 ( .A1(n14435), .A2(n15748), .ZN(n14355) );
  INV_X1 U17614 ( .A(DATAI_11_), .ZN(n14351) );
  MUX2_X1 U17615 ( .A(n14351), .B(n14350), .S(n20001), .Z(n19896) );
  NAND2_X1 U17616 ( .A1(n15744), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n14352) );
  OAI21_X1 U17617 ( .B1(n14389), .B2(n19896), .A(n14352), .ZN(n14353) );
  AOI21_X1 U17618 ( .B1(n15747), .B2(DATAI_27_), .A(n14353), .ZN(n14354) );
  OAI211_X1 U17619 ( .C1(n15751), .C2(n14356), .A(n14355), .B(n14354), .ZN(
        P1_U2877) );
  INV_X1 U17620 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n14359) );
  NAND2_X1 U17621 ( .A1(n15747), .A2(DATAI_26_), .ZN(n14358) );
  AOI22_X1 U17622 ( .A1(n15746), .A2(n19894), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n15744), .ZN(n14357) );
  OAI211_X1 U17623 ( .C1(n15751), .C2(n14359), .A(n14358), .B(n14357), .ZN(
        n14360) );
  INV_X1 U17624 ( .A(n14360), .ZN(n14361) );
  OAI21_X1 U17625 ( .B1(n14441), .B2(n14404), .A(n14361), .ZN(P1_U2878) );
  INV_X1 U17626 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n14366) );
  NAND2_X1 U17627 ( .A1(n14454), .A2(n15748), .ZN(n14365) );
  NAND2_X1 U17628 ( .A1(n15744), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n14362) );
  OAI21_X1 U17629 ( .B1(n14389), .B2(n19891), .A(n14362), .ZN(n14363) );
  AOI21_X1 U17630 ( .B1(n15747), .B2(DATAI_25_), .A(n14363), .ZN(n14364) );
  OAI211_X1 U17631 ( .C1(n15751), .C2(n14366), .A(n14365), .B(n14364), .ZN(
        P1_U2879) );
  INV_X1 U17632 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n14371) );
  NAND2_X1 U17633 ( .A1(n15603), .A2(n15748), .ZN(n14370) );
  NAND2_X1 U17634 ( .A1(n15744), .A2(P1_EAX_REG_24__SCAN_IN), .ZN(n14367) );
  OAI21_X1 U17635 ( .B1(n14389), .B2(n19888), .A(n14367), .ZN(n14368) );
  AOI21_X1 U17636 ( .B1(n15747), .B2(DATAI_24_), .A(n14368), .ZN(n14369) );
  OAI211_X1 U17637 ( .C1(n14371), .C2(n15751), .A(n14370), .B(n14369), .ZN(
        P1_U2880) );
  INV_X1 U17638 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n14375) );
  NAND2_X1 U17639 ( .A1(n15623), .A2(n15748), .ZN(n14374) );
  OAI22_X1 U17640 ( .A1(n20037), .A2(n14389), .B1(n14401), .B2(n13520), .ZN(
        n14372) );
  AOI21_X1 U17641 ( .B1(n15747), .B2(DATAI_22_), .A(n14372), .ZN(n14373) );
  OAI211_X1 U17642 ( .C1(n15751), .C2(n14375), .A(n14374), .B(n14373), .ZN(
        P1_U2882) );
  OAI22_X1 U17643 ( .A1(n20033), .A2(n14389), .B1(n14401), .B2(n13516), .ZN(
        n14376) );
  AOI21_X1 U17644 ( .B1(n15747), .B2(DATAI_21_), .A(n14376), .ZN(n14378) );
  INV_X1 U17645 ( .A(n15751), .ZN(n14386) );
  NAND2_X1 U17646 ( .A1(n14386), .A2(BUF1_REG_21__SCAN_IN), .ZN(n14377) );
  OAI211_X1 U17647 ( .C1(n14379), .C2(n14404), .A(n14378), .B(n14377), .ZN(
        P1_U2883) );
  OAI22_X1 U17648 ( .A1(n20022), .A2(n14389), .B1(n14401), .B2(n14380), .ZN(
        n14381) );
  AOI21_X1 U17649 ( .B1(n15747), .B2(DATAI_18_), .A(n14381), .ZN(n14383) );
  NAND2_X1 U17650 ( .A1(n14386), .A2(BUF1_REG_18__SCAN_IN), .ZN(n14382) );
  OAI211_X1 U17651 ( .C1(n14384), .C2(n14404), .A(n14383), .B(n14382), .ZN(
        P1_U2886) );
  OAI22_X1 U17652 ( .A1(n20019), .A2(n14389), .B1(n14401), .B2(n13518), .ZN(
        n14385) );
  AOI21_X1 U17653 ( .B1(n15747), .B2(DATAI_17_), .A(n14385), .ZN(n14388) );
  NAND2_X1 U17654 ( .A1(n14386), .A2(BUF1_REG_17__SCAN_IN), .ZN(n14387) );
  OAI211_X1 U17655 ( .C1(n15764), .C2(n14404), .A(n14388), .B(n14387), .ZN(
        P1_U2887) );
  INV_X1 U17656 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n14393) );
  NAND2_X1 U17657 ( .A1(n15684), .A2(n15748), .ZN(n14392) );
  OAI22_X1 U17658 ( .A1(n20010), .A2(n14389), .B1(n14401), .B2(n13524), .ZN(
        n14390) );
  AOI21_X1 U17659 ( .B1(n15747), .B2(DATAI_16_), .A(n14390), .ZN(n14391) );
  OAI211_X1 U17660 ( .C1(n15751), .C2(n14393), .A(n14392), .B(n14391), .ZN(
        P1_U2888) );
  OAI222_X1 U17661 ( .A1(n14404), .A2(n14395), .B1(n14403), .B2(n14394), .C1(
        n14401), .C2(n13339), .ZN(P1_U2889) );
  INV_X1 U17662 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14396) );
  OAI222_X1 U17663 ( .A1(n14516), .A2(n14404), .B1(n19904), .B2(n14403), .C1(
        n14396), .C2(n14401), .ZN(P1_U2890) );
  AOI22_X1 U17664 ( .A1(n14397), .A2(n19902), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15744), .ZN(n14398) );
  OAI21_X1 U17665 ( .B1(n15702), .B2(n14404), .A(n14398), .ZN(P1_U2891) );
  OAI222_X1 U17666 ( .A1(n14400), .A2(n14404), .B1(n19899), .B2(n14403), .C1(
        n14399), .C2(n14401), .ZN(P1_U2892) );
  INV_X1 U17667 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14402) );
  OAI222_X1 U17668 ( .A1(n14405), .A2(n14404), .B1(n19896), .B2(n14403), .C1(
        n14402), .C2(n14401), .ZN(P1_U2893) );
  INV_X1 U17669 ( .A(n14428), .ZN(n14407) );
  NOR4_X1 U17670 ( .A1(n14407), .A2(n14406), .A3(n14584), .A4(n14420), .ZN(
        n14409) );
  NOR2_X1 U17671 ( .A1(n14409), .A2(n14408), .ZN(n14411) );
  INV_X1 U17672 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14410) );
  XNOR2_X1 U17673 ( .A(n14411), .B(n14410), .ZN(n14574) );
  NAND2_X1 U17674 ( .A1(n15781), .A2(n14412), .ZN(n14413) );
  NAND2_X1 U17675 ( .A1(n19950), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14570) );
  OAI211_X1 U17676 ( .C1(n19938), .C2(n14414), .A(n14413), .B(n14570), .ZN(
        n14415) );
  AOI21_X1 U17677 ( .B1(n14416), .B2(n19942), .A(n14415), .ZN(n14417) );
  OAI21_X1 U17678 ( .B1(n14574), .B2(n19944), .A(n14417), .ZN(P1_U2969) );
  NAND2_X1 U17679 ( .A1(n14420), .A2(n14419), .ZN(n14421) );
  XNOR2_X1 U17680 ( .A(n14418), .B(n14421), .ZN(n14582) );
  NOR2_X1 U17681 ( .A1(n19823), .A2(n14422), .ZN(n14577) );
  AOI21_X1 U17682 ( .B1(n19925), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14577), .ZN(n14423) );
  OAI21_X1 U17683 ( .B1(n19934), .B2(n14424), .A(n14423), .ZN(n14425) );
  AOI21_X1 U17684 ( .B1(n14426), .B2(n19942), .A(n14425), .ZN(n14427) );
  OAI21_X1 U17685 ( .B1(n19944), .B2(n14582), .A(n14427), .ZN(P1_U2970) );
  MUX2_X1 U17686 ( .A(n9652), .B(n14428), .S(n15785), .Z(n14431) );
  XNOR2_X1 U17687 ( .A(n14431), .B(n14430), .ZN(n14602) );
  NAND2_X1 U17688 ( .A1(n19950), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14596) );
  NAND2_X1 U17689 ( .A1(n19925), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14432) );
  OAI211_X1 U17690 ( .C1(n19934), .C2(n14433), .A(n14596), .B(n14432), .ZN(
        n14434) );
  AOI21_X1 U17691 ( .B1(n14435), .B2(n19942), .A(n14434), .ZN(n14436) );
  OAI21_X1 U17692 ( .B1(n14602), .B2(n19944), .A(n14436), .ZN(P1_U2972) );
  NAND3_X1 U17693 ( .A1(n10013), .A2(n14438), .A3(n14437), .ZN(n14439) );
  XNOR2_X1 U17694 ( .A(n14439), .B(n14608), .ZN(n14616) );
  NAND2_X1 U17695 ( .A1(n19950), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14610) );
  OAI21_X1 U17696 ( .B1(n19938), .B2(n14440), .A(n14610), .ZN(n14443) );
  NOR2_X1 U17697 ( .A1(n14441), .A2(n20003), .ZN(n14442) );
  AOI211_X1 U17698 ( .C1(n15781), .C2(n14444), .A(n14443), .B(n14442), .ZN(
        n14445) );
  OAI21_X1 U17699 ( .B1(n19944), .B2(n14616), .A(n14445), .ZN(P1_U2973) );
  NOR2_X1 U17700 ( .A1(n14013), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14446) );
  MUX2_X1 U17701 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n14446), .S(
        n9590), .Z(n14449) );
  XNOR2_X1 U17702 ( .A(n14479), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14461) );
  NAND2_X1 U17703 ( .A1(n14013), .A2(n14461), .ZN(n14447) );
  NAND2_X1 U17704 ( .A1(n14447), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14448) );
  NAND2_X1 U17705 ( .A1(n14449), .A2(n14448), .ZN(n14450) );
  INV_X1 U17706 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14603) );
  XNOR2_X1 U17707 ( .A(n14450), .B(n14603), .ZN(n14625) );
  NAND2_X1 U17708 ( .A1(n19950), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14617) );
  NAND2_X1 U17709 ( .A1(n19925), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14451) );
  OAI211_X1 U17710 ( .C1(n19934), .C2(n14452), .A(n14617), .B(n14451), .ZN(
        n14453) );
  AOI21_X1 U17711 ( .B1(n14454), .B2(n19942), .A(n14453), .ZN(n14455) );
  OAI21_X1 U17712 ( .B1(n19944), .B2(n14625), .A(n14455), .ZN(P1_U2974) );
  INV_X1 U17713 ( .A(n14013), .ZN(n14456) );
  OAI211_X1 U17714 ( .C1(n14456), .C2(n14479), .A(n10013), .B(n14461), .ZN(
        n14457) );
  XOR2_X1 U17715 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n14457), .Z(
        n14634) );
  INV_X1 U17716 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20631) );
  NOR2_X1 U17717 ( .A1(n19823), .A2(n20631), .ZN(n14628) );
  INV_X1 U17718 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15598) );
  NOR2_X1 U17719 ( .A1(n19938), .A2(n15598), .ZN(n14458) );
  AOI211_X1 U17720 ( .C1(n15781), .C2(n15601), .A(n14628), .B(n14458), .ZN(
        n14460) );
  NAND2_X1 U17721 ( .A1(n15603), .A2(n19942), .ZN(n14459) );
  OAI211_X1 U17722 ( .C1(n14634), .C2(n19944), .A(n14460), .B(n14459), .ZN(
        P1_U2975) );
  XNOR2_X1 U17723 ( .A(n14013), .B(n14461), .ZN(n14646) );
  NAND2_X1 U17724 ( .A1(n14248), .A2(n14462), .ZN(n14463) );
  AND2_X1 U17725 ( .A1(n9716), .A2(n14463), .ZN(n15737) );
  NAND2_X1 U17726 ( .A1(n15737), .A2(n19942), .ZN(n14468) );
  INV_X1 U17727 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14464) );
  NOR2_X1 U17728 ( .A1(n19823), .A2(n14464), .ZN(n14639) );
  INV_X1 U17729 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14465) );
  NOR2_X1 U17730 ( .A1(n19938), .A2(n14465), .ZN(n14466) );
  AOI211_X1 U17731 ( .C1(n15781), .C2(n15607), .A(n14639), .B(n14466), .ZN(
        n14467) );
  OAI211_X1 U17732 ( .C1(n14646), .C2(n19944), .A(n14468), .B(n14467), .ZN(
        P1_U2976) );
  NAND2_X1 U17733 ( .A1(n14470), .A2(n14469), .ZN(n14471) );
  XNOR2_X1 U17734 ( .A(n14471), .B(n14657), .ZN(n14661) );
  NAND2_X1 U17735 ( .A1(n15781), .A2(n15620), .ZN(n14472) );
  NAND2_X1 U17736 ( .A1(n19950), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n14656) );
  OAI211_X1 U17737 ( .C1(n19938), .C2(n15617), .A(n14472), .B(n14656), .ZN(
        n14473) );
  AOI21_X1 U17738 ( .B1(n15623), .B2(n19942), .A(n14473), .ZN(n14474) );
  OAI21_X1 U17739 ( .B1(n14661), .B2(n19944), .A(n14474), .ZN(P1_U2977) );
  OAI21_X1 U17740 ( .B1(n15785), .B2(n15820), .A(n14475), .ZN(n14681) );
  INV_X1 U17741 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14476) );
  NAND2_X1 U17742 ( .A1(n9590), .A2(n14476), .ZN(n14680) );
  NAND2_X1 U17743 ( .A1(n14479), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14679) );
  OAI22_X1 U17744 ( .A1(n14681), .A2(n14680), .B1(n14475), .B2(n14679), .ZN(
        n14485) );
  NAND2_X1 U17745 ( .A1(n14485), .A2(n12012), .ZN(n14484) );
  INV_X1 U17746 ( .A(n14679), .ZN(n14477) );
  NAND2_X1 U17747 ( .A1(n14477), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14478) );
  OAI22_X1 U17748 ( .A1(n14484), .A2(n14479), .B1(n14475), .B2(n14478), .ZN(
        n14480) );
  XNOR2_X1 U17749 ( .A(n14480), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14669) );
  NAND2_X1 U17750 ( .A1(n19950), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14664) );
  NAND2_X1 U17751 ( .A1(n19925), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14481) );
  OAI211_X1 U17752 ( .C1(n19934), .C2(n15627), .A(n14664), .B(n14481), .ZN(
        n14482) );
  AOI21_X1 U17753 ( .B1(n15637), .B2(n19942), .A(n14482), .ZN(n14483) );
  OAI21_X1 U17754 ( .B1(n14669), .B2(n19944), .A(n14483), .ZN(P1_U2978) );
  OAI21_X1 U17755 ( .B1(n14485), .B2(n12012), .A(n14484), .ZN(n14670) );
  NAND2_X1 U17756 ( .A1(n14670), .A2(n19930), .ZN(n14488) );
  NAND2_X1 U17757 ( .A1(n19950), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n14675) );
  OAI21_X1 U17758 ( .B1(n19938), .B2(n15649), .A(n14675), .ZN(n14486) );
  AOI21_X1 U17759 ( .B1(n15781), .B2(n15640), .A(n14486), .ZN(n14487) );
  OAI211_X1 U17760 ( .C1(n20003), .C2(n15641), .A(n14488), .B(n14487), .ZN(
        P1_U2979) );
  OAI21_X1 U17761 ( .B1(n14490), .B2(n14489), .A(n14475), .ZN(n15814) );
  INV_X1 U17762 ( .A(n15663), .ZN(n14492) );
  AOI22_X1 U17763 ( .A1(n19925), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n19950), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14491) );
  OAI21_X1 U17764 ( .B1(n14492), .B2(n19934), .A(n14491), .ZN(n14493) );
  AOI21_X1 U17765 ( .B1(n15667), .B2(n19942), .A(n14493), .ZN(n14494) );
  OAI21_X1 U17766 ( .B1(n19944), .B2(n15814), .A(n14494), .ZN(P1_U2981) );
  AND2_X1 U17767 ( .A1(n14495), .A2(n14496), .ZN(n14508) );
  NOR2_X1 U17768 ( .A1(n14508), .A2(n14497), .ZN(n15770) );
  INV_X1 U17769 ( .A(n14498), .ZN(n14499) );
  OAI21_X1 U17770 ( .B1(n15770), .B2(n14499), .A(n15771), .ZN(n14500) );
  XOR2_X1 U17771 ( .A(n14501), .B(n14500), .Z(n14699) );
  NAND2_X1 U17772 ( .A1(n15781), .A2(n15678), .ZN(n14502) );
  NAND2_X1 U17773 ( .A1(n19950), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n14690) );
  OAI211_X1 U17774 ( .C1(n19938), .C2(n15681), .A(n14502), .B(n14690), .ZN(
        n14503) );
  AOI21_X1 U17775 ( .B1(n15684), .B2(n19942), .A(n14503), .ZN(n14504) );
  OAI21_X1 U17776 ( .B1(n14699), .B2(n19944), .A(n14504), .ZN(P1_U2983) );
  INV_X1 U17777 ( .A(n14505), .ZN(n14507) );
  OAI21_X1 U17778 ( .B1(n14508), .B2(n14507), .A(n14506), .ZN(n14510) );
  MUX2_X1 U17779 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n14068), .S(
        n15785), .Z(n14509) );
  XNOR2_X1 U17780 ( .A(n14510), .B(n14509), .ZN(n14713) );
  NAND2_X1 U17781 ( .A1(n14713), .A2(n19930), .ZN(n14515) );
  OR2_X1 U17782 ( .A1(n19823), .A2(n14219), .ZN(n14709) );
  INV_X1 U17783 ( .A(n14709), .ZN(n14513) );
  NOR2_X1 U17784 ( .A1(n19934), .A2(n14511), .ZN(n14512) );
  AOI211_X1 U17785 ( .C1(n19925), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n14513), .B(n14512), .ZN(n14514) );
  OAI211_X1 U17786 ( .C1(n20003), .C2(n14516), .A(n14515), .B(n14514), .ZN(
        P1_U2985) );
  INV_X1 U17787 ( .A(n14517), .ZN(n14522) );
  OAI21_X1 U17788 ( .B1(n14495), .B2(n14519), .A(n14518), .ZN(n14731) );
  MUX2_X1 U17789 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n14737), .S(
        n15785), .Z(n14732) );
  NOR2_X1 U17790 ( .A1(n14731), .A2(n14732), .ZN(n14730) );
  MUX2_X1 U17791 ( .A(n9736), .B(n14520), .S(n14730), .Z(n14521) );
  AOI21_X1 U17792 ( .B1(n14522), .B2(n14737), .A(n14521), .ZN(n14715) );
  NAND2_X1 U17793 ( .A1(n14715), .A2(n19930), .ZN(n14526) );
  INV_X1 U17794 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14523) );
  OAI22_X1 U17795 ( .A1(n19938), .A2(n14523), .B1(n19823), .B2(n20615), .ZN(
        n14524) );
  AOI21_X1 U17796 ( .B1(n15781), .B2(n15698), .A(n14524), .ZN(n14525) );
  OAI211_X1 U17797 ( .C1(n20003), .C2(n15702), .A(n14526), .B(n14525), .ZN(
        P1_U2986) );
  MUX2_X1 U17798 ( .A(n14527), .B(n14495), .S(n15785), .Z(n14528) );
  XOR2_X1 U17799 ( .A(n13898), .B(n14528), .Z(n15853) );
  NAND2_X1 U17800 ( .A1(n15853), .A2(n19930), .ZN(n14533) );
  INV_X1 U17801 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14529) );
  NOR2_X1 U17802 ( .A1(n19823), .A2(n14529), .ZN(n15848) );
  INV_X1 U17803 ( .A(n15729), .ZN(n14530) );
  NOR2_X1 U17804 ( .A1(n19934), .A2(n14530), .ZN(n14531) );
  AOI211_X1 U17805 ( .C1(n19925), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15848), .B(n14531), .ZN(n14532) );
  OAI211_X1 U17806 ( .C1(n20003), .C2(n15726), .A(n14533), .B(n14532), .ZN(
        P1_U2989) );
  NOR2_X1 U17807 ( .A1(n19957), .A2(n19967), .ZN(n19948) );
  NAND4_X1 U17808 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A4(n19948), .ZN(n15850) );
  NAND2_X1 U17809 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15879) );
  INV_X1 U17810 ( .A(n15879), .ZN(n15847) );
  NAND4_X1 U17811 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A4(n15847), .ZN(n14734) );
  NOR2_X1 U17812 ( .A1(n14535), .A2(n14734), .ZN(n14740) );
  NAND2_X1 U17813 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n14740), .ZN(
        n14537) );
  NOR2_X1 U17814 ( .A1(n15850), .A2(n14537), .ZN(n14718) );
  AND2_X1 U17815 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14718), .ZN(
        n14716) );
  NAND2_X1 U17816 ( .A1(n19969), .A2(n14716), .ZN(n14627) );
  OAI21_X1 U17817 ( .B1(n14536), .B2(n19972), .A(n19984), .ZN(n19945) );
  NAND3_X1 U17818 ( .A1(n19948), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n19945), .ZN(n14733) );
  OR2_X1 U17819 ( .A1(n14537), .A2(n14733), .ZN(n14701) );
  NOR2_X1 U17820 ( .A1(n14727), .A2(n14701), .ZN(n14691) );
  NAND2_X1 U17821 ( .A1(n19987), .A2(n14691), .ZN(n14538) );
  NAND2_X1 U17822 ( .A1(n14627), .A2(n14538), .ZN(n15817) );
  NAND4_X1 U17823 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15812) );
  NOR2_X1 U17824 ( .A1(n15820), .A2(n15812), .ZN(n14542) );
  AND4_X1 U17825 ( .A1(n14542), .A2(n12011), .A3(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14539) );
  NAND2_X1 U17826 ( .A1(n15817), .A2(n14539), .ZN(n14643) );
  NOR3_X1 U17827 ( .A1(n14643), .A2(n14607), .A3(n14608), .ZN(n14586) );
  NAND3_X1 U17828 ( .A1(n14586), .A2(n14541), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14566) );
  NAND2_X1 U17829 ( .A1(n14540), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14561) );
  INV_X1 U17830 ( .A(n14541), .ZN(n14585) );
  AND2_X1 U17831 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14542), .ZN(
        n14684) );
  AND2_X1 U17832 ( .A1(n14718), .A2(n14684), .ZN(n14545) );
  INV_X1 U17833 ( .A(n19970), .ZN(n14547) );
  NAND2_X1 U17834 ( .A1(n14542), .A2(n14691), .ZN(n14543) );
  NAND2_X1 U17835 ( .A1(n19987), .A2(n14543), .ZN(n14544) );
  OAI211_X1 U17836 ( .C1(n15869), .C2(n14545), .A(n14547), .B(n14544), .ZN(
        n14683) );
  NOR2_X1 U17837 ( .A1(n14683), .A2(n14546), .ZN(n14548) );
  AND2_X1 U17838 ( .A1(n14557), .A2(n14547), .ZN(n15851) );
  OR2_X1 U17839 ( .A1(n14548), .A2(n15851), .ZN(n14663) );
  NAND2_X1 U17840 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14654) );
  INV_X1 U17841 ( .A(n14654), .ZN(n14549) );
  OR2_X1 U17842 ( .A1(n14557), .A2(n14549), .ZN(n14550) );
  NAND2_X1 U17843 ( .A1(n14663), .A2(n14550), .ZN(n14640) );
  AND2_X1 U17844 ( .A1(n19987), .A2(n12013), .ZN(n14551) );
  NOR2_X1 U17845 ( .A1(n14640), .A2(n14551), .ZN(n14626) );
  INV_X1 U17846 ( .A(n19990), .ZN(n14671) );
  OR2_X1 U17847 ( .A1(n14671), .A2(n19987), .ZN(n14553) );
  INV_X1 U17848 ( .A(n14704), .ZN(n19988) );
  INV_X1 U17849 ( .A(n14604), .ZN(n14552) );
  AOI22_X1 U17850 ( .A1(n14553), .A2(n14607), .B1(n19988), .B2(n14552), .ZN(
        n14554) );
  NAND2_X1 U17851 ( .A1(n14626), .A2(n14554), .ZN(n14619) );
  NOR2_X1 U17852 ( .A1(n14619), .A2(n15874), .ZN(n14555) );
  INV_X1 U17853 ( .A(n14555), .ZN(n14558) );
  NOR3_X1 U17854 ( .A1(n14619), .A2(n14603), .A3(n14608), .ZN(n14556) );
  NOR2_X1 U17855 ( .A1(n14556), .A2(n14555), .ZN(n14595) );
  AOI21_X1 U17856 ( .B1(n14585), .B2(n14558), .A(n14595), .ZN(n14575) );
  OAI211_X1 U17857 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14557), .A(
        n14575), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14567) );
  NAND3_X1 U17858 ( .A1(n14567), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14558), .ZN(n14559) );
  OAI211_X1 U17859 ( .C1(n14566), .C2(n14561), .A(n14560), .B(n14559), .ZN(
        n14562) );
  AOI21_X1 U17860 ( .B1(n14563), .B2(n19993), .A(n14562), .ZN(n14564) );
  OAI21_X1 U17861 ( .B1(n14565), .B2(n19998), .A(n14564), .ZN(P1_U3000) );
  INV_X1 U17862 ( .A(n14566), .ZN(n14568) );
  OAI21_X1 U17863 ( .B1(n14568), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n14567), .ZN(n14569) );
  OAI211_X1 U17864 ( .C1(n14571), .C2(n19953), .A(n14570), .B(n14569), .ZN(
        n14572) );
  INV_X1 U17865 ( .A(n14572), .ZN(n14573) );
  OAI21_X1 U17866 ( .B1(n14574), .B2(n19998), .A(n14573), .ZN(P1_U3001) );
  INV_X1 U17867 ( .A(n14575), .ZN(n14578) );
  INV_X1 U17868 ( .A(n14586), .ZN(n14598) );
  NOR3_X1 U17869 ( .A1(n14598), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14585), .ZN(n14576) );
  AOI211_X1 U17870 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14578), .A(
        n14577), .B(n14576), .ZN(n14581) );
  NAND2_X1 U17871 ( .A1(n14579), .A2(n19993), .ZN(n14580) );
  OAI211_X1 U17872 ( .C1(n14582), .C2(n19998), .A(n14581), .B(n14580), .ZN(
        P1_U3002) );
  INV_X1 U17873 ( .A(n14583), .ZN(n14592) );
  INV_X1 U17874 ( .A(n14595), .ZN(n14590) );
  NAND3_X1 U17875 ( .A1(n14586), .A2(n14585), .A3(n14584), .ZN(n14588) );
  OAI211_X1 U17876 ( .C1(n14590), .C2(n14589), .A(n14588), .B(n14587), .ZN(
        n14591) );
  AOI21_X1 U17877 ( .B1(n14592), .B2(n19993), .A(n14591), .ZN(n14593) );
  OAI21_X1 U17878 ( .B1(n14594), .B2(n19998), .A(n14593), .ZN(P1_U3003) );
  NAND2_X1 U17879 ( .A1(n14595), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14597) );
  OAI211_X1 U17880 ( .C1(n14598), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14597), .B(n14596), .ZN(n14599) );
  AOI21_X1 U17881 ( .B1(n14600), .B2(n19993), .A(n14599), .ZN(n14601) );
  OAI21_X1 U17882 ( .B1(n14602), .B2(n19998), .A(n14601), .ZN(P1_U3004) );
  NAND2_X1 U17883 ( .A1(n14604), .A2(n14603), .ZN(n14605) );
  OR2_X1 U17884 ( .A1(n14643), .A2(n14605), .ZN(n14620) );
  INV_X1 U17885 ( .A(n14619), .ZN(n14606) );
  AOI21_X1 U17886 ( .B1(n14620), .B2(n14606), .A(n14608), .ZN(n14613) );
  INV_X1 U17887 ( .A(n14607), .ZN(n14609) );
  NAND2_X1 U17888 ( .A1(n14609), .A2(n14608), .ZN(n14611) );
  OAI21_X1 U17889 ( .B1(n14643), .B2(n14611), .A(n14610), .ZN(n14612) );
  AOI211_X1 U17890 ( .C1(n14614), .C2(n19993), .A(n14613), .B(n14612), .ZN(
        n14615) );
  OAI21_X1 U17891 ( .B1(n14616), .B2(n19998), .A(n14615), .ZN(P1_U3005) );
  INV_X1 U17892 ( .A(n14617), .ZN(n14618) );
  AOI21_X1 U17893 ( .B1(n14619), .B2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n14618), .ZN(n14621) );
  OAI211_X1 U17894 ( .C1(n14622), .C2(n19953), .A(n14621), .B(n14620), .ZN(
        n14623) );
  INV_X1 U17895 ( .A(n14623), .ZN(n14624) );
  OAI21_X1 U17896 ( .B1(n14625), .B2(n19998), .A(n14624), .ZN(P1_U3006) );
  OAI21_X1 U17897 ( .B1(n14627), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n14626), .ZN(n14632) );
  NOR3_X1 U17898 ( .A1(n14643), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n12013), .ZN(n14631) );
  INV_X1 U17899 ( .A(n14628), .ZN(n14629) );
  OAI21_X1 U17900 ( .B1(n15606), .B2(n19953), .A(n14629), .ZN(n14630) );
  AOI211_X1 U17901 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n14632), .A(
        n14631), .B(n14630), .ZN(n14633) );
  OAI21_X1 U17902 ( .B1(n14634), .B2(n19998), .A(n14633), .ZN(P1_U3007) );
  AND2_X1 U17903 ( .A1(n14636), .A2(n14635), .ZN(n14637) );
  NOR2_X1 U17904 ( .A1(n14638), .A2(n14637), .ZN(n15734) );
  NAND2_X1 U17905 ( .A1(n15734), .A2(n19993), .ZN(n14642) );
  AOI21_X1 U17906 ( .B1(n14640), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n14639), .ZN(n14641) );
  OAI211_X1 U17907 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n14643), .A(
        n14642), .B(n14641), .ZN(n14644) );
  INV_X1 U17908 ( .A(n14644), .ZN(n14645) );
  OAI21_X1 U17909 ( .B1(n14646), .B2(n19998), .A(n14645), .ZN(P1_U3008) );
  INV_X1 U17910 ( .A(n15626), .ZN(n14659) );
  INV_X1 U17911 ( .A(n14701), .ZN(n14647) );
  NAND2_X1 U17912 ( .A1(n19987), .A2(n14647), .ZN(n14650) );
  NAND2_X1 U17913 ( .A1(n14718), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14648) );
  OR2_X1 U17914 ( .A1(n14704), .A2(n14648), .ZN(n14649) );
  NAND2_X1 U17915 ( .A1(n14650), .A2(n14649), .ZN(n14706) );
  INV_X1 U17916 ( .A(n14718), .ZN(n14651) );
  NOR2_X1 U17917 ( .A1(n19990), .A2(n14651), .ZN(n14652) );
  OR2_X1 U17918 ( .A1(n14706), .A2(n14652), .ZN(n14673) );
  NAND3_X1 U17919 ( .A1(n14673), .A2(n14684), .A3(n12011), .ZN(n14665) );
  AOI21_X1 U17920 ( .B1(n14662), .B2(n14657), .A(n14665), .ZN(n14653) );
  NAND2_X1 U17921 ( .A1(n14654), .A2(n14653), .ZN(n14655) );
  OAI211_X1 U17922 ( .C1(n14663), .C2(n14657), .A(n14656), .B(n14655), .ZN(
        n14658) );
  AOI21_X1 U17923 ( .B1(n14659), .B2(n19993), .A(n14658), .ZN(n14660) );
  OAI21_X1 U17924 ( .B1(n14661), .B2(n19998), .A(n14660), .ZN(P1_U3009) );
  NOR2_X1 U17925 ( .A1(n14663), .A2(n14662), .ZN(n14667) );
  OAI21_X1 U17926 ( .B1(n14665), .B2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n14664), .ZN(n14666) );
  AOI211_X1 U17927 ( .C1(n15636), .C2(n19993), .A(n14667), .B(n14666), .ZN(
        n14668) );
  OAI21_X1 U17928 ( .B1(n14669), .B2(n19998), .A(n14668), .ZN(P1_U3010) );
  NAND2_X1 U17929 ( .A1(n14670), .A2(n19973), .ZN(n14678) );
  NOR2_X1 U17930 ( .A1(n14706), .A2(n14671), .ZN(n14672) );
  NOR2_X1 U17931 ( .A1(n14672), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14685) );
  OAI21_X1 U17932 ( .B1(n14685), .B2(n14683), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14676) );
  NAND4_X1 U17933 ( .A1(n14673), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n14684), .A4(n12012), .ZN(n14674) );
  AND3_X1 U17934 ( .A1(n14676), .A2(n14675), .A3(n14674), .ZN(n14677) );
  OAI211_X1 U17935 ( .C1(n19953), .C2(n15645), .A(n14678), .B(n14677), .ZN(
        P1_U3011) );
  NAND2_X1 U17936 ( .A1(n14680), .A2(n14679), .ZN(n14682) );
  XOR2_X1 U17937 ( .A(n14682), .B(n14681), .Z(n15753) );
  AOI22_X1 U17938 ( .A1(n14683), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n19950), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n14687) );
  OAI211_X1 U17939 ( .C1(n14718), .C2(n14706), .A(n14685), .B(n14684), .ZN(
        n14686) );
  OAI211_X1 U17940 ( .C1(n15662), .C2(n19953), .A(n14687), .B(n14686), .ZN(
        n14688) );
  AOI21_X1 U17941 ( .B1(n15753), .B2(n19973), .A(n14688), .ZN(n14689) );
  INV_X1 U17942 ( .A(n14689), .ZN(P1_U3012) );
  INV_X1 U17943 ( .A(n15688), .ZN(n14697) );
  INV_X1 U17944 ( .A(n14690), .ZN(n14696) );
  INV_X1 U17945 ( .A(n14691), .ZN(n14700) );
  AOI21_X1 U17946 ( .B1(n19987), .B2(n14700), .A(n19970), .ZN(n14692) );
  OAI21_X1 U17947 ( .B1(n15869), .B2(n14716), .A(n14692), .ZN(n15811) );
  AOI21_X1 U17948 ( .B1(n14068), .B2(n15874), .A(n15811), .ZN(n15838) );
  NAND2_X1 U17949 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15817), .ZN(
        n15830) );
  NAND2_X1 U17950 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15823) );
  OAI21_X1 U17951 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n15823), .ZN(n14693) );
  OAI22_X1 U17952 ( .A1(n15838), .A2(n14694), .B1(n15830), .B2(n14693), .ZN(
        n14695) );
  AOI211_X1 U17953 ( .C1(n19993), .C2(n14697), .A(n14696), .B(n14695), .ZN(
        n14698) );
  OAI21_X1 U17954 ( .B1(n14699), .B2(n19998), .A(n14698), .ZN(P1_U3015) );
  NAND3_X1 U17955 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n19969), .ZN(n15873) );
  NAND2_X1 U17956 ( .A1(n14736), .A2(n15873), .ZN(n15895) );
  INV_X1 U17957 ( .A(n15895), .ZN(n14729) );
  NOR3_X1 U17958 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n14729), .A3(
        n14700), .ZN(n14712) );
  NAND2_X1 U17959 ( .A1(n19987), .A2(n14701), .ZN(n14703) );
  OR2_X1 U17960 ( .A1(n19990), .A2(n14716), .ZN(n14702) );
  OAI211_X1 U17961 ( .C1(n14718), .C2(n14704), .A(n14703), .B(n14702), .ZN(
        n14705) );
  NOR2_X1 U17962 ( .A1(n14705), .A2(n19970), .ZN(n14728) );
  NAND2_X1 U17963 ( .A1(n14727), .A2(n14706), .ZN(n14719) );
  AOI21_X1 U17964 ( .B1(n14728), .B2(n14719), .A(n14068), .ZN(n14707) );
  INV_X1 U17965 ( .A(n14707), .ZN(n14708) );
  OAI211_X1 U17966 ( .C1(n14710), .C2(n19953), .A(n14709), .B(n14708), .ZN(
        n14711) );
  AOI211_X1 U17967 ( .C1(n14713), .C2(n19973), .A(n14712), .B(n14711), .ZN(
        n14714) );
  INV_X1 U17968 ( .A(n14714), .ZN(P1_U3017) );
  NAND2_X1 U17969 ( .A1(n14715), .A2(n19973), .ZN(n14726) );
  NOR2_X1 U17970 ( .A1(n14716), .A2(n19990), .ZN(n14717) );
  NAND2_X1 U17971 ( .A1(n14718), .A2(n14717), .ZN(n14723) );
  NOR2_X1 U17972 ( .A1(n19823), .A2(n20615), .ZN(n14721) );
  INV_X1 U17973 ( .A(n14719), .ZN(n14720) );
  NOR2_X1 U17974 ( .A1(n14721), .A2(n14720), .ZN(n14722) );
  NAND2_X1 U17975 ( .A1(n14723), .A2(n14722), .ZN(n14724) );
  AOI21_X1 U17976 ( .B1(n15705), .B2(n19993), .A(n14724), .ZN(n14725) );
  OAI211_X1 U17977 ( .C1(n14728), .C2(n14727), .A(n14726), .B(n14725), .ZN(
        P1_U3018) );
  NOR2_X1 U17978 ( .A1(n15894), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14741) );
  AOI21_X1 U17979 ( .B1(n14732), .B2(n14731), .A(n14730), .ZN(n15784) );
  NOR2_X1 U17980 ( .A1(n14734), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15839) );
  AOI21_X1 U17981 ( .B1(n19987), .B2(n14733), .A(n19970), .ZN(n15870) );
  INV_X1 U17982 ( .A(n15869), .ZN(n19971) );
  OAI21_X1 U17983 ( .B1(n15850), .B2(n14734), .A(n19971), .ZN(n14735) );
  OAI211_X1 U17984 ( .C1(n14740), .C2(n14736), .A(n15870), .B(n14735), .ZN(
        n15843) );
  AOI21_X1 U17985 ( .B1(n19969), .B2(n15839), .A(n15843), .ZN(n14738) );
  INV_X1 U17986 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14737) );
  OAI22_X1 U17987 ( .A1(n15784), .A2(n19998), .B1(n14738), .B2(n14737), .ZN(
        n14739) );
  AOI21_X1 U17988 ( .B1(n14741), .B2(n14740), .A(n14739), .ZN(n14743) );
  AOI22_X1 U17989 ( .A1(n15708), .A2(n19993), .B1(n19950), .B2(
        P1_REIP_REG_12__SCAN_IN), .ZN(n14742) );
  NAND2_X1 U17990 ( .A1(n14743), .A2(n14742), .ZN(P1_U3019) );
  OAI21_X1 U17991 ( .B1(n16004), .B2(n14744), .A(n18882), .ZN(n14746) );
  AOI22_X1 U17992 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18901), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18890), .ZN(n14745) );
  OAI21_X1 U17993 ( .B1(n14747), .B2(n14746), .A(n14745), .ZN(n14748) );
  AOI21_X1 U17994 ( .B1(P2_EBX_REG_22__SCAN_IN), .B2(n18889), .A(n14748), .ZN(
        n14756) );
  INV_X1 U17995 ( .A(n14749), .ZN(n14750) );
  AOI21_X1 U17996 ( .B1(n14751), .B2(n14761), .A(n14750), .ZN(n16084) );
  NOR2_X1 U17997 ( .A1(n14752), .A2(n14764), .ZN(n14753) );
  OR2_X1 U17998 ( .A1(n14754), .A2(n14753), .ZN(n16079) );
  INV_X1 U17999 ( .A(n16079), .ZN(n15977) );
  AOI22_X1 U18000 ( .A1(n16084), .A2(n18896), .B1(n15977), .B2(n18877), .ZN(
        n14755) );
  OAI211_X1 U18001 ( .C1(n14757), .C2(n18888), .A(n14756), .B(n14755), .ZN(
        P2_U2833) );
  AOI21_X1 U18002 ( .B1(n9828), .B2(n14771), .A(n19606), .ZN(n14774) );
  OR2_X1 U18003 ( .A1(n14758), .A2(n14759), .ZN(n14760) );
  NAND2_X1 U18004 ( .A1(n14761), .A2(n14760), .ZN(n15020) );
  INV_X1 U18005 ( .A(n15020), .ZN(n15162) );
  OAI22_X1 U18006 ( .A1(n15019), .A2(n18874), .B1(n19649), .B2(n18849), .ZN(
        n14768) );
  OR2_X1 U18007 ( .A1(n14762), .A2(n14763), .ZN(n14766) );
  INV_X1 U18008 ( .A(n14764), .ZN(n14765) );
  NAND2_X1 U18009 ( .A1(n14766), .A2(n14765), .ZN(n15160) );
  NOR2_X1 U18010 ( .A1(n15160), .A2(n18893), .ZN(n14767) );
  AOI211_X1 U18011 ( .C1(n15162), .C2(n18896), .A(n14768), .B(n14767), .ZN(
        n14769) );
  OAI21_X1 U18012 ( .B1(n14770), .B2(n18888), .A(n14769), .ZN(n14773) );
  NAND2_X1 U18013 ( .A1(n18899), .A2(n14771), .ZN(n14782) );
  OAI22_X1 U18014 ( .A1(n15023), .A2(n14782), .B1(n18857), .B2(n14848), .ZN(
        n14772) );
  AOI211_X1 U18015 ( .C1(n15023), .C2(n14774), .A(n14773), .B(n14772), .ZN(
        n14775) );
  INV_X1 U18016 ( .A(n14775), .ZN(P2_U2834) );
  NOR2_X1 U18017 ( .A1(n14857), .A2(n14776), .ZN(n14777) );
  OR2_X1 U18018 ( .A1(n14758), .A2(n14777), .ZN(n15174) );
  INV_X1 U18019 ( .A(n15034), .ZN(n14778) );
  NAND2_X1 U18020 ( .A1(n18865), .A2(n18882), .ZN(n18886) );
  INV_X1 U18021 ( .A(n18886), .ZN(n18900) );
  AOI22_X1 U18022 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18901), .B1(
        n14778), .B2(n18900), .ZN(n14780) );
  AOI22_X1 U18023 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n18889), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18890), .ZN(n14779) );
  OAI211_X1 U18024 ( .C1(n15174), .C2(n18871), .A(n14780), .B(n14779), .ZN(
        n14781) );
  INV_X1 U18025 ( .A(n14781), .ZN(n14791) );
  INV_X1 U18026 ( .A(n14782), .ZN(n14783) );
  OAI21_X1 U18027 ( .B1(n14784), .B2(n15034), .A(n14783), .ZN(n14790) );
  NOR2_X1 U18028 ( .A1(n14785), .A2(n14786), .ZN(n14787) );
  NOR2_X1 U18029 ( .A1(n14762), .A2(n14787), .ZN(n15983) );
  AOI22_X1 U18030 ( .A1(n14788), .A2(n18876), .B1(n15983), .B2(n18877), .ZN(
        n14789) );
  NAND3_X1 U18031 ( .A1(n14791), .A2(n14790), .A3(n14789), .ZN(P2_U2835) );
  INV_X1 U18032 ( .A(n14792), .ZN(n14793) );
  NAND2_X1 U18033 ( .A1(n14793), .A2(n14796), .ZN(n14794) );
  OAI21_X1 U18034 ( .B1(n14796), .B2(n14795), .A(n14794), .ZN(P2_U2856) );
  NAND2_X1 U18035 ( .A1(n14798), .A2(n14797), .ZN(n14800) );
  XNOR2_X1 U18036 ( .A(n14800), .B(n14799), .ZN(n14880) );
  NOR2_X1 U18037 ( .A1(n15941), .A2(n13122), .ZN(n14801) );
  AOI21_X1 U18038 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n13122), .A(n14801), .ZN(
        n14802) );
  OAI21_X1 U18039 ( .B1(n14880), .B2(n14854), .A(n14802), .ZN(P2_U2859) );
  AOI21_X1 U18040 ( .B1(n14805), .B2(n14804), .A(n14803), .ZN(n14806) );
  INV_X1 U18041 ( .A(n14806), .ZN(n14886) );
  NOR2_X1 U18042 ( .A1(n15108), .A2(n14861), .ZN(n14807) );
  AOI21_X1 U18043 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n14861), .A(n14807), .ZN(
        n14808) );
  OAI21_X1 U18044 ( .B1(n14886), .B2(n14854), .A(n14808), .ZN(P2_U2860) );
  NAND2_X1 U18045 ( .A1(n14809), .A2(n14810), .ZN(n14811) );
  NAND2_X1 U18046 ( .A1(n14812), .A2(n14811), .ZN(n15948) );
  AOI21_X1 U18047 ( .B1(n14815), .B2(n14814), .A(n14813), .ZN(n14887) );
  NAND2_X1 U18048 ( .A1(n14887), .A2(n14860), .ZN(n14817) );
  NAND2_X1 U18049 ( .A1(n14861), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14816) );
  OAI211_X1 U18050 ( .C1(n14861), .C2(n15948), .A(n14817), .B(n14816), .ZN(
        P2_U2861) );
  OAI21_X1 U18051 ( .B1(n14820), .B2(n14819), .A(n14818), .ZN(n14905) );
  OAI21_X1 U18052 ( .B1(n14831), .B2(n14821), .A(n14809), .ZN(n15126) );
  NOR2_X1 U18053 ( .A1(n15126), .A2(n13122), .ZN(n14822) );
  AOI21_X1 U18054 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n13122), .A(n14822), .ZN(
        n14823) );
  OAI21_X1 U18055 ( .B1(n14905), .B2(n14854), .A(n14823), .ZN(P2_U2862) );
  INV_X1 U18056 ( .A(n14824), .ZN(n14828) );
  AOI21_X1 U18057 ( .B1(n14828), .B2(n14827), .A(n14826), .ZN(n14829) );
  XOR2_X1 U18058 ( .A(n14830), .B(n14829), .Z(n14913) );
  AOI21_X1 U18059 ( .B1(n14833), .B2(n14832), .A(n14831), .ZN(n14984) );
  INV_X1 U18060 ( .A(n14984), .ZN(n15975) );
  MUX2_X1 U18061 ( .A(n14834), .B(n15975), .S(n14796), .Z(n14835) );
  OAI21_X1 U18062 ( .B1(n14913), .B2(n14854), .A(n14835), .ZN(P2_U2863) );
  AOI21_X1 U18063 ( .B1(n14838), .B2(n14837), .A(n14836), .ZN(n14839) );
  INV_X1 U18064 ( .A(n14839), .ZN(n14919) );
  MUX2_X1 U18065 ( .A(n15146), .B(n10787), .S(n14861), .Z(n14840) );
  OAI21_X1 U18066 ( .B1(n14919), .B2(n14854), .A(n14840), .ZN(P2_U2864) );
  INV_X1 U18067 ( .A(n16084), .ZN(n14845) );
  AOI21_X1 U18068 ( .B1(n14842), .B2(n14841), .A(n9701), .ZN(n15978) );
  NAND2_X1 U18069 ( .A1(n15978), .A2(n14860), .ZN(n14844) );
  NAND2_X1 U18070 ( .A1(n14861), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14843) );
  OAI211_X1 U18071 ( .C1(n14845), .C2(n14861), .A(n14844), .B(n14843), .ZN(
        P2_U2865) );
  OAI21_X1 U18072 ( .B1(n14846), .B2(n14847), .A(n14841), .ZN(n14925) );
  MUX2_X1 U18073 ( .A(n15020), .B(n14848), .S(n14861), .Z(n14849) );
  OAI21_X1 U18074 ( .B1(n14925), .B2(n14854), .A(n14849), .ZN(P2_U2866) );
  NOR2_X1 U18075 ( .A1(n9723), .A2(n14850), .ZN(n14851) );
  OR2_X1 U18076 ( .A1(n14846), .A2(n14851), .ZN(n15985) );
  MUX2_X1 U18077 ( .A(n15174), .B(n14852), .S(n13122), .Z(n14853) );
  OAI21_X1 U18078 ( .B1(n15985), .B2(n14854), .A(n14853), .ZN(P2_U2867) );
  AND2_X1 U18079 ( .A1(n14856), .A2(n14855), .ZN(n14858) );
  OR2_X1 U18080 ( .A1(n14858), .A2(n14857), .ZN(n18689) );
  AOI21_X1 U18081 ( .B1(n14859), .B2(n13934), .A(n9723), .ZN(n14926) );
  NAND2_X1 U18082 ( .A1(n14926), .A2(n14860), .ZN(n14863) );
  NAND2_X1 U18083 ( .A1(n14861), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n14862) );
  OAI211_X1 U18084 ( .C1(n18689), .C2(n13122), .A(n14863), .B(n14862), .ZN(
        P2_U2868) );
  NAND3_X1 U18085 ( .A1(n14865), .A2(n18945), .A3(n14864), .ZN(n14875) );
  NOR2_X1 U18086 ( .A1(n14867), .A2(n14866), .ZN(n14868) );
  INV_X1 U18087 ( .A(n15092), .ZN(n14872) );
  OAI22_X1 U18088 ( .A1(n14930), .A2(n18924), .B1(n18953), .B2(n14870), .ZN(
        n14871) );
  AOI21_X1 U18089 ( .B1(n14872), .B2(n18964), .A(n14871), .ZN(n14874) );
  AOI22_X1 U18090 ( .A1(n18910), .A2(BUF2_REG_29__SCAN_IN), .B1(n18911), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14873) );
  NAND3_X1 U18091 ( .A1(n14875), .A2(n14874), .A3(n14873), .ZN(P2_U2890) );
  INV_X1 U18092 ( .A(n18926), .ZN(n14876) );
  OAI22_X1 U18093 ( .A1(n14930), .A2(n14876), .B1(n18953), .B2(n13171), .ZN(
        n14877) );
  AOI21_X1 U18094 ( .B1(n15939), .B2(n18964), .A(n14877), .ZN(n14879) );
  AOI22_X1 U18095 ( .A1(n18910), .A2(BUF2_REG_28__SCAN_IN), .B1(n18911), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n14878) );
  OAI211_X1 U18096 ( .C1(n14880), .C2(n18968), .A(n14879), .B(n14878), .ZN(
        P2_U2891) );
  OAI22_X1 U18097 ( .A1(n14930), .A2(n18929), .B1(n18953), .B2(n14882), .ZN(
        n14883) );
  AOI21_X1 U18098 ( .B1(n18964), .B2(n15105), .A(n14883), .ZN(n14885) );
  AOI22_X1 U18099 ( .A1(n18910), .A2(BUF2_REG_27__SCAN_IN), .B1(n18911), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n14884) );
  OAI211_X1 U18100 ( .C1(n14886), .C2(n18968), .A(n14885), .B(n14884), .ZN(
        P2_U2892) );
  NAND2_X1 U18101 ( .A1(n14887), .A2(n18945), .ZN(n14895) );
  AOI22_X1 U18102 ( .A1(n18909), .A2(n18931), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n18963), .ZN(n14894) );
  AOI22_X1 U18103 ( .A1(n18910), .A2(BUF2_REG_26__SCAN_IN), .B1(n18911), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n14893) );
  INV_X1 U18104 ( .A(n14888), .ZN(n14891) );
  INV_X1 U18105 ( .A(n14889), .ZN(n14898) );
  AOI21_X1 U18106 ( .B1(n14891), .B2(n14898), .A(n14890), .ZN(n15951) );
  NAND2_X1 U18107 ( .A1(n18964), .A2(n15951), .ZN(n14892) );
  NAND4_X1 U18108 ( .A1(n14895), .A2(n14894), .A3(n14893), .A4(n14892), .ZN(
        P2_U2893) );
  INV_X1 U18109 ( .A(n14896), .ZN(n14906) );
  INV_X1 U18110 ( .A(n14897), .ZN(n14899) );
  OAI21_X1 U18111 ( .B1(n14906), .B2(n14899), .A(n14898), .ZN(n15964) );
  INV_X1 U18112 ( .A(n15964), .ZN(n14902) );
  OAI22_X1 U18113 ( .A1(n14930), .A2(n18934), .B1(n18953), .B2(n14900), .ZN(
        n14901) );
  AOI21_X1 U18114 ( .B1(n18964), .B2(n14902), .A(n14901), .ZN(n14904) );
  AOI22_X1 U18115 ( .A1(n18910), .A2(BUF2_REG_25__SCAN_IN), .B1(n18911), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n14903) );
  OAI211_X1 U18116 ( .C1(n14905), .C2(n18968), .A(n14904), .B(n14903), .ZN(
        P2_U2894) );
  AOI21_X1 U18117 ( .B1(n14908), .B2(n14907), .A(n14906), .ZN(n15973) );
  INV_X1 U18118 ( .A(n18938), .ZN(n14909) );
  OAI22_X1 U18119 ( .A1(n14930), .A2(n14909), .B1(n18953), .B2(n13169), .ZN(
        n14910) );
  AOI21_X1 U18120 ( .B1(n18964), .B2(n15973), .A(n14910), .ZN(n14912) );
  AOI22_X1 U18121 ( .A1(n18910), .A2(BUF2_REG_24__SCAN_IN), .B1(n18911), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14911) );
  OAI211_X1 U18122 ( .C1(n14913), .C2(n18968), .A(n14912), .B(n14911), .ZN(
        P2_U2895) );
  INV_X1 U18123 ( .A(n15150), .ZN(n14916) );
  OAI22_X1 U18124 ( .A1(n14930), .A2(n19069), .B1(n18953), .B2(n14914), .ZN(
        n14915) );
  AOI21_X1 U18125 ( .B1(n18964), .B2(n14916), .A(n14915), .ZN(n14918) );
  AOI22_X1 U18126 ( .A1(n18910), .A2(BUF2_REG_23__SCAN_IN), .B1(n18911), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n14917) );
  OAI211_X1 U18127 ( .C1(n14919), .C2(n18968), .A(n14918), .B(n14917), .ZN(
        P2_U2896) );
  INV_X1 U18128 ( .A(n15160), .ZN(n14922) );
  OAI22_X1 U18129 ( .A1(n14930), .A2(n19053), .B1(n18953), .B2(n14920), .ZN(
        n14921) );
  AOI21_X1 U18130 ( .B1(n18964), .B2(n14922), .A(n14921), .ZN(n14924) );
  AOI22_X1 U18131 ( .A1(n18910), .A2(BUF2_REG_21__SCAN_IN), .B1(n18911), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n14923) );
  OAI211_X1 U18132 ( .C1(n14925), .C2(n18968), .A(n14924), .B(n14923), .ZN(
        P2_U2898) );
  INV_X1 U18133 ( .A(n14926), .ZN(n14934) );
  NOR2_X1 U18134 ( .A1(n15198), .A2(n14927), .ZN(n14928) );
  OAI22_X1 U18135 ( .A1(n14930), .A2(n19046), .B1(n18953), .B2(n14929), .ZN(
        n14931) );
  AOI21_X1 U18136 ( .B1(n18964), .B2(n10069), .A(n14931), .ZN(n14933) );
  AOI22_X1 U18137 ( .A1(n18910), .A2(BUF2_REG_19__SCAN_IN), .B1(n18911), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n14932) );
  OAI211_X1 U18138 ( .C1(n14934), .C2(n18968), .A(n14933), .B(n14932), .ZN(
        P2_U2900) );
  NAND2_X1 U18139 ( .A1(n14936), .A2(n14935), .ZN(n14938) );
  XOR2_X1 U18140 ( .A(n14938), .B(n14937), .Z(n15104) );
  AOI21_X1 U18141 ( .B1(n15096), .B2(n14940), .A(n14939), .ZN(n15102) );
  NAND2_X1 U18142 ( .A1(n19011), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15091) );
  OAI21_X1 U18143 ( .B1(n16059), .B2(n14941), .A(n15091), .ZN(n14942) );
  AOI21_X1 U18144 ( .B1(n16052), .B2(n15926), .A(n14942), .ZN(n14943) );
  OAI21_X1 U18145 ( .B1(n15930), .B2(n19020), .A(n14943), .ZN(n14944) );
  AOI21_X1 U18146 ( .B1(n15102), .B2(n19015), .A(n14944), .ZN(n14945) );
  OAI21_X1 U18147 ( .B1(n15104), .B2(n16072), .A(n14945), .ZN(P2_U2985) );
  XNOR2_X1 U18148 ( .A(n14946), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15114) );
  AOI21_X1 U18149 ( .B1(n14948), .B2(n14947), .A(n12475), .ZN(n15111) );
  NAND2_X1 U18150 ( .A1(n19011), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15107) );
  OAI21_X1 U18151 ( .B1(n16059), .B2(n14949), .A(n15107), .ZN(n14950) );
  AOI21_X1 U18152 ( .B1(n16052), .B2(n14951), .A(n14950), .ZN(n14952) );
  OAI21_X1 U18153 ( .B1(n15108), .B2(n19020), .A(n14952), .ZN(n14953) );
  AOI21_X1 U18154 ( .B1(n15111), .B2(n19015), .A(n14953), .ZN(n14954) );
  OAI21_X1 U18155 ( .B1(n15114), .B2(n16072), .A(n14954), .ZN(P2_U2987) );
  NAND2_X1 U18156 ( .A1(n14955), .A2(n14966), .ZN(n14956) );
  XOR2_X1 U18157 ( .A(n14957), .B(n14956), .Z(n15125) );
  INV_X1 U18158 ( .A(n15948), .ZN(n14963) );
  NOR2_X1 U18159 ( .A1(n18847), .A2(n14958), .ZN(n15117) );
  AOI21_X1 U18160 ( .B1(n19012), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15117), .ZN(n14959) );
  OAI21_X1 U18161 ( .B1(n19025), .B2(n14960), .A(n14959), .ZN(n14962) );
  OAI21_X1 U18162 ( .B1(n14969), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14947), .ZN(n15119) );
  NOR2_X1 U18163 ( .A1(n15119), .A2(n16073), .ZN(n14961) );
  AOI211_X1 U18164 ( .C1(n14963), .C2(n16067), .A(n14962), .B(n14961), .ZN(
        n14964) );
  OAI21_X1 U18165 ( .B1(n15125), .B2(n16072), .A(n14964), .ZN(P2_U2988) );
  INV_X1 U18166 ( .A(n14966), .ZN(n14968) );
  AND2_X1 U18167 ( .A1(n14966), .A2(n14965), .ZN(n14967) );
  OAI22_X1 U18168 ( .A1(n14955), .A2(n14968), .B1(n9676), .B2(n14967), .ZN(
        n15135) );
  AOI21_X1 U18169 ( .B1(n15116), .B2(n14976), .A(n14969), .ZN(n15133) );
  NAND2_X1 U18170 ( .A1(n19011), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15127) );
  OAI21_X1 U18171 ( .B1(n16059), .B2(n14970), .A(n15127), .ZN(n14971) );
  AOI21_X1 U18172 ( .B1(n16052), .B2(n15959), .A(n14971), .ZN(n14972) );
  OAI21_X1 U18173 ( .B1(n15126), .B2(n19020), .A(n14972), .ZN(n14973) );
  AOI21_X1 U18174 ( .B1(n15133), .B2(n19015), .A(n14973), .ZN(n14974) );
  OAI21_X1 U18175 ( .B1(n15135), .B2(n16072), .A(n14974), .ZN(P2_U2989) );
  INV_X1 U18176 ( .A(n14975), .ZN(n14977) );
  OAI21_X1 U18177 ( .B1(n14977), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n14976), .ZN(n15144) );
  XNOR2_X1 U18178 ( .A(n14979), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14980) );
  XNOR2_X1 U18179 ( .A(n14978), .B(n14980), .ZN(n15136) );
  NAND2_X1 U18180 ( .A1(n15136), .A2(n19013), .ZN(n14986) );
  NAND2_X1 U18181 ( .A1(n19011), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15138) );
  NAND2_X1 U18182 ( .A1(n19012), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14981) );
  OAI211_X1 U18183 ( .C1(n19025), .C2(n14982), .A(n15138), .B(n14981), .ZN(
        n14983) );
  AOI21_X1 U18184 ( .B1(n14984), .B2(n16067), .A(n14983), .ZN(n14985) );
  OAI211_X1 U18185 ( .C1(n16073), .C2(n15144), .A(n14986), .B(n14985), .ZN(
        P2_U2990) );
  OAI21_X1 U18186 ( .B1(n14987), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n14975), .ZN(n15157) );
  XOR2_X1 U18187 ( .A(n14988), .B(n14989), .Z(n15145) );
  NAND2_X1 U18188 ( .A1(n15145), .A2(n19013), .ZN(n14995) );
  OAI22_X1 U18189 ( .A1(n16059), .A2(n14990), .B1(n10377), .B2(n18831), .ZN(
        n14992) );
  NOR2_X1 U18190 ( .A1(n15146), .A2(n19020), .ZN(n14991) );
  AOI211_X1 U18191 ( .C1(n16052), .C2(n14993), .A(n14992), .B(n14991), .ZN(
        n14994) );
  OAI211_X1 U18192 ( .C1(n16073), .C2(n15157), .A(n14995), .B(n14994), .ZN(
        P2_U2991) );
  OAI211_X1 U18193 ( .C1(n14997), .C2(n15285), .A(n14998), .B(n15266), .ZN(
        n15001) );
  INV_X1 U18194 ( .A(n14999), .ZN(n15000) );
  NAND3_X1 U18195 ( .A1(n15001), .A2(n15265), .A3(n15000), .ZN(n15004) );
  INV_X1 U18196 ( .A(n15229), .ZN(n15007) );
  INV_X1 U18197 ( .A(n15005), .ZN(n15006) );
  AOI21_X1 U18198 ( .B1(n15230), .B2(n15007), .A(n15006), .ZN(n15059) );
  INV_X1 U18199 ( .A(n15008), .ZN(n15009) );
  NOR2_X1 U18200 ( .A1(n15010), .A2(n15009), .ZN(n15060) );
  AOI21_X1 U18201 ( .B1(n15059), .B2(n15060), .A(n15010), .ZN(n15052) );
  NOR2_X1 U18202 ( .A1(n15052), .A2(n15050), .ZN(n15042) );
  INV_X1 U18203 ( .A(n15011), .ZN(n15040) );
  NAND2_X1 U18204 ( .A1(n15042), .A2(n15040), .ZN(n15028) );
  INV_X1 U18205 ( .A(n15029), .ZN(n15012) );
  AOI21_X1 U18206 ( .B1(n15028), .B2(n15013), .A(n15012), .ZN(n15018) );
  INV_X1 U18207 ( .A(n15014), .ZN(n15016) );
  NAND2_X1 U18208 ( .A1(n15016), .A2(n15015), .ZN(n15017) );
  XNOR2_X1 U18209 ( .A(n15018), .B(n15017), .ZN(n15170) );
  NAND2_X1 U18210 ( .A1(n19011), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15159) );
  OAI21_X1 U18211 ( .B1(n16059), .B2(n15019), .A(n15159), .ZN(n15022) );
  NOR2_X1 U18212 ( .A1(n15020), .A2(n19020), .ZN(n15021) );
  AOI211_X1 U18213 ( .C1(n16052), .C2(n15023), .A(n15022), .B(n15021), .ZN(
        n15026) );
  NAND2_X1 U18214 ( .A1(n15024), .A2(n9617), .ZN(n15158) );
  NAND3_X1 U18215 ( .A1(n16000), .A2(n19015), .A3(n15158), .ZN(n15025) );
  OAI211_X1 U18216 ( .C1(n15170), .C2(n16072), .A(n15026), .B(n15025), .ZN(
        P2_U2993) );
  NAND2_X1 U18217 ( .A1(n15028), .A2(n15027), .ZN(n15032) );
  NAND2_X1 U18218 ( .A1(n15030), .A2(n15029), .ZN(n15031) );
  XNOR2_X1 U18219 ( .A(n15032), .B(n15031), .ZN(n15183) );
  NAND2_X1 U18220 ( .A1(n12971), .A2(n15173), .ZN(n15055) );
  OAI21_X1 U18221 ( .B1(n15055), .B2(n15189), .A(n15172), .ZN(n15033) );
  AND2_X1 U18222 ( .A1(n15033), .A2(n15024), .ZN(n15181) );
  NOR2_X1 U18223 ( .A1(n18847), .A2(n19647), .ZN(n15176) );
  NOR2_X1 U18224 ( .A1(n19025), .A2(n15034), .ZN(n15035) );
  AOI211_X1 U18225 ( .C1(n19012), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15176), .B(n15035), .ZN(n15036) );
  OAI21_X1 U18226 ( .B1(n19020), .B2(n15174), .A(n15036), .ZN(n15037) );
  AOI21_X1 U18227 ( .B1(n15181), .B2(n19015), .A(n15037), .ZN(n15038) );
  OAI21_X1 U18228 ( .B1(n15183), .B2(n16072), .A(n15038), .ZN(P2_U2994) );
  NAND2_X1 U18229 ( .A1(n15040), .A2(n15039), .ZN(n15044) );
  INV_X1 U18230 ( .A(n15041), .ZN(n15049) );
  NOR2_X1 U18231 ( .A1(n15042), .A2(n15049), .ZN(n15043) );
  XOR2_X1 U18232 ( .A(n15044), .B(n15043), .Z(n15193) );
  XNOR2_X1 U18233 ( .A(n15055), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15191) );
  NAND2_X1 U18234 ( .A1(n19011), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15184) );
  OAI21_X1 U18235 ( .B1(n16059), .B2(n18685), .A(n15184), .ZN(n15045) );
  AOI21_X1 U18236 ( .B1(n18684), .B2(n16052), .A(n15045), .ZN(n15046) );
  OAI21_X1 U18237 ( .B1(n19020), .B2(n18689), .A(n15046), .ZN(n15047) );
  AOI21_X1 U18238 ( .B1(n15191), .B2(n19015), .A(n15047), .ZN(n15048) );
  OAI21_X1 U18239 ( .B1(n15193), .B2(n16072), .A(n15048), .ZN(P2_U2995) );
  NOR2_X1 U18240 ( .A1(n15050), .A2(n15049), .ZN(n15051) );
  XNOR2_X1 U18241 ( .A(n15052), .B(n15051), .ZN(n15210) );
  NAND2_X1 U18242 ( .A1(n19011), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n15199) );
  NAND2_X1 U18243 ( .A1(n19012), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15053) );
  OAI211_X1 U18244 ( .C1(n18695), .C2(n19025), .A(n15199), .B(n15053), .ZN(
        n15057) );
  INV_X1 U18245 ( .A(n15054), .ZN(n15201) );
  NOR2_X1 U18246 ( .A1(n15243), .A2(n15201), .ZN(n15065) );
  OAI21_X1 U18247 ( .B1(n15065), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15055), .ZN(n15194) );
  NOR2_X1 U18248 ( .A1(n15194), .A2(n16073), .ZN(n15056) );
  AOI211_X1 U18249 ( .C1(n16067), .C2(n18701), .A(n15057), .B(n15056), .ZN(
        n15058) );
  OAI21_X1 U18250 ( .B1(n15210), .B2(n16072), .A(n15058), .ZN(P2_U2996) );
  XOR2_X1 U18251 ( .A(n15060), .B(n15059), .Z(n15228) );
  NOR2_X1 U18252 ( .A1(n19641), .A2(n18831), .ZN(n15063) );
  INV_X1 U18253 ( .A(n18707), .ZN(n15061) );
  OAI22_X1 U18254 ( .A1(n16059), .A2(n18709), .B1(n19025), .B2(n15061), .ZN(
        n15062) );
  AOI211_X1 U18255 ( .C1(n16067), .C2(n18713), .A(n15063), .B(n15062), .ZN(
        n15068) );
  NAND2_X1 U18256 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15064) );
  NOR2_X1 U18257 ( .A1(n15243), .A2(n15064), .ZN(n16006) );
  INV_X1 U18258 ( .A(n15065), .ZN(n15066) );
  OAI211_X1 U18259 ( .C1(n16006), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15066), .B(n19015), .ZN(n15067) );
  OAI211_X1 U18260 ( .C1(n15228), .C2(n16072), .A(n15068), .B(n15067), .ZN(
        P2_U2997) );
  XNOR2_X1 U18261 ( .A(n15070), .B(n15069), .ZN(n15071) );
  XNOR2_X1 U18262 ( .A(n9653), .B(n15071), .ZN(n15374) );
  INV_X1 U18263 ( .A(n16063), .ZN(n15073) );
  NOR2_X1 U18264 ( .A1(n15073), .A2(n15072), .ZN(n15075) );
  XOR2_X1 U18265 ( .A(n15075), .B(n15074), .Z(n15372) );
  OAI22_X1 U18266 ( .A1(n16059), .A2(n15076), .B1(n10335), .B2(n18847), .ZN(
        n15077) );
  AOI21_X1 U18267 ( .B1(n16052), .B2(n18821), .A(n15077), .ZN(n15078) );
  OAI21_X1 U18268 ( .B1(n18825), .B2(n19020), .A(n15078), .ZN(n15079) );
  AOI21_X1 U18269 ( .B1(n15372), .B2(n19013), .A(n15079), .ZN(n15080) );
  OAI21_X1 U18270 ( .B1(n16073), .B2(n15374), .A(n15080), .ZN(P2_U3007) );
  INV_X1 U18271 ( .A(n15081), .ZN(n15083) );
  OAI21_X1 U18272 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15083), .A(
        n15082), .ZN(n15086) );
  OAI21_X1 U18273 ( .B1(n15090), .B2(n15405), .A(n15089), .ZN(P2_U3016) );
  OAI21_X1 U18274 ( .B1(n15092), .B2(n16097), .A(n15091), .ZN(n15099) );
  XNOR2_X1 U18275 ( .A(n15096), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15093) );
  NAND2_X1 U18276 ( .A1(n15094), .A2(n15093), .ZN(n15095) );
  OAI21_X1 U18277 ( .B1(n15097), .B2(n15096), .A(n15095), .ZN(n15098) );
  NOR2_X1 U18278 ( .A1(n15099), .A2(n15098), .ZN(n15100) );
  OAI21_X1 U18279 ( .B1(n15104), .B2(n15405), .A(n15103), .ZN(P2_U3017) );
  NAND2_X1 U18280 ( .A1(n15410), .A2(n15105), .ZN(n15106) );
  OAI211_X1 U18281 ( .C1(n15108), .C2(n15404), .A(n15107), .B(n15106), .ZN(
        n15109) );
  AOI211_X1 U18282 ( .C1(n15123), .C2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15110), .B(n15109), .ZN(n15113) );
  NAND2_X1 U18283 ( .A1(n15111), .A2(n16105), .ZN(n15112) );
  OAI211_X1 U18284 ( .C1(n15114), .C2(n15405), .A(n15113), .B(n15112), .ZN(
        P2_U3019) );
  INV_X1 U18285 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15115) );
  OAI21_X1 U18286 ( .B1(n15131), .B2(n15116), .A(n15115), .ZN(n15122) );
  AOI21_X1 U18287 ( .B1(n15410), .B2(n15951), .A(n15117), .ZN(n15118) );
  OAI21_X1 U18288 ( .B1(n15948), .B2(n15404), .A(n15118), .ZN(n15121) );
  NOR2_X1 U18289 ( .A1(n15119), .A2(n15413), .ZN(n15120) );
  AOI211_X1 U18290 ( .C1(n15123), .C2(n15122), .A(n15121), .B(n15120), .ZN(
        n15124) );
  OAI21_X1 U18291 ( .B1(n15125), .B2(n15405), .A(n15124), .ZN(P2_U3020) );
  NAND2_X1 U18292 ( .A1(n15141), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15130) );
  INV_X1 U18293 ( .A(n15126), .ZN(n15961) );
  OAI21_X1 U18294 ( .B1(n16097), .B2(n15964), .A(n15127), .ZN(n15128) );
  AOI21_X1 U18295 ( .B1(n15961), .B2(n16104), .A(n15128), .ZN(n15129) );
  OAI211_X1 U18296 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n15131), .A(
        n15130), .B(n15129), .ZN(n15132) );
  AOI21_X1 U18297 ( .B1(n15133), .B2(n16105), .A(n15132), .ZN(n15134) );
  OAI21_X1 U18298 ( .B1(n15135), .B2(n15405), .A(n15134), .ZN(P2_U3021) );
  NAND2_X1 U18299 ( .A1(n15136), .A2(n16102), .ZN(n15143) );
  INV_X1 U18300 ( .A(n16086), .ZN(n15147) );
  NOR4_X1 U18301 ( .A1(n15147), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15153), .A4(n16001), .ZN(n15140) );
  NAND2_X1 U18302 ( .A1(n15410), .A2(n15973), .ZN(n15137) );
  OAI211_X1 U18303 ( .C1(n15975), .C2(n15404), .A(n15138), .B(n15137), .ZN(
        n15139) );
  AOI211_X1 U18304 ( .C1(n15141), .C2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15140), .B(n15139), .ZN(n15142) );
  OAI211_X1 U18305 ( .C1(n15144), .C2(n15413), .A(n15143), .B(n15142), .ZN(
        P2_U3022) );
  NAND2_X1 U18306 ( .A1(n15145), .A2(n16102), .ZN(n15156) );
  NOR2_X1 U18307 ( .A1(n16001), .A2(n15147), .ZN(n15154) );
  NOR2_X1 U18308 ( .A1(n15146), .A2(n15404), .ZN(n15152) );
  OAI22_X1 U18309 ( .A1(n15315), .A2(n16081), .B1(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15147), .ZN(n15148) );
  AOI22_X1 U18310 ( .A1(n19011), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15148), .ZN(n15149) );
  OAI21_X1 U18311 ( .B1(n16097), .B2(n15150), .A(n15149), .ZN(n15151) );
  AOI211_X1 U18312 ( .C1(n15154), .C2(n15153), .A(n15152), .B(n15151), .ZN(
        n15155) );
  OAI211_X1 U18313 ( .C1(n15157), .C2(n15413), .A(n15156), .B(n15155), .ZN(
        P2_U3023) );
  NAND3_X1 U18314 ( .A1(n16000), .A2(n16105), .A3(n15158), .ZN(n15168) );
  OAI21_X1 U18315 ( .B1(n16097), .B2(n15160), .A(n15159), .ZN(n15161) );
  AOI21_X1 U18316 ( .B1(n15162), .B2(n16104), .A(n15161), .ZN(n15167) );
  OAI21_X1 U18317 ( .B1(n15164), .B2(n15367), .A(n15316), .ZN(n15163) );
  NAND2_X1 U18318 ( .A1(n15163), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15166) );
  NAND3_X1 U18319 ( .A1(n15349), .A2(n15164), .A3(n9617), .ZN(n15165) );
  AND4_X1 U18320 ( .A1(n15168), .A2(n15167), .A3(n15166), .A4(n15165), .ZN(
        n15169) );
  OAI21_X1 U18321 ( .B1(n15170), .B2(n15405), .A(n15169), .ZN(P2_U3025) );
  AOI21_X1 U18322 ( .B1(n15171), .B2(n15366), .A(n15215), .ZN(n15206) );
  NOR2_X1 U18323 ( .A1(n15206), .A2(n15172), .ZN(n15180) );
  XNOR2_X1 U18324 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15178) );
  NAND2_X1 U18325 ( .A1(n15349), .A2(n15173), .ZN(n15185) );
  NOR2_X1 U18326 ( .A1(n15174), .A2(n15404), .ZN(n15175) );
  AOI211_X1 U18327 ( .C1(n15410), .C2(n15983), .A(n15176), .B(n15175), .ZN(
        n15177) );
  OAI21_X1 U18328 ( .B1(n15178), .B2(n15185), .A(n15177), .ZN(n15179) );
  AOI211_X1 U18329 ( .C1(n15181), .C2(n16105), .A(n15180), .B(n15179), .ZN(
        n15182) );
  OAI21_X1 U18330 ( .B1(n15183), .B2(n15405), .A(n15182), .ZN(P2_U3026) );
  OAI21_X1 U18331 ( .B1(n18689), .B2(n15404), .A(n15184), .ZN(n15187) );
  NOR2_X1 U18332 ( .A1(n15185), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15186) );
  AOI211_X1 U18333 ( .C1(n15410), .C2(n10069), .A(n15187), .B(n15186), .ZN(
        n15188) );
  OAI21_X1 U18334 ( .B1(n15206), .B2(n15189), .A(n15188), .ZN(n15190) );
  AOI21_X1 U18335 ( .B1(n15191), .B2(n16105), .A(n15190), .ZN(n15192) );
  OAI21_X1 U18336 ( .B1(n15193), .B2(n15405), .A(n15192), .ZN(P2_U3027) );
  INV_X1 U18337 ( .A(n15194), .ZN(n15208) );
  AND2_X1 U18338 ( .A1(n15196), .A2(n15195), .ZN(n15197) );
  NOR2_X1 U18339 ( .A1(n15198), .A2(n15197), .ZN(n18700) );
  INV_X1 U18340 ( .A(n18700), .ZN(n15200) );
  OAI21_X1 U18341 ( .B1(n16097), .B2(n15200), .A(n15199), .ZN(n15203) );
  NOR3_X1 U18342 ( .A1(n15219), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15201), .ZN(n15202) );
  AOI211_X1 U18343 ( .C1(n18701), .C2(n16104), .A(n15203), .B(n15202), .ZN(
        n15204) );
  OAI21_X1 U18344 ( .B1(n15206), .B2(n15205), .A(n15204), .ZN(n15207) );
  AOI21_X1 U18345 ( .B1(n15208), .B2(n16105), .A(n15207), .ZN(n15209) );
  OAI21_X1 U18346 ( .B1(n15210), .B2(n15405), .A(n15209), .ZN(P2_U3028) );
  NOR2_X1 U18347 ( .A1(n15211), .A2(n16105), .ZN(n15212) );
  OR2_X1 U18348 ( .A1(n16006), .A2(n15212), .ZN(n15217) );
  NOR2_X1 U18349 ( .A1(n15213), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15214) );
  NOR2_X1 U18350 ( .A1(n15215), .A2(n15214), .ZN(n15216) );
  NAND2_X1 U18351 ( .A1(n15217), .A2(n15216), .ZN(n15239) );
  NOR2_X1 U18352 ( .A1(n15367), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15218) );
  OR2_X1 U18353 ( .A1(n15239), .A2(n15218), .ZN(n15226) );
  OAI21_X1 U18354 ( .B1(n15243), .B2(n15413), .A(n15219), .ZN(n15220) );
  NAND2_X1 U18355 ( .A1(n15220), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15236) );
  NAND2_X1 U18356 ( .A1(n15221), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15224) );
  AOI22_X1 U18357 ( .A1(n18713), .A2(n16104), .B1(P2_REIP_REG_17__SCAN_IN), 
        .B2(n19011), .ZN(n15223) );
  NAND2_X1 U18358 ( .A1(n15410), .A2(n18714), .ZN(n15222) );
  OAI211_X1 U18359 ( .C1(n15236), .C2(n15224), .A(n15223), .B(n15222), .ZN(
        n15225) );
  AOI21_X1 U18360 ( .B1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n15226), .A(
        n15225), .ZN(n15227) );
  OAI21_X1 U18361 ( .B1(n15228), .B2(n15405), .A(n15227), .ZN(P2_U3029) );
  XNOR2_X1 U18362 ( .A(n15230), .B(n15229), .ZN(n16010) );
  INV_X1 U18363 ( .A(n16010), .ZN(n15241) );
  OR2_X1 U18364 ( .A1(n15232), .A2(n15231), .ZN(n15234) );
  AND2_X1 U18365 ( .A1(n15234), .A2(n15233), .ZN(n18912) );
  AOI22_X1 U18366 ( .A1(n15410), .A2(n18912), .B1(P2_REIP_REG_16__SCAN_IN), 
        .B2(n19011), .ZN(n15235) );
  OAI21_X1 U18367 ( .B1(n15404), .B2(n18727), .A(n15235), .ZN(n15238) );
  NOR2_X1 U18368 ( .A1(n15236), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15237) );
  AOI211_X1 U18369 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15239), .A(
        n15238), .B(n15237), .ZN(n15240) );
  OAI21_X1 U18370 ( .B1(n15241), .B2(n15405), .A(n15240), .ZN(P2_U3030) );
  NAND2_X1 U18371 ( .A1(n12971), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15341) );
  NAND2_X1 U18372 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15312) );
  INV_X1 U18373 ( .A(n15243), .ZN(n16005) );
  AOI21_X1 U18374 ( .B1(n15269), .B2(n15244), .A(n16005), .ZN(n16020) );
  INV_X1 U18375 ( .A(n16020), .ZN(n15263) );
  AND2_X1 U18376 ( .A1(n15246), .A2(n15245), .ZN(n15247) );
  OR2_X1 U18377 ( .A1(n15248), .A2(n15247), .ZN(n16019) );
  NAND2_X1 U18378 ( .A1(n16019), .A2(n16102), .ZN(n15262) );
  INV_X1 U18379 ( .A(n18751), .ZN(n15260) );
  INV_X1 U18380 ( .A(n15272), .ZN(n15249) );
  OR2_X1 U18381 ( .A1(n15250), .A2(n15249), .ZN(n15252) );
  INV_X1 U18382 ( .A(n12980), .ZN(n15251) );
  NAND2_X1 U18383 ( .A1(n15252), .A2(n15251), .ZN(n18923) );
  OAI22_X1 U18384 ( .A1(n16097), .A2(n18923), .B1(n10729), .B2(n18847), .ZN(
        n15259) );
  NAND2_X1 U18385 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15254) );
  INV_X1 U18386 ( .A(n15275), .ZN(n15253) );
  NOR2_X1 U18387 ( .A1(n15254), .A2(n15253), .ZN(n15257) );
  NAND2_X1 U18388 ( .A1(n15275), .A2(n15300), .ZN(n15294) );
  NAND2_X1 U18389 ( .A1(n15296), .A2(n15294), .ZN(n15276) );
  AOI21_X1 U18390 ( .B1(n15275), .B2(n15274), .A(n15276), .ZN(n15255) );
  INV_X1 U18391 ( .A(n15255), .ZN(n15256) );
  MUX2_X1 U18392 ( .A(n15257), .B(n15256), .S(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n15258) );
  AOI211_X1 U18393 ( .C1(n15260), .C2(n16104), .A(n15259), .B(n15258), .ZN(
        n15261) );
  OAI211_X1 U18394 ( .C1(n15263), .C2(n15413), .A(n15262), .B(n15261), .ZN(
        P2_U3032) );
  INV_X1 U18395 ( .A(n15266), .ZN(n15268) );
  AND2_X1 U18396 ( .A1(n15266), .A2(n15265), .ZN(n15267) );
  OAI22_X1 U18397 ( .A1(n12966), .A2(n15268), .B1(n15264), .B2(n15267), .ZN(
        n16027) );
  NOR2_X1 U18398 ( .A1(n15300), .A2(n15305), .ZN(n15301) );
  INV_X1 U18399 ( .A(n16029), .ZN(n18757) );
  OAI22_X1 U18400 ( .A1(n15413), .A2(n16026), .B1(n15404), .B2(n18757), .ZN(
        n15281) );
  OR2_X1 U18401 ( .A1(n15271), .A2(n15270), .ZN(n15273) );
  NAND2_X1 U18402 ( .A1(n15273), .A2(n15272), .ZN(n18925) );
  AND2_X1 U18403 ( .A1(n15275), .A2(n15274), .ZN(n15277) );
  AOI22_X1 U18404 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15277), .B1(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15276), .ZN(n15279) );
  OR2_X1 U18405 ( .A1(n10711), .A2(n18847), .ZN(n15278) );
  OAI211_X1 U18406 ( .C1(n16097), .C2(n18925), .A(n15279), .B(n15278), .ZN(
        n15280) );
  NOR2_X1 U18407 ( .A1(n15281), .A2(n15280), .ZN(n15282) );
  OAI21_X1 U18408 ( .B1(n16027), .B2(n15405), .A(n15282), .ZN(P2_U3033) );
  NAND2_X1 U18409 ( .A1(n14997), .A2(n15283), .ZN(n15288) );
  INV_X1 U18410 ( .A(n15284), .ZN(n15286) );
  OR2_X1 U18411 ( .A1(n15286), .A2(n15285), .ZN(n15287) );
  XNOR2_X1 U18412 ( .A(n15288), .B(n15287), .ZN(n16033) );
  INV_X1 U18413 ( .A(n16033), .ZN(n15304) );
  INV_X1 U18414 ( .A(n18772), .ZN(n15299) );
  INV_X1 U18415 ( .A(n15289), .ZN(n15290) );
  OR2_X1 U18416 ( .A1(n15291), .A2(n15290), .ZN(n15293) );
  INV_X1 U18417 ( .A(n15270), .ZN(n15292) );
  NAND2_X1 U18418 ( .A1(n15293), .A2(n15292), .ZN(n18928) );
  NAND2_X1 U18419 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19011), .ZN(n15295) );
  OAI211_X1 U18420 ( .C1(n16097), .C2(n18928), .A(n15295), .B(n15294), .ZN(
        n15298) );
  NOR2_X1 U18421 ( .A1(n15296), .A2(n15300), .ZN(n15297) );
  AOI211_X1 U18422 ( .C1(n15299), .C2(n16104), .A(n15298), .B(n15297), .ZN(
        n15303) );
  NAND2_X1 U18423 ( .A1(n15305), .A2(n15300), .ZN(n16035) );
  INV_X1 U18424 ( .A(n15301), .ZN(n16034) );
  NAND3_X1 U18425 ( .A1(n16035), .A2(n16105), .A3(n16034), .ZN(n15302) );
  OAI211_X1 U18426 ( .C1(n15304), .C2(n15405), .A(n15303), .B(n15302), .ZN(
        P2_U3034) );
  NOR2_X1 U18427 ( .A1(n15341), .A2(n15333), .ZN(n15323) );
  OAI21_X1 U18428 ( .B1(n15323), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15305), .ZN(n16042) );
  NAND2_X1 U18429 ( .A1(n15306), .A2(n10093), .ZN(n15311) );
  INV_X1 U18430 ( .A(n15307), .ZN(n15308) );
  NOR2_X1 U18431 ( .A1(n15309), .A2(n15308), .ZN(n15310) );
  XNOR2_X1 U18432 ( .A(n15311), .B(n15310), .ZN(n16041) );
  AND2_X1 U18433 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15349), .ZN(
        n15334) );
  OAI211_X1 U18434 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n15334), .B(n15312), .ZN(
        n15320) );
  OAI21_X1 U18435 ( .B1(n15314), .B2(n15313), .A(n15289), .ZN(n18930) );
  AOI21_X1 U18436 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15316), .A(
        n15315), .ZN(n15335) );
  AOI22_X1 U18437 ( .A1(n19011), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15335), .ZN(n15317) );
  OAI21_X1 U18438 ( .B1(n16097), .B2(n18930), .A(n15317), .ZN(n15318) );
  AOI21_X1 U18439 ( .B1(n16104), .B2(n18773), .A(n15318), .ZN(n15319) );
  OAI211_X1 U18440 ( .C1(n16041), .C2(n15405), .A(n15320), .B(n15319), .ZN(
        n15321) );
  INV_X1 U18441 ( .A(n15321), .ZN(n15322) );
  OAI21_X1 U18442 ( .B1(n16042), .B2(n15413), .A(n15322), .ZN(P2_U3035) );
  AOI21_X1 U18443 ( .B1(n15333), .B2(n15341), .A(n15323), .ZN(n16047) );
  INV_X1 U18444 ( .A(n16047), .ZN(n15340) );
  NAND2_X1 U18445 ( .A1(n15325), .A2(n15324), .ZN(n15329) );
  INV_X1 U18446 ( .A(n15327), .ZN(n15344) );
  NOR2_X1 U18447 ( .A1(n15326), .A2(n15344), .ZN(n15328) );
  XOR2_X1 U18448 ( .A(n15329), .B(n15328), .Z(n16049) );
  INV_X1 U18449 ( .A(n15352), .ZN(n15330) );
  XNOR2_X1 U18450 ( .A(n15331), .B(n15330), .ZN(n18933) );
  NOR2_X1 U18451 ( .A1(n10659), .A2(n18847), .ZN(n15332) );
  AOI221_X1 U18452 ( .B1(n15335), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), 
        .C1(n15334), .C2(n15333), .A(n15332), .ZN(n15337) );
  INV_X1 U18453 ( .A(n18793), .ZN(n16048) );
  NAND2_X1 U18454 ( .A1(n16104), .A2(n16048), .ZN(n15336) );
  OAI211_X1 U18455 ( .C1(n16097), .C2(n18933), .A(n15337), .B(n15336), .ZN(
        n15338) );
  AOI21_X1 U18456 ( .B1(n16049), .B2(n16102), .A(n15338), .ZN(n15339) );
  OAI21_X1 U18457 ( .B1(n15340), .B2(n15413), .A(n15339), .ZN(P2_U3036) );
  OAI21_X1 U18458 ( .B1(n12971), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15341), .ZN(n16054) );
  OR2_X1 U18459 ( .A1(n15344), .A2(n15343), .ZN(n15345) );
  XNOR2_X1 U18460 ( .A(n15342), .B(n15345), .ZN(n16053) );
  NOR2_X1 U18461 ( .A1(n10638), .A2(n18847), .ZN(n15346) );
  AOI221_X1 U18462 ( .B1(n15349), .B2(n15348), .C1(n15347), .C2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15346), .ZN(n15357) );
  INV_X1 U18463 ( .A(n18806), .ZN(n15354) );
  OR2_X1 U18464 ( .A1(n15351), .A2(n15350), .ZN(n15353) );
  NAND2_X1 U18465 ( .A1(n15353), .A2(n15352), .ZN(n18936) );
  OAI22_X1 U18466 ( .A1(n15404), .A2(n15354), .B1(n16097), .B2(n18936), .ZN(
        n15355) );
  INV_X1 U18467 ( .A(n15355), .ZN(n15356) );
  OAI211_X1 U18468 ( .C1(n16053), .C2(n15405), .A(n15357), .B(n15356), .ZN(
        n15358) );
  INV_X1 U18469 ( .A(n15358), .ZN(n15359) );
  OAI21_X1 U18470 ( .B1(n16054), .B2(n15413), .A(n15359), .ZN(P2_U3037) );
  NAND2_X1 U18471 ( .A1(n15396), .A2(n15402), .ZN(n15384) );
  NOR3_X1 U18472 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n15383), .A3(
        n15384), .ZN(n16108) );
  OR2_X1 U18473 ( .A1(n15361), .A2(n15360), .ZN(n15363) );
  NAND2_X1 U18474 ( .A1(n15363), .A2(n15362), .ZN(n18941) );
  AOI21_X1 U18475 ( .B1(n15366), .B2(n15365), .A(n15364), .ZN(n15382) );
  OAI21_X1 U18476 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15367), .A(
        n15382), .ZN(n16107) );
  NAND2_X1 U18477 ( .A1(n16107), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15370) );
  INV_X1 U18478 ( .A(n18825), .ZN(n15368) );
  AOI22_X1 U18479 ( .A1(n15368), .A2(n16104), .B1(n19011), .B2(
        P2_REIP_REG_7__SCAN_IN), .ZN(n15369) );
  OAI211_X1 U18480 ( .C1(n16097), .C2(n18941), .A(n15370), .B(n15369), .ZN(
        n15371) );
  AOI211_X1 U18481 ( .C1(n15372), .C2(n16102), .A(n16108), .B(n15371), .ZN(
        n15373) );
  OAI21_X1 U18482 ( .B1(n15413), .B2(n15374), .A(n15373), .ZN(P2_U3039) );
  OR2_X1 U18483 ( .A1(n15377), .A2(n15376), .ZN(n15378) );
  NAND2_X1 U18484 ( .A1(n15375), .A2(n15378), .ZN(n16071) );
  OAI21_X1 U18485 ( .B1(n15380), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15379), .ZN(n16074) );
  OR2_X1 U18486 ( .A1(n16074), .A2(n15413), .ZN(n15392) );
  NAND2_X1 U18487 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n19011), .ZN(n15381) );
  OAI221_X1 U18488 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15384), .C1(
        n15383), .C2(n15382), .A(n15381), .ZN(n15390) );
  INV_X1 U18489 ( .A(n15385), .ZN(n15386) );
  XNOR2_X1 U18490 ( .A(n15387), .B(n15386), .ZN(n18942) );
  NAND2_X1 U18491 ( .A1(n18942), .A2(n15410), .ZN(n15388) );
  OAI21_X1 U18492 ( .B1(n15404), .B2(n18841), .A(n15388), .ZN(n15389) );
  NOR2_X1 U18493 ( .A1(n15390), .A2(n15389), .ZN(n15391) );
  OAI211_X1 U18494 ( .C1(n16071), .C2(n15405), .A(n15392), .B(n15391), .ZN(
        P2_U3040) );
  OAI21_X1 U18495 ( .B1(n15395), .B2(n15394), .A(n15393), .ZN(n18950) );
  INV_X1 U18496 ( .A(n18950), .ZN(n15409) );
  AOI21_X1 U18497 ( .B1(n15398), .B2(n15397), .A(n15396), .ZN(n15401) );
  OAI22_X1 U18498 ( .A1(n15399), .A2(n15398), .B1(n10328), .B2(n18847), .ZN(
        n15400) );
  AOI21_X1 U18499 ( .B1(n15402), .B2(n15401), .A(n15400), .ZN(n15403) );
  OAI21_X1 U18500 ( .B1(n18850), .B2(n15404), .A(n15403), .ZN(n15408) );
  NOR2_X1 U18501 ( .A1(n15406), .A2(n15405), .ZN(n15407) );
  AOI211_X1 U18502 ( .C1(n15410), .C2(n15409), .A(n15408), .B(n15407), .ZN(
        n15411) );
  OAI21_X1 U18503 ( .B1(n15413), .B2(n15412), .A(n15411), .ZN(P2_U3041) );
  NAND2_X1 U18504 ( .A1(n15414), .A2(n12551), .ZN(n15424) );
  AND2_X1 U18505 ( .A1(n15424), .A2(n15415), .ZN(n15416) );
  AOI21_X1 U18506 ( .B1(n12601), .B2(n16114), .A(n15416), .ZN(n16147) );
  OAI22_X1 U18507 ( .A1(n9828), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n18898), .B2(n18865), .ZN(n15417) );
  INV_X1 U18508 ( .A(n15417), .ZN(n15423) );
  OAI222_X1 U18509 ( .A1(n19678), .A2(n12605), .B1(n16147), .B2(n19685), .C1(
        n19601), .C2(n15423), .ZN(n15419) );
  INV_X1 U18510 ( .A(n16145), .ZN(n15436) );
  OAI21_X1 U18511 ( .B1(n15436), .B2(n19685), .A(n19679), .ZN(n15418) );
  AOI22_X1 U18512 ( .A1(n15419), .A2(n19679), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15418), .ZN(n15420) );
  INV_X1 U18513 ( .A(n15420), .ZN(P2_U3601) );
  INV_X1 U18514 ( .A(n19678), .ZN(n15429) );
  AOI211_X1 U18515 ( .C1(n18898), .C2(n15422), .A(n18865), .B(n15421), .ZN(
        n18883) );
  AOI21_X1 U18516 ( .B1(n18865), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n18883), .ZN(n19676) );
  NAND2_X1 U18517 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15423), .ZN(n19675) );
  INV_X1 U18518 ( .A(n19675), .ZN(n15428) );
  NAND2_X1 U18519 ( .A1(n18872), .A2(n16114), .ZN(n15427) );
  OAI21_X1 U18520 ( .B1(n10435), .B2(n15425), .A(n15424), .ZN(n15426) );
  OAI211_X1 U18521 ( .C1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n15436), .A(
        n15427), .B(n15426), .ZN(n16151) );
  AOI222_X1 U18522 ( .A1(n19706), .A2(n15429), .B1(n19676), .B2(n15428), .C1(
        n16151), .C2(n19600), .ZN(n15432) );
  NAND2_X1 U18523 ( .A1(n15431), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15430) );
  OAI21_X1 U18524 ( .B1(n15432), .B2(n15431), .A(n15430), .ZN(P2_U3600) );
  NAND2_X1 U18525 ( .A1(n15433), .A2(n16114), .ZN(n15444) );
  INV_X1 U18526 ( .A(n15434), .ZN(n16134) );
  NOR2_X1 U18527 ( .A1(n16130), .A2(n16134), .ZN(n16119) );
  NOR2_X1 U18528 ( .A1(n10437), .A2(n19681), .ZN(n16116) );
  INV_X1 U18529 ( .A(n15435), .ZN(n15437) );
  OAI22_X1 U18530 ( .A1(n16119), .A2(n16116), .B1(n15436), .B2(n15437), .ZN(
        n15441) );
  NAND2_X1 U18531 ( .A1(n16145), .A2(n15437), .ZN(n16123) );
  NAND2_X1 U18532 ( .A1(n15438), .A2(n9620), .ZN(n15439) );
  NAND2_X1 U18533 ( .A1(n15439), .A2(n16121), .ZN(n16122) );
  NAND3_X1 U18534 ( .A1(n16120), .A2(n16123), .A3(n16122), .ZN(n15440) );
  MUX2_X1 U18535 ( .A(n15441), .B(n15440), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n15442) );
  NOR2_X1 U18536 ( .A1(n15442), .A2(n10522), .ZN(n15443) );
  NAND2_X1 U18537 ( .A1(n15444), .A2(n15443), .ZN(n16113) );
  NAND2_X1 U18538 ( .A1(n16113), .A2(n19600), .ZN(n15445) );
  OAI21_X1 U18539 ( .B1(n19304), .B2(n19678), .A(n15445), .ZN(n15446) );
  MUX2_X1 U18540 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15446), .S(
        n19679), .Z(P2_U3596) );
  AOI22_X1 U18541 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15450) );
  AOI22_X1 U18542 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15449) );
  AOI22_X1 U18543 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15448) );
  AOI22_X1 U18544 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15510), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15447) );
  NAND4_X1 U18545 ( .A1(n15450), .A2(n15449), .A3(n15448), .A4(n15447), .ZN(
        n15456) );
  AOI22_X1 U18546 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15454) );
  AOI22_X1 U18547 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15453) );
  AOI22_X1 U18548 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n16952), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15452) );
  AOI22_X1 U18549 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15451) );
  NAND4_X1 U18550 ( .A1(n15454), .A2(n15453), .A3(n15452), .A4(n15451), .ZN(
        n15455) );
  NOR2_X1 U18551 ( .A1(n15456), .A2(n15455), .ZN(n16738) );
  AOI22_X1 U18552 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16929), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15460) );
  AOI22_X1 U18553 ( .A1(n16883), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15459) );
  AOI22_X1 U18554 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15458) );
  AOI22_X1 U18555 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15510), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15457) );
  NAND4_X1 U18556 ( .A1(n15460), .A2(n15459), .A3(n15458), .A4(n15457), .ZN(
        n15466) );
  AOI22_X1 U18557 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15464) );
  AOI22_X1 U18558 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15463) );
  AOI22_X1 U18559 ( .A1(n10890), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15462) );
  AOI22_X1 U18560 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15461) );
  NAND4_X1 U18561 ( .A1(n15464), .A2(n15463), .A3(n15462), .A4(n15461), .ZN(
        n15465) );
  NOR2_X1 U18562 ( .A1(n15466), .A2(n15465), .ZN(n16756) );
  AOI22_X1 U18563 ( .A1(n15523), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15470) );
  AOI22_X1 U18564 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15469) );
  AOI22_X1 U18565 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15468) );
  AOI22_X1 U18566 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15510), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15467) );
  NAND4_X1 U18567 ( .A1(n15470), .A2(n15469), .A3(n15468), .A4(n15467), .ZN(
        n15476) );
  AOI22_X1 U18568 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15474) );
  AOI22_X1 U18569 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16844), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15473) );
  AOI22_X1 U18570 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15472) );
  AOI22_X1 U18571 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15471) );
  NAND4_X1 U18572 ( .A1(n15474), .A2(n15473), .A3(n15472), .A4(n15471), .ZN(
        n15475) );
  NOR2_X1 U18573 ( .A1(n15476), .A2(n15475), .ZN(n16749) );
  AOI22_X1 U18574 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15480) );
  AOI22_X1 U18575 ( .A1(n10890), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15479) );
  AOI22_X1 U18576 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15478) );
  AOI22_X1 U18577 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15510), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15477) );
  NAND4_X1 U18578 ( .A1(n15480), .A2(n15479), .A3(n15478), .A4(n15477), .ZN(
        n15486) );
  AOI22_X1 U18579 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15484) );
  AOI22_X1 U18580 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n15483) );
  AOI22_X1 U18581 ( .A1(n16839), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n15482) );
  AOI22_X1 U18582 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15481) );
  NAND4_X1 U18583 ( .A1(n15484), .A2(n15483), .A3(n15482), .A4(n15481), .ZN(
        n15485) );
  OR2_X1 U18584 ( .A1(n15486), .A2(n15485), .ZN(n16761) );
  AOI22_X1 U18585 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15497) );
  AOI22_X1 U18586 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15496) );
  AOI22_X1 U18587 ( .A1(n16955), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15487) );
  OAI21_X1 U18588 ( .B1(n15488), .B2(n16949), .A(n15487), .ZN(n15494) );
  AOI22_X1 U18589 ( .A1(n16839), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15492) );
  AOI22_X1 U18590 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15491) );
  AOI22_X1 U18591 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15490) );
  AOI22_X1 U18592 ( .A1(n10890), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15510), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15489) );
  NAND4_X1 U18593 ( .A1(n15492), .A2(n15491), .A3(n15490), .A4(n15489), .ZN(
        n15493) );
  AOI211_X1 U18594 ( .C1(n16929), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n15494), .B(n15493), .ZN(n15495) );
  NAND3_X1 U18595 ( .A1(n15497), .A2(n15496), .A3(n15495), .ZN(n16767) );
  AOI22_X1 U18596 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15507) );
  AOI22_X1 U18597 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16952), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15506) );
  AOI22_X1 U18598 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n16955), .B1(
        n15510), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15498) );
  OAI21_X1 U18599 ( .B1(n20770), .B2(n10809), .A(n15498), .ZN(n15504) );
  AOI22_X1 U18600 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n15523), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n16947), .ZN(n15502) );
  AOI22_X1 U18601 ( .A1(n16839), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15501) );
  AOI22_X1 U18602 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n16844), .B1(
        n10890), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15500) );
  AOI22_X1 U18603 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n16883), .ZN(n15499) );
  NAND4_X1 U18604 ( .A1(n15502), .A2(n15501), .A3(n15500), .A4(n15499), .ZN(
        n15503) );
  AOI211_X1 U18605 ( .C1(n16945), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n15504), .B(n15503), .ZN(n15505) );
  NAND3_X1 U18606 ( .A1(n15507), .A2(n15506), .A3(n15505), .ZN(n16768) );
  NAND2_X1 U18607 ( .A1(n16767), .A2(n16768), .ZN(n16766) );
  INV_X1 U18608 ( .A(n16766), .ZN(n16762) );
  NAND2_X1 U18609 ( .A1(n16761), .A2(n16762), .ZN(n16760) );
  NOR3_X1 U18610 ( .A1(n16756), .A2(n16749), .A3(n16760), .ZN(n17023) );
  AOI22_X1 U18611 ( .A1(n16839), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15519) );
  AOI22_X1 U18612 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15518) );
  AOI22_X1 U18613 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15508) );
  OAI21_X1 U18614 ( .B1(n15509), .B2(n20846), .A(n15508), .ZN(n15516) );
  AOI22_X1 U18615 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16844), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15514) );
  AOI22_X1 U18616 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15513) );
  AOI22_X1 U18617 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15512) );
  AOI22_X1 U18618 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15510), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15511) );
  NAND4_X1 U18619 ( .A1(n15514), .A2(n15513), .A3(n15512), .A4(n15511), .ZN(
        n15515) );
  AOI211_X1 U18620 ( .C1(n16927), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n15516), .B(n15515), .ZN(n15517) );
  NAND3_X1 U18621 ( .A1(n15519), .A2(n15518), .A3(n15517), .ZN(n17022) );
  NAND2_X1 U18622 ( .A1(n17023), .A2(n17022), .ZN(n17021) );
  XNOR2_X1 U18623 ( .A(n16738), .B(n17021), .ZN(n17020) );
  AND2_X1 U18624 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16742) );
  NAND2_X1 U18625 ( .A1(n18024), .A2(n16994), .ZN(n17000) );
  INV_X1 U18626 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n16836) );
  INV_X1 U18627 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n16854) );
  NOR2_X2 U18628 ( .A1(n17092), .A2(n16783), .ZN(n16808) );
  NAND2_X1 U18629 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16808), .ZN(n16754) );
  INV_X1 U18630 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16416) );
  INV_X1 U18631 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16438) );
  NOR2_X1 U18632 ( .A1(n16416), .A2(n16438), .ZN(n15520) );
  NAND4_X1 U18633 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .A4(n15520), .ZN(n16707) );
  NAND2_X1 U18634 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16758), .ZN(n16748) );
  NAND2_X1 U18635 ( .A1(n16980), .A2(n16748), .ZN(n16746) );
  OAI21_X1 U18636 ( .B1(n16742), .B2(n17000), .A(n16746), .ZN(n16743) );
  INV_X1 U18637 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16747) );
  NOR3_X1 U18638 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16747), .A3(n16748), .ZN(
        n15521) );
  AOI21_X1 U18639 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n16743), .A(n15521), .ZN(
        n15522) );
  OAI21_X1 U18640 ( .B1(n16980), .B2(n17020), .A(n15522), .ZN(P3_U2675) );
  AOI22_X1 U18641 ( .A1(n16946), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15534) );
  AOI22_X1 U18642 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15533) );
  INV_X1 U18643 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n20847) );
  AOI22_X1 U18644 ( .A1(n16928), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15524) );
  OAI21_X1 U18645 ( .B1(n9695), .B2(n20847), .A(n15524), .ZN(n15531) );
  AOI22_X1 U18646 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15529) );
  AOI22_X1 U18647 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15528) );
  AOI22_X1 U18648 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16844), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15527) );
  AOI22_X1 U18649 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15526) );
  NAND4_X1 U18650 ( .A1(n15529), .A2(n15528), .A3(n15527), .A4(n15526), .ZN(
        n15530) );
  AOI211_X1 U18651 ( .C1(n16962), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n15531), .B(n15530), .ZN(n15532) );
  NAND3_X1 U18652 ( .A1(n15534), .A2(n15533), .A3(n15532), .ZN(n17100) );
  INV_X1 U18653 ( .A(n17100), .ZN(n15537) );
  OAI211_X1 U18654 ( .C1(n16895), .C2(P3_EBX_REG_13__SCAN_IN), .A(n16980), .B(
        n15535), .ZN(n15536) );
  OAI21_X1 U18655 ( .B1(n15537), .B2(n16980), .A(n15536), .ZN(P3_U2690) );
  AOI221_X1 U18656 ( .B1(n10936), .B2(n17955), .C1(n20801), .C2(n17955), .A(
        n15538), .ZN(n15544) );
  NOR2_X1 U18657 ( .A1(n15540), .A2(n15539), .ZN(n15541) );
  XOR2_X1 U18658 ( .A(n16193), .B(n15541), .Z(n16203) );
  AOI22_X1 U18659 ( .A1(n17872), .A2(n16203), .B1(n16193), .B2(n15542), .ZN(
        n15543) );
  NAND2_X1 U18660 ( .A1(n17965), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16197) );
  OAI211_X1 U18661 ( .C1(n15544), .C2(n16193), .A(n15543), .B(n16197), .ZN(
        P3_U2833) );
  OAI211_X1 U18662 ( .C1(n15547), .C2(n15546), .A(n15545), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n15550) );
  INV_X1 U18663 ( .A(n15548), .ZN(n15549) );
  OAI21_X1 U18664 ( .B1(n20327), .B2(n15550), .A(n15549), .ZN(n15552) );
  NAND2_X1 U18665 ( .A1(n15550), .A2(n20327), .ZN(n15551) );
  OAI21_X1 U18666 ( .B1(n15553), .B2(n15552), .A(n15551), .ZN(n15554) );
  AOI222_X1 U18667 ( .A1(n15555), .A2(n20407), .B1(n15555), .B2(n15554), .C1(
        n20407), .C2(n15554), .ZN(n15557) );
  AOI21_X1 U18668 ( .B1(n15557), .B2(n15556), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n15559) );
  NOR2_X1 U18669 ( .A1(n15557), .A2(n15556), .ZN(n15558) );
  OAI21_X1 U18670 ( .B1(n15559), .B2(n15558), .A(n20000), .ZN(n15568) );
  NOR2_X1 U18671 ( .A1(P1_MORE_REG_SCAN_IN), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(
        n15563) );
  OAI211_X1 U18672 ( .C1(n15563), .C2(n15562), .A(n15561), .B(n15560), .ZN(
        n15564) );
  INV_X1 U18673 ( .A(n15564), .ZN(n15566) );
  NAND4_X1 U18674 ( .A1(n15568), .A2(n15567), .A3(n15566), .A4(n15565), .ZN(
        n15576) );
  NOR2_X1 U18675 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20581), .ZN(n15569) );
  AND2_X1 U18676 ( .A1(n20585), .A2(n15569), .ZN(n15574) );
  NAND4_X1 U18677 ( .A1(n13378), .A2(n15572), .A3(n15571), .A4(n15570), .ZN(
        n15573) );
  OAI21_X1 U18678 ( .B1(n15577), .B2(n15574), .A(n15573), .ZN(n15917) );
  AOI221_X1 U18679 ( .B1(n20578), .B2(n20577), .C1(n15576), .C2(n20577), .A(
        n15917), .ZN(n15919) );
  NOR2_X1 U18680 ( .A1(n15575), .A2(n15920), .ZN(n20661) );
  AOI21_X1 U18681 ( .B1(n15577), .B2(n15576), .A(n20661), .ZN(n15578) );
  OAI211_X1 U18682 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20677), .A(n15578), 
        .B(n15914), .ZN(n15579) );
  NOR2_X1 U18683 ( .A1(n15919), .A2(n15579), .ZN(n15583) );
  OR2_X1 U18684 ( .A1(n15914), .A2(n15580), .ZN(n15581) );
  NAND2_X1 U18685 ( .A1(n20578), .A2(n15581), .ZN(n15582) );
  OAI22_X1 U18686 ( .A1(n15583), .A2(n20578), .B1(n15919), .B2(n15582), .ZN(
        P1_U3161) );
  INV_X1 U18687 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n15586) );
  INV_X1 U18688 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20584) );
  INV_X1 U18689 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20685) );
  NOR2_X1 U18690 ( .A1(n20584), .A2(n20685), .ZN(n20591) );
  INV_X1 U18691 ( .A(HOLD), .ZN(n20595) );
  NOR2_X1 U18692 ( .A1(n15586), .A2(n20595), .ZN(n20587) );
  INV_X1 U18693 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20599) );
  OAI22_X1 U18694 ( .A1(n20591), .A2(n20587), .B1(n20599), .B2(n20595), .ZN(
        n15584) );
  OAI211_X1 U18695 ( .C1(n20677), .C2(n15586), .A(n15585), .B(n15584), .ZN(
        P1_U3195) );
  AND2_X1 U18696 ( .A1(n19871), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U18697 ( .A(n19740), .ZN(n19738) );
  NOR2_X1 U18698 ( .A1(n19738), .A2(n19741), .ZN(n19599) );
  NAND2_X1 U18699 ( .A1(n19599), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15588) );
  AOI21_X1 U18700 ( .B1(n19702), .B2(n19741), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15587) );
  AOI21_X1 U18701 ( .B1(n15588), .B2(n15587), .A(n16182), .ZN(P2_U3178) );
  AOI221_X1 U18702 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16182), .C1(n15589), .C2(
        n16182), .A(n19544), .ZN(n19711) );
  INV_X1 U18703 ( .A(n19711), .ZN(n19721) );
  NOR2_X1 U18704 ( .A1(n16155), .A2(n19721), .ZN(P2_U3047) );
  NOR2_X1 U18705 ( .A1(n15591), .A2(n15590), .ZN(n15592) );
  NOR2_X1 U18706 ( .A1(n18452), .A2(n17158), .ZN(n17155) );
  NAND2_X1 U18707 ( .A1(n18452), .A2(n17149), .ZN(n17147) );
  AOI22_X1 U18708 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17156), .B1(
        P3_EAX_REG_0__SCAN_IN), .B2(n17158), .ZN(n15594) );
  INV_X1 U18709 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17222) );
  NOR2_X1 U18710 ( .A1(n17092), .A2(n17158), .ZN(n17154) );
  NAND2_X1 U18711 ( .A1(n17222), .A2(n17154), .ZN(n17157) );
  OAI211_X1 U18712 ( .C1(n15595), .C2(n17144), .A(n15594), .B(n17157), .ZN(
        P3_U2735) );
  NOR3_X1 U18713 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n19820), .A3(n15596), 
        .ZN(n15600) );
  OAI22_X1 U18714 ( .A1(n19791), .A2(n15598), .B1(n15597), .B2(n19833), .ZN(
        n15599) );
  AOI211_X1 U18715 ( .C1(n19816), .C2(n15601), .A(n15600), .B(n15599), .ZN(
        n15605) );
  NOR2_X1 U18716 ( .A1(n15602), .A2(n15659), .ZN(n15608) );
  AOI22_X1 U18717 ( .A1(n15603), .A2(n19811), .B1(P1_REIP_REG_24__SCAN_IN), 
        .B2(n15608), .ZN(n15604) );
  OAI211_X1 U18718 ( .C1(n15606), .C2(n19835), .A(n15605), .B(n15604), .ZN(
        P1_U2816) );
  AOI222_X1 U18719 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19832), .B1(
        n19816), .B2(n15607), .C1(n19818), .C2(P1_EBX_REG_23__SCAN_IN), .ZN(
        n15612) );
  AOI22_X1 U18720 ( .A1(n15737), .A2(n19811), .B1(n15734), .B2(n19815), .ZN(
        n15611) );
  NAND2_X1 U18721 ( .A1(n15658), .A2(n15730), .ZN(n15665) );
  NOR2_X1 U18722 ( .A1(n15650), .A2(n15665), .ZN(n15642) );
  OAI221_X1 U18723 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(n15609), .C1(
        P1_REIP_REG_23__SCAN_IN), .C2(n15642), .A(n15608), .ZN(n15610) );
  NAND3_X1 U18724 ( .A1(n15612), .A2(n15611), .A3(n15610), .ZN(P1_U2817) );
  NAND2_X1 U18725 ( .A1(n15613), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15630) );
  AOI21_X1 U18726 ( .B1(n15615), .B2(n15630), .A(n19792), .ZN(n15643) );
  INV_X1 U18727 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15614) );
  NAND2_X1 U18728 ( .A1(n15615), .A2(n15614), .ZN(n15631) );
  AOI21_X1 U18729 ( .B1(n15643), .B2(n15631), .A(n20628), .ZN(n15619) );
  OAI22_X1 U18730 ( .A1(n19791), .A2(n15617), .B1(n15616), .B2(n19833), .ZN(
        n15618) );
  AOI211_X1 U18731 ( .C1(n19816), .C2(n15620), .A(n15619), .B(n15618), .ZN(
        n15625) );
  NOR2_X1 U18732 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n15621), .ZN(n15622) );
  AOI22_X1 U18733 ( .A1(n15623), .A2(n19811), .B1(n15622), .B2(n15642), .ZN(
        n15624) );
  OAI211_X1 U18734 ( .C1(n19835), .C2(n15626), .A(n15625), .B(n15624), .ZN(
        P1_U2818) );
  INV_X1 U18735 ( .A(n15627), .ZN(n15635) );
  INV_X1 U18736 ( .A(n15643), .ZN(n15628) );
  AOI22_X1 U18737 ( .A1(n19818), .A2(P1_EBX_REG_21__SCAN_IN), .B1(n15628), 
        .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15629) );
  OAI21_X1 U18738 ( .B1(n15631), .B2(n15630), .A(n15629), .ZN(n15634) );
  INV_X1 U18739 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15632) );
  NOR2_X1 U18740 ( .A1(n19791), .A2(n15632), .ZN(n15633) );
  AOI211_X1 U18741 ( .C1(n19816), .C2(n15635), .A(n15634), .B(n15633), .ZN(
        n15639) );
  AOI22_X1 U18742 ( .A1(n15637), .A2(n19811), .B1(n15636), .B2(n19815), .ZN(
        n15638) );
  NAND2_X1 U18743 ( .A1(n15639), .A2(n15638), .ZN(P1_U2819) );
  AOI22_X1 U18744 ( .A1(n19816), .A2(n15640), .B1(P1_EBX_REG_20__SCAN_IN), 
        .B2(n19818), .ZN(n15648) );
  INV_X1 U18745 ( .A(n15641), .ZN(n15741) );
  NOR2_X1 U18746 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n15642), .ZN(n15644) );
  OAI22_X1 U18747 ( .A1(n15645), .A2(n19835), .B1(n15644), .B2(n15643), .ZN(
        n15646) );
  AOI21_X1 U18748 ( .B1(n15741), .B2(n19811), .A(n15646), .ZN(n15647) );
  OAI211_X1 U18749 ( .C1(n15649), .C2(n19791), .A(n15648), .B(n15647), .ZN(
        P1_U2820) );
  OAI21_X1 U18750 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(P1_REIP_REG_18__SCAN_IN), 
        .A(n15650), .ZN(n15656) );
  INV_X1 U18751 ( .A(n15756), .ZN(n15653) );
  OAI21_X1 U18752 ( .B1(n19833), .B2(n15651), .A(n19823), .ZN(n15652) );
  AOI21_X1 U18753 ( .B1(n19816), .B2(n15653), .A(n15652), .ZN(n15655) );
  NAND2_X1 U18754 ( .A1(n19832), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15654) );
  OAI211_X1 U18755 ( .C1(n15665), .C2(n15656), .A(n15655), .B(n15654), .ZN(
        n15657) );
  INV_X1 U18756 ( .A(n15657), .ZN(n15661) );
  OAI21_X1 U18757 ( .B1(n15659), .B2(n15658), .A(n19783), .ZN(n15672) );
  AOI22_X1 U18758 ( .A1(n15752), .A2(n19811), .B1(P1_REIP_REG_19__SCAN_IN), 
        .B2(n15672), .ZN(n15660) );
  OAI211_X1 U18759 ( .C1(n19835), .C2(n15662), .A(n15661), .B(n15660), .ZN(
        P1_U2821) );
  AOI22_X1 U18760 ( .A1(n15663), .A2(n19816), .B1(P1_EBX_REG_18__SCAN_IN), 
        .B2(n19818), .ZN(n15664) );
  OAI21_X1 U18761 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n15665), .A(n15664), 
        .ZN(n15666) );
  AOI211_X1 U18762 ( .C1(n19832), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n19950), .B(n15666), .ZN(n15669) );
  AOI22_X1 U18763 ( .A1(n15667), .A2(n19811), .B1(P1_REIP_REG_18__SCAN_IN), 
        .B2(n15672), .ZN(n15668) );
  OAI211_X1 U18764 ( .C1(n19835), .C2(n15813), .A(n15669), .B(n15668), .ZN(
        P1_U2822) );
  AOI22_X1 U18765 ( .A1(n19832), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n19818), .B2(P1_EBX_REG_17__SCAN_IN), .ZN(n15677) );
  AOI21_X1 U18766 ( .B1(n19816), .B2(n15762), .A(n19950), .ZN(n15676) );
  OAI22_X1 U18767 ( .A1(n15764), .A2(n19795), .B1(n19835), .B2(n15824), .ZN(
        n15670) );
  INV_X1 U18768 ( .A(n15670), .ZN(n15675) );
  NOR2_X1 U18769 ( .A1(n20620), .A2(n15831), .ZN(n15673) );
  NOR2_X1 U18770 ( .A1(n15671), .A2(n19781), .ZN(n15685) );
  OAI221_X1 U18771 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n15673), .C1(
        P1_REIP_REG_17__SCAN_IN), .C2(n15685), .A(n15672), .ZN(n15674) );
  NAND4_X1 U18772 ( .A1(n15677), .A2(n15676), .A3(n15675), .A4(n15674), .ZN(
        P1_U2823) );
  NAND2_X1 U18773 ( .A1(n15685), .A2(n15831), .ZN(n15692) );
  AOI21_X1 U18774 ( .B1(n15696), .B2(n15692), .A(n20620), .ZN(n15683) );
  AOI21_X1 U18775 ( .B1(n19818), .B2(P1_EBX_REG_16__SCAN_IN), .A(n19950), .ZN(
        n15680) );
  NAND2_X1 U18776 ( .A1(n19816), .A2(n15678), .ZN(n15679) );
  OAI211_X1 U18777 ( .C1(n19791), .C2(n15681), .A(n15680), .B(n15679), .ZN(
        n15682) );
  AOI211_X1 U18778 ( .C1(n15684), .C2(n19811), .A(n15683), .B(n15682), .ZN(
        n15687) );
  NAND3_X1 U18779 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n15685), .A3(n20620), 
        .ZN(n15686) );
  OAI211_X1 U18780 ( .C1(n15688), .C2(n19835), .A(n15687), .B(n15686), .ZN(
        P1_U2824) );
  INV_X1 U18781 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15693) );
  AOI22_X1 U18782 ( .A1(n15775), .A2(n19816), .B1(n19815), .B2(n15835), .ZN(
        n15689) );
  INV_X1 U18783 ( .A(n15689), .ZN(n15690) );
  AOI211_X1 U18784 ( .C1(n19818), .C2(P1_EBX_REG_15__SCAN_IN), .A(n19950), .B(
        n15690), .ZN(n15691) );
  OAI211_X1 U18785 ( .C1(n15693), .C2(n19791), .A(n15692), .B(n15691), .ZN(
        n15694) );
  AOI21_X1 U18786 ( .B1(n15776), .B2(n19811), .A(n15694), .ZN(n15695) );
  OAI21_X1 U18787 ( .B1(n15831), .B2(n15696), .A(n15695), .ZN(P1_U2825) );
  OAI21_X1 U18788 ( .B1(n15697), .B2(n15715), .A(n19806), .ZN(n15713) );
  NAND2_X1 U18789 ( .A1(n19816), .A2(n15698), .ZN(n15700) );
  AOI21_X1 U18790 ( .B1(n19832), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n19950), .ZN(n15699) );
  OAI211_X1 U18791 ( .C1(n19833), .C2(n15701), .A(n15700), .B(n15699), .ZN(
        n15704) );
  NOR2_X1 U18792 ( .A1(n15702), .A2(n19795), .ZN(n15703) );
  AOI211_X1 U18793 ( .C1(n15705), .C2(n19815), .A(n15704), .B(n15703), .ZN(
        n15706) );
  OAI221_X1 U18794 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15707), .C1(n20615), 
        .C2(n15713), .A(n15706), .ZN(P1_U2827) );
  AOI21_X1 U18795 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15721), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15714) );
  AOI22_X1 U18796 ( .A1(n15780), .A2(n19816), .B1(n19815), .B2(n15708), .ZN(
        n15712) );
  OAI22_X1 U18797 ( .A1(n19791), .A2(n15709), .B1(n20835), .B2(n19833), .ZN(
        n15710) );
  AOI211_X1 U18798 ( .C1(n15779), .C2(n19811), .A(n19950), .B(n15710), .ZN(
        n15711) );
  OAI211_X1 U18799 ( .C1(n15714), .C2(n15713), .A(n15712), .B(n15711), .ZN(
        P1_U2828) );
  INV_X1 U18800 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20613) );
  OAI21_X1 U18801 ( .B1(n15716), .B2(n15715), .A(n19806), .ZN(n15725) );
  OAI22_X1 U18802 ( .A1(n15840), .A2(n19835), .B1(n19833), .B2(n15717), .ZN(
        n15718) );
  INV_X1 U18803 ( .A(n15718), .ZN(n15719) );
  OAI21_X1 U18804 ( .B1(n15792), .B2(n19828), .A(n15719), .ZN(n15720) );
  AOI211_X1 U18805 ( .C1(n19832), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n19950), .B(n15720), .ZN(n15723) );
  AOI22_X1 U18806 ( .A1(n15789), .A2(n19811), .B1(n15721), .B2(n20613), .ZN(
        n15722) );
  OAI211_X1 U18807 ( .C1(n20613), .C2(n15725), .A(n15723), .B(n15722), .ZN(
        P1_U2829) );
  AOI22_X1 U18808 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19832), .B1(
        n19815), .B2(n15849), .ZN(n15733) );
  NOR2_X1 U18809 ( .A1(n19833), .A2(n15724), .ZN(n15728) );
  OAI22_X1 U18810 ( .A1(n15726), .A2(n19795), .B1(n14529), .B2(n15725), .ZN(
        n15727) );
  AOI211_X1 U18811 ( .C1(n19816), .C2(n15729), .A(n15728), .B(n15727), .ZN(
        n15732) );
  NAND3_X1 U18812 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n15730), .A3(n14529), 
        .ZN(n15731) );
  NAND4_X1 U18813 ( .A1(n15733), .A2(n15732), .A3(n19823), .A4(n15731), .ZN(
        P1_U2830) );
  AOI22_X1 U18814 ( .A1(n15737), .A2(n19854), .B1(n15734), .B2(n19853), .ZN(
        n15735) );
  OAI21_X1 U18815 ( .B1(n19858), .B2(n20738), .A(n15735), .ZN(P1_U2849) );
  INV_X1 U18816 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16236) );
  AOI22_X1 U18817 ( .A1(n15746), .A2(n15736), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n15744), .ZN(n15739) );
  AOI22_X1 U18818 ( .A1(n15737), .A2(n15748), .B1(n15747), .B2(DATAI_23_), 
        .ZN(n15738) );
  OAI211_X1 U18819 ( .C1(n15751), .C2(n16236), .A(n15739), .B(n15738), .ZN(
        P1_U2881) );
  INV_X1 U18820 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16241) );
  AOI22_X1 U18821 ( .A1(n15746), .A2(n15740), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n15744), .ZN(n15743) );
  AOI22_X1 U18822 ( .A1(n15741), .A2(n15748), .B1(n15747), .B2(DATAI_20_), 
        .ZN(n15742) );
  OAI211_X1 U18823 ( .C1(n15751), .C2(n16241), .A(n15743), .B(n15742), .ZN(
        P1_U2884) );
  INV_X1 U18824 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16243) );
  AOI22_X1 U18825 ( .A1(n15746), .A2(n15745), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n15744), .ZN(n15750) );
  AOI22_X1 U18826 ( .A1(n15752), .A2(n15748), .B1(n15747), .B2(DATAI_19_), 
        .ZN(n15749) );
  OAI211_X1 U18827 ( .C1(n15751), .C2(n16243), .A(n15750), .B(n15749), .ZN(
        P1_U2885) );
  AOI22_X1 U18828 ( .A1(n19925), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n19950), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15755) );
  AOI22_X1 U18829 ( .A1(n15753), .A2(n19930), .B1(n19942), .B2(n15752), .ZN(
        n15754) );
  OAI211_X1 U18830 ( .C1(n19934), .C2(n15756), .A(n15755), .B(n15754), .ZN(
        P1_U2980) );
  AOI21_X1 U18831 ( .B1(n14495), .B2(n15758), .A(n15757), .ZN(n15760) );
  NOR2_X1 U18832 ( .A1(n15760), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15759) );
  MUX2_X1 U18833 ( .A(n15760), .B(n15759), .S(n9590), .Z(n15761) );
  XNOR2_X1 U18834 ( .A(n15761), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15829) );
  AOI22_X1 U18835 ( .A1(n19925), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n19950), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15767) );
  INV_X1 U18836 ( .A(n15762), .ZN(n15763) );
  OAI22_X1 U18837 ( .A1(n15764), .A2(n20003), .B1(n15763), .B2(n19934), .ZN(
        n15765) );
  INV_X1 U18838 ( .A(n15765), .ZN(n15766) );
  OAI211_X1 U18839 ( .C1(n19944), .C2(n15829), .A(n15767), .B(n15766), .ZN(
        P1_U2982) );
  INV_X1 U18840 ( .A(n15768), .ZN(n15769) );
  NOR2_X1 U18841 ( .A1(n15770), .A2(n15769), .ZN(n15774) );
  NAND2_X1 U18842 ( .A1(n15772), .A2(n15771), .ZN(n15773) );
  XNOR2_X1 U18843 ( .A(n15774), .B(n15773), .ZN(n15832) );
  AOI22_X1 U18844 ( .A1(n19925), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n19950), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15778) );
  AOI22_X1 U18845 ( .A1(n15776), .A2(n19942), .B1(n15775), .B2(n15781), .ZN(
        n15777) );
  OAI211_X1 U18846 ( .C1(n15832), .C2(n19944), .A(n15778), .B(n15777), .ZN(
        P1_U2984) );
  AOI22_X1 U18847 ( .A1(n19925), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n19950), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15783) );
  AOI22_X1 U18848 ( .A1(n15781), .A2(n15780), .B1(n19942), .B2(n15779), .ZN(
        n15782) );
  OAI211_X1 U18849 ( .C1(n15784), .C2(n19944), .A(n15783), .B(n15782), .ZN(
        P1_U2987) );
  AOI22_X1 U18850 ( .A1(n19925), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n19950), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15791) );
  NOR2_X1 U18851 ( .A1(n14527), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15787) );
  NOR2_X1 U18852 ( .A1(n14495), .A2(n13898), .ZN(n15786) );
  MUX2_X1 U18853 ( .A(n15787), .B(n15786), .S(n15785), .Z(n15788) );
  XOR2_X1 U18854 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n15788), .Z(
        n15842) );
  AOI22_X1 U18855 ( .A1(n19930), .A2(n15842), .B1(n19942), .B2(n15789), .ZN(
        n15790) );
  OAI211_X1 U18856 ( .C1(n19934), .C2(n15792), .A(n15791), .B(n15790), .ZN(
        P1_U2988) );
  AOI22_X1 U18857 ( .A1(n19925), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n19950), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15799) );
  NAND2_X1 U18858 ( .A1(n15794), .A2(n15793), .ZN(n15795) );
  XNOR2_X1 U18859 ( .A(n9648), .B(n15795), .ZN(n15884) );
  AOI22_X1 U18860 ( .A1(n15884), .A2(n19930), .B1(n19942), .B2(n15797), .ZN(
        n15798) );
  OAI211_X1 U18861 ( .C1(n19934), .C2(n19803), .A(n15799), .B(n15798), .ZN(
        P1_U2992) );
  AOI22_X1 U18862 ( .A1(n19925), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n19950), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15804) );
  XNOR2_X1 U18863 ( .A(n15800), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15801) );
  XNOR2_X1 U18864 ( .A(n15802), .B(n15801), .ZN(n15891) );
  AOI22_X1 U18865 ( .A1(n15891), .A2(n19930), .B1(n19942), .B2(n19849), .ZN(
        n15803) );
  OAI211_X1 U18866 ( .C1(n19934), .C2(n19804), .A(n15804), .B(n15803), .ZN(
        P1_U2993) );
  AOI22_X1 U18867 ( .A1(n19925), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n19950), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15810) );
  OAI21_X1 U18868 ( .B1(n15807), .B2(n15806), .A(n9655), .ZN(n15808) );
  INV_X1 U18869 ( .A(n15808), .ZN(n15901) );
  AOI22_X1 U18870 ( .A1(n15901), .A2(n19930), .B1(n19942), .B2(n19855), .ZN(
        n15809) );
  OAI211_X1 U18871 ( .C1(n19934), .C2(n19814), .A(n15810), .B(n15809), .ZN(
        P1_U2994) );
  AOI21_X1 U18872 ( .B1(n15874), .B2(n15812), .A(n15811), .ZN(n15821) );
  NOR2_X1 U18873 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15812), .ZN(
        n15818) );
  AND2_X1 U18874 ( .A1(n19950), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15816) );
  OAI22_X1 U18875 ( .A1(n15814), .A2(n19998), .B1(n19953), .B2(n15813), .ZN(
        n15815) );
  AOI211_X1 U18876 ( .C1(n15818), .C2(n15817), .A(n15816), .B(n15815), .ZN(
        n15819) );
  OAI21_X1 U18877 ( .B1(n15821), .B2(n15820), .A(n15819), .ZN(P1_U3013) );
  AOI221_X1 U18878 ( .B1(n15823), .B2(n15822), .C1(n15830), .C2(n15822), .A(
        n15821), .ZN(n15826) );
  NOR2_X1 U18879 ( .A1(n15824), .A2(n19953), .ZN(n15825) );
  NOR2_X1 U18880 ( .A1(n15826), .A2(n15825), .ZN(n15828) );
  NAND2_X1 U18881 ( .A1(n19950), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15827) );
  OAI211_X1 U18882 ( .C1(n15829), .C2(n19998), .A(n15828), .B(n15827), .ZN(
        P1_U3014) );
  INV_X1 U18883 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15837) );
  OAI22_X1 U18884 ( .A1(n19823), .A2(n15831), .B1(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15830), .ZN(n15834) );
  NOR2_X1 U18885 ( .A1(n15832), .A2(n19998), .ZN(n15833) );
  AOI211_X1 U18886 ( .C1(n19993), .C2(n15835), .A(n15834), .B(n15833), .ZN(
        n15836) );
  OAI21_X1 U18887 ( .B1(n15838), .B2(n15837), .A(n15836), .ZN(P1_U3016) );
  INV_X1 U18888 ( .A(n15839), .ZN(n15846) );
  OAI22_X1 U18889 ( .A1(n15840), .A2(n19953), .B1(n19823), .B2(n20613), .ZN(
        n15841) );
  INV_X1 U18890 ( .A(n15841), .ZN(n15845) );
  AOI22_X1 U18891 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15843), .B1(
        n19973), .B2(n15842), .ZN(n15844) );
  OAI211_X1 U18892 ( .C1(n15894), .C2(n15846), .A(n15845), .B(n15844), .ZN(
        P1_U3020) );
  INV_X1 U18893 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15875) );
  NOR2_X1 U18894 ( .A1(n15875), .A2(n15894), .ZN(n15883) );
  NAND2_X1 U18895 ( .A1(n15847), .A2(n15883), .ZN(n15867) );
  AOI22_X1 U18896 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n11999), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n13898), .ZN(n15856) );
  AOI21_X1 U18897 ( .B1(n15849), .B2(n19993), .A(n15848), .ZN(n15855) );
  AOI211_X1 U18898 ( .C1(n19971), .C2(n15850), .A(n15875), .B(n15879), .ZN(
        n15852) );
  AOI21_X1 U18899 ( .B1(n15870), .B2(n15852), .A(n15851), .ZN(n15863) );
  AOI22_X1 U18900 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15863), .B1(
        n19973), .B2(n15853), .ZN(n15854) );
  OAI211_X1 U18901 ( .C1(n15867), .C2(n15856), .A(n15855), .B(n15854), .ZN(
        P1_U3021) );
  NAND2_X1 U18902 ( .A1(n15858), .A2(n15857), .ZN(n15859) );
  AND2_X1 U18903 ( .A1(n15860), .A2(n15859), .ZN(n19842) );
  INV_X1 U18904 ( .A(n15861), .ZN(n15862) );
  AOI21_X1 U18905 ( .B1(n19842), .B2(n19993), .A(n15862), .ZN(n15866) );
  AOI22_X1 U18906 ( .A1(n15864), .A2(n19973), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15863), .ZN(n15865) );
  OAI211_X1 U18907 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n15867), .A(
        n15866), .B(n15865), .ZN(P1_U3022) );
  NAND2_X1 U18908 ( .A1(n19948), .A2(n15868), .ZN(n15905) );
  INV_X1 U18909 ( .A(n19948), .ZN(n15872) );
  AOI21_X1 U18910 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n15869), .ZN(n19947) );
  INV_X1 U18911 ( .A(n15870), .ZN(n15871) );
  AOI211_X1 U18912 ( .C1(n19971), .C2(n15872), .A(n19947), .B(n15871), .ZN(
        n15900) );
  OAI21_X1 U18913 ( .B1(n15873), .B2(n15905), .A(n15900), .ZN(n15890) );
  AOI21_X1 U18914 ( .B1(n15875), .B2(n15874), .A(n15890), .ZN(n15888) );
  INV_X1 U18915 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15882) );
  OAI222_X1 U18916 ( .A1(n15877), .A2(n19953), .B1(n19823), .B2(n13859), .C1(
        n19998), .C2(n15876), .ZN(n15878) );
  INV_X1 U18917 ( .A(n15878), .ZN(n15881) );
  OAI211_X1 U18918 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n15883), .B(n15879), .ZN(n15880) );
  OAI211_X1 U18919 ( .C1(n15888), .C2(n15882), .A(n15881), .B(n15880), .ZN(
        P1_U3023) );
  INV_X1 U18920 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15887) );
  AOI22_X1 U18921 ( .A1(n19800), .A2(n19993), .B1(n19950), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n15886) );
  AOI22_X1 U18922 ( .A1(n15884), .A2(n19973), .B1(n15883), .B2(n15887), .ZN(
        n15885) );
  OAI211_X1 U18923 ( .C1(n15888), .C2(n15887), .A(n15886), .B(n15885), .ZN(
        P1_U3024) );
  XNOR2_X1 U18924 ( .A(n15896), .B(n15889), .ZN(n19848) );
  AOI22_X1 U18925 ( .A1(n19993), .A2(n19848), .B1(n19950), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n15893) );
  AOI22_X1 U18926 ( .A1(n15891), .A2(n19973), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15890), .ZN(n15892) );
  OAI211_X1 U18927 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n15894), .A(
        n15893), .B(n15892), .ZN(P1_U3025) );
  NAND2_X1 U18928 ( .A1(n19945), .A2(n15895), .ZN(n19963) );
  INV_X1 U18929 ( .A(n15896), .ZN(n15897) );
  AOI21_X1 U18930 ( .B1(n15899), .B2(n15898), .A(n15897), .ZN(n19852) );
  AOI22_X1 U18931 ( .A1(n19993), .A2(n19852), .B1(n19950), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n15904) );
  INV_X1 U18932 ( .A(n15900), .ZN(n15902) );
  AOI22_X1 U18933 ( .A1(n15902), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n19973), .B2(n15901), .ZN(n15903) );
  OAI211_X1 U18934 ( .C1(n15905), .C2(n19963), .A(n15904), .B(n15903), .ZN(
        P1_U3026) );
  INV_X1 U18935 ( .A(n15906), .ZN(n20655) );
  NAND3_X1 U18936 ( .A1(n15909), .A2(n15908), .A3(n15907), .ZN(n15910) );
  OAI21_X1 U18937 ( .B1(n20655), .B2(n11469), .A(n15910), .ZN(P1_U3468) );
  NAND4_X1 U18938 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20581), .A4(n20677), .ZN(n15911) );
  NAND2_X1 U18939 ( .A1(n15912), .A2(n15911), .ZN(n20579) );
  OAI21_X1 U18940 ( .B1(n15919), .B2(n20578), .A(n20577), .ZN(n15913) );
  OAI211_X1 U18941 ( .C1(n15915), .C2(n20677), .A(n15914), .B(n15913), .ZN(
        n15916) );
  AOI221_X1 U18942 ( .B1(n15918), .B2(n15917), .C1(n20579), .C2(n15917), .A(
        n15916), .ZN(P1_U3162) );
  NOR2_X1 U18943 ( .A1(n15919), .A2(n20578), .ZN(n15921) );
  OAI22_X1 U18944 ( .A1(n20412), .A2(n15921), .B1(n15920), .B2(n20578), .ZN(
        P1_U3466) );
  AOI22_X1 U18945 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18901), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n18890), .ZN(n15924) );
  AOI22_X1 U18946 ( .A1(n15922), .A2(n18876), .B1(P2_EBX_REG_29__SCAN_IN), 
        .B2(n18889), .ZN(n15923) );
  OAI211_X1 U18947 ( .C1(n15092), .C2(n18893), .A(n15924), .B(n15923), .ZN(
        n15928) );
  NOR2_X1 U18948 ( .A1(n15928), .A2(n15927), .ZN(n15929) );
  OAI21_X1 U18949 ( .B1(n15930), .B2(n18871), .A(n15929), .ZN(P2_U2826) );
  AOI211_X1 U18950 ( .C1(n15933), .C2(n15932), .A(n15931), .B(n19606), .ZN(
        n15938) );
  NAND2_X1 U18951 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n18889), .ZN(n15935) );
  AOI22_X1 U18952 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18901), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n18890), .ZN(n15934) );
  OAI211_X1 U18953 ( .C1(n15936), .C2(n18888), .A(n15935), .B(n15934), .ZN(
        n15937) );
  AOI211_X1 U18954 ( .C1(n18877), .C2(n15939), .A(n15938), .B(n15937), .ZN(
        n15940) );
  OAI21_X1 U18955 ( .B1(n15941), .B2(n18871), .A(n15940), .ZN(P2_U2827) );
  AOI211_X1 U18956 ( .C1(n15944), .C2(n15943), .A(n15942), .B(n19606), .ZN(
        n15950) );
  AOI22_X1 U18957 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18901), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n18890), .ZN(n15947) );
  AOI22_X1 U18958 ( .A1(n15945), .A2(n18876), .B1(P2_EBX_REG_26__SCAN_IN), 
        .B2(n18889), .ZN(n15946) );
  OAI211_X1 U18959 ( .C1(n15948), .C2(n18871), .A(n15947), .B(n15946), .ZN(
        n15949) );
  AOI211_X1 U18960 ( .C1(n18877), .C2(n15951), .A(n15950), .B(n15949), .ZN(
        n15952) );
  INV_X1 U18961 ( .A(n15952), .ZN(P2_U2829) );
  AOI211_X1 U18962 ( .C1(P2_EBX_REG_25__SCAN_IN), .C2(n15968), .A(n18888), .B(
        n15953), .ZN(n15956) );
  INV_X1 U18963 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15954) );
  OAI22_X1 U18964 ( .A1(n18857), .A2(n15954), .B1(n19654), .B2(n18849), .ZN(
        n15955) );
  AOI211_X1 U18965 ( .C1(n18901), .C2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15956), .B(n15955), .ZN(n15963) );
  AOI211_X1 U18966 ( .C1(n15959), .C2(n15958), .A(n15957), .B(n19606), .ZN(
        n15960) );
  AOI21_X1 U18967 ( .B1(n18896), .B2(n15961), .A(n15960), .ZN(n15962) );
  OAI211_X1 U18968 ( .C1(n15964), .C2(n18893), .A(n15963), .B(n15962), .ZN(
        P2_U2830) );
  AOI211_X1 U18969 ( .C1(n15967), .C2(n15966), .A(n15965), .B(n19606), .ZN(
        n15972) );
  AOI22_X1 U18970 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18901), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18890), .ZN(n15970) );
  OAI211_X1 U18971 ( .C1(n9700), .C2(n14834), .A(n18876), .B(n15968), .ZN(
        n15969) );
  OAI211_X1 U18972 ( .C1(n18857), .C2(n14834), .A(n15970), .B(n15969), .ZN(
        n15971) );
  AOI211_X1 U18973 ( .C1(n18877), .C2(n15973), .A(n15972), .B(n15971), .ZN(
        n15974) );
  OAI21_X1 U18974 ( .B1(n15975), .B2(n18871), .A(n15974), .ZN(P2_U2831) );
  AOI22_X1 U18975 ( .A1(n18909), .A2(n15976), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n18963), .ZN(n15981) );
  AOI22_X1 U18976 ( .A1(n18911), .A2(BUF1_REG_22__SCAN_IN), .B1(n18910), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n15980) );
  AOI22_X1 U18977 ( .A1(n15978), .A2(n18945), .B1(n18964), .B2(n15977), .ZN(
        n15979) );
  NAND3_X1 U18978 ( .A1(n15981), .A2(n15980), .A3(n15979), .ZN(P2_U2897) );
  AOI22_X1 U18979 ( .A1(n18909), .A2(n15982), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n18963), .ZN(n15989) );
  AOI22_X1 U18980 ( .A1(n18911), .A2(BUF1_REG_20__SCAN_IN), .B1(n18910), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n15988) );
  INV_X1 U18981 ( .A(n15983), .ZN(n15984) );
  OAI22_X1 U18982 ( .A1(n15985), .A2(n18968), .B1(n18954), .B2(n15984), .ZN(
        n15986) );
  INV_X1 U18983 ( .A(n15986), .ZN(n15987) );
  NAND3_X1 U18984 ( .A1(n15989), .A2(n15988), .A3(n15987), .ZN(P2_U2899) );
  AOI22_X1 U18985 ( .A1(n18909), .A2(n15990), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n18963), .ZN(n15994) );
  AOI22_X1 U18986 ( .A1(n18911), .A2(BUF1_REG_18__SCAN_IN), .B1(n18910), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n15993) );
  AOI22_X1 U18987 ( .A1(n15991), .A2(n18945), .B1(n18964), .B2(n18700), .ZN(
        n15992) );
  NAND3_X1 U18988 ( .A1(n15994), .A2(n15993), .A3(n15992), .ZN(P2_U2901) );
  AOI22_X1 U18989 ( .A1(n19012), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19011), .ZN(n16003) );
  INV_X1 U18990 ( .A(n15996), .ZN(n15998) );
  NAND2_X1 U18991 ( .A1(n15998), .A2(n15997), .ZN(n15999) );
  XNOR2_X1 U18992 ( .A(n15995), .B(n15999), .ZN(n16085) );
  AOI21_X1 U18993 ( .B1(n16001), .B2(n16000), .A(n14987), .ZN(n16083) );
  AOI222_X1 U18994 ( .A1(n16085), .A2(n19013), .B1(n16067), .B2(n16084), .C1(
        n19015), .C2(n16083), .ZN(n16002) );
  OAI211_X1 U18995 ( .C1(n19025), .C2(n16004), .A(n16003), .B(n16002), .ZN(
        P2_U2992) );
  AOI22_X1 U18996 ( .A1(n19012), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n19011), .ZN(n16012) );
  AOI21_X1 U18997 ( .B1(n16005), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16007) );
  NOR3_X1 U18998 ( .A1(n16007), .A2(n16006), .A3(n16073), .ZN(n16009) );
  NOR2_X1 U18999 ( .A1(n19020), .A2(n18727), .ZN(n16008) );
  AOI211_X1 U19000 ( .C1(n16010), .C2(n19013), .A(n16009), .B(n16008), .ZN(
        n16011) );
  OAI211_X1 U19001 ( .C1(n19025), .C2(n18722), .A(n16012), .B(n16011), .ZN(
        P2_U2998) );
  AOI22_X1 U19002 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19011), .B1(n16052), 
        .B2(n18729), .ZN(n16017) );
  OAI22_X1 U19003 ( .A1(n16014), .A2(n16072), .B1(n16073), .B2(n16013), .ZN(
        n16015) );
  AOI21_X1 U19004 ( .B1(n16067), .B2(n18733), .A(n16015), .ZN(n16016) );
  OAI211_X1 U19005 ( .C1(n16059), .C2(n16018), .A(n16017), .B(n16016), .ZN(
        P2_U2999) );
  AOI22_X1 U19006 ( .A1(n19012), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19011), .ZN(n16025) );
  NAND2_X1 U19007 ( .A1(n16019), .A2(n19013), .ZN(n16022) );
  NAND2_X1 U19008 ( .A1(n16020), .A2(n19015), .ZN(n16021) );
  OAI211_X1 U19009 ( .C1(n19020), .C2(n18751), .A(n16022), .B(n16021), .ZN(
        n16023) );
  INV_X1 U19010 ( .A(n16023), .ZN(n16024) );
  OAI211_X1 U19011 ( .C1(n19025), .C2(n18747), .A(n16025), .B(n16024), .ZN(
        P2_U3000) );
  AOI22_X1 U19012 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19011), .B1(n16052), 
        .B2(n18756), .ZN(n16031) );
  OAI22_X1 U19013 ( .A1(n16027), .A2(n16072), .B1(n16026), .B2(n16073), .ZN(
        n16028) );
  AOI21_X1 U19014 ( .B1(n16067), .B2(n16029), .A(n16028), .ZN(n16030) );
  OAI211_X1 U19015 ( .C1(n16059), .C2(n16032), .A(n16031), .B(n16030), .ZN(
        P2_U3001) );
  AOI22_X1 U19016 ( .A1(n19012), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19011), .ZN(n16040) );
  NAND2_X1 U19017 ( .A1(n16033), .A2(n19013), .ZN(n16037) );
  NAND3_X1 U19018 ( .A1(n16035), .A2(n19015), .A3(n16034), .ZN(n16036) );
  OAI211_X1 U19019 ( .C1(n19020), .C2(n18772), .A(n16037), .B(n16036), .ZN(
        n16038) );
  INV_X1 U19020 ( .A(n16038), .ZN(n16039) );
  OAI211_X1 U19021 ( .C1(n19025), .C2(n18766), .A(n16040), .B(n16039), .ZN(
        P2_U3002) );
  AOI22_X1 U19022 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19011), .B1(n16052), 
        .B2(n18780), .ZN(n16045) );
  OAI22_X1 U19023 ( .A1(n16042), .A2(n16073), .B1(n16041), .B2(n16072), .ZN(
        n16043) );
  AOI21_X1 U19024 ( .B1(n16067), .B2(n18773), .A(n16043), .ZN(n16044) );
  OAI211_X1 U19025 ( .C1(n16059), .C2(n16046), .A(n16045), .B(n16044), .ZN(
        P2_U3003) );
  AOI22_X1 U19026 ( .A1(n19012), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19011), .ZN(n16051) );
  AOI222_X1 U19027 ( .A1(n16049), .A2(n19013), .B1(n16067), .B2(n16048), .C1(
        n19015), .C2(n16047), .ZN(n16050) );
  OAI211_X1 U19028 ( .C1(n19025), .C2(n18788), .A(n16051), .B(n16050), .ZN(
        P2_U3004) );
  AOI22_X1 U19029 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19011), .B1(n16052), 
        .B2(n18804), .ZN(n16057) );
  OAI22_X1 U19030 ( .A1(n16054), .A2(n16073), .B1(n16072), .B2(n16053), .ZN(
        n16055) );
  AOI21_X1 U19031 ( .B1(n16067), .B2(n18806), .A(n16055), .ZN(n16056) );
  OAI211_X1 U19032 ( .C1(n16059), .C2(n16058), .A(n16057), .B(n16056), .ZN(
        P2_U3005) );
  AOI22_X1 U19033 ( .A1(n19012), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19011), .ZN(n16069) );
  XOR2_X1 U19034 ( .A(n16060), .B(n16061), .Z(n16106) );
  INV_X1 U19035 ( .A(n18819), .ZN(n16103) );
  NAND2_X1 U19036 ( .A1(n16062), .A2(n16063), .ZN(n16066) );
  XOR2_X1 U19037 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n16064), .Z(
        n16065) );
  XNOR2_X1 U19038 ( .A(n16066), .B(n16065), .ZN(n16101) );
  AOI222_X1 U19039 ( .A1(n16106), .A2(n19015), .B1(n16067), .B2(n16103), .C1(
        n19013), .C2(n16101), .ZN(n16068) );
  OAI211_X1 U19040 ( .C1(n19025), .C2(n18813), .A(n16069), .B(n16068), .ZN(
        P2_U3006) );
  OAI22_X1 U19041 ( .A1(n10332), .A2(n18847), .B1(n19025), .B2(n18836), .ZN(
        n16070) );
  AOI21_X1 U19042 ( .B1(n19012), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16070), .ZN(n16077) );
  OAI22_X1 U19043 ( .A1(n16074), .A2(n16073), .B1(n16072), .B2(n16071), .ZN(
        n16075) );
  INV_X1 U19044 ( .A(n16075), .ZN(n16076) );
  OAI211_X1 U19045 ( .C1(n19020), .C2(n18841), .A(n16077), .B(n16076), .ZN(
        P2_U3008) );
  NAND2_X1 U19046 ( .A1(n16078), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16080) );
  OAI22_X1 U19047 ( .A1(n16081), .A2(n16080), .B1(n16079), .B2(n16097), .ZN(
        n16082) );
  INV_X1 U19048 ( .A(n16082), .ZN(n16090) );
  AOI222_X1 U19049 ( .A1(n16085), .A2(n16102), .B1(n16104), .B2(n16084), .C1(
        n16105), .C2(n16083), .ZN(n16089) );
  NAND2_X1 U19050 ( .A1(n16086), .A2(n16001), .ZN(n16088) );
  NAND2_X1 U19051 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19011), .ZN(n16087) );
  NAND4_X1 U19052 ( .A1(n16090), .A2(n16089), .A3(n16088), .A4(n16087), .ZN(
        P2_U3024) );
  NAND2_X1 U19053 ( .A1(n16092), .A2(n16091), .ZN(n16098) );
  INV_X1 U19054 ( .A(n15362), .ZN(n16093) );
  OR2_X1 U19055 ( .A1(n16094), .A2(n16093), .ZN(n16096) );
  INV_X1 U19056 ( .A(n15350), .ZN(n16095) );
  NAND2_X1 U19057 ( .A1(n16096), .A2(n16095), .ZN(n18940) );
  OAI22_X1 U19058 ( .A1(n16099), .A2(n16098), .B1(n16097), .B2(n18940), .ZN(
        n16100) );
  INV_X1 U19059 ( .A(n16100), .ZN(n16112) );
  AOI222_X1 U19060 ( .A1(n16106), .A2(n16105), .B1(n16104), .B2(n16103), .C1(
        n16102), .C2(n16101), .ZN(n16111) );
  NAND2_X1 U19061 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19011), .ZN(n16110) );
  OAI21_X1 U19062 ( .B1(n16108), .B2(n16107), .A(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16109) );
  NAND4_X1 U19063 ( .A1(n16112), .A2(n16111), .A3(n16110), .A4(n16109), .ZN(
        P2_U3038) );
  INV_X1 U19064 ( .A(n16129), .ZN(n16149) );
  MUX2_X1 U19065 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16113), .S(
        n16149), .Z(n16166) );
  NAND2_X1 U19066 ( .A1(n16115), .A2(n16114), .ZN(n16128) );
  INV_X1 U19067 ( .A(n16122), .ZN(n16117) );
  INV_X1 U19068 ( .A(n16116), .ZN(n16120) );
  NAND2_X1 U19069 ( .A1(n16117), .A2(n16120), .ZN(n16118) );
  NAND2_X1 U19070 ( .A1(n16119), .A2(n16118), .ZN(n16126) );
  NAND3_X1 U19071 ( .A1(n16122), .A2(n16121), .A3(n16120), .ZN(n16125) );
  INV_X1 U19072 ( .A(n16123), .ZN(n16124) );
  AOI22_X1 U19073 ( .A1(n16126), .A2(n16125), .B1(n16124), .B2(n9755), .ZN(
        n16127) );
  NAND2_X1 U19074 ( .A1(n16128), .A2(n16127), .ZN(n19674) );
  MUX2_X1 U19075 ( .A(n19681), .B(n19674), .S(n16149), .Z(n16165) );
  NAND2_X1 U19076 ( .A1(n16129), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n16163) );
  INV_X1 U19077 ( .A(n16130), .ZN(n16137) );
  INV_X1 U19078 ( .A(n16131), .ZN(n16132) );
  NAND2_X1 U19079 ( .A1(n16133), .A2(n16132), .ZN(n16136) );
  NAND2_X1 U19080 ( .A1(n16138), .A2(n16134), .ZN(n16135) );
  OAI211_X1 U19081 ( .C1(n16138), .C2(n16137), .A(n16136), .B(n16135), .ZN(
        n19729) );
  NAND2_X1 U19082 ( .A1(n16140), .A2(n16139), .ZN(n16141) );
  NOR2_X1 U19083 ( .A1(n16142), .A2(n16141), .ZN(n18658) );
  OAI21_X1 U19084 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n18658), .ZN(n16159) );
  INV_X1 U19085 ( .A(n16165), .ZN(n16143) );
  NAND2_X1 U19086 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16143), .ZN(
        n16144) );
  OAI21_X1 U19087 ( .B1(n16166), .B2(n19693), .A(n16144), .ZN(n16154) );
  INV_X1 U19088 ( .A(n16151), .ZN(n16148) );
  AOI21_X1 U19089 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n16145), .A(
        n19720), .ZN(n16146) );
  OAI211_X1 U19090 ( .C1(n16148), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16147), .B(n16146), .ZN(n16150) );
  OAI211_X1 U19091 ( .C1(n19710), .C2(n16151), .A(n16150), .B(n16149), .ZN(
        n16153) );
  AOI21_X1 U19092 ( .B1(n16165), .B2(n19700), .A(n16166), .ZN(n16152) );
  OAI22_X1 U19093 ( .A1(n16154), .A2(n16153), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16152), .ZN(n16156) );
  AOI22_X1 U19094 ( .A1(n16157), .A2(n19742), .B1(n16156), .B2(n16155), .ZN(
        n16158) );
  OAI211_X1 U19095 ( .C1(n13135), .C2(n16160), .A(n16159), .B(n16158), .ZN(
        n16161) );
  NOR2_X1 U19096 ( .A1(n19729), .A2(n16161), .ZN(n16162) );
  NAND2_X1 U19097 ( .A1(n16163), .A2(n16162), .ZN(n16164) );
  AOI21_X1 U19098 ( .B1(n16166), .B2(n16165), .A(n16164), .ZN(n16181) );
  NAND2_X1 U19099 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19733), .ZN(n19602) );
  NOR2_X1 U19100 ( .A1(n19740), .A2(n19602), .ZN(n16168) );
  AOI211_X1 U19101 ( .C1(n19725), .C2(n16182), .A(n16168), .B(n16167), .ZN(
        n16180) );
  NAND2_X1 U19102 ( .A1(n16181), .A2(n19601), .ZN(n16169) );
  NAND2_X1 U19103 ( .A1(n16169), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16176) );
  NAND2_X1 U19104 ( .A1(n10264), .A2(n16170), .ZN(n16172) );
  OAI211_X1 U19105 ( .C1(n16173), .C2(n16172), .A(P2_STATE2_REG_2__SCAN_IN), 
        .B(n16171), .ZN(n16174) );
  INV_X1 U19106 ( .A(n16174), .ZN(n16175) );
  AOI21_X1 U19107 ( .B1(n19741), .B2(n19678), .A(n19739), .ZN(n16177) );
  AOI21_X1 U19108 ( .B1(n19738), .B2(n19608), .A(n16177), .ZN(n16178) );
  AOI21_X1 U19109 ( .B1(n19608), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16178), 
        .ZN(n16179) );
  OAI211_X1 U19110 ( .C1(n16181), .C2(n18657), .A(n16180), .B(n16179), .ZN(
        P2_U3176) );
  AOI221_X1 U19111 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19741), .C1(
        P2_STATE2_REG_3__SCAN_IN), .C2(n19608), .A(n16182), .ZN(n16183) );
  INV_X1 U19112 ( .A(n16183), .ZN(P2_U3593) );
  OR2_X1 U19113 ( .A1(n17454), .A2(n16184), .ZN(n16192) );
  OAI21_X1 U19114 ( .B1(n16185), .B2(n17658), .A(n17633), .ZN(n16206) );
  XNOR2_X1 U19115 ( .A(n9885), .B(n9753), .ZN(n16360) );
  AOI22_X1 U19116 ( .A1(n17965), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n17476), 
        .B2(n16360), .ZN(n16186) );
  OAI221_X1 U19117 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16188), .C1(
        n9885), .C2(n16187), .A(n16186), .ZN(n16189) );
  NOR2_X1 U19118 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16209), .ZN(
        n16207) );
  AOI21_X1 U19119 ( .B1(n16194), .B2(n16193), .A(n16192), .ZN(n16201) );
  AOI21_X1 U19120 ( .B1(n16368), .B2(n16349), .A(n9753), .ZN(n16367) );
  OAI21_X1 U19121 ( .B1(n16195), .B2(n17476), .A(n16367), .ZN(n16196) );
  OAI211_X1 U19122 ( .C1(n16199), .C2(n16198), .A(n16197), .B(n16196), .ZN(
        n16200) );
  AOI211_X1 U19123 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16202), .A(
        n16201), .B(n16200), .ZN(n16205) );
  NAND2_X1 U19124 ( .A1(n17537), .A2(n16203), .ZN(n16204) );
  OAI211_X1 U19125 ( .C1(n16207), .C2(n16206), .A(n16205), .B(n16204), .ZN(
        P3_U2801) );
  INV_X1 U19126 ( .A(n17967), .ZN(n17949) );
  NAND3_X1 U19127 ( .A1(n17431), .A2(n17949), .A3(n20801), .ZN(n16223) );
  NOR2_X1 U19128 ( .A1(n16208), .A2(n16213), .ZN(n17827) );
  INV_X1 U19129 ( .A(n17827), .ZN(n17844) );
  OAI22_X1 U19130 ( .A1(n16210), .A2(n17844), .B1(n16209), .B2(n18426), .ZN(
        n16211) );
  AOI211_X1 U19131 ( .C1(n9768), .C2(n10936), .A(n16212), .B(n16211), .ZN(
        n16217) );
  NOR2_X1 U19132 ( .A1(n17126), .A2(n16213), .ZN(n17794) );
  AOI22_X1 U19133 ( .A1(n17431), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n20801), .B2(n17546), .ZN(n17286) );
  INV_X1 U19134 ( .A(n17290), .ZN(n16214) );
  OAI21_X1 U19135 ( .B1(n16214), .B2(n17546), .A(n17291), .ZN(n17285) );
  NAND2_X1 U19136 ( .A1(n17286), .A2(n17285), .ZN(n17284) );
  OAI211_X1 U19137 ( .C1(n17290), .C2(n16215), .A(n17794), .B(n17284), .ZN(
        n16216) );
  AOI21_X1 U19138 ( .B1(n16217), .B2(n16216), .A(n20801), .ZN(n16220) );
  OAI22_X1 U19139 ( .A1(n18426), .A2(n17788), .B1(n17712), .B2(n17844), .ZN(
        n17754) );
  NOR2_X1 U19140 ( .A1(n16218), .A2(n17754), .ZN(n17687) );
  NOR2_X1 U19141 ( .A1(n17687), .A2(n17717), .ZN(n17723) );
  NAND2_X1 U19142 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17723), .ZN(
        n17703) );
  NOR4_X1 U19143 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17952), .A3(
        n17272), .A4(n17703), .ZN(n16219) );
  AOI221_X1 U19144 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(n17965), .C1(n16220), 
        .C2(n17963), .A(n16219), .ZN(n16222) );
  OR3_X1 U19145 ( .A1(n17891), .A2(n17291), .A3(n17286), .ZN(n16221) );
  OAI211_X1 U19146 ( .C1(n16223), .C2(n17290), .A(n16222), .B(n16221), .ZN(
        P3_U2834) );
  NOR3_X1 U19147 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16225) );
  NOR4_X1 U19148 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16224) );
  NAND4_X1 U19149 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16225), .A3(n16224), .A4(
        U215), .ZN(U213) );
  INV_X1 U19150 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n18974) );
  INV_X2 U19151 ( .A(U214), .ZN(n16273) );
  NOR2_X1 U19152 ( .A1(n16273), .A2(n16226), .ZN(n16270) );
  INV_X1 U19153 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16308) );
  OAI222_X1 U19154 ( .A1(U212), .A2(n18974), .B1(n16275), .B2(n19066), .C1(
        U214), .C2(n16308), .ZN(U216) );
  INV_X1 U19155 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16228) );
  AOI22_X1 U19156 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16272), .ZN(n16227) );
  OAI21_X1 U19157 ( .B1(n16228), .B2(n16275), .A(n16227), .ZN(U217) );
  AOI222_X1 U19158 ( .A1(n16272), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(n16270), 
        .B2(BUF1_REG_29__SCAN_IN), .C1(n16273), .C2(P1_DATAO_REG_29__SCAN_IN), 
        .ZN(n16229) );
  INV_X1 U19159 ( .A(n16229), .ZN(U218) );
  AOI22_X1 U19160 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16272), .ZN(n16230) );
  OAI21_X1 U19161 ( .B1(n14349), .B2(n16275), .A(n16230), .ZN(U219) );
  AOI22_X1 U19162 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16272), .ZN(n16231) );
  OAI21_X1 U19163 ( .B1(n14356), .B2(n16275), .A(n16231), .ZN(U220) );
  AOI22_X1 U19164 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16272), .ZN(n16232) );
  OAI21_X1 U19165 ( .B1(n14359), .B2(n16275), .A(n16232), .ZN(U221) );
  AOI22_X1 U19166 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16272), .ZN(n16233) );
  OAI21_X1 U19167 ( .B1(n14366), .B2(n16275), .A(n16233), .ZN(U222) );
  AOI22_X1 U19168 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16272), .ZN(n16234) );
  OAI21_X1 U19169 ( .B1(n14371), .B2(n16275), .A(n16234), .ZN(U223) );
  AOI22_X1 U19170 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16272), .ZN(n16235) );
  OAI21_X1 U19171 ( .B1(n16236), .B2(n16275), .A(n16235), .ZN(U224) );
  AOI22_X1 U19172 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16272), .ZN(n16237) );
  OAI21_X1 U19173 ( .B1(n14375), .B2(n16275), .A(n16237), .ZN(U225) );
  INV_X1 U19174 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16239) );
  AOI22_X1 U19175 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16272), .ZN(n16238) );
  OAI21_X1 U19176 ( .B1(n16239), .B2(n16275), .A(n16238), .ZN(U226) );
  AOI22_X1 U19177 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16272), .ZN(n16240) );
  OAI21_X1 U19178 ( .B1(n16241), .B2(n16275), .A(n16240), .ZN(U227) );
  AOI22_X1 U19179 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16272), .ZN(n16242) );
  OAI21_X1 U19180 ( .B1(n16243), .B2(n16275), .A(n16242), .ZN(U228) );
  AOI222_X1 U19181 ( .A1(n16272), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n16270), 
        .B2(BUF1_REG_18__SCAN_IN), .C1(n16273), .C2(P1_DATAO_REG_18__SCAN_IN), 
        .ZN(n16244) );
  INV_X1 U19182 ( .A(n16244), .ZN(U229) );
  AOI22_X1 U19183 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n16270), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16273), .ZN(n16245) );
  OAI21_X1 U19184 ( .B1(n16246), .B2(U212), .A(n16245), .ZN(U230) );
  AOI22_X1 U19185 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16272), .ZN(n16247) );
  OAI21_X1 U19186 ( .B1(n14393), .B2(n16275), .A(n16247), .ZN(U231) );
  INV_X1 U19187 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n20706) );
  AOI22_X1 U19188 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16272), .ZN(n16248) );
  OAI21_X1 U19189 ( .B1(n20706), .B2(n16275), .A(n16248), .ZN(U232) );
  INV_X1 U19190 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16250) );
  AOI22_X1 U19191 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16270), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16273), .ZN(n16249) );
  OAI21_X1 U19192 ( .B1(n16250), .B2(U212), .A(n16249), .ZN(U233) );
  INV_X1 U19193 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16252) );
  AOI22_X1 U19194 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n16270), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16273), .ZN(n16251) );
  OAI21_X1 U19195 ( .B1(n16252), .B2(U212), .A(n16251), .ZN(U234) );
  AOI22_X1 U19196 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16272), .ZN(n16253) );
  OAI21_X1 U19197 ( .B1(n16254), .B2(n16275), .A(n16253), .ZN(U235) );
  INV_X1 U19198 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16287) );
  AOI22_X1 U19199 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16270), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16273), .ZN(n16255) );
  OAI21_X1 U19200 ( .B1(n16287), .B2(U212), .A(n16255), .ZN(U236) );
  AOI22_X1 U19201 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16272), .ZN(n16256) );
  OAI21_X1 U19202 ( .B1(n16257), .B2(n16275), .A(n16256), .ZN(U237) );
  AOI222_X1 U19203 ( .A1(n16272), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n16270), 
        .B2(BUF1_REG_9__SCAN_IN), .C1(n16273), .C2(P1_DATAO_REG_9__SCAN_IN), 
        .ZN(n16258) );
  INV_X1 U19204 ( .A(n16258), .ZN(U238) );
  AOI22_X1 U19205 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16272), .ZN(n16259) );
  OAI21_X1 U19206 ( .B1(n16260), .B2(n16275), .A(n16259), .ZN(U239) );
  INV_X1 U19207 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16284) );
  AOI22_X1 U19208 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16270), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16273), .ZN(n16261) );
  OAI21_X1 U19209 ( .B1(n16284), .B2(U212), .A(n16261), .ZN(U240) );
  INV_X1 U19210 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16263) );
  AOI22_X1 U19211 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16272), .ZN(n16262) );
  OAI21_X1 U19212 ( .B1(n16263), .B2(n16275), .A(n16262), .ZN(U241) );
  INV_X1 U19213 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16282) );
  AOI22_X1 U19214 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16270), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16273), .ZN(n16264) );
  OAI21_X1 U19215 ( .B1(n16282), .B2(U212), .A(n16264), .ZN(U242) );
  INV_X1 U19216 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16266) );
  AOI22_X1 U19217 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16272), .ZN(n16265) );
  OAI21_X1 U19218 ( .B1(n16266), .B2(n16275), .A(n16265), .ZN(U243) );
  INV_X1 U19219 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16280) );
  AOI22_X1 U19220 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16270), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16273), .ZN(n16267) );
  OAI21_X1 U19221 ( .B1(n16280), .B2(U212), .A(n16267), .ZN(U244) );
  INV_X1 U19222 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16269) );
  AOI22_X1 U19223 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16272), .ZN(n16268) );
  OAI21_X1 U19224 ( .B1(n16269), .B2(n16275), .A(n16268), .ZN(U245) );
  INV_X1 U19225 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16278) );
  AOI22_X1 U19226 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16270), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16273), .ZN(n16271) );
  OAI21_X1 U19227 ( .B1(n16278), .B2(U212), .A(n16271), .ZN(U246) );
  INV_X1 U19228 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16276) );
  AOI22_X1 U19229 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16273), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16272), .ZN(n16274) );
  OAI21_X1 U19230 ( .B1(n16276), .B2(n16275), .A(n16274), .ZN(U247) );
  OAI22_X1 U19231 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16307), .ZN(n16277) );
  INV_X1 U19232 ( .A(n16277), .ZN(U251) );
  INV_X1 U19233 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n20751) );
  AOI22_X1 U19234 ( .A1(n16307), .A2(n16278), .B1(n20751), .B2(U215), .ZN(U252) );
  OAI22_X1 U19235 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16299), .ZN(n16279) );
  INV_X1 U19236 ( .A(n16279), .ZN(U253) );
  INV_X1 U19237 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n17999) );
  AOI22_X1 U19238 ( .A1(n16307), .A2(n16280), .B1(n17999), .B2(U215), .ZN(U254) );
  OAI22_X1 U19239 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16299), .ZN(n16281) );
  INV_X1 U19240 ( .A(n16281), .ZN(U255) );
  INV_X1 U19241 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18012) );
  AOI22_X1 U19242 ( .A1(n16307), .A2(n16282), .B1(n18012), .B2(U215), .ZN(U256) );
  OAI22_X1 U19243 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16299), .ZN(n16283) );
  INV_X1 U19244 ( .A(n16283), .ZN(U257) );
  INV_X1 U19245 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18021) );
  AOI22_X1 U19246 ( .A1(n16307), .A2(n16284), .B1(n18021), .B2(U215), .ZN(U258) );
  OAI22_X1 U19247 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16299), .ZN(n16285) );
  INV_X1 U19248 ( .A(n16285), .ZN(U259) );
  INV_X1 U19249 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n20735) );
  INV_X1 U19250 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17253) );
  AOI22_X1 U19251 ( .A1(n16307), .A2(n20735), .B1(n17253), .B2(U215), .ZN(U260) );
  OAI22_X1 U19252 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16299), .ZN(n16286) );
  INV_X1 U19253 ( .A(n16286), .ZN(U261) );
  INV_X1 U19254 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17257) );
  AOI22_X1 U19255 ( .A1(n16307), .A2(n16287), .B1(n17257), .B2(U215), .ZN(U262) );
  OAI22_X1 U19256 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16299), .ZN(n16288) );
  INV_X1 U19257 ( .A(n16288), .ZN(U263) );
  OAI22_X1 U19258 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16299), .ZN(n16289) );
  INV_X1 U19259 ( .A(n16289), .ZN(U264) );
  OAI22_X1 U19260 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16307), .ZN(n16290) );
  INV_X1 U19261 ( .A(n16290), .ZN(U265) );
  OAI22_X1 U19262 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16299), .ZN(n16291) );
  INV_X1 U19263 ( .A(n16291), .ZN(U266) );
  OAI22_X1 U19264 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16307), .ZN(n16292) );
  INV_X1 U19265 ( .A(n16292), .ZN(U267) );
  OAI22_X1 U19266 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16299), .ZN(n16293) );
  INV_X1 U19267 ( .A(n16293), .ZN(U268) );
  OAI22_X1 U19268 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16307), .ZN(n16294) );
  INV_X1 U19269 ( .A(n16294), .ZN(U269) );
  OAI22_X1 U19270 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16307), .ZN(n16295) );
  INV_X1 U19271 ( .A(n16295), .ZN(U270) );
  OAI22_X1 U19272 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16307), .ZN(n16296) );
  INV_X1 U19273 ( .A(n16296), .ZN(U271) );
  OAI22_X1 U19274 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16307), .ZN(n16297) );
  INV_X1 U19275 ( .A(n16297), .ZN(U272) );
  OAI22_X1 U19276 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16307), .ZN(n16298) );
  INV_X1 U19277 ( .A(n16298), .ZN(U273) );
  OAI22_X1 U19278 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16299), .ZN(n16300) );
  INV_X1 U19279 ( .A(n16300), .ZN(U274) );
  OAI22_X1 U19280 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16307), .ZN(n16301) );
  INV_X1 U19281 ( .A(n16301), .ZN(U275) );
  OAI22_X1 U19282 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16307), .ZN(n16302) );
  INV_X1 U19283 ( .A(n16302), .ZN(U276) );
  OAI22_X1 U19284 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16307), .ZN(n16303) );
  INV_X1 U19285 ( .A(n16303), .ZN(U277) );
  OAI22_X1 U19286 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16307), .ZN(n16304) );
  INV_X1 U19287 ( .A(n16304), .ZN(U278) );
  OAI22_X1 U19288 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16307), .ZN(n16305) );
  INV_X1 U19289 ( .A(n16305), .ZN(U279) );
  INV_X1 U19290 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n20776) );
  INV_X1 U19291 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18011) );
  AOI22_X1 U19292 ( .A1(n16307), .A2(n20776), .B1(n18011), .B2(U215), .ZN(U280) );
  OAI22_X1 U19293 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16307), .ZN(n16306) );
  INV_X1 U19294 ( .A(n16306), .ZN(U281) );
  INV_X1 U19295 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19064) );
  AOI22_X1 U19296 ( .A1(n16307), .A2(n18974), .B1(n19064), .B2(U215), .ZN(U282) );
  INV_X1 U19297 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17165) );
  AOI222_X1 U19298 ( .A1(n16308), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n18974), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n17165), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16309) );
  INV_X2 U19299 ( .A(n16311), .ZN(n16310) );
  INV_X1 U19300 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18529) );
  INV_X1 U19301 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19634) );
  AOI22_X1 U19302 ( .A1(n16310), .A2(n18529), .B1(n19634), .B2(n16311), .ZN(
        U347) );
  INV_X1 U19303 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18527) );
  INV_X1 U19304 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19633) );
  AOI22_X1 U19305 ( .A1(n16310), .A2(n18527), .B1(n19633), .B2(n16311), .ZN(
        U348) );
  INV_X1 U19306 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18525) );
  INV_X1 U19307 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19632) );
  AOI22_X1 U19308 ( .A1(n16310), .A2(n18525), .B1(n19632), .B2(n16311), .ZN(
        U349) );
  INV_X1 U19309 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18523) );
  INV_X1 U19310 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19631) );
  AOI22_X1 U19311 ( .A1(n16310), .A2(n18523), .B1(n19631), .B2(n16311), .ZN(
        U350) );
  INV_X1 U19312 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18522) );
  INV_X1 U19313 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19630) );
  AOI22_X1 U19314 ( .A1(n16310), .A2(n18522), .B1(n19630), .B2(n16311), .ZN(
        U351) );
  INV_X1 U19315 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18519) );
  INV_X1 U19316 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19629) );
  AOI22_X1 U19317 ( .A1(n16310), .A2(n18519), .B1(n19629), .B2(n16311), .ZN(
        U352) );
  INV_X1 U19318 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18517) );
  INV_X1 U19319 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19628) );
  AOI22_X1 U19320 ( .A1(n16310), .A2(n18517), .B1(n19628), .B2(n16311), .ZN(
        U353) );
  INV_X1 U19321 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18515) );
  AOI22_X1 U19322 ( .A1(n16310), .A2(n18515), .B1(n19627), .B2(n16311), .ZN(
        U354) );
  INV_X1 U19323 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18573) );
  INV_X1 U19324 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19663) );
  AOI22_X1 U19325 ( .A1(n16310), .A2(n18573), .B1(n19663), .B2(n16311), .ZN(
        U355) );
  INV_X1 U19326 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18570) );
  INV_X1 U19327 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19660) );
  AOI22_X1 U19328 ( .A1(n16310), .A2(n18570), .B1(n19660), .B2(n16311), .ZN(
        U356) );
  INV_X1 U19329 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18566) );
  INV_X1 U19330 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20719) );
  AOI22_X1 U19331 ( .A1(n16310), .A2(n18566), .B1(n20719), .B2(n16311), .ZN(
        U357) );
  INV_X1 U19332 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18564) );
  INV_X1 U19333 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19657) );
  AOI22_X1 U19334 ( .A1(n16310), .A2(n18564), .B1(n19657), .B2(n16311), .ZN(
        U358) );
  INV_X1 U19335 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18562) );
  INV_X1 U19336 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19656) );
  AOI22_X1 U19337 ( .A1(n16310), .A2(n18562), .B1(n19656), .B2(n16311), .ZN(
        U359) );
  INV_X1 U19338 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18560) );
  INV_X1 U19339 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19655) );
  AOI22_X1 U19340 ( .A1(n16310), .A2(n18560), .B1(n19655), .B2(n16311), .ZN(
        U360) );
  INV_X1 U19341 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18558) );
  INV_X1 U19342 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19653) );
  AOI22_X1 U19343 ( .A1(n16310), .A2(n18558), .B1(n19653), .B2(n16311), .ZN(
        U361) );
  INV_X1 U19344 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18555) );
  INV_X1 U19345 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19652) );
  AOI22_X1 U19346 ( .A1(n16310), .A2(n18555), .B1(n19652), .B2(n16311), .ZN(
        U362) );
  INV_X1 U19347 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18554) );
  INV_X1 U19348 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19651) );
  AOI22_X1 U19349 ( .A1(n16310), .A2(n18554), .B1(n19651), .B2(n16311), .ZN(
        U363) );
  INV_X1 U19350 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18551) );
  INV_X1 U19351 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19650) );
  AOI22_X1 U19352 ( .A1(n16310), .A2(n18551), .B1(n19650), .B2(n16311), .ZN(
        U364) );
  INV_X1 U19353 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18513) );
  INV_X1 U19354 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19626) );
  AOI22_X1 U19355 ( .A1(n16310), .A2(n18513), .B1(n19626), .B2(n16311), .ZN(
        U365) );
  INV_X1 U19356 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18550) );
  INV_X1 U19357 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19648) );
  AOI22_X1 U19358 ( .A1(n16310), .A2(n18550), .B1(n19648), .B2(n16311), .ZN(
        U366) );
  INV_X1 U19359 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18548) );
  INV_X1 U19360 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19646) );
  AOI22_X1 U19361 ( .A1(n16310), .A2(n18548), .B1(n19646), .B2(n16311), .ZN(
        U367) );
  INV_X1 U19362 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18546) );
  INV_X1 U19363 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19644) );
  AOI22_X1 U19364 ( .A1(n16310), .A2(n18546), .B1(n19644), .B2(n16311), .ZN(
        U368) );
  INV_X1 U19365 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18543) );
  INV_X1 U19366 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19642) );
  AOI22_X1 U19367 ( .A1(n16310), .A2(n18543), .B1(n19642), .B2(n16311), .ZN(
        U369) );
  INV_X1 U19368 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18541) );
  INV_X1 U19369 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19640) );
  AOI22_X1 U19370 ( .A1(n16310), .A2(n18541), .B1(n19640), .B2(n16311), .ZN(
        U370) );
  INV_X1 U19371 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18539) );
  INV_X1 U19372 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19639) );
  AOI22_X1 U19373 ( .A1(n16310), .A2(n18539), .B1(n19639), .B2(n16311), .ZN(
        U371) );
  INV_X1 U19374 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18537) );
  INV_X1 U19375 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19638) );
  AOI22_X1 U19376 ( .A1(n16310), .A2(n18537), .B1(n19638), .B2(n16311), .ZN(
        U372) );
  INV_X1 U19377 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18536) );
  INV_X1 U19378 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19637) );
  AOI22_X1 U19379 ( .A1(n16310), .A2(n18536), .B1(n19637), .B2(n16311), .ZN(
        U373) );
  INV_X1 U19380 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18533) );
  INV_X1 U19381 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19636) );
  AOI22_X1 U19382 ( .A1(n16310), .A2(n18533), .B1(n19636), .B2(n16311), .ZN(
        U374) );
  INV_X1 U19383 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18531) );
  INV_X1 U19384 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19635) );
  AOI22_X1 U19385 ( .A1(n16310), .A2(n18531), .B1(n19635), .B2(n16311), .ZN(
        U375) );
  INV_X1 U19386 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18512) );
  INV_X1 U19387 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19625) );
  AOI22_X1 U19388 ( .A1(n16310), .A2(n18512), .B1(n19625), .B2(n16311), .ZN(
        U376) );
  INV_X1 U19389 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18511) );
  NAND2_X1 U19390 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18511), .ZN(n18499) );
  AOI22_X1 U19391 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18499), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18509), .ZN(n18583) );
  AOI21_X1 U19392 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18583), .ZN(n16312) );
  INV_X1 U19393 ( .A(n16312), .ZN(P3_U2633) );
  INV_X1 U19394 ( .A(n16317), .ZN(n18424) );
  NOR2_X1 U19395 ( .A1(n16318), .A2(n17224), .ZN(n16313) );
  OAI21_X1 U19396 ( .B1(n17164), .B2(n16313), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16314) );
  INV_X1 U19397 ( .A(n18593), .ZN(n18647) );
  NAND3_X1 U19398 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18647), .A3(n18646), 
        .ZN(n18489) );
  NAND2_X1 U19399 ( .A1(n16314), .A2(n18489), .ZN(P3_U2634) );
  AOI21_X1 U19400 ( .B1(n18509), .B2(n18511), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16315) );
  AOI22_X1 U19401 ( .A1(n18640), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16315), 
        .B2(n18641), .ZN(P3_U2635) );
  OAI21_X1 U19402 ( .B1(n18496), .B2(BS16), .A(n18583), .ZN(n18581) );
  OAI21_X1 U19403 ( .B1(n18583), .B2(n18630), .A(n18581), .ZN(P3_U2636) );
  OAI211_X1 U19404 ( .C1(n16318), .C2(n17224), .A(n16317), .B(n16316), .ZN(
        n16319) );
  INV_X1 U19405 ( .A(n16319), .ZN(n18429) );
  NOR2_X1 U19406 ( .A1(n18429), .A2(n18490), .ZN(n18623) );
  OAI21_X1 U19407 ( .B1(n18623), .B2(n17972), .A(n16320), .ZN(P3_U2637) );
  NOR4_X1 U19408 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16324) );
  NOR4_X1 U19409 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16323) );
  NOR4_X1 U19410 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16322) );
  NOR4_X1 U19411 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16321) );
  NAND4_X1 U19412 ( .A1(n16324), .A2(n16323), .A3(n16322), .A4(n16321), .ZN(
        n16330) );
  NOR4_X1 U19413 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n16328) );
  AOI211_X1 U19414 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_9__SCAN_IN), .B(
        P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(n16327) );
  NOR4_X1 U19415 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16326) );
  NOR4_X1 U19416 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16325) );
  NAND4_X1 U19417 ( .A1(n16328), .A2(n16327), .A3(n16326), .A4(n16325), .ZN(
        n16329) );
  NOR2_X1 U19418 ( .A1(n16330), .A2(n16329), .ZN(n18621) );
  INV_X1 U19419 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16332) );
  NOR3_X1 U19420 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16333) );
  OAI21_X1 U19421 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16333), .A(n18621), .ZN(
        n16331) );
  OAI21_X1 U19422 ( .B1(n18621), .B2(n16332), .A(n16331), .ZN(P3_U2638) );
  INV_X1 U19423 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18614) );
  INV_X1 U19424 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18582) );
  AOI21_X1 U19425 ( .B1(n18614), .B2(n18582), .A(n16333), .ZN(n16335) );
  INV_X1 U19426 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16334) );
  INV_X1 U19427 ( .A(n18621), .ZN(n18616) );
  AOI22_X1 U19428 ( .A1(n18621), .A2(n16335), .B1(n16334), .B2(n18616), .ZN(
        P3_U2639) );
  NOR2_X1 U19429 ( .A1(n18586), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18358) );
  INV_X1 U19430 ( .A(n18358), .ZN(n18250) );
  NOR2_X1 U19431 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18250), .ZN(n18479) );
  NOR3_X1 U19432 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n18494) );
  NAND2_X1 U19433 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18494), .ZN(n20816) );
  INV_X1 U19434 ( .A(n20816), .ZN(n18487) );
  AOI211_X1 U19435 ( .C1(P3_STATE2_REG_0__SCAN_IN), .C2(n18479), .A(n18487), 
        .B(n18651), .ZN(n16336) );
  INV_X1 U19436 ( .A(n18632), .ZN(n18504) );
  AOI211_X1 U19437 ( .C1(n18631), .C2(n18629), .A(n18504), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18474) );
  INV_X1 U19438 ( .A(n18651), .ZN(n18643) );
  INV_X1 U19439 ( .A(n16337), .ZN(n18648) );
  AOI211_X4 U19440 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n17991), .A(n18474), .B(
        n18648), .ZN(n20834) );
  INV_X1 U19441 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18574) );
  INV_X1 U19442 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18559) );
  INV_X1 U19443 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18556) );
  INV_X1 U19444 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18552) );
  INV_X1 U19445 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18547) );
  NAND3_X1 U19446 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .A3(P3_REIP_REG_3__SCAN_IN), .ZN(n16650) );
  INV_X1 U19447 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18518) );
  INV_X1 U19448 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18520) );
  NOR3_X1 U19449 ( .A1(n16650), .A2(n18518), .A3(n18520), .ZN(n16566) );
  NAND2_X1 U19450 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n16598) );
  INV_X1 U19451 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18526) );
  NOR2_X1 U19452 ( .A1(n16598), .A2(n18526), .ZN(n16555) );
  NAND2_X1 U19453 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n16577) );
  INV_X1 U19454 ( .A(n16577), .ZN(n16556) );
  NAND4_X1 U19455 ( .A1(n16566), .A2(n16555), .A3(n16556), .A4(
        P3_REIP_REG_11__SCAN_IN), .ZN(n16549) );
  INV_X1 U19456 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18534) );
  NOR2_X1 U19457 ( .A1(n16549), .A2(n18534), .ZN(n16521) );
  NAND3_X1 U19458 ( .A1(n16521), .A2(P3_REIP_REG_14__SCAN_IN), .A3(
        P3_REIP_REG_13__SCAN_IN), .ZN(n16522) );
  INV_X1 U19459 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18540) );
  NOR2_X1 U19460 ( .A1(n16522), .A2(n18540), .ZN(n16497) );
  NAND2_X1 U19461 ( .A1(n16497), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n16483) );
  INV_X1 U19462 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18544) );
  NOR2_X1 U19463 ( .A1(n16483), .A2(n18544), .ZN(n16463) );
  NAND2_X1 U19464 ( .A1(n16463), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n16464) );
  NOR2_X1 U19465 ( .A1(n18547), .A2(n16464), .ZN(n20828) );
  NAND2_X1 U19466 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n20828), .ZN(n20826) );
  NOR2_X1 U19467 ( .A1(n18552), .A2(n20826), .ZN(n16443) );
  NAND2_X1 U19468 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16443), .ZN(n16434) );
  NOR2_X1 U19469 ( .A1(n18556), .A2(n16434), .ZN(n16432) );
  NAND2_X1 U19470 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16432), .ZN(n16411) );
  NOR2_X1 U19471 ( .A1(n18559), .A2(n16411), .ZN(n16399) );
  NAND2_X1 U19472 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16399), .ZN(n16351) );
  NOR2_X1 U19473 ( .A1(n16691), .A2(n16351), .ZN(n16393) );
  NAND4_X1 U19474 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16393), .ZN(n16353) );
  NOR3_X1 U19475 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18574), .A3(n16353), 
        .ZN(n16338) );
  AOI21_X1 U19476 ( .B1(n20834), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16338), .ZN(
        n16357) );
  NAND2_X1 U19477 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n17991), .ZN(n16339) );
  AOI211_X4 U19478 ( .C1(n18630), .C2(n18632), .A(n18648), .B(n16339), .ZN(
        n16696) );
  NOR3_X1 U19479 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n16685) );
  NAND2_X1 U19480 ( .A1(n16685), .A2(n16668), .ZN(n16667) );
  NOR2_X1 U19481 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16667), .ZN(n16645) );
  INV_X1 U19482 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16639) );
  NAND2_X1 U19483 ( .A1(n16645), .A2(n16639), .ZN(n16638) );
  NAND2_X1 U19484 ( .A1(n16624), .A2(n16610), .ZN(n16609) );
  NAND2_X1 U19485 ( .A1(n16584), .A2(n16587), .ZN(n16572) );
  NAND2_X1 U19486 ( .A1(n16571), .A2(n16563), .ZN(n16562) );
  INV_X1 U19487 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16539) );
  NAND2_X1 U19488 ( .A1(n16543), .A2(n16539), .ZN(n16536) );
  INV_X1 U19489 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16518) );
  NAND2_X1 U19490 ( .A1(n16520), .A2(n16518), .ZN(n16512) );
  INV_X1 U19491 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16494) );
  NAND2_X1 U19492 ( .A1(n16496), .A2(n16494), .ZN(n16487) );
  INV_X1 U19493 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16822) );
  NAND2_X1 U19494 ( .A1(n16477), .A2(n16822), .ZN(n20822) );
  INV_X1 U19495 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16797) );
  NAND2_X1 U19496 ( .A1(n20821), .A2(n16797), .ZN(n16457) );
  NAND2_X1 U19497 ( .A1(n16444), .A2(n16438), .ZN(n16437) );
  NAND2_X1 U19498 ( .A1(n16421), .A2(n16416), .ZN(n16415) );
  NOR2_X1 U19499 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16415), .ZN(n16400) );
  NAND2_X1 U19500 ( .A1(n16400), .A2(n16747), .ZN(n16394) );
  NOR2_X1 U19501 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16394), .ZN(n16378) );
  INV_X1 U19502 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16374) );
  NAND2_X1 U19503 ( .A1(n16378), .A2(n16374), .ZN(n16358) );
  NOR2_X1 U19504 ( .A1(n20820), .A2(n16358), .ZN(n16362) );
  INV_X1 U19505 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16712) );
  AOI21_X1 U19506 ( .B1(n16340), .B2(n16390), .A(n16350), .ZN(n17293) );
  NOR2_X1 U19507 ( .A1(n17639), .A2(n17339), .ZN(n16343) );
  NAND2_X1 U19508 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n16343), .ZN(
        n16348) );
  INV_X1 U19509 ( .A(n16348), .ZN(n16342) );
  NAND3_X1 U19510 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(n16342), .ZN(n17278) );
  AOI21_X1 U19511 ( .B1(n17304), .B2(n17278), .A(n16341), .ZN(n17306) );
  INV_X1 U19512 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17317) );
  NOR2_X1 U19513 ( .A1(n17317), .A2(n16348), .ZN(n16347) );
  OAI21_X1 U19514 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16347), .A(
        n17278), .ZN(n17319) );
  INV_X1 U19515 ( .A(n17319), .ZN(n16410) );
  INV_X1 U19516 ( .A(n16343), .ZN(n17344) );
  AOI21_X1 U19517 ( .B1(n17341), .B2(n17344), .A(n16342), .ZN(n17348) );
  INV_X1 U19518 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17361) );
  NOR3_X1 U19519 ( .A1(n17639), .A2(n17422), .A3(n17421), .ZN(n17393) );
  NAND3_X1 U19520 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A3(n17393), .ZN(n17358) );
  NOR2_X1 U19521 ( .A1(n20831), .A2(n17358), .ZN(n16346) );
  NAND2_X1 U19522 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16346), .ZN(
        n16344) );
  AOI21_X1 U19523 ( .B1(n17361), .B2(n16344), .A(n16343), .ZN(n17359) );
  AOI21_X1 U19524 ( .B1(n20831), .B2(n17358), .A(n16346), .ZN(n20819) );
  INV_X1 U19525 ( .A(n17358), .ZN(n16345) );
  NOR2_X1 U19526 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17639), .ZN(
        n16674) );
  AND2_X1 U19527 ( .A1(n17433), .A2(n16674), .ZN(n16509) );
  NAND2_X1 U19528 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n16509), .ZN(
        n16503) );
  INV_X1 U19529 ( .A(n16503), .ZN(n16474) );
  AOI21_X1 U19530 ( .B1(n16345), .B2(n16474), .A(n16659), .ZN(n20818) );
  NOR2_X1 U19531 ( .A1(n20819), .A2(n20818), .ZN(n20817) );
  NOR2_X1 U19532 ( .A1(n20817), .A2(n16659), .ZN(n16452) );
  INV_X1 U19533 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17360) );
  XOR2_X1 U19534 ( .A(n17360), .B(n16346), .Z(n17373) );
  INV_X1 U19535 ( .A(n17373), .ZN(n16453) );
  NOR2_X1 U19536 ( .A1(n16430), .A2(n16659), .ZN(n16424) );
  AOI21_X1 U19537 ( .B1(n17317), .B2(n16348), .A(n16347), .ZN(n17331) );
  NOR2_X1 U19538 ( .A1(n16410), .A2(n16409), .ZN(n16408) );
  NOR2_X1 U19539 ( .A1(n16408), .A2(n16659), .ZN(n16402) );
  OAI21_X1 U19540 ( .B1(n16350), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16349), .ZN(n17281) );
  INV_X1 U19541 ( .A(n17281), .ZN(n16382) );
  NOR2_X1 U19542 ( .A1(n16659), .A2(n20816), .ZN(n16689) );
  INV_X1 U19543 ( .A(n16689), .ZN(n16605) );
  NOR3_X1 U19544 ( .A1(n16360), .A2(n16359), .A3(n16605), .ZN(n16355) );
  NAND3_X1 U19545 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16352) );
  AND2_X1 U19546 ( .A1(n20827), .A2(n16351), .ZN(n16398) );
  NOR2_X1 U19547 ( .A1(n20825), .A2(n16398), .ZN(n16397) );
  INV_X1 U19548 ( .A(n16397), .ZN(n16405) );
  AOI21_X1 U19549 ( .B1(n20827), .B2(n16352), .A(n16405), .ZN(n16377) );
  AOI21_X1 U19550 ( .B1(n16377), .B2(n9729), .A(n18572), .ZN(n16354) );
  AOI211_X1 U19551 ( .C1(n16362), .C2(n16712), .A(n16355), .B(n16354), .ZN(
        n16356) );
  OAI211_X1 U19552 ( .C1(n9880), .C2(n20832), .A(n16357), .B(n16356), .ZN(
        P3_U2640) );
  NAND2_X1 U19553 ( .A1(n16696), .A2(n16358), .ZN(n16372) );
  OAI22_X1 U19554 ( .A1(n16377), .A2(n18574), .B1(n9885), .B2(n20832), .ZN(
        n16361) );
  OAI21_X1 U19555 ( .B1(n20834), .B2(n16362), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16363) );
  OAI211_X1 U19556 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16372), .A(n16364), .B(
        n16363), .ZN(P3_U2641) );
  INV_X1 U19557 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18569) );
  AOI211_X1 U19558 ( .C1(n16367), .C2(n16366), .A(n16365), .B(n20816), .ZN(
        n16371) );
  NAND3_X1 U19559 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16393), .ZN(n16369) );
  OAI22_X1 U19560 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16369), .B1(n16368), 
        .B2(n20832), .ZN(n16370) );
  AOI211_X1 U19561 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n20834), .A(n16371), .B(
        n16370), .ZN(n16376) );
  INV_X1 U19562 ( .A(n16372), .ZN(n16373) );
  OAI21_X1 U19563 ( .B1(n16378), .B2(n16374), .A(n16373), .ZN(n16375) );
  OAI211_X1 U19564 ( .C1(n16377), .C2(n18569), .A(n16376), .B(n16375), .ZN(
        P3_U2642) );
  AOI22_X1 U19565 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16688), .B1(
        n20834), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16388) );
  AOI211_X1 U19566 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16394), .A(n16378), .B(
        n20820), .ZN(n16384) );
  INV_X1 U19567 ( .A(n16379), .ZN(n16380) );
  AOI211_X1 U19568 ( .C1(n16382), .C2(n16381), .A(n16380), .B(n20816), .ZN(
        n16383) );
  AOI211_X1 U19569 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16405), .A(n16384), 
        .B(n16383), .ZN(n16387) );
  NAND2_X1 U19570 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16385) );
  OAI211_X1 U19571 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16393), .B(n16385), .ZN(n16386) );
  NAND3_X1 U19572 ( .A1(n16388), .A2(n16387), .A3(n16386), .ZN(P3_U2643) );
  INV_X1 U19573 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18563) );
  AOI211_X1 U19574 ( .C1(n17293), .C2(n16389), .A(n9740), .B(n20816), .ZN(
        n16392) );
  OAI22_X1 U19575 ( .A1(n16390), .A2(n20832), .B1(n16700), .B2(n16747), .ZN(
        n16391) );
  AOI211_X1 U19576 ( .C1(n16393), .C2(n18563), .A(n16392), .B(n16391), .ZN(
        n16396) );
  OAI211_X1 U19577 ( .C1(n16400), .C2(n16747), .A(n16696), .B(n16394), .ZN(
        n16395) );
  OAI211_X1 U19578 ( .C1(n16397), .C2(n18563), .A(n16396), .B(n16395), .ZN(
        P3_U2644) );
  AOI22_X1 U19579 ( .A1(n20834), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n16399), 
        .B2(n16398), .ZN(n16407) );
  AOI211_X1 U19580 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16415), .A(n16400), .B(
        n20820), .ZN(n16404) );
  AOI211_X1 U19581 ( .C1(n17306), .C2(n16402), .A(n16401), .B(n20816), .ZN(
        n16403) );
  AOI211_X1 U19582 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16405), .A(n16404), 
        .B(n16403), .ZN(n16406) );
  OAI211_X1 U19583 ( .C1(n17304), .C2(n20832), .A(n16407), .B(n16406), .ZN(
        P3_U2645) );
  INV_X1 U19584 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18557) );
  OAI21_X1 U19585 ( .B1(n16432), .B2(n16691), .A(n16703), .ZN(n16429) );
  AOI21_X1 U19586 ( .B1(n20827), .B2(n18557), .A(n16429), .ZN(n16419) );
  AOI211_X1 U19587 ( .C1(n16410), .C2(n16409), .A(n16408), .B(n20816), .ZN(
        n16414) );
  NOR3_X1 U19588 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16691), .A3(n16411), 
        .ZN(n16413) );
  INV_X1 U19589 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17318) );
  OAI22_X1 U19590 ( .A1(n17318), .A2(n20832), .B1(n16700), .B2(n16416), .ZN(
        n16412) );
  NOR3_X1 U19591 ( .A1(n16414), .A2(n16413), .A3(n16412), .ZN(n16418) );
  OAI211_X1 U19592 ( .C1(n16421), .C2(n16416), .A(n16696), .B(n16415), .ZN(
        n16417) );
  OAI211_X1 U19593 ( .C1(n16419), .C2(n18559), .A(n16418), .B(n16417), .ZN(
        P3_U2646) );
  NOR2_X1 U19594 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16691), .ZN(n16420) );
  AOI22_X1 U19595 ( .A1(n20834), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16432), 
        .B2(n16420), .ZN(n16428) );
  AOI211_X1 U19596 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16437), .A(n16421), .B(
        n20820), .ZN(n16426) );
  INV_X1 U19597 ( .A(n16422), .ZN(n16423) );
  AOI211_X1 U19598 ( .C1(n17331), .C2(n16424), .A(n16423), .B(n20816), .ZN(
        n16425) );
  AOI211_X1 U19599 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16429), .A(n16426), 
        .B(n16425), .ZN(n16427) );
  OAI211_X1 U19600 ( .C1(n17317), .C2(n20832), .A(n16428), .B(n16427), .ZN(
        P3_U2647) );
  INV_X1 U19601 ( .A(n16429), .ZN(n16441) );
  AOI211_X1 U19602 ( .C1(n17348), .C2(n16431), .A(n16430), .B(n20816), .ZN(
        n16436) );
  OR2_X1 U19603 ( .A1(n16691), .A2(n16432), .ZN(n16433) );
  OAI22_X1 U19604 ( .A1(n16700), .A2(n16438), .B1(n16434), .B2(n16433), .ZN(
        n16435) );
  AOI211_X1 U19605 ( .C1(n16688), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16436), .B(n16435), .ZN(n16440) );
  OAI211_X1 U19606 ( .C1(n16444), .C2(n16438), .A(n16696), .B(n16437), .ZN(
        n16439) );
  OAI211_X1 U19607 ( .C1(n16441), .C2(n18556), .A(n16440), .B(n16439), .ZN(
        P3_U2648) );
  NOR4_X1 U19608 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16691), .A3(n18552), 
        .A4(n20826), .ZN(n16442) );
  AOI21_X1 U19609 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n20834), .A(n16442), .ZN(
        n16449) );
  OAI21_X1 U19610 ( .B1(n16443), .B2(n16691), .A(n16703), .ZN(n16456) );
  AOI211_X1 U19611 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16457), .A(n16444), .B(
        n20820), .ZN(n16447) );
  AOI211_X1 U19612 ( .C1(n17359), .C2(n16445), .A(n9749), .B(n20816), .ZN(
        n16446) );
  AOI211_X1 U19613 ( .C1(n16456), .C2(P3_REIP_REG_22__SCAN_IN), .A(n16447), 
        .B(n16446), .ZN(n16448) );
  OAI211_X1 U19614 ( .C1(n17361), .C2(n20832), .A(n16449), .B(n16448), .ZN(
        P3_U2649) );
  AOI22_X1 U19615 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16688), .B1(
        n20834), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n16460) );
  NOR2_X1 U19616 ( .A1(n16691), .A2(n20826), .ZN(n16455) );
  INV_X1 U19617 ( .A(n16450), .ZN(n16451) );
  AOI211_X1 U19618 ( .C1(n16453), .C2(n16452), .A(n16451), .B(n20816), .ZN(
        n16454) );
  AOI221_X1 U19619 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16456), .C1(n16455), 
        .C2(n16456), .A(n16454), .ZN(n16459) );
  OAI211_X1 U19620 ( .C1(n20821), .C2(n16797), .A(n16696), .B(n16457), .ZN(
        n16458) );
  NAND3_X1 U19621 ( .A1(n16460), .A2(n16459), .A3(n16458), .ZN(P3_U2650) );
  NAND2_X1 U19622 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17393), .ZN(
        n16473) );
  INV_X1 U19623 ( .A(n16473), .ZN(n16461) );
  OAI21_X1 U19624 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16461), .A(
        n17358), .ZN(n17394) );
  AOI21_X1 U19625 ( .B1(n16461), .B2(n16474), .A(n16659), .ZN(n16462) );
  XOR2_X1 U19626 ( .A(n17394), .B(n16462), .Z(n16471) );
  NOR4_X1 U19627 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16483), .A3(n16691), 
        .A4(n18544), .ZN(n16472) );
  OAI21_X1 U19628 ( .B1(n16463), .B2(n16691), .A(n16703), .ZN(n16492) );
  INV_X1 U19629 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16468) );
  NOR3_X1 U19630 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16691), .A3(n16464), 
        .ZN(n16465) );
  AOI211_X1 U19631 ( .C1(n20834), .C2(P3_EBX_REG_19__SCAN_IN), .A(n17965), .B(
        n16465), .ZN(n16467) );
  OAI211_X1 U19632 ( .C1(n16477), .C2(n16822), .A(n16696), .B(n20822), .ZN(
        n16466) );
  OAI211_X1 U19633 ( .C1(n20832), .C2(n16468), .A(n16467), .B(n16466), .ZN(
        n16469) );
  AOI221_X1 U19634 ( .B1(n16472), .B2(P3_REIP_REG_19__SCAN_IN), .C1(n16492), 
        .C2(P3_REIP_REG_19__SCAN_IN), .A(n16469), .ZN(n16470) );
  OAI21_X1 U19635 ( .B1(n20816), .B2(n16471), .A(n16470), .ZN(P3_U2652) );
  INV_X1 U19636 ( .A(n16492), .ZN(n16482) );
  INV_X1 U19637 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18545) );
  AOI211_X1 U19638 ( .C1(n20834), .C2(P3_EBX_REG_18__SCAN_IN), .A(n11114), .B(
        n16472), .ZN(n16481) );
  OAI21_X1 U19639 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17393), .A(
        n16473), .ZN(n17409) );
  AOI21_X1 U19640 ( .B1(n17393), .B2(n16474), .A(n16659), .ZN(n16486) );
  INV_X1 U19641 ( .A(n16486), .ZN(n16476) );
  OAI21_X1 U19642 ( .B1(n17409), .B2(n16476), .A(n18487), .ZN(n16475) );
  AOI21_X1 U19643 ( .B1(n17409), .B2(n16476), .A(n16475), .ZN(n16479) );
  AOI211_X1 U19644 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16487), .A(n16477), .B(
        n20820), .ZN(n16478) );
  AOI211_X1 U19645 ( .C1(n16688), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16479), .B(n16478), .ZN(n16480) );
  OAI211_X1 U19646 ( .C1(n16482), .C2(n18545), .A(n16481), .B(n16480), .ZN(
        P3_U2653) );
  NOR2_X1 U19647 ( .A1(n16691), .A2(n16483), .ZN(n16491) );
  OR2_X1 U19648 ( .A1(n17639), .A2(n17422), .ZN(n16484) );
  AOI21_X1 U19649 ( .B1(n17421), .B2(n16484), .A(n17393), .ZN(n17424) );
  NOR2_X1 U19650 ( .A1(n20816), .A2(n9732), .ZN(n16686) );
  AOI221_X1 U19651 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n17424), .C1(
        n16503), .C2(n17424), .A(n20816), .ZN(n16485) );
  OAI22_X1 U19652 ( .A1(n17424), .A2(n16486), .B1(n16686), .B2(n16485), .ZN(
        n16489) );
  OAI211_X1 U19653 ( .C1(n16496), .C2(n16494), .A(n16696), .B(n16487), .ZN(
        n16488) );
  OAI211_X1 U19654 ( .C1(n20832), .C2(n17421), .A(n16489), .B(n16488), .ZN(
        n16490) );
  AOI221_X1 U19655 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n16492), .C1(n16491), 
        .C2(n16492), .A(n16490), .ZN(n16493) );
  OAI211_X1 U19656 ( .C1(n16700), .C2(n16494), .A(n16493), .B(n17963), .ZN(
        P3_U2654) );
  OAI21_X1 U19657 ( .B1(n16691), .B2(n16497), .A(n16703), .ZN(n16495) );
  INV_X1 U19658 ( .A(n16495), .ZN(n16508) );
  INV_X1 U19659 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18542) );
  AOI211_X1 U19660 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16512), .A(n16496), .B(
        n20820), .ZN(n16500) );
  NAND3_X1 U19661 ( .A1(n16497), .A2(n20827), .A3(n18542), .ZN(n16498) );
  OAI211_X1 U19662 ( .C1(n16700), .C2(n16854), .A(n17963), .B(n16498), .ZN(
        n16499) );
  AOI211_X1 U19663 ( .C1(n16688), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16500), .B(n16499), .ZN(n16507) );
  INV_X1 U19664 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17448) );
  AND2_X1 U19665 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17572), .ZN(
        n16633) );
  NAND2_X1 U19666 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16633), .ZN(
        n16622) );
  NOR2_X1 U19667 ( .A1(n16501), .A2(n16622), .ZN(n16568) );
  NAND2_X1 U19668 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n16568), .ZN(
        n17472) );
  NOR2_X1 U19669 ( .A1(n17487), .A2(n17472), .ZN(n16531) );
  NAND2_X1 U19670 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16531), .ZN(
        n16519) );
  NOR2_X1 U19671 ( .A1(n17448), .A2(n16519), .ZN(n16502) );
  OAI22_X1 U19672 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16502), .B1(
        n17639), .B2(n17422), .ZN(n17440) );
  INV_X1 U19673 ( .A(n17440), .ZN(n16505) );
  NAND2_X1 U19674 ( .A1(n16503), .A2(n9732), .ZN(n16511) );
  INV_X1 U19675 ( .A(n16511), .ZN(n16504) );
  OAI221_X1 U19676 ( .B1(n16505), .B2(n16504), .C1(n17440), .C2(n16511), .A(
        n18487), .ZN(n16506) );
  OAI211_X1 U19677 ( .C1(n16508), .C2(n18542), .A(n16507), .B(n16506), .ZN(
        P3_U2655) );
  AOI221_X1 U19678 ( .B1(n16691), .B2(n18540), .C1(n16522), .C2(n18540), .A(
        n16508), .ZN(n16516) );
  INV_X1 U19679 ( .A(n16519), .ZN(n17435) );
  AOI22_X1 U19680 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n16519), .B1(
        n17435), .B2(n17448), .ZN(n17445) );
  INV_X1 U19681 ( .A(n16686), .ZN(n16675) );
  OAI21_X1 U19682 ( .B1(n16509), .B2(n17445), .A(n18487), .ZN(n16510) );
  AOI22_X1 U19683 ( .A1(n17445), .A2(n16511), .B1(n16675), .B2(n16510), .ZN(
        n16515) );
  OAI211_X1 U19684 ( .C1(n16520), .C2(n16518), .A(n16696), .B(n16512), .ZN(
        n16513) );
  OAI21_X1 U19685 ( .B1(n20832), .B2(n17448), .A(n16513), .ZN(n16514) );
  NOR3_X1 U19686 ( .A1(n16516), .A2(n16515), .A3(n16514), .ZN(n16517) );
  OAI211_X1 U19687 ( .C1(n16700), .C2(n16518), .A(n16517), .B(n17963), .ZN(
        P3_U2656) );
  INV_X1 U19688 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16606) );
  AOI21_X1 U19689 ( .B1(n16531), .B2(n16606), .A(n16659), .ZN(n16535) );
  OAI21_X1 U19690 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16531), .A(
        n16519), .ZN(n17465) );
  XOR2_X1 U19691 ( .A(n16535), .B(n17465), .Z(n16529) );
  AOI21_X1 U19692 ( .B1(n20834), .B2(P3_EBX_REG_14__SCAN_IN), .A(n17965), .ZN(
        n16528) );
  AOI211_X1 U19693 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16536), .A(n16520), .B(
        n20820), .ZN(n16526) );
  NAND2_X1 U19694 ( .A1(n20827), .A2(n16521), .ZN(n16530) );
  NAND2_X1 U19695 ( .A1(n16703), .A2(n16691), .ZN(n16701) );
  NAND2_X1 U19696 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16701), .ZN(n16524) );
  INV_X1 U19697 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18535) );
  NOR2_X1 U19698 ( .A1(n20825), .A2(n16522), .ZN(n16523) );
  AOI221_X1 U19699 ( .B1(n16530), .B2(n16524), .C1(n18535), .C2(n16524), .A(
        n16523), .ZN(n16525) );
  AOI211_X1 U19700 ( .C1(n16688), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16526), .B(n16525), .ZN(n16527) );
  OAI211_X1 U19701 ( .C1(n20816), .C2(n16529), .A(n16528), .B(n16527), .ZN(
        P3_U2657) );
  AOI21_X1 U19702 ( .B1(n20827), .B2(n16549), .A(n20825), .ZN(n16559) );
  NAND2_X1 U19703 ( .A1(n20827), .A2(n18534), .ZN(n16548) );
  AOI21_X1 U19704 ( .B1(n16559), .B2(n16548), .A(n18535), .ZN(n16542) );
  INV_X1 U19705 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16532) );
  OAI22_X1 U19706 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16530), .B1(n16532), 
        .B2(n20832), .ZN(n16541) );
  INV_X1 U19707 ( .A(n17472), .ZN(n16546) );
  NAND2_X1 U19708 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16546), .ZN(
        n16545) );
  AOI21_X1 U19709 ( .B1(n16532), .B2(n16545), .A(n16531), .ZN(n17475) );
  OAI211_X1 U19710 ( .C1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n16545), .A(
        n9732), .B(n17475), .ZN(n16534) );
  OAI211_X1 U19711 ( .C1(n17475), .C2(n16535), .A(n18487), .B(n16534), .ZN(
        n16538) );
  OAI211_X1 U19712 ( .C1(n16543), .C2(n16539), .A(n16696), .B(n16536), .ZN(
        n16537) );
  OAI211_X1 U19713 ( .C1(n16539), .C2(n16700), .A(n16538), .B(n16537), .ZN(
        n16540) );
  OR4_X1 U19714 ( .A1(n17965), .A2(n16542), .A3(n16541), .A4(n16540), .ZN(
        P3_U2658) );
  AOI211_X1 U19715 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16562), .A(n16543), .B(
        n20820), .ZN(n16544) );
  AOI21_X1 U19716 ( .B1(n16688), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16544), .ZN(n16554) );
  AOI21_X1 U19717 ( .B1(n16546), .B2(n16606), .A(n16659), .ZN(n16547) );
  OAI21_X1 U19718 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n16546), .A(
        n16545), .ZN(n17503) );
  XNOR2_X1 U19719 ( .A(n16547), .B(n17503), .ZN(n16552) );
  OAI22_X1 U19720 ( .A1(n16700), .A2(n16550), .B1(n16549), .B2(n16548), .ZN(
        n16551) );
  AOI211_X1 U19721 ( .C1(n18487), .C2(n16552), .A(n17965), .B(n16551), .ZN(
        n16553) );
  OAI211_X1 U19722 ( .C1(n18534), .C2(n16559), .A(n16554), .B(n16553), .ZN(
        P3_U2659) );
  INV_X1 U19723 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17508) );
  INV_X1 U19724 ( .A(n16555), .ZN(n16567) );
  NAND2_X1 U19725 ( .A1(n20827), .A2(n16566), .ZN(n16617) );
  NOR2_X1 U19726 ( .A1(n16567), .A2(n16617), .ZN(n16582) );
  AOI21_X1 U19727 ( .B1(n16556), .B2(n16582), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16560) );
  INV_X1 U19728 ( .A(n16622), .ZN(n16608) );
  NAND4_X1 U19729 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A4(n16608), .ZN(n16580) );
  NOR2_X1 U19730 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16580), .ZN(
        n16591) );
  AOI21_X1 U19731 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16591), .A(
        n16659), .ZN(n16557) );
  OAI21_X1 U19732 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16568), .A(
        n17472), .ZN(n17510) );
  XOR2_X1 U19733 ( .A(n16557), .B(n17510), .Z(n16558) );
  OAI22_X1 U19734 ( .A1(n16560), .A2(n16559), .B1(n20816), .B2(n16558), .ZN(
        n16561) );
  AOI211_X1 U19735 ( .C1(n20834), .C2(P3_EBX_REG_11__SCAN_IN), .A(n11114), .B(
        n16561), .ZN(n16565) );
  OAI211_X1 U19736 ( .C1(n16571), .C2(n16563), .A(n16696), .B(n16562), .ZN(
        n16564) );
  OAI211_X1 U19737 ( .C1(n20832), .C2(n17508), .A(n16565), .B(n16564), .ZN(
        P3_U2660) );
  NAND2_X1 U19738 ( .A1(n16566), .A2(n16703), .ZN(n16618) );
  OAI21_X1 U19739 ( .B1(n16567), .B2(n16618), .A(n16701), .ZN(n16604) );
  INV_X1 U19740 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18530) );
  INV_X1 U19741 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16573) );
  AOI21_X1 U19742 ( .B1(n16573), .B2(n16580), .A(n16568), .ZN(n17517) );
  NOR2_X1 U19743 ( .A1(n16591), .A2(n16659), .ZN(n16570) );
  OAI21_X1 U19744 ( .B1(n17517), .B2(n16570), .A(n18487), .ZN(n16569) );
  AOI21_X1 U19745 ( .B1(n17517), .B2(n16570), .A(n16569), .ZN(n16576) );
  AOI211_X1 U19746 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16572), .A(n16571), .B(
        n20820), .ZN(n16575) );
  OAI22_X1 U19747 ( .A1(n16573), .A2(n20832), .B1(n16700), .B2(n16921), .ZN(
        n16574) );
  NOR4_X1 U19748 ( .A1(n17965), .A2(n16576), .A3(n16575), .A4(n16574), .ZN(
        n16579) );
  OAI211_X1 U19749 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(P3_REIP_REG_10__SCAN_IN), 
        .A(n16582), .B(n16577), .ZN(n16578) );
  OAI211_X1 U19750 ( .C1(n16604), .C2(n18530), .A(n16579), .B(n16578), .ZN(
        P3_U2661) );
  INV_X1 U19751 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17543) );
  INV_X1 U19752 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20849) );
  NOR2_X1 U19753 ( .A1(n20849), .A2(n16622), .ZN(n16594) );
  INV_X1 U19754 ( .A(n16594), .ZN(n16607) );
  NOR2_X1 U19755 ( .A1(n17543), .A2(n16607), .ZN(n16595) );
  OAI21_X1 U19756 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16595), .A(
        n16580), .ZN(n17534) );
  NOR2_X1 U19757 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20816), .ZN(
        n16687) );
  AOI22_X1 U19758 ( .A1(n16689), .A2(n17534), .B1(n16595), .B2(n16687), .ZN(
        n16590) );
  AOI21_X1 U19759 ( .B1(n16696), .B2(n16584), .A(n20834), .ZN(n16581) );
  INV_X1 U19760 ( .A(n16581), .ZN(n16583) );
  INV_X1 U19761 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18528) );
  AOI22_X1 U19762 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n16583), .B1(n16582), .B2(
        n18528), .ZN(n16589) );
  NOR2_X1 U19763 ( .A1(n16584), .A2(n20820), .ZN(n16593) );
  OAI22_X1 U19764 ( .A1(n18528), .A2(n16604), .B1(n17534), .B2(n16675), .ZN(
        n16586) );
  INV_X1 U19765 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17532) );
  OAI21_X1 U19766 ( .B1(n17532), .B2(n20832), .A(n17963), .ZN(n16585) );
  AOI211_X1 U19767 ( .C1(n16593), .C2(n16587), .A(n16586), .B(n16585), .ZN(
        n16588) );
  OAI211_X1 U19768 ( .C1(n16591), .C2(n16590), .A(n16589), .B(n16588), .ZN(
        P3_U2662) );
  NAND2_X1 U19769 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16609), .ZN(n16592) );
  AOI22_X1 U19770 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n20834), .B1(n16593), .B2(
        n16592), .ZN(n16603) );
  AOI21_X1 U19771 ( .B1(n16594), .B2(n16606), .A(n16659), .ZN(n16597) );
  AOI21_X1 U19772 ( .B1(n17543), .B2(n16607), .A(n16595), .ZN(n16596) );
  INV_X1 U19773 ( .A(n16596), .ZN(n17555) );
  XNOR2_X1 U19774 ( .A(n16597), .B(n17555), .ZN(n16601) );
  NOR3_X1 U19775 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16598), .A3(n16617), .ZN(
        n16600) );
  OAI21_X1 U19776 ( .B1(n17543), .B2(n20832), .A(n17963), .ZN(n16599) );
  AOI211_X1 U19777 ( .C1(n16601), .C2(n18487), .A(n16600), .B(n16599), .ZN(
        n16602) );
  OAI211_X1 U19778 ( .C1(n18526), .C2(n16604), .A(n16603), .B(n16602), .ZN(
        P3_U2663) );
  AOI21_X1 U19779 ( .B1(n16608), .B2(n16606), .A(n16605), .ZN(n16629) );
  OAI21_X1 U19780 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16608), .A(
        n16607), .ZN(n16615) );
  INV_X1 U19781 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18521) );
  NOR3_X1 U19782 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n18521), .A3(n16617), .ZN(
        n16614) );
  AOI22_X1 U19783 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16688), .B1(
        n20834), .B2(P3_EBX_REG_7__SCAN_IN), .ZN(n16612) );
  OAI211_X1 U19784 ( .C1(n16624), .C2(n16610), .A(n16696), .B(n16609), .ZN(
        n16611) );
  NAND3_X1 U19785 ( .A1(n16612), .A2(n17963), .A3(n16611), .ZN(n16613) );
  AOI211_X1 U19786 ( .C1(n16629), .C2(n16615), .A(n16614), .B(n16613), .ZN(
        n16621) );
  NOR2_X1 U19787 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16622), .ZN(
        n16616) );
  INV_X1 U19788 ( .A(n16615), .ZN(n17566) );
  OAI211_X1 U19789 ( .C1(n16616), .C2(n16659), .A(n18487), .B(n17566), .ZN(
        n16620) );
  NOR2_X1 U19790 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16617), .ZN(n16623) );
  NAND2_X1 U19791 ( .A1(n16701), .A2(n16618), .ZN(n16635) );
  INV_X1 U19792 ( .A(n16635), .ZN(n16625) );
  OAI21_X1 U19793 ( .B1(n16623), .B2(n16625), .A(P3_REIP_REG_7__SCAN_IN), .ZN(
        n16619) );
  NAND3_X1 U19794 ( .A1(n16621), .A2(n16620), .A3(n16619), .ZN(P3_U2664) );
  OAI21_X1 U19795 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16633), .A(
        n16622), .ZN(n17575) );
  AOI21_X1 U19796 ( .B1(n16633), .B2(n16687), .A(n16686), .ZN(n16632) );
  AOI211_X1 U19797 ( .C1(n20834), .C2(P3_EBX_REG_6__SCAN_IN), .A(n11114), .B(
        n16623), .ZN(n16631) );
  AOI211_X1 U19798 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16638), .A(n16624), .B(
        n20820), .ZN(n16628) );
  AOI22_X1 U19799 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16688), .B1(
        P3_REIP_REG_6__SCAN_IN), .B2(n16625), .ZN(n16626) );
  INV_X1 U19800 ( .A(n16626), .ZN(n16627) );
  AOI211_X1 U19801 ( .C1(n16629), .C2(n17575), .A(n16628), .B(n16627), .ZN(
        n16630) );
  OAI211_X1 U19802 ( .C1(n17575), .C2(n16632), .A(n16631), .B(n16630), .ZN(
        P3_U2665) );
  NOR2_X1 U19803 ( .A1(n16691), .A2(n16650), .ZN(n16654) );
  AOI21_X1 U19804 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n16654), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n16636) );
  NAND2_X1 U19805 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9898), .ZN(
        n16643) );
  AOI21_X1 U19806 ( .B1(n17587), .B2(n16643), .A(n16633), .ZN(n17589) );
  AOI21_X1 U19807 ( .B1(n9898), .B2(n16674), .A(n16659), .ZN(n16644) );
  XNOR2_X1 U19808 ( .A(n17589), .B(n16644), .ZN(n16634) );
  OAI22_X1 U19809 ( .A1(n16636), .A2(n16635), .B1(n20816), .B2(n16634), .ZN(
        n16637) );
  AOI211_X1 U19810 ( .C1(n20834), .C2(P3_EBX_REG_5__SCAN_IN), .A(n11114), .B(
        n16637), .ZN(n16641) );
  OAI211_X1 U19811 ( .C1(n16645), .C2(n16639), .A(n16696), .B(n16638), .ZN(
        n16640) );
  OAI211_X1 U19812 ( .C1(n20832), .C2(n17587), .A(n16641), .B(n16640), .ZN(
        P3_U2666) );
  NOR2_X1 U19813 ( .A1(n16642), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17597) );
  NOR2_X1 U19814 ( .A1(n17639), .A2(n16642), .ZN(n16658) );
  OAI21_X1 U19815 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16658), .A(
        n16643), .ZN(n17607) );
  AOI22_X1 U19816 ( .A1(n16674), .A2(n17597), .B1(n16644), .B2(n17607), .ZN(
        n16657) );
  INV_X1 U19817 ( .A(n17607), .ZN(n16649) );
  AOI211_X1 U19818 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16667), .A(n16645), .B(
        n20820), .ZN(n16648) );
  NAND2_X1 U19819 ( .A1(n16646), .A2(n18651), .ZN(n16706) );
  OAI221_X1 U19820 ( .B1(n16706), .B2(n9694), .C1(n16706), .C2(n18478), .A(
        n17963), .ZN(n16647) );
  AOI211_X1 U19821 ( .C1(n16686), .C2(n16649), .A(n16648), .B(n16647), .ZN(
        n16656) );
  AOI21_X1 U19822 ( .B1(n16650), .B2(n20827), .A(n20825), .ZN(n16651) );
  INV_X1 U19823 ( .A(n16651), .ZN(n16666) );
  AOI22_X1 U19824 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16688), .B1(
        n20834), .B2(P3_EBX_REG_4__SCAN_IN), .ZN(n16652) );
  INV_X1 U19825 ( .A(n16652), .ZN(n16653) );
  AOI221_X1 U19826 ( .B1(n16666), .B2(P3_REIP_REG_4__SCAN_IN), .C1(n16654), 
        .C2(n18518), .A(n16653), .ZN(n16655) );
  OAI211_X1 U19827 ( .C1(n16657), .C2(n20816), .A(n16656), .B(n16655), .ZN(
        P3_U2667) );
  INV_X1 U19828 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17613) );
  NAND2_X1 U19829 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16681) );
  INV_X1 U19830 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18516) );
  OAI21_X1 U19831 ( .B1(n16681), .B2(n16691), .A(n18516), .ZN(n16665) );
  NAND2_X1 U19832 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16673) );
  AOI21_X1 U19833 ( .B1(n17613), .B2(n16673), .A(n16658), .ZN(n17617) );
  NOR2_X1 U19834 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16673), .ZN(
        n16677) );
  NOR2_X1 U19835 ( .A1(n16677), .A2(n16659), .ZN(n16661) );
  OAI21_X1 U19836 ( .B1(n17617), .B2(n16661), .A(n18487), .ZN(n16660) );
  AOI21_X1 U19837 ( .B1(n17617), .B2(n16661), .A(n16660), .ZN(n16664) );
  NOR2_X1 U19838 ( .A1(n11052), .A2(n18604), .ZN(n18440) );
  NAND2_X1 U19839 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18440), .ZN(
        n16672) );
  AOI21_X1 U19840 ( .B1(n18590), .B2(n16672), .A(n16945), .ZN(n18587) );
  INV_X1 U19841 ( .A(n18587), .ZN(n16662) );
  OAI22_X1 U19842 ( .A1(n16700), .A2(n16668), .B1(n16706), .B2(n16662), .ZN(
        n16663) );
  AOI211_X1 U19843 ( .C1(n16666), .C2(n16665), .A(n16664), .B(n16663), .ZN(
        n16670) );
  OAI211_X1 U19844 ( .C1(n16685), .C2(n16668), .A(n16696), .B(n16667), .ZN(
        n16669) );
  OAI211_X1 U19845 ( .C1(n20832), .C2(n17613), .A(n16670), .B(n16669), .ZN(
        P3_U2668) );
  NOR2_X1 U19846 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n16690) );
  OAI21_X1 U19847 ( .B1(n16690), .B2(n16671), .A(n16696), .ZN(n16684) );
  INV_X1 U19848 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17631) );
  OAI22_X1 U19849 ( .A1(n17631), .A2(n20832), .B1(n16700), .B2(n16671), .ZN(
        n16680) );
  INV_X1 U19850 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18514) );
  NAND2_X1 U19851 ( .A1(n11052), .A2(n16693), .ZN(n18442) );
  NAND2_X1 U19852 ( .A1(n18442), .A2(n16672), .ZN(n18592) );
  OAI22_X1 U19853 ( .A1(n16703), .A2(n18514), .B1(n18592), .B2(n16706), .ZN(
        n16679) );
  OAI21_X1 U19854 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16673), .ZN(n17626) );
  OAI21_X1 U19855 ( .B1(n16674), .B2(n17626), .A(n16689), .ZN(n16676) );
  OAI22_X1 U19856 ( .A1(n16677), .A2(n16676), .B1(n17626), .B2(n16675), .ZN(
        n16678) );
  NOR3_X1 U19857 ( .A1(n16680), .A2(n16679), .A3(n16678), .ZN(n16683) );
  OAI211_X1 U19858 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n20827), .B(n16681), .ZN(n16682) );
  OAI211_X1 U19859 ( .C1(n16685), .C2(n16684), .A(n16683), .B(n16682), .ZN(
        P3_U2669) );
  NOR2_X1 U19860 ( .A1(n16687), .A2(n16686), .ZN(n16699) );
  AOI21_X1 U19861 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16689), .A(
        n16688), .ZN(n16698) );
  AOI21_X1 U19862 ( .B1(P3_EBX_REG_1__SCAN_IN), .B2(P3_EBX_REG_0__SCAN_IN), 
        .A(n16690), .ZN(n16992) );
  INV_X1 U19863 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n16995) );
  OAI22_X1 U19864 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16691), .B1(n16700), 
        .B2(n16995), .ZN(n16695) );
  NAND2_X1 U19865 ( .A1(n16693), .A2(n16692), .ZN(n18598) );
  OAI22_X1 U19866 ( .A1(n16703), .A2(n18614), .B1(n18598), .B2(n16706), .ZN(
        n16694) );
  AOI211_X1 U19867 ( .C1(n16696), .C2(n16992), .A(n16695), .B(n16694), .ZN(
        n16697) );
  OAI221_X1 U19868 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16699), .C1(
        n17639), .C2(n16698), .A(n16697), .ZN(P3_U2670) );
  NAND2_X1 U19869 ( .A1(n16700), .A2(n20820), .ZN(n16702) );
  AOI22_X1 U19870 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n16702), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n16701), .ZN(n16705) );
  NAND3_X1 U19871 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18593), .A3(
        n16703), .ZN(n16704) );
  OAI211_X1 U19872 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n16706), .A(
        n16705), .B(n16704), .ZN(P3_U2671) );
  INV_X1 U19873 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16784) );
  NOR3_X1 U19874 ( .A1(n16784), .A2(n16783), .A3(n16707), .ZN(n16708) );
  NAND4_X1 U19875 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_26__SCAN_IN), 
        .A3(n16742), .A4(n16708), .ZN(n16711) );
  NOR2_X1 U19876 ( .A1(n16712), .A2(n16711), .ZN(n16737) );
  NAND2_X1 U19877 ( .A1(n16980), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16710) );
  NAND2_X1 U19878 ( .A1(n16737), .A2(n18024), .ZN(n16709) );
  OAI22_X1 U19879 ( .A1(n16737), .A2(n16710), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16709), .ZN(P3_U2672) );
  NAND2_X1 U19880 ( .A1(n16712), .A2(n16711), .ZN(n16713) );
  NAND2_X1 U19881 ( .A1(n16713), .A2(n16980), .ZN(n16736) );
  AOI22_X1 U19882 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16844), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16723) );
  AOI22_X1 U19883 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n15523), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16722) );
  AOI22_X1 U19884 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n16955), .ZN(n16714) );
  OAI21_X1 U19885 ( .B1(n20770), .B2(n9694), .A(n16714), .ZN(n16720) );
  AOI22_X1 U19886 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n15525), .B1(
        n16952), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16718) );
  AOI22_X1 U19887 ( .A1(n16946), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n16944), .ZN(n16717) );
  AOI22_X1 U19888 ( .A1(n16927), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n9588), .ZN(n16716) );
  AOI22_X1 U19889 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n16883), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16715) );
  NAND4_X1 U19890 ( .A1(n16718), .A2(n16717), .A3(n16716), .A4(n16715), .ZN(
        n16719) );
  AOI211_X1 U19891 ( .C1(n16962), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n16720), .B(n16719), .ZN(n16721) );
  NAND3_X1 U19892 ( .A1(n16723), .A2(n16722), .A3(n16721), .ZN(n16735) );
  AOI22_X1 U19893 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16727) );
  AOI22_X1 U19894 ( .A1(n16946), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16726) );
  AOI22_X1 U19895 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16725) );
  AOI22_X1 U19896 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16724) );
  NAND4_X1 U19897 ( .A1(n16727), .A2(n16726), .A3(n16725), .A4(n16724), .ZN(
        n16733) );
  AOI22_X1 U19898 ( .A1(n16883), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16731) );
  AOI22_X1 U19899 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16730) );
  AOI22_X1 U19900 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16729) );
  AOI22_X1 U19901 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16728) );
  NAND4_X1 U19902 ( .A1(n16731), .A2(n16730), .A3(n16729), .A4(n16728), .ZN(
        n16732) );
  NOR2_X1 U19903 ( .A1(n16733), .A2(n16732), .ZN(n16740) );
  NOR3_X1 U19904 ( .A1(n16740), .A2(n16738), .A3(n17021), .ZN(n16734) );
  XNOR2_X1 U19905 ( .A(n16735), .B(n16734), .ZN(n17008) );
  OAI22_X1 U19906 ( .A1(n16737), .A2(n16736), .B1(n17008), .B2(n16980), .ZN(
        P3_U2673) );
  NOR2_X1 U19907 ( .A1(n16738), .A2(n17021), .ZN(n16739) );
  XOR2_X1 U19908 ( .A(n16740), .B(n16739), .Z(n17015) );
  NOR2_X1 U19909 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16748), .ZN(n16741) );
  AOI22_X1 U19910 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16743), .B1(n16742), 
        .B2(n16741), .ZN(n16744) );
  OAI21_X1 U19911 ( .B1(n16980), .B2(n17015), .A(n16744), .ZN(P3_U2674) );
  OAI211_X1 U19912 ( .C1(n17023), .C2(n17022), .A(n16998), .B(n17021), .ZN(
        n16745) );
  OAI221_X1 U19913 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n16748), .C1(n16747), 
        .C2(n16746), .A(n16745), .ZN(P3_U2676) );
  INV_X1 U19914 ( .A(n16748), .ZN(n16753) );
  AOI21_X1 U19915 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n16980), .A(n16758), .ZN(
        n16752) );
  OAI21_X1 U19916 ( .B1(n16760), .B2(n16756), .A(n16749), .ZN(n16751) );
  INV_X1 U19917 ( .A(n17023), .ZN(n16750) );
  NAND2_X1 U19918 ( .A1(n16751), .A2(n16750), .ZN(n17032) );
  OAI22_X1 U19919 ( .A1(n16753), .A2(n16752), .B1(n16980), .B2(n17032), .ZN(
        P3_U2677) );
  INV_X1 U19920 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n20795) );
  INV_X1 U19921 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16755) );
  INV_X1 U19922 ( .A(n16754), .ZN(n16795) );
  NAND2_X1 U19923 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16795), .ZN(n16782) );
  NOR2_X1 U19924 ( .A1(n16755), .A2(n16782), .ZN(n16765) );
  NAND2_X1 U19925 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n16765), .ZN(n16759) );
  NOR2_X1 U19926 ( .A1(n20795), .A2(n16759), .ZN(n16764) );
  AOI21_X1 U19927 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n16980), .A(n16764), .ZN(
        n16757) );
  XNOR2_X1 U19928 ( .A(n16760), .B(n16756), .ZN(n17037) );
  OAI22_X1 U19929 ( .A1(n16758), .A2(n16757), .B1(n17037), .B2(n16980), .ZN(
        P3_U2678) );
  INV_X1 U19930 ( .A(n16759), .ZN(n16770) );
  AOI21_X1 U19931 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16980), .A(n16770), .ZN(
        n16763) );
  OAI21_X1 U19932 ( .B1(n16762), .B2(n16761), .A(n16760), .ZN(n17042) );
  OAI22_X1 U19933 ( .A1(n16764), .A2(n16763), .B1(n16980), .B2(n17042), .ZN(
        P3_U2679) );
  AOI21_X1 U19934 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n16980), .A(n16765), .ZN(
        n16769) );
  OAI21_X1 U19935 ( .B1(n16768), .B2(n16767), .A(n16766), .ZN(n17047) );
  OAI22_X1 U19936 ( .A1(n16770), .A2(n16769), .B1(n16980), .B2(n17047), .ZN(
        P3_U2680) );
  AOI22_X1 U19937 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16883), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16774) );
  AOI22_X1 U19938 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16773) );
  AOI22_X1 U19939 ( .A1(n16946), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16772) );
  AOI22_X1 U19940 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16771) );
  NAND4_X1 U19941 ( .A1(n16774), .A2(n16773), .A3(n16772), .A4(n16771), .ZN(
        n16780) );
  AOI22_X1 U19942 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16778) );
  AOI22_X1 U19943 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16777) );
  AOI22_X1 U19944 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16776) );
  AOI22_X1 U19945 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n16844), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16775) );
  NAND4_X1 U19946 ( .A1(n16778), .A2(n16777), .A3(n16776), .A4(n16775), .ZN(
        n16779) );
  NOR2_X1 U19947 ( .A1(n16780), .A2(n16779), .ZN(n17051) );
  NAND3_X1 U19948 ( .A1(n16782), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n16980), 
        .ZN(n16781) );
  OAI221_X1 U19949 ( .B1(n16782), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n16980), 
        .C2(n17051), .A(n16781), .ZN(P3_U2681) );
  OAI21_X1 U19950 ( .B1(n16784), .B2(n16783), .A(n16980), .ZN(n16809) );
  AOI22_X1 U19951 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16794) );
  AOI22_X1 U19952 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16793) );
  AOI22_X1 U19953 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16785) );
  OAI21_X1 U19954 ( .B1(n10090), .B2(n20847), .A(n16785), .ZN(n16791) );
  AOI22_X1 U19955 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16883), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16789) );
  AOI22_X1 U19956 ( .A1(n16955), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16788) );
  AOI22_X1 U19957 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16787) );
  AOI22_X1 U19958 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16786) );
  NAND4_X1 U19959 ( .A1(n16789), .A2(n16788), .A3(n16787), .A4(n16786), .ZN(
        n16790) );
  AOI211_X1 U19960 ( .C1(n16946), .C2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n16791), .B(n16790), .ZN(n16792) );
  NAND3_X1 U19961 ( .A1(n16794), .A2(n16793), .A3(n16792), .ZN(n17056) );
  AOI22_X1 U19962 ( .A1(n16998), .A2(n17056), .B1(n16795), .B2(n16797), .ZN(
        n16796) );
  OAI21_X1 U19963 ( .B1(n16797), .B2(n16809), .A(n16796), .ZN(P3_U2682) );
  AOI22_X1 U19964 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16883), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16801) );
  AOI22_X1 U19965 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16872), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16800) );
  AOI22_X1 U19966 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16799) );
  AOI22_X1 U19967 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16798) );
  NAND4_X1 U19968 ( .A1(n16801), .A2(n16800), .A3(n16799), .A4(n16798), .ZN(
        n16807) );
  AOI22_X1 U19969 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16805) );
  AOI22_X1 U19970 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16804) );
  AOI22_X1 U19971 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16803) );
  AOI22_X1 U19972 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16802) );
  NAND4_X1 U19973 ( .A1(n16805), .A2(n16804), .A3(n16803), .A4(n16802), .ZN(
        n16806) );
  NOR2_X1 U19974 ( .A1(n16807), .A2(n16806), .ZN(n17065) );
  NOR2_X1 U19975 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16808), .ZN(n16810) );
  OAI22_X1 U19976 ( .A1(n17065), .A2(n16980), .B1(n16810), .B2(n16809), .ZN(
        P3_U2683) );
  AOI22_X1 U19977 ( .A1(n16927), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16814) );
  AOI22_X1 U19978 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n16883), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16813) );
  AOI22_X1 U19979 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16952), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16812) );
  AOI22_X1 U19980 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16811) );
  NAND4_X1 U19981 ( .A1(n16814), .A2(n16813), .A3(n16812), .A4(n16811), .ZN(
        n16820) );
  AOI22_X1 U19982 ( .A1(n15523), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16818) );
  AOI22_X1 U19983 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16844), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16817) );
  AOI22_X1 U19984 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16816) );
  AOI22_X1 U19985 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16815) );
  NAND4_X1 U19986 ( .A1(n16818), .A2(n16817), .A3(n16816), .A4(n16815), .ZN(
        n16819) );
  NOR2_X1 U19987 ( .A1(n16820), .A2(n16819), .ZN(n17069) );
  INV_X1 U19988 ( .A(n16821), .ZN(n16823) );
  OAI33_X1 U19989 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17092), .A3(n16823), 
        .B1(n16822), .B2(n16998), .B3(n16821), .ZN(n16824) );
  INV_X1 U19990 ( .A(n16824), .ZN(n16825) );
  OAI21_X1 U19991 ( .B1(n17069), .B2(n16980), .A(n16825), .ZN(P3_U2684) );
  AOI22_X1 U19992 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16829) );
  AOI22_X1 U19993 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16828) );
  AOI22_X1 U19994 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16827) );
  AOI22_X1 U19995 ( .A1(n16883), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16826) );
  NAND4_X1 U19996 ( .A1(n16829), .A2(n16828), .A3(n16827), .A4(n16826), .ZN(
        n16835) );
  AOI22_X1 U19997 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16952), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16833) );
  AOI22_X1 U19998 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n16832) );
  AOI22_X1 U19999 ( .A1(n16927), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16831) );
  AOI22_X1 U20000 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16830) );
  NAND4_X1 U20001 ( .A1(n16833), .A2(n16832), .A3(n16831), .A4(n16830), .ZN(
        n16834) );
  NOR2_X1 U20002 ( .A1(n16835), .A2(n16834), .ZN(n17070) );
  NAND4_X1 U20003 ( .A1(n18024), .A2(P3_EBX_REG_17__SCAN_IN), .A3(n16867), 
        .A4(n16836), .ZN(n16838) );
  NAND3_X1 U20004 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16980), .A3(n16851), 
        .ZN(n16837) );
  OAI211_X1 U20005 ( .C1(n17070), .C2(n16980), .A(n16838), .B(n16837), .ZN(
        P3_U2685) );
  AOI22_X1 U20006 ( .A1(n16839), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16843) );
  AOI22_X1 U20007 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n16883), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16842) );
  AOI22_X1 U20008 ( .A1(n15523), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16841) );
  AOI22_X1 U20009 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n16840) );
  NAND4_X1 U20010 ( .A1(n16843), .A2(n16842), .A3(n16841), .A4(n16840), .ZN(
        n16850) );
  AOI22_X1 U20011 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16848) );
  AOI22_X1 U20012 ( .A1(n16927), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n16844), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n16847) );
  AOI22_X1 U20013 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16846) );
  AOI22_X1 U20014 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16845) );
  NAND4_X1 U20015 ( .A1(n16848), .A2(n16847), .A3(n16846), .A4(n16845), .ZN(
        n16849) );
  NOR2_X1 U20016 ( .A1(n16850), .A2(n16849), .ZN(n17080) );
  NOR2_X1 U20017 ( .A1(n16867), .A2(P3_EBX_REG_17__SCAN_IN), .ZN(n16853) );
  NAND2_X1 U20018 ( .A1(n16980), .A2(n16851), .ZN(n16852) );
  OAI22_X1 U20019 ( .A1(n17080), .A2(n16980), .B1(n16853), .B2(n16852), .ZN(
        P3_U2686) );
  AOI21_X1 U20020 ( .B1(n16854), .B2(n16879), .A(n16998), .ZN(n16855) );
  INV_X1 U20021 ( .A(n16855), .ZN(n16866) );
  AOI22_X1 U20022 ( .A1(n15523), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16859) );
  AOI22_X1 U20023 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16858) );
  AOI22_X1 U20024 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16857) );
  AOI22_X1 U20025 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16856) );
  NAND4_X1 U20026 ( .A1(n16859), .A2(n16858), .A3(n16857), .A4(n16856), .ZN(
        n16865) );
  AOI22_X1 U20027 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16883), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16863) );
  AOI22_X1 U20028 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16862) );
  AOI22_X1 U20029 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16861) );
  AOI22_X1 U20030 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16860) );
  NAND4_X1 U20031 ( .A1(n16863), .A2(n16862), .A3(n16861), .A4(n16860), .ZN(
        n16864) );
  NOR2_X1 U20032 ( .A1(n16865), .A2(n16864), .ZN(n17086) );
  OAI22_X1 U20033 ( .A1(n16867), .A2(n16866), .B1(n17086), .B2(n16980), .ZN(
        P3_U2687) );
  AOI22_X1 U20034 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n16883), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16871) );
  AOI22_X1 U20035 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n16910), .ZN(n16870) );
  AOI22_X1 U20036 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n15523), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n16944), .ZN(n16869) );
  AOI22_X1 U20037 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n9588), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n16928), .ZN(n16868) );
  NAND4_X1 U20038 ( .A1(n16871), .A2(n16870), .A3(n16869), .A4(n16868), .ZN(
        n16878) );
  AOI22_X1 U20039 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n16872), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16876) );
  AOI22_X1 U20040 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16875) );
  AOI22_X1 U20041 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n15525), .ZN(n16874) );
  AOI22_X1 U20042 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n16955), .ZN(n16873) );
  NAND4_X1 U20043 ( .A1(n16876), .A2(n16875), .A3(n16874), .A4(n16873), .ZN(
        n16877) );
  NOR2_X1 U20044 ( .A1(n16878), .A2(n16877), .ZN(n17091) );
  OAI21_X1 U20045 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n16880), .A(n16879), .ZN(
        n16881) );
  AOI22_X1 U20046 ( .A1(n16998), .A2(n17091), .B1(n16881), .B2(n16980), .ZN(
        P3_U2688) );
  INV_X1 U20047 ( .A(n16882), .ZN(n16907) );
  AOI21_X1 U20048 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n16980), .A(n16907), .ZN(
        n16894) );
  AOI22_X1 U20049 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16883), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16887) );
  AOI22_X1 U20050 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16886) );
  AOI22_X1 U20051 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16926), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16885) );
  AOI22_X1 U20052 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16884) );
  NAND4_X1 U20053 ( .A1(n16887), .A2(n16886), .A3(n16885), .A4(n16884), .ZN(
        n16893) );
  AOI22_X1 U20054 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16891) );
  AOI22_X1 U20055 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16890) );
  AOI22_X1 U20056 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16889) );
  AOI22_X1 U20057 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16888) );
  NAND4_X1 U20058 ( .A1(n16891), .A2(n16890), .A3(n16889), .A4(n16888), .ZN(
        n16892) );
  NOR2_X1 U20059 ( .A1(n16893), .A2(n16892), .ZN(n17104) );
  OAI22_X1 U20060 ( .A1(n16895), .A2(n16894), .B1(n17104), .B2(n16980), .ZN(
        P3_U2691) );
  AOI22_X1 U20061 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16899) );
  AOI22_X1 U20062 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16898) );
  AOI22_X1 U20063 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16897) );
  AOI22_X1 U20064 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16896) );
  NAND4_X1 U20065 ( .A1(n16899), .A2(n16898), .A3(n16897), .A4(n16896), .ZN(
        n16905) );
  AOI22_X1 U20066 ( .A1(n10858), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16903) );
  AOI22_X1 U20067 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16902) );
  AOI22_X1 U20068 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16901) );
  AOI22_X1 U20069 ( .A1(n15523), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16900) );
  NAND4_X1 U20070 ( .A1(n16903), .A2(n16902), .A3(n16901), .A4(n16900), .ZN(
        n16904) );
  NOR2_X1 U20071 ( .A1(n16905), .A2(n16904), .ZN(n17108) );
  AOI211_X1 U20072 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16922), .A(
        P3_EBX_REG_11__SCAN_IN), .B(n16998), .ZN(n16906) );
  AOI211_X1 U20073 ( .C1(n16998), .C2(n17108), .A(n16907), .B(n16906), .ZN(
        P3_U2692) );
  AOI22_X1 U20074 ( .A1(n16945), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16920) );
  AOI22_X1 U20075 ( .A1(n16927), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16919) );
  AOI22_X1 U20076 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16909) );
  OAI21_X1 U20077 ( .B1(n10944), .B2(n20848), .A(n16909), .ZN(n16917) );
  AOI22_X1 U20078 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16915) );
  AOI22_X1 U20079 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16911), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16914) );
  AOI22_X1 U20080 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n16944), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16913) );
  AOI22_X1 U20081 ( .A1(n16951), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16912) );
  NAND4_X1 U20082 ( .A1(n16915), .A2(n16914), .A3(n16913), .A4(n16912), .ZN(
        n16916) );
  AOI211_X1 U20083 ( .C1(n16962), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n16917), .B(n16916), .ZN(n16918) );
  NAND3_X1 U20084 ( .A1(n16920), .A2(n16919), .A3(n16918), .ZN(n17111) );
  INV_X1 U20085 ( .A(n17111), .ZN(n16925) );
  NOR2_X1 U20086 ( .A1(n16998), .A2(n16922), .ZN(n16940) );
  NOR2_X1 U20087 ( .A1(n16940), .A2(n16921), .ZN(n16924) );
  AOI21_X1 U20088 ( .B1(n18024), .B2(n16922), .A(P3_EBX_REG_10__SCAN_IN), .ZN(
        n16923) );
  OAI22_X1 U20089 ( .A1(n16925), .A2(n16980), .B1(n16924), .B2(n16923), .ZN(
        P3_U2693) );
  AOI22_X1 U20090 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16933) );
  AOI22_X1 U20091 ( .A1(n16962), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n16927), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n16932) );
  AOI22_X1 U20092 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n16931) );
  AOI22_X1 U20093 ( .A1(n16929), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n16928), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n16930) );
  NAND4_X1 U20094 ( .A1(n16933), .A2(n16932), .A3(n16931), .A4(n16930), .ZN(
        n16939) );
  AOI22_X1 U20095 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15525), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16937) );
  AOI22_X1 U20096 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16936) );
  AOI22_X1 U20097 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n16935) );
  AOI22_X1 U20098 ( .A1(n10858), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16934) );
  NAND4_X1 U20099 ( .A1(n16937), .A2(n16936), .A3(n16935), .A4(n16934), .ZN(
        n16938) );
  NOR2_X1 U20100 ( .A1(n16939), .A2(n16938), .ZN(n17116) );
  INV_X1 U20101 ( .A(n16966), .ZN(n16941) );
  OAI21_X1 U20102 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n16941), .A(n16940), .ZN(
        n16942) );
  OAI21_X1 U20103 ( .B1(n17116), .B2(n16980), .A(n16942), .ZN(P3_U2694) );
  AOI22_X1 U20104 ( .A1(n16944), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16943), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16965) );
  AOI22_X1 U20105 ( .A1(n16946), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16945), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16964) );
  AOI22_X1 U20106 ( .A1(n16926), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16947), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16948) );
  OAI21_X1 U20107 ( .B1(n16950), .B2(n16949), .A(n16948), .ZN(n16961) );
  AOI22_X1 U20108 ( .A1(n16952), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16951), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16959) );
  AOI22_X1 U20109 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16953), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16958) );
  AOI22_X1 U20110 ( .A1(n16954), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15523), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16957) );
  AOI22_X1 U20111 ( .A1(n16911), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16955), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16956) );
  NAND4_X1 U20112 ( .A1(n16959), .A2(n16958), .A3(n16957), .A4(n16956), .ZN(
        n16960) );
  AOI211_X1 U20113 ( .C1(n16962), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n16961), .B(n16960), .ZN(n16963) );
  NAND3_X1 U20114 ( .A1(n16965), .A2(n16964), .A3(n16963), .ZN(n17120) );
  INV_X1 U20115 ( .A(n17120), .ZN(n16968) );
  OAI21_X1 U20116 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n16971), .A(n16966), .ZN(
        n16967) );
  AOI22_X1 U20117 ( .A1(n16998), .A2(n16968), .B1(n16967), .B2(n16980), .ZN(
        P3_U2695) );
  NOR2_X1 U20118 ( .A1(n17092), .A2(n16972), .ZN(n16973) );
  AOI22_X1 U20119 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n16980), .B1(
        P3_EBX_REG_6__SCAN_IN), .B2(n16973), .ZN(n16970) );
  INV_X1 U20120 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16969) );
  OAI22_X1 U20121 ( .A1(n16971), .A2(n16970), .B1(n16969), .B2(n16980), .ZN(
        P3_U2696) );
  NAND2_X1 U20122 ( .A1(n16980), .A2(n16972), .ZN(n16977) );
  AOI22_X1 U20123 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n16998), .B1(
        n16973), .B2(n16975), .ZN(n16974) );
  OAI21_X1 U20124 ( .B1(n16975), .B2(n16977), .A(n16974), .ZN(P3_U2697) );
  NOR2_X1 U20125 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n16983), .ZN(n16978) );
  INV_X1 U20126 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16976) );
  OAI22_X1 U20127 ( .A1(n16978), .A2(n16977), .B1(n16976), .B2(n16980), .ZN(
        P3_U2698) );
  OAI21_X1 U20128 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n16979), .A(n16980), .ZN(
        n16982) );
  INV_X1 U20129 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16981) );
  OAI22_X1 U20130 ( .A1(n16983), .A2(n16982), .B1(n16981), .B2(n16980), .ZN(
        P3_U2699) );
  NAND2_X1 U20131 ( .A1(n18024), .A2(n16984), .ZN(n16986) );
  NOR2_X1 U20132 ( .A1(n16998), .A2(n16984), .ZN(n16988) );
  AOI22_X1 U20133 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n16998), .B1(
        P3_EBX_REG_3__SCAN_IN), .B2(n16988), .ZN(n16985) );
  OAI21_X1 U20134 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n16986), .A(n16985), .ZN(
        P3_U2700) );
  INV_X1 U20135 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16991) );
  INV_X1 U20136 ( .A(n16987), .ZN(n16989) );
  OAI21_X1 U20137 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n16989), .A(n16988), .ZN(
        n16990) );
  OAI21_X1 U20138 ( .B1(n16980), .B2(n16991), .A(n16990), .ZN(P3_U2701) );
  INV_X1 U20139 ( .A(n16992), .ZN(n16996) );
  OAI222_X1 U20140 ( .A1(n16996), .A2(n17000), .B1(n16995), .B2(n16994), .C1(
        n16993), .C2(n16980), .ZN(P3_U2702) );
  AOI22_X1 U20141 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n16998), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n16997), .ZN(n16999) );
  OAI21_X1 U20142 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17000), .A(n16999), .ZN(
        P3_U2703) );
  INV_X1 U20143 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17169) );
  INV_X1 U20144 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17173) );
  INV_X1 U20145 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17181) );
  INV_X1 U20146 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17270) );
  AND4_X1 U20147 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_3__SCAN_IN), 
        .A3(P3_EAX_REG_2__SCAN_IN), .A4(P3_EAX_REG_1__SCAN_IN), .ZN(n17001) );
  NAND4_X1 U20148 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_5__SCAN_IN), .A4(n17001), .ZN(n17129) );
  NOR2_X2 U20149 ( .A1(n17158), .A2(n17129), .ZN(n17123) );
  INV_X1 U20150 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n20711) );
  INV_X1 U20151 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17262) );
  INV_X1 U20152 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17198) );
  INV_X1 U20153 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17200) );
  NOR4_X1 U20154 ( .A1(n20711), .A2(n17262), .A3(n17198), .A4(n17200), .ZN(
        n17002) );
  NAND3_X1 U20155 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(n17002), .ZN(n17093) );
  NAND2_X1 U20156 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17095), .ZN(n17088) );
  NOR2_X2 U20157 ( .A1(n17270), .A2(n17088), .ZN(n17087) );
  INV_X1 U20158 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17189) );
  INV_X1 U20159 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17191) );
  NOR2_X1 U20160 ( .A1(n17189), .A2(n17191), .ZN(n17050) );
  NAND4_X1 U20161 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .A4(n17050), .ZN(n17048) );
  NAND2_X1 U20162 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17044), .ZN(n17043) );
  NAND2_X1 U20163 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17039), .ZN(n17038) );
  NAND2_X1 U20164 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17016), .ZN(n17012) );
  INV_X1 U20165 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17241) );
  OR2_X1 U20166 ( .A1(n17012), .A2(n17241), .ZN(n17005) );
  NOR2_X2 U20167 ( .A1(n18017), .A2(n17142), .ZN(n17081) );
  INV_X1 U20168 ( .A(n17154), .ZN(n17128) );
  NAND2_X1 U20169 ( .A1(n17142), .A2(n17012), .ZN(n17011) );
  OAI21_X1 U20170 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17128), .A(n17011), .ZN(
        n17003) );
  AOI22_X1 U20171 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17081), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17003), .ZN(n17004) );
  OAI21_X1 U20172 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17005), .A(n17004), .ZN(
        P3_U2704) );
  NAND2_X1 U20173 ( .A1(n17006), .A2(n17149), .ZN(n17075) );
  INV_X1 U20174 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n17007) );
  INV_X1 U20175 ( .A(n17081), .ZN(n17060) );
  OAI22_X1 U20176 ( .A1(n17008), .A2(n17144), .B1(n17007), .B2(n17060), .ZN(
        n17009) );
  AOI21_X1 U20177 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17082), .A(n17009), .ZN(
        n17010) );
  OAI221_X1 U20178 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17012), .C1(n17241), 
        .C2(n17011), .A(n17010), .ZN(P3_U2705) );
  AOI22_X1 U20179 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17082), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17081), .ZN(n17014) );
  OAI211_X1 U20180 ( .C1(n17016), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17142), .B(
        n17012), .ZN(n17013) );
  OAI211_X1 U20181 ( .C1(n17144), .C2(n17015), .A(n17014), .B(n17013), .ZN(
        P3_U2706) );
  AOI22_X1 U20182 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17082), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17081), .ZN(n17019) );
  AOI211_X1 U20183 ( .C1(n17169), .C2(n17024), .A(n17016), .B(n17149), .ZN(
        n17017) );
  INV_X1 U20184 ( .A(n17017), .ZN(n17018) );
  OAI211_X1 U20185 ( .C1(n17144), .C2(n17020), .A(n17019), .B(n17018), .ZN(
        P3_U2707) );
  OAI21_X1 U20186 ( .B1(n17023), .B2(n17022), .A(n17021), .ZN(n17027) );
  AOI22_X1 U20187 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17082), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17081), .ZN(n17026) );
  OAI211_X1 U20188 ( .C1(n17028), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17142), .B(
        n17024), .ZN(n17025) );
  OAI211_X1 U20189 ( .C1(n17027), .C2(n17144), .A(n17026), .B(n17025), .ZN(
        P3_U2708) );
  AOI22_X1 U20190 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17082), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17081), .ZN(n17031) );
  AOI211_X1 U20191 ( .C1(n17173), .C2(n17033), .A(n17028), .B(n17149), .ZN(
        n17029) );
  INV_X1 U20192 ( .A(n17029), .ZN(n17030) );
  OAI211_X1 U20193 ( .C1(n17032), .C2(n17144), .A(n17031), .B(n17030), .ZN(
        P3_U2709) );
  AOI22_X1 U20194 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17082), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17081), .ZN(n17036) );
  OAI211_X1 U20195 ( .C1(n17034), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17142), .B(
        n17033), .ZN(n17035) );
  OAI211_X1 U20196 ( .C1(n17144), .C2(n17037), .A(n17036), .B(n17035), .ZN(
        P3_U2710) );
  AOI22_X1 U20197 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17082), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17081), .ZN(n17041) );
  OAI211_X1 U20198 ( .C1(n17039), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17142), .B(
        n17038), .ZN(n17040) );
  OAI211_X1 U20199 ( .C1(n17144), .C2(n17042), .A(n17041), .B(n17040), .ZN(
        P3_U2711) );
  AOI22_X1 U20200 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17082), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17081), .ZN(n17046) );
  OAI211_X1 U20201 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17044), .A(n17142), .B(
        n17043), .ZN(n17045) );
  OAI211_X1 U20202 ( .C1(n17047), .C2(n17144), .A(n17046), .B(n17045), .ZN(
        P3_U2712) );
  INV_X1 U20203 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18016) );
  INV_X1 U20204 ( .A(n17048), .ZN(n17049) );
  NOR2_X1 U20205 ( .A1(n17092), .A2(n17083), .ZN(n17077) );
  NAND2_X1 U20206 ( .A1(n17049), .A2(n17077), .ZN(n17057) );
  INV_X1 U20207 ( .A(n17057), .ZN(n17054) );
  INV_X1 U20208 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17185) );
  NAND2_X1 U20209 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17072), .ZN(n17066) );
  NOR2_X1 U20210 ( .A1(n17185), .A2(n17066), .ZN(n17061) );
  OAI22_X1 U20211 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17128), .B1(n17149), 
        .B2(n17061), .ZN(n17053) );
  INV_X1 U20212 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n19056) );
  OAI22_X1 U20213 ( .A1(n17051), .A2(n17144), .B1(n19056), .B2(n17060), .ZN(
        n17052) );
  AOI221_X1 U20214 ( .B1(n17054), .B2(n17181), .C1(n17053), .C2(
        P3_EAX_REG_22__SCAN_IN), .A(n17052), .ZN(n17055) );
  OAI21_X1 U20215 ( .B1(n18016), .B2(n17075), .A(n17055), .ZN(P3_U2713) );
  INV_X1 U20216 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18013) );
  AOI22_X1 U20217 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17082), .B1(n17155), .B2(
        n17056), .ZN(n17059) );
  OAI211_X1 U20218 ( .C1(n17061), .C2(P3_EAX_REG_21__SCAN_IN), .A(n17142), .B(
        n17057), .ZN(n17058) );
  OAI211_X1 U20219 ( .C1(n17060), .C2(n18013), .A(n17059), .B(n17058), .ZN(
        P3_U2714) );
  AOI22_X1 U20220 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17082), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17081), .ZN(n17064) );
  AOI211_X1 U20221 ( .C1(n17185), .C2(n17066), .A(n17061), .B(n17149), .ZN(
        n17062) );
  INV_X1 U20222 ( .A(n17062), .ZN(n17063) );
  OAI211_X1 U20223 ( .C1(n17065), .C2(n17144), .A(n17064), .B(n17063), .ZN(
        P3_U2715) );
  AOI22_X1 U20224 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17082), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17081), .ZN(n17068) );
  OAI211_X1 U20225 ( .C1(n17072), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17142), .B(
        n17066), .ZN(n17067) );
  OAI211_X1 U20226 ( .C1(n17069), .C2(n17144), .A(n17068), .B(n17067), .ZN(
        P3_U2716) );
  INV_X1 U20227 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n17994) );
  AOI22_X1 U20228 ( .A1(n17077), .A2(P3_EAX_REG_17__SCAN_IN), .B1(
        P3_EAX_REG_18__SCAN_IN), .B2(n17142), .ZN(n17071) );
  OAI22_X1 U20229 ( .A1(n17072), .A2(n17071), .B1(n17070), .B2(n17144), .ZN(
        n17073) );
  AOI21_X1 U20230 ( .B1(BUF2_REG_18__SCAN_IN), .B2(n17081), .A(n17073), .ZN(
        n17074) );
  OAI21_X1 U20231 ( .B1(n17994), .B2(n17075), .A(n17074), .ZN(P3_U2717) );
  AOI22_X1 U20232 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17082), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17081), .ZN(n17079) );
  NAND2_X1 U20233 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17077), .ZN(n17076) );
  OAI211_X1 U20234 ( .C1(n17077), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17142), .B(
        n17076), .ZN(n17078) );
  OAI211_X1 U20235 ( .C1(n17080), .C2(n17144), .A(n17079), .B(n17078), .ZN(
        P3_U2718) );
  AOI22_X1 U20236 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17082), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17081), .ZN(n17085) );
  OAI211_X1 U20237 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17087), .A(n17142), .B(
        n17083), .ZN(n17084) );
  OAI211_X1 U20238 ( .C1(n17086), .C2(n17144), .A(n17085), .B(n17084), .ZN(
        P3_U2719) );
  AOI211_X1 U20239 ( .C1(n17270), .C2(n17088), .A(n17149), .B(n17087), .ZN(
        n17089) );
  AOI21_X1 U20240 ( .B1(n17156), .B2(BUF2_REG_15__SCAN_IN), .A(n17089), .ZN(
        n17090) );
  OAI21_X1 U20241 ( .B1(n17091), .B2(n17144), .A(n17090), .ZN(P3_U2720) );
  NOR2_X1 U20242 ( .A1(n17092), .A2(n17119), .ZN(n17099) );
  NOR2_X1 U20243 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17093), .ZN(n17094) );
  AOI22_X1 U20244 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17156), .B1(n17099), .B2(
        n17094), .ZN(n17097) );
  INV_X1 U20245 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17265) );
  OR3_X1 U20246 ( .A1(n17265), .A2(n17149), .A3(n17095), .ZN(n17096) );
  OAI211_X1 U20247 ( .C1(n17098), .C2(n17144), .A(n17097), .B(n17096), .ZN(
        P3_U2721) );
  INV_X1 U20248 ( .A(n17099), .ZN(n17122) );
  NOR2_X1 U20249 ( .A1(n20711), .A2(n17122), .ZN(n17115) );
  NAND2_X1 U20250 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17118), .ZN(n17112) );
  NOR2_X1 U20251 ( .A1(n17200), .A2(n17112), .ZN(n17110) );
  NAND2_X1 U20252 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17110), .ZN(n17103) );
  NAND2_X1 U20253 ( .A1(n17103), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n17102) );
  AOI22_X1 U20254 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17156), .B1(n17155), .B2(
        n17100), .ZN(n17101) );
  OAI221_X1 U20255 ( .B1(n17103), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n17102), 
        .C2(n17149), .A(n17101), .ZN(P3_U2722) );
  INV_X1 U20256 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n20725) );
  INV_X1 U20257 ( .A(n17103), .ZN(n17106) );
  AOI21_X1 U20258 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17142), .A(n17110), .ZN(
        n17105) );
  OAI222_X1 U20259 ( .A1(n17147), .A2(n20725), .B1(n17106), .B2(n17105), .C1(
        n17144), .C2(n17104), .ZN(P3_U2723) );
  OAI21_X1 U20260 ( .B1(n17200), .B2(n17149), .A(n17112), .ZN(n17107) );
  INV_X1 U20261 ( .A(n17107), .ZN(n17109) );
  OAI222_X1 U20262 ( .A1(n17147), .A2(n17257), .B1(n17110), .B2(n17109), .C1(
        n17144), .C2(n17108), .ZN(P3_U2724) );
  AOI22_X1 U20263 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17156), .B1(n17155), .B2(
        n17111), .ZN(n17114) );
  OAI211_X1 U20264 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17118), .A(n17142), .B(
        n17112), .ZN(n17113) );
  NAND2_X1 U20265 ( .A1(n17114), .A2(n17113), .ZN(P3_U2725) );
  AOI21_X1 U20266 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17142), .A(n17115), .ZN(
        n17117) );
  OAI222_X1 U20267 ( .A1(n17147), .A2(n17253), .B1(n17118), .B2(n17117), .C1(
        n17144), .C2(n17116), .ZN(P3_U2726) );
  NAND2_X1 U20268 ( .A1(n17142), .A2(n17119), .ZN(n17125) );
  AOI22_X1 U20269 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17156), .B1(n17155), .B2(
        n17120), .ZN(n17121) );
  OAI221_X1 U20270 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n17122), .C1(n20711), 
        .C2(n17125), .A(n17121), .ZN(P3_U2727) );
  NOR2_X1 U20271 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17123), .ZN(n17124) );
  OAI222_X1 U20272 ( .A1(n17147), .A2(n18021), .B1(n17144), .B2(n17126), .C1(
        n17125), .C2(n17124), .ZN(P3_U2728) );
  NAND2_X1 U20273 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .ZN(n17127) );
  INV_X1 U20274 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17213) );
  INV_X1 U20275 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17215) );
  NAND3_X1 U20276 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .A3(n17154), .ZN(n17148) );
  NOR2_X1 U20277 ( .A1(n17215), .A2(n17148), .ZN(n17141) );
  INV_X1 U20278 ( .A(n17141), .ZN(n17152) );
  NOR2_X1 U20279 ( .A1(n17213), .A2(n17152), .ZN(n17146) );
  INV_X1 U20280 ( .A(n17146), .ZN(n17136) );
  NOR2_X1 U20281 ( .A1(n17127), .A2(n17136), .ZN(n17135) );
  AOI21_X1 U20282 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17142), .A(n17135), .ZN(
        n17132) );
  NOR2_X1 U20283 ( .A1(n17129), .A2(n17128), .ZN(n17131) );
  OAI222_X1 U20284 ( .A1(n18016), .A2(n17147), .B1(n17132), .B2(n17131), .C1(
        n17144), .C2(n17130), .ZN(P3_U2729) );
  AOI22_X1 U20285 ( .A1(n17146), .A2(P3_EAX_REG_4__SCAN_IN), .B1(
        P3_EAX_REG_5__SCAN_IN), .B2(n17142), .ZN(n17134) );
  OAI222_X1 U20286 ( .A1(n18012), .A2(n17147), .B1(n17135), .B2(n17134), .C1(
        n17144), .C2(n17133), .ZN(P3_U2730) );
  INV_X1 U20287 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18004) );
  INV_X1 U20288 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n20752) );
  NOR2_X1 U20289 ( .A1(n20752), .A2(n17136), .ZN(n17140) );
  AOI21_X1 U20290 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17142), .A(n17146), .ZN(
        n17139) );
  INV_X1 U20291 ( .A(n17137), .ZN(n17138) );
  OAI222_X1 U20292 ( .A1(n18004), .A2(n17147), .B1(n17140), .B2(n17139), .C1(
        n17144), .C2(n17138), .ZN(P3_U2731) );
  AOI21_X1 U20293 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17142), .A(n17141), .ZN(
        n17145) );
  OAI222_X1 U20294 ( .A1(n17999), .A2(n17147), .B1(n17146), .B2(n17145), .C1(
        n17144), .C2(n17143), .ZN(P3_U2732) );
  OAI21_X1 U20295 ( .B1(n17215), .B2(n17149), .A(n17148), .ZN(n17151) );
  AOI222_X1 U20296 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17156), .B1(n17152), .B2(
        n17151), .C1(n17155), .C2(n17150), .ZN(n17153) );
  INV_X1 U20297 ( .A(n17153), .ZN(P3_U2733) );
  NAND2_X1 U20298 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17154), .ZN(n17162) );
  AOI22_X1 U20299 ( .A1(n17156), .A2(BUF2_REG_1__SCAN_IN), .B1(n17155), .B2(
        n10905), .ZN(n17161) );
  INV_X1 U20300 ( .A(n17157), .ZN(n17159) );
  OAI21_X1 U20301 ( .B1(n17159), .B2(n17158), .A(P3_EAX_REG_1__SCAN_IN), .ZN(
        n17160) );
  OAI211_X1 U20302 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n17162), .A(n17161), .B(
        n17160), .ZN(P3_U2734) );
  NOR2_X1 U20303 ( .A1(n18605), .A2(n17644), .ZN(n18628) );
  NOR2_X1 U20304 ( .A1(n17218), .A2(n17165), .ZN(P3_U2736) );
  NAND2_X1 U20305 ( .A1(n17216), .A2(n17988), .ZN(n17193) );
  INV_X2 U20306 ( .A(n17218), .ZN(n17219) );
  AOI22_X1 U20307 ( .A1(n18628), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17166) );
  OAI21_X1 U20308 ( .B1(n17241), .B2(n17193), .A(n17166), .ZN(P3_U2737) );
  INV_X1 U20309 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17239) );
  AOI22_X1 U20310 ( .A1(n18628), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17167) );
  OAI21_X1 U20311 ( .B1(n17239), .B2(n17193), .A(n17167), .ZN(P3_U2738) );
  AOI22_X1 U20312 ( .A1(n18628), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17168) );
  OAI21_X1 U20313 ( .B1(n17169), .B2(n17193), .A(n17168), .ZN(P3_U2739) );
  INV_X1 U20314 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17171) );
  AOI22_X1 U20315 ( .A1(n18628), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17170) );
  OAI21_X1 U20316 ( .B1(n17171), .B2(n17193), .A(n17170), .ZN(P3_U2740) );
  AOI22_X1 U20317 ( .A1(n18628), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17172) );
  OAI21_X1 U20318 ( .B1(n17173), .B2(n17193), .A(n17172), .ZN(P3_U2741) );
  INV_X1 U20319 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17175) );
  AOI22_X1 U20320 ( .A1(n18628), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17174) );
  OAI21_X1 U20321 ( .B1(n17175), .B2(n17193), .A(n17174), .ZN(P3_U2742) );
  INV_X1 U20322 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17177) );
  AOI22_X1 U20323 ( .A1(n18628), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17176) );
  OAI21_X1 U20324 ( .B1(n17177), .B2(n17193), .A(n17176), .ZN(P3_U2743) );
  INV_X1 U20325 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17179) );
  CLKBUF_X1 U20326 ( .A(n18628), .Z(n18480) );
  AOI22_X1 U20327 ( .A1(n18480), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17178) );
  OAI21_X1 U20328 ( .B1(n17179), .B2(n17193), .A(n17178), .ZN(P3_U2744) );
  AOI22_X1 U20329 ( .A1(n18480), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17180) );
  OAI21_X1 U20330 ( .B1(n17181), .B2(n17193), .A(n17180), .ZN(P3_U2745) );
  INV_X1 U20331 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17183) );
  AOI22_X1 U20332 ( .A1(n18480), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17182) );
  OAI21_X1 U20333 ( .B1(n17183), .B2(n17193), .A(n17182), .ZN(P3_U2746) );
  AOI22_X1 U20334 ( .A1(n18480), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17184) );
  OAI21_X1 U20335 ( .B1(n17185), .B2(n17193), .A(n17184), .ZN(P3_U2747) );
  INV_X1 U20336 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17187) );
  AOI22_X1 U20337 ( .A1(n18480), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17186) );
  OAI21_X1 U20338 ( .B1(n17187), .B2(n17193), .A(n17186), .ZN(P3_U2748) );
  AOI22_X1 U20339 ( .A1(n18480), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17188) );
  OAI21_X1 U20340 ( .B1(n17189), .B2(n17193), .A(n17188), .ZN(P3_U2749) );
  AOI22_X1 U20341 ( .A1(n18480), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17190) );
  OAI21_X1 U20342 ( .B1(n17191), .B2(n17193), .A(n17190), .ZN(P3_U2750) );
  INV_X1 U20343 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n20708) );
  AOI22_X1 U20344 ( .A1(n18480), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17192) );
  OAI21_X1 U20345 ( .B1(n20708), .B2(n17193), .A(n17192), .ZN(P3_U2751) );
  INV_X1 U20346 ( .A(n17216), .ZN(n17221) );
  AOI22_X1 U20347 ( .A1(n18480), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17194) );
  OAI21_X1 U20348 ( .B1(n17270), .B2(n17221), .A(n17194), .ZN(P3_U2752) );
  AOI22_X1 U20349 ( .A1(n18480), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17195) );
  OAI21_X1 U20350 ( .B1(n17265), .B2(n17221), .A(n17195), .ZN(P3_U2753) );
  AOI22_X1 U20351 ( .A1(n18480), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17196) );
  OAI21_X1 U20352 ( .B1(n17262), .B2(n17221), .A(n17196), .ZN(P3_U2754) );
  AOI22_X1 U20353 ( .A1(n18480), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17197) );
  OAI21_X1 U20354 ( .B1(n17198), .B2(n17221), .A(n17197), .ZN(P3_U2755) );
  AOI22_X1 U20355 ( .A1(n18480), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17199) );
  OAI21_X1 U20356 ( .B1(n17200), .B2(n17221), .A(n17199), .ZN(P3_U2756) );
  INV_X1 U20357 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17202) );
  AOI22_X1 U20358 ( .A1(n18480), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17201) );
  OAI21_X1 U20359 ( .B1(n17202), .B2(n17221), .A(n17201), .ZN(P3_U2757) );
  INV_X1 U20360 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17204) );
  AOI22_X1 U20361 ( .A1(n18480), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17203) );
  OAI21_X1 U20362 ( .B1(n17204), .B2(n17221), .A(n17203), .ZN(P3_U2758) );
  AOI22_X1 U20363 ( .A1(n18480), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17205) );
  OAI21_X1 U20364 ( .B1(n20711), .B2(n17221), .A(n17205), .ZN(P3_U2759) );
  INV_X1 U20365 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n20740) );
  AOI22_X1 U20366 ( .A1(n18480), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17206) );
  OAI21_X1 U20367 ( .B1(n20740), .B2(n17221), .A(n17206), .ZN(P3_U2760) );
  INV_X1 U20368 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17208) );
  AOI22_X1 U20369 ( .A1(n18480), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17207) );
  OAI21_X1 U20370 ( .B1(n17208), .B2(n17221), .A(n17207), .ZN(P3_U2761) );
  INV_X1 U20371 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17210) );
  AOI22_X1 U20372 ( .A1(n18480), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17209) );
  OAI21_X1 U20373 ( .B1(n17210), .B2(n17221), .A(n17209), .ZN(P3_U2762) );
  AOI22_X1 U20374 ( .A1(n18480), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17211) );
  OAI21_X1 U20375 ( .B1(n20752), .B2(n17221), .A(n17211), .ZN(P3_U2763) );
  AOI22_X1 U20376 ( .A1(n18480), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17212) );
  OAI21_X1 U20377 ( .B1(n17213), .B2(n17221), .A(n17212), .ZN(P3_U2764) );
  AOI22_X1 U20378 ( .A1(n18480), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17214) );
  OAI21_X1 U20379 ( .B1(n17215), .B2(n17221), .A(n17214), .ZN(P3_U2765) );
  INV_X1 U20380 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n20705) );
  AOI22_X1 U20381 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17216), .B1(n18628), .B2(
        P3_LWORD_REG_1__SCAN_IN), .ZN(n17217) );
  OAI21_X1 U20382 ( .B1(n20705), .B2(n17218), .A(n17217), .ZN(P3_U2766) );
  AOI22_X1 U20383 ( .A1(n18480), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17219), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17220) );
  OAI21_X1 U20384 ( .B1(n17222), .B2(n17221), .A(n17220), .ZN(P3_U2767) );
  INV_X1 U20385 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n17983) );
  OAI211_X1 U20386 ( .C1(n18632), .C2(n18631), .A(n17224), .B(n17223), .ZN(
        n17263) );
  INV_X2 U20387 ( .A(n17267), .ZN(n17260) );
  NAND3_X1 U20388 ( .A1(n18631), .A2(n17224), .A3(n17223), .ZN(n17269) );
  INV_X2 U20389 ( .A(n17269), .ZN(n17258) );
  AOI22_X1 U20390 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17258), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17266), .ZN(n17225) );
  OAI21_X1 U20391 ( .B1(n17983), .B2(n17260), .A(n17225), .ZN(P3_U2768) );
  AOI22_X1 U20392 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17258), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17266), .ZN(n17226) );
  OAI21_X1 U20393 ( .B1(n20751), .B2(n17260), .A(n17226), .ZN(P3_U2769) );
  AOI22_X1 U20394 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17258), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17266), .ZN(n17227) );
  OAI21_X1 U20395 ( .B1(n17994), .B2(n17260), .A(n17227), .ZN(P3_U2770) );
  AOI22_X1 U20396 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17258), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17266), .ZN(n17228) );
  OAI21_X1 U20397 ( .B1(n17999), .B2(n17260), .A(n17228), .ZN(P3_U2771) );
  AOI22_X1 U20398 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17258), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17266), .ZN(n17229) );
  OAI21_X1 U20399 ( .B1(n18004), .B2(n17260), .A(n17229), .ZN(P3_U2772) );
  AOI22_X1 U20400 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17258), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17266), .ZN(n17230) );
  OAI21_X1 U20401 ( .B1(n18012), .B2(n17260), .A(n17230), .ZN(P3_U2773) );
  AOI22_X1 U20402 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17258), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17266), .ZN(n17231) );
  OAI21_X1 U20403 ( .B1(n18016), .B2(n17260), .A(n17231), .ZN(P3_U2774) );
  AOI22_X1 U20404 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17258), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17266), .ZN(n17232) );
  OAI21_X1 U20405 ( .B1(n18021), .B2(n17260), .A(n17232), .ZN(P3_U2775) );
  INV_X1 U20406 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17251) );
  AOI22_X1 U20407 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17258), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17266), .ZN(n17233) );
  OAI21_X1 U20408 ( .B1(n17251), .B2(n17260), .A(n17233), .ZN(P3_U2776) );
  AOI22_X1 U20409 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17258), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17266), .ZN(n17234) );
  OAI21_X1 U20410 ( .B1(n17253), .B2(n17260), .A(n17234), .ZN(P3_U2777) );
  INV_X1 U20411 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17255) );
  AOI22_X1 U20412 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17258), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17266), .ZN(n17235) );
  OAI21_X1 U20413 ( .B1(n17255), .B2(n17260), .A(n17235), .ZN(P3_U2778) );
  AOI22_X1 U20414 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17258), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17266), .ZN(n17236) );
  OAI21_X1 U20415 ( .B1(n17257), .B2(n17260), .A(n17236), .ZN(P3_U2779) );
  AOI22_X1 U20416 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17258), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17266), .ZN(n17237) );
  OAI21_X1 U20417 ( .B1(n20725), .B2(n17260), .A(n17237), .ZN(P3_U2780) );
  AOI22_X1 U20418 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17267), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17266), .ZN(n17238) );
  OAI21_X1 U20419 ( .B1(n17239), .B2(n17269), .A(n17238), .ZN(P3_U2781) );
  AOI22_X1 U20420 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17267), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17266), .ZN(n17240) );
  OAI21_X1 U20421 ( .B1(n17241), .B2(n17269), .A(n17240), .ZN(P3_U2782) );
  AOI22_X1 U20422 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17258), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17266), .ZN(n17242) );
  OAI21_X1 U20423 ( .B1(n17983), .B2(n17260), .A(n17242), .ZN(P3_U2783) );
  AOI22_X1 U20424 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17258), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17266), .ZN(n17243) );
  OAI21_X1 U20425 ( .B1(n20751), .B2(n17260), .A(n17243), .ZN(P3_U2784) );
  AOI22_X1 U20426 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17258), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17266), .ZN(n17244) );
  OAI21_X1 U20427 ( .B1(n17994), .B2(n17260), .A(n17244), .ZN(P3_U2785) );
  AOI22_X1 U20428 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17258), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17263), .ZN(n17245) );
  OAI21_X1 U20429 ( .B1(n17999), .B2(n17260), .A(n17245), .ZN(P3_U2786) );
  AOI22_X1 U20430 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17258), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17263), .ZN(n17246) );
  OAI21_X1 U20431 ( .B1(n18004), .B2(n17260), .A(n17246), .ZN(P3_U2787) );
  AOI22_X1 U20432 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17258), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17263), .ZN(n17247) );
  OAI21_X1 U20433 ( .B1(n18012), .B2(n17260), .A(n17247), .ZN(P3_U2788) );
  AOI22_X1 U20434 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17258), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17263), .ZN(n17248) );
  OAI21_X1 U20435 ( .B1(n18016), .B2(n17260), .A(n17248), .ZN(P3_U2789) );
  AOI22_X1 U20436 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17258), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17263), .ZN(n17249) );
  OAI21_X1 U20437 ( .B1(n18021), .B2(n17260), .A(n17249), .ZN(P3_U2790) );
  AOI22_X1 U20438 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17258), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17263), .ZN(n17250) );
  OAI21_X1 U20439 ( .B1(n17251), .B2(n17260), .A(n17250), .ZN(P3_U2791) );
  AOI22_X1 U20440 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17258), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17263), .ZN(n17252) );
  OAI21_X1 U20441 ( .B1(n17253), .B2(n17260), .A(n17252), .ZN(P3_U2792) );
  AOI22_X1 U20442 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17258), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17263), .ZN(n17254) );
  OAI21_X1 U20443 ( .B1(n17255), .B2(n17260), .A(n17254), .ZN(P3_U2793) );
  AOI22_X1 U20444 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17258), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17266), .ZN(n17256) );
  OAI21_X1 U20445 ( .B1(n17257), .B2(n17260), .A(n17256), .ZN(P3_U2794) );
  AOI22_X1 U20446 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17258), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17266), .ZN(n17259) );
  OAI21_X1 U20447 ( .B1(n20725), .B2(n17260), .A(n17259), .ZN(P3_U2795) );
  AOI22_X1 U20448 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17267), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17263), .ZN(n17261) );
  OAI21_X1 U20449 ( .B1(n17262), .B2(n17269), .A(n17261), .ZN(P3_U2796) );
  AOI22_X1 U20450 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17267), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17263), .ZN(n17264) );
  OAI21_X1 U20451 ( .B1(n17265), .B2(n17269), .A(n17264), .ZN(P3_U2797) );
  AOI22_X1 U20452 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17267), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17266), .ZN(n17268) );
  OAI21_X1 U20453 ( .B1(n17270), .B2(n17269), .A(n17268), .ZN(P3_U2798) );
  NAND2_X1 U20454 ( .A1(n17271), .A2(n17372), .ZN(n17356) );
  OR2_X1 U20455 ( .A1(n17272), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17289) );
  NOR2_X1 U20456 ( .A1(n17552), .A2(n17633), .ZN(n17388) );
  INV_X1 U20457 ( .A(n17273), .ZN(n17656) );
  OAI22_X1 U20458 ( .A1(n17656), .A2(n17454), .B1(n17274), .B2(n17648), .ZN(
        n17309) );
  NOR2_X1 U20459 ( .A1(n10936), .A2(n17309), .ZN(n17294) );
  NOR3_X1 U20460 ( .A1(n17388), .A2(n17294), .A3(n20801), .ZN(n17283) );
  NAND3_X1 U20461 ( .A1(n17275), .A2(n9884), .A3(n17407), .ZN(n17280) );
  NOR3_X1 U20462 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17486), .A3(
        n12194), .ZN(n17297) );
  INV_X1 U20463 ( .A(n17644), .ZN(n17473) );
  INV_X1 U20464 ( .A(n17541), .ZN(n17603) );
  OAI21_X1 U20465 ( .B1(n17276), .B2(n17603), .A(n17643), .ZN(n17277) );
  AOI21_X1 U20466 ( .B1(n17473), .B2(n17278), .A(n17277), .ZN(n17303) );
  OAI21_X1 U20467 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17384), .A(
        n17303), .ZN(n17298) );
  OAI21_X1 U20468 ( .B1(n17297), .B2(n17298), .A(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17279) );
  OAI211_X1 U20469 ( .C1(n17504), .C2(n17281), .A(n17280), .B(n17279), .ZN(
        n17282) );
  AOI211_X1 U20470 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17965), .A(n17283), 
        .B(n17282), .ZN(n17288) );
  OAI211_X1 U20471 ( .C1(n17286), .C2(n17285), .A(n17537), .B(n17284), .ZN(
        n17287) );
  OAI211_X1 U20472 ( .C1(n17356), .C2(n17289), .A(n17288), .B(n17287), .ZN(
        P3_U2802) );
  NAND2_X1 U20473 ( .A1(n17291), .A2(n17290), .ZN(n17292) );
  XOR2_X1 U20474 ( .A(n17546), .B(n17292), .Z(n17664) );
  AOI22_X1 U20475 ( .A1(n17965), .A2(P3_REIP_REG_27__SCAN_IN), .B1(n17476), 
        .B2(n17293), .ZN(n17300) );
  OR2_X1 U20476 ( .A1(n17649), .A2(n17444), .ZN(n17295) );
  AOI21_X1 U20477 ( .B1(n10936), .B2(n17295), .A(n17294), .ZN(n17296) );
  AOI211_X1 U20478 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17298), .A(
        n17297), .B(n17296), .ZN(n17299) );
  OAI211_X1 U20479 ( .C1(n17664), .C2(n17549), .A(n17300), .B(n17299), .ZN(
        P3_U2803) );
  AOI21_X1 U20480 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17302), .A(
        n17301), .ZN(n17671) );
  AOI221_X1 U20481 ( .B1(n17305), .B2(n17304), .C1(n18006), .C2(n17304), .A(
        n17303), .ZN(n17308) );
  AOI21_X1 U20482 ( .B1(n17504), .B2(n17384), .A(n9893), .ZN(n17307) );
  AOI211_X1 U20483 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n17965), .A(n17308), 
        .B(n17307), .ZN(n17312) );
  OAI21_X1 U20484 ( .B1(n17667), .B2(n17356), .A(n17666), .ZN(n17310) );
  NAND2_X1 U20485 ( .A1(n17310), .A2(n17309), .ZN(n17311) );
  OAI211_X1 U20486 ( .C1(n17671), .C2(n17549), .A(n17312), .B(n17311), .ZN(
        P3_U2804) );
  OAI21_X1 U20487 ( .B1(n17546), .B2(n17314), .A(n17313), .ZN(n17315) );
  XOR2_X1 U20488 ( .A(n17315), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17686) );
  OAI21_X1 U20489 ( .B1(n17330), .B2(n18006), .A(n17643), .ZN(n17316) );
  AOI21_X1 U20490 ( .B1(n17473), .B2(n17344), .A(n17316), .ZN(n17346) );
  OAI21_X1 U20491 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17384), .A(
        n17346), .ZN(n17335) );
  NOR2_X1 U20492 ( .A1(n17963), .A2(n18559), .ZN(n17681) );
  NOR2_X1 U20493 ( .A1(n17318), .A2(n17317), .ZN(n17321) );
  OAI211_X1 U20494 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17330), .B(n17407), .ZN(n17320) );
  OAI22_X1 U20495 ( .A1(n17321), .A2(n17320), .B1(n17319), .B2(n17504), .ZN(
        n17322) );
  AOI211_X1 U20496 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17335), .A(
        n17681), .B(n17322), .ZN(n17327) );
  AOI21_X1 U20497 ( .B1(n17678), .B2(n17324), .A(n17323), .ZN(n17682) );
  INV_X1 U20498 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17695) );
  NOR3_X1 U20499 ( .A1(n17788), .A2(n17336), .A3(n17695), .ZN(n17325) );
  XOR2_X1 U20500 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17325), .Z(
        n17683) );
  AOI22_X1 U20501 ( .A1(n17552), .A2(n17682), .B1(n17633), .B2(n17683), .ZN(
        n17326) );
  OAI211_X1 U20502 ( .C1(n17549), .C2(n17686), .A(n17327), .B(n17326), .ZN(
        P3_U2805) );
  AOI21_X1 U20503 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17329), .A(
        n17328), .ZN(n17701) );
  NOR2_X1 U20504 ( .A1(n17963), .A2(n18557), .ZN(n17698) );
  NAND2_X1 U20505 ( .A1(n17330), .A2(n17407), .ZN(n17333) );
  INV_X1 U20506 ( .A(n17331), .ZN(n17332) );
  OAI22_X1 U20507 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17333), .B1(
        n17332), .B2(n17504), .ZN(n17334) );
  AOI211_X1 U20508 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n17335), .A(
        n17698), .B(n17334), .ZN(n17338) );
  NOR2_X1 U20509 ( .A1(n17336), .A2(n17788), .ZN(n17688) );
  OAI22_X1 U20510 ( .A1(n17690), .A2(n17454), .B1(n17688), .B2(n17648), .ZN(
        n17353) );
  NOR2_X1 U20511 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17336), .ZN(
        n17699) );
  AOI22_X1 U20512 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17353), .B1(
        n17372), .B2(n17699), .ZN(n17337) );
  OAI211_X1 U20513 ( .C1(n17701), .C2(n17549), .A(n17338), .B(n17337), .ZN(
        P3_U2806) );
  NOR2_X1 U20514 ( .A1(n17963), .A2(n18556), .ZN(n17705) );
  INV_X1 U20515 ( .A(n17339), .ZN(n17340) );
  AOI21_X1 U20516 ( .B1(n17340), .B2(n18364), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17345) );
  NAND2_X1 U20517 ( .A1(n17342), .A2(n17341), .ZN(n17343) );
  OAI22_X1 U20518 ( .A1(n17346), .A2(n17345), .B1(n17344), .B2(n17343), .ZN(
        n17347) );
  AOI211_X1 U20519 ( .C1(n17476), .C2(n17348), .A(n17705), .B(n17347), .ZN(
        n17355) );
  AOI22_X1 U20520 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17546), .B1(
        n17350), .B2(n17363), .ZN(n17351) );
  NAND2_X1 U20521 ( .A1(n17349), .A2(n17351), .ZN(n17352) );
  XOR2_X1 U20522 ( .A(n17352), .B(n17702), .Z(n17706) );
  AOI22_X1 U20523 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17353), .B1(
        n17537), .B2(n17706), .ZN(n17354) );
  OAI211_X1 U20524 ( .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n17356), .A(
        n17355), .B(n17354), .ZN(P3_U2807) );
  OAI21_X1 U20525 ( .B1(n9756), .B2(n17603), .A(n17643), .ZN(n17357) );
  AOI21_X1 U20526 ( .B1(n17473), .B2(n17358), .A(n17357), .ZN(n17385) );
  OAI21_X1 U20527 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17384), .A(
        n17385), .ZN(n17376) );
  AOI22_X1 U20528 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17376), .B1(
        n17476), .B2(n17359), .ZN(n17371) );
  NAND2_X1 U20529 ( .A1(n9756), .A2(n17407), .ZN(n17374) );
  AOI221_X1 U20530 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C1(n17361), .C2(n17360), .A(
        n17374), .ZN(n17362) );
  AOI21_X1 U20531 ( .B1(P3_REIP_REG_22__SCAN_IN), .B2(n17965), .A(n17362), 
        .ZN(n17370) );
  AOI22_X1 U20532 ( .A1(n17552), .A2(n17712), .B1(n17633), .B2(n17788), .ZN(
        n17443) );
  OAI21_X1 U20533 ( .B1(n17651), .B2(n17388), .A(n17443), .ZN(n17381) );
  INV_X1 U20534 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17726) );
  INV_X1 U20535 ( .A(n17363), .ZN(n17366) );
  INV_X1 U20536 ( .A(n17377), .ZN(n17365) );
  OAI221_X1 U20537 ( .B1(n17366), .B2(n17365), .C1(n17366), .C2(n17364), .A(
        n17349), .ZN(n17367) );
  XOR2_X1 U20538 ( .A(n17726), .B(n17367), .Z(n17710) );
  AOI22_X1 U20539 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17381), .B1(
        n17537), .B2(n17710), .ZN(n17369) );
  NAND3_X1 U20540 ( .A1(n17651), .A2(n17372), .A3(n17726), .ZN(n17368) );
  NAND4_X1 U20541 ( .A1(n17371), .A2(n17370), .A3(n17369), .A4(n17368), .ZN(
        P3_U2808) );
  NAND2_X1 U20542 ( .A1(n17732), .A2(n17718), .ZN(n17736) );
  NAND2_X1 U20543 ( .A1(n17730), .A2(n17372), .ZN(n17405) );
  NOR2_X1 U20544 ( .A1(n17963), .A2(n18552), .ZN(n17728) );
  OAI22_X1 U20545 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17374), .B1(
        n17373), .B2(n17504), .ZN(n17375) );
  AOI211_X1 U20546 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n17376), .A(
        n17728), .B(n17375), .ZN(n17383) );
  NOR3_X1 U20547 ( .A1(n17546), .A2(n17406), .A3(n17377), .ZN(n17399) );
  INV_X1 U20548 ( .A(n17378), .ZN(n17415) );
  AOI22_X1 U20549 ( .A1(n17732), .A2(n17399), .B1(n17415), .B2(n17379), .ZN(
        n17380) );
  XOR2_X1 U20550 ( .A(n17718), .B(n17380), .Z(n17729) );
  AOI22_X1 U20551 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17381), .B1(
        n17537), .B2(n17729), .ZN(n17382) );
  OAI211_X1 U20552 ( .C1(n17736), .C2(n17405), .A(n17383), .B(n17382), .ZN(
        P3_U2809) );
  OR2_X1 U20553 ( .A1(n17401), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17747) );
  NAND2_X1 U20554 ( .A1(n17504), .A2(n17384), .ZN(n17419) );
  INV_X1 U20555 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18549) );
  NOR2_X1 U20556 ( .A1(n17963), .A2(n18549), .ZN(n17737) );
  AOI221_X1 U20557 ( .B1(n17386), .B2(n20831), .C1(n18006), .C2(n20831), .A(
        n17385), .ZN(n17387) );
  AOI211_X1 U20558 ( .C1(n20819), .C2(n17419), .A(n17737), .B(n17387), .ZN(
        n17391) );
  NAND2_X1 U20559 ( .A1(n17730), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17741) );
  INV_X1 U20560 ( .A(n17741), .ZN(n17713) );
  OAI21_X1 U20561 ( .B1(n17388), .B2(n17713), .A(n17443), .ZN(n17402) );
  OAI221_X1 U20562 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17414), 
        .C1(n17401), .C2(n17399), .A(n17349), .ZN(n17389) );
  XNOR2_X1 U20563 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17389), .ZN(
        n17738) );
  AOI22_X1 U20564 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17402), .B1(
        n17537), .B2(n17738), .ZN(n17390) );
  OAI211_X1 U20565 ( .C1(n17405), .C2(n17747), .A(n17391), .B(n17390), .ZN(
        P3_U2810) );
  INV_X1 U20566 ( .A(n17408), .ZN(n17392) );
  INV_X1 U20567 ( .A(n17640), .ZN(n17524) );
  OAI21_X1 U20568 ( .B1(n17614), .B2(n17392), .A(n17524), .ZN(n17420) );
  OAI21_X1 U20569 ( .B1(n17393), .B2(n17644), .A(n17420), .ZN(n17413) );
  NAND2_X1 U20570 ( .A1(n17965), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17750) );
  INV_X1 U20571 ( .A(n17750), .ZN(n17398) );
  AND2_X1 U20572 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17396) );
  OAI211_X1 U20573 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17408), .B(n17407), .ZN(n17395) );
  OAI22_X1 U20574 ( .A1(n17396), .A2(n17395), .B1(n17394), .B2(n17504), .ZN(
        n17397) );
  AOI211_X1 U20575 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n17413), .A(
        n17398), .B(n17397), .ZN(n17404) );
  AOI21_X1 U20576 ( .B1(n17414), .B2(n17415), .A(n17399), .ZN(n17400) );
  XOR2_X1 U20577 ( .A(n17401), .B(n17400), .Z(n17748) );
  AOI22_X1 U20578 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17402), .B1(
        n17537), .B2(n17748), .ZN(n17403) );
  OAI211_X1 U20579 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17405), .A(
        n17404), .B(n17403), .ZN(P3_U2811) );
  NAND2_X1 U20580 ( .A1(n17759), .A2(n17406), .ZN(n17768) );
  NAND2_X1 U20581 ( .A1(n17965), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17766) );
  INV_X1 U20582 ( .A(n17766), .ZN(n17412) );
  NAND2_X1 U20583 ( .A1(n17408), .A2(n17407), .ZN(n17410) );
  OAI22_X1 U20584 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17410), .B1(
        n17409), .B2(n17504), .ZN(n17411) );
  AOI211_X1 U20585 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n17413), .A(
        n17412), .B(n17411), .ZN(n17418) );
  OAI21_X1 U20586 ( .B1(n17759), .B2(n17444), .A(n17443), .ZN(n17426) );
  AOI21_X1 U20587 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17431), .A(
        n17414), .ZN(n17416) );
  XOR2_X1 U20588 ( .A(n17416), .B(n17415), .Z(n17764) );
  AOI22_X1 U20589 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17426), .B1(
        n17537), .B2(n17764), .ZN(n17417) );
  OAI211_X1 U20590 ( .C1(n17444), .C2(n17768), .A(n17418), .B(n17417), .ZN(
        P3_U2812) );
  NAND2_X1 U20591 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17769), .ZN(
        n17775) );
  INV_X1 U20592 ( .A(n17419), .ZN(n17627) );
  NOR2_X1 U20593 ( .A1(n17963), .A2(n18544), .ZN(n17772) );
  AOI221_X1 U20594 ( .B1(n17422), .B2(n17421), .C1(n18006), .C2(n17421), .A(
        n17420), .ZN(n17423) );
  AOI211_X1 U20595 ( .C1(n17424), .C2(n17419), .A(n17772), .B(n17423), .ZN(
        n17428) );
  OAI21_X1 U20596 ( .B1(n9738), .B2(n17769), .A(n17425), .ZN(n17773) );
  AOI22_X1 U20597 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17426), .B1(
        n17537), .B2(n17773), .ZN(n17427) );
  OAI211_X1 U20598 ( .C1(n17444), .C2(n17775), .A(n17428), .B(n17427), .ZN(
        P3_U2813) );
  NOR2_X1 U20599 ( .A1(n17546), .A2(n17820), .ZN(n17529) );
  INV_X1 U20600 ( .A(n17529), .ZN(n17519) );
  OAI22_X1 U20601 ( .A1(n17431), .A2(n17430), .B1(n17519), .B2(n17429), .ZN(
        n17432) );
  XOR2_X1 U20602 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17432), .Z(
        n17783) );
  INV_X1 U20603 ( .A(n17433), .ZN(n17434) );
  AOI21_X1 U20604 ( .B1(n17541), .B2(n17434), .A(n17614), .ZN(n17464) );
  OAI21_X1 U20605 ( .B1(n17435), .B2(n17644), .A(n17464), .ZN(n17447) );
  AOI22_X1 U20606 ( .A1(n17965), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17447), .ZN(n17439) );
  INV_X1 U20607 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17437) );
  NOR3_X1 U20608 ( .A1(n17486), .A2(n17485), .A3(n17436), .ZN(n17449) );
  OAI221_X1 U20609 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C1(n17437), .C2(n17448), .A(
        n17449), .ZN(n17438) );
  OAI211_X1 U20610 ( .C1(n17504), .C2(n17440), .A(n17439), .B(n17438), .ZN(
        n17441) );
  AOI21_X1 U20611 ( .B1(n17537), .B2(n17783), .A(n17441), .ZN(n17442) );
  OAI221_X1 U20612 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17444), 
        .C1(n17786), .C2(n17443), .A(n17442), .ZN(P3_U2814) );
  NAND2_X1 U20613 ( .A1(n17843), .A2(n17481), .ZN(n17482) );
  AOI21_X1 U20614 ( .B1(n17459), .B2(n17830), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17801) );
  NAND2_X1 U20615 ( .A1(n17633), .A2(n17788), .ZN(n17458) );
  OAI22_X1 U20616 ( .A1(n17963), .A2(n18540), .B1(n17504), .B2(n17445), .ZN(
        n17446) );
  AOI221_X1 U20617 ( .B1(n17449), .B2(n17448), .C1(n17447), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17446), .ZN(n17457) );
  AND2_X1 U20618 ( .A1(n17825), .A2(n17459), .ZN(n17451) );
  AOI21_X1 U20619 ( .B1(n17478), .B2(n17451), .A(n17450), .ZN(n17452) );
  AOI221_X1 U20620 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17842), 
        .C1(n17546), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17452), .ZN(
        n17453) );
  XOR2_X1 U20621 ( .A(n17453), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Z(
        n17793) );
  NOR2_X1 U20622 ( .A1(n17790), .A2(n17454), .ZN(n17455) );
  OAI21_X1 U20623 ( .B1(n17778), .B2(n17820), .A(n17804), .ZN(n17791) );
  AOI22_X1 U20624 ( .A1(n17537), .A2(n17793), .B1(n17455), .B2(n17791), .ZN(
        n17456) );
  OAI211_X1 U20625 ( .C1(n17801), .C2(n17458), .A(n17457), .B(n17456), .ZN(
        P3_U2815) );
  NAND2_X1 U20626 ( .A1(n17459), .A2(n17830), .ZN(n17460) );
  OAI221_X1 U20627 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17830), .A(n17460), .ZN(
        n17819) );
  NAND2_X1 U20628 ( .A1(n17461), .A2(n18364), .ZN(n17523) );
  NOR2_X1 U20629 ( .A1(n17508), .A2(n17523), .ZN(n17512) );
  AOI21_X1 U20630 ( .B1(n17462), .B2(n17512), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17463) );
  OAI22_X1 U20631 ( .A1(n17627), .A2(n17465), .B1(n17464), .B2(n17463), .ZN(
        n17466) );
  AOI21_X1 U20632 ( .B1(n17965), .B2(P3_REIP_REG_14__SCAN_IN), .A(n17466), 
        .ZN(n17471) );
  NAND2_X1 U20633 ( .A1(n17845), .A2(n17481), .ZN(n17826) );
  NOR2_X1 U20634 ( .A1(n17820), .A2(n17778), .ZN(n17467) );
  AOI221_X1 U20635 ( .B1(n17483), .B2(n17811), .C1(n17826), .C2(n17811), .A(
        n17467), .ZN(n17815) );
  NAND2_X1 U20636 ( .A1(n17481), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17808) );
  OAI21_X1 U20637 ( .B1(n17519), .B2(n17808), .A(n17468), .ZN(n17469) );
  XOR2_X1 U20638 ( .A(n17469), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n17814) );
  AOI22_X1 U20639 ( .A1(n17552), .A2(n17815), .B1(n17537), .B2(n17814), .ZN(
        n17470) );
  OAI211_X1 U20640 ( .C1(n17648), .C2(n17819), .A(n17471), .B(n17470), .ZN(
        P3_U2816) );
  AOI22_X1 U20641 ( .A1(n17473), .A2(n17472), .B1(n17541), .B2(n17485), .ZN(
        n17474) );
  NAND2_X1 U20642 ( .A1(n17474), .A2(n17643), .ZN(n17493) );
  AOI22_X1 U20643 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17493), .B1(
        n17476), .B2(n17475), .ZN(n17491) );
  AOI22_X1 U20644 ( .A1(n17478), .A2(n17481), .B1(n17546), .B2(n17842), .ZN(
        n17479) );
  AOI21_X1 U20645 ( .B1(n17477), .B2(n17546), .A(n17479), .ZN(n17480) );
  XOR2_X1 U20646 ( .A(n17480), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n17824) );
  NAND2_X1 U20647 ( .A1(n17481), .A2(n17483), .ZN(n17835) );
  AOI22_X1 U20648 ( .A1(n17552), .A2(n17826), .B1(n17633), .B2(n17482), .ZN(
        n17497) );
  OAI22_X1 U20649 ( .A1(n17540), .A2(n17835), .B1(n17497), .B2(n17483), .ZN(
        n17484) );
  AOI21_X1 U20650 ( .B1(n17537), .B2(n17824), .A(n17484), .ZN(n17490) );
  NAND2_X1 U20651 ( .A1(n17965), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17489) );
  NOR2_X1 U20652 ( .A1(n17486), .A2(n17485), .ZN(n17495) );
  OAI211_X1 U20653 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17495), .B(n17487), .ZN(n17488) );
  NAND4_X1 U20654 ( .A1(n17491), .A2(n17490), .A3(n17489), .A4(n17488), .ZN(
        P3_U2817) );
  INV_X1 U20655 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17494) );
  NOR2_X1 U20656 ( .A1(n17963), .A2(n18534), .ZN(n17492) );
  AOI221_X1 U20657 ( .B1(n17495), .B2(n17494), .C1(n17493), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17492), .ZN(n17502) );
  INV_X1 U20658 ( .A(n17825), .ZN(n17837) );
  OAI21_X1 U20659 ( .B1(n17837), .B2(n17519), .A(n17477), .ZN(n17496) );
  XOR2_X1 U20660 ( .A(n17496), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n17836) );
  NOR2_X1 U20661 ( .A1(n17540), .A2(n17837), .ZN(n17499) );
  INV_X1 U20662 ( .A(n17497), .ZN(n17498) );
  MUX2_X1 U20663 ( .A(n17499), .B(n17498), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n17500) );
  AOI21_X1 U20664 ( .B1(n17537), .B2(n17836), .A(n17500), .ZN(n17501) );
  OAI211_X1 U20665 ( .C1(n17504), .C2(n17503), .A(n17502), .B(n17501), .ZN(
        P3_U2818) );
  INV_X1 U20666 ( .A(n17507), .ZN(n17849) );
  AOI21_X1 U20667 ( .B1(n17529), .B2(n17849), .A(n17505), .ZN(n17506) );
  XOR2_X1 U20668 ( .A(n17506), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n17857) );
  NOR2_X1 U20669 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17507), .ZN(
        n17855) );
  INV_X1 U20670 ( .A(n17540), .ZN(n17514) );
  INV_X1 U20671 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18532) );
  NOR2_X1 U20672 ( .A1(n17963), .A2(n18532), .ZN(n17854) );
  OAI21_X1 U20673 ( .B1(n17508), .B2(n17640), .A(n17523), .ZN(n17509) );
  INV_X1 U20674 ( .A(n17509), .ZN(n17511) );
  OAI22_X1 U20675 ( .A1(n17512), .A2(n17511), .B1(n17627), .B2(n17510), .ZN(
        n17513) );
  AOI211_X1 U20676 ( .C1(n17855), .C2(n17514), .A(n17854), .B(n17513), .ZN(
        n17516) );
  NOR2_X1 U20677 ( .A1(n17849), .A2(n17540), .ZN(n17522) );
  INV_X1 U20678 ( .A(n17843), .ZN(n17821) );
  AOI22_X1 U20679 ( .A1(n17820), .A2(n17552), .B1(n17633), .B2(n17821), .ZN(
        n17539) );
  INV_X1 U20680 ( .A(n17539), .ZN(n17521) );
  OAI21_X1 U20681 ( .B1(n17522), .B2(n17521), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17515) );
  OAI211_X1 U20682 ( .C1(n17857), .C2(n17549), .A(n17516), .B(n17515), .ZN(
        P3_U2819) );
  AOI22_X1 U20683 ( .A1(n17965), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17517), 
        .B2(n17419), .ZN(n17528) );
  OAI21_X1 U20684 ( .B1(n17859), .B2(n17519), .A(n17518), .ZN(n17520) );
  XOR2_X1 U20685 ( .A(n17520), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .Z(
        n17861) );
  AOI22_X1 U20686 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17521), .B1(
        n17537), .B2(n17861), .ZN(n17527) );
  OAI21_X1 U20687 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n17522), .ZN(n17526) );
  NOR3_X1 U20688 ( .A1(n20849), .A2(n17561), .A3(n18006), .ZN(n17544) );
  NAND2_X1 U20689 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17544), .ZN(
        n17533) );
  NOR2_X1 U20690 ( .A1(n17532), .A2(n17533), .ZN(n17531) );
  OAI211_X1 U20691 ( .C1(n17531), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n17524), .B(n17523), .ZN(n17525) );
  NAND4_X1 U20692 ( .A1(n17528), .A2(n17527), .A3(n17526), .A4(n17525), .ZN(
        P3_U2820) );
  NOR2_X1 U20693 ( .A1(n17529), .A2(n9748), .ZN(n17530) );
  XOR2_X1 U20694 ( .A(n17530), .B(n17859), .Z(n17871) );
  AOI211_X1 U20695 ( .C1(n17533), .C2(n17532), .A(n17640), .B(n17531), .ZN(
        n17536) );
  OAI22_X1 U20696 ( .A1(n17627), .A2(n17534), .B1(n17963), .B2(n18528), .ZN(
        n17535) );
  AOI211_X1 U20697 ( .C1(n17537), .C2(n17871), .A(n17536), .B(n17535), .ZN(
        n17538) );
  OAI221_X1 U20698 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17540), .C1(
        n17859), .C2(n17539), .A(n17538), .ZN(P3_U2821) );
  AOI21_X1 U20699 ( .B1(n17541), .B2(n17561), .A(n17614), .ZN(n17562) );
  OAI21_X1 U20700 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18006), .A(
        n17562), .ZN(n17542) );
  NOR2_X1 U20701 ( .A1(n17963), .A2(n18526), .ZN(n17889) );
  AOI221_X1 U20702 ( .B1(n17544), .B2(n17543), .C1(n17542), .C2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(n17889), .ZN(n17554) );
  INV_X1 U20703 ( .A(n17551), .ZN(n17886) );
  AOI21_X1 U20704 ( .B1(n17546), .B2(n17886), .A(n17545), .ZN(n17892) );
  OAI21_X1 U20705 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17548), .A(
        n17547), .ZN(n17884) );
  OAI22_X1 U20706 ( .A1(n17892), .A2(n17549), .B1(n17648), .B2(n17884), .ZN(
        n17550) );
  AOI21_X1 U20707 ( .B1(n17552), .B2(n17551), .A(n17550), .ZN(n17553) );
  OAI211_X1 U20708 ( .C1(n17627), .C2(n17555), .A(n17554), .B(n17553), .ZN(
        P3_U2822) );
  OAI21_X1 U20709 ( .B1(n17558), .B2(n17557), .A(n17556), .ZN(n17559) );
  XOR2_X1 U20710 ( .A(n17559), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n17900) );
  NAND2_X1 U20711 ( .A1(n18364), .A2(n20849), .ZN(n17560) );
  OAI22_X1 U20712 ( .A1(n17562), .A2(n20849), .B1(n17561), .B2(n17560), .ZN(
        n17563) );
  AOI21_X1 U20713 ( .B1(n17965), .B2(P3_REIP_REG_7__SCAN_IN), .A(n17563), .ZN(
        n17568) );
  AOI21_X1 U20714 ( .B1(n17565), .B2(n17894), .A(n17564), .ZN(n17897) );
  AOI22_X1 U20715 ( .A1(n17636), .A2(n17897), .B1(n17566), .B2(n17419), .ZN(
        n17567) );
  OAI211_X1 U20716 ( .C1(n17648), .C2(n17900), .A(n17568), .B(n17567), .ZN(
        P3_U2823) );
  NAND2_X1 U20717 ( .A1(n17572), .A2(n18364), .ZN(n17579) );
  AOI21_X1 U20718 ( .B1(n17571), .B2(n17570), .A(n17569), .ZN(n17904) );
  AOI22_X1 U20719 ( .A1(n17636), .A2(n17904), .B1(n17965), .B2(
        P3_REIP_REG_6__SCAN_IN), .ZN(n17578) );
  AOI21_X1 U20720 ( .B1(n18364), .B2(n17572), .A(n17640), .ZN(n17591) );
  OAI21_X1 U20721 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17574), .A(
        n17573), .ZN(n17907) );
  OAI22_X1 U20722 ( .A1(n17627), .A2(n17575), .B1(n17648), .B2(n17907), .ZN(
        n17576) );
  AOI21_X1 U20723 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17591), .A(
        n17576), .ZN(n17577) );
  OAI211_X1 U20724 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n17579), .A(
        n17578), .B(n17577), .ZN(P3_U2824) );
  OAI21_X1 U20725 ( .B1(n17582), .B2(n17581), .A(n17580), .ZN(n17583) );
  XOR2_X1 U20726 ( .A(n17583), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n17913) );
  OAI21_X1 U20727 ( .B1(n17585), .B2(n9751), .A(n17584), .ZN(n17586) );
  XOR2_X1 U20728 ( .A(n17586), .B(n10917), .Z(n17910) );
  AOI22_X1 U20729 ( .A1(n17636), .A2(n17910), .B1(n17965), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17593) );
  OAI21_X1 U20730 ( .B1(n17614), .B2(n17588), .A(n17587), .ZN(n17590) );
  AOI22_X1 U20731 ( .A1(n17591), .A2(n17590), .B1(n17589), .B2(n17419), .ZN(
        n17592) );
  OAI211_X1 U20732 ( .C1(n17648), .C2(n17913), .A(n17593), .B(n17592), .ZN(
        P3_U2825) );
  AOI21_X1 U20733 ( .B1(n17596), .B2(n17595), .A(n17594), .ZN(n17924) );
  INV_X1 U20734 ( .A(n17597), .ZN(n17598) );
  OAI22_X1 U20735 ( .A1(n17924), .A2(n17648), .B1(n18006), .B2(n17598), .ZN(
        n17599) );
  AOI21_X1 U20736 ( .B1(n17965), .B2(P3_REIP_REG_4__SCAN_IN), .A(n17599), .ZN(
        n17606) );
  AOI21_X1 U20737 ( .B1(n17602), .B2(n17601), .A(n17600), .ZN(n17922) );
  OAI21_X1 U20738 ( .B1(n17604), .B2(n17603), .A(n17643), .ZN(n17616) );
  AOI22_X1 U20739 ( .A1(n17636), .A2(n17922), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17616), .ZN(n17605) );
  OAI211_X1 U20740 ( .C1(n17627), .C2(n17607), .A(n17606), .B(n17605), .ZN(
        P3_U2826) );
  OAI21_X1 U20741 ( .B1(n17610), .B2(n17609), .A(n17608), .ZN(n17933) );
  AOI21_X1 U20742 ( .B1(n17926), .B2(n17612), .A(n17611), .ZN(n17928) );
  AOI22_X1 U20743 ( .A1(n17636), .A2(n17928), .B1(n17965), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17619) );
  OAI21_X1 U20744 ( .B1(n17614), .B2(n17631), .A(n17613), .ZN(n17615) );
  AOI22_X1 U20745 ( .A1(n17617), .A2(n17419), .B1(n17616), .B2(n17615), .ZN(
        n17618) );
  OAI211_X1 U20746 ( .C1(n17648), .C2(n17933), .A(n17619), .B(n17618), .ZN(
        P3_U2827) );
  AOI21_X1 U20747 ( .B1(n17622), .B2(n17621), .A(n17620), .ZN(n17940) );
  NAND2_X1 U20748 ( .A1(n17965), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n17945) );
  INV_X1 U20749 ( .A(n17945), .ZN(n17629) );
  OAI21_X1 U20750 ( .B1(n17625), .B2(n17624), .A(n17623), .ZN(n17947) );
  OAI22_X1 U20751 ( .A1(n17627), .A2(n17626), .B1(n17648), .B2(n17947), .ZN(
        n17628) );
  AOI211_X1 U20752 ( .C1(n17636), .C2(n17940), .A(n17629), .B(n17628), .ZN(
        n17630) );
  OAI221_X1 U20753 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18006), .C1(
        n17631), .C2(n17643), .A(n17630), .ZN(P3_U2828) );
  NOR2_X1 U20754 ( .A1(n17642), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17632) );
  XNOR2_X1 U20755 ( .A(n17632), .B(n17635), .ZN(n17950) );
  AOI22_X1 U20756 ( .A1(n17633), .A2(n17950), .B1(n17965), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17638) );
  AOI21_X1 U20757 ( .B1(n17641), .B2(n17635), .A(n17634), .ZN(n17948) );
  AOI22_X1 U20758 ( .A1(n17636), .A2(n17948), .B1(n17639), .B2(n17419), .ZN(
        n17637) );
  OAI211_X1 U20759 ( .C1(n17640), .C2(n17639), .A(n17638), .B(n17637), .ZN(
        P3_U2829) );
  OAI21_X1 U20760 ( .B1(n17642), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17641), .ZN(n17968) );
  INV_X1 U20761 ( .A(n17968), .ZN(n17970) );
  NAND3_X1 U20762 ( .A1(n18605), .A2(n17644), .A3(n17643), .ZN(n17645) );
  AOI22_X1 U20763 ( .A1(n17965), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17645), .ZN(n17646) );
  OAI221_X1 U20764 ( .B1(n17970), .B2(n17648), .C1(n17968), .C2(n17647), .A(
        n17646), .ZN(P3_U2830) );
  NOR2_X1 U20765 ( .A1(n17687), .A2(n17649), .ZN(n17660) );
  NAND2_X1 U20766 ( .A1(n18453), .A2(n18451), .ZN(n17934) );
  INV_X1 U20767 ( .A(n17934), .ZN(n17763) );
  OAI21_X1 U20768 ( .B1(n17726), .B2(n18438), .A(n17650), .ZN(n17720) );
  NAND2_X1 U20769 ( .A1(n17651), .A2(n17720), .ZN(n17652) );
  OAI21_X1 U20770 ( .B1(n17711), .B2(n17652), .A(n17934), .ZN(n17689) );
  OAI21_X1 U20771 ( .B1(n17673), .B2(n17763), .A(n17689), .ZN(n17675) );
  NAND2_X1 U20772 ( .A1(n17653), .A2(n17934), .ZN(n17655) );
  OAI211_X1 U20773 ( .C1(n17656), .C2(n17844), .A(n17655), .B(n17654), .ZN(
        n17657) );
  AOI211_X1 U20774 ( .C1(n17789), .C2(n17658), .A(n17675), .B(n17657), .ZN(
        n17665) );
  INV_X1 U20775 ( .A(n17665), .ZN(n17659) );
  MUX2_X1 U20776 ( .A(n17660), .B(n17659), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n17661) );
  AOI22_X1 U20777 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17954), .B1(
        n17961), .B2(n17661), .ZN(n17663) );
  NAND2_X1 U20778 ( .A1(n17965), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17662) );
  OAI211_X1 U20779 ( .C1(n17664), .C2(n17891), .A(n17663), .B(n17662), .ZN(
        P3_U2835) );
  AOI221_X1 U20780 ( .B1(n17667), .B2(n17666), .C1(n17703), .C2(n17666), .A(
        n17665), .ZN(n17668) );
  AOI22_X1 U20781 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17954), .B1(
        n17961), .B2(n17668), .ZN(n17670) );
  NAND2_X1 U20782 ( .A1(n17965), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17669) );
  OAI211_X1 U20783 ( .C1(n17671), .C2(n17891), .A(n17670), .B(n17669), .ZN(
        P3_U2836) );
  NOR2_X1 U20784 ( .A1(n17672), .A2(n17757), .ZN(n17693) );
  OAI221_X1 U20785 ( .B1(n18427), .B2(n17673), .C1(n18427), .C2(n17693), .A(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17674) );
  OAI21_X1 U20786 ( .B1(n17675), .B2(n17674), .A(n17961), .ZN(n17676) );
  AOI221_X1 U20787 ( .B1(n17679), .B2(n17678), .C1(n17677), .C2(n17678), .A(
        n17676), .ZN(n17680) );
  AOI211_X1 U20788 ( .C1(n17954), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17681), .B(n17680), .ZN(n17685) );
  AOI22_X1 U20789 ( .A1(n17951), .A2(n17683), .B1(n17816), .B2(n17682), .ZN(
        n17684) );
  OAI211_X1 U20790 ( .C1(n17891), .C2(n17686), .A(n17685), .B(n17684), .ZN(
        P3_U2837) );
  NOR2_X1 U20791 ( .A1(n17687), .A2(n17952), .ZN(n17727) );
  INV_X1 U20792 ( .A(n17688), .ZN(n17692) );
  OAI211_X1 U20793 ( .C1(n17690), .C2(n17844), .A(n17689), .B(n17925), .ZN(
        n17691) );
  AOI21_X1 U20794 ( .B1(n17789), .B2(n17692), .A(n17691), .ZN(n17696) );
  OAI211_X1 U20795 ( .C1(n17693), .C2(n18427), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n17696), .ZN(n17694) );
  NAND2_X1 U20796 ( .A1(n17963), .A2(n17694), .ZN(n17708) );
  AOI211_X1 U20797 ( .C1(n17880), .C2(n17696), .A(n17695), .B(n17708), .ZN(
        n17697) );
  AOI211_X1 U20798 ( .C1(n17699), .C2(n17727), .A(n17698), .B(n17697), .ZN(
        n17700) );
  OAI21_X1 U20799 ( .B1(n17701), .B2(n17891), .A(n17700), .ZN(P3_U2838) );
  OAI21_X1 U20800 ( .B1(n17703), .B2(n17954), .A(n17702), .ZN(n17704) );
  INV_X1 U20801 ( .A(n17704), .ZN(n17709) );
  AOI21_X1 U20802 ( .B1(n17706), .B2(n17872), .A(n17705), .ZN(n17707) );
  OAI21_X1 U20803 ( .B1(n17709), .B2(n17708), .A(n17707), .ZN(P3_U2839) );
  AOI22_X1 U20804 ( .A1(n17965), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n17872), 
        .B2(n17710), .ZN(n17725) );
  NOR2_X1 U20805 ( .A1(n17789), .A2(n17827), .ZN(n17848) );
  INV_X1 U20806 ( .A(n17848), .ZN(n17740) );
  INV_X1 U20807 ( .A(n17711), .ZN(n17756) );
  AOI22_X1 U20808 ( .A1(n17789), .A2(n17788), .B1(n17827), .B2(n17712), .ZN(
        n17760) );
  OAI221_X1 U20809 ( .B1(n18453), .B2(n17756), .C1(n18453), .C2(n17713), .A(
        n17760), .ZN(n17714) );
  AOI221_X1 U20810 ( .B1(n17715), .B2(n18449), .C1(n17757), .C2(n18449), .A(
        n17714), .ZN(n17743) );
  OAI21_X1 U20811 ( .B1(n18453), .B2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n17743), .ZN(n17716) );
  AOI21_X1 U20812 ( .B1(n17717), .B2(n17740), .A(n17716), .ZN(n17731) );
  AOI22_X1 U20813 ( .A1(n18449), .A2(n17719), .B1(n9768), .B2(n17718), .ZN(
        n17721) );
  NAND3_X1 U20814 ( .A1(n17731), .A2(n17721), .A3(n17720), .ZN(n17722) );
  OAI211_X1 U20815 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17723), .A(
        n17961), .B(n17722), .ZN(n17724) );
  OAI211_X1 U20816 ( .C1(n17925), .C2(n17726), .A(n17725), .B(n17724), .ZN(
        P3_U2840) );
  NAND2_X1 U20817 ( .A1(n17730), .A2(n17727), .ZN(n17752) );
  AOI21_X1 U20818 ( .B1(n17872), .B2(n17729), .A(n17728), .ZN(n17735) );
  OAI221_X1 U20819 ( .B1(n18451), .B2(n17730), .C1(n18451), .C2(n17780), .A(
        n17961), .ZN(n17739) );
  NOR2_X1 U20820 ( .A1(n18449), .A2(n18438), .ZN(n17953) );
  OAI21_X1 U20821 ( .B1(n17732), .B2(n17953), .A(n17731), .ZN(n17733) );
  OAI211_X1 U20822 ( .C1(n17739), .C2(n17733), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17963), .ZN(n17734) );
  OAI211_X1 U20823 ( .C1(n17736), .C2(n17752), .A(n17735), .B(n17734), .ZN(
        P3_U2841) );
  AOI21_X1 U20824 ( .B1(n17738), .B2(n17872), .A(n17737), .ZN(n17746) );
  AOI21_X1 U20825 ( .B1(n17741), .B2(n17740), .A(n17739), .ZN(n17742) );
  AOI21_X1 U20826 ( .B1(n17743), .B2(n17742), .A(n11114), .ZN(n17749) );
  NOR3_X1 U20827 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17953), .A3(
        n18646), .ZN(n17744) );
  OAI21_X1 U20828 ( .B1(n17749), .B2(n17744), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17745) );
  OAI211_X1 U20829 ( .C1(n17752), .C2(n17747), .A(n17746), .B(n17745), .ZN(
        P3_U2842) );
  AOI22_X1 U20830 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17749), .B1(
        n17872), .B2(n17748), .ZN(n17751) );
  OAI211_X1 U20831 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17752), .A(
        n17751), .B(n17750), .ZN(P3_U2843) );
  OAI22_X1 U20832 ( .A1(n17915), .A2(n18427), .B1(n17937), .B2(n17914), .ZN(
        n17930) );
  NAND2_X1 U20833 ( .A1(n17753), .A2(n17930), .ZN(n17893) );
  NOR2_X1 U20834 ( .A1(n17952), .A2(n17893), .ZN(n17903) );
  NAND3_X1 U20835 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n17903), .ZN(n17882) );
  NOR2_X1 U20836 ( .A1(n17881), .A2(n17882), .ZN(n17823) );
  AOI22_X1 U20837 ( .A1(n17755), .A2(n17823), .B1(n17961), .B2(n17754), .ZN(
        n17787) );
  NAND2_X1 U20838 ( .A1(n18438), .A2(n17960), .ZN(n17942) );
  NAND3_X1 U20839 ( .A1(n17756), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n17942), .ZN(n17762) );
  NAND2_X1 U20840 ( .A1(n18449), .A2(n17757), .ZN(n17758) );
  AOI22_X1 U20841 ( .A1(n17759), .A2(n17758), .B1(n17848), .B2(n18427), .ZN(
        n17761) );
  NAND2_X1 U20842 ( .A1(n17961), .A2(n17760), .ZN(n17782) );
  AOI211_X1 U20843 ( .C1(n17934), .C2(n17762), .A(n17761), .B(n17782), .ZN(
        n17770) );
  AOI221_X1 U20844 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17770), 
        .C1(n17763), .C2(n17770), .A(n17965), .ZN(n17765) );
  AOI22_X1 U20845 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17765), .B1(
        n17872), .B2(n17764), .ZN(n17767) );
  OAI211_X1 U20846 ( .C1(n17787), .C2(n17768), .A(n17767), .B(n17766), .ZN(
        P3_U2844) );
  NOR3_X1 U20847 ( .A1(n17965), .A2(n17770), .A3(n17769), .ZN(n17771) );
  AOI211_X1 U20848 ( .C1(n17872), .C2(n17773), .A(n17772), .B(n17771), .ZN(
        n17774) );
  OAI21_X1 U20849 ( .B1(n17787), .B2(n17775), .A(n17774), .ZN(P3_U2845) );
  OAI22_X1 U20850 ( .A1(n18453), .A2(n17777), .B1(n17776), .B2(n18427), .ZN(
        n17867) );
  AOI21_X1 U20851 ( .B1(n9768), .B2(n17778), .A(n17867), .ZN(n17779) );
  OAI211_X1 U20852 ( .C1(n17780), .C2(n18451), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17779), .ZN(n17797) );
  OAI221_X1 U20853 ( .B1(n17782), .B2(n17781), .C1(n17782), .C2(n17797), .A(
        n17963), .ZN(n17785) );
  AOI22_X1 U20854 ( .A1(n17965), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n17872), 
        .B2(n17783), .ZN(n17784) );
  OAI221_X1 U20855 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17787), 
        .C1(n17786), .C2(n17785), .A(n17784), .ZN(P3_U2846) );
  NAND2_X1 U20856 ( .A1(n17789), .A2(n17788), .ZN(n17800) );
  NOR2_X1 U20857 ( .A1(n17790), .A2(n17844), .ZN(n17792) );
  AOI22_X1 U20858 ( .A1(n17794), .A2(n17793), .B1(n17792), .B2(n17791), .ZN(
        n17799) );
  NOR3_X1 U20859 ( .A1(n17795), .A2(n17893), .A3(n17808), .ZN(n17805) );
  OAI211_X1 U20860 ( .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n17805), .A(
        n17797), .B(n17796), .ZN(n17798) );
  OAI211_X1 U20861 ( .C1(n17801), .C2(n17800), .A(n17799), .B(n17798), .ZN(
        n17802) );
  AOI22_X1 U20862 ( .A1(n17965), .A2(P3_REIP_REG_15__SCAN_IN), .B1(n17961), 
        .B2(n17802), .ZN(n17803) );
  OAI21_X1 U20863 ( .B1(n17804), .B2(n17925), .A(n17803), .ZN(P3_U2847) );
  INV_X1 U20864 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18538) );
  NOR2_X1 U20865 ( .A1(n17963), .A2(n18538), .ZN(n17813) );
  INV_X1 U20866 ( .A(n17805), .ZN(n17810) );
  OAI21_X1 U20867 ( .B1(n17806), .B2(n17866), .A(n18438), .ZN(n17828) );
  OAI211_X1 U20868 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n17953), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17828), .ZN(n17807) );
  AOI211_X1 U20869 ( .C1(n9768), .C2(n17808), .A(n17867), .B(n17807), .ZN(
        n17809) );
  AOI211_X1 U20870 ( .C1(n17811), .C2(n17810), .A(n17809), .B(n17952), .ZN(
        n17812) );
  AOI211_X1 U20871 ( .C1(n17954), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17813), .B(n17812), .ZN(n17818) );
  AOI22_X1 U20872 ( .A1(n17816), .A2(n17815), .B1(n17872), .B2(n17814), .ZN(
        n17817) );
  OAI211_X1 U20873 ( .C1(n17969), .C2(n17819), .A(n17818), .B(n17817), .ZN(
        P3_U2848) );
  OAI22_X1 U20874 ( .A1(n17821), .A2(n17969), .B1(n17820), .B2(n17885), .ZN(
        n17822) );
  NOR2_X1 U20875 ( .A1(n17823), .A2(n17822), .ZN(n17876) );
  AOI22_X1 U20876 ( .A1(n17965), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n17872), 
        .B2(n17824), .ZN(n17834) );
  NOR2_X1 U20877 ( .A1(n17831), .A2(n17825), .ZN(n17850) );
  AOI211_X1 U20878 ( .C1(n17827), .C2(n17826), .A(n17850), .B(n17867), .ZN(
        n17829) );
  OAI211_X1 U20879 ( .C1(n17830), .C2(n18426), .A(n17829), .B(n17828), .ZN(
        n17839) );
  OAI21_X1 U20880 ( .B1(n17831), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n17961), .ZN(n17832) );
  OAI211_X1 U20881 ( .C1(n17839), .C2(n17832), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17963), .ZN(n17833) );
  OAI211_X1 U20882 ( .C1(n17876), .C2(n17835), .A(n17834), .B(n17833), .ZN(
        P3_U2849) );
  AOI22_X1 U20883 ( .A1(n17965), .A2(P3_REIP_REG_12__SCAN_IN), .B1(n17872), 
        .B2(n17836), .ZN(n17841) );
  OAI22_X1 U20884 ( .A1(n17876), .A2(n17837), .B1(n17842), .B2(n17952), .ZN(
        n17838) );
  OAI21_X1 U20885 ( .B1(n17839), .B2(n17842), .A(n17838), .ZN(n17840) );
  OAI211_X1 U20886 ( .C1(n17925), .C2(n17842), .A(n17841), .B(n17840), .ZN(
        P3_U2850) );
  INV_X1 U20887 ( .A(n17876), .ZN(n17858) );
  INV_X1 U20888 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17864) );
  OAI22_X1 U20889 ( .A1(n17845), .A2(n17844), .B1(n18426), .B2(n17843), .ZN(
        n17846) );
  NOR2_X1 U20890 ( .A1(n17952), .A2(n17846), .ZN(n17869) );
  OAI22_X1 U20891 ( .A1(n18438), .A2(n17867), .B1(n17859), .B2(n17866), .ZN(
        n17847) );
  OAI211_X1 U20892 ( .C1(n17849), .C2(n17848), .A(n17869), .B(n17847), .ZN(
        n17860) );
  AOI211_X1 U20893 ( .C1(n18438), .C2(n17864), .A(n17850), .B(n17860), .ZN(
        n17852) );
  NOR3_X1 U20894 ( .A1(n17965), .A2(n17852), .A3(n17851), .ZN(n17853) );
  AOI211_X1 U20895 ( .C1(n17855), .C2(n17858), .A(n17854), .B(n17853), .ZN(
        n17856) );
  OAI21_X1 U20896 ( .B1(n17857), .B2(n17891), .A(n17856), .ZN(P3_U2851) );
  NAND2_X1 U20897 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17858), .ZN(
        n17865) );
  OAI221_X1 U20898 ( .B1(n17860), .B2(n9768), .C1(n17860), .C2(n17859), .A(
        n17963), .ZN(n17863) );
  AOI22_X1 U20899 ( .A1(n17965), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17872), 
        .B2(n17861), .ZN(n17862) );
  OAI221_X1 U20900 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n17865), 
        .C1(n17864), .C2(n17863), .A(n17862), .ZN(P3_U2852) );
  INV_X1 U20901 ( .A(n17866), .ZN(n17870) );
  NOR2_X1 U20902 ( .A1(n18438), .A2(n17867), .ZN(n17868) );
  AOI221_X1 U20903 ( .B1(n17870), .B2(n17869), .C1(n17868), .C2(n17869), .A(
        n17965), .ZN(n17873) );
  AOI22_X1 U20904 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17873), .B1(
        n17872), .B2(n17871), .ZN(n17875) );
  NAND2_X1 U20905 ( .A1(n17965), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n17874) );
  OAI211_X1 U20906 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n17876), .A(
        n17875), .B(n17874), .ZN(P3_U2853) );
  AOI22_X1 U20907 ( .A1(n18449), .A2(n17878), .B1(n17934), .B2(n17877), .ZN(
        n17879) );
  AND2_X1 U20908 ( .A1(n17879), .A2(n17942), .ZN(n17901) );
  OAI211_X1 U20909 ( .C1(n17880), .C2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n17901), .ZN(n17895) );
  AOI21_X1 U20910 ( .B1(n17955), .B2(n17895), .A(n17954), .ZN(n17883) );
  AOI22_X1 U20911 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17883), .B1(
        n17882), .B2(n17881), .ZN(n17888) );
  OAI22_X1 U20912 ( .A1(n17886), .A2(n17885), .B1(n17969), .B2(n17884), .ZN(
        n17887) );
  NOR3_X1 U20913 ( .A1(n17889), .A2(n17888), .A3(n17887), .ZN(n17890) );
  OAI21_X1 U20914 ( .B1(n17892), .B2(n17891), .A(n17890), .ZN(P3_U2854) );
  AOI22_X1 U20915 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17954), .B1(
        n17965), .B2(P3_REIP_REG_7__SCAN_IN), .ZN(n17899) );
  AOI221_X1 U20916 ( .B1(n17902), .B2(n17894), .C1(n17893), .C2(n17894), .A(
        n17952), .ZN(n17896) );
  AOI22_X1 U20917 ( .A1(n17949), .A2(n17897), .B1(n17896), .B2(n17895), .ZN(
        n17898) );
  OAI211_X1 U20918 ( .C1(n17969), .C2(n17900), .A(n17899), .B(n17898), .ZN(
        P3_U2855) );
  OAI21_X1 U20919 ( .B1(n17901), .B2(n17952), .A(n17925), .ZN(n17908) );
  AOI22_X1 U20920 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17908), .B1(
        n17965), .B2(P3_REIP_REG_6__SCAN_IN), .ZN(n17906) );
  AOI22_X1 U20921 ( .A1(n17904), .A2(n17949), .B1(n17903), .B2(n17902), .ZN(
        n17905) );
  OAI211_X1 U20922 ( .C1(n17969), .C2(n17907), .A(n17906), .B(n17905), .ZN(
        P3_U2856) );
  AOI22_X1 U20923 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17908), .B1(
        n17965), .B2(P3_REIP_REG_5__SCAN_IN), .ZN(n17912) );
  NAND3_X1 U20924 ( .A1(n17961), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n17930), .ZN(n17918) );
  NOR3_X1 U20925 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17917), .A3(
        n17918), .ZN(n17909) );
  AOI21_X1 U20926 ( .B1(n17910), .B2(n17949), .A(n17909), .ZN(n17911) );
  OAI211_X1 U20927 ( .C1(n17969), .C2(n17913), .A(n17912), .B(n17911), .ZN(
        P3_U2857) );
  NOR2_X1 U20928 ( .A1(n17963), .A2(n18518), .ZN(n17921) );
  AOI22_X1 U20929 ( .A1(n18449), .A2(n17915), .B1(n17934), .B2(n17914), .ZN(
        n17916) );
  NAND3_X1 U20930 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17916), .A3(
        n17942), .ZN(n17929) );
  AOI21_X1 U20931 ( .B1(n17955), .B2(n17929), .A(n17954), .ZN(n17919) );
  AOI22_X1 U20932 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n17919), .B1(
        n17918), .B2(n17917), .ZN(n17920) );
  AOI211_X1 U20933 ( .C1(n17922), .C2(n17949), .A(n17921), .B(n17920), .ZN(
        n17923) );
  OAI21_X1 U20934 ( .B1(n17924), .B2(n17969), .A(n17923), .ZN(P3_U2858) );
  OAI22_X1 U20935 ( .A1(n17926), .A2(n17925), .B1(n17963), .B2(n18516), .ZN(
        n17927) );
  AOI21_X1 U20936 ( .B1(n17949), .B2(n17928), .A(n17927), .ZN(n17932) );
  OAI211_X1 U20937 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n17930), .A(
        n17961), .B(n17929), .ZN(n17931) );
  OAI211_X1 U20938 ( .C1(n17933), .C2(n17969), .A(n17932), .B(n17931), .ZN(
        P3_U2859) );
  NOR2_X1 U20939 ( .A1(n10903), .A2(n17960), .ZN(n17935) );
  AOI22_X1 U20940 ( .A1(n18449), .A2(n17935), .B1(n10903), .B2(n17934), .ZN(
        n17943) );
  NOR2_X1 U20941 ( .A1(n18427), .A2(n17936), .ZN(n17939) );
  NOR3_X1 U20942 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10903), .A3(
        n17937), .ZN(n17938) );
  AOI211_X1 U20943 ( .C1(n17940), .C2(n18422), .A(n17939), .B(n17938), .ZN(
        n17941) );
  OAI221_X1 U20944 ( .B1(n10906), .B2(n17943), .C1(n10906), .C2(n17942), .A(
        n17941), .ZN(n17944) );
  AOI22_X1 U20945 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n17954), .B1(
        n17961), .B2(n17944), .ZN(n17946) );
  OAI211_X1 U20946 ( .C1(n17947), .C2(n17969), .A(n17946), .B(n17945), .ZN(
        P3_U2860) );
  AOI22_X1 U20947 ( .A1(n17951), .A2(n17950), .B1(n17949), .B2(n17948), .ZN(
        n17959) );
  NAND2_X1 U20948 ( .A1(n17965), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n17958) );
  NOR3_X1 U20949 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17953), .A3(
        n17952), .ZN(n17962) );
  OAI21_X1 U20950 ( .B1(n17954), .B2(n17962), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17957) );
  OAI211_X1 U20951 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18437), .A(
        n17955), .B(n10903), .ZN(n17956) );
  NAND4_X1 U20952 ( .A1(n17959), .A2(n17958), .A3(n17957), .A4(n17956), .ZN(
        P3_U2861) );
  AOI21_X1 U20953 ( .B1(n18453), .B2(n17961), .A(n17960), .ZN(n17964) );
  AOI221_X1 U20954 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n17965), .C1(n17964), 
        .C2(n17963), .A(n17962), .ZN(n17966) );
  OAI221_X1 U20955 ( .B1(n17970), .B2(n17969), .C1(n17968), .C2(n17967), .A(
        n17966), .ZN(P3_U2862) );
  AOI211_X1 U20956 ( .C1(n17972), .C2(n17971), .A(n18646), .B(n18605), .ZN(
        n18477) );
  OAI21_X1 U20957 ( .B1(n18477), .B2(n18028), .A(n17982), .ZN(n17973) );
  OAI221_X1 U20958 ( .B1(n18272), .B2(n18625), .C1(n18272), .C2(n17982), .A(
        n17973), .ZN(P3_U2863) );
  AOI221_X1 U20959 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18457), .C1(n17975), 
        .C2(n18457), .A(n17974), .ZN(n17981) );
  NOR2_X1 U20960 ( .A1(n17976), .A2(n18457), .ZN(n17978) );
  OAI21_X1 U20961 ( .B1(n17978), .B2(n17977), .A(n17982), .ZN(n17979) );
  AOI22_X1 U20962 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17981), .B1(
        n17979), .B2(n18463), .ZN(P3_U2865) );
  INV_X1 U20963 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18466) );
  NOR2_X1 U20964 ( .A1(n18466), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18201) );
  NOR2_X1 U20965 ( .A1(n18463), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18156) );
  NOR2_X1 U20966 ( .A1(n18201), .A2(n18156), .ZN(n17980) );
  OAI22_X1 U20967 ( .A1(n17981), .A2(n18466), .B1(n17980), .B2(n17979), .ZN(
        P3_U2866) );
  NOR2_X1 U20968 ( .A1(n18467), .A2(n17982), .ZN(P3_U2867) );
  NAND2_X1 U20969 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18364), .ZN(n18330) );
  NOR2_X1 U20970 ( .A1(n18463), .A2(n18466), .ZN(n18301) );
  NAND2_X1 U20971 ( .A1(n18301), .A2(n18457), .ZN(n18299) );
  NOR2_X2 U20972 ( .A1(n18272), .A2(n18299), .ZN(n18410) );
  INV_X1 U20973 ( .A(n18410), .ZN(n18406) );
  NAND2_X1 U20974 ( .A1(n18364), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18368) );
  INV_X1 U20975 ( .A(n18368), .ZN(n18323) );
  NAND2_X1 U20976 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18301), .ZN(
        n18357) );
  NOR2_X2 U20977 ( .A1(n18357), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18352) );
  NOR2_X2 U20978 ( .A1(n18178), .A2(n17983), .ZN(n18359) );
  INV_X1 U20979 ( .A(n18357), .ZN(n18362) );
  NAND2_X1 U20980 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18362), .ZN(
        n18399) );
  INV_X1 U20981 ( .A(n18399), .ZN(n18413) );
  NAND2_X1 U20982 ( .A1(n18457), .A2(n18272), .ZN(n18459) );
  NAND2_X1 U20983 ( .A1(n18463), .A2(n18466), .ZN(n18047) );
  NOR2_X2 U20984 ( .A1(n18459), .A2(n18047), .ZN(n18086) );
  NOR2_X1 U20985 ( .A1(n18413), .A2(n18086), .ZN(n18048) );
  NOR2_X1 U20986 ( .A1(n18358), .A2(n18048), .ZN(n18022) );
  AOI22_X1 U20987 ( .A1(n18323), .A2(n18352), .B1(n18359), .B2(n18022), .ZN(
        n17990) );
  INV_X1 U20988 ( .A(n18352), .ZN(n18343) );
  NAND2_X1 U20989 ( .A1(n18343), .A2(n18406), .ZN(n17985) );
  AOI211_X1 U20990 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18048), .B(n18178), .ZN(
        n17984) );
  AOI21_X1 U20991 ( .B1(n18364), .B2(n17985), .A(n17984), .ZN(n18025) );
  NAND2_X1 U20992 ( .A1(n17987), .A2(n17986), .ZN(n18023) );
  INV_X1 U20993 ( .A(n18023), .ZN(n18010) );
  NAND2_X1 U20994 ( .A1(n17988), .A2(n18010), .ZN(n18231) );
  INV_X1 U20995 ( .A(n18231), .ZN(n18365) );
  AOI22_X1 U20996 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18025), .B1(
        n18086), .B2(n18365), .ZN(n17989) );
  OAI211_X1 U20997 ( .C1(n18330), .C2(n18406), .A(n17990), .B(n17989), .ZN(
        P3_U2868) );
  NAND2_X1 U20998 ( .A1(n18364), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18281) );
  NOR2_X2 U20999 ( .A1(n18178), .A2(n20751), .ZN(n18369) );
  NAND2_X1 U21000 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18364), .ZN(n18374) );
  INV_X1 U21001 ( .A(n18374), .ZN(n18278) );
  AOI22_X1 U21002 ( .A1(n18369), .A2(n18022), .B1(n18278), .B2(n18410), .ZN(
        n17993) );
  NAND2_X1 U21003 ( .A1(n17991), .A2(n18010), .ZN(n18209) );
  INV_X1 U21004 ( .A(n18209), .ZN(n18371) );
  AOI22_X1 U21005 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18025), .B1(
        n18086), .B2(n18371), .ZN(n17992) );
  OAI211_X1 U21006 ( .C1(n18281), .C2(n18343), .A(n17993), .B(n17992), .ZN(
        P3_U2869) );
  NAND2_X1 U21007 ( .A1(n18364), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18380) );
  NOR2_X2 U21008 ( .A1(n18178), .A2(n17994), .ZN(n18376) );
  AND2_X1 U21009 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18364), .ZN(n18375) );
  AOI22_X1 U21010 ( .A1(n18376), .A2(n18022), .B1(n18375), .B2(n18410), .ZN(
        n17997) );
  NAND2_X1 U21011 ( .A1(n17995), .A2(n18010), .ZN(n18285) );
  INV_X1 U21012 ( .A(n18285), .ZN(n18377) );
  AOI22_X1 U21013 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18025), .B1(
        n18086), .B2(n18377), .ZN(n17996) );
  OAI211_X1 U21014 ( .C1(n18380), .C2(n18343), .A(n17997), .B(n17996), .ZN(
        P3_U2870) );
  INV_X1 U21015 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n17998) );
  NOR2_X1 U21016 ( .A1(n18006), .A2(n17998), .ZN(n18382) );
  INV_X1 U21017 ( .A(n18382), .ZN(n18338) );
  AND2_X1 U21018 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18364), .ZN(n18383) );
  NOR2_X2 U21019 ( .A1(n18178), .A2(n17999), .ZN(n18381) );
  AOI22_X1 U21020 ( .A1(n18383), .A2(n18410), .B1(n18381), .B2(n18022), .ZN(
        n18002) );
  NAND2_X1 U21021 ( .A1(n18000), .A2(n18010), .ZN(n18386) );
  INV_X1 U21022 ( .A(n18386), .ZN(n18335) );
  AOI22_X1 U21023 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18025), .B1(
        n18086), .B2(n18335), .ZN(n18001) );
  OAI211_X1 U21024 ( .C1(n18338), .C2(n18343), .A(n18002), .B(n18001), .ZN(
        P3_U2871) );
  INV_X1 U21025 ( .A(n18086), .ZN(n18068) );
  NAND2_X1 U21026 ( .A1(n18010), .A2(n18003), .ZN(n18392) );
  NOR2_X2 U21027 ( .A1(n18178), .A2(n18004), .ZN(n18387) );
  INV_X1 U21028 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n18005) );
  NOR2_X2 U21029 ( .A1(n18006), .A2(n18005), .ZN(n18389) );
  AOI22_X1 U21030 ( .A1(n18387), .A2(n18022), .B1(n18389), .B2(n18352), .ZN(
        n18008) );
  AND2_X1 U21031 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18364), .ZN(n18388) );
  AOI22_X1 U21032 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18025), .B1(
        n18388), .B2(n18410), .ZN(n18007) );
  OAI211_X1 U21033 ( .C1(n18068), .C2(n18392), .A(n18008), .B(n18007), .ZN(
        P3_U2872) );
  NAND2_X1 U21034 ( .A1(n18010), .A2(n18009), .ZN(n18398) );
  NOR2_X2 U21035 ( .A1(n18011), .A2(n18006), .ZN(n18395) );
  NOR2_X2 U21036 ( .A1(n18178), .A2(n18012), .ZN(n18393) );
  AOI22_X1 U21037 ( .A1(n18395), .A2(n18410), .B1(n18393), .B2(n18022), .ZN(
        n18015) );
  NOR2_X2 U21038 ( .A1(n18006), .A2(n18013), .ZN(n18394) );
  AOI22_X1 U21039 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18025), .B1(
        n18394), .B2(n18352), .ZN(n18014) );
  OAI211_X1 U21040 ( .C1(n18068), .C2(n18398), .A(n18015), .B(n18014), .ZN(
        P3_U2873) );
  NOR2_X1 U21041 ( .A1(n18006), .A2(n19056), .ZN(n18344) );
  INV_X1 U21042 ( .A(n18344), .ZN(n18407) );
  NAND2_X1 U21043 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18364), .ZN(n18348) );
  INV_X1 U21044 ( .A(n18348), .ZN(n18402) );
  NOR2_X2 U21045 ( .A1(n18178), .A2(n18016), .ZN(n18400) );
  AOI22_X1 U21046 ( .A1(n18402), .A2(n18410), .B1(n18400), .B2(n18022), .ZN(
        n18019) );
  NOR2_X2 U21047 ( .A1(n18017), .A2(n18023), .ZN(n18403) );
  AOI22_X1 U21048 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18025), .B1(
        n18086), .B2(n18403), .ZN(n18018) );
  OAI211_X1 U21049 ( .C1(n18407), .C2(n18343), .A(n18019), .B(n18018), .ZN(
        P3_U2874) );
  NAND2_X1 U21050 ( .A1(n18364), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18418) );
  INV_X1 U21051 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n18020) );
  NOR2_X1 U21052 ( .A1(n18020), .A2(n18006), .ZN(n18411) );
  NOR2_X2 U21053 ( .A1(n18021), .A2(n18178), .ZN(n18409) );
  AOI22_X1 U21054 ( .A1(n18411), .A2(n18352), .B1(n18409), .B2(n18022), .ZN(
        n18027) );
  NOR2_X2 U21055 ( .A1(n18024), .A2(n18023), .ZN(n18412) );
  AOI22_X1 U21056 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18025), .B1(
        n18086), .B2(n18412), .ZN(n18026) );
  OAI211_X1 U21057 ( .C1(n18418), .C2(n18406), .A(n18027), .B(n18026), .ZN(
        P3_U2875) );
  INV_X1 U21058 ( .A(n18047), .ZN(n18070) );
  NOR2_X1 U21059 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18272), .ZN(
        n18202) );
  NAND2_X1 U21060 ( .A1(n18070), .A2(n18202), .ZN(n18111) );
  INV_X1 U21061 ( .A(n18330), .ZN(n18360) );
  NAND2_X1 U21062 ( .A1(n18457), .A2(n18250), .ZN(n18203) );
  NOR2_X1 U21063 ( .A1(n18047), .A2(n18203), .ZN(n18043) );
  AOI22_X1 U21064 ( .A1(n18360), .A2(n18352), .B1(n18359), .B2(n18043), .ZN(
        n18030) );
  NOR2_X1 U21065 ( .A1(n18178), .A2(n18028), .ZN(n18361) );
  INV_X1 U21066 ( .A(n18361), .ZN(n18069) );
  NOR2_X1 U21067 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18069), .ZN(
        n18300) );
  AOI22_X1 U21068 ( .A1(n18364), .A2(n18362), .B1(n18070), .B2(n18300), .ZN(
        n18044) );
  AOI22_X1 U21069 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18044), .B1(
        n18413), .B2(n18323), .ZN(n18029) );
  OAI211_X1 U21070 ( .C1(n18111), .C2(n18231), .A(n18030), .B(n18029), .ZN(
        P3_U2876) );
  AOI22_X1 U21071 ( .A1(n18369), .A2(n18043), .B1(n18278), .B2(n18352), .ZN(
        n18032) );
  INV_X1 U21072 ( .A(n18281), .ZN(n18370) );
  AOI22_X1 U21073 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18044), .B1(
        n18413), .B2(n18370), .ZN(n18031) );
  OAI211_X1 U21074 ( .C1(n18111), .C2(n18209), .A(n18032), .B(n18031), .ZN(
        P3_U2877) );
  INV_X1 U21075 ( .A(n18380), .ZN(n18282) );
  AOI22_X1 U21076 ( .A1(n18413), .A2(n18282), .B1(n18376), .B2(n18043), .ZN(
        n18034) );
  AOI22_X1 U21077 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18044), .B1(
        n18375), .B2(n18352), .ZN(n18033) );
  OAI211_X1 U21078 ( .C1(n18111), .C2(n18285), .A(n18034), .B(n18033), .ZN(
        P3_U2878) );
  AOI22_X1 U21079 ( .A1(n18383), .A2(n18352), .B1(n18381), .B2(n18043), .ZN(
        n18036) );
  INV_X1 U21080 ( .A(n18111), .ZN(n18104) );
  AOI22_X1 U21081 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18044), .B1(
        n18104), .B2(n18335), .ZN(n18035) );
  OAI211_X1 U21082 ( .C1(n18399), .C2(n18338), .A(n18036), .B(n18035), .ZN(
        P3_U2879) );
  AOI22_X1 U21083 ( .A1(n18413), .A2(n18389), .B1(n18387), .B2(n18043), .ZN(
        n18038) );
  AOI22_X1 U21084 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18044), .B1(
        n18388), .B2(n18352), .ZN(n18037) );
  OAI211_X1 U21085 ( .C1(n18111), .C2(n18392), .A(n18038), .B(n18037), .ZN(
        P3_U2880) );
  AOI22_X1 U21086 ( .A1(n18413), .A2(n18394), .B1(n18393), .B2(n18043), .ZN(
        n18040) );
  AOI22_X1 U21087 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18044), .B1(
        n18395), .B2(n18352), .ZN(n18039) );
  OAI211_X1 U21088 ( .C1(n18111), .C2(n18398), .A(n18040), .B(n18039), .ZN(
        P3_U2881) );
  AOI22_X1 U21089 ( .A1(n18402), .A2(n18352), .B1(n18400), .B2(n18043), .ZN(
        n18042) );
  AOI22_X1 U21090 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18044), .B1(
        n18104), .B2(n18403), .ZN(n18041) );
  OAI211_X1 U21091 ( .C1(n18399), .C2(n18407), .A(n18042), .B(n18041), .ZN(
        P3_U2882) );
  AOI22_X1 U21092 ( .A1(n18413), .A2(n18411), .B1(n18409), .B2(n18043), .ZN(
        n18046) );
  AOI22_X1 U21093 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18044), .B1(
        n18104), .B2(n18412), .ZN(n18045) );
  OAI211_X1 U21094 ( .C1(n18418), .C2(n18343), .A(n18046), .B(n18045), .ZN(
        P3_U2883) );
  NOR2_X1 U21095 ( .A1(n18457), .A2(n18047), .ZN(n18112) );
  NAND2_X1 U21096 ( .A1(n18112), .A2(n18272), .ZN(n18127) );
  AOI21_X1 U21097 ( .B1(n18127), .B2(n18111), .A(n18358), .ZN(n18064) );
  AOI22_X1 U21098 ( .A1(n18413), .A2(n18360), .B1(n18359), .B2(n18064), .ZN(
        n18051) );
  INV_X1 U21099 ( .A(n18127), .ZN(n18129) );
  AOI221_X1 U21100 ( .B1(n18048), .B2(n18111), .C1(n18324), .C2(n18111), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18049) );
  INV_X1 U21101 ( .A(n18178), .ZN(n18326) );
  OAI21_X1 U21102 ( .B1(n18129), .B2(n18049), .A(n18326), .ZN(n18065) );
  AOI22_X1 U21103 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18065), .B1(
        n18129), .B2(n18365), .ZN(n18050) );
  OAI211_X1 U21104 ( .C1(n18068), .C2(n18368), .A(n18051), .B(n18050), .ZN(
        P3_U2884) );
  AOI22_X1 U21105 ( .A1(n18413), .A2(n18278), .B1(n18064), .B2(n18369), .ZN(
        n18053) );
  AOI22_X1 U21106 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18065), .B1(
        n18129), .B2(n18371), .ZN(n18052) );
  OAI211_X1 U21107 ( .C1(n18068), .C2(n18281), .A(n18053), .B(n18052), .ZN(
        P3_U2885) );
  AOI22_X1 U21108 ( .A1(n18413), .A2(n18375), .B1(n18064), .B2(n18376), .ZN(
        n18055) );
  AOI22_X1 U21109 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18065), .B1(
        n18129), .B2(n18377), .ZN(n18054) );
  OAI211_X1 U21110 ( .C1(n18068), .C2(n18380), .A(n18055), .B(n18054), .ZN(
        P3_U2886) );
  AOI22_X1 U21111 ( .A1(n18413), .A2(n18383), .B1(n18064), .B2(n18381), .ZN(
        n18057) );
  AOI22_X1 U21112 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18065), .B1(
        n18129), .B2(n18335), .ZN(n18056) );
  OAI211_X1 U21113 ( .C1(n18068), .C2(n18338), .A(n18057), .B(n18056), .ZN(
        P3_U2887) );
  AOI22_X1 U21114 ( .A1(n18086), .A2(n18389), .B1(n18064), .B2(n18387), .ZN(
        n18059) );
  AOI22_X1 U21115 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18065), .B1(
        n18413), .B2(n18388), .ZN(n18058) );
  OAI211_X1 U21116 ( .C1(n18127), .C2(n18392), .A(n18059), .B(n18058), .ZN(
        P3_U2888) );
  AOI22_X1 U21117 ( .A1(n18086), .A2(n18394), .B1(n18064), .B2(n18393), .ZN(
        n18061) );
  AOI22_X1 U21118 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18065), .B1(
        n18413), .B2(n18395), .ZN(n18060) );
  OAI211_X1 U21119 ( .C1(n18127), .C2(n18398), .A(n18061), .B(n18060), .ZN(
        P3_U2889) );
  AOI22_X1 U21120 ( .A1(n18413), .A2(n18402), .B1(n18064), .B2(n18400), .ZN(
        n18063) );
  AOI22_X1 U21121 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18065), .B1(
        n18129), .B2(n18403), .ZN(n18062) );
  OAI211_X1 U21122 ( .C1(n18068), .C2(n18407), .A(n18063), .B(n18062), .ZN(
        P3_U2890) );
  INV_X1 U21123 ( .A(n18411), .ZN(n18356) );
  INV_X1 U21124 ( .A(n18418), .ZN(n18351) );
  AOI22_X1 U21125 ( .A1(n18413), .A2(n18351), .B1(n18064), .B2(n18409), .ZN(
        n18067) );
  AOI22_X1 U21126 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18065), .B1(
        n18129), .B2(n18412), .ZN(n18066) );
  OAI211_X1 U21127 ( .C1(n18068), .C2(n18356), .A(n18067), .B(n18066), .ZN(
        P3_U2891) );
  NAND2_X1 U21128 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18112), .ZN(
        n18140) );
  AND2_X1 U21129 ( .A1(n18250), .A2(n18112), .ZN(n18085) );
  AOI22_X1 U21130 ( .A1(n18086), .A2(n18360), .B1(n18359), .B2(n18085), .ZN(
        n18072) );
  AOI21_X1 U21131 ( .B1(n18457), .B2(n18324), .A(n18069), .ZN(n18157) );
  NAND2_X1 U21132 ( .A1(n18070), .A2(n18157), .ZN(n18087) );
  AOI22_X1 U21133 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18087), .B1(
        n18104), .B2(n18323), .ZN(n18071) );
  OAI211_X1 U21134 ( .C1(n18231), .C2(n18140), .A(n18072), .B(n18071), .ZN(
        P3_U2892) );
  AOI22_X1 U21135 ( .A1(n18086), .A2(n18278), .B1(n18369), .B2(n18085), .ZN(
        n18074) );
  AOI22_X1 U21136 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18087), .B1(
        n18104), .B2(n18370), .ZN(n18073) );
  OAI211_X1 U21137 ( .C1(n18209), .C2(n18140), .A(n18074), .B(n18073), .ZN(
        P3_U2893) );
  AOI22_X1 U21138 ( .A1(n18086), .A2(n18375), .B1(n18376), .B2(n18085), .ZN(
        n18076) );
  AOI22_X1 U21139 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18087), .B1(
        n18104), .B2(n18282), .ZN(n18075) );
  OAI211_X1 U21140 ( .C1(n18285), .C2(n18140), .A(n18076), .B(n18075), .ZN(
        P3_U2894) );
  AOI22_X1 U21141 ( .A1(n18104), .A2(n18382), .B1(n18381), .B2(n18085), .ZN(
        n18078) );
  AOI22_X1 U21142 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18087), .B1(
        n18086), .B2(n18383), .ZN(n18077) );
  OAI211_X1 U21143 ( .C1(n18386), .C2(n18140), .A(n18078), .B(n18077), .ZN(
        P3_U2895) );
  AOI22_X1 U21144 ( .A1(n18104), .A2(n18389), .B1(n18387), .B2(n18085), .ZN(
        n18080) );
  AOI22_X1 U21145 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18087), .B1(
        n18086), .B2(n18388), .ZN(n18079) );
  OAI211_X1 U21146 ( .C1(n18392), .C2(n18140), .A(n18080), .B(n18079), .ZN(
        P3_U2896) );
  AOI22_X1 U21147 ( .A1(n18086), .A2(n18395), .B1(n18393), .B2(n18085), .ZN(
        n18082) );
  AOI22_X1 U21148 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18087), .B1(
        n18104), .B2(n18394), .ZN(n18081) );
  OAI211_X1 U21149 ( .C1(n18398), .C2(n18140), .A(n18082), .B(n18081), .ZN(
        P3_U2897) );
  AOI22_X1 U21150 ( .A1(n18086), .A2(n18402), .B1(n18400), .B2(n18085), .ZN(
        n18084) );
  INV_X1 U21151 ( .A(n18140), .ZN(n18152) );
  AOI22_X1 U21152 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18087), .B1(
        n18403), .B2(n18152), .ZN(n18083) );
  OAI211_X1 U21153 ( .C1(n18111), .C2(n18407), .A(n18084), .B(n18083), .ZN(
        P3_U2898) );
  AOI22_X1 U21154 ( .A1(n18086), .A2(n18351), .B1(n18409), .B2(n18085), .ZN(
        n18089) );
  AOI22_X1 U21155 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18087), .B1(
        n18412), .B2(n18152), .ZN(n18088) );
  OAI211_X1 U21156 ( .C1(n18111), .C2(n18356), .A(n18089), .B(n18088), .ZN(
        P3_U2899) );
  INV_X1 U21157 ( .A(n18156), .ZN(n18133) );
  NOR2_X2 U21158 ( .A1(n18459), .A2(n18133), .ZN(n18168) );
  NOR2_X1 U21159 ( .A1(n18152), .A2(n18168), .ZN(n18134) );
  NOR2_X1 U21160 ( .A1(n18358), .A2(n18134), .ZN(n18107) );
  AOI22_X1 U21161 ( .A1(n18104), .A2(n18360), .B1(n18359), .B2(n18107), .ZN(
        n18093) );
  NOR2_X1 U21162 ( .A1(n18129), .A2(n18104), .ZN(n18090) );
  OAI21_X1 U21163 ( .B1(n18090), .B2(n18324), .A(n18134), .ZN(n18091) );
  OAI211_X1 U21164 ( .C1(n18168), .C2(n18586), .A(n18326), .B(n18091), .ZN(
        n18108) );
  AOI22_X1 U21165 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18108), .B1(
        n18365), .B2(n18168), .ZN(n18092) );
  OAI211_X1 U21166 ( .C1(n18127), .C2(n18368), .A(n18093), .B(n18092), .ZN(
        P3_U2900) );
  AOI22_X1 U21167 ( .A1(n18104), .A2(n18278), .B1(n18369), .B2(n18107), .ZN(
        n18095) );
  AOI22_X1 U21168 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18108), .B1(
        n18371), .B2(n18168), .ZN(n18094) );
  OAI211_X1 U21169 ( .C1(n18127), .C2(n18281), .A(n18095), .B(n18094), .ZN(
        P3_U2901) );
  INV_X1 U21170 ( .A(n18168), .ZN(n18177) );
  AOI22_X1 U21171 ( .A1(n18129), .A2(n18282), .B1(n18376), .B2(n18107), .ZN(
        n18097) );
  AOI22_X1 U21172 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18108), .B1(
        n18104), .B2(n18375), .ZN(n18096) );
  OAI211_X1 U21173 ( .C1(n18285), .C2(n18177), .A(n18097), .B(n18096), .ZN(
        P3_U2902) );
  AOI22_X1 U21174 ( .A1(n18104), .A2(n18383), .B1(n18381), .B2(n18107), .ZN(
        n18099) );
  AOI22_X1 U21175 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18108), .B1(
        n18335), .B2(n18168), .ZN(n18098) );
  OAI211_X1 U21176 ( .C1(n18127), .C2(n18338), .A(n18099), .B(n18098), .ZN(
        P3_U2903) );
  AOI22_X1 U21177 ( .A1(n18129), .A2(n18389), .B1(n18387), .B2(n18107), .ZN(
        n18101) );
  AOI22_X1 U21178 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18108), .B1(
        n18104), .B2(n18388), .ZN(n18100) );
  OAI211_X1 U21179 ( .C1(n18392), .C2(n18177), .A(n18101), .B(n18100), .ZN(
        P3_U2904) );
  AOI22_X1 U21180 ( .A1(n18129), .A2(n18394), .B1(n18393), .B2(n18107), .ZN(
        n18103) );
  AOI22_X1 U21181 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18108), .B1(
        n18104), .B2(n18395), .ZN(n18102) );
  OAI211_X1 U21182 ( .C1(n18398), .C2(n18177), .A(n18103), .B(n18102), .ZN(
        P3_U2905) );
  AOI22_X1 U21183 ( .A1(n18104), .A2(n18402), .B1(n18400), .B2(n18107), .ZN(
        n18106) );
  AOI22_X1 U21184 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18108), .B1(
        n18403), .B2(n18168), .ZN(n18105) );
  OAI211_X1 U21185 ( .C1(n18127), .C2(n18407), .A(n18106), .B(n18105), .ZN(
        P3_U2906) );
  AOI22_X1 U21186 ( .A1(n18129), .A2(n18411), .B1(n18409), .B2(n18107), .ZN(
        n18110) );
  AOI22_X1 U21187 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18108), .B1(
        n18412), .B2(n18168), .ZN(n18109) );
  OAI211_X1 U21188 ( .C1(n18111), .C2(n18418), .A(n18110), .B(n18109), .ZN(
        P3_U2907) );
  NAND2_X1 U21189 ( .A1(n18202), .A2(n18156), .ZN(n18200) );
  NOR2_X1 U21190 ( .A1(n18203), .A2(n18133), .ZN(n18128) );
  AOI22_X1 U21191 ( .A1(n18129), .A2(n18360), .B1(n18359), .B2(n18128), .ZN(
        n18114) );
  AOI22_X1 U21192 ( .A1(n18364), .A2(n18112), .B1(n18300), .B2(n18156), .ZN(
        n18130) );
  AOI22_X1 U21193 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18130), .B1(
        n18323), .B2(n18152), .ZN(n18113) );
  OAI211_X1 U21194 ( .C1(n18231), .C2(n18200), .A(n18114), .B(n18113), .ZN(
        P3_U2908) );
  AOI22_X1 U21195 ( .A1(n18370), .A2(n18152), .B1(n18369), .B2(n18128), .ZN(
        n18116) );
  AOI22_X1 U21196 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18130), .B1(
        n18129), .B2(n18278), .ZN(n18115) );
  OAI211_X1 U21197 ( .C1(n18209), .C2(n18200), .A(n18116), .B(n18115), .ZN(
        P3_U2909) );
  AOI22_X1 U21198 ( .A1(n18129), .A2(n18375), .B1(n18376), .B2(n18128), .ZN(
        n18118) );
  AOI22_X1 U21199 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18130), .B1(
        n18282), .B2(n18152), .ZN(n18117) );
  OAI211_X1 U21200 ( .C1(n18285), .C2(n18200), .A(n18118), .B(n18117), .ZN(
        P3_U2910) );
  AOI22_X1 U21201 ( .A1(n18129), .A2(n18383), .B1(n18381), .B2(n18128), .ZN(
        n18120) );
  AOI22_X1 U21202 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18130), .B1(
        n18382), .B2(n18152), .ZN(n18119) );
  OAI211_X1 U21203 ( .C1(n18386), .C2(n18200), .A(n18120), .B(n18119), .ZN(
        P3_U2911) );
  AOI22_X1 U21204 ( .A1(n18387), .A2(n18128), .B1(n18389), .B2(n18152), .ZN(
        n18122) );
  AOI22_X1 U21205 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18130), .B1(
        n18129), .B2(n18388), .ZN(n18121) );
  OAI211_X1 U21206 ( .C1(n18392), .C2(n18200), .A(n18122), .B(n18121), .ZN(
        P3_U2912) );
  AOI22_X1 U21207 ( .A1(n18394), .A2(n18152), .B1(n18393), .B2(n18128), .ZN(
        n18124) );
  AOI22_X1 U21208 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18130), .B1(
        n18129), .B2(n18395), .ZN(n18123) );
  OAI211_X1 U21209 ( .C1(n18398), .C2(n18200), .A(n18124), .B(n18123), .ZN(
        P3_U2913) );
  AOI22_X1 U21210 ( .A1(n18344), .A2(n18152), .B1(n18400), .B2(n18128), .ZN(
        n18126) );
  INV_X1 U21211 ( .A(n18200), .ZN(n18193) );
  AOI22_X1 U21212 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18130), .B1(
        n18403), .B2(n18193), .ZN(n18125) );
  OAI211_X1 U21213 ( .C1(n18127), .C2(n18348), .A(n18126), .B(n18125), .ZN(
        P3_U2914) );
  AOI22_X1 U21214 ( .A1(n18129), .A2(n18351), .B1(n18409), .B2(n18128), .ZN(
        n18132) );
  AOI22_X1 U21215 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18130), .B1(
        n18412), .B2(n18193), .ZN(n18131) );
  OAI211_X1 U21216 ( .C1(n18356), .C2(n18140), .A(n18132), .B(n18131), .ZN(
        P3_U2915) );
  NOR2_X1 U21217 ( .A1(n18457), .A2(n18133), .ZN(n18204) );
  NAND2_X1 U21218 ( .A1(n18272), .A2(n18204), .ZN(n18225) );
  INV_X1 U21219 ( .A(n18225), .ZN(n18218) );
  NOR2_X1 U21220 ( .A1(n18193), .A2(n18218), .ZN(n18179) );
  NOR2_X1 U21221 ( .A1(n18358), .A2(n18179), .ZN(n18151) );
  AOI22_X1 U21222 ( .A1(n18360), .A2(n18152), .B1(n18359), .B2(n18151), .ZN(
        n18137) );
  OAI21_X1 U21223 ( .B1(n18134), .B2(n18324), .A(n18179), .ZN(n18135) );
  OAI211_X1 U21224 ( .C1(n18218), .C2(n18586), .A(n18326), .B(n18135), .ZN(
        n18153) );
  AOI22_X1 U21225 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18153), .B1(
        n18365), .B2(n18218), .ZN(n18136) );
  OAI211_X1 U21226 ( .C1(n18368), .C2(n18177), .A(n18137), .B(n18136), .ZN(
        P3_U2916) );
  AOI22_X1 U21227 ( .A1(n18370), .A2(n18168), .B1(n18369), .B2(n18151), .ZN(
        n18139) );
  AOI22_X1 U21228 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18153), .B1(
        n18371), .B2(n18218), .ZN(n18138) );
  OAI211_X1 U21229 ( .C1(n18374), .C2(n18140), .A(n18139), .B(n18138), .ZN(
        P3_U2917) );
  AOI22_X1 U21230 ( .A1(n18282), .A2(n18168), .B1(n18376), .B2(n18151), .ZN(
        n18142) );
  AOI22_X1 U21231 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18153), .B1(
        n18375), .B2(n18152), .ZN(n18141) );
  OAI211_X1 U21232 ( .C1(n18285), .C2(n18225), .A(n18142), .B(n18141), .ZN(
        P3_U2918) );
  AOI22_X1 U21233 ( .A1(n18382), .A2(n18168), .B1(n18381), .B2(n18151), .ZN(
        n18144) );
  AOI22_X1 U21234 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18153), .B1(
        n18383), .B2(n18152), .ZN(n18143) );
  OAI211_X1 U21235 ( .C1(n18386), .C2(n18225), .A(n18144), .B(n18143), .ZN(
        P3_U2919) );
  AOI22_X1 U21236 ( .A1(n18388), .A2(n18152), .B1(n18387), .B2(n18151), .ZN(
        n18146) );
  AOI22_X1 U21237 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18153), .B1(
        n18389), .B2(n18168), .ZN(n18145) );
  OAI211_X1 U21238 ( .C1(n18392), .C2(n18225), .A(n18146), .B(n18145), .ZN(
        P3_U2920) );
  AOI22_X1 U21239 ( .A1(n18394), .A2(n18168), .B1(n18393), .B2(n18151), .ZN(
        n18148) );
  AOI22_X1 U21240 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18153), .B1(
        n18395), .B2(n18152), .ZN(n18147) );
  OAI211_X1 U21241 ( .C1(n18398), .C2(n18225), .A(n18148), .B(n18147), .ZN(
        P3_U2921) );
  AOI22_X1 U21242 ( .A1(n18402), .A2(n18152), .B1(n18400), .B2(n18151), .ZN(
        n18150) );
  AOI22_X1 U21243 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18153), .B1(
        n18403), .B2(n18218), .ZN(n18149) );
  OAI211_X1 U21244 ( .C1(n18407), .C2(n18177), .A(n18150), .B(n18149), .ZN(
        P3_U2922) );
  AOI22_X1 U21245 ( .A1(n18351), .A2(n18152), .B1(n18409), .B2(n18151), .ZN(
        n18155) );
  AOI22_X1 U21246 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18153), .B1(
        n18412), .B2(n18218), .ZN(n18154) );
  OAI211_X1 U21247 ( .C1(n18356), .C2(n18177), .A(n18155), .B(n18154), .ZN(
        P3_U2923) );
  AND2_X1 U21248 ( .A1(n18250), .A2(n18204), .ZN(n18173) );
  AOI22_X1 U21249 ( .A1(n18323), .A2(n18193), .B1(n18359), .B2(n18173), .ZN(
        n18159) );
  NAND2_X1 U21250 ( .A1(n18157), .A2(n18156), .ZN(n18174) );
  NAND2_X1 U21251 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18204), .ZN(
        n18249) );
  AOI22_X1 U21252 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18174), .B1(
        n18365), .B2(n18242), .ZN(n18158) );
  OAI211_X1 U21253 ( .C1(n18330), .C2(n18177), .A(n18159), .B(n18158), .ZN(
        P3_U2924) );
  AOI22_X1 U21254 ( .A1(n18370), .A2(n18193), .B1(n18369), .B2(n18173), .ZN(
        n18161) );
  AOI22_X1 U21255 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18174), .B1(
        n18371), .B2(n18242), .ZN(n18160) );
  OAI211_X1 U21256 ( .C1(n18374), .C2(n18177), .A(n18161), .B(n18160), .ZN(
        P3_U2925) );
  AOI22_X1 U21257 ( .A1(n18282), .A2(n18193), .B1(n18376), .B2(n18173), .ZN(
        n18163) );
  AOI22_X1 U21258 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18174), .B1(
        n18375), .B2(n18168), .ZN(n18162) );
  OAI211_X1 U21259 ( .C1(n18285), .C2(n18249), .A(n18163), .B(n18162), .ZN(
        P3_U2926) );
  AOI22_X1 U21260 ( .A1(n18383), .A2(n18168), .B1(n18381), .B2(n18173), .ZN(
        n18165) );
  AOI22_X1 U21261 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18174), .B1(
        n18335), .B2(n18242), .ZN(n18164) );
  OAI211_X1 U21262 ( .C1(n18338), .C2(n18200), .A(n18165), .B(n18164), .ZN(
        P3_U2927) );
  AOI22_X1 U21263 ( .A1(n18387), .A2(n18173), .B1(n18389), .B2(n18193), .ZN(
        n18167) );
  AOI22_X1 U21264 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18174), .B1(
        n18388), .B2(n18168), .ZN(n18166) );
  OAI211_X1 U21265 ( .C1(n18392), .C2(n18249), .A(n18167), .B(n18166), .ZN(
        P3_U2928) );
  AOI22_X1 U21266 ( .A1(n18394), .A2(n18193), .B1(n18393), .B2(n18173), .ZN(
        n18170) );
  AOI22_X1 U21267 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18174), .B1(
        n18395), .B2(n18168), .ZN(n18169) );
  OAI211_X1 U21268 ( .C1(n18398), .C2(n18249), .A(n18170), .B(n18169), .ZN(
        P3_U2929) );
  AOI22_X1 U21269 ( .A1(n18344), .A2(n18193), .B1(n18400), .B2(n18173), .ZN(
        n18172) );
  AOI22_X1 U21270 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18174), .B1(
        n18403), .B2(n18242), .ZN(n18171) );
  OAI211_X1 U21271 ( .C1(n18348), .C2(n18177), .A(n18172), .B(n18171), .ZN(
        P3_U2930) );
  AOI22_X1 U21272 ( .A1(n18411), .A2(n18193), .B1(n18409), .B2(n18173), .ZN(
        n18176) );
  AOI22_X1 U21273 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18174), .B1(
        n18412), .B2(n18242), .ZN(n18175) );
  OAI211_X1 U21274 ( .C1(n18418), .C2(n18177), .A(n18176), .B(n18175), .ZN(
        P3_U2931) );
  INV_X1 U21275 ( .A(n18201), .ZN(n18226) );
  NOR2_X2 U21276 ( .A1(n18459), .A2(n18226), .ZN(n18264) );
  NOR2_X1 U21277 ( .A1(n18242), .A2(n18264), .ZN(n18227) );
  NOR2_X1 U21278 ( .A1(n18358), .A2(n18227), .ZN(n18196) );
  AOI22_X1 U21279 ( .A1(n18360), .A2(n18193), .B1(n18359), .B2(n18196), .ZN(
        n18182) );
  OAI22_X1 U21280 ( .A1(n18179), .A2(n18006), .B1(n18227), .B2(n18178), .ZN(
        n18180) );
  OAI21_X1 U21281 ( .B1(n18264), .B2(n18586), .A(n18180), .ZN(n18197) );
  AOI22_X1 U21282 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18197), .B1(
        n18365), .B2(n18264), .ZN(n18181) );
  OAI211_X1 U21283 ( .C1(n18368), .C2(n18225), .A(n18182), .B(n18181), .ZN(
        P3_U2932) );
  AOI22_X1 U21284 ( .A1(n18369), .A2(n18196), .B1(n18278), .B2(n18193), .ZN(
        n18184) );
  AOI22_X1 U21285 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18197), .B1(
        n18371), .B2(n18264), .ZN(n18183) );
  OAI211_X1 U21286 ( .C1(n18281), .C2(n18225), .A(n18184), .B(n18183), .ZN(
        P3_U2933) );
  INV_X1 U21287 ( .A(n18264), .ZN(n18271) );
  AOI22_X1 U21288 ( .A1(n18282), .A2(n18218), .B1(n18376), .B2(n18196), .ZN(
        n18186) );
  AOI22_X1 U21289 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18197), .B1(
        n18375), .B2(n18193), .ZN(n18185) );
  OAI211_X1 U21290 ( .C1(n18285), .C2(n18271), .A(n18186), .B(n18185), .ZN(
        P3_U2934) );
  AOI22_X1 U21291 ( .A1(n18383), .A2(n18193), .B1(n18381), .B2(n18196), .ZN(
        n18188) );
  AOI22_X1 U21292 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18197), .B1(
        n18335), .B2(n18264), .ZN(n18187) );
  OAI211_X1 U21293 ( .C1(n18338), .C2(n18225), .A(n18188), .B(n18187), .ZN(
        P3_U2935) );
  AOI22_X1 U21294 ( .A1(n18387), .A2(n18196), .B1(n18389), .B2(n18218), .ZN(
        n18190) );
  AOI22_X1 U21295 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18197), .B1(
        n18388), .B2(n18193), .ZN(n18189) );
  OAI211_X1 U21296 ( .C1(n18392), .C2(n18271), .A(n18190), .B(n18189), .ZN(
        P3_U2936) );
  AOI22_X1 U21297 ( .A1(n18395), .A2(n18193), .B1(n18393), .B2(n18196), .ZN(
        n18192) );
  AOI22_X1 U21298 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18197), .B1(
        n18394), .B2(n18218), .ZN(n18191) );
  OAI211_X1 U21299 ( .C1(n18398), .C2(n18271), .A(n18192), .B(n18191), .ZN(
        P3_U2937) );
  AOI22_X1 U21300 ( .A1(n18402), .A2(n18193), .B1(n18400), .B2(n18196), .ZN(
        n18195) );
  AOI22_X1 U21301 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18197), .B1(
        n18403), .B2(n18264), .ZN(n18194) );
  OAI211_X1 U21302 ( .C1(n18407), .C2(n18225), .A(n18195), .B(n18194), .ZN(
        P3_U2938) );
  AOI22_X1 U21303 ( .A1(n18411), .A2(n18218), .B1(n18409), .B2(n18196), .ZN(
        n18199) );
  AOI22_X1 U21304 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18197), .B1(
        n18412), .B2(n18264), .ZN(n18198) );
  OAI211_X1 U21305 ( .C1(n18418), .C2(n18200), .A(n18199), .B(n18198), .ZN(
        P3_U2939) );
  NAND2_X1 U21306 ( .A1(n18202), .A2(n18201), .ZN(n18277) );
  NOR2_X1 U21307 ( .A1(n18226), .A2(n18203), .ZN(n18221) );
  AOI22_X1 U21308 ( .A1(n18323), .A2(n18242), .B1(n18359), .B2(n18221), .ZN(
        n18206) );
  NOR2_X1 U21309 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18226), .ZN(
        n18251) );
  AOI22_X1 U21310 ( .A1(n18364), .A2(n18204), .B1(n18361), .B2(n18251), .ZN(
        n18222) );
  AOI22_X1 U21311 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18222), .B1(
        n18360), .B2(n18218), .ZN(n18205) );
  OAI211_X1 U21312 ( .C1(n18231), .C2(n18277), .A(n18206), .B(n18205), .ZN(
        P3_U2940) );
  AOI22_X1 U21313 ( .A1(n18369), .A2(n18221), .B1(n18278), .B2(n18218), .ZN(
        n18208) );
  AOI22_X1 U21314 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18222), .B1(
        n18370), .B2(n18242), .ZN(n18207) );
  OAI211_X1 U21315 ( .C1(n18209), .C2(n18277), .A(n18208), .B(n18207), .ZN(
        P3_U2941) );
  AOI22_X1 U21316 ( .A1(n18376), .A2(n18221), .B1(n18375), .B2(n18218), .ZN(
        n18211) );
  AOI22_X1 U21317 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18222), .B1(
        n18282), .B2(n18242), .ZN(n18210) );
  OAI211_X1 U21318 ( .C1(n18285), .C2(n18277), .A(n18211), .B(n18210), .ZN(
        P3_U2942) );
  AOI22_X1 U21319 ( .A1(n18382), .A2(n18242), .B1(n18381), .B2(n18221), .ZN(
        n18213) );
  AOI22_X1 U21320 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18222), .B1(
        n18383), .B2(n18218), .ZN(n18212) );
  OAI211_X1 U21321 ( .C1(n18386), .C2(n18277), .A(n18213), .B(n18212), .ZN(
        P3_U2943) );
  AOI22_X1 U21322 ( .A1(n18388), .A2(n18218), .B1(n18387), .B2(n18221), .ZN(
        n18215) );
  AOI22_X1 U21323 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18222), .B1(
        n18389), .B2(n18242), .ZN(n18214) );
  OAI211_X1 U21324 ( .C1(n18392), .C2(n18277), .A(n18215), .B(n18214), .ZN(
        P3_U2944) );
  AOI22_X1 U21325 ( .A1(n18395), .A2(n18218), .B1(n18393), .B2(n18221), .ZN(
        n18217) );
  AOI22_X1 U21326 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18222), .B1(
        n18394), .B2(n18242), .ZN(n18216) );
  OAI211_X1 U21327 ( .C1(n18398), .C2(n18277), .A(n18217), .B(n18216), .ZN(
        P3_U2945) );
  AOI22_X1 U21328 ( .A1(n18402), .A2(n18218), .B1(n18400), .B2(n18221), .ZN(
        n18220) );
  INV_X1 U21329 ( .A(n18277), .ZN(n18295) );
  AOI22_X1 U21330 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18222), .B1(
        n18403), .B2(n18295), .ZN(n18219) );
  OAI211_X1 U21331 ( .C1(n18407), .C2(n18249), .A(n18220), .B(n18219), .ZN(
        P3_U2946) );
  AOI22_X1 U21332 ( .A1(n18411), .A2(n18242), .B1(n18409), .B2(n18221), .ZN(
        n18224) );
  AOI22_X1 U21333 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18222), .B1(
        n18412), .B2(n18295), .ZN(n18223) );
  OAI211_X1 U21334 ( .C1(n18418), .C2(n18225), .A(n18224), .B(n18223), .ZN(
        P3_U2947) );
  NOR2_X1 U21335 ( .A1(n18457), .A2(n18226), .ZN(n18302) );
  NAND2_X1 U21336 ( .A1(n18302), .A2(n18272), .ZN(n18317) );
  NOR2_X1 U21337 ( .A1(n18295), .A2(n18319), .ZN(n18273) );
  NOR2_X1 U21338 ( .A1(n18358), .A2(n18273), .ZN(n18245) );
  AOI22_X1 U21339 ( .A1(n18360), .A2(n18242), .B1(n18359), .B2(n18245), .ZN(
        n18230) );
  OAI21_X1 U21340 ( .B1(n18227), .B2(n18324), .A(n18273), .ZN(n18228) );
  OAI211_X1 U21341 ( .C1(n18319), .C2(n18586), .A(n18326), .B(n18228), .ZN(
        n18246) );
  AOI22_X1 U21342 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18246), .B1(
        n18323), .B2(n18264), .ZN(n18229) );
  OAI211_X1 U21343 ( .C1(n18231), .C2(n18317), .A(n18230), .B(n18229), .ZN(
        P3_U2948) );
  AOI22_X1 U21344 ( .A1(n18370), .A2(n18264), .B1(n18369), .B2(n18245), .ZN(
        n18233) );
  AOI22_X1 U21345 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18246), .B1(
        n18371), .B2(n18319), .ZN(n18232) );
  OAI211_X1 U21346 ( .C1(n18374), .C2(n18249), .A(n18233), .B(n18232), .ZN(
        P3_U2949) );
  AOI22_X1 U21347 ( .A1(n18282), .A2(n18264), .B1(n18376), .B2(n18245), .ZN(
        n18235) );
  AOI22_X1 U21348 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18246), .B1(
        n18375), .B2(n18242), .ZN(n18234) );
  OAI211_X1 U21349 ( .C1(n18285), .C2(n18317), .A(n18235), .B(n18234), .ZN(
        P3_U2950) );
  AOI22_X1 U21350 ( .A1(n18383), .A2(n18242), .B1(n18381), .B2(n18245), .ZN(
        n18237) );
  AOI22_X1 U21351 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18246), .B1(
        n18335), .B2(n18319), .ZN(n18236) );
  OAI211_X1 U21352 ( .C1(n18338), .C2(n18271), .A(n18237), .B(n18236), .ZN(
        P3_U2951) );
  AOI22_X1 U21353 ( .A1(n18387), .A2(n18245), .B1(n18389), .B2(n18264), .ZN(
        n18239) );
  AOI22_X1 U21354 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18246), .B1(
        n18388), .B2(n18242), .ZN(n18238) );
  OAI211_X1 U21355 ( .C1(n18392), .C2(n18317), .A(n18239), .B(n18238), .ZN(
        P3_U2952) );
  AOI22_X1 U21356 ( .A1(n18395), .A2(n18242), .B1(n18393), .B2(n18245), .ZN(
        n18241) );
  AOI22_X1 U21357 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18246), .B1(
        n18394), .B2(n18264), .ZN(n18240) );
  OAI211_X1 U21358 ( .C1(n18398), .C2(n18317), .A(n18241), .B(n18240), .ZN(
        P3_U2953) );
  AOI22_X1 U21359 ( .A1(n18402), .A2(n18242), .B1(n18400), .B2(n18245), .ZN(
        n18244) );
  AOI22_X1 U21360 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18246), .B1(
        n18403), .B2(n18319), .ZN(n18243) );
  OAI211_X1 U21361 ( .C1(n18407), .C2(n18271), .A(n18244), .B(n18243), .ZN(
        P3_U2954) );
  AOI22_X1 U21362 ( .A1(n18411), .A2(n18264), .B1(n18409), .B2(n18245), .ZN(
        n18248) );
  AOI22_X1 U21363 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18246), .B1(
        n18412), .B2(n18319), .ZN(n18247) );
  OAI211_X1 U21364 ( .C1(n18418), .C2(n18249), .A(n18248), .B(n18247), .ZN(
        P3_U2955) );
  AND2_X1 U21365 ( .A1(n18250), .A2(n18302), .ZN(n18267) );
  AOI22_X1 U21366 ( .A1(n18323), .A2(n18295), .B1(n18359), .B2(n18267), .ZN(
        n18253) );
  AOI22_X1 U21367 ( .A1(n18364), .A2(n18251), .B1(n18302), .B2(n18361), .ZN(
        n18268) );
  NAND2_X1 U21368 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18302), .ZN(
        n18347) );
  INV_X1 U21369 ( .A(n18347), .ZN(n18350) );
  AOI22_X1 U21370 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18268), .B1(
        n18365), .B2(n18350), .ZN(n18252) );
  OAI211_X1 U21371 ( .C1(n18330), .C2(n18271), .A(n18253), .B(n18252), .ZN(
        P3_U2956) );
  AOI22_X1 U21372 ( .A1(n18370), .A2(n18295), .B1(n18369), .B2(n18267), .ZN(
        n18255) );
  AOI22_X1 U21373 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18268), .B1(
        n18371), .B2(n18350), .ZN(n18254) );
  OAI211_X1 U21374 ( .C1(n18374), .C2(n18271), .A(n18255), .B(n18254), .ZN(
        P3_U2957) );
  AOI22_X1 U21375 ( .A1(n18376), .A2(n18267), .B1(n18375), .B2(n18264), .ZN(
        n18257) );
  AOI22_X1 U21376 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18268), .B1(
        n18377), .B2(n18350), .ZN(n18256) );
  OAI211_X1 U21377 ( .C1(n18380), .C2(n18277), .A(n18257), .B(n18256), .ZN(
        P3_U2958) );
  AOI22_X1 U21378 ( .A1(n18383), .A2(n18264), .B1(n18381), .B2(n18267), .ZN(
        n18259) );
  AOI22_X1 U21379 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18268), .B1(
        n18335), .B2(n18350), .ZN(n18258) );
  OAI211_X1 U21380 ( .C1(n18338), .C2(n18277), .A(n18259), .B(n18258), .ZN(
        P3_U2959) );
  AOI22_X1 U21381 ( .A1(n18388), .A2(n18264), .B1(n18387), .B2(n18267), .ZN(
        n18261) );
  AOI22_X1 U21382 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18268), .B1(
        n18389), .B2(n18295), .ZN(n18260) );
  OAI211_X1 U21383 ( .C1(n18392), .C2(n18347), .A(n18261), .B(n18260), .ZN(
        P3_U2960) );
  AOI22_X1 U21384 ( .A1(n18394), .A2(n18295), .B1(n18393), .B2(n18267), .ZN(
        n18263) );
  AOI22_X1 U21385 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18268), .B1(
        n18395), .B2(n18264), .ZN(n18262) );
  OAI211_X1 U21386 ( .C1(n18398), .C2(n18347), .A(n18263), .B(n18262), .ZN(
        P3_U2961) );
  AOI22_X1 U21387 ( .A1(n18402), .A2(n18264), .B1(n18400), .B2(n18267), .ZN(
        n18266) );
  AOI22_X1 U21388 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18268), .B1(
        n18403), .B2(n18350), .ZN(n18265) );
  OAI211_X1 U21389 ( .C1(n18407), .C2(n18277), .A(n18266), .B(n18265), .ZN(
        P3_U2962) );
  AOI22_X1 U21390 ( .A1(n18411), .A2(n18295), .B1(n18409), .B2(n18267), .ZN(
        n18270) );
  AOI22_X1 U21391 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18268), .B1(
        n18412), .B2(n18350), .ZN(n18269) );
  OAI211_X1 U21392 ( .C1(n18418), .C2(n18271), .A(n18270), .B(n18269), .ZN(
        P3_U2963) );
  INV_X1 U21393 ( .A(n18299), .ZN(n18363) );
  NAND2_X1 U21394 ( .A1(n18272), .A2(n18363), .ZN(n18417) );
  INV_X1 U21395 ( .A(n18417), .ZN(n18401) );
  NOR2_X1 U21396 ( .A1(n18350), .A2(n18401), .ZN(n18325) );
  NOR2_X1 U21397 ( .A1(n18358), .A2(n18325), .ZN(n18294) );
  AOI22_X1 U21398 ( .A1(n18323), .A2(n18319), .B1(n18359), .B2(n18294), .ZN(
        n18276) );
  OAI21_X1 U21399 ( .B1(n18273), .B2(n18324), .A(n18325), .ZN(n18274) );
  OAI211_X1 U21400 ( .C1(n18401), .C2(n18586), .A(n18326), .B(n18274), .ZN(
        n18296) );
  AOI22_X1 U21401 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18296), .B1(
        n18365), .B2(n18401), .ZN(n18275) );
  OAI211_X1 U21402 ( .C1(n18330), .C2(n18277), .A(n18276), .B(n18275), .ZN(
        P3_U2964) );
  AOI22_X1 U21403 ( .A1(n18369), .A2(n18294), .B1(n18278), .B2(n18295), .ZN(
        n18280) );
  AOI22_X1 U21404 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18296), .B1(
        n18371), .B2(n18401), .ZN(n18279) );
  OAI211_X1 U21405 ( .C1(n18281), .C2(n18317), .A(n18280), .B(n18279), .ZN(
        P3_U2965) );
  AOI22_X1 U21406 ( .A1(n18282), .A2(n18319), .B1(n18376), .B2(n18294), .ZN(
        n18284) );
  AOI22_X1 U21407 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18296), .B1(
        n18375), .B2(n18295), .ZN(n18283) );
  OAI211_X1 U21408 ( .C1(n18285), .C2(n18417), .A(n18284), .B(n18283), .ZN(
        P3_U2966) );
  AOI22_X1 U21409 ( .A1(n18383), .A2(n18295), .B1(n18381), .B2(n18294), .ZN(
        n18287) );
  AOI22_X1 U21410 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18296), .B1(
        n18335), .B2(n18401), .ZN(n18286) );
  OAI211_X1 U21411 ( .C1(n18338), .C2(n18317), .A(n18287), .B(n18286), .ZN(
        P3_U2967) );
  AOI22_X1 U21412 ( .A1(n18388), .A2(n18295), .B1(n18387), .B2(n18294), .ZN(
        n18289) );
  AOI22_X1 U21413 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18296), .B1(
        n18389), .B2(n18319), .ZN(n18288) );
  OAI211_X1 U21414 ( .C1(n18392), .C2(n18417), .A(n18289), .B(n18288), .ZN(
        P3_U2968) );
  AOI22_X1 U21415 ( .A1(n18395), .A2(n18295), .B1(n18393), .B2(n18294), .ZN(
        n18291) );
  AOI22_X1 U21416 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18296), .B1(
        n18394), .B2(n18319), .ZN(n18290) );
  OAI211_X1 U21417 ( .C1(n18398), .C2(n18417), .A(n18291), .B(n18290), .ZN(
        P3_U2969) );
  AOI22_X1 U21418 ( .A1(n18402), .A2(n18295), .B1(n18400), .B2(n18294), .ZN(
        n18293) );
  AOI22_X1 U21419 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18296), .B1(
        n18403), .B2(n18401), .ZN(n18292) );
  OAI211_X1 U21420 ( .C1(n18407), .C2(n18317), .A(n18293), .B(n18292), .ZN(
        P3_U2970) );
  AOI22_X1 U21421 ( .A1(n18351), .A2(n18295), .B1(n18409), .B2(n18294), .ZN(
        n18298) );
  AOI22_X1 U21422 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18296), .B1(
        n18412), .B2(n18401), .ZN(n18297) );
  OAI211_X1 U21423 ( .C1(n18356), .C2(n18317), .A(n18298), .B(n18297), .ZN(
        P3_U2971) );
  NOR2_X1 U21424 ( .A1(n18358), .A2(n18299), .ZN(n18318) );
  AOI22_X1 U21425 ( .A1(n18360), .A2(n18319), .B1(n18359), .B2(n18318), .ZN(
        n18304) );
  AOI22_X1 U21426 ( .A1(n18364), .A2(n18302), .B1(n18301), .B2(n18300), .ZN(
        n18320) );
  AOI22_X1 U21427 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18320), .B1(
        n18365), .B2(n18410), .ZN(n18303) );
  OAI211_X1 U21428 ( .C1(n18368), .C2(n18347), .A(n18304), .B(n18303), .ZN(
        P3_U2972) );
  AOI22_X1 U21429 ( .A1(n18370), .A2(n18350), .B1(n18369), .B2(n18318), .ZN(
        n18306) );
  AOI22_X1 U21430 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18320), .B1(
        n18371), .B2(n18410), .ZN(n18305) );
  OAI211_X1 U21431 ( .C1(n18374), .C2(n18317), .A(n18306), .B(n18305), .ZN(
        P3_U2973) );
  AOI22_X1 U21432 ( .A1(n18376), .A2(n18318), .B1(n18375), .B2(n18319), .ZN(
        n18308) );
  AOI22_X1 U21433 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18320), .B1(
        n18377), .B2(n18410), .ZN(n18307) );
  OAI211_X1 U21434 ( .C1(n18380), .C2(n18347), .A(n18308), .B(n18307), .ZN(
        P3_U2974) );
  AOI22_X1 U21435 ( .A1(n18383), .A2(n18319), .B1(n18381), .B2(n18318), .ZN(
        n18310) );
  AOI22_X1 U21436 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18320), .B1(
        n18335), .B2(n18410), .ZN(n18309) );
  OAI211_X1 U21437 ( .C1(n18338), .C2(n18347), .A(n18310), .B(n18309), .ZN(
        P3_U2975) );
  AOI22_X1 U21438 ( .A1(n18387), .A2(n18318), .B1(n18389), .B2(n18350), .ZN(
        n18312) );
  AOI22_X1 U21439 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18320), .B1(
        n18388), .B2(n18319), .ZN(n18311) );
  OAI211_X1 U21440 ( .C1(n18392), .C2(n18406), .A(n18312), .B(n18311), .ZN(
        P3_U2976) );
  AOI22_X1 U21441 ( .A1(n18394), .A2(n18350), .B1(n18393), .B2(n18318), .ZN(
        n18314) );
  AOI22_X1 U21442 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18320), .B1(
        n18395), .B2(n18319), .ZN(n18313) );
  OAI211_X1 U21443 ( .C1(n18398), .C2(n18406), .A(n18314), .B(n18313), .ZN(
        P3_U2977) );
  AOI22_X1 U21444 ( .A1(n18344), .A2(n18350), .B1(n18400), .B2(n18318), .ZN(
        n18316) );
  AOI22_X1 U21445 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18320), .B1(
        n18403), .B2(n18410), .ZN(n18315) );
  OAI211_X1 U21446 ( .C1(n18348), .C2(n18317), .A(n18316), .B(n18315), .ZN(
        P3_U2978) );
  AOI22_X1 U21447 ( .A1(n18351), .A2(n18319), .B1(n18409), .B2(n18318), .ZN(
        n18322) );
  AOI22_X1 U21448 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18320), .B1(
        n18412), .B2(n18410), .ZN(n18321) );
  OAI211_X1 U21449 ( .C1(n18356), .C2(n18347), .A(n18322), .B(n18321), .ZN(
        P3_U2979) );
  AOI21_X1 U21450 ( .B1(n18343), .B2(n18406), .A(n18358), .ZN(n18349) );
  AOI22_X1 U21451 ( .A1(n18323), .A2(n18401), .B1(n18359), .B2(n18349), .ZN(
        n18329) );
  AOI221_X1 U21452 ( .B1(n18325), .B2(n18406), .C1(n18324), .C2(n18406), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18327) );
  OAI21_X1 U21453 ( .B1(n18352), .B2(n18327), .A(n18326), .ZN(n18353) );
  AOI22_X1 U21454 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18353), .B1(
        n18365), .B2(n18352), .ZN(n18328) );
  OAI211_X1 U21455 ( .C1(n18330), .C2(n18347), .A(n18329), .B(n18328), .ZN(
        P3_U2980) );
  AOI22_X1 U21456 ( .A1(n18370), .A2(n18401), .B1(n18369), .B2(n18349), .ZN(
        n18332) );
  AOI22_X1 U21457 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18353), .B1(
        n18371), .B2(n18352), .ZN(n18331) );
  OAI211_X1 U21458 ( .C1(n18374), .C2(n18347), .A(n18332), .B(n18331), .ZN(
        P3_U2981) );
  AOI22_X1 U21459 ( .A1(n18376), .A2(n18349), .B1(n18375), .B2(n18350), .ZN(
        n18334) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18353), .B1(
        n18377), .B2(n18352), .ZN(n18333) );
  OAI211_X1 U21461 ( .C1(n18380), .C2(n18417), .A(n18334), .B(n18333), .ZN(
        P3_U2982) );
  AOI22_X1 U21462 ( .A1(n18383), .A2(n18350), .B1(n18381), .B2(n18349), .ZN(
        n18337) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18353), .B1(
        n18335), .B2(n18352), .ZN(n18336) );
  OAI211_X1 U21464 ( .C1(n18338), .C2(n18417), .A(n18337), .B(n18336), .ZN(
        P3_U2983) );
  AOI22_X1 U21465 ( .A1(n18387), .A2(n18349), .B1(n18389), .B2(n18401), .ZN(
        n18340) );
  AOI22_X1 U21466 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18353), .B1(
        n18388), .B2(n18350), .ZN(n18339) );
  OAI211_X1 U21467 ( .C1(n18392), .C2(n18343), .A(n18340), .B(n18339), .ZN(
        P3_U2984) );
  AOI22_X1 U21468 ( .A1(n18394), .A2(n18401), .B1(n18393), .B2(n18349), .ZN(
        n18342) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18353), .B1(
        n18395), .B2(n18350), .ZN(n18341) );
  OAI211_X1 U21470 ( .C1(n18398), .C2(n18343), .A(n18342), .B(n18341), .ZN(
        P3_U2985) );
  AOI22_X1 U21471 ( .A1(n18344), .A2(n18401), .B1(n18400), .B2(n18349), .ZN(
        n18346) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18353), .B1(
        n18403), .B2(n18352), .ZN(n18345) );
  OAI211_X1 U21473 ( .C1(n18348), .C2(n18347), .A(n18346), .B(n18345), .ZN(
        P3_U2986) );
  AOI22_X1 U21474 ( .A1(n18351), .A2(n18350), .B1(n18409), .B2(n18349), .ZN(
        n18355) );
  AOI22_X1 U21475 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18353), .B1(
        n18412), .B2(n18352), .ZN(n18354) );
  OAI211_X1 U21476 ( .C1(n18356), .C2(n18417), .A(n18355), .B(n18354), .ZN(
        P3_U2987) );
  NOR2_X1 U21477 ( .A1(n18358), .A2(n18357), .ZN(n18408) );
  AOI22_X1 U21478 ( .A1(n18360), .A2(n18401), .B1(n18359), .B2(n18408), .ZN(
        n18367) );
  AOI22_X1 U21479 ( .A1(n18364), .A2(n18363), .B1(n18362), .B2(n18361), .ZN(
        n18414) );
  AOI22_X1 U21480 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18414), .B1(
        n18413), .B2(n18365), .ZN(n18366) );
  OAI211_X1 U21481 ( .C1(n18368), .C2(n18406), .A(n18367), .B(n18366), .ZN(
        P3_U2988) );
  AOI22_X1 U21482 ( .A1(n18370), .A2(n18410), .B1(n18369), .B2(n18408), .ZN(
        n18373) );
  AOI22_X1 U21483 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18414), .B1(
        n18413), .B2(n18371), .ZN(n18372) );
  OAI211_X1 U21484 ( .C1(n18374), .C2(n18417), .A(n18373), .B(n18372), .ZN(
        P3_U2989) );
  AOI22_X1 U21485 ( .A1(n18376), .A2(n18408), .B1(n18375), .B2(n18401), .ZN(
        n18379) );
  AOI22_X1 U21486 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18414), .B1(
        n18413), .B2(n18377), .ZN(n18378) );
  OAI211_X1 U21487 ( .C1(n18380), .C2(n18406), .A(n18379), .B(n18378), .ZN(
        P3_U2990) );
  AOI22_X1 U21488 ( .A1(n18382), .A2(n18410), .B1(n18381), .B2(n18408), .ZN(
        n18385) );
  AOI22_X1 U21489 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18414), .B1(
        n18383), .B2(n18401), .ZN(n18384) );
  OAI211_X1 U21490 ( .C1(n18399), .C2(n18386), .A(n18385), .B(n18384), .ZN(
        P3_U2991) );
  AOI22_X1 U21491 ( .A1(n18388), .A2(n18401), .B1(n18387), .B2(n18408), .ZN(
        n18391) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18414), .B1(
        n18389), .B2(n18410), .ZN(n18390) );
  OAI211_X1 U21493 ( .C1(n18399), .C2(n18392), .A(n18391), .B(n18390), .ZN(
        P3_U2992) );
  AOI22_X1 U21494 ( .A1(n18394), .A2(n18410), .B1(n18393), .B2(n18408), .ZN(
        n18397) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18414), .B1(
        n18395), .B2(n18401), .ZN(n18396) );
  OAI211_X1 U21496 ( .C1(n18399), .C2(n18398), .A(n18397), .B(n18396), .ZN(
        P3_U2993) );
  AOI22_X1 U21497 ( .A1(n18402), .A2(n18401), .B1(n18400), .B2(n18408), .ZN(
        n18405) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18414), .B1(
        n18413), .B2(n18403), .ZN(n18404) );
  OAI211_X1 U21499 ( .C1(n18407), .C2(n18406), .A(n18405), .B(n18404), .ZN(
        P3_U2994) );
  AOI22_X1 U21500 ( .A1(n18411), .A2(n18410), .B1(n18409), .B2(n18408), .ZN(
        n18416) );
  AOI22_X1 U21501 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18414), .B1(
        n18413), .B2(n18412), .ZN(n18415) );
  OAI211_X1 U21502 ( .C1(n18418), .C2(n18417), .A(n18416), .B(n18415), .ZN(
        P3_U2995) );
  NAND2_X1 U21503 ( .A1(n18420), .A2(n18419), .ZN(n18423) );
  AOI22_X1 U21504 ( .A1(n18424), .A2(n18423), .B1(n18422), .B2(n18421), .ZN(
        n18425) );
  OAI221_X1 U21505 ( .B1(n18428), .B2(n18427), .C1(n18428), .C2(n18426), .A(
        n18425), .ZN(n18624) );
  OAI21_X1 U21506 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18429), .ZN(n18431) );
  OAI211_X1 U21507 ( .C1(n18450), .C2(n18478), .A(n18431), .B(n18430), .ZN(
        n18472) );
  INV_X1 U21508 ( .A(n18450), .ZN(n18461) );
  NAND3_X1 U21509 ( .A1(n18433), .A2(n18432), .A3(n18453), .ZN(n18444) );
  INV_X1 U21510 ( .A(n18440), .ZN(n18436) );
  OAI21_X1 U21511 ( .B1(n18434), .B2(n18433), .A(n18432), .ZN(n18435) );
  AND2_X1 U21512 ( .A1(n18612), .A2(n18435), .ZN(n18445) );
  AOI211_X1 U21513 ( .C1(n18444), .C2(n18436), .A(n18445), .B(n18590), .ZN(
        n18443) );
  AOI21_X1 U21514 ( .B1(n18438), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n18437), .ZN(n18454) );
  INV_X1 U21515 ( .A(n18454), .ZN(n18439) );
  AOI22_X1 U21516 ( .A1(n18449), .A2(n18442), .B1(n18440), .B2(n18439), .ZN(
        n18441) );
  AOI22_X1 U21517 ( .A1(n18443), .A2(n18442), .B1(n18441), .B2(n18590), .ZN(
        n18588) );
  AOI22_X1 U21518 ( .A1(n18461), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n18588), .B2(n18450), .ZN(n18470) );
  NOR3_X1 U21519 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18604), .A3(
        n18454), .ZN(n18448) );
  OAI211_X1 U21520 ( .C1(n18604), .C2(n18445), .A(n18444), .B(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18446) );
  INV_X1 U21521 ( .A(n18446), .ZN(n18447) );
  AOI211_X1 U21522 ( .C1(n18449), .C2(n18592), .A(n18448), .B(n18447), .ZN(
        n18594) );
  AOI22_X1 U21523 ( .A1(n18461), .A2(n11052), .B1(n18594), .B2(n18450), .ZN(
        n18465) );
  AND2_X1 U21524 ( .A1(n18452), .A2(n18451), .ZN(n18455) );
  AOI22_X1 U21525 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18453), .B1(
        n18455), .B2(n18612), .ZN(n18458) );
  OAI22_X1 U21526 ( .A1(n18455), .A2(n18598), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18454), .ZN(n18602) );
  INV_X1 U21527 ( .A(n18458), .ZN(n18606) );
  NAND3_X1 U21528 ( .A1(n18606), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18456) );
  AOI22_X1 U21529 ( .A1(n18458), .A2(n18457), .B1(n18602), .B2(n18456), .ZN(
        n18460) );
  OAI21_X1 U21530 ( .B1(n18461), .B2(n18460), .A(n18459), .ZN(n18464) );
  AND2_X1 U21531 ( .A1(n18465), .A2(n18464), .ZN(n18462) );
  OAI221_X1 U21532 ( .B1(n18465), .B2(n18464), .C1(n18463), .C2(n18462), .A(
        n18467), .ZN(n18469) );
  AOI21_X1 U21533 ( .B1(n18467), .B2(n18466), .A(n18465), .ZN(n18468) );
  AOI222_X1 U21534 ( .A1(n18470), .A2(n18469), .B1(n18470), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18469), .C2(n18468), .ZN(
        n18471) );
  OR4_X1 U21535 ( .A1(n18473), .A2(n18624), .A3(n18472), .A4(n18471), .ZN(
        n18482) );
  AOI211_X1 U21536 ( .C1(n18475), .C2(n18474), .A(n18490), .B(n18482), .ZN(
        n18476) );
  INV_X1 U21537 ( .A(n18476), .ZN(n18585) );
  OAI21_X1 U21538 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18632), .A(n18585), 
        .ZN(n18491) );
  NOR3_X1 U21539 ( .A1(n18479), .A2(n18477), .A3(n18491), .ZN(n18485) );
  AOI22_X1 U21540 ( .A1(n18480), .A2(n18504), .B1(n18479), .B2(n18478), .ZN(
        n18481) );
  AOI22_X1 U21541 ( .A1(n18483), .A2(n18482), .B1(n18481), .B2(n18486), .ZN(
        n18484) );
  OAI21_X1 U21542 ( .B1(n18485), .B2(n18486), .A(n18484), .ZN(P3_U2996) );
  NOR4_X1 U21543 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18605), .A3(n18486), 
        .A4(n18632), .ZN(n18493) );
  AOI211_X1 U21544 ( .C1(n18504), .C2(n18628), .A(n18487), .B(n18493), .ZN(
        n18488) );
  OAI221_X1 U21545 ( .B1(n18491), .B2(n18490), .C1(n18491), .C2(n18489), .A(
        n18488), .ZN(P3_U2997) );
  NOR2_X1 U21546 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18635) );
  INV_X1 U21547 ( .A(n18584), .ZN(n18492) );
  NOR4_X1 U21548 ( .A1(n18635), .A2(n18494), .A3(n18493), .A4(n18492), .ZN(
        P3_U2998) );
  AND2_X1 U21549 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18495), .ZN(
        P3_U2999) );
  AND2_X1 U21550 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18495), .ZN(
        P3_U3000) );
  AND2_X1 U21551 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18495), .ZN(
        P3_U3001) );
  AND2_X1 U21552 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18495), .ZN(
        P3_U3002) );
  AND2_X1 U21553 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18495), .ZN(
        P3_U3003) );
  AND2_X1 U21554 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18495), .ZN(
        P3_U3004) );
  AND2_X1 U21555 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18495), .ZN(
        P3_U3005) );
  AND2_X1 U21556 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18495), .ZN(
        P3_U3006) );
  AND2_X1 U21557 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18495), .ZN(
        P3_U3007) );
  INV_X1 U21558 ( .A(P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20784) );
  NOR2_X1 U21559 ( .A1(n20784), .A2(n18583), .ZN(P3_U3008) );
  AND2_X1 U21560 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18495), .ZN(
        P3_U3009) );
  AND2_X1 U21561 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18495), .ZN(
        P3_U3010) );
  AND2_X1 U21562 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18495), .ZN(
        P3_U3011) );
  AND2_X1 U21563 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18495), .ZN(
        P3_U3012) );
  AND2_X1 U21564 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18495), .ZN(
        P3_U3013) );
  AND2_X1 U21565 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18495), .ZN(
        P3_U3014) );
  AND2_X1 U21566 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18495), .ZN(
        P3_U3015) );
  AND2_X1 U21567 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18495), .ZN(
        P3_U3016) );
  AND2_X1 U21568 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18495), .ZN(
        P3_U3017) );
  AND2_X1 U21569 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18495), .ZN(
        P3_U3018) );
  AND2_X1 U21570 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18495), .ZN(
        P3_U3019) );
  AND2_X1 U21571 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18495), .ZN(
        P3_U3020) );
  INV_X1 U21572 ( .A(P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20767) );
  NOR2_X1 U21573 ( .A1(n20767), .A2(n18583), .ZN(P3_U3021) );
  AND2_X1 U21574 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18495), .ZN(P3_U3022) );
  AND2_X1 U21575 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18495), .ZN(P3_U3023) );
  AND2_X1 U21576 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18495), .ZN(P3_U3024) );
  AND2_X1 U21577 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18495), .ZN(P3_U3025) );
  INV_X1 U21578 ( .A(P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(n20758) );
  NOR2_X1 U21579 ( .A1(n20758), .A2(n18583), .ZN(P3_U3026) );
  AND2_X1 U21580 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18495), .ZN(P3_U3027) );
  AND2_X1 U21581 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18495), .ZN(P3_U3028) );
  OAI21_X1 U21582 ( .B1(n18496), .B2(n20595), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18497) );
  AOI22_X1 U21583 ( .A1(n18509), .A2(n18511), .B1(n18641), .B2(n18497), .ZN(
        n18498) );
  INV_X1 U21584 ( .A(NA), .ZN(n20592) );
  OR3_X1 U21585 ( .A1(n20592), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n18503) );
  OAI211_X1 U21586 ( .C1(n18499), .C2(n18632), .A(n18498), .B(n18503), .ZN(
        P3_U3029) );
  AOI21_X1 U21587 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(HOLD), .A(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18500) );
  AOI21_X1 U21588 ( .B1(HOLD), .B2(P3_STATE_REG_2__SCAN_IN), .A(n18500), .ZN(
        n18501) );
  AOI22_X1 U21589 ( .A1(n18504), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n18501), .ZN(n18502) );
  NAND2_X1 U21590 ( .A1(n18502), .A2(n18629), .ZN(P3_U3030) );
  AOI22_X1 U21591 ( .A1(n18504), .A2(P3_STATE_REG_1__SCAN_IN), .B1(n18509), 
        .B2(n18503), .ZN(n18510) );
  NOR2_X1 U21592 ( .A1(n18511), .A2(n20595), .ZN(n18507) );
  NAND2_X1 U21593 ( .A1(n18504), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18505) );
  OAI22_X1 U21594 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18505), .ZN(n18506) );
  OAI22_X1 U21595 ( .A1(n18507), .A2(n18506), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18508) );
  OAI22_X1 U21596 ( .A1(n18510), .A2(n18511), .B1(n18509), .B2(n18508), .ZN(
        P3_U3031) );
  NAND2_X1 U21597 ( .A1(n18640), .A2(n18511), .ZN(n18565) );
  OAI222_X1 U21598 ( .A1(n18614), .A2(n18575), .B1(n18512), .B2(n18640), .C1(
        n18514), .C2(n18571), .ZN(P3_U3032) );
  OAI222_X1 U21599 ( .A1(n18514), .A2(n18575), .B1(n18513), .B2(n18640), .C1(
        n18516), .C2(n18571), .ZN(P3_U3033) );
  OAI222_X1 U21600 ( .A1(n18516), .A2(n18575), .B1(n18515), .B2(n18640), .C1(
        n18518), .C2(n18571), .ZN(P3_U3034) );
  OAI222_X1 U21601 ( .A1(n18518), .A2(n18575), .B1(n18517), .B2(n18640), .C1(
        n18520), .C2(n18571), .ZN(P3_U3035) );
  OAI222_X1 U21602 ( .A1(n18520), .A2(n18575), .B1(n18519), .B2(n18640), .C1(
        n18521), .C2(n18571), .ZN(P3_U3036) );
  INV_X1 U21603 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18524) );
  OAI222_X1 U21604 ( .A1(n18565), .A2(n18524), .B1(n18522), .B2(n18640), .C1(
        n18521), .C2(n18568), .ZN(P3_U3037) );
  OAI222_X1 U21605 ( .A1(n18524), .A2(n18575), .B1(n18523), .B2(n18640), .C1(
        n18526), .C2(n18571), .ZN(P3_U3038) );
  OAI222_X1 U21606 ( .A1(n18526), .A2(n18575), .B1(n18525), .B2(n18640), .C1(
        n18528), .C2(n18565), .ZN(P3_U3039) );
  OAI222_X1 U21607 ( .A1(n18528), .A2(n18568), .B1(n18527), .B2(n18640), .C1(
        n18530), .C2(n18565), .ZN(P3_U3040) );
  OAI222_X1 U21608 ( .A1(n18530), .A2(n18568), .B1(n18529), .B2(n18640), .C1(
        n18532), .C2(n18571), .ZN(P3_U3041) );
  OAI222_X1 U21609 ( .A1(n18532), .A2(n18568), .B1(n18531), .B2(n18640), .C1(
        n18534), .C2(n18571), .ZN(P3_U3042) );
  OAI222_X1 U21610 ( .A1(n18534), .A2(n18568), .B1(n18533), .B2(n18640), .C1(
        n18535), .C2(n18571), .ZN(P3_U3043) );
  OAI222_X1 U21611 ( .A1(n18565), .A2(n18538), .B1(n18536), .B2(n18640), .C1(
        n18535), .C2(n18568), .ZN(P3_U3044) );
  OAI222_X1 U21612 ( .A1(n18538), .A2(n18568), .B1(n18537), .B2(n18640), .C1(
        n18540), .C2(n18571), .ZN(P3_U3045) );
  OAI222_X1 U21613 ( .A1(n18540), .A2(n18568), .B1(n18539), .B2(n18640), .C1(
        n18542), .C2(n18571), .ZN(P3_U3046) );
  OAI222_X1 U21614 ( .A1(n18542), .A2(n18568), .B1(n18541), .B2(n18640), .C1(
        n18544), .C2(n18571), .ZN(P3_U3047) );
  OAI222_X1 U21615 ( .A1(n18544), .A2(n18568), .B1(n18543), .B2(n18640), .C1(
        n18545), .C2(n18571), .ZN(P3_U3048) );
  OAI222_X1 U21616 ( .A1(n18565), .A2(n18547), .B1(n18546), .B2(n18640), .C1(
        n18545), .C2(n18568), .ZN(P3_U3049) );
  OAI222_X1 U21617 ( .A1(n18565), .A2(n18549), .B1(n18548), .B2(n18640), .C1(
        n18547), .C2(n18568), .ZN(P3_U3050) );
  OAI222_X1 U21618 ( .A1(n18565), .A2(n18552), .B1(n18550), .B2(n18640), .C1(
        n18549), .C2(n18568), .ZN(P3_U3051) );
  INV_X1 U21619 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18553) );
  OAI222_X1 U21620 ( .A1(n18552), .A2(n18568), .B1(n18551), .B2(n18640), .C1(
        n18553), .C2(n18571), .ZN(P3_U3052) );
  OAI222_X1 U21621 ( .A1(n18565), .A2(n18556), .B1(n18554), .B2(n18640), .C1(
        n18553), .C2(n18568), .ZN(P3_U3053) );
  OAI222_X1 U21622 ( .A1(n18556), .A2(n18575), .B1(n18555), .B2(n18640), .C1(
        n18557), .C2(n18571), .ZN(P3_U3054) );
  OAI222_X1 U21623 ( .A1(n18571), .A2(n18559), .B1(n18558), .B2(n18640), .C1(
        n18557), .C2(n18568), .ZN(P3_U3055) );
  INV_X1 U21624 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18561) );
  OAI222_X1 U21625 ( .A1(n18565), .A2(n18561), .B1(n18560), .B2(n18640), .C1(
        n18559), .C2(n18568), .ZN(P3_U3056) );
  OAI222_X1 U21626 ( .A1(n18571), .A2(n18563), .B1(n18562), .B2(n18640), .C1(
        n18561), .C2(n18568), .ZN(P3_U3057) );
  INV_X1 U21627 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18567) );
  OAI222_X1 U21628 ( .A1(n18565), .A2(n18567), .B1(n18564), .B2(n18640), .C1(
        n18563), .C2(n18568), .ZN(P3_U3058) );
  OAI222_X1 U21629 ( .A1(n18567), .A2(n18575), .B1(n18566), .B2(n18640), .C1(
        n18569), .C2(n18571), .ZN(P3_U3059) );
  OAI222_X1 U21630 ( .A1(n18571), .A2(n18574), .B1(n18570), .B2(n18640), .C1(
        n18569), .C2(n18568), .ZN(P3_U3060) );
  OAI222_X1 U21631 ( .A1(n18575), .A2(n18574), .B1(n18573), .B2(n18640), .C1(
        n18572), .C2(n18571), .ZN(P3_U3061) );
  OAI22_X1 U21632 ( .A1(n18641), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18640), .ZN(n18576) );
  INV_X1 U21633 ( .A(n18576), .ZN(P3_U3274) );
  OAI22_X1 U21634 ( .A1(n18641), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18640), .ZN(n18577) );
  INV_X1 U21635 ( .A(n18577), .ZN(P3_U3275) );
  OAI22_X1 U21636 ( .A1(n18641), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18640), .ZN(n18578) );
  INV_X1 U21637 ( .A(n18578), .ZN(P3_U3276) );
  OAI22_X1 U21638 ( .A1(n18641), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18640), .ZN(n18579) );
  INV_X1 U21639 ( .A(n18579), .ZN(P3_U3277) );
  OAI21_X1 U21640 ( .B1(n18583), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18581), 
        .ZN(n18580) );
  INV_X1 U21641 ( .A(n18580), .ZN(P3_U3280) );
  OAI21_X1 U21642 ( .B1(n18583), .B2(n18582), .A(n18581), .ZN(P3_U3281) );
  OAI221_X1 U21643 ( .B1(n18586), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18586), 
        .C2(n18585), .A(n18584), .ZN(P3_U3282) );
  INV_X1 U21644 ( .A(n18599), .ZN(n18609) );
  AOI22_X1 U21645 ( .A1(n18647), .A2(n18588), .B1(n18609), .B2(n18587), .ZN(
        n18589) );
  INV_X1 U21646 ( .A(n18613), .ZN(n18610) );
  AOI22_X1 U21647 ( .A1(n18613), .A2(n18590), .B1(n18589), .B2(n18610), .ZN(
        P3_U3285) );
  NAND2_X1 U21648 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18608) );
  INV_X1 U21649 ( .A(n18608), .ZN(n18596) );
  AOI22_X1 U21650 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n18591), .B2(n10903), .ZN(
        n18600) );
  OAI22_X1 U21651 ( .A1(n18594), .A2(n18593), .B1(n18599), .B2(n18592), .ZN(
        n18595) );
  AOI21_X1 U21652 ( .B1(n18596), .B2(n18600), .A(n18595), .ZN(n18597) );
  AOI22_X1 U21653 ( .A1(n18613), .A2(n11052), .B1(n18597), .B2(n18610), .ZN(
        P3_U3288) );
  OAI22_X1 U21654 ( .A1(n18600), .A2(n18608), .B1(n18599), .B2(n18598), .ZN(
        n18601) );
  AOI21_X1 U21655 ( .B1(n18647), .B2(n18602), .A(n18601), .ZN(n18603) );
  AOI22_X1 U21656 ( .A1(n18613), .A2(n18604), .B1(n18603), .B2(n18610), .ZN(
        P3_U3289) );
  OAI21_X1 U21657 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18606), .A(n18605), 
        .ZN(n18607) );
  AOI22_X1 U21658 ( .A1(n18609), .A2(n18612), .B1(n18608), .B2(n18607), .ZN(
        n18611) );
  AOI22_X1 U21659 ( .A1(n18613), .A2(n18612), .B1(n18611), .B2(n18610), .ZN(
        P3_U3290) );
  AOI21_X1 U21660 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18615) );
  AOI22_X1 U21661 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18615), .B2(n18614), .ZN(n18618) );
  INV_X1 U21662 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18617) );
  AOI22_X1 U21663 ( .A1(n18621), .A2(n18618), .B1(n18617), .B2(n18616), .ZN(
        P3_U3292) );
  INV_X1 U21664 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18620) );
  OAI21_X1 U21665 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18621), .ZN(n18619) );
  OAI21_X1 U21666 ( .B1(n18621), .B2(n18620), .A(n18619), .ZN(P3_U3293) );
  INV_X1 U21667 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18622) );
  AOI22_X1 U21668 ( .A1(n18640), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18622), 
        .B2(n18641), .ZN(P3_U3294) );
  MUX2_X1 U21669 ( .A(P3_MORE_REG_SCAN_IN), .B(n18624), .S(n18623), .Z(
        P3_U3295) );
  NOR2_X1 U21670 ( .A1(n18626), .A2(n18625), .ZN(n18627) );
  AOI211_X1 U21671 ( .C1(n18628), .C2(n18632), .A(n18627), .B(n18651), .ZN(
        n18639) );
  AOI21_X1 U21672 ( .B1(n18631), .B2(n18630), .A(n18629), .ZN(n18633) );
  OAI211_X1 U21673 ( .C1(n18634), .C2(n18633), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18632), .ZN(n18636) );
  AOI21_X1 U21674 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18636), .A(n18635), 
        .ZN(n18638) );
  NAND2_X1 U21675 ( .A1(n18639), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18637) );
  OAI21_X1 U21676 ( .B1(n18639), .B2(n18638), .A(n18637), .ZN(P3_U3296) );
  OAI22_X1 U21677 ( .A1(n18641), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18640), .ZN(n18642) );
  INV_X1 U21678 ( .A(n18642), .ZN(P3_U3297) );
  AOI21_X1 U21679 ( .B1(n18647), .B2(n18646), .A(P3_READREQUEST_REG_SCAN_IN), 
        .ZN(n18644) );
  AOI22_X1 U21680 ( .A1(n18651), .A2(n18645), .B1(n18644), .B2(n18643), .ZN(
        P3_U3298) );
  INV_X1 U21681 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18650) );
  NAND2_X1 U21682 ( .A1(n18647), .A2(n18646), .ZN(n18649) );
  OAI211_X1 U21683 ( .C1(n18651), .C2(n18650), .A(n18649), .B(n18648), .ZN(
        P3_U3299) );
  INV_X1 U21684 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19624) );
  NAND2_X1 U21685 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19624), .ZN(n19617) );
  OR2_X1 U21686 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19614) );
  OAI21_X1 U21687 ( .B1(n20805), .B2(n19617), .A(n19614), .ZN(n19673) );
  AOI21_X1 U21688 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19673), .ZN(n18652) );
  INV_X1 U21689 ( .A(n18652), .ZN(P2_U2815) );
  INV_X1 U21690 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18654) );
  OAI22_X1 U21691 ( .A1(n18653), .A2(n18654), .B1(n19685), .B2(n19602), .ZN(
        P2_U2816) );
  AOI22_X1 U21692 ( .A1(n19752), .A2(n18654), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n19753), .ZN(n18655) );
  OAI21_X1 U21693 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n19614), .A(n18655), 
        .ZN(P2_U2817) );
  OAI21_X1 U21694 ( .B1(n18656), .B2(BS16), .A(n19673), .ZN(n19671) );
  OAI21_X1 U21695 ( .B1(n19673), .B2(n19682), .A(n19671), .ZN(P2_U2818) );
  NOR2_X1 U21696 ( .A1(n18658), .A2(n18657), .ZN(n19730) );
  INV_X1 U21697 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n18660) );
  OAI21_X1 U21698 ( .B1(n19730), .B2(n18660), .A(n18659), .ZN(P2_U2819) );
  NOR4_X1 U21699 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18664) );
  NOR4_X1 U21700 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18663) );
  NOR4_X1 U21701 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18662) );
  NOR4_X1 U21702 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18661) );
  NAND4_X1 U21703 ( .A1(n18664), .A2(n18663), .A3(n18662), .A4(n18661), .ZN(
        n18670) );
  NOR4_X1 U21704 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18668) );
  AOI211_X1 U21705 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_29__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18667) );
  NOR4_X1 U21706 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18666) );
  NOR4_X1 U21707 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18665) );
  NAND4_X1 U21708 ( .A1(n18668), .A2(n18667), .A3(n18666), .A4(n18665), .ZN(
        n18669) );
  NOR2_X1 U21709 ( .A1(n18670), .A2(n18669), .ZN(n18681) );
  INV_X1 U21710 ( .A(n18681), .ZN(n18679) );
  NOR2_X1 U21711 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18679), .ZN(n18673) );
  INV_X1 U21712 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18671) );
  AOI22_X1 U21713 ( .A1(n18673), .A2(n18674), .B1(n18679), .B2(n18671), .ZN(
        P2_U2820) );
  OR3_X1 U21714 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18678) );
  INV_X1 U21715 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18672) );
  AOI22_X1 U21716 ( .A1(n18673), .A2(n18678), .B1(n18679), .B2(n18672), .ZN(
        P2_U2821) );
  INV_X1 U21717 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19672) );
  NAND2_X1 U21718 ( .A1(n18673), .A2(n19672), .ZN(n18677) );
  OAI21_X1 U21719 ( .B1(n10247), .B2(n18674), .A(n18681), .ZN(n18675) );
  OAI21_X1 U21720 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18681), .A(n18675), 
        .ZN(n18676) );
  OAI221_X1 U21721 ( .B1(n18677), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18677), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18676), .ZN(P2_U2822) );
  INV_X1 U21722 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18680) );
  OAI221_X1 U21723 ( .B1(n18681), .B2(n18680), .C1(n18679), .C2(n18678), .A(
        n18677), .ZN(P2_U2823) );
  NAND2_X1 U21724 ( .A1(n9828), .A2(n18682), .ZN(n18683) );
  XOR2_X1 U21725 ( .A(n18684), .B(n18683), .Z(n18693) );
  OAI21_X1 U21726 ( .B1(n19645), .B2(n18849), .A(n18831), .ZN(n18688) );
  OAI22_X1 U21727 ( .A1(n18686), .A2(n18888), .B1(n18874), .B2(n18685), .ZN(
        n18687) );
  AOI211_X1 U21728 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n18889), .A(n18688), .B(
        n18687), .ZN(n18692) );
  INV_X1 U21729 ( .A(n18689), .ZN(n18690) );
  AOI22_X1 U21730 ( .A1(n18690), .A2(n18896), .B1(n10069), .B2(n18877), .ZN(
        n18691) );
  OAI211_X1 U21731 ( .C1(n19606), .C2(n18693), .A(n18692), .B(n18691), .ZN(
        P2_U2836) );
  NOR2_X1 U21732 ( .A1(n18865), .A2(n18694), .ZN(n18696) );
  XOR2_X1 U21733 ( .A(n18696), .B(n18695), .Z(n18704) );
  AOI22_X1 U21734 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(n18889), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18901), .ZN(n18697) );
  OAI21_X1 U21735 ( .B1(n18698), .B2(n18888), .A(n18697), .ZN(n18699) );
  AOI211_X1 U21736 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n18890), .A(n19011), 
        .B(n18699), .ZN(n18703) );
  AOI22_X1 U21737 ( .A1(n18701), .A2(n18896), .B1(n18700), .B2(n18877), .ZN(
        n18702) );
  OAI211_X1 U21738 ( .C1(n19606), .C2(n18704), .A(n18703), .B(n18702), .ZN(
        P2_U2837) );
  NAND2_X1 U21739 ( .A1(n9828), .A2(n18705), .ZN(n18706) );
  XOR2_X1 U21740 ( .A(n18707), .B(n18706), .Z(n18717) );
  OAI21_X1 U21741 ( .B1(n19641), .B2(n18849), .A(n18847), .ZN(n18712) );
  INV_X1 U21742 ( .A(n18708), .ZN(n18710) );
  OAI22_X1 U21743 ( .A1(n18710), .A2(n18888), .B1(n18874), .B2(n18709), .ZN(
        n18711) );
  AOI211_X1 U21744 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n18889), .A(n18712), .B(
        n18711), .ZN(n18716) );
  AOI22_X1 U21745 ( .A1(n18714), .A2(n18877), .B1(n18713), .B2(n18896), .ZN(
        n18715) );
  OAI211_X1 U21746 ( .C1(n19606), .C2(n18717), .A(n18716), .B(n18715), .ZN(
        P2_U2838) );
  AOI22_X1 U21747 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n18901), .B1(
        P2_EBX_REG_16__SCAN_IN), .B2(n18889), .ZN(n18718) );
  OAI21_X1 U21748 ( .B1(n18719), .B2(n18888), .A(n18718), .ZN(n18720) );
  AOI211_X1 U21749 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n18890), .A(n19011), 
        .B(n18720), .ZN(n18726) );
  NOR2_X1 U21750 ( .A1(n18865), .A2(n18721), .ZN(n18723) );
  XNOR2_X1 U21751 ( .A(n18723), .B(n18722), .ZN(n18724) );
  AOI22_X1 U21752 ( .A1(n18912), .A2(n18877), .B1(n18882), .B2(n18724), .ZN(
        n18725) );
  OAI211_X1 U21753 ( .C1(n18727), .C2(n18871), .A(n18726), .B(n18725), .ZN(
        P2_U2839) );
  NAND2_X1 U21754 ( .A1(n9828), .A2(n18728), .ZN(n18730) );
  XOR2_X1 U21755 ( .A(n18730), .B(n18729), .Z(n18738) );
  AOI22_X1 U21756 ( .A1(n18731), .A2(n18876), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18901), .ZN(n18732) );
  OAI211_X1 U21757 ( .C1(n10456), .C2(n18849), .A(n18732), .B(n18847), .ZN(
        n18736) );
  INV_X1 U21758 ( .A(n18733), .ZN(n18734) );
  OAI22_X1 U21759 ( .A1(n18734), .A2(n18871), .B1(n18920), .B2(n18893), .ZN(
        n18735) );
  AOI211_X1 U21760 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n18889), .A(n18736), .B(
        n18735), .ZN(n18737) );
  OAI21_X1 U21761 ( .B1(n18738), .B2(n19606), .A(n18737), .ZN(P2_U2840) );
  NOR2_X1 U21762 ( .A1(n18865), .A2(n18746), .ZN(n18739) );
  NOR3_X1 U21763 ( .A1(n18739), .A2(n19606), .A3(n18747), .ZN(n18745) );
  NAND2_X1 U21764 ( .A1(n18740), .A2(n18876), .ZN(n18743) );
  AOI22_X1 U21765 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18901), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n18890), .ZN(n18742) );
  NAND2_X1 U21766 ( .A1(n18889), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n18741) );
  NAND4_X1 U21767 ( .A1(n18743), .A2(n18742), .A3(n18847), .A4(n18741), .ZN(
        n18744) );
  NOR2_X1 U21768 ( .A1(n18745), .A2(n18744), .ZN(n18750) );
  INV_X1 U21769 ( .A(n18923), .ZN(n18748) );
  NOR3_X1 U21770 ( .A1(n18865), .A2(n18746), .A3(n19606), .ZN(n18760) );
  AOI22_X1 U21771 ( .A1(n18877), .A2(n18748), .B1(n18760), .B2(n18747), .ZN(
        n18749) );
  OAI211_X1 U21772 ( .C1(n18751), .C2(n18871), .A(n18750), .B(n18749), .ZN(
        P2_U2841) );
  AOI22_X1 U21773 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n18901), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n18890), .ZN(n18752) );
  OAI211_X1 U21774 ( .C1(n18753), .C2(n18888), .A(n18752), .B(n18831), .ZN(
        n18754) );
  AOI21_X1 U21775 ( .B1(n18756), .B2(n18900), .A(n18754), .ZN(n18762) );
  NAND2_X1 U21776 ( .A1(n18756), .A2(n18755), .ZN(n18759) );
  OAI22_X1 U21777 ( .A1(n18757), .A2(n18871), .B1(n18925), .B2(n18893), .ZN(
        n18758) );
  AOI21_X1 U21778 ( .B1(n18760), .B2(n18759), .A(n18758), .ZN(n18761) );
  OAI211_X1 U21779 ( .C1(n18857), .C2(n10779), .A(n18762), .B(n18761), .ZN(
        P2_U2842) );
  AOI22_X1 U21780 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18901), .B1(
        P2_EBX_REG_12__SCAN_IN), .B2(n18889), .ZN(n18763) );
  OAI21_X1 U21781 ( .B1(n18764), .B2(n18888), .A(n18763), .ZN(n18765) );
  AOI211_X1 U21782 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n18890), .A(n19011), 
        .B(n18765), .ZN(n18771) );
  INV_X1 U21783 ( .A(n18928), .ZN(n18769) );
  NOR2_X1 U21784 ( .A1(n18865), .A2(n18779), .ZN(n18767) );
  XNOR2_X1 U21785 ( .A(n18767), .B(n18766), .ZN(n18768) );
  AOI22_X1 U21786 ( .A1(n18769), .A2(n18877), .B1(n18882), .B2(n18768), .ZN(
        n18770) );
  OAI211_X1 U21787 ( .C1(n18772), .C2(n18871), .A(n18771), .B(n18770), .ZN(
        P2_U2843) );
  INV_X1 U21788 ( .A(n18773), .ZN(n18785) );
  AOI22_X1 U21789 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18901), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n18890), .ZN(n18774) );
  OAI211_X1 U21790 ( .C1(n18930), .C2(n18893), .A(n18774), .B(n18847), .ZN(
        n18778) );
  INV_X1 U21791 ( .A(n18775), .ZN(n18776) );
  OAI22_X1 U21792 ( .A1(n18776), .A2(n18888), .B1(n18857), .B2(n10001), .ZN(
        n18777) );
  AOI211_X1 U21793 ( .C1(n18780), .C2(n18900), .A(n18778), .B(n18777), .ZN(
        n18784) );
  AOI21_X1 U21794 ( .B1(n18781), .B2(n18780), .A(n18779), .ZN(n18782) );
  NAND2_X1 U21795 ( .A1(n18899), .A2(n18782), .ZN(n18783) );
  OAI211_X1 U21796 ( .C1(n18871), .C2(n18785), .A(n18784), .B(n18783), .ZN(
        P2_U2844) );
  NOR2_X1 U21797 ( .A1(n18865), .A2(n18786), .ZN(n18787) );
  XOR2_X1 U21798 ( .A(n18788), .B(n18787), .Z(n18797) );
  INV_X1 U21799 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18789) );
  OAI22_X1 U21800 ( .A1(n18790), .A2(n18888), .B1(n18874), .B2(n18789), .ZN(
        n18791) );
  INV_X1 U21801 ( .A(n18791), .ZN(n18792) );
  OAI211_X1 U21802 ( .C1(n10659), .C2(n18849), .A(n18792), .B(n18847), .ZN(
        n18795) );
  OAI22_X1 U21803 ( .A1(n18793), .A2(n18871), .B1(n18933), .B2(n18893), .ZN(
        n18794) );
  AOI211_X1 U21804 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n18889), .A(n18795), .B(
        n18794), .ZN(n18796) );
  OAI21_X1 U21805 ( .B1(n19606), .B2(n18797), .A(n18796), .ZN(P2_U2845) );
  OAI21_X1 U21806 ( .B1(n10638), .B2(n18849), .A(n18847), .ZN(n18801) );
  INV_X1 U21807 ( .A(n18798), .ZN(n18799) );
  OAI22_X1 U21808 ( .A1(n18799), .A2(n18888), .B1(n18857), .B2(n10777), .ZN(
        n18800) );
  AOI211_X1 U21809 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n18901), .A(
        n18801), .B(n18800), .ZN(n18808) );
  NAND2_X1 U21810 ( .A1(n9828), .A2(n18802), .ZN(n18803) );
  XNOR2_X1 U21811 ( .A(n18804), .B(n18803), .ZN(n18805) );
  AOI22_X1 U21812 ( .A1(n18806), .A2(n18896), .B1(n18882), .B2(n18805), .ZN(
        n18807) );
  OAI211_X1 U21813 ( .C1(n18936), .C2(n18893), .A(n18808), .B(n18807), .ZN(
        P2_U2846) );
  AOI22_X1 U21814 ( .A1(n18809), .A2(n18876), .B1(P2_EBX_REG_8__SCAN_IN), .B2(
        n18889), .ZN(n18810) );
  OAI211_X1 U21815 ( .C1(n10620), .C2(n18849), .A(n18810), .B(n18831), .ZN(
        n18811) );
  AOI21_X1 U21816 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18901), .A(
        n18811), .ZN(n18818) );
  NOR2_X1 U21817 ( .A1(n18865), .A2(n18812), .ZN(n18814) );
  XNOR2_X1 U21818 ( .A(n18814), .B(n18813), .ZN(n18816) );
  INV_X1 U21819 ( .A(n18940), .ZN(n18815) );
  AOI22_X1 U21820 ( .A1(n18882), .A2(n18816), .B1(n18877), .B2(n18815), .ZN(
        n18817) );
  OAI211_X1 U21821 ( .C1(n18871), .C2(n18819), .A(n18818), .B(n18817), .ZN(
        P2_U2847) );
  NAND2_X1 U21822 ( .A1(n9828), .A2(n18820), .ZN(n18822) );
  XOR2_X1 U21823 ( .A(n18822), .B(n18821), .Z(n18829) );
  AOI22_X1 U21824 ( .A1(n18823), .A2(n18876), .B1(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18901), .ZN(n18824) );
  OAI211_X1 U21825 ( .C1(n10335), .C2(n18849), .A(n18824), .B(n18847), .ZN(
        n18827) );
  OAI22_X1 U21826 ( .A1(n18893), .A2(n18941), .B1(n18871), .B2(n18825), .ZN(
        n18826) );
  AOI211_X1 U21827 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n18889), .A(n18827), .B(
        n18826), .ZN(n18828) );
  OAI21_X1 U21828 ( .B1(n18829), .B2(n19606), .A(n18828), .ZN(P2_U2848) );
  INV_X1 U21829 ( .A(n18830), .ZN(n18834) );
  AOI22_X1 U21830 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18901), .B1(
        P2_EBX_REG_6__SCAN_IN), .B2(n18889), .ZN(n18832) );
  OAI211_X1 U21831 ( .C1(n18849), .C2(n10332), .A(n18832), .B(n18831), .ZN(
        n18833) );
  AOI21_X1 U21832 ( .B1(n18834), .B2(n18876), .A(n18833), .ZN(n18840) );
  NOR2_X1 U21833 ( .A1(n18865), .A2(n18835), .ZN(n18837) );
  XNOR2_X1 U21834 ( .A(n18837), .B(n18836), .ZN(n18838) );
  AOI22_X1 U21835 ( .A1(n18882), .A2(n18838), .B1(n18877), .B2(n18942), .ZN(
        n18839) );
  OAI211_X1 U21836 ( .C1(n18871), .C2(n18841), .A(n18840), .B(n18839), .ZN(
        P2_U2849) );
  NAND2_X1 U21837 ( .A1(n9828), .A2(n18842), .ZN(n18844) );
  XOR2_X1 U21838 ( .A(n18844), .B(n18843), .Z(n18854) );
  INV_X1 U21839 ( .A(n18845), .ZN(n18846) );
  AOI22_X1 U21840 ( .A1(n18846), .A2(n18876), .B1(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18901), .ZN(n18848) );
  OAI211_X1 U21841 ( .C1(n10328), .C2(n18849), .A(n18848), .B(n18847), .ZN(
        n18852) );
  OAI22_X1 U21842 ( .A1(n18893), .A2(n18950), .B1(n18871), .B2(n18850), .ZN(
        n18851) );
  AOI211_X1 U21843 ( .C1(P2_EBX_REG_5__SCAN_IN), .C2(n18889), .A(n18852), .B(
        n18851), .ZN(n18853) );
  OAI21_X1 U21844 ( .B1(n18854), .B2(n19606), .A(n18853), .ZN(P2_U2850) );
  INV_X1 U21845 ( .A(n18855), .ZN(n18946) );
  NOR2_X1 U21846 ( .A1(n18857), .A2(n18856), .ZN(n18858) );
  AOI211_X1 U21847 ( .C1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n18901), .A(
        n19011), .B(n18858), .ZN(n18861) );
  AOI22_X1 U21848 ( .A1(n18877), .A2(n18859), .B1(n18890), .B2(
        P2_REIP_REG_4__SCAN_IN), .ZN(n18860) );
  OAI211_X1 U21849 ( .C1(n18862), .C2(n18888), .A(n18861), .B(n18860), .ZN(
        n18863) );
  AOI21_X1 U21850 ( .B1(n18946), .B2(n18897), .A(n18863), .ZN(n18870) );
  INV_X1 U21851 ( .A(n19024), .ZN(n18868) );
  NOR2_X1 U21852 ( .A1(n18865), .A2(n18864), .ZN(n18867) );
  AOI21_X1 U21853 ( .B1(n18868), .B2(n18867), .A(n19606), .ZN(n18866) );
  OAI21_X1 U21854 ( .B1(n18868), .B2(n18867), .A(n18866), .ZN(n18869) );
  OAI211_X1 U21855 ( .C1(n19019), .C2(n18871), .A(n18870), .B(n18869), .ZN(
        P2_U2851) );
  NAND2_X1 U21856 ( .A1(n18872), .A2(n18896), .ZN(n18881) );
  NOR2_X1 U21857 ( .A1(n18874), .A2(n18873), .ZN(n18875) );
  AOI21_X1 U21858 ( .B1(n18889), .B2(P2_EBX_REG_1__SCAN_IN), .A(n18875), .ZN(
        n18880) );
  AOI22_X1 U21859 ( .A1(n18876), .A2(n10079), .B1(n18890), .B2(
        P2_REIP_REG_1__SCAN_IN), .ZN(n18879) );
  NAND2_X1 U21860 ( .A1(n19708), .A2(n18877), .ZN(n18878) );
  AND4_X1 U21861 ( .A1(n18881), .A2(n18880), .A3(n18879), .A4(n18878), .ZN(
        n18885) );
  AOI22_X1 U21862 ( .A1(n18883), .A2(n18882), .B1(n18897), .B2(n19706), .ZN(
        n18884) );
  OAI211_X1 U21863 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n18886), .A(
        n18885), .B(n18884), .ZN(P2_U2854) );
  NOR2_X1 U21864 ( .A1(n18888), .A2(n18887), .ZN(n18895) );
  AOI22_X1 U21865 ( .A1(n18890), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n18889), 
        .B2(P2_EBX_REG_0__SCAN_IN), .ZN(n18891) );
  OAI21_X1 U21866 ( .B1(n18893), .B2(n18892), .A(n18891), .ZN(n18894) );
  AOI211_X1 U21867 ( .C1(n18896), .C2(n12601), .A(n18895), .B(n18894), .ZN(
        n18904) );
  AOI22_X1 U21868 ( .A1(n18899), .A2(n18898), .B1(n19303), .B2(n18897), .ZN(
        n18903) );
  OAI21_X1 U21869 ( .B1(n18901), .B2(n18900), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18902) );
  NAND3_X1 U21870 ( .A1(n18904), .A2(n18903), .A3(n18902), .ZN(P2_U2855) );
  AOI22_X1 U21871 ( .A1(n18905), .A2(n18964), .B1(n18911), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n18907) );
  AOI22_X1 U21872 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n18963), .B1(n18910), 
        .B2(BUF2_REG_31__SCAN_IN), .ZN(n18906) );
  NAND2_X1 U21873 ( .A1(n18907), .A2(n18906), .ZN(P2_U2888) );
  INV_X1 U21874 ( .A(n19033), .ZN(n18908) );
  AOI22_X1 U21875 ( .A1(n18909), .A2(n18908), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n18963), .ZN(n18918) );
  AOI22_X1 U21876 ( .A1(n18911), .A2(BUF1_REG_16__SCAN_IN), .B1(n18910), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n18917) );
  INV_X1 U21877 ( .A(n18912), .ZN(n18913) );
  OAI22_X1 U21878 ( .A1(n18914), .A2(n18968), .B1(n18954), .B2(n18913), .ZN(
        n18915) );
  INV_X1 U21879 ( .A(n18915), .ZN(n18916) );
  NAND3_X1 U21880 ( .A1(n18918), .A2(n18917), .A3(n18916), .ZN(P2_U2903) );
  OAI222_X1 U21881 ( .A1(n18920), .A2(n18951), .B1(n13041), .B2(n18953), .C1(
        n18919), .C2(n18972), .ZN(P2_U2904) );
  AOI22_X1 U21882 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n18963), .B1(n18921), 
        .B2(n18937), .ZN(n18922) );
  OAI21_X1 U21883 ( .B1(n18951), .B2(n18923), .A(n18922), .ZN(P2_U2905) );
  INV_X1 U21884 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n18983) );
  OAI222_X1 U21885 ( .A1(n18925), .A2(n18951), .B1(n18983), .B2(n18953), .C1(
        n18972), .C2(n18924), .ZN(P2_U2906) );
  AOI22_X1 U21886 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n18963), .B1(n18926), 
        .B2(n18937), .ZN(n18927) );
  OAI21_X1 U21887 ( .B1(n18951), .B2(n18928), .A(n18927), .ZN(P2_U2907) );
  INV_X1 U21888 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n18987) );
  OAI222_X1 U21889 ( .A1(n18930), .A2(n18951), .B1(n18987), .B2(n18953), .C1(
        n18972), .C2(n18929), .ZN(P2_U2908) );
  AOI22_X1 U21890 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n18963), .B1(n18931), 
        .B2(n18937), .ZN(n18932) );
  OAI21_X1 U21891 ( .B1(n18951), .B2(n18933), .A(n18932), .ZN(P2_U2909) );
  INV_X1 U21892 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n18935) );
  OAI222_X1 U21893 ( .A1(n18936), .A2(n18951), .B1(n18935), .B2(n18953), .C1(
        n18972), .C2(n18934), .ZN(P2_U2910) );
  AOI22_X1 U21894 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n18963), .B1(n18938), .B2(
        n18937), .ZN(n18939) );
  OAI21_X1 U21895 ( .B1(n18951), .B2(n18940), .A(n18939), .ZN(P2_U2911) );
  INV_X1 U21896 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n18995) );
  OAI222_X1 U21897 ( .A1(n18941), .A2(n18951), .B1(n18995), .B2(n18953), .C1(
        n18972), .C2(n19069), .ZN(P2_U2912) );
  INV_X1 U21898 ( .A(n18942), .ZN(n18943) );
  INV_X1 U21899 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n18997) );
  OAI222_X1 U21900 ( .A1(n18943), .A2(n18951), .B1(n18997), .B2(n18953), .C1(
        n18972), .C2(n19058), .ZN(P2_U2913) );
  INV_X1 U21901 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n18999) );
  OAI22_X1 U21902 ( .A1(n18999), .A2(n18953), .B1(n19053), .B2(n18972), .ZN(
        n18944) );
  INV_X1 U21903 ( .A(n18944), .ZN(n18949) );
  NAND3_X1 U21904 ( .A1(n18947), .A2(n18946), .A3(n18945), .ZN(n18948) );
  OAI211_X1 U21905 ( .C1(n18951), .C2(n18950), .A(n18949), .B(n18948), .ZN(
        P2_U2914) );
  INV_X1 U21906 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n18952) );
  OAI22_X1 U21907 ( .A1(n18955), .A2(n18954), .B1(n18953), .B2(n18952), .ZN(
        n18956) );
  INV_X1 U21908 ( .A(n18956), .ZN(n18962) );
  AOI21_X1 U21909 ( .B1(n18959), .B2(n18958), .A(n18957), .ZN(n18960) );
  OR2_X1 U21910 ( .A1(n18960), .A2(n18968), .ZN(n18961) );
  OAI211_X1 U21911 ( .C1(n19046), .C2(n18972), .A(n18962), .B(n18961), .ZN(
        P2_U2916) );
  AOI22_X1 U21912 ( .A1(n18964), .A2(n19708), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n18963), .ZN(n18971) );
  AOI21_X1 U21913 ( .B1(n18967), .B2(n18966), .A(n18965), .ZN(n18969) );
  OR2_X1 U21914 ( .A1(n18969), .A2(n18968), .ZN(n18970) );
  OAI211_X1 U21915 ( .C1(n18973), .C2(n18972), .A(n18971), .B(n18970), .ZN(
        P2_U2918) );
  NOR2_X1 U21916 ( .A1(n18978), .A2(n18974), .ZN(P2_U2920) );
  INV_X1 U21917 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n20787) );
  INV_X1 U21918 ( .A(n18975), .ZN(n18976) );
  AOI22_X1 U21919 ( .A1(n18976), .A2(P2_EAX_REG_18__SCAN_IN), .B1(
        P2_UWORD_REG_2__SCAN_IN), .B2(n19008), .ZN(n18977) );
  OAI21_X1 U21920 ( .B1(n20787), .B2(n18978), .A(n18977), .ZN(P2_U2933) );
  AOI22_X1 U21921 ( .A1(n19008), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n18979) );
  OAI21_X1 U21922 ( .B1(n13041), .B2(n19010), .A(n18979), .ZN(P2_U2936) );
  AOI22_X1 U21923 ( .A1(n19008), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n18980) );
  OAI21_X1 U21924 ( .B1(n18981), .B2(n19010), .A(n18980), .ZN(P2_U2937) );
  AOI22_X1 U21925 ( .A1(n19008), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n18982) );
  OAI21_X1 U21926 ( .B1(n18983), .B2(n19010), .A(n18982), .ZN(P2_U2938) );
  AOI22_X1 U21927 ( .A1(n19008), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n18984) );
  OAI21_X1 U21928 ( .B1(n18985), .B2(n19010), .A(n18984), .ZN(P2_U2939) );
  AOI22_X1 U21929 ( .A1(n19008), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n18986) );
  OAI21_X1 U21930 ( .B1(n18987), .B2(n19010), .A(n18986), .ZN(P2_U2940) );
  AOI22_X1 U21931 ( .A1(n19008), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n18988) );
  OAI21_X1 U21932 ( .B1(n18989), .B2(n19010), .A(n18988), .ZN(P2_U2941) );
  AOI222_X1 U21933 ( .A1(n19007), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n18990), 
        .B2(P2_EAX_REG_9__SCAN_IN), .C1(n19008), .C2(P2_LWORD_REG_9__SCAN_IN), 
        .ZN(n18991) );
  INV_X1 U21934 ( .A(n18991), .ZN(P2_U2942) );
  AOI22_X1 U21935 ( .A1(n19008), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n18992) );
  OAI21_X1 U21936 ( .B1(n18993), .B2(n19010), .A(n18992), .ZN(P2_U2943) );
  AOI22_X1 U21937 ( .A1(n19008), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n18994) );
  OAI21_X1 U21938 ( .B1(n18995), .B2(n19010), .A(n18994), .ZN(P2_U2944) );
  AOI22_X1 U21939 ( .A1(n19008), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n18996) );
  OAI21_X1 U21940 ( .B1(n18997), .B2(n19010), .A(n18996), .ZN(P2_U2945) );
  AOI22_X1 U21941 ( .A1(n19008), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n18998) );
  OAI21_X1 U21942 ( .B1(n18999), .B2(n19010), .A(n18998), .ZN(P2_U2946) );
  INV_X1 U21943 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19001) );
  AOI22_X1 U21944 ( .A1(n19008), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19000) );
  OAI21_X1 U21945 ( .B1(n19001), .B2(n19010), .A(n19000), .ZN(P2_U2947) );
  AOI22_X1 U21946 ( .A1(n19008), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19002) );
  OAI21_X1 U21947 ( .B1(n18952), .B2(n19010), .A(n19002), .ZN(P2_U2948) );
  INV_X1 U21948 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19004) );
  AOI22_X1 U21949 ( .A1(n19008), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19003) );
  OAI21_X1 U21950 ( .B1(n19004), .B2(n19010), .A(n19003), .ZN(P2_U2949) );
  INV_X1 U21951 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19006) );
  AOI22_X1 U21952 ( .A1(n19008), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19005) );
  OAI21_X1 U21953 ( .B1(n19006), .B2(n19010), .A(n19005), .ZN(P2_U2950) );
  AOI22_X1 U21954 ( .A1(n19008), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19007), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19009) );
  OAI21_X1 U21955 ( .B1(n13039), .B2(n19010), .A(n19009), .ZN(P2_U2951) );
  AOI22_X1 U21956 ( .A1(n19012), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19011), .ZN(n19023) );
  NAND3_X1 U21957 ( .A1(n19014), .A2(n19013), .A3(n13839), .ZN(n19018) );
  NAND2_X1 U21958 ( .A1(n19016), .A2(n19015), .ZN(n19017) );
  OAI211_X1 U21959 ( .C1(n19020), .C2(n19019), .A(n19018), .B(n19017), .ZN(
        n19021) );
  INV_X1 U21960 ( .A(n19021), .ZN(n19022) );
  OAI211_X1 U21961 ( .C1(n19025), .C2(n19024), .A(n19023), .B(n19022), .ZN(
        P2_U3010) );
  AOI22_X1 U21962 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19062), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19061), .ZN(n19511) );
  AOI22_X1 U21963 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19062), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19061), .ZN(n19550) );
  NOR2_X2 U21964 ( .A1(n19027), .A2(n19049), .ZN(n19539) );
  NAND2_X1 U21965 ( .A1(n19693), .A2(n19700), .ZN(n19157) );
  NOR2_X1 U21966 ( .A1(n19306), .A2(n19157), .ZN(n19068) );
  AOI22_X1 U21967 ( .A1(n19592), .A2(n19499), .B1(n19539), .B2(n19068), .ZN(
        n19039) );
  OAI21_X1 U21968 ( .B1(n19592), .B2(n19124), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19028) );
  NAND2_X1 U21969 ( .A1(n19028), .A2(n19688), .ZN(n19037) );
  INV_X1 U21970 ( .A(n19534), .ZN(n19588) );
  NOR2_X1 U21971 ( .A1(n19037), .A2(n19588), .ZN(n19031) );
  OAI21_X1 U21972 ( .B1(n12290), .B2(n19733), .A(n19732), .ZN(n19030) );
  INV_X1 U21973 ( .A(n19068), .ZN(n19029) );
  OAI21_X1 U21974 ( .B1(n19031), .B2(n19030), .A(n19029), .ZN(n19032) );
  NAND2_X1 U21975 ( .A1(n19032), .A2(n19544), .ZN(n19071) );
  NOR2_X1 U21976 ( .A1(n19588), .A2(n19068), .ZN(n19036) );
  OAI21_X1 U21977 ( .B1(n12290), .B2(n19068), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19035) );
  AOI22_X1 U21978 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19071), .B1(
        n19034), .B2(n19070), .ZN(n19038) );
  OAI211_X1 U21979 ( .C1(n19511), .C2(n19103), .A(n19039), .B(n19038), .ZN(
        P2_U3048) );
  AOI22_X1 U21980 ( .A1(n19592), .A2(n19438), .B1(n19551), .B2(n19068), .ZN(
        n19041) );
  AOI22_X1 U21981 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19071), .B1(
        n19552), .B2(n19070), .ZN(n19040) );
  OAI211_X1 U21982 ( .C1(n19441), .C2(n19103), .A(n19041), .B(n19040), .ZN(
        P2_U3049) );
  AOI22_X1 U21983 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19062), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19061), .ZN(n19445) );
  AOI22_X1 U21984 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19061), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19062), .ZN(n19562) );
  NOR2_X2 U21985 ( .A1(n12515), .A2(n19049), .ZN(n19557) );
  AOI22_X1 U21986 ( .A1(n19592), .A2(n19442), .B1(n19557), .B2(n19068), .ZN(
        n19044) );
  NOR2_X2 U21987 ( .A1(n19042), .A2(n19338), .ZN(n19558) );
  AOI22_X1 U21988 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19071), .B1(
        n19558), .B2(n19070), .ZN(n19043) );
  OAI211_X1 U21989 ( .C1(n19445), .C2(n19103), .A(n19044), .B(n19043), .ZN(
        P2_U3050) );
  AOI22_X1 U21990 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19062), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19061), .ZN(n19449) );
  AOI22_X1 U21991 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19062), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19061), .ZN(n19568) );
  AND2_X1 U21992 ( .A1(n19045), .A2(n19067), .ZN(n19563) );
  AOI22_X1 U21993 ( .A1(n19592), .A2(n19446), .B1(n19563), .B2(n19068), .ZN(
        n19048) );
  NOR2_X2 U21994 ( .A1(n19046), .A2(n19338), .ZN(n19564) );
  AOI22_X1 U21995 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19071), .B1(
        n19564), .B2(n19070), .ZN(n19047) );
  OAI211_X1 U21996 ( .C1(n19449), .C2(n19103), .A(n19048), .B(n19047), .ZN(
        P2_U3051) );
  AOI22_X1 U21997 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19062), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19061), .ZN(n19453) );
  AOI22_X1 U21998 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19061), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19062), .ZN(n19574) );
  NOR2_X2 U21999 ( .A1(n10259), .A2(n19049), .ZN(n19569) );
  AOI22_X1 U22000 ( .A1(n19592), .A2(n19450), .B1(n19569), .B2(n19068), .ZN(
        n19052) );
  NOR2_X2 U22001 ( .A1(n19050), .A2(n19338), .ZN(n19570) );
  AOI22_X1 U22002 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19071), .B1(
        n19570), .B2(n19070), .ZN(n19051) );
  OAI211_X1 U22003 ( .C1(n19453), .C2(n19103), .A(n19052), .B(n19051), .ZN(
        P2_U3052) );
  AOI22_X1 U22004 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19062), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19061), .ZN(n19524) );
  AOI22_X1 U22005 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19062), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19061), .ZN(n19580) );
  AOI22_X1 U22006 ( .A1(n19592), .A2(n19520), .B1(n19575), .B2(n19068), .ZN(
        n19055) );
  NOR2_X2 U22007 ( .A1(n19053), .A2(n19338), .ZN(n19576) );
  AOI22_X1 U22008 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19071), .B1(
        n19576), .B2(n19070), .ZN(n19054) );
  OAI211_X1 U22009 ( .C1(n19524), .C2(n19103), .A(n19055), .B(n19054), .ZN(
        P2_U3053) );
  INV_X1 U22010 ( .A(n19062), .ZN(n19065) );
  INV_X1 U22011 ( .A(n19061), .ZN(n19063) );
  AOI22_X1 U22012 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19062), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19061), .ZN(n19586) );
  AOI22_X1 U22013 ( .A1(n19592), .A2(n19456), .B1(n19581), .B2(n19068), .ZN(
        n19060) );
  NOR2_X2 U22014 ( .A1(n19058), .A2(n19338), .ZN(n19582) );
  AOI22_X1 U22015 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19071), .B1(
        n19582), .B2(n19070), .ZN(n19059) );
  OAI211_X1 U22016 ( .C1(n19459), .C2(n19103), .A(n19060), .B(n19059), .ZN(
        P2_U3054) );
  AOI22_X1 U22017 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19062), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19061), .ZN(n19467) );
  AND2_X1 U22018 ( .A1(n10271), .A2(n19067), .ZN(n19587) );
  AOI22_X1 U22019 ( .A1(n19462), .A2(n19592), .B1(n19587), .B2(n19068), .ZN(
        n19073) );
  NOR2_X2 U22020 ( .A1(n19069), .A2(n19338), .ZN(n19589) );
  AOI22_X1 U22021 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19071), .B1(
        n19589), .B2(n19070), .ZN(n19072) );
  OAI211_X1 U22022 ( .C1(n19467), .C2(n19103), .A(n19073), .B(n19072), .ZN(
        P2_U3055) );
  NOR3_X1 U22023 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19720), .A3(
        n19157), .ZN(n19085) );
  INV_X1 U22024 ( .A(n19085), .ZN(n19119) );
  NAND2_X1 U22025 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19119), .ZN(n19074) );
  NOR2_X1 U22026 ( .A1(n12289), .A2(n19074), .ZN(n19081) );
  OR2_X1 U22027 ( .A1(n19157), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19082) );
  INV_X1 U22028 ( .A(n19082), .ZN(n19075) );
  AOI21_X1 U22029 ( .B1(n19732), .B2(n19075), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19076) );
  INV_X1 U22030 ( .A(n19034), .ZN(n19078) );
  INV_X1 U22031 ( .A(n19539), .ZN(n19077) );
  OAI22_X1 U22032 ( .A1(n19122), .A2(n19078), .B1(n19077), .B2(n19119), .ZN(
        n19079) );
  INV_X1 U22033 ( .A(n19079), .ZN(n19087) );
  NAND2_X1 U22034 ( .A1(n19304), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19268) );
  INV_X1 U22035 ( .A(n19268), .ZN(n19080) );
  NAND2_X1 U22036 ( .A1(n19080), .A2(n19305), .ZN(n19083) );
  AOI21_X1 U22037 ( .B1(n19083), .B2(n19082), .A(n19081), .ZN(n19084) );
  OAI211_X1 U22038 ( .C1(n19085), .C2(n19732), .A(n19084), .B(n19544), .ZN(
        n19125) );
  INV_X1 U22039 ( .A(n19511), .ZN(n19547) );
  AOI22_X1 U22040 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19125), .B1(
        n19153), .B2(n19547), .ZN(n19086) );
  OAI211_X1 U22041 ( .C1(n19550), .C2(n19103), .A(n19087), .B(n19086), .ZN(
        P2_U3056) );
  INV_X1 U22042 ( .A(n19552), .ZN(n19089) );
  INV_X1 U22043 ( .A(n19551), .ZN(n19088) );
  OAI22_X1 U22044 ( .A1(n19122), .A2(n19089), .B1(n19088), .B2(n19119), .ZN(
        n19090) );
  INV_X1 U22045 ( .A(n19090), .ZN(n19092) );
  AOI22_X1 U22046 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19125), .B1(
        n19124), .B2(n19438), .ZN(n19091) );
  OAI211_X1 U22047 ( .C1(n19441), .C2(n19130), .A(n19092), .B(n19091), .ZN(
        P2_U3057) );
  INV_X1 U22048 ( .A(n19558), .ZN(n19094) );
  INV_X1 U22049 ( .A(n19557), .ZN(n19093) );
  OAI22_X1 U22050 ( .A1(n19122), .A2(n19094), .B1(n19093), .B2(n19119), .ZN(
        n19095) );
  INV_X1 U22051 ( .A(n19095), .ZN(n19097) );
  AOI22_X1 U22052 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19125), .B1(
        n19124), .B2(n19442), .ZN(n19096) );
  OAI211_X1 U22053 ( .C1(n19445), .C2(n19130), .A(n19097), .B(n19096), .ZN(
        P2_U3058) );
  INV_X1 U22054 ( .A(n19564), .ZN(n19099) );
  INV_X1 U22055 ( .A(n19563), .ZN(n19098) );
  OAI22_X1 U22056 ( .A1(n19122), .A2(n19099), .B1(n19098), .B2(n19119), .ZN(
        n19100) );
  INV_X1 U22057 ( .A(n19100), .ZN(n19102) );
  INV_X1 U22058 ( .A(n19449), .ZN(n19565) );
  AOI22_X1 U22059 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19125), .B1(
        n19153), .B2(n19565), .ZN(n19101) );
  OAI211_X1 U22060 ( .C1(n19568), .C2(n19103), .A(n19102), .B(n19101), .ZN(
        P2_U3059) );
  INV_X1 U22061 ( .A(n19570), .ZN(n19105) );
  INV_X1 U22062 ( .A(n19569), .ZN(n19104) );
  OAI22_X1 U22063 ( .A1(n19122), .A2(n19105), .B1(n19104), .B2(n19119), .ZN(
        n19106) );
  INV_X1 U22064 ( .A(n19106), .ZN(n19108) );
  AOI22_X1 U22065 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19125), .B1(
        n19124), .B2(n19450), .ZN(n19107) );
  OAI211_X1 U22066 ( .C1(n19453), .C2(n19130), .A(n19108), .B(n19107), .ZN(
        P2_U3060) );
  INV_X1 U22067 ( .A(n19576), .ZN(n19110) );
  INV_X1 U22068 ( .A(n19575), .ZN(n19109) );
  OAI22_X1 U22069 ( .A1(n19122), .A2(n19110), .B1(n19109), .B2(n19119), .ZN(
        n19111) );
  INV_X1 U22070 ( .A(n19111), .ZN(n19113) );
  AOI22_X1 U22071 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19125), .B1(
        n19124), .B2(n19520), .ZN(n19112) );
  OAI211_X1 U22072 ( .C1(n19524), .C2(n19130), .A(n19113), .B(n19112), .ZN(
        P2_U3061) );
  INV_X1 U22073 ( .A(n19582), .ZN(n19115) );
  INV_X1 U22074 ( .A(n19581), .ZN(n19114) );
  OAI22_X1 U22075 ( .A1(n19122), .A2(n19115), .B1(n19114), .B2(n19119), .ZN(
        n19116) );
  INV_X1 U22076 ( .A(n19116), .ZN(n19118) );
  AOI22_X1 U22077 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19125), .B1(
        n19124), .B2(n19456), .ZN(n19117) );
  OAI211_X1 U22078 ( .C1(n19459), .C2(n19130), .A(n19118), .B(n19117), .ZN(
        P2_U3062) );
  INV_X1 U22079 ( .A(n19589), .ZN(n19121) );
  INV_X1 U22080 ( .A(n19587), .ZN(n19120) );
  OAI22_X1 U22081 ( .A1(n19122), .A2(n19121), .B1(n19120), .B2(n19119), .ZN(
        n19123) );
  INV_X1 U22082 ( .A(n19123), .ZN(n19127) );
  AOI22_X1 U22083 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19125), .B1(
        n19124), .B2(n19462), .ZN(n19126) );
  OAI211_X1 U22084 ( .C1(n19467), .C2(n19130), .A(n19127), .B(n19126), .ZN(
        P2_U3063) );
  NOR3_X2 U22085 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19710), .A3(
        n19157), .ZN(n19151) );
  OAI21_X1 U22086 ( .B1(n19133), .B2(n19151), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19129) );
  NOR2_X1 U22087 ( .A1(n19370), .A2(n19157), .ZN(n19131) );
  INV_X1 U22088 ( .A(n19131), .ZN(n19128) );
  NAND2_X1 U22089 ( .A1(n19129), .A2(n19128), .ZN(n19152) );
  AOI22_X1 U22090 ( .A1(n19152), .A2(n19034), .B1(n19539), .B2(n19151), .ZN(
        n19138) );
  NAND2_X1 U22091 ( .A1(n19186), .A2(n19130), .ZN(n19132) );
  AOI21_X1 U22092 ( .B1(n19132), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19131), 
        .ZN(n19135) );
  AOI21_X1 U22093 ( .B1(n19133), .B2(n19732), .A(n19151), .ZN(n19134) );
  INV_X1 U22094 ( .A(n19688), .ZN(n19683) );
  MUX2_X1 U22095 ( .A(n19135), .B(n19134), .S(n19683), .Z(n19136) );
  AOI22_X1 U22096 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19154), .B1(
        n19153), .B2(n19499), .ZN(n19137) );
  OAI211_X1 U22097 ( .C1(n19511), .C2(n19186), .A(n19138), .B(n19137), .ZN(
        P2_U3064) );
  AOI22_X1 U22098 ( .A1(n19152), .A2(n19552), .B1(n19551), .B2(n19151), .ZN(
        n19140) );
  AOI22_X1 U22099 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19154), .B1(
        n19153), .B2(n19438), .ZN(n19139) );
  OAI211_X1 U22100 ( .C1(n19441), .C2(n19186), .A(n19140), .B(n19139), .ZN(
        P2_U3065) );
  AOI22_X1 U22101 ( .A1(n19152), .A2(n19558), .B1(n19557), .B2(n19151), .ZN(
        n19142) );
  AOI22_X1 U22102 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19154), .B1(
        n19153), .B2(n19442), .ZN(n19141) );
  OAI211_X1 U22103 ( .C1(n19445), .C2(n19186), .A(n19142), .B(n19141), .ZN(
        P2_U3066) );
  AOI22_X1 U22104 ( .A1(n19152), .A2(n19564), .B1(n19563), .B2(n19151), .ZN(
        n19144) );
  AOI22_X1 U22105 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19154), .B1(
        n19153), .B2(n19446), .ZN(n19143) );
  OAI211_X1 U22106 ( .C1(n19449), .C2(n19186), .A(n19144), .B(n19143), .ZN(
        P2_U3067) );
  AOI22_X1 U22107 ( .A1(n19152), .A2(n19570), .B1(n19569), .B2(n19151), .ZN(
        n19146) );
  AOI22_X1 U22108 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19154), .B1(
        n19153), .B2(n19450), .ZN(n19145) );
  OAI211_X1 U22109 ( .C1(n19453), .C2(n19186), .A(n19146), .B(n19145), .ZN(
        P2_U3068) );
  AOI22_X1 U22110 ( .A1(n19152), .A2(n19576), .B1(n19575), .B2(n19151), .ZN(
        n19148) );
  AOI22_X1 U22111 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19154), .B1(
        n19153), .B2(n19520), .ZN(n19147) );
  OAI211_X1 U22112 ( .C1(n19524), .C2(n19186), .A(n19148), .B(n19147), .ZN(
        P2_U3069) );
  AOI22_X1 U22113 ( .A1(n19152), .A2(n19582), .B1(n19581), .B2(n19151), .ZN(
        n19150) );
  AOI22_X1 U22114 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19154), .B1(
        n19153), .B2(n19456), .ZN(n19149) );
  OAI211_X1 U22115 ( .C1(n19459), .C2(n19186), .A(n19150), .B(n19149), .ZN(
        P2_U3070) );
  AOI22_X1 U22116 ( .A1(n19152), .A2(n19589), .B1(n19587), .B2(n19151), .ZN(
        n19156) );
  AOI22_X1 U22117 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19154), .B1(
        n19153), .B2(n19462), .ZN(n19155) );
  OAI211_X1 U22118 ( .C1(n19467), .C2(n19186), .A(n19156), .B(n19155), .ZN(
        P2_U3071) );
  INV_X1 U22119 ( .A(n19213), .ZN(n19178) );
  INV_X1 U22120 ( .A(n19186), .ZN(n19175) );
  NOR2_X1 U22121 ( .A1(n19397), .A2(n19157), .ZN(n19181) );
  AOI22_X1 U22122 ( .A1(n19175), .A2(n19499), .B1(n19181), .B2(n19539), .ZN(
        n19166) );
  OAI21_X1 U22123 ( .B1(n19268), .B2(n19403), .A(n19688), .ZN(n19164) );
  NOR2_X1 U22124 ( .A1(n19710), .A2(n19157), .ZN(n19161) );
  INV_X1 U22125 ( .A(n12279), .ZN(n19159) );
  INV_X1 U22126 ( .A(n19181), .ZN(n19158) );
  OAI211_X1 U22127 ( .C1(n19159), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19158), 
        .B(n19683), .ZN(n19160) );
  OAI211_X1 U22128 ( .C1(n19164), .C2(n19161), .A(n19544), .B(n19160), .ZN(
        n19183) );
  INV_X1 U22129 ( .A(n19161), .ZN(n19163) );
  OAI21_X1 U22130 ( .B1(n12279), .B2(n19181), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19162) );
  OAI21_X1 U22131 ( .B1(n19164), .B2(n19163), .A(n19162), .ZN(n19182) );
  AOI22_X1 U22132 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19183), .B1(
        n19034), .B2(n19182), .ZN(n19165) );
  OAI211_X1 U22133 ( .C1(n19511), .C2(n19178), .A(n19166), .B(n19165), .ZN(
        P2_U3072) );
  AOI22_X1 U22134 ( .A1(n19553), .A2(n19213), .B1(n19551), .B2(n19181), .ZN(
        n19168) );
  AOI22_X1 U22135 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19183), .B1(
        n19552), .B2(n19182), .ZN(n19167) );
  OAI211_X1 U22136 ( .C1(n19556), .C2(n19186), .A(n19168), .B(n19167), .ZN(
        P2_U3073) );
  INV_X1 U22137 ( .A(n19445), .ZN(n19559) );
  AOI22_X1 U22138 ( .A1(n19559), .A2(n19213), .B1(n19181), .B2(n19557), .ZN(
        n19170) );
  AOI22_X1 U22139 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19183), .B1(
        n19558), .B2(n19182), .ZN(n19169) );
  OAI211_X1 U22140 ( .C1(n19562), .C2(n19186), .A(n19170), .B(n19169), .ZN(
        P2_U3074) );
  AOI22_X1 U22141 ( .A1(n19175), .A2(n19446), .B1(n19181), .B2(n19563), .ZN(
        n19172) );
  AOI22_X1 U22142 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19183), .B1(
        n19564), .B2(n19182), .ZN(n19171) );
  OAI211_X1 U22143 ( .C1(n19449), .C2(n19178), .A(n19172), .B(n19171), .ZN(
        P2_U3075) );
  AOI22_X1 U22144 ( .A1(n19175), .A2(n19450), .B1(n19181), .B2(n19569), .ZN(
        n19174) );
  AOI22_X1 U22145 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19183), .B1(
        n19570), .B2(n19182), .ZN(n19173) );
  OAI211_X1 U22146 ( .C1(n19453), .C2(n19178), .A(n19174), .B(n19173), .ZN(
        P2_U3076) );
  AOI22_X1 U22147 ( .A1(n19175), .A2(n19520), .B1(n19181), .B2(n19575), .ZN(
        n19177) );
  AOI22_X1 U22148 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19183), .B1(
        n19576), .B2(n19182), .ZN(n19176) );
  OAI211_X1 U22149 ( .C1(n19524), .C2(n19178), .A(n19177), .B(n19176), .ZN(
        P2_U3077) );
  AOI22_X1 U22150 ( .A1(n19583), .A2(n19213), .B1(n19181), .B2(n19581), .ZN(
        n19180) );
  AOI22_X1 U22151 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19183), .B1(
        n19582), .B2(n19182), .ZN(n19179) );
  OAI211_X1 U22152 ( .C1(n19586), .C2(n19186), .A(n19180), .B(n19179), .ZN(
        P2_U3078) );
  INV_X1 U22153 ( .A(n19467), .ZN(n19591) );
  AOI22_X1 U22154 ( .A1(n19591), .A2(n19213), .B1(n19181), .B2(n19587), .ZN(
        n19185) );
  AOI22_X1 U22155 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19183), .B1(
        n19589), .B2(n19182), .ZN(n19184) );
  OAI211_X1 U22156 ( .C1(n19597), .C2(n19186), .A(n19185), .B(n19184), .ZN(
        P2_U3079) );
  INV_X1 U22157 ( .A(n19476), .ZN(n19218) );
  INV_X1 U22158 ( .A(n19188), .ZN(n19190) );
  NOR2_X1 U22159 ( .A1(n19190), .A2(n19189), .ZN(n19434) );
  NAND2_X1 U22160 ( .A1(n19434), .A2(n19693), .ZN(n19195) );
  NOR2_X1 U22161 ( .A1(n19306), .A2(n19217), .ZN(n19211) );
  OAI21_X1 U22162 ( .B1(n19192), .B2(n19211), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19191) );
  OAI21_X1 U22163 ( .B1(n19195), .B2(n19683), .A(n19191), .ZN(n19212) );
  AOI22_X1 U22164 ( .A1(n19212), .A2(n19034), .B1(n19539), .B2(n19211), .ZN(
        n19198) );
  OAI21_X1 U22165 ( .B1(n19213), .B2(n19236), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19194) );
  AOI211_X1 U22166 ( .C1(n19192), .C2(n19732), .A(n19211), .B(n19688), .ZN(
        n19193) );
  AOI211_X1 U22167 ( .C1(n19195), .C2(n19194), .A(n19338), .B(n19193), .ZN(
        n19196) );
  AOI22_X1 U22168 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19214), .B1(
        n19213), .B2(n19499), .ZN(n19197) );
  OAI211_X1 U22169 ( .C1(n19511), .C2(n19246), .A(n19198), .B(n19197), .ZN(
        P2_U3080) );
  AOI22_X1 U22170 ( .A1(n19212), .A2(n19552), .B1(n19551), .B2(n19211), .ZN(
        n19200) );
  AOI22_X1 U22171 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19214), .B1(
        n19213), .B2(n19438), .ZN(n19199) );
  OAI211_X1 U22172 ( .C1(n19441), .C2(n19246), .A(n19200), .B(n19199), .ZN(
        P2_U3081) );
  AOI22_X1 U22173 ( .A1(n19212), .A2(n19558), .B1(n19557), .B2(n19211), .ZN(
        n19202) );
  AOI22_X1 U22174 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19214), .B1(
        n19213), .B2(n19442), .ZN(n19201) );
  OAI211_X1 U22175 ( .C1(n19445), .C2(n19246), .A(n19202), .B(n19201), .ZN(
        P2_U3082) );
  AOI22_X1 U22176 ( .A1(n19212), .A2(n19564), .B1(n19563), .B2(n19211), .ZN(
        n19204) );
  AOI22_X1 U22177 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19214), .B1(
        n19213), .B2(n19446), .ZN(n19203) );
  OAI211_X1 U22178 ( .C1(n19449), .C2(n19246), .A(n19204), .B(n19203), .ZN(
        P2_U3083) );
  AOI22_X1 U22179 ( .A1(n19212), .A2(n19570), .B1(n19569), .B2(n19211), .ZN(
        n19206) );
  AOI22_X1 U22180 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19214), .B1(
        n19213), .B2(n19450), .ZN(n19205) );
  OAI211_X1 U22181 ( .C1(n19453), .C2(n19246), .A(n19206), .B(n19205), .ZN(
        P2_U3084) );
  AOI22_X1 U22182 ( .A1(n19212), .A2(n19576), .B1(n19575), .B2(n19211), .ZN(
        n19208) );
  AOI22_X1 U22183 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19214), .B1(
        n19213), .B2(n19520), .ZN(n19207) );
  OAI211_X1 U22184 ( .C1(n19524), .C2(n19246), .A(n19208), .B(n19207), .ZN(
        P2_U3085) );
  AOI22_X1 U22185 ( .A1(n19212), .A2(n19582), .B1(n19581), .B2(n19211), .ZN(
        n19210) );
  AOI22_X1 U22186 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19214), .B1(
        n19213), .B2(n19456), .ZN(n19209) );
  OAI211_X1 U22187 ( .C1(n19459), .C2(n19246), .A(n19210), .B(n19209), .ZN(
        P2_U3086) );
  AOI22_X1 U22188 ( .A1(n19212), .A2(n19589), .B1(n19587), .B2(n19211), .ZN(
        n19216) );
  AOI22_X1 U22189 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19214), .B1(
        n19213), .B2(n19462), .ZN(n19215) );
  OAI211_X1 U22190 ( .C1(n19467), .C2(n19246), .A(n19216), .B(n19215), .ZN(
        P2_U3087) );
  NOR2_X1 U22191 ( .A1(n19217), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19222) );
  INV_X1 U22192 ( .A(n19222), .ZN(n19224) );
  NOR2_X1 U22193 ( .A1(n19720), .A2(n19224), .ZN(n19241) );
  AOI22_X1 U22194 ( .A1(n19547), .A2(n19247), .B1(n19539), .B2(n19241), .ZN(
        n19227) );
  OAI21_X1 U22195 ( .B1(n19268), .B2(n19218), .A(n19688), .ZN(n19225) );
  INV_X1 U22196 ( .A(n12291), .ZN(n19220) );
  INV_X1 U22197 ( .A(n19241), .ZN(n19219) );
  OAI211_X1 U22198 ( .C1(n19220), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19219), 
        .B(n19683), .ZN(n19221) );
  OAI211_X1 U22199 ( .C1(n19225), .C2(n19222), .A(n19544), .B(n19221), .ZN(
        n19243) );
  OAI21_X1 U22200 ( .B1(n12291), .B2(n19241), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19223) );
  OAI21_X1 U22201 ( .B1(n19225), .B2(n19224), .A(n19223), .ZN(n19242) );
  AOI22_X1 U22202 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19243), .B1(
        n19034), .B2(n19242), .ZN(n19226) );
  OAI211_X1 U22203 ( .C1(n19550), .C2(n19246), .A(n19227), .B(n19226), .ZN(
        P2_U3088) );
  AOI22_X1 U22204 ( .A1(n19553), .A2(n19247), .B1(n19551), .B2(n19241), .ZN(
        n19229) );
  AOI22_X1 U22205 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19243), .B1(
        n19552), .B2(n19242), .ZN(n19228) );
  OAI211_X1 U22206 ( .C1(n19556), .C2(n19246), .A(n19229), .B(n19228), .ZN(
        P2_U3089) );
  AOI22_X1 U22207 ( .A1(n19236), .A2(n19442), .B1(n19557), .B2(n19241), .ZN(
        n19231) );
  AOI22_X1 U22208 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19243), .B1(
        n19558), .B2(n19242), .ZN(n19230) );
  OAI211_X1 U22209 ( .C1(n19445), .C2(n19267), .A(n19231), .B(n19230), .ZN(
        P2_U3090) );
  AOI22_X1 U22210 ( .A1(n19236), .A2(n19446), .B1(n19563), .B2(n19241), .ZN(
        n19233) );
  AOI22_X1 U22211 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19243), .B1(
        n19564), .B2(n19242), .ZN(n19232) );
  OAI211_X1 U22212 ( .C1(n19449), .C2(n19267), .A(n19233), .B(n19232), .ZN(
        P2_U3091) );
  AOI22_X1 U22213 ( .A1(n19236), .A2(n19450), .B1(n19569), .B2(n19241), .ZN(
        n19235) );
  AOI22_X1 U22214 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19243), .B1(
        n19570), .B2(n19242), .ZN(n19234) );
  OAI211_X1 U22215 ( .C1(n19453), .C2(n19267), .A(n19235), .B(n19234), .ZN(
        P2_U3092) );
  AOI22_X1 U22216 ( .A1(n19236), .A2(n19520), .B1(n19575), .B2(n19241), .ZN(
        n19238) );
  AOI22_X1 U22217 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19243), .B1(
        n19576), .B2(n19242), .ZN(n19237) );
  OAI211_X1 U22218 ( .C1(n19524), .C2(n19267), .A(n19238), .B(n19237), .ZN(
        P2_U3093) );
  AOI22_X1 U22219 ( .A1(n19583), .A2(n19247), .B1(n19581), .B2(n19241), .ZN(
        n19240) );
  AOI22_X1 U22220 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19243), .B1(
        n19582), .B2(n19242), .ZN(n19239) );
  OAI211_X1 U22221 ( .C1(n19586), .C2(n19246), .A(n19240), .B(n19239), .ZN(
        P2_U3094) );
  AOI22_X1 U22222 ( .A1(n19591), .A2(n19247), .B1(n19587), .B2(n19241), .ZN(
        n19245) );
  AOI22_X1 U22223 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19243), .B1(
        n19589), .B2(n19242), .ZN(n19244) );
  OAI211_X1 U22224 ( .C1(n19597), .C2(n19246), .A(n19245), .B(n19244), .ZN(
        P2_U3095) );
  AOI22_X1 U22225 ( .A1(n19263), .A2(n19034), .B1(n19262), .B2(n19539), .ZN(
        n19249) );
  AOI22_X1 U22226 ( .A1(n19247), .A2(n19499), .B1(n19299), .B2(n19547), .ZN(
        n19248) );
  OAI211_X1 U22227 ( .C1(n19251), .C2(n19250), .A(n19249), .B(n19248), .ZN(
        P2_U3096) );
  AOI22_X1 U22228 ( .A1(n19263), .A2(n19558), .B1(n19262), .B2(n19557), .ZN(
        n19253) );
  AOI22_X1 U22229 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19264), .B1(
        n19299), .B2(n19559), .ZN(n19252) );
  OAI211_X1 U22230 ( .C1(n19562), .C2(n19267), .A(n19253), .B(n19252), .ZN(
        P2_U3098) );
  AOI22_X1 U22231 ( .A1(n19263), .A2(n19564), .B1(n19262), .B2(n19563), .ZN(
        n19255) );
  AOI22_X1 U22232 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19264), .B1(
        n19299), .B2(n19565), .ZN(n19254) );
  OAI211_X1 U22233 ( .C1(n19568), .C2(n19267), .A(n19255), .B(n19254), .ZN(
        P2_U3099) );
  AOI22_X1 U22234 ( .A1(n19263), .A2(n19570), .B1(n19262), .B2(n19569), .ZN(
        n19257) );
  INV_X1 U22235 ( .A(n19453), .ZN(n19571) );
  AOI22_X1 U22236 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19264), .B1(
        n19299), .B2(n19571), .ZN(n19256) );
  OAI211_X1 U22237 ( .C1(n19574), .C2(n19267), .A(n19257), .B(n19256), .ZN(
        P2_U3100) );
  AOI22_X1 U22238 ( .A1(n19263), .A2(n19576), .B1(n19262), .B2(n19575), .ZN(
        n19259) );
  INV_X1 U22239 ( .A(n19524), .ZN(n19577) );
  AOI22_X1 U22240 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19264), .B1(
        n19299), .B2(n19577), .ZN(n19258) );
  OAI211_X1 U22241 ( .C1(n19580), .C2(n19267), .A(n19259), .B(n19258), .ZN(
        P2_U3101) );
  AOI22_X1 U22242 ( .A1(n19263), .A2(n19582), .B1(n19262), .B2(n19581), .ZN(
        n19261) );
  AOI22_X1 U22243 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19264), .B1(
        n19299), .B2(n19583), .ZN(n19260) );
  OAI211_X1 U22244 ( .C1(n19586), .C2(n19267), .A(n19261), .B(n19260), .ZN(
        P2_U3102) );
  AOI22_X1 U22245 ( .A1(n19263), .A2(n19589), .B1(n19262), .B2(n19587), .ZN(
        n19266) );
  AOI22_X1 U22246 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19264), .B1(
        n19299), .B2(n19591), .ZN(n19265) );
  OAI211_X1 U22247 ( .C1(n19597), .C2(n19267), .A(n19266), .B(n19265), .ZN(
        P2_U3103) );
  NAND2_X1 U22248 ( .A1(n19693), .A2(n19536), .ZN(n19275) );
  INV_X1 U22249 ( .A(n19275), .ZN(n19269) );
  NOR2_X1 U22250 ( .A1(n19268), .A2(n19540), .ZN(n19687) );
  OAI21_X1 U22251 ( .B1(n19269), .B2(n19687), .A(n19544), .ZN(n19274) );
  INV_X1 U22252 ( .A(n19397), .ZN(n19271) );
  NAND2_X1 U22253 ( .A1(n19271), .A2(n19270), .ZN(n19309) );
  INV_X1 U22254 ( .A(n19309), .ZN(n19312) );
  NAND2_X1 U22255 ( .A1(n19309), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19272) );
  OR2_X1 U22256 ( .A1(n12278), .A2(n19272), .ZN(n19277) );
  OAI21_X1 U22257 ( .B1(n19312), .B2(n19732), .A(n19277), .ZN(n19273) );
  INV_X1 U22258 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n19281) );
  OAI21_X1 U22259 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19275), .A(n19733), 
        .ZN(n19276) );
  AND2_X1 U22260 ( .A1(n19277), .A2(n19276), .ZN(n19298) );
  AOI22_X1 U22261 ( .A1(n19298), .A2(n19034), .B1(n19312), .B2(n19539), .ZN(
        n19280) );
  AOI22_X1 U22262 ( .A1(n19328), .A2(n19547), .B1(n19299), .B2(n19499), .ZN(
        n19279) );
  OAI211_X1 U22263 ( .C1(n19293), .C2(n19281), .A(n19280), .B(n19279), .ZN(
        P2_U3104) );
  INV_X1 U22264 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n19284) );
  AOI22_X1 U22265 ( .A1(n19298), .A2(n19552), .B1(n19551), .B2(n19312), .ZN(
        n19283) );
  AOI22_X1 U22266 ( .A1(n19328), .A2(n19553), .B1(n19299), .B2(n19438), .ZN(
        n19282) );
  OAI211_X1 U22267 ( .C1(n19293), .C2(n19284), .A(n19283), .B(n19282), .ZN(
        P2_U3105) );
  INV_X1 U22268 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n19287) );
  AOI22_X1 U22269 ( .A1(n19298), .A2(n19558), .B1(n19312), .B2(n19557), .ZN(
        n19286) );
  AOI22_X1 U22270 ( .A1(n19328), .A2(n19559), .B1(n19299), .B2(n19442), .ZN(
        n19285) );
  OAI211_X1 U22271 ( .C1(n19293), .C2(n19287), .A(n19286), .B(n19285), .ZN(
        P2_U3106) );
  AOI22_X1 U22272 ( .A1(n19298), .A2(n19564), .B1(n19312), .B2(n19563), .ZN(
        n19289) );
  AOI22_X1 U22273 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19300), .B1(
        n19299), .B2(n19446), .ZN(n19288) );
  OAI211_X1 U22274 ( .C1(n19449), .C2(n19336), .A(n19289), .B(n19288), .ZN(
        P2_U3107) );
  INV_X1 U22275 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n19292) );
  AOI22_X1 U22276 ( .A1(n19298), .A2(n19570), .B1(n19312), .B2(n19569), .ZN(
        n19291) );
  AOI22_X1 U22277 ( .A1(n19328), .A2(n19571), .B1(n19299), .B2(n19450), .ZN(
        n19290) );
  OAI211_X1 U22278 ( .C1(n19293), .C2(n19292), .A(n19291), .B(n19290), .ZN(
        P2_U3108) );
  AOI22_X1 U22279 ( .A1(n19298), .A2(n19576), .B1(n19312), .B2(n19575), .ZN(
        n19295) );
  AOI22_X1 U22280 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19300), .B1(
        n19299), .B2(n19520), .ZN(n19294) );
  OAI211_X1 U22281 ( .C1(n19524), .C2(n19336), .A(n19295), .B(n19294), .ZN(
        P2_U3109) );
  AOI22_X1 U22282 ( .A1(n19298), .A2(n19582), .B1(n19312), .B2(n19581), .ZN(
        n19297) );
  AOI22_X1 U22283 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19300), .B1(
        n19299), .B2(n19456), .ZN(n19296) );
  OAI211_X1 U22284 ( .C1(n19459), .C2(n19336), .A(n19297), .B(n19296), .ZN(
        P2_U3110) );
  AOI22_X1 U22285 ( .A1(n19298), .A2(n19589), .B1(n19312), .B2(n19587), .ZN(
        n19302) );
  AOI22_X1 U22286 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19300), .B1(
        n19299), .B2(n19462), .ZN(n19301) );
  OAI211_X1 U22287 ( .C1(n19467), .C2(n19336), .A(n19302), .B(n19301), .ZN(
        P2_U3111) );
  NAND2_X1 U22288 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19700), .ZN(
        n19396) );
  NOR2_X1 U22289 ( .A1(n19306), .A2(n19396), .ZN(n19331) );
  AOI22_X1 U22290 ( .A1(n19328), .A2(n19499), .B1(n19331), .B2(n19539), .ZN(
        n19317) );
  NAND2_X1 U22291 ( .A1(n19361), .A2(n19336), .ZN(n19307) );
  AOI21_X1 U22292 ( .B1(n19307), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19683), 
        .ZN(n19311) );
  AOI21_X1 U22293 ( .B1(n19313), .B2(n19732), .A(n19688), .ZN(n19308) );
  AOI21_X1 U22294 ( .B1(n19311), .B2(n19309), .A(n19308), .ZN(n19310) );
  OAI21_X1 U22295 ( .B1(n19331), .B2(n19310), .A(n19544), .ZN(n19333) );
  OAI21_X1 U22296 ( .B1(n19312), .B2(n19331), .A(n19311), .ZN(n19315) );
  OAI21_X1 U22297 ( .B1(n19313), .B2(n19331), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19314) );
  NAND2_X1 U22298 ( .A1(n19315), .A2(n19314), .ZN(n19332) );
  AOI22_X1 U22299 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19333), .B1(
        n19034), .B2(n19332), .ZN(n19316) );
  OAI211_X1 U22300 ( .C1(n19511), .C2(n19361), .A(n19317), .B(n19316), .ZN(
        P2_U3112) );
  AOI22_X1 U22301 ( .A1(n19328), .A2(n19438), .B1(n19551), .B2(n19331), .ZN(
        n19319) );
  AOI22_X1 U22302 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19333), .B1(
        n19332), .B2(n19552), .ZN(n19318) );
  OAI211_X1 U22303 ( .C1(n19441), .C2(n19361), .A(n19319), .B(n19318), .ZN(
        P2_U3113) );
  AOI22_X1 U22304 ( .A1(n19362), .A2(n19559), .B1(n19557), .B2(n19331), .ZN(
        n19321) );
  AOI22_X1 U22305 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19333), .B1(
        n19332), .B2(n19558), .ZN(n19320) );
  OAI211_X1 U22306 ( .C1(n19562), .C2(n19336), .A(n19321), .B(n19320), .ZN(
        P2_U3114) );
  AOI22_X1 U22307 ( .A1(n19362), .A2(n19565), .B1(n19331), .B2(n19563), .ZN(
        n19323) );
  AOI22_X1 U22308 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19333), .B1(
        n19332), .B2(n19564), .ZN(n19322) );
  OAI211_X1 U22309 ( .C1(n19568), .C2(n19336), .A(n19323), .B(n19322), .ZN(
        P2_U3115) );
  AOI22_X1 U22310 ( .A1(n19362), .A2(n19571), .B1(n19331), .B2(n19569), .ZN(
        n19325) );
  AOI22_X1 U22311 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19333), .B1(
        n19332), .B2(n19570), .ZN(n19324) );
  OAI211_X1 U22312 ( .C1(n19574), .C2(n19336), .A(n19325), .B(n19324), .ZN(
        P2_U3116) );
  AOI22_X1 U22313 ( .A1(n19362), .A2(n19577), .B1(n19331), .B2(n19575), .ZN(
        n19327) );
  AOI22_X1 U22314 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19333), .B1(
        n19332), .B2(n19576), .ZN(n19326) );
  OAI211_X1 U22315 ( .C1(n19580), .C2(n19336), .A(n19327), .B(n19326), .ZN(
        P2_U3117) );
  AOI22_X1 U22316 ( .A1(n19328), .A2(n19456), .B1(n19331), .B2(n19581), .ZN(
        n19330) );
  AOI22_X1 U22317 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19333), .B1(
        n19332), .B2(n19582), .ZN(n19329) );
  OAI211_X1 U22318 ( .C1(n19459), .C2(n19361), .A(n19330), .B(n19329), .ZN(
        P2_U3118) );
  AOI22_X1 U22319 ( .A1(n19362), .A2(n19591), .B1(n19331), .B2(n19587), .ZN(
        n19335) );
  AOI22_X1 U22320 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19333), .B1(
        n19332), .B2(n19589), .ZN(n19334) );
  OAI211_X1 U22321 ( .C1(n19597), .C2(n19336), .A(n19335), .B(n19334), .ZN(
        P2_U3119) );
  NOR3_X2 U22322 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19720), .A3(
        n19396), .ZN(n19371) );
  AOI22_X1 U22323 ( .A1(n19392), .A2(n19547), .B1(n19371), .B2(n19539), .ZN(
        n19348) );
  NAND2_X1 U22324 ( .A1(n19690), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19541) );
  OAI21_X1 U22325 ( .B1(n19541), .B2(n19337), .A(n19688), .ZN(n19346) );
  NOR2_X1 U22326 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19396), .ZN(
        n19342) );
  OAI21_X1 U22327 ( .B1(n19343), .B2(n19733), .A(n19732), .ZN(n19340) );
  INV_X1 U22328 ( .A(n19371), .ZN(n19339) );
  AOI21_X1 U22329 ( .B1(n19340), .B2(n19339), .A(n19338), .ZN(n19341) );
  OAI21_X1 U22330 ( .B1(n19346), .B2(n19342), .A(n19341), .ZN(n19364) );
  INV_X1 U22331 ( .A(n19342), .ZN(n19345) );
  OAI21_X1 U22332 ( .B1(n19343), .B2(n19371), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19344) );
  OAI21_X1 U22333 ( .B1(n19346), .B2(n19345), .A(n19344), .ZN(n19363) );
  AOI22_X1 U22334 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19364), .B1(
        n19034), .B2(n19363), .ZN(n19347) );
  OAI211_X1 U22335 ( .C1(n19550), .C2(n19361), .A(n19348), .B(n19347), .ZN(
        P2_U3120) );
  AOI22_X1 U22336 ( .A1(n19392), .A2(n19553), .B1(n19551), .B2(n19371), .ZN(
        n19350) );
  AOI22_X1 U22337 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19364), .B1(
        n19552), .B2(n19363), .ZN(n19349) );
  OAI211_X1 U22338 ( .C1(n19556), .C2(n19361), .A(n19350), .B(n19349), .ZN(
        P2_U3121) );
  INV_X1 U22339 ( .A(n19392), .ZN(n19367) );
  AOI22_X1 U22340 ( .A1(n19362), .A2(n19442), .B1(n19557), .B2(n19371), .ZN(
        n19352) );
  AOI22_X1 U22341 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19364), .B1(
        n19558), .B2(n19363), .ZN(n19351) );
  OAI211_X1 U22342 ( .C1(n19445), .C2(n19367), .A(n19352), .B(n19351), .ZN(
        P2_U3122) );
  AOI22_X1 U22343 ( .A1(n19565), .A2(n19392), .B1(n19563), .B2(n19371), .ZN(
        n19354) );
  AOI22_X1 U22344 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19364), .B1(
        n19564), .B2(n19363), .ZN(n19353) );
  OAI211_X1 U22345 ( .C1(n19568), .C2(n19361), .A(n19354), .B(n19353), .ZN(
        P2_U3123) );
  AOI22_X1 U22346 ( .A1(n19362), .A2(n19450), .B1(n19569), .B2(n19371), .ZN(
        n19356) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19364), .B1(
        n19570), .B2(n19363), .ZN(n19355) );
  OAI211_X1 U22348 ( .C1(n19453), .C2(n19367), .A(n19356), .B(n19355), .ZN(
        P2_U3124) );
  AOI22_X1 U22349 ( .A1(n19577), .A2(n19392), .B1(n19575), .B2(n19371), .ZN(
        n19358) );
  AOI22_X1 U22350 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19364), .B1(
        n19576), .B2(n19363), .ZN(n19357) );
  OAI211_X1 U22351 ( .C1(n19580), .C2(n19361), .A(n19358), .B(n19357), .ZN(
        P2_U3125) );
  AOI22_X1 U22352 ( .A1(n19583), .A2(n19392), .B1(n19371), .B2(n19581), .ZN(
        n19360) );
  AOI22_X1 U22353 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19364), .B1(
        n19582), .B2(n19363), .ZN(n19359) );
  OAI211_X1 U22354 ( .C1(n19586), .C2(n19361), .A(n19360), .B(n19359), .ZN(
        P2_U3126) );
  AOI22_X1 U22355 ( .A1(n19362), .A2(n19462), .B1(n19587), .B2(n19371), .ZN(
        n19366) );
  AOI22_X1 U22356 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19364), .B1(
        n19589), .B2(n19363), .ZN(n19365) );
  OAI211_X1 U22357 ( .C1(n19467), .C2(n19367), .A(n19366), .B(n19365), .ZN(
        P2_U3127) );
  NOR3_X2 U22358 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19710), .A3(
        n19396), .ZN(n19390) );
  OAI21_X1 U22359 ( .B1(n19368), .B2(n19390), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19369) );
  OAI21_X1 U22360 ( .B1(n19396), .B2(n19370), .A(n19369), .ZN(n19391) );
  AOI22_X1 U22361 ( .A1(n19391), .A2(n19034), .B1(n19539), .B2(n19390), .ZN(
        n19377) );
  AOI221_X1 U22362 ( .B1(n19416), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19392), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19371), .ZN(n19373) );
  MUX2_X1 U22363 ( .A(n19373), .B(n19372), .S(P2_STATE2_REG_2__SCAN_IN), .Z(
        n19374) );
  NOR2_X1 U22364 ( .A1(n19374), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19375) );
  AOI22_X1 U22365 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19393), .B1(
        n19392), .B2(n19499), .ZN(n19376) );
  OAI211_X1 U22366 ( .C1(n19511), .C2(n19424), .A(n19377), .B(n19376), .ZN(
        P2_U3128) );
  AOI22_X1 U22367 ( .A1(n19391), .A2(n19552), .B1(n19551), .B2(n19390), .ZN(
        n19379) );
  AOI22_X1 U22368 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19393), .B1(
        n19392), .B2(n19438), .ZN(n19378) );
  OAI211_X1 U22369 ( .C1(n19441), .C2(n19424), .A(n19379), .B(n19378), .ZN(
        P2_U3129) );
  AOI22_X1 U22370 ( .A1(n19391), .A2(n19558), .B1(n19557), .B2(n19390), .ZN(
        n19381) );
  AOI22_X1 U22371 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19393), .B1(
        n19392), .B2(n19442), .ZN(n19380) );
  OAI211_X1 U22372 ( .C1(n19445), .C2(n19424), .A(n19381), .B(n19380), .ZN(
        P2_U3130) );
  AOI22_X1 U22373 ( .A1(n19391), .A2(n19564), .B1(n19563), .B2(n19390), .ZN(
        n19383) );
  AOI22_X1 U22374 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19393), .B1(
        n19392), .B2(n19446), .ZN(n19382) );
  OAI211_X1 U22375 ( .C1(n19449), .C2(n19424), .A(n19383), .B(n19382), .ZN(
        P2_U3131) );
  AOI22_X1 U22376 ( .A1(n19391), .A2(n19570), .B1(n19569), .B2(n19390), .ZN(
        n19385) );
  AOI22_X1 U22377 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19393), .B1(
        n19392), .B2(n19450), .ZN(n19384) );
  OAI211_X1 U22378 ( .C1(n19453), .C2(n19424), .A(n19385), .B(n19384), .ZN(
        P2_U3132) );
  AOI22_X1 U22379 ( .A1(n19391), .A2(n19576), .B1(n19575), .B2(n19390), .ZN(
        n19387) );
  AOI22_X1 U22380 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19393), .B1(
        n19392), .B2(n19520), .ZN(n19386) );
  OAI211_X1 U22381 ( .C1(n19524), .C2(n19424), .A(n19387), .B(n19386), .ZN(
        P2_U3133) );
  AOI22_X1 U22382 ( .A1(n19391), .A2(n19582), .B1(n19581), .B2(n19390), .ZN(
        n19389) );
  AOI22_X1 U22383 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19393), .B1(
        n19392), .B2(n19456), .ZN(n19388) );
  OAI211_X1 U22384 ( .C1(n19459), .C2(n19424), .A(n19389), .B(n19388), .ZN(
        P2_U3134) );
  AOI22_X1 U22385 ( .A1(n19391), .A2(n19589), .B1(n19587), .B2(n19390), .ZN(
        n19395) );
  AOI22_X1 U22386 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19393), .B1(
        n19392), .B2(n19462), .ZN(n19394) );
  OAI211_X1 U22387 ( .C1(n19467), .C2(n19424), .A(n19395), .B(n19394), .ZN(
        P2_U3135) );
  OR2_X1 U22388 ( .A1(n19710), .A2(n19396), .ZN(n19400) );
  OR2_X1 U22389 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19400), .ZN(n19398) );
  NOR2_X1 U22390 ( .A1(n19397), .A2(n19396), .ZN(n19419) );
  NOR3_X1 U22391 ( .A1(n12245), .A2(n19419), .A3(n19733), .ZN(n19399) );
  AOI21_X1 U22392 ( .B1(n19733), .B2(n19398), .A(n19399), .ZN(n19420) );
  AOI22_X1 U22393 ( .A1(n19420), .A2(n19034), .B1(n19539), .B2(n19419), .ZN(
        n19405) );
  INV_X1 U22394 ( .A(n19541), .ZN(n19470) );
  NAND2_X1 U22395 ( .A1(n19470), .A2(n19684), .ZN(n19401) );
  AOI21_X1 U22396 ( .B1(n19401), .B2(n19400), .A(n19399), .ZN(n19402) );
  OAI211_X1 U22397 ( .C1(n19419), .C2(n19732), .A(n19402), .B(n19544), .ZN(
        n19421) );
  NOR2_X2 U22398 ( .A1(n19475), .A2(n19403), .ZN(n19463) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19421), .B1(
        n19463), .B2(n19547), .ZN(n19404) );
  OAI211_X1 U22400 ( .C1(n19550), .C2(n19424), .A(n19405), .B(n19404), .ZN(
        P2_U3136) );
  AOI22_X1 U22401 ( .A1(n19420), .A2(n19552), .B1(n19551), .B2(n19419), .ZN(
        n19407) );
  AOI22_X1 U22402 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19421), .B1(
        n19416), .B2(n19438), .ZN(n19406) );
  OAI211_X1 U22403 ( .C1(n19441), .C2(n19429), .A(n19407), .B(n19406), .ZN(
        P2_U3137) );
  AOI22_X1 U22404 ( .A1(n19420), .A2(n19558), .B1(n19557), .B2(n19419), .ZN(
        n19409) );
  AOI22_X1 U22405 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19421), .B1(
        n19463), .B2(n19559), .ZN(n19408) );
  OAI211_X1 U22406 ( .C1(n19562), .C2(n19424), .A(n19409), .B(n19408), .ZN(
        P2_U3138) );
  AOI22_X1 U22407 ( .A1(n19420), .A2(n19564), .B1(n19563), .B2(n19419), .ZN(
        n19411) );
  AOI22_X1 U22408 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19421), .B1(
        n19416), .B2(n19446), .ZN(n19410) );
  OAI211_X1 U22409 ( .C1(n19449), .C2(n19429), .A(n19411), .B(n19410), .ZN(
        P2_U3139) );
  AOI22_X1 U22410 ( .A1(n19420), .A2(n19570), .B1(n19569), .B2(n19419), .ZN(
        n19413) );
  AOI22_X1 U22411 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19421), .B1(
        n19416), .B2(n19450), .ZN(n19412) );
  OAI211_X1 U22412 ( .C1(n19453), .C2(n19429), .A(n19413), .B(n19412), .ZN(
        P2_U3140) );
  AOI22_X1 U22413 ( .A1(n19420), .A2(n19576), .B1(n19575), .B2(n19419), .ZN(
        n19415) );
  AOI22_X1 U22414 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19421), .B1(
        n19463), .B2(n19577), .ZN(n19414) );
  OAI211_X1 U22415 ( .C1(n19580), .C2(n19424), .A(n19415), .B(n19414), .ZN(
        P2_U3141) );
  AOI22_X1 U22416 ( .A1(n19420), .A2(n19582), .B1(n19581), .B2(n19419), .ZN(
        n19418) );
  AOI22_X1 U22417 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19421), .B1(
        n19416), .B2(n19456), .ZN(n19417) );
  OAI211_X1 U22418 ( .C1(n19459), .C2(n19429), .A(n19418), .B(n19417), .ZN(
        P2_U3142) );
  AOI22_X1 U22419 ( .A1(n19420), .A2(n19589), .B1(n19587), .B2(n19419), .ZN(
        n19423) );
  AOI22_X1 U22420 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19421), .B1(
        n19463), .B2(n19591), .ZN(n19422) );
  OAI211_X1 U22421 ( .C1(n19597), .C2(n19424), .A(n19423), .B(n19422), .ZN(
        P2_U3143) );
  INV_X1 U22422 ( .A(n19425), .ZN(n19428) );
  INV_X1 U22423 ( .A(n19434), .ZN(n19427) );
  NAND3_X1 U22424 ( .A1(n19710), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19472) );
  NOR2_X1 U22425 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19472), .ZN(
        n19460) );
  OAI21_X1 U22426 ( .B1(n12305), .B2(n19460), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19426) );
  OAI21_X1 U22427 ( .B1(n19428), .B2(n19427), .A(n19426), .ZN(n19461) );
  AOI22_X1 U22428 ( .A1(n19461), .A2(n19034), .B1(n19539), .B2(n19460), .ZN(
        n19437) );
  AOI21_X1 U22429 ( .B1(n19429), .B2(n19496), .A(n19682), .ZN(n19435) );
  INV_X1 U22430 ( .A(n12305), .ZN(n19431) );
  INV_X1 U22431 ( .A(n19460), .ZN(n19430) );
  OAI211_X1 U22432 ( .C1(n19431), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19430), 
        .B(n19683), .ZN(n19432) );
  AND2_X1 U22433 ( .A1(n19432), .A2(n19544), .ZN(n19433) );
  OAI211_X1 U22434 ( .C1(n19435), .C2(n19434), .A(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n19433), .ZN(n19464) );
  AOI22_X1 U22435 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19464), .B1(
        n19463), .B2(n19499), .ZN(n19436) );
  OAI211_X1 U22436 ( .C1(n19511), .C2(n19496), .A(n19437), .B(n19436), .ZN(
        P2_U3144) );
  AOI22_X1 U22437 ( .A1(n19461), .A2(n19552), .B1(n19551), .B2(n19460), .ZN(
        n19440) );
  AOI22_X1 U22438 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19464), .B1(
        n19463), .B2(n19438), .ZN(n19439) );
  OAI211_X1 U22439 ( .C1(n19441), .C2(n19496), .A(n19440), .B(n19439), .ZN(
        P2_U3145) );
  AOI22_X1 U22440 ( .A1(n19461), .A2(n19558), .B1(n19557), .B2(n19460), .ZN(
        n19444) );
  AOI22_X1 U22441 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19464), .B1(
        n19463), .B2(n19442), .ZN(n19443) );
  OAI211_X1 U22442 ( .C1(n19445), .C2(n19496), .A(n19444), .B(n19443), .ZN(
        P2_U3146) );
  AOI22_X1 U22443 ( .A1(n19461), .A2(n19564), .B1(n19563), .B2(n19460), .ZN(
        n19448) );
  AOI22_X1 U22444 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19464), .B1(
        n19463), .B2(n19446), .ZN(n19447) );
  OAI211_X1 U22445 ( .C1(n19449), .C2(n19496), .A(n19448), .B(n19447), .ZN(
        P2_U3147) );
  AOI22_X1 U22446 ( .A1(n19461), .A2(n19570), .B1(n19569), .B2(n19460), .ZN(
        n19452) );
  AOI22_X1 U22447 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19464), .B1(
        n19463), .B2(n19450), .ZN(n19451) );
  OAI211_X1 U22448 ( .C1(n19453), .C2(n19496), .A(n19452), .B(n19451), .ZN(
        P2_U3148) );
  AOI22_X1 U22449 ( .A1(n19461), .A2(n19576), .B1(n19575), .B2(n19460), .ZN(
        n19455) );
  AOI22_X1 U22450 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19464), .B1(
        n19463), .B2(n19520), .ZN(n19454) );
  OAI211_X1 U22451 ( .C1(n19524), .C2(n19496), .A(n19455), .B(n19454), .ZN(
        P2_U3149) );
  AOI22_X1 U22452 ( .A1(n19461), .A2(n19582), .B1(n19581), .B2(n19460), .ZN(
        n19458) );
  AOI22_X1 U22453 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19464), .B1(
        n19463), .B2(n19456), .ZN(n19457) );
  OAI211_X1 U22454 ( .C1(n19459), .C2(n19496), .A(n19458), .B(n19457), .ZN(
        P2_U3150) );
  AOI22_X1 U22455 ( .A1(n19461), .A2(n19589), .B1(n19587), .B2(n19460), .ZN(
        n19466) );
  AOI22_X1 U22456 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19464), .B1(
        n19463), .B2(n19462), .ZN(n19465) );
  OAI211_X1 U22457 ( .C1(n19467), .C2(n19496), .A(n19466), .B(n19465), .ZN(
        P2_U3151) );
  NOR2_X1 U22458 ( .A1(n19720), .A2(n19472), .ZN(n19502) );
  NOR3_X1 U22459 ( .A1(n12288), .A2(n19502), .A3(n19733), .ZN(n19471) );
  INV_X1 U22460 ( .A(n19472), .ZN(n19468) );
  AOI21_X1 U22461 ( .B1(n19732), .B2(n19468), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19469) );
  NOR2_X1 U22462 ( .A1(n19471), .A2(n19469), .ZN(n19492) );
  AOI22_X1 U22463 ( .A1(n19492), .A2(n19034), .B1(n19539), .B2(n19502), .ZN(
        n19479) );
  NAND2_X1 U22464 ( .A1(n19470), .A2(n19476), .ZN(n19473) );
  AOI21_X1 U22465 ( .B1(n19473), .B2(n19472), .A(n19471), .ZN(n19474) );
  OAI211_X1 U22466 ( .C1(n19502), .C2(n19732), .A(n19474), .B(n19544), .ZN(
        n19493) );
  INV_X1 U22467 ( .A(n19475), .ZN(n19477) );
  AOI22_X1 U22468 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19493), .B1(
        n19521), .B2(n19547), .ZN(n19478) );
  OAI211_X1 U22469 ( .C1(n19550), .C2(n19496), .A(n19479), .B(n19478), .ZN(
        P2_U3152) );
  AOI22_X1 U22470 ( .A1(n19492), .A2(n19552), .B1(n19551), .B2(n19502), .ZN(
        n19481) );
  AOI22_X1 U22471 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19493), .B1(
        n19521), .B2(n19553), .ZN(n19480) );
  OAI211_X1 U22472 ( .C1(n19556), .C2(n19496), .A(n19481), .B(n19480), .ZN(
        P2_U3153) );
  AOI22_X1 U22473 ( .A1(n19492), .A2(n19558), .B1(n19557), .B2(n19502), .ZN(
        n19483) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19493), .B1(
        n19521), .B2(n19559), .ZN(n19482) );
  OAI211_X1 U22475 ( .C1(n19562), .C2(n19496), .A(n19483), .B(n19482), .ZN(
        P2_U3154) );
  AOI22_X1 U22476 ( .A1(n19492), .A2(n19564), .B1(n19563), .B2(n19502), .ZN(
        n19485) );
  AOI22_X1 U22477 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19493), .B1(
        n19521), .B2(n19565), .ZN(n19484) );
  OAI211_X1 U22478 ( .C1(n19568), .C2(n19496), .A(n19485), .B(n19484), .ZN(
        P2_U3155) );
  AOI22_X1 U22479 ( .A1(n19492), .A2(n19570), .B1(n19569), .B2(n19502), .ZN(
        n19487) );
  AOI22_X1 U22480 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19493), .B1(
        n19521), .B2(n19571), .ZN(n19486) );
  OAI211_X1 U22481 ( .C1(n19574), .C2(n19496), .A(n19487), .B(n19486), .ZN(
        P2_U3156) );
  AOI22_X1 U22482 ( .A1(n19492), .A2(n19576), .B1(n19575), .B2(n19502), .ZN(
        n19489) );
  AOI22_X1 U22483 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19493), .B1(
        n19521), .B2(n19577), .ZN(n19488) );
  OAI211_X1 U22484 ( .C1(n19580), .C2(n19496), .A(n19489), .B(n19488), .ZN(
        P2_U3157) );
  AOI22_X1 U22485 ( .A1(n19492), .A2(n19582), .B1(n19581), .B2(n19502), .ZN(
        n19491) );
  AOI22_X1 U22486 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19493), .B1(
        n19521), .B2(n19583), .ZN(n19490) );
  OAI211_X1 U22487 ( .C1(n19586), .C2(n19496), .A(n19491), .B(n19490), .ZN(
        P2_U3158) );
  AOI22_X1 U22488 ( .A1(n19492), .A2(n19589), .B1(n19587), .B2(n19502), .ZN(
        n19495) );
  AOI22_X1 U22489 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19493), .B1(
        n19521), .B2(n19591), .ZN(n19494) );
  OAI211_X1 U22490 ( .C1(n19597), .C2(n19496), .A(n19495), .B(n19494), .ZN(
        P2_U3159) );
  NOR3_X2 U22491 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19693), .A3(
        n19542), .ZN(n19527) );
  AOI22_X1 U22492 ( .A1(n19521), .A2(n19499), .B1(n19527), .B2(n19539), .ZN(
        n19510) );
  INV_X1 U22493 ( .A(n12281), .ZN(n19500) );
  AOI21_X1 U22494 ( .B1(n19500), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19504) );
  AOI21_X1 U22495 ( .B1(n19596), .B2(n19533), .A(n19682), .ZN(n19501) );
  NOR2_X1 U22496 ( .A1(n19501), .A2(n19683), .ZN(n19505) );
  NOR2_X1 U22497 ( .A1(n19527), .A2(n19502), .ZN(n19507) );
  NAND2_X1 U22498 ( .A1(n19505), .A2(n19507), .ZN(n19503) );
  OAI211_X1 U22499 ( .C1(n19527), .C2(n19504), .A(n19503), .B(n19544), .ZN(
        n19530) );
  INV_X1 U22500 ( .A(n19505), .ZN(n19508) );
  OAI21_X1 U22501 ( .B1(n12281), .B2(n19527), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19506) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19530), .B1(
        n19034), .B2(n19529), .ZN(n19509) );
  OAI211_X1 U22503 ( .C1(n19511), .C2(n19596), .A(n19510), .B(n19509), .ZN(
        P2_U3160) );
  AOI22_X1 U22504 ( .A1(n19528), .A2(n19553), .B1(n19551), .B2(n19527), .ZN(
        n19513) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19530), .B1(
        n19552), .B2(n19529), .ZN(n19512) );
  OAI211_X1 U22506 ( .C1(n19556), .C2(n19533), .A(n19513), .B(n19512), .ZN(
        P2_U3161) );
  AOI22_X1 U22507 ( .A1(n19528), .A2(n19559), .B1(n19557), .B2(n19527), .ZN(
        n19515) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19530), .B1(
        n19558), .B2(n19529), .ZN(n19514) );
  OAI211_X1 U22509 ( .C1(n19562), .C2(n19533), .A(n19515), .B(n19514), .ZN(
        P2_U3162) );
  AOI22_X1 U22510 ( .A1(n19528), .A2(n19565), .B1(n19563), .B2(n19527), .ZN(
        n19517) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19530), .B1(
        n19564), .B2(n19529), .ZN(n19516) );
  OAI211_X1 U22512 ( .C1(n19568), .C2(n19533), .A(n19517), .B(n19516), .ZN(
        P2_U3163) );
  AOI22_X1 U22513 ( .A1(n19528), .A2(n19571), .B1(n19569), .B2(n19527), .ZN(
        n19519) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19530), .B1(
        n19570), .B2(n19529), .ZN(n19518) );
  OAI211_X1 U22515 ( .C1(n19574), .C2(n19533), .A(n19519), .B(n19518), .ZN(
        P2_U3164) );
  AOI22_X1 U22516 ( .A1(n19521), .A2(n19520), .B1(n19575), .B2(n19527), .ZN(
        n19523) );
  AOI22_X1 U22517 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19530), .B1(
        n19576), .B2(n19529), .ZN(n19522) );
  OAI211_X1 U22518 ( .C1(n19524), .C2(n19596), .A(n19523), .B(n19522), .ZN(
        P2_U3165) );
  AOI22_X1 U22519 ( .A1(n19528), .A2(n19583), .B1(n19527), .B2(n19581), .ZN(
        n19526) );
  AOI22_X1 U22520 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19530), .B1(
        n19582), .B2(n19529), .ZN(n19525) );
  OAI211_X1 U22521 ( .C1(n19586), .C2(n19533), .A(n19526), .B(n19525), .ZN(
        P2_U3166) );
  AOI22_X1 U22522 ( .A1(n19528), .A2(n19591), .B1(n19587), .B2(n19527), .ZN(
        n19532) );
  AOI22_X1 U22523 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19530), .B1(
        n19589), .B2(n19529), .ZN(n19531) );
  OAI211_X1 U22524 ( .C1(n19597), .C2(n19533), .A(n19532), .B(n19531), .ZN(
        P2_U3167) );
  NAND3_X1 U22525 ( .A1(n19535), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19534), 
        .ZN(n19543) );
  NAND2_X1 U22526 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19536), .ZN(
        n19537) );
  OAI21_X1 U22527 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19537), .A(n19733), 
        .ZN(n19538) );
  AND2_X1 U22528 ( .A1(n19543), .A2(n19538), .ZN(n19590) );
  AOI22_X1 U22529 ( .A1(n19590), .A2(n19034), .B1(n19588), .B2(n19539), .ZN(
        n19549) );
  NOR3_X1 U22530 ( .A1(n19541), .A2(P2_STATE2_REG_3__SCAN_IN), .A3(n19540), 
        .ZN(n19546) );
  NOR3_X1 U22531 ( .A1(n19717), .A2(n19693), .A3(n19542), .ZN(n19545) );
  OAI211_X1 U22532 ( .C1(n19546), .C2(n19545), .A(n19544), .B(n19543), .ZN(
        n19593) );
  AOI22_X1 U22533 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19593), .B1(
        n19592), .B2(n19547), .ZN(n19548) );
  OAI211_X1 U22534 ( .C1(n19550), .C2(n19596), .A(n19549), .B(n19548), .ZN(
        P2_U3168) );
  AOI22_X1 U22535 ( .A1(n19590), .A2(n19552), .B1(n19588), .B2(n19551), .ZN(
        n19555) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19593), .B1(
        n19592), .B2(n19553), .ZN(n19554) );
  OAI211_X1 U22537 ( .C1(n19556), .C2(n19596), .A(n19555), .B(n19554), .ZN(
        P2_U3169) );
  AOI22_X1 U22538 ( .A1(n19590), .A2(n19558), .B1(n19588), .B2(n19557), .ZN(
        n19561) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19593), .B1(
        n19592), .B2(n19559), .ZN(n19560) );
  OAI211_X1 U22540 ( .C1(n19562), .C2(n19596), .A(n19561), .B(n19560), .ZN(
        P2_U3170) );
  AOI22_X1 U22541 ( .A1(n19590), .A2(n19564), .B1(n19588), .B2(n19563), .ZN(
        n19567) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19593), .B1(
        n19592), .B2(n19565), .ZN(n19566) );
  OAI211_X1 U22543 ( .C1(n19568), .C2(n19596), .A(n19567), .B(n19566), .ZN(
        P2_U3171) );
  AOI22_X1 U22544 ( .A1(n19590), .A2(n19570), .B1(n19588), .B2(n19569), .ZN(
        n19573) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19593), .B1(
        n19592), .B2(n19571), .ZN(n19572) );
  OAI211_X1 U22546 ( .C1(n19574), .C2(n19596), .A(n19573), .B(n19572), .ZN(
        P2_U3172) );
  AOI22_X1 U22547 ( .A1(n19590), .A2(n19576), .B1(n19588), .B2(n19575), .ZN(
        n19579) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19593), .B1(
        n19592), .B2(n19577), .ZN(n19578) );
  OAI211_X1 U22549 ( .C1(n19580), .C2(n19596), .A(n19579), .B(n19578), .ZN(
        P2_U3173) );
  AOI22_X1 U22550 ( .A1(n19590), .A2(n19582), .B1(n19588), .B2(n19581), .ZN(
        n19585) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19593), .B1(
        n19592), .B2(n19583), .ZN(n19584) );
  OAI211_X1 U22552 ( .C1(n19586), .C2(n19596), .A(n19585), .B(n19584), .ZN(
        P2_U3174) );
  AOI22_X1 U22553 ( .A1(n19590), .A2(n19589), .B1(n19588), .B2(n19587), .ZN(
        n19595) );
  AOI22_X1 U22554 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19593), .B1(
        n19592), .B2(n19591), .ZN(n19594) );
  OAI211_X1 U22555 ( .C1(n19597), .C2(n19596), .A(n19595), .B(n19594), .ZN(
        P2_U3175) );
  AOI21_X1 U22556 ( .B1(n19600), .B2(n19599), .A(n19598), .ZN(n19607) );
  INV_X1 U22557 ( .A(n19608), .ZN(n19603) );
  AOI211_X1 U22558 ( .C1(n19603), .C2(n19602), .A(n19740), .B(n19601), .ZN(
        n19604) );
  INV_X1 U22559 ( .A(n19604), .ZN(n19605) );
  OAI211_X1 U22560 ( .C1(n19608), .C2(n19607), .A(n19606), .B(n19605), .ZN(
        P2_U3177) );
  AND2_X1 U22561 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19609), .ZN(
        P2_U3179) );
  AND2_X1 U22562 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19609), .ZN(
        P2_U3180) );
  INV_X1 U22563 ( .A(P2_DATAWIDTH_REG_29__SCAN_IN), .ZN(n20723) );
  NOR2_X1 U22564 ( .A1(n20723), .A2(n19673), .ZN(P2_U3181) );
  AND2_X1 U22565 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19609), .ZN(
        P2_U3182) );
  AND2_X1 U22566 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19609), .ZN(
        P2_U3183) );
  AND2_X1 U22567 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19609), .ZN(
        P2_U3184) );
  AND2_X1 U22568 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19609), .ZN(
        P2_U3185) );
  AND2_X1 U22569 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19609), .ZN(
        P2_U3186) );
  AND2_X1 U22570 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19609), .ZN(
        P2_U3187) );
  AND2_X1 U22571 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19609), .ZN(
        P2_U3188) );
  AND2_X1 U22572 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19609), .ZN(
        P2_U3189) );
  AND2_X1 U22573 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19609), .ZN(
        P2_U3190) );
  AND2_X1 U22574 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19609), .ZN(
        P2_U3191) );
  AND2_X1 U22575 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19609), .ZN(
        P2_U3192) );
  AND2_X1 U22576 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19609), .ZN(
        P2_U3193) );
  AND2_X1 U22577 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19609), .ZN(
        P2_U3194) );
  AND2_X1 U22578 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19609), .ZN(
        P2_U3195) );
  AND2_X1 U22579 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19609), .ZN(
        P2_U3196) );
  AND2_X1 U22580 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19609), .ZN(
        P2_U3197) );
  AND2_X1 U22581 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19609), .ZN(
        P2_U3198) );
  AND2_X1 U22582 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19609), .ZN(
        P2_U3199) );
  AND2_X1 U22583 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19609), .ZN(
        P2_U3200) );
  AND2_X1 U22584 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19609), .ZN(P2_U3201) );
  AND2_X1 U22585 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19609), .ZN(P2_U3202) );
  AND2_X1 U22586 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19609), .ZN(P2_U3203) );
  AND2_X1 U22587 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19609), .ZN(P2_U3204) );
  AND2_X1 U22588 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19609), .ZN(P2_U3205) );
  AND2_X1 U22589 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19609), .ZN(P2_U3206) );
  AND2_X1 U22590 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19609), .ZN(P2_U3207) );
  AND2_X1 U22591 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19609), .ZN(P2_U3208) );
  OAI21_X1 U22592 ( .B1(n20592), .B2(n19614), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19623) );
  INV_X1 U22593 ( .A(n19623), .ZN(n19612) );
  NAND2_X1 U22594 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19738), .ZN(n19621) );
  INV_X1 U22595 ( .A(n19621), .ZN(n19613) );
  INV_X1 U22596 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19750) );
  NOR3_X1 U22597 ( .A1(n19613), .A2(n19750), .A3(n20805), .ZN(n19611) );
  OAI21_X1 U22598 ( .B1(HOLD), .B2(n19750), .A(n19618), .ZN(n19610) );
  OAI22_X1 U22599 ( .A1(n19612), .A2(n19611), .B1(n19752), .B2(n19610), .ZN(
        P2_U3209) );
  NOR2_X1 U22600 ( .A1(n19744), .A2(n19613), .ZN(n19616) );
  NOR2_X1 U22601 ( .A1(HOLD), .A2(n20805), .ZN(n19622) );
  OAI211_X1 U22602 ( .C1(n19622), .C2(n19624), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .B(n19614), .ZN(n19615) );
  OAI211_X1 U22603 ( .C1(n19617), .C2(n20595), .A(n19616), .B(n19615), .ZN(
        P2_U3210) );
  OAI22_X1 U22604 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19618), .B1(NA), 
        .B2(n19621), .ZN(n19619) );
  OAI211_X1 U22605 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19619), .ZN(n19620) );
  OAI221_X1 U22606 ( .B1(n19623), .B2(n19622), .C1(n19623), .C2(n19621), .A(
        n19620), .ZN(P2_U3211) );
  NAND2_X1 U22607 ( .A1(n19752), .A2(n19624), .ZN(n19665) );
  CLKBUF_X1 U22608 ( .A(n19665), .Z(n19661) );
  OAI222_X1 U22609 ( .A1(n19661), .A2(n13818), .B1(n19625), .B2(n19752), .C1(
        n10247), .C2(n19662), .ZN(P2_U3212) );
  OAI222_X1 U22610 ( .A1(n19665), .A2(n10536), .B1(n19626), .B2(n19752), .C1(
        n13818), .C2(n19662), .ZN(P2_U3213) );
  OAI222_X1 U22611 ( .A1(n19665), .A2(n10551), .B1(n19627), .B2(n19752), .C1(
        n10536), .C2(n19662), .ZN(P2_U3214) );
  OAI222_X1 U22612 ( .A1(n19665), .A2(n10328), .B1(n19628), .B2(n19752), .C1(
        n10551), .C2(n19662), .ZN(P2_U3215) );
  OAI222_X1 U22613 ( .A1(n19665), .A2(n10332), .B1(n19629), .B2(n19752), .C1(
        n10328), .C2(n19662), .ZN(P2_U3216) );
  OAI222_X1 U22614 ( .A1(n19665), .A2(n10335), .B1(n19630), .B2(n19752), .C1(
        n10332), .C2(n19662), .ZN(P2_U3217) );
  OAI222_X1 U22615 ( .A1(n19661), .A2(n10620), .B1(n19631), .B2(n19752), .C1(
        n10335), .C2(n19662), .ZN(P2_U3218) );
  OAI222_X1 U22616 ( .A1(n19661), .A2(n10638), .B1(n19632), .B2(n19752), .C1(
        n10620), .C2(n19662), .ZN(P2_U3219) );
  OAI222_X1 U22617 ( .A1(n19661), .A2(n10659), .B1(n19633), .B2(n19752), .C1(
        n10638), .C2(n19662), .ZN(P2_U3220) );
  OAI222_X1 U22618 ( .A1(n19661), .A2(n10676), .B1(n19634), .B2(n19752), .C1(
        n10659), .C2(n19662), .ZN(P2_U3221) );
  OAI222_X1 U22619 ( .A1(n19661), .A2(n10693), .B1(n19635), .B2(n19752), .C1(
        n10676), .C2(n19662), .ZN(P2_U3222) );
  OAI222_X1 U22620 ( .A1(n19661), .A2(n10711), .B1(n19636), .B2(n19752), .C1(
        n10693), .C2(n19662), .ZN(P2_U3223) );
  OAI222_X1 U22621 ( .A1(n19665), .A2(n10729), .B1(n19637), .B2(n19752), .C1(
        n10711), .C2(n19662), .ZN(P2_U3224) );
  OAI222_X1 U22622 ( .A1(n19665), .A2(n10456), .B1(n19638), .B2(n19752), .C1(
        n10729), .C2(n19662), .ZN(P2_U3225) );
  OAI222_X1 U22623 ( .A1(n19665), .A2(n10732), .B1(n19639), .B2(n19752), .C1(
        n10456), .C2(n19662), .ZN(P2_U3226) );
  OAI222_X1 U22624 ( .A1(n19665), .A2(n19641), .B1(n19640), .B2(n19752), .C1(
        n10732), .C2(n19662), .ZN(P2_U3227) );
  OAI222_X1 U22625 ( .A1(n19665), .A2(n19643), .B1(n19642), .B2(n19752), .C1(
        n19641), .C2(n19662), .ZN(P2_U3228) );
  OAI222_X1 U22626 ( .A1(n19665), .A2(n19645), .B1(n19644), .B2(n19752), .C1(
        n19643), .C2(n19662), .ZN(P2_U3229) );
  OAI222_X1 U22627 ( .A1(n19661), .A2(n19647), .B1(n19646), .B2(n19752), .C1(
        n19645), .C2(n19662), .ZN(P2_U3230) );
  OAI222_X1 U22628 ( .A1(n19661), .A2(n19649), .B1(n19648), .B2(n19752), .C1(
        n19647), .C2(n19662), .ZN(P2_U3231) );
  OAI222_X1 U22629 ( .A1(n19661), .A2(n10741), .B1(n19650), .B2(n19752), .C1(
        n19649), .C2(n19662), .ZN(P2_U3232) );
  OAI222_X1 U22630 ( .A1(n19661), .A2(n10377), .B1(n19651), .B2(n19752), .C1(
        n10741), .C2(n19662), .ZN(P2_U3233) );
  OAI222_X1 U22631 ( .A1(n19661), .A2(n10381), .B1(n19652), .B2(n19752), .C1(
        n10377), .C2(n19662), .ZN(P2_U3234) );
  OAI222_X1 U22632 ( .A1(n19661), .A2(n19654), .B1(n19653), .B2(n19752), .C1(
        n10381), .C2(n19662), .ZN(P2_U3235) );
  OAI222_X1 U22633 ( .A1(n19661), .A2(n14958), .B1(n19655), .B2(n19752), .C1(
        n19654), .C2(n19662), .ZN(P2_U3236) );
  OAI222_X1 U22634 ( .A1(n19661), .A2(n19658), .B1(n19656), .B2(n19752), .C1(
        n14958), .C2(n19662), .ZN(P2_U3237) );
  OAI222_X1 U22635 ( .A1(n19662), .A2(n19658), .B1(n19657), .B2(n19752), .C1(
        n10398), .C2(n19661), .ZN(P2_U3238) );
  OAI222_X1 U22636 ( .A1(n19661), .A2(n19659), .B1(n20719), .B2(n19752), .C1(
        n10398), .C2(n19662), .ZN(P2_U3239) );
  OAI222_X1 U22637 ( .A1(n19661), .A2(n14007), .B1(n19660), .B2(n19752), .C1(
        n19659), .C2(n19662), .ZN(P2_U3240) );
  OAI222_X1 U22638 ( .A1(n19665), .A2(n19664), .B1(n19663), .B2(n19752), .C1(
        n14007), .C2(n19662), .ZN(P2_U3241) );
  OAI22_X1 U22639 ( .A1(n19753), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19752), .ZN(n19666) );
  INV_X1 U22640 ( .A(n19666), .ZN(P2_U3585) );
  OAI22_X1 U22641 ( .A1(n19753), .A2(P2_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P2_BE_N_REG_2__SCAN_IN), .B2(n19752), .ZN(n19667) );
  INV_X1 U22642 ( .A(n19667), .ZN(P2_U3586) );
  OAI22_X1 U22643 ( .A1(n19753), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19752), .ZN(n19668) );
  INV_X1 U22644 ( .A(n19668), .ZN(P2_U3587) );
  OAI22_X1 U22645 ( .A1(n19753), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19752), .ZN(n19669) );
  INV_X1 U22646 ( .A(n19669), .ZN(P2_U3588) );
  OAI21_X1 U22647 ( .B1(n19673), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19671), 
        .ZN(n19670) );
  INV_X1 U22648 ( .A(n19670), .ZN(P2_U3591) );
  OAI21_X1 U22649 ( .B1(n19673), .B2(n19672), .A(n19671), .ZN(P2_U3592) );
  INV_X1 U22650 ( .A(n19674), .ZN(n19677) );
  OAI222_X1 U22651 ( .A1(n19696), .A2(n19678), .B1(n19685), .B2(n19677), .C1(
        n19676), .C2(n19675), .ZN(n19680) );
  MUX2_X1 U22652 ( .A(n19681), .B(n19680), .S(n19679), .Z(P2_U3599) );
  NOR2_X1 U22653 ( .A1(n19683), .A2(n19682), .ZN(n19701) );
  NAND2_X1 U22654 ( .A1(n19684), .A2(n19701), .ZN(n19694) );
  NAND3_X1 U22655 ( .A1(n19706), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19685), 
        .ZN(n19686) );
  NAND2_X1 U22656 ( .A1(n19686), .A2(n19712), .ZN(n19695) );
  NAND2_X1 U22657 ( .A1(n19694), .A2(n19695), .ZN(n19691) );
  AOI222_X1 U22658 ( .A1(n19691), .A2(n19690), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19689), .C1(n19688), .C2(n19687), .ZN(n19692) );
  AOI22_X1 U22659 ( .A1(n19711), .A2(n19693), .B1(n19692), .B2(n19721), .ZN(
        P2_U3602) );
  OAI21_X1 U22660 ( .B1(n19696), .B2(n19695), .A(n19694), .ZN(n19697) );
  AOI21_X1 U22661 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19698), .A(n19697), 
        .ZN(n19699) );
  AOI22_X1 U22662 ( .A1(n19711), .A2(n19700), .B1(n19699), .B2(n19721), .ZN(
        P2_U3603) );
  INV_X1 U22663 ( .A(n19701), .ZN(n19705) );
  INV_X1 U22664 ( .A(n19702), .ZN(n19703) );
  NAND3_X1 U22665 ( .A1(n19706), .A2(n19712), .A3(n19703), .ZN(n19704) );
  OAI21_X1 U22666 ( .B1(n19706), .B2(n19705), .A(n19704), .ZN(n19707) );
  AOI21_X1 U22667 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19708), .A(n19707), 
        .ZN(n19709) );
  AOI22_X1 U22668 ( .A1(n19711), .A2(n19710), .B1(n19709), .B2(n19721), .ZN(
        P2_U3604) );
  INV_X1 U22669 ( .A(n19712), .ZN(n19715) );
  OAI22_X1 U22670 ( .A1(n19716), .A2(n19715), .B1(n19714), .B2(n19713), .ZN(
        n19718) );
  OAI21_X1 U22671 ( .B1(n19718), .B2(n19717), .A(n19721), .ZN(n19719) );
  OAI21_X1 U22672 ( .B1(n19721), .B2(n19720), .A(n19719), .ZN(P2_U3605) );
  INV_X1 U22673 ( .A(P2_READREQUEST_REG_SCAN_IN), .ZN(n20712) );
  OAI22_X1 U22674 ( .A1(n19753), .A2(n20712), .B1(P2_W_R_N_REG_SCAN_IN), .B2(
        n19752), .ZN(n19722) );
  INV_X1 U22675 ( .A(n19722), .ZN(P2_U3608) );
  INV_X1 U22676 ( .A(n19723), .ZN(n19726) );
  OAI22_X1 U22677 ( .A1(n19727), .A2(n19726), .B1(n19725), .B2(n19724), .ZN(
        n19728) );
  OR2_X1 U22678 ( .A1(n19729), .A2(n19728), .ZN(n19731) );
  MUX2_X1 U22679 ( .A(P2_MORE_REG_SCAN_IN), .B(n19731), .S(n19730), .Z(
        P2_U3609) );
  OAI21_X1 U22680 ( .B1(n19734), .B2(n19733), .A(n19732), .ZN(n19736) );
  OAI211_X1 U22681 ( .C1(n19738), .C2(n19737), .A(n19736), .B(n19735), .ZN(
        n19751) );
  AOI21_X1 U22682 ( .B1(n19740), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n19739), 
        .ZN(n19748) );
  NOR3_X1 U22683 ( .A1(n19744), .A2(n19742), .A3(n19741), .ZN(n19746) );
  AOI21_X1 U22684 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19744), .A(n19743), 
        .ZN(n19745) );
  MUX2_X1 U22685 ( .A(n19746), .B(n19745), .S(n10264), .Z(n19747) );
  OAI21_X1 U22686 ( .B1(n19748), .B2(n19747), .A(n19751), .ZN(n19749) );
  OAI21_X1 U22687 ( .B1(n19751), .B2(n19750), .A(n19749), .ZN(P2_U3610) );
  OAI22_X1 U22688 ( .A1(n19753), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19752), .ZN(n19754) );
  INV_X1 U22689 ( .A(n19754), .ZN(P2_U3611) );
  AOI21_X1 U22690 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20599), .A(n20584), 
        .ZN(n19761) );
  INV_X1 U22691 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19755) );
  NAND2_X1 U22692 ( .A1(n20584), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20687) );
  INV_X1 U22693 ( .A(n20687), .ZN(n20598) );
  AOI21_X1 U22694 ( .B1(n19761), .B2(n19755), .A(n20598), .ZN(P1_U2802) );
  OAI21_X1 U22695 ( .B1(n19757), .B2(n19756), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19758) );
  OAI21_X1 U22696 ( .B1(n19759), .B2(n20578), .A(n19758), .ZN(P1_U2803) );
  NOR2_X1 U22697 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19762) );
  OAI21_X1 U22698 ( .B1(n19762), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20673), .ZN(
        n19760) );
  OAI21_X1 U22699 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20673), .A(n19760), 
        .ZN(P1_U2804) );
  NOR2_X1 U22700 ( .A1(n20598), .A2(n19761), .ZN(n20648) );
  OAI21_X1 U22701 ( .B1(BS16), .B2(n19762), .A(n20648), .ZN(n20646) );
  OAI21_X1 U22702 ( .B1(n20648), .B2(n20468), .A(n20646), .ZN(P1_U2805) );
  AOI21_X1 U22703 ( .B1(n19763), .B2(P1_FLUSH_REG_SCAN_IN), .A(n19930), .ZN(
        n19764) );
  INV_X1 U22704 ( .A(n19764), .ZN(P1_U2806) );
  NOR4_X1 U22705 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19768) );
  NOR4_X1 U22706 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19767) );
  NOR4_X1 U22707 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19766) );
  NOR4_X1 U22708 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19765) );
  NAND4_X1 U22709 ( .A1(n19768), .A2(n19767), .A3(n19766), .A4(n19765), .ZN(
        n19774) );
  NOR4_X1 U22710 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n19772) );
  AOI211_X1 U22711 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_15__SCAN_IN), .B(
        P1_DATAWIDTH_REG_20__SCAN_IN), .ZN(n19771) );
  NOR4_X1 U22712 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_11__SCAN_IN), .A3(P1_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n19770) );
  NOR4_X1 U22713 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n19769) );
  NAND4_X1 U22714 ( .A1(n19772), .A2(n19771), .A3(n19770), .A4(n19769), .ZN(
        n19773) );
  NOR2_X1 U22715 ( .A1(n19774), .A2(n19773), .ZN(n20672) );
  INV_X1 U22716 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19776) );
  NOR3_X1 U22717 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19777) );
  OAI21_X1 U22718 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19777), .A(n20672), .ZN(
        n19775) );
  OAI21_X1 U22719 ( .B1(n20672), .B2(n19776), .A(n19775), .ZN(P1_U2807) );
  INV_X1 U22720 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20647) );
  AOI21_X1 U22721 ( .B1(n13624), .B2(n20647), .A(n19777), .ZN(n19778) );
  INV_X1 U22722 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20641) );
  INV_X1 U22723 ( .A(n20672), .ZN(n20667) );
  AOI22_X1 U22724 ( .A1(n20672), .A2(n19778), .B1(n20641), .B2(n20667), .ZN(
        P1_U2808) );
  AOI22_X1 U22725 ( .A1(n19816), .A2(n19779), .B1(n19818), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n19788) );
  OAI22_X1 U22726 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19781), .B1(n19780), 
        .B2(n19791), .ZN(n19782) );
  AOI211_X1 U22727 ( .C1(n19815), .C2(n19842), .A(n19950), .B(n19782), .ZN(
        n19787) );
  INV_X1 U22728 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n19784) );
  OAI22_X1 U22729 ( .A1(n19844), .A2(n19795), .B1(n19784), .B2(n19783), .ZN(
        n19785) );
  INV_X1 U22730 ( .A(n19785), .ZN(n19786) );
  NAND3_X1 U22731 ( .A1(n19788), .A2(n19787), .A3(n19786), .ZN(P1_U2831) );
  NOR4_X1 U22732 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19820), .A3(n19819), .A4(
        n19793), .ZN(n19799) );
  INV_X1 U22733 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19790) );
  OAI22_X1 U22734 ( .A1(n19791), .A2(n19790), .B1(n19833), .B2(n19789), .ZN(
        n19798) );
  OR2_X1 U22735 ( .A1(n19819), .A2(n19792), .ZN(n19805) );
  OAI21_X1 U22736 ( .B1(n19805), .B2(n19793), .A(n19806), .ZN(n19807) );
  OAI22_X1 U22737 ( .A1(n19796), .A2(n19795), .B1(n19794), .B2(n19807), .ZN(
        n19797) );
  NOR4_X1 U22738 ( .A1(n19950), .A2(n19799), .A3(n19798), .A4(n19797), .ZN(
        n19802) );
  NAND2_X1 U22739 ( .A1(n19815), .A2(n19800), .ZN(n19801) );
  OAI211_X1 U22740 ( .C1(n19828), .C2(n19803), .A(n19802), .B(n19801), .ZN(
        P1_U2833) );
  AOI22_X1 U22741 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n19832), .B1(
        n19815), .B2(n19848), .ZN(n19813) );
  INV_X1 U22742 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n19851) );
  OAI22_X1 U22743 ( .A1(n19828), .A2(n19804), .B1(n19851), .B2(n19833), .ZN(
        n19810) );
  INV_X1 U22744 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n19808) );
  NAND2_X1 U22745 ( .A1(n19806), .A2(n19805), .ZN(n19840) );
  NAND2_X1 U22746 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19840), .ZN(n19822) );
  AOI21_X1 U22747 ( .B1(n19808), .B2(n19822), .A(n19807), .ZN(n19809) );
  AOI211_X1 U22748 ( .C1(n19811), .C2(n19849), .A(n19810), .B(n19809), .ZN(
        n19812) );
  NAND3_X1 U22749 ( .A1(n19813), .A2(n19812), .A3(n19823), .ZN(P1_U2834) );
  INV_X1 U22750 ( .A(n19814), .ZN(n19817) );
  AOI22_X1 U22751 ( .A1(n19817), .A2(n19816), .B1(n19815), .B2(n19852), .ZN(
        n19826) );
  AOI22_X1 U22752 ( .A1(n19832), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n19818), .B2(P1_EBX_REG_5__SCAN_IN), .ZN(n19825) );
  INV_X1 U22753 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20605) );
  OAI21_X1 U22754 ( .B1(n19820), .B2(n19819), .A(n20605), .ZN(n19821) );
  AOI22_X1 U22755 ( .A1(n19855), .A2(n19837), .B1(n19822), .B2(n19821), .ZN(
        n19824) );
  NAND4_X1 U22756 ( .A1(n19826), .A2(n19825), .A3(n19824), .A4(n19823), .ZN(
        P1_U2835) );
  AOI21_X1 U22757 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(n19827), .A(
        P1_REIP_REG_4__SCAN_IN), .ZN(n19841) );
  OAI22_X1 U22758 ( .A1(n19830), .A2(n19829), .B1(n19933), .B2(n19828), .ZN(
        n19831) );
  AOI211_X1 U22759 ( .C1(n19832), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n19950), .B(n19831), .ZN(n19839) );
  OAI22_X1 U22760 ( .A1(n19952), .A2(n19835), .B1(n19834), .B2(n19833), .ZN(
        n19836) );
  AOI21_X1 U22761 ( .B1(n19929), .B2(n19837), .A(n19836), .ZN(n19838) );
  OAI211_X1 U22762 ( .C1(n19841), .C2(n19840), .A(n19839), .B(n19838), .ZN(
        P1_U2836) );
  INV_X1 U22763 ( .A(n19842), .ZN(n19843) );
  OAI22_X1 U22764 ( .A1(n19844), .A2(n14322), .B1(n14329), .B2(n19843), .ZN(
        n19845) );
  INV_X1 U22765 ( .A(n19845), .ZN(n19846) );
  OAI21_X1 U22766 ( .B1(n19858), .B2(n19847), .A(n19846), .ZN(P1_U2863) );
  AOI22_X1 U22767 ( .A1(n19849), .A2(n19854), .B1(n19853), .B2(n19848), .ZN(
        n19850) );
  OAI21_X1 U22768 ( .B1(n19858), .B2(n19851), .A(n19850), .ZN(P1_U2866) );
  AOI22_X1 U22769 ( .A1(n19855), .A2(n19854), .B1(n19853), .B2(n19852), .ZN(
        n19856) );
  OAI21_X1 U22770 ( .B1(n19858), .B2(n19857), .A(n19856), .ZN(P1_U2867) );
  AOI22_X1 U22771 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19859) );
  OAI21_X1 U22772 ( .B1(n13339), .B2(n19886), .A(n19859), .ZN(P1_U2921) );
  AOI22_X1 U22773 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19860) );
  OAI21_X1 U22774 ( .B1(n14396), .B2(n19886), .A(n19860), .ZN(P1_U2922) );
  INV_X1 U22775 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n19862) );
  AOI22_X1 U22776 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19861) );
  OAI21_X1 U22777 ( .B1(n19862), .B2(n19886), .A(n19861), .ZN(P1_U2923) );
  AOI22_X1 U22778 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19863) );
  OAI21_X1 U22779 ( .B1(n14399), .B2(n19886), .A(n19863), .ZN(P1_U2924) );
  AOI22_X1 U22780 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19864) );
  OAI21_X1 U22781 ( .B1(n14402), .B2(n19886), .A(n19864), .ZN(P1_U2925) );
  INV_X1 U22782 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n19866) );
  AOI22_X1 U22783 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19865) );
  OAI21_X1 U22784 ( .B1(n19866), .B2(n19886), .A(n19865), .ZN(P1_U2926) );
  INV_X1 U22785 ( .A(P1_LWORD_REG_9__SCAN_IN), .ZN(n20769) );
  AOI22_X1 U22786 ( .A1(P1_EAX_REG_9__SCAN_IN), .A2(n19867), .B1(n19871), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n19868) );
  OAI21_X1 U22787 ( .B1(n20769), .B2(n19869), .A(n19868), .ZN(P1_U2927) );
  AOI22_X1 U22788 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19870) );
  OAI21_X1 U22789 ( .B1(n13866), .B2(n19886), .A(n19870), .ZN(P1_U2928) );
  AOI22_X1 U22790 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19872) );
  OAI21_X1 U22791 ( .B1(n11533), .B2(n19886), .A(n19872), .ZN(P1_U2929) );
  AOI22_X1 U22792 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19873) );
  OAI21_X1 U22793 ( .B1(n19874), .B2(n19886), .A(n19873), .ZN(P1_U2930) );
  AOI22_X1 U22794 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19875) );
  OAI21_X1 U22795 ( .B1(n13766), .B2(n19886), .A(n19875), .ZN(P1_U2931) );
  AOI22_X1 U22796 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19876) );
  OAI21_X1 U22797 ( .B1(n19877), .B2(n19886), .A(n19876), .ZN(P1_U2932) );
  AOI22_X1 U22798 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19878) );
  OAI21_X1 U22799 ( .B1(n19879), .B2(n19886), .A(n19878), .ZN(P1_U2933) );
  AOI22_X1 U22800 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19880) );
  OAI21_X1 U22801 ( .B1(n19881), .B2(n19886), .A(n19880), .ZN(P1_U2934) );
  AOI22_X1 U22802 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19882) );
  OAI21_X1 U22803 ( .B1(n19883), .B2(n19886), .A(n19882), .ZN(P1_U2935) );
  AOI22_X1 U22804 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n19884), .B1(n19871), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19885) );
  OAI21_X1 U22805 ( .B1(n19887), .B2(n19886), .A(n19885), .ZN(P1_U2936) );
  AOI22_X1 U22806 ( .A1(n19922), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n19916), .ZN(n19890) );
  INV_X1 U22807 ( .A(n19888), .ZN(n19889) );
  NAND2_X1 U22808 ( .A1(n19906), .A2(n19889), .ZN(n19908) );
  NAND2_X1 U22809 ( .A1(n19890), .A2(n19908), .ZN(P1_U2945) );
  AOI22_X1 U22810 ( .A1(n19922), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n19916), .ZN(n19893) );
  INV_X1 U22811 ( .A(n19891), .ZN(n19892) );
  NAND2_X1 U22812 ( .A1(n19906), .A2(n19892), .ZN(n19910) );
  NAND2_X1 U22813 ( .A1(n19893), .A2(n19910), .ZN(P1_U2946) );
  AOI22_X1 U22814 ( .A1(n19922), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n19916), .ZN(n19895) );
  NAND2_X1 U22815 ( .A1(n19906), .A2(n19894), .ZN(n19912) );
  NAND2_X1 U22816 ( .A1(n19895), .A2(n19912), .ZN(P1_U2947) );
  AOI22_X1 U22817 ( .A1(n19922), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n19916), .ZN(n19898) );
  INV_X1 U22818 ( .A(n19896), .ZN(n19897) );
  NAND2_X1 U22819 ( .A1(n19906), .A2(n19897), .ZN(n19914) );
  NAND2_X1 U22820 ( .A1(n19898), .A2(n19914), .ZN(P1_U2948) );
  AOI22_X1 U22821 ( .A1(n19922), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n19916), .ZN(n19901) );
  INV_X1 U22822 ( .A(n19899), .ZN(n19900) );
  NAND2_X1 U22823 ( .A1(n19906), .A2(n19900), .ZN(n19917) );
  NAND2_X1 U22824 ( .A1(n19901), .A2(n19917), .ZN(P1_U2949) );
  AOI22_X1 U22825 ( .A1(n19922), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n19916), .ZN(n19903) );
  NAND2_X1 U22826 ( .A1(n19906), .A2(n19902), .ZN(n19919) );
  NAND2_X1 U22827 ( .A1(n19903), .A2(n19919), .ZN(P1_U2950) );
  AOI22_X1 U22828 ( .A1(n19922), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n19916), .ZN(n19907) );
  INV_X1 U22829 ( .A(n19904), .ZN(n19905) );
  NAND2_X1 U22830 ( .A1(n19906), .A2(n19905), .ZN(n19923) );
  NAND2_X1 U22831 ( .A1(n19907), .A2(n19923), .ZN(P1_U2951) );
  AOI22_X1 U22832 ( .A1(n19922), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n19916), .ZN(n19909) );
  NAND2_X1 U22833 ( .A1(n19909), .A2(n19908), .ZN(P1_U2960) );
  AOI22_X1 U22834 ( .A1(n19922), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n19916), .ZN(n19911) );
  NAND2_X1 U22835 ( .A1(n19911), .A2(n19910), .ZN(P1_U2961) );
  AOI22_X1 U22836 ( .A1(n19922), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n19916), .ZN(n19913) );
  NAND2_X1 U22837 ( .A1(n19913), .A2(n19912), .ZN(P1_U2962) );
  AOI22_X1 U22838 ( .A1(n19922), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n19916), .ZN(n19915) );
  NAND2_X1 U22839 ( .A1(n19915), .A2(n19914), .ZN(P1_U2963) );
  AOI22_X1 U22840 ( .A1(n19922), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n19916), .ZN(n19918) );
  NAND2_X1 U22841 ( .A1(n19918), .A2(n19917), .ZN(P1_U2964) );
  AOI22_X1 U22842 ( .A1(n19922), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n19921), .ZN(n19920) );
  NAND2_X1 U22843 ( .A1(n19920), .A2(n19919), .ZN(P1_U2965) );
  AOI22_X1 U22844 ( .A1(n19922), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n19921), .ZN(n19924) );
  NAND2_X1 U22845 ( .A1(n19924), .A2(n19923), .ZN(P1_U2966) );
  AOI22_X1 U22846 ( .A1(n19925), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n19950), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n19932) );
  OAI21_X1 U22847 ( .B1(n19927), .B2(n19926), .A(n9649), .ZN(n19928) );
  INV_X1 U22848 ( .A(n19928), .ZN(n19955) );
  AOI22_X1 U22849 ( .A1(n19955), .A2(n19930), .B1(n19942), .B2(n19929), .ZN(
        n19931) );
  OAI211_X1 U22850 ( .C1(n19934), .C2(n19933), .A(n19932), .B(n19931), .ZN(
        P1_U2995) );
  OAI21_X1 U22851 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19936), .A(
        n19935), .ZN(n19997) );
  INV_X1 U22852 ( .A(n19937), .ZN(n19941) );
  NAND2_X1 U22853 ( .A1(n19939), .A2(n19938), .ZN(n19940) );
  AOI22_X1 U22854 ( .A1(n19942), .A2(n19941), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n19940), .ZN(n19943) );
  NAND2_X1 U22855 ( .A1(n19950), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n19995) );
  OAI211_X1 U22856 ( .C1(n19944), .C2(n19997), .A(n19943), .B(n19995), .ZN(
        P1_U2999) );
  INV_X1 U22857 ( .A(n19945), .ZN(n19946) );
  AND2_X1 U22858 ( .A1(n19987), .A2(n19946), .ZN(n19977) );
  NOR3_X1 U22859 ( .A1(n19947), .A2(n19977), .A3(n19970), .ZN(n19968) );
  AOI211_X1 U22860 ( .C1(n19957), .C2(n19967), .A(n19948), .B(n19963), .ZN(
        n19949) );
  AOI21_X1 U22861 ( .B1(n19950), .B2(P1_REIP_REG_4__SCAN_IN), .A(n19949), .ZN(
        n19951) );
  OAI21_X1 U22862 ( .B1(n19953), .B2(n19952), .A(n19951), .ZN(n19954) );
  AOI21_X1 U22863 ( .B1(n19955), .B2(n19973), .A(n19954), .ZN(n19956) );
  OAI21_X1 U22864 ( .B1(n19968), .B2(n19957), .A(n19956), .ZN(P1_U3027) );
  INV_X1 U22865 ( .A(n19958), .ZN(n19961) );
  INV_X1 U22866 ( .A(n19959), .ZN(n19960) );
  AOI21_X1 U22867 ( .B1(n19993), .B2(n19961), .A(n19960), .ZN(n19966) );
  OAI22_X1 U22868 ( .A1(n19963), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        n19962), .B2(n19998), .ZN(n19964) );
  INV_X1 U22869 ( .A(n19964), .ZN(n19965) );
  OAI211_X1 U22870 ( .C1(n19968), .C2(n19967), .A(n19966), .B(n19965), .ZN(
        P1_U3028) );
  NAND2_X1 U22871 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19969), .ZN(
        n19985) );
  AOI21_X1 U22872 ( .B1(n19972), .B2(n19971), .A(n19970), .ZN(n19983) );
  NAND3_X1 U22873 ( .A1(n19974), .A2(n13356), .A3(n19973), .ZN(n19981) );
  AOI21_X1 U22874 ( .B1(n19993), .B2(n19976), .A(n19975), .ZN(n19980) );
  INV_X1 U22875 ( .A(n19977), .ZN(n19979) );
  NAND4_X1 U22876 ( .A1(n19987), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19978) );
  AND4_X1 U22877 ( .A1(n19981), .A2(n19980), .A3(n19979), .A4(n19978), .ZN(
        n19982) );
  OAI221_X1 U22878 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n19985), .C1(
        n19984), .C2(n19983), .A(n19982), .ZN(P1_U3029) );
  INV_X1 U22879 ( .A(n19986), .ZN(n19994) );
  NOR3_X1 U22880 ( .A1(n19988), .A2(n19987), .A3(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19989) );
  AOI21_X1 U22881 ( .B1(n19991), .B2(n19990), .A(n19989), .ZN(n19992) );
  AOI21_X1 U22882 ( .B1(n19994), .B2(n19993), .A(n19992), .ZN(n19996) );
  OAI211_X1 U22883 ( .C1(n19998), .C2(n19997), .A(n19996), .B(n19995), .ZN(
        P1_U3031) );
  NOR2_X1 U22884 ( .A1(n20000), .A2(n19999), .ZN(P1_U3032) );
  NOR2_X2 U22885 ( .A1(n20001), .A2(n20003), .ZN(n20041) );
  NOR2_X2 U22886 ( .A1(n20003), .A2(n20002), .ZN(n20040) );
  AOI22_X1 U22887 ( .A1(DATAI_16_), .A2(n20041), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20040), .ZN(n20480) );
  INV_X1 U22888 ( .A(n20078), .ZN(n20658) );
  AOI22_X1 U22889 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20040), .B1(DATAI_24_), 
        .B2(n20041), .ZN(n20529) );
  INV_X1 U22890 ( .A(n20529), .ZN(n20477) );
  AND2_X1 U22891 ( .A1(n20005), .A2(n20042), .ZN(n20519) );
  NOR3_X1 U22892 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20055) );
  NAND2_X1 U22893 ( .A1(n20665), .A2(n20055), .ZN(n20008) );
  INV_X1 U22894 ( .A(n20008), .ZN(n20044) );
  AOI22_X1 U22895 ( .A1(n20571), .A2(n20477), .B1(n20519), .B2(n20044), .ZN(
        n20018) );
  AND2_X1 U22896 ( .A1(n20332), .A2(n20273), .ZN(n20014) );
  NAND2_X1 U22897 ( .A1(n20012), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20466) );
  OAI21_X1 U22898 ( .B1(n20074), .B2(n20571), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20006) );
  NOR2_X1 U22899 ( .A1(n9664), .A2(n20007), .ZN(n20117) );
  NAND2_X1 U22900 ( .A1(n20117), .A2(n13459), .ZN(n20015) );
  AOI22_X1 U22901 ( .A1(n20011), .A2(n20015), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20008), .ZN(n20009) );
  NOR2_X2 U22902 ( .A1(n20010), .A2(n20052), .ZN(n20520) );
  INV_X1 U22903 ( .A(n20011), .ZN(n20016) );
  INV_X1 U22904 ( .A(n20012), .ZN(n20013) );
  NAND2_X1 U22905 ( .A1(n20013), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20338) );
  INV_X1 U22906 ( .A(n20014), .ZN(n20155) );
  AOI22_X1 U22907 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20047), .B1(
        n20520), .B2(n20046), .ZN(n20017) );
  OAI211_X1 U22908 ( .C1(n20480), .C2(n20067), .A(n20018), .B(n20017), .ZN(
        P1_U3033) );
  AOI22_X1 U22909 ( .A1(DATAI_17_), .A2(n20041), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20040), .ZN(n20484) );
  AOI22_X1 U22910 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20040), .B1(DATAI_25_), 
        .B2(n20041), .ZN(n20535) );
  INV_X1 U22911 ( .A(n20535), .ZN(n20481) );
  AOI22_X1 U22912 ( .A1(n20571), .A2(n20481), .B1(n20530), .B2(n20044), .ZN(
        n20021) );
  NOR2_X2 U22913 ( .A1(n20019), .A2(n20052), .ZN(n20531) );
  AOI22_X1 U22914 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20047), .B1(
        n20531), .B2(n20046), .ZN(n20020) );
  OAI211_X1 U22915 ( .C1(n20484), .C2(n20067), .A(n20021), .B(n20020), .ZN(
        P1_U3034) );
  AOI22_X1 U22916 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20040), .B1(DATAI_26_), 
        .B2(n20041), .ZN(n20541) );
  INV_X1 U22917 ( .A(n20541), .ZN(n20485) );
  AOI22_X1 U22918 ( .A1(n20571), .A2(n20485), .B1(n20536), .B2(n20044), .ZN(
        n20024) );
  NOR2_X2 U22919 ( .A1(n20022), .A2(n20052), .ZN(n20537) );
  AOI22_X1 U22920 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20047), .B1(
        n20537), .B2(n20046), .ZN(n20023) );
  OAI211_X1 U22921 ( .C1(n20488), .C2(n20067), .A(n20024), .B(n20023), .ZN(
        P1_U3035) );
  AOI22_X1 U22922 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20040), .B1(DATAI_19_), 
        .B2(n20041), .ZN(n20492) );
  AOI22_X1 U22923 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20040), .B1(DATAI_27_), 
        .B2(n20041), .ZN(n20547) );
  INV_X1 U22924 ( .A(n20547), .ZN(n20489) );
  AOI22_X1 U22925 ( .A1(n20571), .A2(n20489), .B1(n20542), .B2(n20044), .ZN(
        n20028) );
  NOR2_X2 U22926 ( .A1(n20026), .A2(n20052), .ZN(n20543) );
  AOI22_X1 U22927 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20047), .B1(
        n20543), .B2(n20046), .ZN(n20027) );
  OAI211_X1 U22928 ( .C1(n20492), .C2(n20067), .A(n20028), .B(n20027), .ZN(
        P1_U3036) );
  AOI22_X1 U22929 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20040), .B1(DATAI_20_), 
        .B2(n20041), .ZN(n20496) );
  AOI22_X1 U22930 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20040), .B1(DATAI_28_), 
        .B2(n20041), .ZN(n20553) );
  INV_X1 U22931 ( .A(n20553), .ZN(n20493) );
  AOI22_X1 U22932 ( .A1(n20571), .A2(n20493), .B1(n20548), .B2(n20044), .ZN(
        n20031) );
  NOR2_X2 U22933 ( .A1(n20029), .A2(n20052), .ZN(n20549) );
  AOI22_X1 U22934 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20047), .B1(
        n20549), .B2(n20046), .ZN(n20030) );
  OAI211_X1 U22935 ( .C1(n20496), .C2(n20067), .A(n20031), .B(n20030), .ZN(
        P1_U3037) );
  AOI22_X1 U22936 ( .A1(DATAI_21_), .A2(n20041), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20040), .ZN(n20500) );
  AOI22_X1 U22937 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20040), .B1(DATAI_29_), 
        .B2(n20041), .ZN(n20559) );
  INV_X1 U22938 ( .A(n20559), .ZN(n20497) );
  AOI22_X1 U22939 ( .A1(n20571), .A2(n20497), .B1(n20554), .B2(n20044), .ZN(
        n20035) );
  NOR2_X2 U22940 ( .A1(n20033), .A2(n20052), .ZN(n20555) );
  AOI22_X1 U22941 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20047), .B1(
        n20555), .B2(n20046), .ZN(n20034) );
  OAI211_X1 U22942 ( .C1(n20500), .C2(n20067), .A(n20035), .B(n20034), .ZN(
        P1_U3038) );
  AOI22_X1 U22943 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20040), .B1(DATAI_22_), 
        .B2(n20041), .ZN(n20504) );
  AOI22_X1 U22944 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20040), .B1(DATAI_30_), 
        .B2(n20041), .ZN(n20565) );
  INV_X1 U22945 ( .A(n20565), .ZN(n20501) );
  AOI22_X1 U22946 ( .A1(n20571), .A2(n20501), .B1(n20560), .B2(n20044), .ZN(
        n20039) );
  NOR2_X2 U22947 ( .A1(n20037), .A2(n20052), .ZN(n20561) );
  AOI22_X1 U22948 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20047), .B1(
        n20561), .B2(n20046), .ZN(n20038) );
  OAI211_X1 U22949 ( .C1(n20504), .C2(n20067), .A(n20039), .B(n20038), .ZN(
        P1_U3039) );
  AOI22_X1 U22950 ( .A1(DATAI_31_), .A2(n20041), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20040), .ZN(n20576) );
  INV_X1 U22951 ( .A(n20576), .ZN(n20507) );
  AOI22_X1 U22952 ( .A1(n20571), .A2(n20507), .B1(n20567), .B2(n20044), .ZN(
        n20049) );
  NOR2_X2 U22953 ( .A1(n20045), .A2(n20052), .ZN(n20569) );
  AOI22_X1 U22954 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20047), .B1(
        n20569), .B2(n20046), .ZN(n20048) );
  OAI211_X1 U22955 ( .C1(n20512), .C2(n20067), .A(n20049), .B(n20048), .ZN(
        P1_U3040) );
  INV_X1 U22956 ( .A(n20050), .ZN(n20299) );
  INV_X1 U22957 ( .A(n20055), .ZN(n20051) );
  NOR2_X1 U22958 ( .A1(n20665), .A2(n20051), .ZN(n20072) );
  AOI21_X1 U22959 ( .B1(n20117), .B2(n20299), .A(n20072), .ZN(n20053) );
  OAI22_X1 U22960 ( .A1(n20053), .A2(n20515), .B1(n20051), .B2(n20581), .ZN(
        n20073) );
  AOI22_X1 U22961 ( .A1(n20520), .A2(n20073), .B1(n20519), .B2(n20072), .ZN(
        n20057) );
  OAI211_X1 U22962 ( .C1(n20118), .C2(n20302), .A(n20657), .B(n20053), .ZN(
        n20054) );
  OAI211_X1 U22963 ( .C1(n20657), .C2(n20055), .A(n20523), .B(n20054), .ZN(
        n20075) );
  INV_X1 U22964 ( .A(n20111), .ZN(n20064) );
  INV_X1 U22965 ( .A(n20480), .ZN(n20526) );
  AOI22_X1 U22966 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20075), .B1(
        n20064), .B2(n20526), .ZN(n20056) );
  OAI211_X1 U22967 ( .C1(n20529), .C2(n20067), .A(n20057), .B(n20056), .ZN(
        P1_U3041) );
  AOI22_X1 U22968 ( .A1(n20531), .A2(n20073), .B1(n20530), .B2(n20072), .ZN(
        n20059) );
  INV_X1 U22969 ( .A(n20484), .ZN(n20532) );
  AOI22_X1 U22970 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20075), .B1(
        n20064), .B2(n20532), .ZN(n20058) );
  OAI211_X1 U22971 ( .C1(n20535), .C2(n20067), .A(n20059), .B(n20058), .ZN(
        P1_U3042) );
  AOI22_X1 U22972 ( .A1(n20537), .A2(n20073), .B1(n20536), .B2(n20072), .ZN(
        n20061) );
  INV_X1 U22973 ( .A(n20488), .ZN(n20538) );
  AOI22_X1 U22974 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20075), .B1(
        n20064), .B2(n20538), .ZN(n20060) );
  OAI211_X1 U22975 ( .C1(n20541), .C2(n20067), .A(n20061), .B(n20060), .ZN(
        P1_U3043) );
  AOI22_X1 U22976 ( .A1(n20543), .A2(n20073), .B1(n20542), .B2(n20072), .ZN(
        n20063) );
  INV_X1 U22977 ( .A(n20492), .ZN(n20544) );
  AOI22_X1 U22978 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20075), .B1(
        n20064), .B2(n20544), .ZN(n20062) );
  OAI211_X1 U22979 ( .C1(n20547), .C2(n20067), .A(n20063), .B(n20062), .ZN(
        P1_U3044) );
  AOI22_X1 U22980 ( .A1(n20549), .A2(n20073), .B1(n20548), .B2(n20072), .ZN(
        n20066) );
  INV_X1 U22981 ( .A(n20496), .ZN(n20550) );
  AOI22_X1 U22982 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20075), .B1(
        n20064), .B2(n20550), .ZN(n20065) );
  OAI211_X1 U22983 ( .C1(n20553), .C2(n20067), .A(n20066), .B(n20065), .ZN(
        P1_U3045) );
  AOI22_X1 U22984 ( .A1(n20555), .A2(n20073), .B1(n20554), .B2(n20072), .ZN(
        n20069) );
  AOI22_X1 U22985 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20075), .B1(
        n20074), .B2(n20497), .ZN(n20068) );
  OAI211_X1 U22986 ( .C1(n20500), .C2(n20111), .A(n20069), .B(n20068), .ZN(
        P1_U3046) );
  AOI22_X1 U22987 ( .A1(n20561), .A2(n20073), .B1(n20560), .B2(n20072), .ZN(
        n20071) );
  AOI22_X1 U22988 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20075), .B1(
        n20074), .B2(n20501), .ZN(n20070) );
  OAI211_X1 U22989 ( .C1(n20504), .C2(n20111), .A(n20071), .B(n20070), .ZN(
        P1_U3047) );
  AOI22_X1 U22990 ( .A1(n20569), .A2(n20073), .B1(n20567), .B2(n20072), .ZN(
        n20077) );
  AOI22_X1 U22991 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20075), .B1(
        n20074), .B2(n20507), .ZN(n20076) );
  OAI211_X1 U22992 ( .C1(n20512), .C2(n20111), .A(n20077), .B(n20076), .ZN(
        P1_U3048) );
  NAND2_X1 U22993 ( .A1(n13657), .A2(n20078), .ZN(n20326) );
  INV_X1 U22994 ( .A(n20519), .ZN(n20328) );
  NAND3_X1 U22995 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20406), .A3(
        n20407), .ZN(n20122) );
  OR2_X1 U22996 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20122), .ZN(
        n20105) );
  OAI22_X1 U22997 ( .A1(n20151), .A2(n20480), .B1(n20328), .B2(n20105), .ZN(
        n20079) );
  INV_X1 U22998 ( .A(n20079), .ZN(n20086) );
  NAND2_X1 U22999 ( .A1(n20151), .A2(n20111), .ZN(n20080) );
  AOI21_X1 U23000 ( .B1(n20080), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20515), 
        .ZN(n20082) );
  NAND2_X1 U23001 ( .A1(n20117), .A2(n20470), .ZN(n20083) );
  AOI22_X1 U23002 ( .A1(n20082), .A2(n20083), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20105), .ZN(n20081) );
  OR2_X1 U23003 ( .A1(n20332), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20212) );
  NAND2_X1 U23004 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20212), .ZN(n20209) );
  NAND3_X1 U23005 ( .A1(n20335), .A2(n20081), .A3(n20209), .ZN(n20108) );
  INV_X1 U23006 ( .A(n20082), .ZN(n20084) );
  AOI22_X1 U23007 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20108), .B1(
        n20520), .B2(n20107), .ZN(n20085) );
  OAI211_X1 U23008 ( .C1(n20529), .C2(n20111), .A(n20086), .B(n20085), .ZN(
        P1_U3049) );
  INV_X1 U23009 ( .A(n20530), .ZN(n20343) );
  OAI22_X1 U23010 ( .A1(n20151), .A2(n20484), .B1(n20105), .B2(n20343), .ZN(
        n20087) );
  INV_X1 U23011 ( .A(n20087), .ZN(n20089) );
  AOI22_X1 U23012 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20108), .B1(
        n20531), .B2(n20107), .ZN(n20088) );
  OAI211_X1 U23013 ( .C1(n20535), .C2(n20111), .A(n20089), .B(n20088), .ZN(
        P1_U3050) );
  INV_X1 U23014 ( .A(n20536), .ZN(n20347) );
  OAI22_X1 U23015 ( .A1(n20111), .A2(n20541), .B1(n20105), .B2(n20347), .ZN(
        n20090) );
  INV_X1 U23016 ( .A(n20090), .ZN(n20092) );
  AOI22_X1 U23017 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20108), .B1(
        n20537), .B2(n20107), .ZN(n20091) );
  OAI211_X1 U23018 ( .C1(n20488), .C2(n20151), .A(n20092), .B(n20091), .ZN(
        P1_U3051) );
  INV_X1 U23019 ( .A(n20542), .ZN(n20351) );
  OAI22_X1 U23020 ( .A1(n20111), .A2(n20547), .B1(n20105), .B2(n20351), .ZN(
        n20093) );
  INV_X1 U23021 ( .A(n20093), .ZN(n20095) );
  AOI22_X1 U23022 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20108), .B1(
        n20543), .B2(n20107), .ZN(n20094) );
  OAI211_X1 U23023 ( .C1(n20492), .C2(n20151), .A(n20095), .B(n20094), .ZN(
        P1_U3052) );
  OAI22_X1 U23024 ( .A1(n20111), .A2(n20553), .B1(n20105), .B2(n20355), .ZN(
        n20096) );
  INV_X1 U23025 ( .A(n20096), .ZN(n20098) );
  AOI22_X1 U23026 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20108), .B1(
        n20549), .B2(n20107), .ZN(n20097) );
  OAI211_X1 U23027 ( .C1(n20496), .C2(n20151), .A(n20098), .B(n20097), .ZN(
        P1_U3053) );
  INV_X1 U23028 ( .A(n20554), .ZN(n20359) );
  OAI22_X1 U23029 ( .A1(n20151), .A2(n20500), .B1(n20105), .B2(n20359), .ZN(
        n20099) );
  INV_X1 U23030 ( .A(n20099), .ZN(n20101) );
  AOI22_X1 U23031 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20108), .B1(
        n20555), .B2(n20107), .ZN(n20100) );
  OAI211_X1 U23032 ( .C1(n20559), .C2(n20111), .A(n20101), .B(n20100), .ZN(
        P1_U3054) );
  INV_X1 U23033 ( .A(n20560), .ZN(n20363) );
  OAI22_X1 U23034 ( .A1(n20151), .A2(n20504), .B1(n20105), .B2(n20363), .ZN(
        n20102) );
  INV_X1 U23035 ( .A(n20102), .ZN(n20104) );
  AOI22_X1 U23036 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20108), .B1(
        n20561), .B2(n20107), .ZN(n20103) );
  OAI211_X1 U23037 ( .C1(n20565), .C2(n20111), .A(n20104), .B(n20103), .ZN(
        P1_U3055) );
  INV_X1 U23038 ( .A(n20567), .ZN(n20368) );
  OAI22_X1 U23039 ( .A1(n20151), .A2(n20512), .B1(n20105), .B2(n20368), .ZN(
        n20106) );
  INV_X1 U23040 ( .A(n20106), .ZN(n20110) );
  AOI22_X1 U23041 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20108), .B1(
        n20569), .B2(n20107), .ZN(n20109) );
  OAI211_X1 U23042 ( .C1(n20576), .C2(n20111), .A(n20110), .B(n20109), .ZN(
        P1_U3056) );
  INV_X1 U23043 ( .A(n20248), .ZN(n20375) );
  INV_X1 U23044 ( .A(n20376), .ZN(n20112) );
  NAND2_X1 U23045 ( .A1(n20112), .A2(n20406), .ZN(n20145) );
  OAI22_X1 U23046 ( .A1(n20151), .A2(n20529), .B1(n20328), .B2(n20145), .ZN(
        n20113) );
  INV_X1 U23047 ( .A(n20113), .ZN(n20126) );
  NOR2_X1 U23048 ( .A1(n20115), .A2(n20114), .ZN(n20513) );
  INV_X1 U23049 ( .A(n20145), .ZN(n20116) );
  AOI21_X1 U23050 ( .B1(n20117), .B2(n20513), .A(n20116), .ZN(n20124) );
  OR2_X1 U23051 ( .A1(n20118), .A2(n20521), .ZN(n20119) );
  AND2_X1 U23052 ( .A1(n20119), .A2(n20657), .ZN(n20121) );
  AOI22_X1 U23053 ( .A1(n20124), .A2(n20121), .B1(n20515), .B2(n20122), .ZN(
        n20120) );
  NAND2_X1 U23054 ( .A1(n20523), .A2(n20120), .ZN(n20148) );
  INV_X1 U23055 ( .A(n20121), .ZN(n20123) );
  OAI22_X1 U23056 ( .A1(n20124), .A2(n20123), .B1(n20581), .B2(n20122), .ZN(
        n20147) );
  AOI22_X1 U23057 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20148), .B1(
        n20520), .B2(n20147), .ZN(n20125) );
  OAI211_X1 U23058 ( .C1(n20480), .C2(n20156), .A(n20126), .B(n20125), .ZN(
        P1_U3057) );
  OAI22_X1 U23059 ( .A1(n20151), .A2(n20535), .B1(n20343), .B2(n20145), .ZN(
        n20127) );
  INV_X1 U23060 ( .A(n20127), .ZN(n20129) );
  AOI22_X1 U23061 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20148), .B1(
        n20531), .B2(n20147), .ZN(n20128) );
  OAI211_X1 U23062 ( .C1(n20484), .C2(n20156), .A(n20129), .B(n20128), .ZN(
        P1_U3058) );
  OAI22_X1 U23063 ( .A1(n20156), .A2(n20488), .B1(n20145), .B2(n20347), .ZN(
        n20130) );
  INV_X1 U23064 ( .A(n20130), .ZN(n20132) );
  AOI22_X1 U23065 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20148), .B1(
        n20537), .B2(n20147), .ZN(n20131) );
  OAI211_X1 U23066 ( .C1(n20541), .C2(n20151), .A(n20132), .B(n20131), .ZN(
        P1_U3059) );
  OAI22_X1 U23067 ( .A1(n20151), .A2(n20547), .B1(n20145), .B2(n20351), .ZN(
        n20133) );
  INV_X1 U23068 ( .A(n20133), .ZN(n20135) );
  AOI22_X1 U23069 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20148), .B1(
        n20543), .B2(n20147), .ZN(n20134) );
  OAI211_X1 U23070 ( .C1(n20492), .C2(n20156), .A(n20135), .B(n20134), .ZN(
        P1_U3060) );
  OAI22_X1 U23071 ( .A1(n20156), .A2(n20496), .B1(n20145), .B2(n20355), .ZN(
        n20136) );
  INV_X1 U23072 ( .A(n20136), .ZN(n20138) );
  AOI22_X1 U23073 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20148), .B1(
        n20549), .B2(n20147), .ZN(n20137) );
  OAI211_X1 U23074 ( .C1(n20553), .C2(n20151), .A(n20138), .B(n20137), .ZN(
        P1_U3061) );
  OAI22_X1 U23075 ( .A1(n20151), .A2(n20559), .B1(n20359), .B2(n20145), .ZN(
        n20139) );
  INV_X1 U23076 ( .A(n20139), .ZN(n20141) );
  AOI22_X1 U23077 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20148), .B1(
        n20555), .B2(n20147), .ZN(n20140) );
  OAI211_X1 U23078 ( .C1(n20500), .C2(n20156), .A(n20141), .B(n20140), .ZN(
        P1_U3062) );
  OAI22_X1 U23079 ( .A1(n20151), .A2(n20565), .B1(n20363), .B2(n20145), .ZN(
        n20142) );
  INV_X1 U23080 ( .A(n20142), .ZN(n20144) );
  AOI22_X1 U23081 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20148), .B1(
        n20561), .B2(n20147), .ZN(n20143) );
  OAI211_X1 U23082 ( .C1(n20504), .C2(n20156), .A(n20144), .B(n20143), .ZN(
        P1_U3063) );
  OAI22_X1 U23083 ( .A1(n20156), .A2(n20512), .B1(n20368), .B2(n20145), .ZN(
        n20146) );
  INV_X1 U23084 ( .A(n20146), .ZN(n20150) );
  AOI22_X1 U23085 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20148), .B1(
        n20569), .B2(n20147), .ZN(n20149) );
  OAI211_X1 U23086 ( .C1(n20576), .C2(n20151), .A(n20150), .B(n20149), .ZN(
        P1_U3064) );
  NOR2_X1 U23087 ( .A1(n13424), .A2(n20153), .ZN(n20242) );
  NAND3_X1 U23088 ( .A1(n20242), .A2(n20657), .A3(n13459), .ZN(n20154) );
  OAI21_X1 U23089 ( .B1(n20466), .B2(n20155), .A(n20154), .ZN(n20177) );
  NOR3_X1 U23090 ( .A1(n20407), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20185) );
  INV_X1 U23091 ( .A(n20185), .ZN(n20182) );
  NOR2_X1 U23092 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20182), .ZN(
        n20176) );
  AOI22_X1 U23093 ( .A1(n20520), .A2(n20177), .B1(n20519), .B2(n20176), .ZN(
        n20163) );
  INV_X1 U23094 ( .A(n20242), .ZN(n20159) );
  INV_X1 U23095 ( .A(n20206), .ZN(n20157) );
  OAI21_X1 U23096 ( .B1(n20178), .B2(n20157), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20158) );
  OAI21_X1 U23097 ( .B1(n20470), .B2(n20159), .A(n20158), .ZN(n20161) );
  AOI22_X1 U23098 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20179), .B1(
        n20178), .B2(n20477), .ZN(n20162) );
  OAI211_X1 U23099 ( .C1(n20480), .C2(n20206), .A(n20163), .B(n20162), .ZN(
        P1_U3065) );
  AOI22_X1 U23100 ( .A1(n20531), .A2(n20177), .B1(n20530), .B2(n20176), .ZN(
        n20165) );
  AOI22_X1 U23101 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20179), .B1(
        n20178), .B2(n20481), .ZN(n20164) );
  OAI211_X1 U23102 ( .C1(n20484), .C2(n20206), .A(n20165), .B(n20164), .ZN(
        P1_U3066) );
  AOI22_X1 U23103 ( .A1(n20537), .A2(n20177), .B1(n20536), .B2(n20176), .ZN(
        n20167) );
  AOI22_X1 U23104 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20179), .B1(
        n20178), .B2(n20485), .ZN(n20166) );
  OAI211_X1 U23105 ( .C1(n20488), .C2(n20206), .A(n20167), .B(n20166), .ZN(
        P1_U3067) );
  AOI22_X1 U23106 ( .A1(n20543), .A2(n20177), .B1(n20542), .B2(n20176), .ZN(
        n20169) );
  AOI22_X1 U23107 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20179), .B1(
        n20178), .B2(n20489), .ZN(n20168) );
  OAI211_X1 U23108 ( .C1(n20492), .C2(n20206), .A(n20169), .B(n20168), .ZN(
        P1_U3068) );
  AOI22_X1 U23109 ( .A1(n20549), .A2(n20177), .B1(n20548), .B2(n20176), .ZN(
        n20171) );
  AOI22_X1 U23110 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20179), .B1(
        n20178), .B2(n20493), .ZN(n20170) );
  OAI211_X1 U23111 ( .C1(n20496), .C2(n20206), .A(n20171), .B(n20170), .ZN(
        P1_U3069) );
  AOI22_X1 U23112 ( .A1(n20555), .A2(n20177), .B1(n20554), .B2(n20176), .ZN(
        n20173) );
  AOI22_X1 U23113 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20179), .B1(
        n20178), .B2(n20497), .ZN(n20172) );
  OAI211_X1 U23114 ( .C1(n20500), .C2(n20206), .A(n20173), .B(n20172), .ZN(
        P1_U3070) );
  AOI22_X1 U23115 ( .A1(n20561), .A2(n20177), .B1(n20560), .B2(n20176), .ZN(
        n20175) );
  AOI22_X1 U23116 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20179), .B1(
        n20178), .B2(n20501), .ZN(n20174) );
  OAI211_X1 U23117 ( .C1(n20504), .C2(n20206), .A(n20175), .B(n20174), .ZN(
        P1_U3071) );
  AOI22_X1 U23118 ( .A1(n20569), .A2(n20177), .B1(n20567), .B2(n20176), .ZN(
        n20181) );
  AOI22_X1 U23119 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20179), .B1(
        n20178), .B2(n20507), .ZN(n20180) );
  OAI211_X1 U23120 ( .C1(n20512), .C2(n20206), .A(n20181), .B(n20180), .ZN(
        P1_U3072) );
  NOR2_X1 U23121 ( .A1(n20665), .A2(n20182), .ZN(n20200) );
  AOI21_X1 U23122 ( .B1(n20242), .B2(n20299), .A(n20200), .ZN(n20183) );
  OAI22_X1 U23123 ( .A1(n20183), .A2(n20515), .B1(n20182), .B2(n20581), .ZN(
        n20201) );
  AOI22_X1 U23124 ( .A1(n20520), .A2(n20201), .B1(n20519), .B2(n20200), .ZN(
        n20187) );
  INV_X1 U23125 ( .A(n20249), .ZN(n20245) );
  OAI21_X1 U23126 ( .B1(n20245), .B2(n20302), .A(n20183), .ZN(n20184) );
  OAI221_X1 U23127 ( .B1(n20657), .B2(n20185), .C1(n20515), .C2(n20184), .A(
        n20523), .ZN(n20203) );
  INV_X1 U23128 ( .A(n20305), .ZN(n20437) );
  AOI22_X1 U23129 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20526), .ZN(n20186) );
  OAI211_X1 U23130 ( .C1(n20529), .C2(n20206), .A(n20187), .B(n20186), .ZN(
        P1_U3073) );
  AOI22_X1 U23131 ( .A1(n20531), .A2(n20201), .B1(n20530), .B2(n20200), .ZN(
        n20189) );
  AOI22_X1 U23132 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20532), .ZN(n20188) );
  OAI211_X1 U23133 ( .C1(n20535), .C2(n20206), .A(n20189), .B(n20188), .ZN(
        P1_U3074) );
  AOI22_X1 U23134 ( .A1(n20537), .A2(n20201), .B1(n20536), .B2(n20200), .ZN(
        n20191) );
  AOI22_X1 U23135 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20538), .ZN(n20190) );
  OAI211_X1 U23136 ( .C1(n20541), .C2(n20206), .A(n20191), .B(n20190), .ZN(
        P1_U3075) );
  AOI22_X1 U23137 ( .A1(n20543), .A2(n20201), .B1(n20542), .B2(n20200), .ZN(
        n20193) );
  AOI22_X1 U23138 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20544), .ZN(n20192) );
  OAI211_X1 U23139 ( .C1(n20547), .C2(n20206), .A(n20193), .B(n20192), .ZN(
        P1_U3076) );
  AOI22_X1 U23140 ( .A1(n20549), .A2(n20201), .B1(n20548), .B2(n20200), .ZN(
        n20195) );
  AOI22_X1 U23141 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20550), .ZN(n20194) );
  OAI211_X1 U23142 ( .C1(n20553), .C2(n20206), .A(n20195), .B(n20194), .ZN(
        P1_U3077) );
  AOI22_X1 U23143 ( .A1(n20555), .A2(n20201), .B1(n20554), .B2(n20200), .ZN(
        n20197) );
  INV_X1 U23144 ( .A(n20500), .ZN(n20556) );
  AOI22_X1 U23145 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20556), .ZN(n20196) );
  OAI211_X1 U23146 ( .C1(n20559), .C2(n20206), .A(n20197), .B(n20196), .ZN(
        P1_U3078) );
  AOI22_X1 U23147 ( .A1(n20561), .A2(n20201), .B1(n20560), .B2(n20200), .ZN(
        n20199) );
  INV_X1 U23148 ( .A(n20504), .ZN(n20562) );
  AOI22_X1 U23149 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20562), .ZN(n20198) );
  OAI211_X1 U23150 ( .C1(n20565), .C2(n20206), .A(n20199), .B(n20198), .ZN(
        P1_U3079) );
  AOI22_X1 U23151 ( .A1(n20569), .A2(n20201), .B1(n20567), .B2(n20200), .ZN(
        n20205) );
  INV_X1 U23152 ( .A(n20512), .ZN(n20570) );
  AOI22_X1 U23153 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20570), .ZN(n20204) );
  OAI211_X1 U23154 ( .C1(n20576), .C2(n20206), .A(n20205), .B(n20204), .ZN(
        P1_U3080) );
  INV_X1 U23155 ( .A(n20326), .ZN(n20464) );
  INV_X1 U23156 ( .A(n20243), .ZN(n20246) );
  NAND2_X1 U23157 ( .A1(n20665), .A2(n20246), .ZN(n20235) );
  OAI22_X1 U23158 ( .A1(n20264), .A2(n20480), .B1(n20328), .B2(n20235), .ZN(
        n20207) );
  INV_X1 U23159 ( .A(n20207), .ZN(n20216) );
  NAND2_X1 U23160 ( .A1(n20264), .A2(n20241), .ZN(n20208) );
  AOI21_X1 U23161 ( .B1(n20208), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20515), 
        .ZN(n20211) );
  NAND2_X1 U23162 ( .A1(n20242), .A2(n20470), .ZN(n20213) );
  AOI22_X1 U23163 ( .A1(n20211), .A2(n20213), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20235), .ZN(n20210) );
  NAND3_X1 U23164 ( .A1(n20474), .A2(n20210), .A3(n20209), .ZN(n20238) );
  INV_X1 U23165 ( .A(n20211), .ZN(n20214) );
  OAI22_X1 U23166 ( .A1(n20214), .A2(n20213), .B1(n20212), .B2(n20466), .ZN(
        n20237) );
  AOI22_X1 U23167 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20238), .B1(
        n20520), .B2(n20237), .ZN(n20215) );
  OAI211_X1 U23168 ( .C1(n20529), .C2(n20241), .A(n20216), .B(n20215), .ZN(
        P1_U3081) );
  OAI22_X1 U23169 ( .A1(n20264), .A2(n20484), .B1(n20343), .B2(n20235), .ZN(
        n20217) );
  INV_X1 U23170 ( .A(n20217), .ZN(n20219) );
  AOI22_X1 U23171 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20238), .B1(
        n20531), .B2(n20237), .ZN(n20218) );
  OAI211_X1 U23172 ( .C1(n20535), .C2(n20241), .A(n20219), .B(n20218), .ZN(
        P1_U3082) );
  OAI22_X1 U23173 ( .A1(n20264), .A2(n20488), .B1(n20347), .B2(n20235), .ZN(
        n20220) );
  INV_X1 U23174 ( .A(n20220), .ZN(n20222) );
  AOI22_X1 U23175 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20238), .B1(
        n20537), .B2(n20237), .ZN(n20221) );
  OAI211_X1 U23176 ( .C1(n20541), .C2(n20241), .A(n20222), .B(n20221), .ZN(
        P1_U3083) );
  OAI22_X1 U23177 ( .A1(n20264), .A2(n20492), .B1(n20351), .B2(n20235), .ZN(
        n20223) );
  INV_X1 U23178 ( .A(n20223), .ZN(n20225) );
  AOI22_X1 U23179 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20238), .B1(
        n20543), .B2(n20237), .ZN(n20224) );
  OAI211_X1 U23180 ( .C1(n20547), .C2(n20241), .A(n20225), .B(n20224), .ZN(
        P1_U3084) );
  OAI22_X1 U23181 ( .A1(n20264), .A2(n20496), .B1(n20355), .B2(n20235), .ZN(
        n20226) );
  INV_X1 U23182 ( .A(n20226), .ZN(n20228) );
  AOI22_X1 U23183 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20238), .B1(
        n20549), .B2(n20237), .ZN(n20227) );
  OAI211_X1 U23184 ( .C1(n20553), .C2(n20241), .A(n20228), .B(n20227), .ZN(
        P1_U3085) );
  OAI22_X1 U23185 ( .A1(n20264), .A2(n20500), .B1(n20359), .B2(n20235), .ZN(
        n20229) );
  INV_X1 U23186 ( .A(n20229), .ZN(n20231) );
  AOI22_X1 U23187 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20238), .B1(
        n20555), .B2(n20237), .ZN(n20230) );
  OAI211_X1 U23188 ( .C1(n20559), .C2(n20241), .A(n20231), .B(n20230), .ZN(
        P1_U3086) );
  OAI22_X1 U23189 ( .A1(n20241), .A2(n20565), .B1(n20363), .B2(n20235), .ZN(
        n20232) );
  INV_X1 U23190 ( .A(n20232), .ZN(n20234) );
  AOI22_X1 U23191 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20238), .B1(
        n20561), .B2(n20237), .ZN(n20233) );
  OAI211_X1 U23192 ( .C1(n20504), .C2(n20264), .A(n20234), .B(n20233), .ZN(
        P1_U3087) );
  OAI22_X1 U23193 ( .A1(n20264), .A2(n20512), .B1(n20368), .B2(n20235), .ZN(
        n20236) );
  INV_X1 U23194 ( .A(n20236), .ZN(n20240) );
  AOI22_X1 U23195 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20238), .B1(
        n20569), .B2(n20237), .ZN(n20239) );
  OAI211_X1 U23196 ( .C1(n20576), .C2(n20241), .A(n20240), .B(n20239), .ZN(
        P1_U3088) );
  AOI21_X1 U23197 ( .B1(n20242), .B2(n20513), .A(n20265), .ZN(n20244) );
  OAI22_X1 U23198 ( .A1(n20244), .A2(n20515), .B1(n20243), .B2(n20581), .ZN(
        n20266) );
  AOI22_X1 U23199 ( .A1(n20520), .A2(n20266), .B1(n20519), .B2(n20265), .ZN(
        n20251) );
  NOR3_X1 U23200 ( .A1(n20245), .A2(n20515), .A3(n20521), .ZN(n20247) );
  OAI21_X1 U23201 ( .B1(n20247), .B2(n20246), .A(n20523), .ZN(n20268) );
  NAND2_X1 U23202 ( .A1(n20249), .A2(n20248), .ZN(n20271) );
  AOI22_X1 U23203 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20268), .B1(
        n20295), .B2(n20526), .ZN(n20250) );
  OAI211_X1 U23204 ( .C1(n20529), .C2(n20264), .A(n20251), .B(n20250), .ZN(
        P1_U3089) );
  AOI22_X1 U23205 ( .A1(n20531), .A2(n20266), .B1(n20530), .B2(n20265), .ZN(
        n20253) );
  INV_X1 U23206 ( .A(n20264), .ZN(n20267) );
  AOI22_X1 U23207 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20268), .B1(
        n20267), .B2(n20481), .ZN(n20252) );
  OAI211_X1 U23208 ( .C1(n20484), .C2(n20271), .A(n20253), .B(n20252), .ZN(
        P1_U3090) );
  AOI22_X1 U23209 ( .A1(n20537), .A2(n20266), .B1(n20536), .B2(n20265), .ZN(
        n20255) );
  AOI22_X1 U23210 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20268), .B1(
        n20267), .B2(n20485), .ZN(n20254) );
  OAI211_X1 U23211 ( .C1(n20488), .C2(n20271), .A(n20255), .B(n20254), .ZN(
        P1_U3091) );
  AOI22_X1 U23212 ( .A1(n20543), .A2(n20266), .B1(n20542), .B2(n20265), .ZN(
        n20257) );
  AOI22_X1 U23213 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20268), .B1(
        n20267), .B2(n20489), .ZN(n20256) );
  OAI211_X1 U23214 ( .C1(n20492), .C2(n20271), .A(n20257), .B(n20256), .ZN(
        P1_U3092) );
  AOI22_X1 U23215 ( .A1(n20549), .A2(n20266), .B1(n20548), .B2(n20265), .ZN(
        n20259) );
  AOI22_X1 U23216 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20268), .B1(
        n20295), .B2(n20550), .ZN(n20258) );
  OAI211_X1 U23217 ( .C1(n20553), .C2(n20264), .A(n20259), .B(n20258), .ZN(
        P1_U3093) );
  AOI22_X1 U23218 ( .A1(n20555), .A2(n20266), .B1(n20554), .B2(n20265), .ZN(
        n20261) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20268), .B1(
        n20295), .B2(n20556), .ZN(n20260) );
  OAI211_X1 U23220 ( .C1(n20559), .C2(n20264), .A(n20261), .B(n20260), .ZN(
        P1_U3094) );
  AOI22_X1 U23221 ( .A1(n20561), .A2(n20266), .B1(n20560), .B2(n20265), .ZN(
        n20263) );
  AOI22_X1 U23222 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20268), .B1(
        n20295), .B2(n20562), .ZN(n20262) );
  OAI211_X1 U23223 ( .C1(n20565), .C2(n20264), .A(n20263), .B(n20262), .ZN(
        P1_U3095) );
  AOI22_X1 U23224 ( .A1(n20569), .A2(n20266), .B1(n20567), .B2(n20265), .ZN(
        n20270) );
  AOI22_X1 U23225 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20268), .B1(
        n20267), .B2(n20507), .ZN(n20269) );
  OAI211_X1 U23226 ( .C1(n20512), .C2(n20271), .A(n20270), .B(n20269), .ZN(
        P1_U3096) );
  INV_X1 U23227 ( .A(n20380), .ZN(n20272) );
  AND2_X1 U23228 ( .A1(n9664), .A2(n13424), .ZN(n20377) );
  NOR3_X1 U23229 ( .A1(n20406), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20304) );
  INV_X1 U23230 ( .A(n20304), .ZN(n20300) );
  NOR2_X1 U23231 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20300), .ZN(
        n20293) );
  AOI21_X1 U23232 ( .B1(n20377), .B2(n13459), .A(n20293), .ZN(n20276) );
  INV_X1 U23233 ( .A(n20273), .ZN(n20274) );
  NAND2_X1 U23234 ( .A1(n20274), .A2(n20332), .ZN(n20414) );
  OAI22_X1 U23235 ( .A1(n20276), .A2(n20515), .B1(n20338), .B2(n20414), .ZN(
        n20294) );
  AOI22_X1 U23236 ( .A1(n20520), .A2(n20294), .B1(n20519), .B2(n20293), .ZN(
        n20280) );
  INV_X1 U23237 ( .A(n20325), .ZN(n20275) );
  OAI21_X1 U23238 ( .B1(n20275), .B2(n20295), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20277) );
  NAND2_X1 U23239 ( .A1(n20277), .A2(n20276), .ZN(n20278) );
  AOI22_X1 U23240 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20296), .B1(
        n20295), .B2(n20477), .ZN(n20279) );
  OAI211_X1 U23241 ( .C1(n20480), .C2(n20325), .A(n20280), .B(n20279), .ZN(
        P1_U3097) );
  AOI22_X1 U23242 ( .A1(n20531), .A2(n20294), .B1(n20530), .B2(n20293), .ZN(
        n20282) );
  AOI22_X1 U23243 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20296), .B1(
        n20295), .B2(n20481), .ZN(n20281) );
  OAI211_X1 U23244 ( .C1(n20484), .C2(n20325), .A(n20282), .B(n20281), .ZN(
        P1_U3098) );
  AOI22_X1 U23245 ( .A1(n20537), .A2(n20294), .B1(n20536), .B2(n20293), .ZN(
        n20284) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20296), .B1(
        n20295), .B2(n20485), .ZN(n20283) );
  OAI211_X1 U23247 ( .C1(n20488), .C2(n20325), .A(n20284), .B(n20283), .ZN(
        P1_U3099) );
  AOI22_X1 U23248 ( .A1(n20543), .A2(n20294), .B1(n20542), .B2(n20293), .ZN(
        n20286) );
  AOI22_X1 U23249 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20296), .B1(
        n20295), .B2(n20489), .ZN(n20285) );
  OAI211_X1 U23250 ( .C1(n20492), .C2(n20325), .A(n20286), .B(n20285), .ZN(
        P1_U3100) );
  AOI22_X1 U23251 ( .A1(n20549), .A2(n20294), .B1(n20548), .B2(n20293), .ZN(
        n20288) );
  AOI22_X1 U23252 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20296), .B1(
        n20295), .B2(n20493), .ZN(n20287) );
  OAI211_X1 U23253 ( .C1(n20496), .C2(n20325), .A(n20288), .B(n20287), .ZN(
        P1_U3101) );
  AOI22_X1 U23254 ( .A1(n20555), .A2(n20294), .B1(n20554), .B2(n20293), .ZN(
        n20290) );
  AOI22_X1 U23255 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20296), .B1(
        n20295), .B2(n20497), .ZN(n20289) );
  OAI211_X1 U23256 ( .C1(n20500), .C2(n20325), .A(n20290), .B(n20289), .ZN(
        P1_U3102) );
  AOI22_X1 U23257 ( .A1(n20561), .A2(n20294), .B1(n20560), .B2(n20293), .ZN(
        n20292) );
  AOI22_X1 U23258 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20296), .B1(
        n20295), .B2(n20501), .ZN(n20291) );
  OAI211_X1 U23259 ( .C1(n20504), .C2(n20325), .A(n20292), .B(n20291), .ZN(
        P1_U3103) );
  AOI22_X1 U23260 ( .A1(n20569), .A2(n20294), .B1(n20567), .B2(n20293), .ZN(
        n20298) );
  AOI22_X1 U23261 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20296), .B1(
        n20295), .B2(n20507), .ZN(n20297) );
  OAI211_X1 U23262 ( .C1(n20512), .C2(n20325), .A(n20298), .B(n20297), .ZN(
        P1_U3104) );
  NOR2_X1 U23263 ( .A1(n20665), .A2(n20300), .ZN(n20320) );
  AOI21_X1 U23264 ( .B1(n20377), .B2(n20299), .A(n20320), .ZN(n20301) );
  OAI22_X1 U23265 ( .A1(n20301), .A2(n20515), .B1(n20300), .B2(n20581), .ZN(
        n20321) );
  AOI22_X1 U23266 ( .A1(n20520), .A2(n20321), .B1(n20519), .B2(n20320), .ZN(
        n20307) );
  OAI211_X1 U23267 ( .C1(n20380), .C2(n20302), .A(n20657), .B(n20301), .ZN(
        n20303) );
  OAI211_X1 U23268 ( .C1(n20657), .C2(n20304), .A(n20523), .B(n20303), .ZN(
        n20322) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20322), .B1(
        n20330), .B2(n20526), .ZN(n20306) );
  OAI211_X1 U23270 ( .C1(n20529), .C2(n20325), .A(n20307), .B(n20306), .ZN(
        P1_U3105) );
  AOI22_X1 U23271 ( .A1(n20531), .A2(n20321), .B1(n20530), .B2(n20320), .ZN(
        n20309) );
  AOI22_X1 U23272 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20322), .B1(
        n20330), .B2(n20532), .ZN(n20308) );
  OAI211_X1 U23273 ( .C1(n20535), .C2(n20325), .A(n20309), .B(n20308), .ZN(
        P1_U3106) );
  AOI22_X1 U23274 ( .A1(n20537), .A2(n20321), .B1(n20536), .B2(n20320), .ZN(
        n20311) );
  AOI22_X1 U23275 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20322), .B1(
        n20330), .B2(n20538), .ZN(n20310) );
  OAI211_X1 U23276 ( .C1(n20541), .C2(n20325), .A(n20311), .B(n20310), .ZN(
        P1_U3107) );
  AOI22_X1 U23277 ( .A1(n20543), .A2(n20321), .B1(n20542), .B2(n20320), .ZN(
        n20313) );
  AOI22_X1 U23278 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20322), .B1(
        n20330), .B2(n20544), .ZN(n20312) );
  OAI211_X1 U23279 ( .C1(n20547), .C2(n20325), .A(n20313), .B(n20312), .ZN(
        P1_U3108) );
  AOI22_X1 U23280 ( .A1(n20549), .A2(n20321), .B1(n20548), .B2(n20320), .ZN(
        n20315) );
  AOI22_X1 U23281 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20322), .B1(
        n20330), .B2(n20550), .ZN(n20314) );
  OAI211_X1 U23282 ( .C1(n20553), .C2(n20325), .A(n20315), .B(n20314), .ZN(
        P1_U3109) );
  AOI22_X1 U23283 ( .A1(n20555), .A2(n20321), .B1(n20554), .B2(n20320), .ZN(
        n20317) );
  AOI22_X1 U23284 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20322), .B1(
        n20330), .B2(n20556), .ZN(n20316) );
  OAI211_X1 U23285 ( .C1(n20559), .C2(n20325), .A(n20317), .B(n20316), .ZN(
        P1_U3110) );
  AOI22_X1 U23286 ( .A1(n20561), .A2(n20321), .B1(n20560), .B2(n20320), .ZN(
        n20319) );
  AOI22_X1 U23287 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20322), .B1(
        n20330), .B2(n20562), .ZN(n20318) );
  OAI211_X1 U23288 ( .C1(n20565), .C2(n20325), .A(n20319), .B(n20318), .ZN(
        P1_U3111) );
  AOI22_X1 U23289 ( .A1(n20569), .A2(n20321), .B1(n20567), .B2(n20320), .ZN(
        n20324) );
  AOI22_X1 U23290 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20322), .B1(
        n20330), .B2(n20570), .ZN(n20323) );
  OAI211_X1 U23291 ( .C1(n20576), .C2(n20325), .A(n20324), .B(n20323), .ZN(
        P1_U3112) );
  NOR3_X1 U23292 ( .A1(n20406), .A2(n20327), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20382) );
  INV_X1 U23293 ( .A(n20382), .ZN(n20378) );
  NOR2_X1 U23294 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20378), .ZN(
        n20333) );
  INV_X1 U23295 ( .A(n20333), .ZN(n20367) );
  OAI22_X1 U23296 ( .A1(n20369), .A2(n20529), .B1(n20328), .B2(n20367), .ZN(
        n20329) );
  INV_X1 U23297 ( .A(n20329), .ZN(n20342) );
  OAI21_X1 U23298 ( .B1(n20391), .B2(n20330), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20331) );
  NAND2_X1 U23299 ( .A1(n20331), .A2(n20657), .ZN(n20340) );
  AND2_X1 U23300 ( .A1(n20377), .A2(n20470), .ZN(n20337) );
  OR2_X1 U23301 ( .A1(n20332), .A2(n20406), .ZN(n20467) );
  NAND2_X1 U23302 ( .A1(n20467), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20473) );
  OAI21_X1 U23303 ( .B1(n20412), .B2(n20333), .A(n20473), .ZN(n20334) );
  INV_X1 U23304 ( .A(n20334), .ZN(n20336) );
  OAI211_X1 U23305 ( .C1(n20340), .C2(n20337), .A(n20336), .B(n20335), .ZN(
        n20372) );
  INV_X1 U23306 ( .A(n20337), .ZN(n20339) );
  AOI22_X1 U23307 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20372), .B1(
        n20520), .B2(n20371), .ZN(n20341) );
  OAI211_X1 U23308 ( .C1(n20480), .C2(n20404), .A(n20342), .B(n20341), .ZN(
        P1_U3113) );
  OAI22_X1 U23309 ( .A1(n20404), .A2(n20484), .B1(n20343), .B2(n20367), .ZN(
        n20344) );
  INV_X1 U23310 ( .A(n20344), .ZN(n20346) );
  AOI22_X1 U23311 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20372), .B1(
        n20531), .B2(n20371), .ZN(n20345) );
  OAI211_X1 U23312 ( .C1(n20535), .C2(n20369), .A(n20346), .B(n20345), .ZN(
        P1_U3114) );
  OAI22_X1 U23313 ( .A1(n20369), .A2(n20541), .B1(n20347), .B2(n20367), .ZN(
        n20348) );
  INV_X1 U23314 ( .A(n20348), .ZN(n20350) );
  AOI22_X1 U23315 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20372), .B1(
        n20537), .B2(n20371), .ZN(n20349) );
  OAI211_X1 U23316 ( .C1(n20488), .C2(n20404), .A(n20350), .B(n20349), .ZN(
        P1_U3115) );
  OAI22_X1 U23317 ( .A1(n20369), .A2(n20547), .B1(n20351), .B2(n20367), .ZN(
        n20352) );
  INV_X1 U23318 ( .A(n20352), .ZN(n20354) );
  AOI22_X1 U23319 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20372), .B1(
        n20543), .B2(n20371), .ZN(n20353) );
  OAI211_X1 U23320 ( .C1(n20492), .C2(n20404), .A(n20354), .B(n20353), .ZN(
        P1_U3116) );
  OAI22_X1 U23321 ( .A1(n20404), .A2(n20496), .B1(n20355), .B2(n20367), .ZN(
        n20356) );
  INV_X1 U23322 ( .A(n20356), .ZN(n20358) );
  AOI22_X1 U23323 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20372), .B1(
        n20549), .B2(n20371), .ZN(n20357) );
  OAI211_X1 U23324 ( .C1(n20553), .C2(n20369), .A(n20358), .B(n20357), .ZN(
        P1_U3117) );
  OAI22_X1 U23325 ( .A1(n20369), .A2(n20559), .B1(n20359), .B2(n20367), .ZN(
        n20360) );
  INV_X1 U23326 ( .A(n20360), .ZN(n20362) );
  AOI22_X1 U23327 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20372), .B1(
        n20555), .B2(n20371), .ZN(n20361) );
  OAI211_X1 U23328 ( .C1(n20500), .C2(n20404), .A(n20362), .B(n20361), .ZN(
        P1_U3118) );
  OAI22_X1 U23329 ( .A1(n20369), .A2(n20565), .B1(n20363), .B2(n20367), .ZN(
        n20364) );
  INV_X1 U23330 ( .A(n20364), .ZN(n20366) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20372), .B1(
        n20561), .B2(n20371), .ZN(n20365) );
  OAI211_X1 U23332 ( .C1(n20504), .C2(n20404), .A(n20366), .B(n20365), .ZN(
        P1_U3119) );
  OAI22_X1 U23333 ( .A1(n20369), .A2(n20576), .B1(n20368), .B2(n20367), .ZN(
        n20370) );
  INV_X1 U23334 ( .A(n20370), .ZN(n20374) );
  AOI22_X1 U23335 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20372), .B1(
        n20569), .B2(n20371), .ZN(n20373) );
  OAI211_X1 U23336 ( .C1(n20512), .C2(n20404), .A(n20374), .B(n20373), .ZN(
        P1_U3120) );
  NOR2_X1 U23337 ( .A1(n20376), .A2(n20406), .ZN(n20398) );
  AOI21_X1 U23338 ( .B1(n20377), .B2(n20513), .A(n20398), .ZN(n20379) );
  OAI22_X1 U23339 ( .A1(n20379), .A2(n20515), .B1(n20378), .B2(n20581), .ZN(
        n20399) );
  AOI22_X1 U23340 ( .A1(n20520), .A2(n20399), .B1(n20519), .B2(n20398), .ZN(
        n20384) );
  OAI211_X1 U23341 ( .C1(n20380), .C2(n20521), .A(n20657), .B(n20379), .ZN(
        n20381) );
  OAI211_X1 U23342 ( .C1(n20657), .C2(n20382), .A(n20523), .B(n20381), .ZN(
        n20401) );
  AOI22_X1 U23343 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20401), .B1(
        n20391), .B2(n20477), .ZN(n20383) );
  OAI211_X1 U23344 ( .C1(n20480), .C2(n20436), .A(n20384), .B(n20383), .ZN(
        P1_U3121) );
  AOI22_X1 U23345 ( .A1(n20531), .A2(n20399), .B1(n20530), .B2(n20398), .ZN(
        n20386) );
  INV_X1 U23346 ( .A(n20436), .ZN(n20400) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20401), .B1(
        n20400), .B2(n20532), .ZN(n20385) );
  OAI211_X1 U23348 ( .C1(n20535), .C2(n20404), .A(n20386), .B(n20385), .ZN(
        P1_U3122) );
  AOI22_X1 U23349 ( .A1(n20537), .A2(n20399), .B1(n20536), .B2(n20398), .ZN(
        n20388) );
  AOI22_X1 U23350 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20401), .B1(
        n20391), .B2(n20485), .ZN(n20387) );
  OAI211_X1 U23351 ( .C1(n20488), .C2(n20436), .A(n20388), .B(n20387), .ZN(
        P1_U3123) );
  AOI22_X1 U23352 ( .A1(n20543), .A2(n20399), .B1(n20542), .B2(n20398), .ZN(
        n20390) );
  AOI22_X1 U23353 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20401), .B1(
        n20400), .B2(n20544), .ZN(n20389) );
  OAI211_X1 U23354 ( .C1(n20547), .C2(n20404), .A(n20390), .B(n20389), .ZN(
        P1_U3124) );
  AOI22_X1 U23355 ( .A1(n20549), .A2(n20399), .B1(n20548), .B2(n20398), .ZN(
        n20393) );
  AOI22_X1 U23356 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20401), .B1(
        n20391), .B2(n20493), .ZN(n20392) );
  OAI211_X1 U23357 ( .C1(n20496), .C2(n20436), .A(n20393), .B(n20392), .ZN(
        P1_U3125) );
  AOI22_X1 U23358 ( .A1(n20555), .A2(n20399), .B1(n20554), .B2(n20398), .ZN(
        n20395) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20401), .B1(
        n20400), .B2(n20556), .ZN(n20394) );
  OAI211_X1 U23360 ( .C1(n20559), .C2(n20404), .A(n20395), .B(n20394), .ZN(
        P1_U3126) );
  AOI22_X1 U23361 ( .A1(n20561), .A2(n20399), .B1(n20560), .B2(n20398), .ZN(
        n20397) );
  AOI22_X1 U23362 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20401), .B1(
        n20400), .B2(n20562), .ZN(n20396) );
  OAI211_X1 U23363 ( .C1(n20565), .C2(n20404), .A(n20397), .B(n20396), .ZN(
        P1_U3127) );
  AOI22_X1 U23364 ( .A1(n20569), .A2(n20399), .B1(n20567), .B2(n20398), .ZN(
        n20403) );
  AOI22_X1 U23365 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20401), .B1(
        n20400), .B2(n20570), .ZN(n20402) );
  OAI211_X1 U23366 ( .C1(n20576), .C2(n20404), .A(n20403), .B(n20402), .ZN(
        P1_U3128) );
  NOR3_X1 U23367 ( .A1(n20407), .A2(n20406), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20442) );
  INV_X1 U23368 ( .A(n20442), .ZN(n20439) );
  NOR2_X1 U23369 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20439), .ZN(
        n20431) );
  AOI22_X1 U23370 ( .A1(n20460), .A2(n20526), .B1(n20519), .B2(n20431), .ZN(
        n20418) );
  INV_X1 U23371 ( .A(n20460), .ZN(n20408) );
  AOI21_X1 U23372 ( .B1(n20408), .B2(n20436), .A(n20468), .ZN(n20409) );
  NOR2_X1 U23373 ( .A1(n20409), .A2(n20515), .ZN(n20413) );
  OR2_X1 U23374 ( .A1(n13424), .A2(n20410), .ZN(n20438) );
  OR2_X1 U23375 ( .A1(n20438), .A2(n20470), .ZN(n20415) );
  AOI22_X1 U23376 ( .A1(n20413), .A2(n20415), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20414), .ZN(n20411) );
  INV_X1 U23377 ( .A(n20413), .ZN(n20416) );
  AOI22_X1 U23378 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20433), .B1(
        n20520), .B2(n20432), .ZN(n20417) );
  OAI211_X1 U23379 ( .C1(n20529), .C2(n20436), .A(n20418), .B(n20417), .ZN(
        P1_U3129) );
  AOI22_X1 U23380 ( .A1(n20460), .A2(n20532), .B1(n20530), .B2(n20431), .ZN(
        n20420) );
  AOI22_X1 U23381 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20433), .B1(
        n20531), .B2(n20432), .ZN(n20419) );
  OAI211_X1 U23382 ( .C1(n20535), .C2(n20436), .A(n20420), .B(n20419), .ZN(
        P1_U3130) );
  AOI22_X1 U23383 ( .A1(n20460), .A2(n20538), .B1(n20536), .B2(n20431), .ZN(
        n20422) );
  AOI22_X1 U23384 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20433), .B1(
        n20537), .B2(n20432), .ZN(n20421) );
  OAI211_X1 U23385 ( .C1(n20541), .C2(n20436), .A(n20422), .B(n20421), .ZN(
        P1_U3131) );
  AOI22_X1 U23386 ( .A1(n20460), .A2(n20544), .B1(n20542), .B2(n20431), .ZN(
        n20424) );
  AOI22_X1 U23387 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20433), .B1(
        n20543), .B2(n20432), .ZN(n20423) );
  OAI211_X1 U23388 ( .C1(n20547), .C2(n20436), .A(n20424), .B(n20423), .ZN(
        P1_U3132) );
  AOI22_X1 U23389 ( .A1(n20460), .A2(n20550), .B1(n20548), .B2(n20431), .ZN(
        n20426) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20433), .B1(
        n20549), .B2(n20432), .ZN(n20425) );
  OAI211_X1 U23391 ( .C1(n20553), .C2(n20436), .A(n20426), .B(n20425), .ZN(
        P1_U3133) );
  AOI22_X1 U23392 ( .A1(n20460), .A2(n20556), .B1(n20554), .B2(n20431), .ZN(
        n20428) );
  AOI22_X1 U23393 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20433), .B1(
        n20555), .B2(n20432), .ZN(n20427) );
  OAI211_X1 U23394 ( .C1(n20559), .C2(n20436), .A(n20428), .B(n20427), .ZN(
        P1_U3134) );
  AOI22_X1 U23395 ( .A1(n20460), .A2(n20562), .B1(n20560), .B2(n20431), .ZN(
        n20430) );
  AOI22_X1 U23396 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20433), .B1(
        n20561), .B2(n20432), .ZN(n20429) );
  OAI211_X1 U23397 ( .C1(n20565), .C2(n20436), .A(n20430), .B(n20429), .ZN(
        P1_U3135) );
  AOI22_X1 U23398 ( .A1(n20460), .A2(n20570), .B1(n20567), .B2(n20431), .ZN(
        n20435) );
  AOI22_X1 U23399 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20433), .B1(
        n20569), .B2(n20432), .ZN(n20434) );
  OAI211_X1 U23400 ( .C1(n20576), .C2(n20436), .A(n20435), .B(n20434), .ZN(
        P1_U3136) );
  NOR2_X1 U23401 ( .A1(n20665), .A2(n20439), .ZN(n20458) );
  INV_X1 U23402 ( .A(n20458), .ZN(n20440) );
  INV_X1 U23403 ( .A(n20438), .ZN(n20471) );
  NAND2_X1 U23404 ( .A1(n20471), .A2(n20657), .ZN(n20518) );
  OAI222_X1 U23405 ( .A1(n20440), .A2(n20515), .B1(n20581), .B2(n20439), .C1(
        n20050), .C2(n20518), .ZN(n20459) );
  AOI22_X1 U23406 ( .A1(n20520), .A2(n20459), .B1(n20519), .B2(n20458), .ZN(
        n20445) );
  NAND2_X1 U23407 ( .A1(n20465), .A2(n20657), .ZN(n20522) );
  NOR2_X1 U23408 ( .A1(n20522), .A2(n20441), .ZN(n20443) );
  OAI21_X1 U23409 ( .B1(n20443), .B2(n20442), .A(n20523), .ZN(n20461) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20461), .B1(
        n20460), .B2(n20477), .ZN(n20444) );
  OAI211_X1 U23411 ( .C1(n20480), .C2(n20476), .A(n20445), .B(n20444), .ZN(
        P1_U3137) );
  AOI22_X1 U23412 ( .A1(n20531), .A2(n20459), .B1(n20530), .B2(n20458), .ZN(
        n20447) );
  AOI22_X1 U23413 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20461), .B1(
        n20460), .B2(n20481), .ZN(n20446) );
  OAI211_X1 U23414 ( .C1(n20484), .C2(n20476), .A(n20447), .B(n20446), .ZN(
        P1_U3138) );
  AOI22_X1 U23415 ( .A1(n20537), .A2(n20459), .B1(n20536), .B2(n20458), .ZN(
        n20449) );
  AOI22_X1 U23416 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20461), .B1(
        n20460), .B2(n20485), .ZN(n20448) );
  OAI211_X1 U23417 ( .C1(n20488), .C2(n20476), .A(n20449), .B(n20448), .ZN(
        P1_U3139) );
  AOI22_X1 U23418 ( .A1(n20543), .A2(n20459), .B1(n20542), .B2(n20458), .ZN(
        n20451) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20461), .B1(
        n20460), .B2(n20489), .ZN(n20450) );
  OAI211_X1 U23420 ( .C1(n20492), .C2(n20476), .A(n20451), .B(n20450), .ZN(
        P1_U3140) );
  AOI22_X1 U23421 ( .A1(n20549), .A2(n20459), .B1(n20548), .B2(n20458), .ZN(
        n20453) );
  AOI22_X1 U23422 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20461), .B1(
        n20460), .B2(n20493), .ZN(n20452) );
  OAI211_X1 U23423 ( .C1(n20496), .C2(n20476), .A(n20453), .B(n20452), .ZN(
        P1_U3141) );
  AOI22_X1 U23424 ( .A1(n20555), .A2(n20459), .B1(n20554), .B2(n20458), .ZN(
        n20455) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20461), .B1(
        n20460), .B2(n20497), .ZN(n20454) );
  OAI211_X1 U23426 ( .C1(n20500), .C2(n20476), .A(n20455), .B(n20454), .ZN(
        P1_U3142) );
  AOI22_X1 U23427 ( .A1(n20561), .A2(n20459), .B1(n20560), .B2(n20458), .ZN(
        n20457) );
  AOI22_X1 U23428 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20461), .B1(
        n20460), .B2(n20501), .ZN(n20456) );
  OAI211_X1 U23429 ( .C1(n20504), .C2(n20476), .A(n20457), .B(n20456), .ZN(
        P1_U3143) );
  AOI22_X1 U23430 ( .A1(n20569), .A2(n20459), .B1(n20567), .B2(n20458), .ZN(
        n20463) );
  AOI22_X1 U23431 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20461), .B1(
        n20460), .B2(n20507), .ZN(n20462) );
  OAI211_X1 U23432 ( .C1(n20512), .C2(n20476), .A(n20463), .B(n20462), .ZN(
        P1_U3144) );
  OAI22_X1 U23433 ( .A1(n20518), .A2(n13459), .B1(n20467), .B2(n20466), .ZN(
        n20506) );
  NOR2_X1 U23434 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20516), .ZN(
        n20505) );
  AOI22_X1 U23435 ( .A1(n20520), .A2(n20506), .B1(n20519), .B2(n20505), .ZN(
        n20479) );
  AOI21_X1 U23436 ( .B1(n20476), .B2(n20575), .A(n20468), .ZN(n20469) );
  AOI21_X1 U23437 ( .B1(n20471), .B2(n20470), .A(n20469), .ZN(n20472) );
  NOR2_X1 U23438 ( .A1(n20472), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20475) );
  AOI22_X1 U23439 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20477), .ZN(n20478) );
  OAI211_X1 U23440 ( .C1(n20480), .C2(n20575), .A(n20479), .B(n20478), .ZN(
        P1_U3145) );
  AOI22_X1 U23441 ( .A1(n20531), .A2(n20506), .B1(n20530), .B2(n20505), .ZN(
        n20483) );
  AOI22_X1 U23442 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20481), .ZN(n20482) );
  OAI211_X1 U23443 ( .C1(n20484), .C2(n20575), .A(n20483), .B(n20482), .ZN(
        P1_U3146) );
  AOI22_X1 U23444 ( .A1(n20537), .A2(n20506), .B1(n20536), .B2(n20505), .ZN(
        n20487) );
  AOI22_X1 U23445 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20485), .ZN(n20486) );
  OAI211_X1 U23446 ( .C1(n20488), .C2(n20575), .A(n20487), .B(n20486), .ZN(
        P1_U3147) );
  AOI22_X1 U23447 ( .A1(n20543), .A2(n20506), .B1(n20542), .B2(n20505), .ZN(
        n20491) );
  AOI22_X1 U23448 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20489), .ZN(n20490) );
  OAI211_X1 U23449 ( .C1(n20492), .C2(n20575), .A(n20491), .B(n20490), .ZN(
        P1_U3148) );
  AOI22_X1 U23450 ( .A1(n20549), .A2(n20506), .B1(n20548), .B2(n20505), .ZN(
        n20495) );
  AOI22_X1 U23451 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20493), .ZN(n20494) );
  OAI211_X1 U23452 ( .C1(n20496), .C2(n20575), .A(n20495), .B(n20494), .ZN(
        P1_U3149) );
  AOI22_X1 U23453 ( .A1(n20555), .A2(n20506), .B1(n20554), .B2(n20505), .ZN(
        n20499) );
  AOI22_X1 U23454 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20497), .ZN(n20498) );
  OAI211_X1 U23455 ( .C1(n20500), .C2(n20575), .A(n20499), .B(n20498), .ZN(
        P1_U3150) );
  AOI22_X1 U23456 ( .A1(n20561), .A2(n20506), .B1(n20560), .B2(n20505), .ZN(
        n20503) );
  AOI22_X1 U23457 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20501), .ZN(n20502) );
  OAI211_X1 U23458 ( .C1(n20504), .C2(n20575), .A(n20503), .B(n20502), .ZN(
        P1_U3151) );
  AOI22_X1 U23459 ( .A1(n20569), .A2(n20506), .B1(n20567), .B2(n20505), .ZN(
        n20511) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20509), .B1(
        n20508), .B2(n20507), .ZN(n20510) );
  OAI211_X1 U23461 ( .C1(n20512), .C2(n20575), .A(n20511), .B(n20510), .ZN(
        P1_U3152) );
  INV_X1 U23462 ( .A(n20513), .ZN(n20517) );
  OAI222_X1 U23463 ( .A1(n20518), .A2(n20517), .B1(n20581), .B2(n20516), .C1(
        n20515), .C2(n20514), .ZN(n20568) );
  AOI22_X1 U23464 ( .A1(n20520), .A2(n20568), .B1(n20519), .B2(n20566), .ZN(
        n20528) );
  NOR2_X1 U23465 ( .A1(n20522), .A2(n20521), .ZN(n20524) );
  OAI21_X1 U23466 ( .B1(n20525), .B2(n20524), .A(n20523), .ZN(n20572) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20572), .B1(
        n20571), .B2(n20526), .ZN(n20527) );
  OAI211_X1 U23468 ( .C1(n20529), .C2(n20575), .A(n20528), .B(n20527), .ZN(
        P1_U3153) );
  AOI22_X1 U23469 ( .A1(n20531), .A2(n20568), .B1(n20530), .B2(n20566), .ZN(
        n20534) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20572), .B1(
        n20571), .B2(n20532), .ZN(n20533) );
  OAI211_X1 U23471 ( .C1(n20535), .C2(n20575), .A(n20534), .B(n20533), .ZN(
        P1_U3154) );
  AOI22_X1 U23472 ( .A1(n20537), .A2(n20568), .B1(n20536), .B2(n20566), .ZN(
        n20540) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20572), .B1(
        n20571), .B2(n20538), .ZN(n20539) );
  OAI211_X1 U23474 ( .C1(n20541), .C2(n20575), .A(n20540), .B(n20539), .ZN(
        P1_U3155) );
  AOI22_X1 U23475 ( .A1(n20543), .A2(n20568), .B1(n20542), .B2(n20566), .ZN(
        n20546) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20572), .B1(
        n20571), .B2(n20544), .ZN(n20545) );
  OAI211_X1 U23477 ( .C1(n20547), .C2(n20575), .A(n20546), .B(n20545), .ZN(
        P1_U3156) );
  AOI22_X1 U23478 ( .A1(n20549), .A2(n20568), .B1(n20548), .B2(n20566), .ZN(
        n20552) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20572), .B1(
        n20571), .B2(n20550), .ZN(n20551) );
  OAI211_X1 U23480 ( .C1(n20553), .C2(n20575), .A(n20552), .B(n20551), .ZN(
        P1_U3157) );
  AOI22_X1 U23481 ( .A1(n20555), .A2(n20568), .B1(n20554), .B2(n20566), .ZN(
        n20558) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20572), .B1(
        n20571), .B2(n20556), .ZN(n20557) );
  OAI211_X1 U23483 ( .C1(n20559), .C2(n20575), .A(n20558), .B(n20557), .ZN(
        P1_U3158) );
  AOI22_X1 U23484 ( .A1(n20561), .A2(n20568), .B1(n20560), .B2(n20566), .ZN(
        n20564) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20572), .B1(
        n20571), .B2(n20562), .ZN(n20563) );
  OAI211_X1 U23486 ( .C1(n20565), .C2(n20575), .A(n20564), .B(n20563), .ZN(
        P1_U3159) );
  AOI22_X1 U23487 ( .A1(n20569), .A2(n20568), .B1(n20567), .B2(n20566), .ZN(
        n20574) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20572), .B1(
        n20571), .B2(n20570), .ZN(n20573) );
  OAI211_X1 U23489 ( .C1(n20576), .C2(n20575), .A(n20574), .B(n20573), .ZN(
        P1_U3160) );
  NOR2_X1 U23490 ( .A1(n20578), .A2(n20577), .ZN(n20582) );
  INV_X1 U23491 ( .A(n20579), .ZN(n20580) );
  OAI21_X1 U23492 ( .B1(n20582), .B2(n20581), .A(n20580), .ZN(P1_U3163) );
  AND2_X1 U23493 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20583), .ZN(
        P1_U3164) );
  AND2_X1 U23494 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20583), .ZN(
        P1_U3165) );
  AND2_X1 U23495 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20583), .ZN(
        P1_U3166) );
  AND2_X1 U23496 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20583), .ZN(
        P1_U3167) );
  AND2_X1 U23497 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20583), .ZN(
        P1_U3168) );
  AND2_X1 U23498 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20583), .ZN(
        P1_U3169) );
  AND2_X1 U23499 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20583), .ZN(
        P1_U3170) );
  AND2_X1 U23500 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20583), .ZN(
        P1_U3171) );
  AND2_X1 U23501 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20583), .ZN(
        P1_U3172) );
  AND2_X1 U23502 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20583), .ZN(
        P1_U3173) );
  AND2_X1 U23503 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20583), .ZN(
        P1_U3174) );
  INV_X1 U23504 ( .A(P1_DATAWIDTH_REG_20__SCAN_IN), .ZN(n20697) );
  NOR2_X1 U23505 ( .A1(n20648), .A2(n20697), .ZN(P1_U3175) );
  AND2_X1 U23506 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20583), .ZN(
        P1_U3176) );
  AND2_X1 U23507 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20583), .ZN(
        P1_U3177) );
  AND2_X1 U23508 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20583), .ZN(
        P1_U3178) );
  AND2_X1 U23509 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20583), .ZN(
        P1_U3179) );
  INV_X1 U23510 ( .A(P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20732) );
  NOR2_X1 U23511 ( .A1(n20648), .A2(n20732), .ZN(P1_U3180) );
  AND2_X1 U23512 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20583), .ZN(
        P1_U3181) );
  AND2_X1 U23513 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20583), .ZN(
        P1_U3182) );
  AND2_X1 U23514 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20583), .ZN(
        P1_U3183) );
  AND2_X1 U23515 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20583), .ZN(
        P1_U3184) );
  AND2_X1 U23516 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20583), .ZN(
        P1_U3185) );
  AND2_X1 U23517 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20583), .ZN(P1_U3186) );
  AND2_X1 U23518 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20583), .ZN(P1_U3187) );
  AND2_X1 U23519 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20583), .ZN(P1_U3188) );
  AND2_X1 U23520 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20583), .ZN(P1_U3189) );
  AND2_X1 U23521 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20583), .ZN(P1_U3190) );
  AND2_X1 U23522 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20583), .ZN(P1_U3191) );
  AND2_X1 U23523 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20583), .ZN(P1_U3192) );
  AND2_X1 U23524 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20583), .ZN(P1_U3193) );
  AOI21_X1 U23525 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20585), .A(n20584), 
        .ZN(n20597) );
  OAI22_X1 U23526 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20592), .B1(n20599), 
        .B2(n20595), .ZN(n20586) );
  NOR3_X1 U23527 ( .A1(n20587), .A2(n20685), .A3(n20586), .ZN(n20588) );
  OAI22_X1 U23528 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20597), .B1(n20598), 
        .B2(n20588), .ZN(P1_U3194) );
  INV_X1 U23529 ( .A(n20589), .ZN(n20590) );
  AOI221_X1 U23530 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20592), .C1(n20591), 
        .C2(n20592), .A(n20590), .ZN(n20596) );
  OAI211_X1 U23531 ( .C1(NA), .C2(n20677), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n20599), .ZN(n20593) );
  OAI211_X1 U23532 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20685), .A(
        P1_STATE_REG_0__SCAN_IN), .B(n20593), .ZN(n20594) );
  OAI22_X1 U23533 ( .A1(n20597), .A2(n20596), .B1(n20595), .B2(n20594), .ZN(
        P1_U3196) );
  OR2_X1 U23534 ( .A1(n20599), .A2(n20673), .ZN(n20627) );
  NAND2_X1 U23535 ( .A1(n20599), .A2(n20598), .ZN(n20630) );
  INV_X1 U23536 ( .A(n20630), .ZN(n20638) );
  AOI22_X1 U23537 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n20673), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20638), .ZN(n20600) );
  OAI21_X1 U23538 ( .B1(n13624), .B2(n20627), .A(n20600), .ZN(P1_U3197) );
  AOI22_X1 U23539 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20673), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20639), .ZN(n20601) );
  OAI21_X1 U23540 ( .B1(n20602), .B2(n20630), .A(n20601), .ZN(P1_U3198) );
  INV_X1 U23541 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20695) );
  INV_X1 U23542 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20603) );
  OAI222_X1 U23543 ( .A1(n20627), .A2(n20602), .B1(n20695), .B2(n20598), .C1(
        n20603), .C2(n20630), .ZN(P1_U3199) );
  OAI222_X1 U23544 ( .A1(n20630), .A2(n20605), .B1(n20604), .B2(n20598), .C1(
        n20603), .C2(n20627), .ZN(P1_U3200) );
  AOI222_X1 U23545 ( .A1(n20639), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20687), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20638), .ZN(n20606) );
  INV_X1 U23546 ( .A(n20606), .ZN(P1_U3201) );
  AOI222_X1 U23547 ( .A1(n20639), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20687), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20638), .ZN(n20607) );
  INV_X1 U23548 ( .A(n20607), .ZN(P1_U3202) );
  AOI222_X1 U23549 ( .A1(n20639), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20687), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20638), .ZN(n20608) );
  INV_X1 U23550 ( .A(n20608), .ZN(P1_U3203) );
  AOI22_X1 U23551 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n20673), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20638), .ZN(n20609) );
  OAI21_X1 U23552 ( .B1(n13859), .B2(n20627), .A(n20609), .ZN(P1_U3204) );
  AOI22_X1 U23553 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n20673), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20639), .ZN(n20610) );
  OAI21_X1 U23554 ( .B1(n14529), .B2(n20630), .A(n20610), .ZN(P1_U3205) );
  AOI222_X1 U23555 ( .A1(n20638), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20687), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20639), .ZN(n20611) );
  INV_X1 U23556 ( .A(n20611), .ZN(P1_U3206) );
  AOI22_X1 U23557 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20673), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20638), .ZN(n20612) );
  OAI21_X1 U23558 ( .B1(n20613), .B2(n20627), .A(n20612), .ZN(P1_U3207) );
  AOI22_X1 U23559 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20673), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20639), .ZN(n20614) );
  OAI21_X1 U23560 ( .B1(n20615), .B2(n20630), .A(n20614), .ZN(P1_U3208) );
  AOI222_X1 U23561 ( .A1(n20639), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20687), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20638), .ZN(n20616) );
  INV_X1 U23562 ( .A(n20616), .ZN(P1_U3209) );
  AOI222_X1 U23563 ( .A1(n20638), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20687), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20639), .ZN(n20617) );
  INV_X1 U23564 ( .A(n20617), .ZN(P1_U3210) );
  AOI222_X1 U23565 ( .A1(n20639), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20687), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20638), .ZN(n20618) );
  INV_X1 U23566 ( .A(n20618), .ZN(P1_U3211) );
  INV_X1 U23567 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n20741) );
  OAI222_X1 U23568 ( .A1(n20627), .A2(n20620), .B1(n20741), .B2(n20598), .C1(
        n20619), .C2(n20630), .ZN(P1_U3212) );
  AOI222_X1 U23569 ( .A1(n20638), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20687), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20639), .ZN(n20621) );
  INV_X1 U23570 ( .A(n20621), .ZN(P1_U3213) );
  AOI222_X1 U23571 ( .A1(n20639), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20687), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20638), .ZN(n20622) );
  INV_X1 U23572 ( .A(n20622), .ZN(P1_U3214) );
  AOI222_X1 U23573 ( .A1(n20638), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20687), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20639), .ZN(n20623) );
  INV_X1 U23574 ( .A(n20623), .ZN(P1_U3215) );
  AOI222_X1 U23575 ( .A1(n20639), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20687), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20638), .ZN(n20624) );
  INV_X1 U23576 ( .A(n20624), .ZN(P1_U3216) );
  AOI222_X1 U23577 ( .A1(n20638), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20687), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20639), .ZN(n20625) );
  INV_X1 U23578 ( .A(n20625), .ZN(P1_U3217) );
  AOI22_X1 U23579 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20673), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20638), .ZN(n20626) );
  OAI21_X1 U23580 ( .B1(n20628), .B2(n20627), .A(n20626), .ZN(P1_U3218) );
  AOI22_X1 U23581 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20673), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20639), .ZN(n20629) );
  OAI21_X1 U23582 ( .B1(n20631), .B2(n20630), .A(n20629), .ZN(P1_U3219) );
  AOI222_X1 U23583 ( .A1(n20639), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20687), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20638), .ZN(n20632) );
  INV_X1 U23584 ( .A(n20632), .ZN(P1_U3220) );
  AOI222_X1 U23585 ( .A1(n20638), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20687), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20639), .ZN(n20633) );
  INV_X1 U23586 ( .A(n20633), .ZN(P1_U3221) );
  AOI222_X1 U23587 ( .A1(n20639), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20673), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20638), .ZN(n20634) );
  INV_X1 U23588 ( .A(n20634), .ZN(P1_U3222) );
  AOI222_X1 U23589 ( .A1(n20638), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20687), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20639), .ZN(n20635) );
  INV_X1 U23590 ( .A(n20635), .ZN(P1_U3223) );
  AOI222_X1 U23591 ( .A1(n20639), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20687), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20638), .ZN(n20636) );
  INV_X1 U23592 ( .A(n20636), .ZN(P1_U3224) );
  AOI222_X1 U23593 ( .A1(n20639), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20687), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n20638), .ZN(n20637) );
  INV_X1 U23594 ( .A(n20637), .ZN(P1_U3225) );
  AOI222_X1 U23595 ( .A1(n20639), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20687), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20638), .ZN(n20640) );
  INV_X1 U23596 ( .A(n20640), .ZN(P1_U3226) );
  INV_X1 U23597 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20709) );
  AOI22_X1 U23598 ( .A1(n20598), .A2(n20641), .B1(n20709), .B2(n20673), .ZN(
        P1_U3458) );
  OAI22_X1 U23599 ( .A1(n20687), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20598), .ZN(n20642) );
  INV_X1 U23600 ( .A(n20642), .ZN(P1_U3459) );
  OAI22_X1 U23601 ( .A1(n20673), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20598), .ZN(n20643) );
  INV_X1 U23602 ( .A(n20643), .ZN(P1_U3460) );
  OAI22_X1 U23603 ( .A1(n20673), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20598), .ZN(n20644) );
  INV_X1 U23604 ( .A(n20644), .ZN(P1_U3461) );
  OAI21_X1 U23605 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20648), .A(n20646), 
        .ZN(n20645) );
  INV_X1 U23606 ( .A(n20645), .ZN(P1_U3464) );
  OAI21_X1 U23607 ( .B1(n20648), .B2(n20647), .A(n20646), .ZN(P1_U3465) );
  INV_X1 U23608 ( .A(n20649), .ZN(n20654) );
  INV_X1 U23609 ( .A(n20650), .ZN(n20653) );
  OAI22_X1 U23610 ( .A1(n20654), .A2(n20653), .B1(n20652), .B2(n20651), .ZN(
        n20656) );
  MUX2_X1 U23611 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20656), .S(
        n20655), .Z(P1_U3469) );
  AOI22_X1 U23612 ( .A1(n20660), .A2(n20659), .B1(n20658), .B2(n20657), .ZN(
        n20663) );
  NOR2_X1 U23613 ( .A1(n20664), .A2(n20661), .ZN(n20662) );
  AOI22_X1 U23614 ( .A1(n20665), .A2(n20664), .B1(n20663), .B2(n20662), .ZN(
        P1_U3478) );
  AOI21_X1 U23615 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20666) );
  AOI22_X1 U23616 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20666), .B2(n13624), .ZN(n20669) );
  INV_X1 U23617 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20668) );
  AOI22_X1 U23618 ( .A1(n20672), .A2(n20669), .B1(n20668), .B2(n20667), .ZN(
        P1_U3481) );
  INV_X1 U23619 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20671) );
  OAI21_X1 U23620 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20672), .ZN(n20670) );
  OAI21_X1 U23621 ( .B1(n20672), .B2(n20671), .A(n20670), .ZN(P1_U3482) );
  AOI22_X1 U23622 ( .A1(n20598), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20674), 
        .B2(n20673), .ZN(P1_U3483) );
  AOI211_X1 U23623 ( .C1(n20677), .C2(n19884), .A(n20676), .B(n20675), .ZN(
        n20679) );
  NAND2_X1 U23624 ( .A1(n20679), .A2(n20678), .ZN(n20686) );
  NOR2_X1 U23625 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20680), .ZN(n20684) );
  OAI211_X1 U23626 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n11295), .A(n20681), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20682) );
  NAND2_X1 U23627 ( .A1(n20686), .A2(n20682), .ZN(n20683) );
  OAI22_X1 U23628 ( .A1(n20686), .A2(n20685), .B1(n20684), .B2(n20683), .ZN(
        P1_U3485) );
  OAI22_X1 U23629 ( .A1(n20687), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n20598), .ZN(n20688) );
  INV_X1 U23630 ( .A(n20688), .ZN(P1_U3486) );
  INV_X1 U23631 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n20691) );
  AOI22_X1 U23632 ( .A1(n20691), .A2(keyinput43), .B1(keyinput17), .B2(n20690), 
        .ZN(n20689) );
  OAI221_X1 U23633 ( .B1(n20691), .B2(keyinput43), .C1(n20690), .C2(keyinput17), .A(n20689), .ZN(n20702) );
  AOI22_X1 U23634 ( .A1(n20846), .A2(keyinput29), .B1(n20693), .B2(keyinput12), 
        .ZN(n20692) );
  OAI221_X1 U23635 ( .B1(n20846), .B2(keyinput29), .C1(n20693), .C2(keyinput12), .A(n20692), .ZN(n20701) );
  AOI22_X1 U23636 ( .A1(n20695), .A2(keyinput28), .B1(n10389), .B2(keyinput62), 
        .ZN(n20694) );
  OAI221_X1 U23637 ( .B1(n20695), .B2(keyinput28), .C1(n10389), .C2(keyinput62), .A(n20694), .ZN(n20700) );
  AOI22_X1 U23638 ( .A1(n20698), .A2(keyinput37), .B1(keyinput36), .B2(n20697), 
        .ZN(n20696) );
  OAI221_X1 U23639 ( .B1(n20698), .B2(keyinput37), .C1(n20697), .C2(keyinput36), .A(n20696), .ZN(n20699) );
  NOR4_X1 U23640 ( .A1(n20702), .A2(n20701), .A3(n20700), .A4(n20699), .ZN(
        n20749) );
  AOI22_X1 U23641 ( .A1(n20847), .A2(keyinput21), .B1(n20848), .B2(keyinput59), 
        .ZN(n20703) );
  OAI221_X1 U23642 ( .B1(n20847), .B2(keyinput21), .C1(n20848), .C2(keyinput59), .A(n20703), .ZN(n20716) );
  AOI22_X1 U23643 ( .A1(n20706), .A2(keyinput4), .B1(keyinput54), .B2(n20705), 
        .ZN(n20704) );
  OAI221_X1 U23644 ( .B1(n20706), .B2(keyinput4), .C1(n20705), .C2(keyinput54), 
        .A(n20704), .ZN(n20715) );
  AOI22_X1 U23645 ( .A1(n20709), .A2(keyinput53), .B1(n20708), .B2(keyinput57), 
        .ZN(n20707) );
  OAI221_X1 U23646 ( .B1(n20709), .B2(keyinput53), .C1(n20708), .C2(keyinput57), .A(n20707), .ZN(n20714) );
  AOI22_X1 U23647 ( .A1(n20712), .A2(keyinput60), .B1(n20711), .B2(keyinput10), 
        .ZN(n20710) );
  OAI221_X1 U23648 ( .B1(n20712), .B2(keyinput60), .C1(n20711), .C2(keyinput10), .A(n20710), .ZN(n20713) );
  NOR4_X1 U23649 ( .A1(n20716), .A2(n20715), .A3(n20714), .A4(n20713), .ZN(
        n20748) );
  INV_X1 U23650 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n20718) );
  AOI22_X1 U23651 ( .A1(n20719), .A2(keyinput33), .B1(keyinput38), .B2(n20718), 
        .ZN(n20717) );
  OAI221_X1 U23652 ( .B1(n20719), .B2(keyinput33), .C1(n20718), .C2(keyinput38), .A(n20717), .ZN(n20730) );
  INV_X1 U23653 ( .A(P3_MORE_REG_SCAN_IN), .ZN(n20721) );
  AOI22_X1 U23654 ( .A1(n20721), .A2(keyinput20), .B1(n12714), .B2(keyinput44), 
        .ZN(n20720) );
  OAI221_X1 U23655 ( .B1(n20721), .B2(keyinput20), .C1(n12714), .C2(keyinput44), .A(n20720), .ZN(n20729) );
  AOI22_X1 U23656 ( .A1(n20723), .A2(keyinput30), .B1(n10551), .B2(keyinput31), 
        .ZN(n20722) );
  OAI221_X1 U23657 ( .B1(n20723), .B2(keyinput30), .C1(n10551), .C2(keyinput31), .A(n20722), .ZN(n20728) );
  INV_X1 U23658 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20726) );
  AOI22_X1 U23659 ( .A1(n20726), .A2(keyinput13), .B1(n20725), .B2(keyinput39), 
        .ZN(n20724) );
  OAI221_X1 U23660 ( .B1(n20726), .B2(keyinput13), .C1(n20725), .C2(keyinput39), .A(n20724), .ZN(n20727) );
  NOR4_X1 U23661 ( .A1(n20730), .A2(n20729), .A3(n20728), .A4(n20727), .ZN(
        n20747) );
  INV_X1 U23662 ( .A(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n20837) );
  AOI22_X1 U23663 ( .A1(n20732), .A2(keyinput63), .B1(n20837), .B2(keyinput58), 
        .ZN(n20731) );
  OAI221_X1 U23664 ( .B1(n20732), .B2(keyinput63), .C1(n20837), .C2(keyinput58), .A(n20731), .ZN(n20745) );
  AOI22_X1 U23665 ( .A1(n20735), .A2(keyinput14), .B1(n20734), .B2(keyinput35), 
        .ZN(n20733) );
  OAI221_X1 U23666 ( .B1(n20735), .B2(keyinput14), .C1(n20734), .C2(keyinput35), .A(n20733), .ZN(n20744) );
  INV_X1 U23667 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n20737) );
  AOI22_X1 U23668 ( .A1(n20738), .A2(keyinput2), .B1(keyinput48), .B2(n20737), 
        .ZN(n20736) );
  OAI221_X1 U23669 ( .B1(n20738), .B2(keyinput2), .C1(n20737), .C2(keyinput48), 
        .A(n20736), .ZN(n20743) );
  AOI22_X1 U23670 ( .A1(n20741), .A2(keyinput0), .B1(keyinput8), .B2(n20740), 
        .ZN(n20739) );
  OAI221_X1 U23671 ( .B1(n20741), .B2(keyinput0), .C1(n20740), .C2(keyinput8), 
        .A(n20739), .ZN(n20742) );
  NOR4_X1 U23672 ( .A1(n20745), .A2(n20744), .A3(n20743), .A4(n20742), .ZN(
        n20746) );
  NAND4_X1 U23673 ( .A1(n20749), .A2(n20748), .A3(n20747), .A4(n20746), .ZN(
        n20815) );
  AOI22_X1 U23674 ( .A1(n20752), .A2(keyinput25), .B1(n20751), .B2(keyinput55), 
        .ZN(n20750) );
  OAI221_X1 U23675 ( .B1(n20752), .B2(keyinput25), .C1(n20751), .C2(keyinput55), .A(n20750), .ZN(n20765) );
  INV_X1 U23676 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n20754) );
  AOI22_X1 U23677 ( .A1(n20755), .A2(keyinput56), .B1(keyinput19), .B2(n20754), 
        .ZN(n20753) );
  OAI221_X1 U23678 ( .B1(n20755), .B2(keyinput56), .C1(n20754), .C2(keyinput19), .A(n20753), .ZN(n20764) );
  INV_X1 U23679 ( .A(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n20757) );
  AOI22_X1 U23680 ( .A1(n20758), .A2(keyinput6), .B1(n20757), .B2(keyinput18), 
        .ZN(n20756) );
  OAI221_X1 U23681 ( .B1(n20758), .B2(keyinput6), .C1(n20757), .C2(keyinput18), 
        .A(n20756), .ZN(n20763) );
  XOR2_X1 U23682 ( .A(n20759), .B(keyinput41), .Z(n20761) );
  XNOR2_X1 U23683 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B(keyinput42), .ZN(
        n20760) );
  NAND2_X1 U23684 ( .A1(n20761), .A2(n20760), .ZN(n20762) );
  NOR4_X1 U23685 ( .A1(n20765), .A2(n20764), .A3(n20763), .A4(n20762), .ZN(
        n20813) );
  AOI22_X1 U23686 ( .A1(n20849), .A2(keyinput22), .B1(keyinput16), .B2(n20767), 
        .ZN(n20766) );
  OAI221_X1 U23687 ( .B1(n20849), .B2(keyinput22), .C1(n20767), .C2(keyinput16), .A(n20766), .ZN(n20780) );
  AOI22_X1 U23688 ( .A1(n20770), .A2(keyinput40), .B1(keyinput50), .B2(n20769), 
        .ZN(n20768) );
  OAI221_X1 U23689 ( .B1(n20770), .B2(keyinput40), .C1(n20769), .C2(keyinput50), .A(n20768), .ZN(n20779) );
  INV_X1 U23690 ( .A(P1_LWORD_REG_4__SCAN_IN), .ZN(n20773) );
  INV_X1 U23691 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n20772) );
  AOI22_X1 U23692 ( .A1(n20773), .A2(keyinput23), .B1(n20772), .B2(keyinput3), 
        .ZN(n20771) );
  OAI221_X1 U23693 ( .B1(n20773), .B2(keyinput23), .C1(n20772), .C2(keyinput3), 
        .A(n20771), .ZN(n20778) );
  AOI22_X1 U23694 ( .A1(n20776), .A2(keyinput11), .B1(keyinput34), .B2(n20775), 
        .ZN(n20774) );
  OAI221_X1 U23695 ( .B1(n20776), .B2(keyinput11), .C1(n20775), .C2(keyinput34), .A(n20774), .ZN(n20777) );
  NOR4_X1 U23696 ( .A1(n20780), .A2(n20779), .A3(n20778), .A4(n20777), .ZN(
        n20812) );
  INV_X1 U23697 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20782) );
  AOI22_X1 U23698 ( .A1(n20836), .A2(keyinput45), .B1(keyinput7), .B2(n20782), 
        .ZN(n20781) );
  OAI221_X1 U23699 ( .B1(n20836), .B2(keyinput45), .C1(n20782), .C2(keyinput7), 
        .A(n20781), .ZN(n20793) );
  AOI22_X1 U23700 ( .A1(n20838), .A2(keyinput51), .B1(keyinput9), .B2(n20784), 
        .ZN(n20783) );
  OAI221_X1 U23701 ( .B1(n20838), .B2(keyinput51), .C1(n20784), .C2(keyinput9), 
        .A(n20783), .ZN(n20792) );
  INV_X1 U23702 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n20786) );
  AOI22_X1 U23703 ( .A1(n20787), .A2(keyinput26), .B1(n20786), .B2(keyinput24), 
        .ZN(n20785) );
  OAI221_X1 U23704 ( .B1(n20787), .B2(keyinput26), .C1(n20786), .C2(keyinput24), .A(n20785), .ZN(n20791) );
  XOR2_X1 U23705 ( .A(n20835), .B(keyinput47), .Z(n20789) );
  XNOR2_X1 U23706 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B(keyinput5), .ZN(
        n20788) );
  NAND2_X1 U23707 ( .A1(n20789), .A2(n20788), .ZN(n20790) );
  NOR4_X1 U23708 ( .A1(n20793), .A2(n20792), .A3(n20791), .A4(n20790), .ZN(
        n20811) );
  AOI22_X1 U23709 ( .A1(n20796), .A2(keyinput46), .B1(keyinput52), .B2(n20795), 
        .ZN(n20794) );
  OAI221_X1 U23710 ( .B1(n20796), .B2(keyinput46), .C1(n20795), .C2(keyinput52), .A(n20794), .ZN(n20809) );
  INV_X1 U23711 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n20799) );
  AOI22_X1 U23712 ( .A1(n20799), .A2(keyinput32), .B1(keyinput61), .B2(n20798), 
        .ZN(n20797) );
  OAI221_X1 U23713 ( .B1(n20799), .B2(keyinput32), .C1(n20798), .C2(keyinput61), .A(n20797), .ZN(n20808) );
  INV_X1 U23714 ( .A(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n20802) );
  AOI22_X1 U23715 ( .A1(n20802), .A2(keyinput49), .B1(keyinput27), .B2(n20801), 
        .ZN(n20800) );
  OAI221_X1 U23716 ( .B1(n20802), .B2(keyinput49), .C1(n20801), .C2(keyinput27), .A(n20800), .ZN(n20807) );
  INV_X1 U23717 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n20804) );
  AOI22_X1 U23718 ( .A1(n20805), .A2(keyinput15), .B1(keyinput1), .B2(n20804), 
        .ZN(n20803) );
  OAI221_X1 U23719 ( .B1(n20805), .B2(keyinput15), .C1(n20804), .C2(keyinput1), 
        .A(n20803), .ZN(n20806) );
  NOR4_X1 U23720 ( .A1(n20809), .A2(n20808), .A3(n20807), .A4(n20806), .ZN(
        n20810) );
  NAND4_X1 U23721 ( .A1(n20813), .A2(n20812), .A3(n20811), .A4(n20810), .ZN(
        n20814) );
  NOR2_X1 U23722 ( .A1(n20815), .A2(n20814), .ZN(n20867) );
  AOI211_X1 U23723 ( .C1(n20819), .C2(n20818), .A(n20817), .B(n20816), .ZN(
        n20824) );
  AOI211_X1 U23724 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n20822), .A(n20821), .B(
        n20820), .ZN(n20823) );
  AOI211_X1 U23725 ( .C1(n20825), .C2(P3_REIP_REG_20__SCAN_IN), .A(n20824), 
        .B(n20823), .ZN(n20830) );
  OAI211_X1 U23726 ( .C1(P3_REIP_REG_20__SCAN_IN), .C2(n20828), .A(n20827), 
        .B(n20826), .ZN(n20829) );
  OAI211_X1 U23727 ( .C1(n20832), .C2(n20831), .A(n20830), .B(n20829), .ZN(
        n20833) );
  AOI21_X1 U23728 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n20834), .A(n20833), .ZN(
        n20865) );
  NOR4_X1 U23729 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .A3(P2_INSTQUEUE_REG_4__6__SCAN_IN), 
        .A4(P2_EBX_REG_1__SCAN_IN), .ZN(n20863) );
  NAND4_X1 U23730 ( .A1(n20838), .A2(n20837), .A3(n20836), .A4(n20835), .ZN(
        n20841) );
  NAND4_X1 U23731 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P1_ADDRESS_REG_15__SCAN_IN), .A3(P1_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P2_UWORD_REG_1__SCAN_IN), .ZN(n20840) );
  NAND4_X1 U23732 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20839) );
  NOR3_X1 U23733 ( .A1(n20841), .A2(n20840), .A3(n20839), .ZN(n20862) );
  NAND4_X1 U23734 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(P3_MORE_REG_SCAN_IN), .A4(P3_DATAO_REG_1__SCAN_IN), .ZN(n20845) );
  NAND4_X1 U23735 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_EBX_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_27__SCAN_IN), .A4(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n20844) );
  NAND4_X1 U23736 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_8__3__SCAN_IN), .A3(P1_INSTQUEUE_REG_2__3__SCAN_IN), 
        .A4(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n20843) );
  NAND4_X1 U23737 ( .A1(P1_EBX_REG_18__SCAN_IN), .A2(P1_EBX_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_19__SCAN_IN), .A4(P3_INSTADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n20842) );
  NOR4_X1 U23738 ( .A1(n20845), .A2(n20844), .A3(n20843), .A4(n20842), .ZN(
        n20861) );
  NAND3_X1 U23739 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_7__4__SCAN_IN), .A3(n20846), .ZN(n20859) );
  NOR4_X1 U23740 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_9__6__SCAN_IN), .A3(n20848), .A4(n20847), .ZN(n20852)
         );
  NOR4_X1 U23741 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_READREQUEST_REG_SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        n20849), .ZN(n20851) );
  NOR4_X1 U23742 ( .A1(P1_EBX_REG_23__SCAN_IN), .A2(P1_LWORD_REG_4__SCAN_IN), 
        .A3(P1_LWORD_REG_9__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n20850)
         );
  NAND3_X1 U23743 ( .A1(n20852), .A2(n20851), .A3(n20850), .ZN(n20858) );
  NOR4_X1 U23744 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_REIP_REG_4__SCAN_IN), .A3(P1_EBX_REG_3__SCAN_IN), .A4(
        BUF1_REG_15__SCAN_IN), .ZN(n20856) );
  NOR4_X1 U23745 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        BUF2_REG_1__SCAN_IN), .A3(P2_BYTEENABLE_REG_2__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20855) );
  NOR4_X1 U23746 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EAX_REG_16__SCAN_IN), 
        .A3(P3_EAX_REG_4__SCAN_IN), .A4(P2_DATAO_REG_18__SCAN_IN), .ZN(n20854)
         );
  NOR4_X1 U23747 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        BUF2_REG_12__SCAN_IN), .A3(P2_DATAO_REG_9__SCAN_IN), .A4(
        P2_DATAO_REG_29__SCAN_IN), .ZN(n20853) );
  NAND4_X1 U23748 ( .A1(n20856), .A2(n20855), .A3(n20854), .A4(n20853), .ZN(
        n20857) );
  NOR4_X1 U23749 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20859), .A3(
        n20858), .A4(n20857), .ZN(n20860) );
  NAND4_X1 U23750 ( .A1(n20863), .A2(n20862), .A3(n20861), .A4(n20860), .ZN(
        n20864) );
  XNOR2_X1 U23751 ( .A(n20865), .B(n20864), .ZN(n20866) );
  XNOR2_X1 U23752 ( .A(n20867), .B(n20866), .ZN(P3_U2651) );
  CLKBUF_X2 U13864 ( .A(n10888), .Z(n16911) );
  CLKBUF_X3 U12683 ( .A(n10877), .Z(n16952) );
  NAND2_X1 U14415 ( .A1(n11305), .A2(n11304), .ZN(n11371) );
  AOI21_X1 U14460 ( .B1(n11934), .B2(n11398), .A(n11357), .ZN(n11391) );
  NOR2_X1 U14628 ( .A1(n13793), .A2(n13796), .ZN(n13794) );
  CLKBUF_X2 U11038 ( .A(n11310), .Z(n9666) );
  CLKBUF_X1 U11057 ( .A(n11458), .Z(n11319) );
  CLKBUF_X1 U11063 ( .A(n16908), .Z(n9587) );
  INV_X1 U11090 ( .A(n12515), .ZN(n12509) );
  NAND2_X1 U11132 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18604), .ZN(
        n10808) );
  CLKBUF_X1 U11146 ( .A(n10888), .Z(n16844) );
  NOR2_X2 U11148 ( .A1(n10808), .A2(n9791), .ZN(n10890) );
  CLKBUF_X1 U11363 ( .A(n18575), .Z(n18568) );
  CLKBUF_X1 U11424 ( .A(n16299), .Z(n16307) );
endmodule

