

module b15_C_gen_AntiSAT_k_128_1 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, 
        U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, 
        U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, 
        U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, 
        U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, 
        U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, 
        U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, 
        U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, 
        U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, 
        U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, 
        U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, 
        U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, 
        U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, 
        U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, 
        U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, 
        U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, 
        U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, 
        U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, 
        U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, 
        U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, 
        U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, 
        U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, 
        U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, 
        U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, 
        U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, 
        U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, 
        U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, 
        U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, 
        U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, 
        U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, 
        U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, 
        U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, 
        U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, 
        U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, 
        U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, 
        U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, 
        U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, 
        U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, 
        U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, 
        U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, 
        U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, 
        U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, 
        U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, 
        U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, 
        U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, 
        U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788;

  OAI21_X1 U3434 ( .B1(n5357), .B2(n5356), .A(n5355), .ZN(n5361) );
  NAND2_X1 U3435 ( .A1(n5693), .A2(n5692), .ZN(n5695) );
  INV_X2 U3436 ( .A(n3903), .ZN(n3904) );
  XNOR2_X1 U3437 ( .A(n3416), .B(n3415), .ZN(n4481) );
  XNOR2_X1 U3438 ( .A(n3066), .B(n3414), .ZN(n3416) );
  CLKBUF_X1 U3439 ( .A(n4183), .Z(n3015) );
  CLKBUF_X2 U3440 ( .A(n3185), .Z(n4145) );
  AND4_X1 U3441 ( .A1(n3223), .A2(n3222), .A3(n3221), .A4(n3220), .ZN(n4511)
         );
  AND2_X1 U3442 ( .A1(n4393), .A2(n3095), .ZN(n3245) );
  AND2_X1 U3443 ( .A1(n4392), .A2(n4393), .ZN(n3395) );
  AND2_X1 U3444 ( .A1(n4340), .A2(n4422), .ZN(n3368) );
  AND3_X1 U34450 ( .A1(n3284), .A2(n3295), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3877) );
  AND2_X1 U34460 ( .A1(n4339), .A2(n4422), .ZN(n3389) );
  NOR2_X1 U34470 ( .A1(n3159), .A2(n3158), .ZN(n3006) );
  NAND2_X1 U34480 ( .A1(n3019), .A2(n5272), .ZN(n5416) );
  NAND4_X2 U3449 ( .A1(n3280), .A2(n3279), .A3(n3278), .A4(n3277), .ZN(n3295)
         );
  INV_X1 U3450 ( .A(n6071), .ZN(n6047) );
  OR2_X1 U34510 ( .A1(n5695), .A2(n4276), .ZN(n2986) );
  AOI21_X2 U34520 ( .B1(n3283), .B2(n4511), .A(n4246), .ZN(n3258) );
  AND2_X4 U34530 ( .A1(n4371), .A2(n3295), .ZN(n4989) );
  OAI22_X2 U3454 ( .A1(n5579), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5587), .B2(n5572), .ZN(n5573) );
  NAND2_X1 U34550 ( .A1(n3502), .A2(n3501), .ZN(n4448) );
  NAND2_X1 U34560 ( .A1(n3439), .A2(n4382), .ZN(n4384) );
  CLKBUF_X1 U3457 ( .A(n4477), .Z(n4478) );
  AND2_X1 U3458 ( .A1(n5186), .A2(n5185), .ZN(n3019) );
  CLKBUF_X1 U34590 ( .A(n3323), .Z(n3000) );
  CLKBUF_X1 U34600 ( .A(n3417), .Z(n4207) );
  BUF_X2 U34610 ( .A(n3244), .Z(n5338) );
  NAND4_X2 U34620 ( .A1(n3243), .A2(n3242), .A3(n3241), .A4(n3240), .ZN(n4371)
         );
  CLKBUF_X2 U34630 ( .A(n3368), .Z(n3790) );
  CLKBUF_X2 U34640 ( .A(n3395), .Z(n3369) );
  CLKBUF_X2 U34650 ( .A(n3592), .Z(n4188) );
  CLKBUF_X2 U3466 ( .A(n3451), .Z(n3337) );
  CLKBUF_X2 U3467 ( .A(n3250), .Z(n4151) );
  BUF_X2 U34680 ( .A(n3367), .Z(n3354) );
  BUF_X2 U34690 ( .A(n3245), .Z(n3785) );
  BUF_X2 U34700 ( .A(n4182), .Z(n4146) );
  AOI22_X1 U34710 ( .A1(n5541), .A2(n5550), .B1(
        INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5540), .ZN(n5542) );
  AND2_X1 U34720 ( .A1(n4227), .A2(n4226), .ZN(n2988) );
  CLKBUF_X1 U34730 ( .A(n2992), .Z(n5578) );
  NAND2_X1 U34740 ( .A1(n4273), .A2(n4272), .ZN(n5543) );
  AND2_X1 U3475 ( .A1(n5555), .A2(n5554), .ZN(n5879) );
  OR2_X1 U3476 ( .A1(n4271), .A2(n4270), .ZN(n4272) );
  AOI21_X1 U3477 ( .B1(n3832), .B2(n3021), .A(n4132), .ZN(n5565) );
  AND2_X1 U3478 ( .A1(n5462), .A2(n5477), .ZN(n5905) );
  CLKBUF_X1 U3479 ( .A(n5439), .Z(n5440) );
  NOR2_X1 U3481 ( .A1(n3022), .A2(n3057), .ZN(n3056) );
  CLKBUF_X1 U3482 ( .A(n4452), .Z(n4914) );
  INV_X2 U3483 ( .A(n5571), .ZN(n5618) );
  INV_X4 U3484 ( .A(n5571), .ZN(n5606) );
  NAND2_X1 U3485 ( .A1(n4081), .A2(n4083), .ZN(n4090) );
  NAND2_X1 U3486 ( .A1(n3545), .A2(n3544), .ZN(n4081) );
  AND2_X1 U3487 ( .A1(n3542), .A2(n3519), .ZN(n4053) );
  AOI21_X1 U3488 ( .B1(n4014), .B2(n3674), .A(n3500), .ZN(n4565) );
  AND2_X1 U3489 ( .A1(n3518), .A2(n3491), .ZN(n4014) );
  AND2_X1 U3490 ( .A1(n5466), .A2(n5465), .ZN(n5457) );
  XNOR2_X1 U3491 ( .A(n3351), .B(n3350), .ZN(n3412) );
  NAND2_X1 U3492 ( .A1(n3041), .A2(n3027), .ZN(n5496) );
  NOR2_X1 U3493 ( .A1(n6129), .A2(n6097), .ZN(n6128) );
  INV_X1 U3494 ( .A(n5416), .ZN(n3041) );
  AND2_X1 U3495 ( .A1(n4306), .A2(n4304), .ZN(n4309) );
  AND2_X1 U3496 ( .A1(n3001), .A2(n3002), .ZN(n3385) );
  NAND2_X1 U3497 ( .A1(n3292), .A2(n3291), .ZN(n3325) );
  OR2_X1 U3498 ( .A1(n4995), .A2(n4994), .ZN(n4997) );
  AND4_X1 U3499 ( .A1(n3321), .A2(n3320), .A3(n4529), .A4(n3319), .ZN(n3322)
         );
  AND2_X1 U3500 ( .A1(n3281), .A2(n4531), .ZN(n3321) );
  NOR2_X1 U3501 ( .A1(n4240), .A2(n4235), .ZN(n4110) );
  NAND2_X1 U3502 ( .A1(n3286), .A2(n3285), .ZN(n4240) );
  INV_X4 U3503 ( .A(n3904), .ZN(n4296) );
  NAND2_X1 U3504 ( .A1(n3282), .A2(n3296), .ZN(n3283) );
  INV_X1 U3505 ( .A(n3244), .ZN(n3282) );
  INV_X1 U3506 ( .A(n4019), .ZN(n4586) );
  OR2_X1 U3507 ( .A1(n3295), .A2(n4371), .ZN(n3298) );
  NAND2_X1 U3508 ( .A1(n3192), .A2(n3006), .ZN(n3202) );
  OR2_X1 U3509 ( .A1(n3380), .A2(n3379), .ZN(n4085) );
  NAND2_X2 U3510 ( .A1(n2996), .A2(n2997), .ZN(n3192) );
  NAND4_X2 U3511 ( .A1(n3180), .A2(n3179), .A3(n3178), .A4(n3177), .ZN(n3284)
         );
  OR2_X1 U3512 ( .A1(n3159), .A2(n3158), .ZN(n3296) );
  AND4_X1 U3513 ( .A1(n3207), .A2(n3206), .A3(n3205), .A4(n3204), .ZN(n3223)
         );
  AND3_X1 U3514 ( .A1(n3160), .A2(n3163), .A3(n3010), .ZN(n3180) );
  AND4_X1 U3515 ( .A1(n3149), .A2(n3146), .A3(n3147), .A4(n3148), .ZN(n2997)
         );
  AND4_X1 U3516 ( .A1(n3263), .A2(n3262), .A3(n3261), .A4(n3260), .ZN(n3280)
         );
  AND4_X1 U3517 ( .A1(n3231), .A2(n3230), .A3(n3229), .A4(n3228), .ZN(n3242)
         );
  AND4_X1 U3518 ( .A1(n3267), .A2(n3266), .A3(n3265), .A4(n3264), .ZN(n3279)
         );
  AND4_X1 U3519 ( .A1(n3235), .A2(n3234), .A3(n3233), .A4(n3232), .ZN(n3241)
         );
  AND4_X1 U3520 ( .A1(n3276), .A2(n3275), .A3(n3274), .A4(n3273), .ZN(n3277)
         );
  AND4_X1 U3521 ( .A1(n3271), .A2(n3270), .A3(n3269), .A4(n3268), .ZN(n3278)
         );
  AND4_X1 U3522 ( .A1(n3239), .A2(n3238), .A3(n3237), .A4(n3236), .ZN(n3240)
         );
  AND4_X1 U3523 ( .A1(n3227), .A2(n3226), .A3(n3225), .A4(n3224), .ZN(n3243)
         );
  AND4_X1 U3524 ( .A1(n3219), .A2(n3218), .A3(n3217), .A4(n3216), .ZN(n3220)
         );
  AND4_X1 U3525 ( .A1(n3171), .A2(n3170), .A3(n3169), .A4(n3168), .ZN(n3178)
         );
  AND4_X1 U3526 ( .A1(n3215), .A2(n3214), .A3(n3213), .A4(n3212), .ZN(n3221)
         );
  AND4_X1 U3527 ( .A1(n3211), .A2(n3210), .A3(n3209), .A4(n3208), .ZN(n3222)
         );
  AND2_X1 U3528 ( .A1(n3161), .A2(n3162), .ZN(n3010) );
  AND4_X1 U3529 ( .A1(n3167), .A2(n3166), .A3(n3165), .A4(n3164), .ZN(n3179)
         );
  AND4_X1 U3530 ( .A1(n3176), .A2(n3175), .A3(n3174), .A4(n3173), .ZN(n3177)
         );
  CLKBUF_X2 U3531 ( .A(n3389), .Z(n3016) );
  INV_X2 U3532 ( .A(n4395), .ZN(n3185) );
  AND2_X4 U3533 ( .A1(n4393), .A2(n4339), .ZN(n4183) );
  INV_X2 U3534 ( .A(n6786), .ZN(n6598) );
  AND2_X2 U3535 ( .A1(n4393), .A2(n4340), .ZN(n3374) );
  AND2_X2 U3536 ( .A1(n3094), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4393)
         );
  NOR2_X2 U3537 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3089) );
  NOR2_X2 U3538 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3095) );
  AND2_X2 U3539 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4392) );
  NAND2_X1 U3540 ( .A1(n5120), .A2(n5184), .ZN(n2987) );
  INV_X1 U3541 ( .A(n5499), .ZN(n2989) );
  NAND2_X1 U3542 ( .A1(n5120), .A2(n5184), .ZN(n5183) );
  NAND2_X1 U3543 ( .A1(n2991), .A2(n3047), .ZN(n2990) );
  INV_X1 U3544 ( .A(n3049), .ZN(n2991) );
  NOR2_X2 U3545 ( .A1(n5599), .A2(n5600), .ZN(n2992) );
  OR2_X2 U3546 ( .A1(n2992), .A2(n2993), .ZN(n5593) );
  OR2_X1 U3547 ( .A1(n2994), .A2(n3080), .ZN(n2993) );
  INV_X1 U3548 ( .A(n5594), .ZN(n2994) );
  NAND2_X1 U3549 ( .A1(n4092), .A2(n4091), .ZN(n5241) );
  OR2_X1 U3550 ( .A1(n3385), .A2(n3384), .ZN(n3386) );
  NAND2_X1 U3551 ( .A1(n4062), .A2(n4061), .ZN(n2995) );
  NAND2_X1 U3552 ( .A1(n4062), .A2(n4061), .ZN(n4691) );
  AOI21_X1 U3553 ( .B1(n3297), .B2(n4501), .A(n4371), .ZN(n3259) );
  AND4_X1 U3554 ( .A1(n3145), .A2(n3144), .A3(n3143), .A4(n3142), .ZN(n2996)
         );
  XOR2_X1 U3555 ( .A(n5571), .B(n2999), .Z(n2998) );
  INV_X1 U3556 ( .A(n2998), .ZN(n5279) );
  INV_X1 U3557 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n2999) );
  NAND2_X1 U3558 ( .A1(n3304), .A2(n3303), .ZN(n3323) );
  CLKBUF_X1 U3559 ( .A(n4390), .Z(n3017) );
  NAND2_X1 U3560 ( .A1(n3292), .A2(n3004), .ZN(n3001) );
  OR2_X1 U3561 ( .A1(n3003), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3002)
         );
  INV_X1 U3562 ( .A(n3310), .ZN(n3003) );
  AND2_X1 U3563 ( .A1(n3291), .A2(n3310), .ZN(n3004) );
  INV_X1 U3564 ( .A(n3284), .ZN(n3005) );
  INV_X1 U3565 ( .A(n3284), .ZN(n4620) );
  NAND2_X1 U3566 ( .A1(n4052), .A2(n4051), .ZN(n3008) );
  AND2_X1 U3567 ( .A1(n3488), .A2(n3487), .ZN(n3009) );
  NAND2_X1 U3568 ( .A1(n4052), .A2(n4051), .ZN(n4547) );
  AND2_X1 U3569 ( .A1(n3044), .A2(n4094), .ZN(n3014) );
  XNOR2_X1 U3570 ( .A(n4081), .B(n3548), .ZN(n4071) );
  NAND2_X1 U3571 ( .A1(n3043), .A2(n3014), .ZN(n3011) );
  OR2_X1 U3573 ( .A1(n3013), .A2(n5311), .ZN(n3012) );
  INV_X1 U3574 ( .A(n4094), .ZN(n3013) );
  AOI21_X2 U3576 ( .B1(n4477), .B2(n3674), .A(n4206), .ZN(n3439) );
  NAND2_X1 U3577 ( .A1(n4070), .A2(n4069), .ZN(n5083) );
  INV_X2 U3578 ( .A(n4912), .ZN(n3571) );
  XNOR2_X2 U3579 ( .A(n5183), .B(n3647), .ZN(n5264) );
  NOR2_X2 U3580 ( .A1(n4448), .A2(n4449), .ZN(n4450) );
  AND2_X2 U3581 ( .A1(n3088), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4339)
         );
  AND2_X2 U3582 ( .A1(n4333), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4340)
         );
  XNOR2_X1 U3583 ( .A(n4050), .B(n4541), .ZN(n4525) );
  AND2_X1 U3584 ( .A1(n3413), .A2(n3473), .ZN(n4477) );
  AOI21_X1 U3585 ( .B1(n3325), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3331), 
        .ZN(n3334) );
  NAND2_X1 U3586 ( .A1(n5758), .A2(n3083), .ZN(n5539) );
  AND2_X2 U3587 ( .A1(n5567), .A2(n4100), .ZN(n5758) );
  NAND2_X1 U3588 ( .A1(n4018), .A2(n4017), .ZN(n4050) );
  NAND2_X2 U3589 ( .A1(n3387), .A2(n3386), .ZN(n3428) );
  NAND2_X2 U3590 ( .A1(n3333), .A2(n3332), .ZN(n3444) );
  XNOR2_X1 U3591 ( .A(n4047), .B(n6188), .ZN(n4455) );
  NAND2_X1 U3592 ( .A1(n4046), .A2(n4045), .ZN(n4047) );
  NOR2_X2 U3593 ( .A1(n3202), .A2(n4620), .ZN(n3257) );
  NOR2_X2 U3594 ( .A1(n5487), .A2(n5488), .ZN(n5399) );
  INV_X2 U3595 ( .A(n3192), .ZN(n4246) );
  XNOR2_X1 U3596 ( .A(n3444), .B(n5008), .ZN(n4390) );
  NOR2_X4 U3597 ( .A1(n5439), .A2(n5442), .ZN(n5382) );
  NAND2_X1 U3598 ( .A1(n3089), .A2(n4392), .ZN(n4395) );
  NOR2_X2 U3599 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4202) );
  NOR2_X2 U3600 ( .A1(n3296), .A2(n4124), .ZN(n3674) );
  NAND2_X1 U3601 ( .A1(n3005), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3450) );
  AND2_X1 U3602 ( .A1(n4573), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4206) );
  AND2_X1 U3603 ( .A1(n5382), .A2(n3074), .ZN(n4234) );
  NOR2_X1 U3604 ( .A1(n4178), .A2(n3076), .ZN(n3074) );
  OR2_X1 U3605 ( .A1(n4225), .A2(n4224), .ZN(n4178) );
  AND2_X1 U3606 ( .A1(n3681), .A2(n5320), .ZN(n3073) );
  AND2_X1 U3607 ( .A1(n5693), .A2(n3038), .ZN(n4297) );
  NOR2_X1 U3608 ( .A1(n4299), .A2(n3039), .ZN(n3038) );
  NAND2_X1 U3609 ( .A1(n3040), .A2(n5692), .ZN(n3039) );
  INV_X1 U3610 ( .A(n4276), .ZN(n3040) );
  NAND2_X1 U3611 ( .A1(n4258), .A2(n4296), .ZN(n5355) );
  INV_X1 U3612 ( .A(n4297), .ZN(n4258) );
  NAND2_X1 U3613 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6430), .ZN(n3847) );
  NAND2_X1 U3614 ( .A1(n3861), .A2(n3837), .ZN(n3844) );
  XNOR2_X1 U3615 ( .A(n4406), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3843)
         );
  OR2_X1 U3616 ( .A1(n3882), .A2(n3537), .ZN(n3539) );
  OR2_X1 U3617 ( .A1(n3882), .A2(n3513), .ZN(n3515) );
  CLKBUF_X1 U3618 ( .A(n3390), .Z(n3750) );
  BUF_X1 U3619 ( .A(n3172), .Z(n4181) );
  OR2_X1 U3620 ( .A1(n3882), .A2(n4054), .ZN(n3486) );
  NAND2_X1 U3621 ( .A1(n4511), .A2(n4019), .ZN(n4235) );
  INV_X1 U3622 ( .A(n3348), .ZN(n4034) );
  NAND2_X1 U3623 ( .A1(n4580), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3449) );
  AOI21_X1 U3624 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6572), .A(n3839), 
        .ZN(n3841) );
  NOR2_X1 U3625 ( .A1(n3838), .A2(n3843), .ZN(n3839) );
  INV_X1 U3626 ( .A(n3844), .ZN(n3838) );
  AND2_X1 U3627 ( .A1(n3071), .A2(n5448), .ZN(n3070) );
  AND2_X1 U3628 ( .A1(n3072), .A2(n5460), .ZN(n3071) );
  AND2_X1 U3629 ( .A1(n3025), .A2(n5111), .ZN(n3068) );
  NAND2_X1 U3630 ( .A1(n4019), .A2(n4371), .ZN(n3903) );
  AOI21_X1 U3631 ( .B1(n5900), .B2(n3063), .A(n3028), .ZN(n3062) );
  INV_X1 U3632 ( .A(n5900), .ZN(n3064) );
  NAND2_X1 U3633 ( .A1(n5605), .A2(n3024), .ZN(n5567) );
  INV_X1 U3634 ( .A(n3978), .ZN(n4250) );
  NAND2_X1 U3635 ( .A1(n4989), .A2(n4296), .ZN(n3978) );
  NAND2_X1 U3636 ( .A1(n3904), .A2(n4989), .ZN(n4294) );
  AND2_X1 U3637 ( .A1(n3302), .A2(n3301), .ZN(n3305) );
  NAND2_X1 U3638 ( .A1(n3426), .A2(n3408), .ZN(n3066) );
  NOR2_X1 U3639 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4489), .ZN(n5132) );
  NAND2_X1 U3640 ( .A1(n3877), .A2(n4082), .ZN(n3883) );
  INV_X1 U3641 ( .A(n3314), .ZN(n6592) );
  INV_X1 U3642 ( .A(n3298), .ZN(n5958) );
  NOR2_X1 U3643 ( .A1(n5478), .A2(n3035), .ZN(n3034) );
  INV_X1 U3644 ( .A(n5490), .ZN(n3035) );
  NOR2_X1 U3645 ( .A1(n4514), .A2(n4370), .ZN(n4444) );
  OR2_X1 U3646 ( .A1(n5956), .A2(READY_N), .ZN(n4370) );
  AND2_X1 U3647 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n3898), .ZN(n4129)
         );
  INV_X1 U3648 ( .A(n5500), .ZN(n3696) );
  INV_X1 U3649 ( .A(n3551), .ZN(n3552) );
  NAND2_X1 U3650 ( .A1(n3919), .A2(n4296), .ZN(n5359) );
  INV_X1 U3651 ( .A(n4989), .ZN(n5358) );
  NOR2_X2 U3652 ( .A1(n5453), .A2(n3988), .ZN(n5388) );
  NAND2_X1 U3653 ( .A1(n5539), .A2(n4103), .ZN(n5899) );
  INV_X1 U3654 ( .A(n5241), .ZN(n3049) );
  INV_X1 U3655 ( .A(n3085), .ZN(n3046) );
  NOR2_X1 U3656 ( .A1(n5180), .A2(n5124), .ZN(n5186) );
  OR2_X1 U3657 ( .A1(n5178), .A2(n5177), .ZN(n5180) );
  NAND2_X1 U3658 ( .A1(n5075), .A2(n5056), .ZN(n5178) );
  AND2_X1 U3659 ( .A1(n4516), .A2(n4515), .ZN(n4533) );
  INV_X1 U3660 ( .A(n4533), .ZN(n4536) );
  INV_X1 U3661 ( .A(n6477), .ZN(n4506) );
  OR2_X1 U3662 ( .A1(n5377), .A2(n3033), .ZN(n3032) );
  AND2_X1 U3663 ( .A1(n6050), .A2(EBX_REG_30__SCAN_IN), .ZN(n3033) );
  INV_X1 U3664 ( .A(n5370), .ZN(n4292) );
  NAND2_X1 U3665 ( .A1(n4290), .A2(n4289), .ZN(n4293) );
  NOR2_X1 U3666 ( .A1(n4281), .A2(n4280), .ZN(n4282) );
  NAND2_X1 U3667 ( .A1(n4000), .A2(n5814), .ZN(n4011) );
  AND2_X1 U3668 ( .A1(n5362), .A2(n3902), .ZN(n6066) );
  INV_X1 U3669 ( .A(n5485), .ZN(n6086) );
  AND2_X1 U3670 ( .A1(n5507), .A2(n4377), .ZN(n6091) );
  INV_X1 U3671 ( .A(n5507), .ZN(n6093) );
  AND2_X1 U3672 ( .A1(n5507), .A2(n4378), .ZN(n5522) );
  INV_X1 U3673 ( .A(n4232), .ZN(n4233) );
  NAND2_X1 U3674 ( .A1(n4265), .A2(n4264), .ZN(n5669) );
  OR2_X1 U3675 ( .A1(n3845), .A2(n3835), .ZN(n3860) );
  AND2_X1 U3676 ( .A1(n3837), .A2(n3836), .ZN(n3859) );
  NAND2_X1 U3677 ( .A1(n3860), .A2(n3859), .ZN(n3861) );
  NAND2_X1 U3678 ( .A1(n3488), .A2(n3487), .ZN(n3518) );
  OR2_X1 U3679 ( .A1(n3365), .A2(n3364), .ZN(n4023) );
  INV_X1 U3680 ( .A(n4103), .ZN(n3063) );
  OR2_X1 U3681 ( .A1(n3536), .A2(n3535), .ZN(n4073) );
  OR2_X1 U3682 ( .A1(n3512), .A2(n3511), .ZN(n4056) );
  OR2_X1 U3683 ( .A1(n3484), .A2(n3483), .ZN(n4015) );
  OR2_X1 U3684 ( .A1(n3461), .A2(n3460), .ZN(n4044) );
  AOI22_X1 U3685 ( .A1(n4182), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3185), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3246) );
  NOR2_X1 U3686 ( .A1(n4235), .A2(n5338), .ZN(n4310) );
  NAND2_X1 U3687 ( .A1(n3203), .A2(n3192), .ZN(n4312) );
  INV_X1 U3688 ( .A(n4312), .ZN(n3293) );
  AND2_X1 U3689 ( .A1(n4310), .A2(n3295), .ZN(n3052) );
  AOI22_X1 U3690 ( .A1(n3390), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3146) );
  AOI22_X1 U3691 ( .A1(n3592), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3148) );
  NOR2_X1 U3692 ( .A1(n3832), .A2(n5384), .ZN(n3077) );
  NOR2_X1 U3693 ( .A1(n3784), .A2(n5476), .ZN(n3072) );
  OR2_X1 U3694 ( .A1(n5470), .A2(n5464), .ZN(n3784) );
  NAND2_X1 U3695 ( .A1(n3659), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3665)
         );
  INV_X1 U3696 ( .A(n5053), .ZN(n3069) );
  NOR2_X1 U3697 ( .A1(n3061), .A2(n4097), .ZN(n3060) );
  AND2_X1 U3698 ( .A1(n5606), .A2(n5780), .ZN(n4097) );
  INV_X1 U3699 ( .A(n4096), .ZN(n3061) );
  AND2_X1 U3700 ( .A1(n4082), .A2(n4085), .ZN(n4083) );
  INV_X1 U3701 ( .A(n4089), .ZN(n3057) );
  NAND2_X1 U3702 ( .A1(n3907), .A2(n3042), .ZN(n3910) );
  AND2_X1 U3703 ( .A1(n3306), .A2(n3305), .ZN(n3303) );
  AND2_X1 U3704 ( .A1(n4245), .A2(n4244), .ZN(n4530) );
  AND4_X1 U3705 ( .A1(n4243), .A2(n4314), .A3(n4242), .A4(n4241), .ZN(n4244)
         );
  AOI21_X1 U3706 ( .B1(n6483), .B2(n4433), .A(n5327), .ZN(n4489) );
  AND2_X2 U3707 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4422) );
  INV_X1 U3708 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6441) );
  INV_X1 U3709 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6437) );
  AND2_X1 U3710 ( .A1(n4418), .A2(n4417), .ZN(n6442) );
  AND2_X2 U3711 ( .A1(n3450), .A2(n3449), .ZN(n3882) );
  OAI21_X1 U3712 ( .B1(n3879), .B2(n3883), .A(n3878), .ZN(n3880) );
  INV_X1 U3713 ( .A(n3891), .ZN(n3879) );
  AOI222_X1 U3714 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n3840), .B1(
        INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6461), .C1(n3840), .C2(n6461), 
        .ZN(n3889) );
  NAND2_X1 U3715 ( .A1(n3293), .A2(n3052), .ZN(n5956) );
  NOR2_X1 U3716 ( .A1(n6528), .A2(n5429), .ZN(n5412) );
  INV_X1 U3717 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6023) );
  AND2_X1 U3718 ( .A1(n6590), .A2(EBX_REG_31__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U3719 ( .A1(n6590), .A2(n3996), .ZN(n6069) );
  OR2_X1 U3720 ( .A1(n4287), .A2(n3524), .ZN(n4166) );
  AND2_X1 U3721 ( .A1(n3957), .A2(n3956), .ZN(n5490) );
  NAND2_X1 U3722 ( .A1(n3917), .A2(n3916), .ZN(n4995) );
  INV_X1 U3723 ( .A(n4984), .ZN(n3916) );
  INV_X1 U3724 ( .A(n4985), .ZN(n3917) );
  OR2_X1 U3725 ( .A1(n6453), .A2(n4527), .ZN(n4322) );
  AOI21_X1 U3726 ( .B1(n4053), .B2(n3674), .A(n3523), .ZN(n4449) );
  AND2_X1 U3727 ( .A1(n4352), .A2(n4502), .ZN(n6097) );
  AOI21_X1 U3728 ( .B1(n4205), .B2(n4204), .A(n4203), .ZN(n4232) );
  NOR2_X1 U3729 ( .A1(n4175), .A2(n4170), .ZN(n4162) );
  INV_X1 U3730 ( .A(n5554), .ZN(n4271) );
  AND2_X1 U3731 ( .A1(n4131), .A2(n4130), .ZN(n5553) );
  NOR2_X1 U3732 ( .A1(n3816), .A2(n3199), .ZN(n3827) );
  NAND2_X1 U3733 ( .A1(n3827), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3897)
         );
  NAND2_X1 U3734 ( .A1(n3808), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3816)
         );
  AND2_X1 U3735 ( .A1(n3802), .A2(n3801), .ZN(n5460) );
  AND2_X1 U3736 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n3198), .ZN(n3781)
         );
  INV_X1 U3737 ( .A(n3764), .ZN(n3198) );
  NAND2_X1 U3738 ( .A1(n3781), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3800)
         );
  NOR2_X1 U3739 ( .A1(n3728), .A2(n3197), .ZN(n3731) );
  NAND2_X1 U3740 ( .A1(n3731), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3764)
         );
  AND2_X1 U3741 ( .A1(n3682), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3712)
         );
  NOR2_X1 U3742 ( .A1(n3665), .A2(n5413), .ZN(n3682) );
  NOR2_X1 U3743 ( .A1(n3630), .A2(n3631), .ZN(n3659) );
  CLKBUF_X1 U3744 ( .A(n5265), .Z(n5266) );
  NAND2_X1 U3745 ( .A1(n3616), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3630)
         );
  INV_X1 U3746 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3631) );
  NOR2_X1 U3747 ( .A1(n3612), .A2(n5170), .ZN(n3616) );
  CLKBUF_X1 U3748 ( .A(n5120), .Z(n5121) );
  NAND2_X1 U3749 ( .A1(n3587), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3612)
         );
  NOR2_X1 U3750 ( .A1(n3572), .A2(n5107), .ZN(n3587) );
  NAND2_X1 U3751 ( .A1(n3555), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3572)
         );
  NOR2_X1 U3752 ( .A1(n3520), .A2(n6038), .ZN(n3525) );
  NAND2_X1 U3753 ( .A1(n3525), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3549)
         );
  NAND2_X1 U3754 ( .A1(n3196), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3520)
         );
  INV_X1 U3755 ( .A(n3494), .ZN(n3196) );
  INV_X1 U3756 ( .A(n3436), .ZN(n3467) );
  NAND2_X1 U3757 ( .A1(n3467), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3494)
         );
  NAND2_X1 U3758 ( .A1(n3472), .A2(n3471), .ZN(n4389) );
  NAND2_X1 U3759 ( .A1(n4438), .A2(n4031), .ZN(n6136) );
  NAND2_X1 U3760 ( .A1(n6453), .A2(n4506), .ZN(n4514) );
  NAND2_X1 U3761 ( .A1(n3065), .A2(n4221), .ZN(n5526) );
  NOR2_X2 U3762 ( .A1(n5551), .A2(n5656), .ZN(n5529) );
  NOR2_X2 U3763 ( .A1(n5471), .A2(n3969), .ZN(n5466) );
  OR2_X1 U3764 ( .A1(n5606), .A2(n4099), .ZN(n4100) );
  NAND2_X1 U3765 ( .A1(n5497), .A2(n5490), .ZN(n5492) );
  OAI21_X1 U3766 ( .B1(n5631), .B2(n5633), .A(n5632), .ZN(n4095) );
  AND3_X1 U3767 ( .A1(n3951), .A2(n3975), .A3(n3950), .ZN(n5415) );
  AOI21_X1 U3768 ( .B1(n3047), .B2(n3045), .A(n3023), .ZN(n3044) );
  INV_X1 U3769 ( .A(n3081), .ZN(n3045) );
  AND3_X1 U3770 ( .A1(n3939), .A2(n3975), .A3(n3938), .ZN(n5177) );
  AND2_X1 U3771 ( .A1(n3937), .A2(n3936), .ZN(n5056) );
  NAND2_X1 U3772 ( .A1(n3079), .A2(n3037), .ZN(n3036) );
  INV_X1 U3773 ( .A(n5073), .ZN(n3037) );
  NAND2_X1 U3774 ( .A1(n3930), .A2(n3079), .ZN(n5074) );
  INV_X1 U3775 ( .A(n4919), .ZN(n3930) );
  OAI211_X1 U3776 ( .C1(n3406), .C2(n3295), .A(n3405), .B(n3404), .ZN(n3424)
         );
  INV_X1 U3777 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4406) );
  NOR2_X1 U3778 ( .A1(n3299), .A2(n3298), .ZN(n3054) );
  AND2_X1 U3779 ( .A1(n4478), .A2(n4480), .ZN(n6281) );
  INV_X1 U3780 ( .A(n4752), .ZN(n4746) );
  OR2_X1 U3781 ( .A1(n6311), .A2(n4482), .ZN(n4752) );
  INV_X1 U3782 ( .A(n4853), .ZN(n4782) );
  NOR2_X1 U3783 ( .A1(n6370), .A2(n4482), .ZN(n4854) );
  INV_X1 U3784 ( .A(n3295), .ZN(n4580) );
  INV_X1 U3785 ( .A(n5006), .ZN(n5198) );
  INV_X1 U3786 ( .A(n4575), .ZN(n6377) );
  INV_X1 U3787 ( .A(n5132), .ZN(n4667) );
  OR2_X1 U3788 ( .A1(n6560), .A2(n4489), .ZN(n4668) );
  OR2_X1 U3789 ( .A1(n4323), .A2(n4111), .ZN(n6457) );
  NAND2_X2 U3790 ( .A1(n3885), .A2(n3884), .ZN(n6453) );
  OR2_X1 U3791 ( .A1(n3889), .A2(n3883), .ZN(n3884) );
  OAI21_X1 U3792 ( .B1(n3889), .B2(n3882), .A(n3881), .ZN(n3885) );
  AOI21_X1 U3793 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6474), .A(n3880), 
        .ZN(n3881) );
  NOR2_X1 U3794 ( .A1(n5836), .A2(n5847), .ZN(n5831) );
  INV_X1 U3795 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6038) );
  INV_X1 U3796 ( .A(n6050), .ZN(n6078) );
  INV_X1 U3797 ( .A(n4342), .ZN(n4763) );
  AND2_X1 U3798 ( .A1(n6068), .A2(n4005), .ZN(n6071) );
  AND2_X1 U3799 ( .A1(n6590), .A2(n4004), .ZN(n6050) );
  OAI21_X1 U3800 ( .B1(n4375), .B2(n4374), .A(n4506), .ZN(n4376) );
  INV_X1 U3801 ( .A(n6091), .ZN(n5524) );
  INV_X1 U3802 ( .A(n5522), .ZN(n5299) );
  NAND2_X1 U3804 ( .A1(n4444), .A2(n4371), .ZN(n4607) );
  AOI21_X1 U3805 ( .B1(n5441), .B2(n5384), .A(n5383), .ZN(n5901) );
  INV_X1 U3807 ( .A(n6145), .ZN(n6137) );
  INV_X1 U3808 ( .A(n6148), .ZN(n5610) );
  INV_X1 U3809 ( .A(n6143), .ZN(n5613) );
  XNOR2_X1 U3810 ( .A(n5361), .B(n5360), .ZN(n5659) );
  AND2_X1 U3811 ( .A1(n5280), .A2(n5929), .ZN(n5782) );
  INV_X1 U3812 ( .A(n5920), .ZN(n5712) );
  AND2_X1 U3813 ( .A1(n5732), .A2(n5738), .ZN(n5730) );
  NAND2_X1 U3814 ( .A1(n3048), .A2(n3047), .ZN(n5278) );
  NAND2_X1 U3815 ( .A1(n3049), .A2(n3081), .ZN(n3048) );
  NAND2_X1 U3816 ( .A1(n4536), .A2(n6454), .ZN(n5929) );
  INV_X1 U3817 ( .A(n6218), .ZN(n6170) );
  OR2_X1 U3818 ( .A1(n5280), .A2(n6204), .ZN(n6198) );
  AND2_X1 U3819 ( .A1(n6225), .A2(n6227), .ZN(n6204) );
  NAND2_X1 U3820 ( .A1(n4536), .A2(n4535), .ZN(n6218) );
  INV_X1 U3821 ( .A(n6206), .ZN(n6223) );
  CLKBUF_X1 U3822 ( .A(n4481), .Z(n4482) );
  CLKBUF_X1 U3823 ( .A(n4407), .Z(n4408) );
  INV_X1 U3824 ( .A(n4478), .ZN(n5801) );
  INV_X1 U3825 ( .A(n6568), .ZN(n6587) );
  INV_X1 U3826 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6461) );
  NOR2_X1 U3827 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n4346) );
  CLKBUF_X1 U3828 ( .A(n3094), .Z(n5336) );
  INV_X1 U3829 ( .A(n6467), .ZN(n5327) );
  OAI21_X1 U3830 ( .B1(n5168), .B2(n6562), .A(n5141), .ZN(n5163) );
  NAND2_X1 U3831 ( .A1(n4492), .A2(n4782), .ZN(n5047) );
  INV_X1 U3832 ( .A(n6306), .ZN(n4899) );
  NOR2_X2 U3833 ( .A1(n4752), .A2(n4853), .ZN(n5236) );
  INV_X1 U3834 ( .A(n6325), .ZN(n6356) );
  INV_X1 U3835 ( .A(n6368), .ZN(n6328) );
  INV_X1 U3836 ( .A(n6383), .ZN(n6332) );
  INV_X1 U3837 ( .A(n6395), .ZN(n6340) );
  INV_X1 U3838 ( .A(n6401), .ZN(n6344) );
  INV_X1 U3839 ( .A(n6407), .ZN(n6348) );
  INV_X1 U3840 ( .A(n6413), .ZN(n6352) );
  AND2_X1 U3841 ( .A1(n4861), .A2(n4860), .ZN(n4906) );
  NOR2_X1 U3842 ( .A1(n4488), .A2(n4667), .ZN(n6389) );
  NOR2_X1 U3843 ( .A1(n4584), .A2(n4667), .ZN(n6395) );
  NOR2_X1 U3844 ( .A1(n6770), .A2(n4667), .ZN(n6407) );
  NOR2_X1 U3845 ( .A1(n4609), .A2(n4667), .ZN(n6413) );
  AND2_X1 U3846 ( .A1(n4419), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U3847 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6453), .ZN(n6467) );
  INV_X1 U3848 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6474) );
  NAND2_X1 U3849 ( .A1(n6470), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6477) );
  OAI211_X1 U3850 ( .C1(n5669), .C2(n6061), .A(n5381), .B(n3031), .ZN(U2797)
         );
  AOI21_X1 U3851 ( .B1(n5536), .B2(n6033), .A(n3032), .ZN(n3031) );
  OR2_X1 U3852 ( .A1(n5674), .A2(n6061), .ZN(n4301) );
  NOR2_X1 U3853 ( .A1(n4293), .A2(n4292), .ZN(n4302) );
  NAND2_X1 U3854 ( .A1(n4285), .A2(n4284), .ZN(U2799) );
  AND2_X1 U3855 ( .A1(n4283), .A2(n4282), .ZN(n4284) );
  OR2_X1 U3856 ( .A1(n5682), .A2(n6061), .ZN(n4283) );
  NAND2_X1 U3857 ( .A1(n4011), .A2(n4010), .ZN(n4012) );
  AND2_X1 U3858 ( .A1(n4267), .A2(n4266), .ZN(n4268) );
  NAND2_X1 U3859 ( .A1(n3749), .A2(n3748), .ZN(n5462) );
  NAND2_X1 U3860 ( .A1(n3664), .A2(n5320), .ZN(n5322) );
  AND2_X1 U3861 ( .A1(n3571), .A2(n3068), .ZN(n3018) );
  AND2_X1 U3862 ( .A1(n3749), .A2(n3072), .ZN(n5458) );
  AND2_X1 U3863 ( .A1(n3749), .A2(n3071), .ZN(n5447) );
  NAND2_X1 U3864 ( .A1(n3553), .A2(n3552), .ZN(n4911) );
  INV_X1 U3865 ( .A(n3067), .ZN(n5054) );
  NAND2_X2 U3866 ( .A1(n4586), .A2(n3295), .ZN(n3919) );
  AND2_X2 U3867 ( .A1(n4615), .A2(n3295), .ZN(n3314) );
  AND2_X1 U3868 ( .A1(n3059), .A2(n3060), .ZN(n5604) );
  NAND2_X1 U3869 ( .A1(n5899), .A2(n5900), .ZN(n3020) );
  INV_X1 U3870 ( .A(n3065), .ZN(n5559) );
  OAI21_X1 U3871 ( .B1(n5539), .B2(n3064), .A(n3062), .ZN(n3065) );
  NAND2_X1 U3872 ( .A1(n5382), .A2(n3831), .ZN(n3021) );
  NAND2_X1 U3873 ( .A1(n3059), .A2(n4096), .ZN(n5617) );
  NOR2_X1 U3874 ( .A1(n5618), .A2(n6167), .ZN(n3022) );
  AND2_X1 U3875 ( .A1(n5618), .A2(n2999), .ZN(n3023) );
  AND2_X1 U3876 ( .A1(n3060), .A2(n4098), .ZN(n3024) );
  NAND2_X1 U3877 ( .A1(n3203), .A2(n3202), .ZN(n3297) );
  AND2_X1 U3878 ( .A1(n6086), .A2(n4246), .ZN(n6081) );
  INV_X1 U3879 ( .A(n5856), .ZN(n6033) );
  AND2_X2 U3880 ( .A1(n4397), .A2(n4339), .ZN(n3390) );
  NAND2_X1 U3881 ( .A1(n5497), .A2(n3034), .ZN(n5471) );
  BUF_X1 U3882 ( .A(n3355), .Z(n3733) );
  NAND2_X1 U3883 ( .A1(n3466), .A2(n3465), .ZN(n4479) );
  NAND2_X1 U3884 ( .A1(n3571), .A2(n3570), .ZN(n5052) );
  AND2_X1 U3885 ( .A1(n3570), .A2(n3069), .ZN(n3025) );
  NAND2_X1 U3886 ( .A1(n3058), .A2(n4089), .ZN(n5113) );
  AND2_X1 U3887 ( .A1(n3048), .A2(n3046), .ZN(n3026) );
  AND2_X1 U3888 ( .A1(n5338), .A2(n4371), .ZN(n4082) );
  NAND2_X1 U3889 ( .A1(n3571), .A2(n3025), .ZN(n3067) );
  NOR2_X1 U3890 ( .A1(n5414), .A2(n5415), .ZN(n3027) );
  INV_X1 U3891 ( .A(n3076), .ZN(n3075) );
  NAND2_X1 U3892 ( .A1(n3077), .A2(n5553), .ZN(n3076) );
  NAND2_X1 U3893 ( .A1(n5457), .A2(n5456), .ZN(n5450) );
  AND2_X1 U3894 ( .A1(n5606), .A2(n5919), .ZN(n3028) );
  AND2_X1 U3895 ( .A1(n5122), .A2(n3068), .ZN(n3029) );
  NAND2_X1 U3896 ( .A1(n3055), .A2(n3054), .ZN(n4324) );
  AND3_X1 U3897 ( .A1(n4586), .A2(n3282), .A3(n4511), .ZN(n3030) );
  XNOR2_X1 U3898 ( .A(n4923), .B(n3910), .ZN(n4756) );
  INV_X1 U3899 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4333) );
  NOR2_X2 U3900 ( .A1(n4919), .A2(n3036), .ZN(n5075) );
  NAND3_X1 U3901 ( .A1(n3904), .A2(n4989), .A3(n4990), .ZN(n3042) );
  NAND2_X1 U3902 ( .A1(n5241), .A2(n3047), .ZN(n3043) );
  NAND2_X1 U3903 ( .A1(n2990), .A2(n3044), .ZN(n5310) );
  NOR2_X2 U3904 ( .A1(n3085), .A2(n2998), .ZN(n3047) );
  INV_X1 U3905 ( .A(n3297), .ZN(n3055) );
  NAND2_X1 U3906 ( .A1(n3050), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3306) );
  NAND3_X1 U3907 ( .A1(n4519), .A2(n4324), .A3(n3051), .ZN(n3050) );
  NAND3_X1 U3908 ( .A1(n3052), .A2(n3293), .A3(n3294), .ZN(n3051) );
  NAND2_X1 U3909 ( .A1(n3053), .A2(n5339), .ZN(n4519) );
  INV_X1 U3910 ( .A(n4373), .ZN(n3053) );
  NAND2_X1 U3911 ( .A1(n5067), .A2(n5068), .ZN(n3058) );
  NAND2_X1 U3912 ( .A1(n3058), .A2(n3056), .ZN(n4092) );
  NAND2_X1 U3913 ( .A1(n5623), .A2(n5624), .ZN(n5605) );
  CLKBUF_X1 U3914 ( .A(n5605), .Z(n3059) );
  OAI21_X1 U3915 ( .B1(n3415), .B2(n3414), .A(n3066), .ZN(n3410) );
  AND2_X2 U3916 ( .A1(n3571), .A2(n3029), .ZN(n5120) );
  NAND2_X1 U3917 ( .A1(n3749), .A2(n3070), .ZN(n5439) );
  NAND2_X1 U3918 ( .A1(n3664), .A2(n3073), .ZN(n5410) );
  INV_X1 U3919 ( .A(n5410), .ZN(n3697) );
  AND2_X1 U3920 ( .A1(n5382), .A2(n3077), .ZN(n4132) );
  NAND2_X1 U3921 ( .A1(n5382), .A2(n3075), .ZN(n5554) );
  NAND2_X1 U3922 ( .A1(n4273), .A2(n4225), .ZN(n4227) );
  NAND2_X1 U3923 ( .A1(n4271), .A2(n4270), .ZN(n4273) );
  NAND2_X1 U3924 ( .A1(n4227), .A2(n4226), .ZN(n4286) );
  INV_X1 U3925 ( .A(n5529), .ZN(n4222) );
  OR2_X1 U3926 ( .A1(n5539), .A2(n5538), .ZN(n5550) );
  INV_X1 U3927 ( .A(n4275), .ZN(n4285) );
  NAND2_X1 U3928 ( .A1(n4477), .A2(n4082), .ZN(n4039) );
  NAND2_X1 U3929 ( .A1(n3444), .A2(n3336), .ZN(n4407) );
  NOR2_X1 U3930 ( .A1(n5567), .A2(n3959), .ZN(n5568) );
  NAND2_X1 U3931 ( .A1(n3407), .A2(n3424), .ZN(n3426) );
  INV_X1 U3932 ( .A(n4565), .ZN(n3501) );
  OAI21_X1 U3933 ( .B1(n3428), .B2(STATE2_REG_0__SCAN_IN), .A(n3422), .ZN(
        n3407) );
  OR2_X1 U3934 ( .A1(n3411), .A2(n3412), .ZN(n3413) );
  INV_X1 U3935 ( .A(n5536), .ZN(n5514) );
  NAND2_X1 U3936 ( .A1(n5536), .A2(n6082), .ZN(n4269) );
  INV_X1 U3937 ( .A(n3543), .ZN(n3544) );
  NAND2_X1 U3938 ( .A1(n6144), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4029)
         );
  INV_X1 U3939 ( .A(n4482), .ZN(n4676) );
  NAND2_X1 U3940 ( .A1(n4039), .A2(n4038), .ZN(n6134) );
  NOR2_X1 U3941 ( .A1(n4478), .A2(n4042), .ZN(n3078) );
  AND2_X1 U3942 ( .A1(n3929), .A2(n4916), .ZN(n3079) );
  AND2_X1 U3943 ( .A1(n5571), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3080)
         );
  NAND2_X1 U3944 ( .A1(n5606), .A2(n4093), .ZN(n3081) );
  AND2_X1 U3945 ( .A1(n5606), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3082)
         );
  OR2_X1 U3946 ( .A1(n5618), .A2(n4102), .ZN(n3083) );
  INV_X1 U3947 ( .A(n6082), .ZN(n5506) );
  AND2_X1 U3948 ( .A1(n6086), .A2(n3192), .ZN(n6082) );
  NOR2_X1 U3949 ( .A1(n5205), .A2(n5128), .ZN(n3084) );
  INV_X1 U3950 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U3951 ( .A1(n5252), .A2(n5254), .ZN(n3085) );
  NAND2_X1 U3952 ( .A1(n4211), .A2(n6568), .ZN(n6371) );
  AND2_X1 U3953 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3086) );
  INV_X1 U3954 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5107) );
  AOI21_X1 U3955 ( .B1(n4322), .B2(n4249), .A(n6477), .ZN(n5504) );
  AND3_X1 U3956 ( .A1(n6572), .A2(n5014), .A3(n5013), .ZN(n3087) );
  INV_X1 U3957 ( .A(n6133), .ZN(n6190) );
  INV_X2 U3958 ( .A(n4090), .ZN(n5571) );
  AND2_X2 U3959 ( .A1(n4340), .A2(n4397), .ZN(n3451) );
  AND2_X2 U3960 ( .A1(n4392), .A2(n4397), .ZN(n3367) );
  INV_X1 U3961 ( .A(n5382), .ZN(n5441) );
  NOR2_X1 U3962 ( .A1(n5958), .A2(n3848), .ZN(n3870) );
  NAND2_X1 U3963 ( .A1(n6437), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3834) );
  NAND2_X1 U3964 ( .A1(n6441), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3837) );
  INV_X1 U3965 ( .A(n4023), .ZN(n3383) );
  INV_X1 U3966 ( .A(n4015), .ZN(n4054) );
  NOR2_X1 U3967 ( .A1(n3846), .A2(n3847), .ZN(n3845) );
  INV_X1 U3968 ( .A(n5384), .ZN(n3831) );
  AND2_X1 U3969 ( .A1(n3486), .A2(n3485), .ZN(n3489) );
  OR2_X1 U3970 ( .A1(n3347), .A2(n3346), .ZN(n3348) );
  INV_X1 U3971 ( .A(n4085), .ZN(n3547) );
  OAI21_X1 U3972 ( .B1(n3877), .B2(n3879), .A(n3876), .ZN(n3878) );
  NAND2_X1 U3973 ( .A1(n3515), .A2(n3514), .ZN(n3516) );
  INV_X1 U3974 ( .A(n5411), .ZN(n3681) );
  INV_X1 U3975 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n4124) );
  INV_X1 U3976 ( .A(n5092), .ZN(n3570) );
  OR2_X1 U3977 ( .A1(n3401), .A2(n3400), .ZN(n4022) );
  NOR2_X1 U3978 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n3842), .ZN(n3891)
         );
  AND2_X1 U3979 ( .A1(n3539), .A2(n3538), .ZN(n3543) );
  NAND2_X1 U3980 ( .A1(n3244), .A2(n3006), .ZN(n3290) );
  INV_X1 U3981 ( .A(n5476), .ZN(n3748) );
  OR2_X1 U3982 ( .A1(n2987), .A2(n3648), .ZN(n5319) );
  OR2_X1 U3983 ( .A1(n5606), .A2(n5945), .ZN(n5632) );
  AND2_X1 U3984 ( .A1(n3934), .A2(n3933), .ZN(n5073) );
  NAND2_X1 U3985 ( .A1(n4245), .A2(n3322), .ZN(n3384) );
  OR2_X1 U3986 ( .A1(n4111), .A2(n3903), .ZN(n4531) );
  NOR2_X1 U3987 ( .A1(n3800), .A2(n5588), .ZN(n3808) );
  INV_X1 U3988 ( .A(n6068), .ZN(n4758) );
  OR2_X1 U3989 ( .A1(n4201), .A2(n5376), .ZN(n3900) );
  NAND2_X1 U3990 ( .A1(n4129), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4175)
         );
  OR2_X1 U3991 ( .A1(n5904), .A2(n3524), .ZN(n3829) );
  OR2_X1 U3992 ( .A1(n4344), .A2(n6474), .ZN(n4173) );
  INV_X1 U3993 ( .A(n4202), .ZN(n3524) );
  INV_X1 U3994 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5527) );
  AND2_X1 U3995 ( .A1(n4679), .A2(n6568), .ZN(n4681) );
  NOR2_X1 U3996 ( .A1(n4491), .A2(n4482), .ZN(n4492) );
  AND2_X1 U3997 ( .A1(n3017), .A2(n6315), .ZN(n6363) );
  NAND2_X1 U3998 ( .A1(n3448), .A2(n3447), .ZN(n5008) );
  NOR2_X1 U3999 ( .A1(n6662), .A2(n4291), .ZN(n5378) );
  NOR2_X1 U4000 ( .A1(n6039), .A2(n4007), .ZN(n4008) );
  INV_X1 U4001 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5413) );
  NOR3_X1 U4002 ( .A1(n4758), .A2(n3993), .A3(n5174), .ZN(n5269) );
  NOR2_X1 U4003 ( .A1(n3549), .A2(n6023), .ZN(n3555) );
  AND2_X1 U4004 ( .A1(n4217), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4005) );
  AND3_X1 U4005 ( .A1(n3954), .A2(n3975), .A3(n3953), .ZN(n5495) );
  XNOR2_X1 U4006 ( .A(n3900), .B(n3899), .ZN(n4217) );
  AND2_X1 U4007 ( .A1(n3730), .A2(n3729), .ZN(n5400) );
  OR2_X1 U4008 ( .A1(n3020), .A2(n4105), .ZN(n4106) );
  OR2_X1 U4009 ( .A1(n5704), .A2(n5706), .ZN(n5699) );
  INV_X1 U4010 ( .A(n5758), .ZN(n5760) );
  AND2_X1 U4011 ( .A1(n6225), .A2(n5930), .ZN(n5280) );
  OR2_X1 U4012 ( .A1(n4514), .A2(n4513), .ZN(n4515) );
  OR2_X1 U4013 ( .A1(n3017), .A2(n4744), .ZN(n6233) );
  NAND2_X1 U4014 ( .A1(n4492), .A2(n4853), .ZN(n5166) );
  AND2_X1 U4015 ( .A1(n4482), .A2(n4853), .ZN(n5006) );
  OR2_X1 U4016 ( .A1(n3424), .A2(n3423), .ZN(n3425) );
  OR2_X1 U4017 ( .A1(n6311), .A2(n5198), .ZN(n6325) );
  NAND2_X1 U4018 ( .A1(n4854), .A2(n4853), .ZN(n4978) );
  INV_X1 U4019 ( .A(n4980), .ZN(n4821) );
  INV_X1 U4020 ( .A(n4309), .ZN(n6590) );
  INV_X1 U4021 ( .A(n5659), .ZN(n5369) );
  NOR2_X1 U4022 ( .A1(n4009), .A2(n4008), .ZN(n4010) );
  AND2_X1 U4023 ( .A1(n3973), .A2(n3972), .ZN(n5465) );
  NAND2_X1 U4024 ( .A1(n4309), .A2(n3896), .ZN(n6068) );
  AND2_X1 U4025 ( .A1(n6068), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6062) );
  INV_X1 U4026 ( .A(n6069), .ZN(n6054) );
  OR2_X1 U4027 ( .A1(n5669), .A2(n5503), .ZN(n4267) );
  INV_X1 U4028 ( .A(n5504), .ZN(n5485) );
  INV_X1 U4029 ( .A(n4625), .ZN(n4660) );
  INV_X1 U4030 ( .A(n4607), .ZN(n4649) );
  INV_X1 U4031 ( .A(n4625), .ZN(n4606) );
  NAND2_X1 U4032 ( .A1(n3712), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3728)
         );
  NAND2_X1 U4033 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3436) );
  NAND2_X1 U4034 ( .A1(n5526), .A2(n4222), .ZN(n4223) );
  NOR2_X1 U4035 ( .A1(n6152), .A2(n5646), .ZN(n5923) );
  NOR2_X1 U4036 ( .A1(n5286), .A2(n6198), .ZN(n5747) );
  INV_X1 U4037 ( .A(n5782), .ZN(n6212) );
  INV_X1 U4038 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4419) );
  INV_X1 U4039 ( .A(n4933), .ZN(n4888) );
  INV_X1 U4040 ( .A(n4930), .ZN(n6275) );
  AND2_X1 U4041 ( .A1(n6281), .A2(n4714), .ZN(n6306) );
  AND2_X1 U4042 ( .A1(n6281), .A2(n5006), .ZN(n6304) );
  OAI21_X1 U4043 ( .B1(n4718), .B2(n4719), .A(n4717), .ZN(n4897) );
  AND2_X1 U4044 ( .A1(n5202), .A2(n3017), .ZN(n6316) );
  INV_X1 U4045 ( .A(n6319), .ZN(n6355) );
  OR4_X1 U4046 ( .A1(n4858), .A2(n4857), .A3(n5203), .A4(n4856), .ZN(n4905) );
  NAND2_X1 U4047 ( .A1(n4042), .A2(n5801), .ZN(n6311) );
  AND2_X1 U4048 ( .A1(n4854), .A2(n4782), .ZN(n4980) );
  NOR2_X1 U4049 ( .A1(n6749), .A2(n4667), .ZN(n6368) );
  NOR2_X1 U4050 ( .A1(n4614), .A2(n4667), .ZN(n6383) );
  NOR2_X1 U4051 ( .A1(n6751), .A2(n4667), .ZN(n6401) );
  NOR2_X1 U4052 ( .A1(n6617), .A2(n4667), .ZN(n6420) );
  OR2_X1 U4053 ( .A1(n4520), .A2(n6592), .ZN(n6465) );
  OR2_X1 U4054 ( .A1(n4514), .A2(n5956), .ZN(n4306) );
  AND2_X1 U4055 ( .A1(n4302), .A2(n4301), .ZN(n4303) );
  INV_X1 U4056 ( .A(n6062), .ZN(n6039) );
  NAND2_X1 U4057 ( .A1(n6068), .A2(n3901), .ZN(n5856) );
  INV_X1 U4058 ( .A(n6066), .ZN(n6061) );
  NAND2_X1 U4059 ( .A1(n4607), .A2(n4376), .ZN(n5507) );
  INV_X1 U4060 ( .A(n6097), .ZN(n6131) );
  OR2_X1 U4061 ( .A1(n4514), .A2(n6465), .ZN(n4445) );
  OR2_X2 U4062 ( .A1(n4514), .A2(n6457), .ZN(n6145) );
  AND2_X1 U4063 ( .A1(n5730), .A2(n5653), .ZN(n5920) );
  NOR2_X1 U4064 ( .A1(n5936), .A2(n5747), .ZN(n6152) );
  NAND2_X1 U4065 ( .A1(n4536), .A2(n4524), .ZN(n6206) );
  INV_X1 U4066 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6430) );
  INV_X1 U4067 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6572) );
  NAND2_X1 U4068 ( .A1(n4677), .A2(n4782), .ZN(n4933) );
  AOI21_X1 U4069 ( .B1(n4701), .B2(n4700), .A(n4699), .ZN(n4927) );
  NAND2_X1 U4070 ( .A1(n3078), .A2(n4714), .ZN(n6280) );
  NAND2_X1 U4071 ( .A1(n4746), .A2(n4853), .ZN(n4904) );
  AOI22_X1 U4072 ( .A1(n5207), .A2(n6316), .B1(n5205), .B2(n5204), .ZN(n5238)
         );
  INV_X1 U4073 ( .A(n6389), .ZN(n6336) );
  INV_X1 U4074 ( .A(n6420), .ZN(n6360) );
  OR2_X1 U4075 ( .A1(n6311), .A2(n6228), .ZN(n6319) );
  AND3_X1 U4076 ( .A1(n4788), .A2(n5013), .A3(n4787), .ZN(n4826) );
  OR2_X1 U4077 ( .A1(n6370), .A2(n6228), .ZN(n6428) );
  INV_X1 U4078 ( .A(n6558), .ZN(n6554) );
  INV_X1 U4079 ( .A(n6550), .ZN(n6549) );
  OAI21_X1 U4080 ( .B1(n4286), .B2(n5856), .A(n4303), .ZN(U2798) );
  NAND2_X1 U4081 ( .A1(n4269), .A2(n4268), .ZN(U2829) );
  INV_X1 U4082 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3088) );
  AND2_X2 U4083 ( .A1(n4339), .A2(n3089), .ZN(n3250) );
  AOI22_X1 U4084 ( .A1(n4151), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3093) );
  AND2_X2 U4085 ( .A1(n4340), .A2(n3089), .ZN(n3592) );
  BUF_X1 U4086 ( .A(n3374), .Z(n3388) );
  AOI22_X1 U4087 ( .A1(n3592), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3092) );
  AOI22_X1 U4088 ( .A1(n3790), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3091) );
  AND2_X2 U4089 ( .A1(n3089), .A2(n3095), .ZN(n3172) );
  AOI22_X1 U4090 ( .A1(n4181), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3090) );
  NAND4_X1 U4091 ( .A1(n3093), .A2(n3092), .A3(n3091), .A4(n3090), .ZN(n3101)
         );
  INV_X2 U4092 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3094) );
  NOR2_X4 U4093 ( .A1(n3094), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4397)
         );
  AOI22_X1 U4094 ( .A1(n3354), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3015), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3099) );
  AOI22_X1 U4095 ( .A1(n3337), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3098) );
  AND2_X4 U4096 ( .A1(n4392), .A2(n4422), .ZN(n3272) );
  INV_X1 U4097 ( .A(n3272), .ZN(n4400) );
  AOI22_X1 U4098 ( .A1(n3750), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3097) );
  AND2_X2 U4099 ( .A1(n4397), .A2(n3095), .ZN(n3355) );
  AND2_X2 U4100 ( .A1(n3095), .A2(n4422), .ZN(n4182) );
  AOI22_X1 U4101 ( .A1(n3733), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3096) );
  NAND4_X1 U4102 ( .A1(n3099), .A2(n3098), .A3(n3097), .A4(n3096), .ZN(n3100)
         );
  NOR2_X1 U4103 ( .A1(n3101), .A2(n3100), .ZN(n3821) );
  AOI22_X1 U4104 ( .A1(n3592), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3105) );
  AOI22_X1 U4105 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n3337), .B1(n3790), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3104) );
  AOI22_X1 U4106 ( .A1(n4181), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3103) );
  AOI22_X1 U4107 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n3015), .B1(n4145), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3102) );
  NAND4_X1 U4108 ( .A1(n3105), .A2(n3104), .A3(n3103), .A4(n3102), .ZN(n3111)
         );
  AOI22_X1 U4109 ( .A1(n4151), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3109) );
  AOI22_X1 U4110 ( .A1(n3388), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3108) );
  AOI22_X1 U4111 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n3369), .B1(n3785), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3107) );
  AOI22_X1 U4112 ( .A1(n3733), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3106) );
  NAND4_X1 U4113 ( .A1(n3109), .A2(n3108), .A3(n3107), .A4(n3106), .ZN(n3110)
         );
  NOR2_X1 U4114 ( .A1(n3111), .A2(n3110), .ZN(n3803) );
  AOI22_X1 U4115 ( .A1(n3592), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3115) );
  AOI22_X1 U4116 ( .A1(n3337), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3114) );
  AOI22_X1 U4117 ( .A1(n3750), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4181), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3113) );
  AOI22_X1 U4118 ( .A1(n4146), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3112) );
  NAND4_X1 U4119 ( .A1(n3115), .A2(n3114), .A3(n3113), .A4(n3112), .ZN(n3121)
         );
  AOI22_X1 U4120 ( .A1(n3374), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3119) );
  AOI22_X1 U4121 ( .A1(n3354), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3118) );
  AOI22_X1 U4122 ( .A1(n3790), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3117) );
  AOI22_X1 U4123 ( .A1(n3733), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3116) );
  NAND4_X1 U4124 ( .A1(n3119), .A2(n3118), .A3(n3117), .A4(n3116), .ZN(n3120)
         );
  NOR2_X1 U4125 ( .A1(n3121), .A2(n3120), .ZN(n3804) );
  OR2_X1 U4126 ( .A1(n3803), .A2(n3804), .ZN(n3815) );
  AOI22_X1 U4127 ( .A1(n3337), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3125) );
  AOI22_X1 U4128 ( .A1(n3592), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3124) );
  AOI22_X1 U4129 ( .A1(n3354), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3123) );
  AOI22_X1 U4130 ( .A1(n4151), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3122) );
  NAND4_X1 U4131 ( .A1(n3125), .A2(n3124), .A3(n3123), .A4(n3122), .ZN(n3131)
         );
  AOI22_X1 U4132 ( .A1(n3733), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3129) );
  AOI22_X1 U4133 ( .A1(n3790), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4181), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3128) );
  AOI22_X1 U4134 ( .A1(n4146), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3127) );
  AOI22_X1 U4135 ( .A1(n3785), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3126) );
  NAND4_X1 U4136 ( .A1(n3129), .A2(n3128), .A3(n3127), .A4(n3126), .ZN(n3130)
         );
  NOR2_X1 U4137 ( .A1(n3131), .A2(n3130), .ZN(n3813) );
  OR2_X1 U4138 ( .A1(n3815), .A2(n3813), .ZN(n3822) );
  NOR2_X1 U4139 ( .A1(n3821), .A2(n3822), .ZN(n4123) );
  AOI22_X1 U4140 ( .A1(n3355), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3135) );
  AOI22_X1 U4141 ( .A1(n3790), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3134) );
  AOI22_X1 U4142 ( .A1(n3337), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3133) );
  AOI22_X1 U4143 ( .A1(n4146), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3132) );
  NAND4_X1 U4144 ( .A1(n3135), .A2(n3134), .A3(n3133), .A4(n3132), .ZN(n3141)
         );
  AOI22_X1 U4145 ( .A1(n3592), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3139) );
  AOI22_X1 U4146 ( .A1(n4151), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3138) );
  AOI22_X1 U4147 ( .A1(n3390), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3137) );
  AOI22_X1 U4148 ( .A1(n3015), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3136) );
  NAND4_X1 U4149 ( .A1(n3139), .A2(n3138), .A3(n3137), .A4(n3136), .ZN(n3140)
         );
  OR2_X1 U4150 ( .A1(n3141), .A2(n3140), .ZN(n4122) );
  XNOR2_X1 U4151 ( .A(n4123), .B(n4122), .ZN(n3195) );
  AOI22_X1 U4152 ( .A1(n3355), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3145) );
  AOI22_X1 U4153 ( .A1(n3368), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3245), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3144) );
  AOI22_X1 U4154 ( .A1(n3451), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3143) );
  AOI22_X1 U4155 ( .A1(n4182), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3185), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3142) );
  AOI22_X1 U4156 ( .A1(n4183), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3149) );
  AOI22_X1 U4157 ( .A1(n3250), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3389), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3147) );
  AOI22_X1 U4158 ( .A1(n3355), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3153) );
  AOI22_X1 U4159 ( .A1(n3368), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3245), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3152) );
  AOI22_X1 U4160 ( .A1(n3451), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U4161 ( .A1(n4182), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3185), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3150) );
  NAND4_X1 U4162 ( .A1(n3153), .A2(n3152), .A3(n3151), .A4(n3150), .ZN(n3159)
         );
  AOI22_X1 U4163 ( .A1(n3592), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3157) );
  AOI22_X1 U4164 ( .A1(n3250), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3389), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3156) );
  AOI22_X1 U4165 ( .A1(n3390), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3155) );
  AOI22_X1 U4166 ( .A1(n4183), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3154) );
  NAND4_X1 U4167 ( .A1(n3157), .A2(n3156), .A3(n3155), .A4(n3154), .ZN(n3158)
         );
  NAND2_X1 U4168 ( .A1(n3592), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3163) );
  NAND2_X1 U4169 ( .A1(n3374), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3162)
         );
  NAND2_X1 U4170 ( .A1(n3250), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3161) );
  NAND2_X1 U4171 ( .A1(n3389), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3160)
         );
  NAND2_X1 U4172 ( .A1(n3368), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3167)
         );
  NAND2_X1 U4173 ( .A1(n3451), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3166) );
  NAND2_X1 U4174 ( .A1(n3245), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3165) );
  NAND2_X1 U4175 ( .A1(n3395), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3164)
         );
  NAND2_X1 U4176 ( .A1(n3355), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3171) );
  NAND2_X1 U4177 ( .A1(n3367), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3170) );
  NAND2_X1 U4178 ( .A1(n4182), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3169)
         );
  NAND2_X1 U4179 ( .A1(n3185), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3168) );
  NAND2_X1 U4180 ( .A1(n3390), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3176) );
  NAND2_X1 U4181 ( .A1(n4183), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3175) );
  NAND2_X1 U4182 ( .A1(n3172), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3174) );
  NAND2_X1 U4183 ( .A1(n3272), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3173)
         );
  AOI22_X1 U4184 ( .A1(n3374), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3389), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3184) );
  AOI22_X1 U4185 ( .A1(n3355), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3183) );
  AOI22_X1 U4186 ( .A1(n3245), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3182) );
  AOI22_X1 U4187 ( .A1(n4183), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3181) );
  NAND4_X1 U4188 ( .A1(n3184), .A2(n3183), .A3(n3182), .A4(n3181), .ZN(n3191)
         );
  AOI22_X1 U4189 ( .A1(n3390), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3189) );
  AOI22_X1 U4190 ( .A1(n3592), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3188) );
  AOI22_X1 U4191 ( .A1(n4182), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3185), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3187) );
  AOI22_X1 U4192 ( .A1(n3451), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3368), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3186) );
  NAND4_X1 U4193 ( .A1(n3189), .A2(n3188), .A3(n3187), .A4(n3186), .ZN(n3190)
         );
  OR2_X2 U4194 ( .A1(n3191), .A2(n3190), .ZN(n3244) );
  NAND2_X1 U4195 ( .A1(n3257), .A2(n5338), .ZN(n4344) );
  NOR2_X2 U4196 ( .A1(n3192), .A2(n4124), .ZN(n3417) );
  INV_X1 U4197 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4007) );
  OAI21_X1 U4198 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4007), .A(n3524), .ZN(
        n3193) );
  AOI21_X1 U4199 ( .B1(n3417), .B2(EAX_REG_26__SCAN_IN), .A(n3193), .ZN(n3194)
         );
  OAI21_X1 U4200 ( .B1(n3195), .B2(n4173), .A(n3194), .ZN(n3201) );
  INV_X1 U4201 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3197) );
  INV_X1 U4202 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5588) );
  INV_X1 U4203 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3199) );
  XNOR2_X1 U4204 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .B(n3897), .ZN(n5561)
         );
  NAND2_X1 U4205 ( .A1(n5561), .A2(n4202), .ZN(n3200) );
  NAND2_X1 U4206 ( .A1(n3201), .A2(n3200), .ZN(n3832) );
  NAND2_X1 U4207 ( .A1(n3283), .A2(n4620), .ZN(n4237) );
  INV_X1 U4208 ( .A(n4237), .ZN(n3203) );
  NAND2_X1 U4209 ( .A1(n3592), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3207) );
  NAND2_X1 U4210 ( .A1(n3374), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3206)
         );
  NAND2_X1 U4211 ( .A1(n3250), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3205) );
  NAND2_X1 U4212 ( .A1(n3389), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3204)
         );
  NAND2_X1 U4213 ( .A1(n3368), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3211)
         );
  NAND2_X1 U4214 ( .A1(n3451), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3210) );
  NAND2_X1 U4215 ( .A1(n3245), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3209) );
  NAND2_X1 U4216 ( .A1(n3395), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3208)
         );
  NAND2_X1 U4217 ( .A1(n3355), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3215) );
  NAND2_X1 U4218 ( .A1(n3367), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3214) );
  NAND2_X1 U4219 ( .A1(n4182), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3213)
         );
  NAND2_X1 U4220 ( .A1(n3185), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3212) );
  NAND2_X1 U4221 ( .A1(n3390), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3219) );
  NAND2_X1 U4222 ( .A1(n4183), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3218) );
  NAND2_X1 U4223 ( .A1(n3172), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3217) );
  NAND2_X1 U4224 ( .A1(n3272), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3216)
         );
  INV_X1 U4225 ( .A(n4511), .ZN(n4501) );
  NAND2_X1 U4226 ( .A1(n3451), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3227) );
  NAND2_X1 U4227 ( .A1(n3368), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3226)
         );
  NAND2_X1 U4228 ( .A1(n3245), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3225) );
  NAND2_X1 U4229 ( .A1(n3185), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3224) );
  NAND2_X1 U4230 ( .A1(n3250), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3231) );
  NAND2_X1 U4231 ( .A1(n3592), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3230) );
  NAND2_X1 U4232 ( .A1(n4183), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3229) );
  NAND2_X1 U4233 ( .A1(n3389), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3228)
         );
  NAND2_X1 U4234 ( .A1(n3355), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3235) );
  NAND2_X1 U4235 ( .A1(n3367), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3234) );
  NAND2_X1 U4236 ( .A1(n3395), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3233)
         );
  NAND2_X1 U4237 ( .A1(n4182), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3232)
         );
  NAND2_X1 U4238 ( .A1(n3390), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3239) );
  NAND2_X1 U4239 ( .A1(n3374), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3238)
         );
  NAND2_X1 U4240 ( .A1(n3272), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3237)
         );
  NAND2_X1 U4241 ( .A1(n3172), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3236) );
  AOI22_X1 U4242 ( .A1(n3355), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3249) );
  AOI22_X1 U4243 ( .A1(n3368), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3245), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3248) );
  AOI22_X1 U4244 ( .A1(n3451), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3395), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3247) );
  NAND4_X1 U4245 ( .A1(n3249), .A2(n3248), .A3(n3247), .A4(n3246), .ZN(n3256)
         );
  AOI22_X1 U4246 ( .A1(n3592), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3254) );
  AOI22_X1 U4247 ( .A1(n3250), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3389), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4248 ( .A1(n3390), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U4249 ( .A1(n4183), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3251) );
  NAND4_X1 U4250 ( .A1(n3254), .A2(n3253), .A3(n3252), .A4(n3251), .ZN(n3255)
         );
  OR2_X2 U4251 ( .A1(n3256), .A2(n3255), .ZN(n4019) );
  NAND2_X1 U4252 ( .A1(n3290), .A2(n4019), .ZN(n3315) );
  OAI21_X1 U4253 ( .B1(n3258), .B2(n3257), .A(n3315), .ZN(n3299) );
  INV_X1 U4254 ( .A(n3299), .ZN(n3892) );
  NAND2_X1 U4255 ( .A1(n3259), .A2(n3892), .ZN(n3312) );
  NAND2_X1 U4256 ( .A1(n3592), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3263) );
  NAND2_X1 U4257 ( .A1(n3374), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3262)
         );
  NAND2_X1 U4258 ( .A1(n3250), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3261) );
  NAND2_X1 U4259 ( .A1(n3389), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3260)
         );
  NAND2_X1 U4260 ( .A1(n3368), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3267)
         );
  NAND2_X1 U4261 ( .A1(n3451), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3266) );
  NAND2_X1 U4262 ( .A1(n3245), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3265) );
  NAND2_X1 U4263 ( .A1(n3395), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3264)
         );
  NAND2_X1 U4264 ( .A1(n3355), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3271) );
  NAND2_X1 U4265 ( .A1(n3367), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3270) );
  NAND2_X1 U4266 ( .A1(n4182), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3269)
         );
  NAND2_X1 U4267 ( .A1(n3185), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3268) );
  NAND2_X1 U4268 ( .A1(n3390), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3276) );
  NAND2_X1 U4269 ( .A1(n4183), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3275) );
  NAND2_X1 U4270 ( .A1(n3172), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3274) );
  NAND2_X1 U4271 ( .A1(n3272), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3273)
         );
  NAND2_X1 U4272 ( .A1(n3312), .A2(n4580), .ZN(n3288) );
  INV_X2 U4273 ( .A(n4371), .ZN(n4615) );
  NAND2_X1 U4274 ( .A1(n3314), .A2(n4312), .ZN(n3281) );
  NAND2_X1 U4275 ( .A1(n4620), .A2(n5338), .ZN(n4111) );
  NAND2_X1 U4276 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6489) );
  OAI21_X1 U4277 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6489), .ZN(n3995) );
  NAND2_X1 U4278 ( .A1(n4615), .A2(n3995), .ZN(n3294) );
  NAND2_X1 U4279 ( .A1(n3294), .A2(n3282), .ZN(n3287) );
  AND2_X1 U4280 ( .A1(n3283), .A2(n3192), .ZN(n3286) );
  OR2_X1 U4281 ( .A1(n3290), .A2(n3284), .ZN(n3285) );
  NAND4_X1 U4282 ( .A1(n3288), .A2(n3321), .A3(n3287), .A4(n4110), .ZN(n3289)
         );
  NAND2_X1 U4283 ( .A1(n3289), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3292) );
  NAND2_X1 U4284 ( .A1(n3290), .A2(n3877), .ZN(n3291) );
  NAND2_X1 U4285 ( .A1(n3325), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3304) );
  NAND2_X1 U4286 ( .A1(n3030), .A2(n5958), .ZN(n4373) );
  AND2_X1 U4287 ( .A1(n3296), .A2(n3192), .ZN(n5339) );
  NAND2_X1 U4288 ( .A1(n4346), .A2(n6474), .ZN(n6586) );
  INV_X1 U4289 ( .A(n6586), .ZN(n3329) );
  XNOR2_X1 U4290 ( .A(n6430), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5205)
         );
  NAND2_X1 U4291 ( .A1(n3329), .A2(n5205), .ZN(n3302) );
  INV_X1 U4292 ( .A(n6470), .ZN(n3300) );
  NAND2_X1 U4293 ( .A1(n3300), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3301) );
  INV_X1 U4294 ( .A(n3305), .ZN(n3308) );
  INV_X1 U4295 ( .A(n3306), .ZN(n3307) );
  OAI21_X1 U4296 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n3308), .A(n3307), 
        .ZN(n3309) );
  AND2_X2 U4297 ( .A1(n3323), .A2(n3309), .ZN(n3352) );
  MUX2_X1 U4298 ( .A(n6470), .B(n6586), .S(n6430), .Z(n3310) );
  NAND2_X1 U4299 ( .A1(n4082), .A2(n3005), .ZN(n3311) );
  NAND2_X1 U4300 ( .A1(n3312), .A2(n3311), .ZN(n3313) );
  MUX2_X1 U4301 ( .A(n4511), .B(n3313), .S(n4580), .Z(n4245) );
  NAND2_X1 U4302 ( .A1(n4346), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6478) );
  AOI21_X1 U4303 ( .B1(n3315), .B2(n3314), .A(n6478), .ZN(n3320) );
  AND3_X1 U4304 ( .A1(n4586), .A2(n4580), .A3(n4511), .ZN(n3316) );
  NAND2_X1 U4305 ( .A1(n3257), .A2(n3316), .ZN(n4529) );
  NAND2_X1 U4306 ( .A1(n3290), .A2(n3284), .ZN(n3317) );
  NAND2_X1 U4307 ( .A1(n3317), .A2(n4019), .ZN(n3318) );
  OAI21_X1 U4308 ( .B1(n4240), .B2(n3318), .A(n4371), .ZN(n3319) );
  NAND2_X2 U4309 ( .A1(n3385), .A2(n3384), .ZN(n3387) );
  NAND2_X1 U4310 ( .A1(n3352), .A2(n3387), .ZN(n3324) );
  NAND2_X1 U4311 ( .A1(n3324), .A2(n3000), .ZN(n3335) );
  INV_X1 U4312 ( .A(n3335), .ZN(n3333) );
  AND2_X1 U4313 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3326) );
  NAND2_X1 U4314 ( .A1(n3326), .A2(n6441), .ZN(n6314) );
  INV_X1 U4315 ( .A(n3326), .ZN(n3327) );
  NAND2_X1 U4316 ( .A1(n3327), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3328) );
  NAND2_X1 U4317 ( .A1(n6314), .A2(n3328), .ZN(n4703) );
  NAND2_X1 U4318 ( .A1(n3329), .A2(n4703), .ZN(n3330) );
  OAI21_X1 U4319 ( .B1(n6470), .B2(n6441), .A(n3330), .ZN(n3331) );
  INV_X1 U4320 ( .A(n3334), .ZN(n3332) );
  NAND2_X1 U4321 ( .A1(n3335), .A2(n3334), .ZN(n3336) );
  AOI22_X1 U4322 ( .A1(n3733), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3341) );
  AOI22_X1 U4323 ( .A1(n3790), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4324 ( .A1(n3337), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4325 ( .A1(n4182), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3338) );
  NAND4_X1 U4326 ( .A1(n3341), .A2(n3340), .A3(n3339), .A4(n3338), .ZN(n3347)
         );
  AOI22_X1 U4327 ( .A1(n4188), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3345) );
  AOI22_X1 U4328 ( .A1(n4151), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3344) );
  AOI22_X1 U4329 ( .A1(n3390), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3343) );
  AOI22_X1 U4330 ( .A1(n4183), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3342) );
  NAND4_X1 U4331 ( .A1(n3345), .A2(n3344), .A3(n3343), .A4(n3342), .ZN(n3346)
         );
  OAI22_X2 U4332 ( .A1(n4407), .A2(STATE2_REG_0__SCAN_IN), .B1(n4034), .B2(
        n3450), .ZN(n3351) );
  INV_X1 U4333 ( .A(n3449), .ZN(n3349) );
  AOI22_X1 U4334 ( .A1(n3349), .A2(n3348), .B1(n3877), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3350) );
  INV_X1 U4335 ( .A(n3352), .ZN(n3353) );
  XNOR2_X2 U4336 ( .A(n3387), .B(n3353), .ZN(n4342) );
  AOI22_X1 U4337 ( .A1(n3354), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4338 ( .A1(n3337), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3790), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4339 ( .A1(n3390), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3357) );
  AOI22_X1 U4340 ( .A1(n3733), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3356) );
  NAND4_X1 U4341 ( .A1(n3359), .A2(n3358), .A3(n3357), .A4(n3356), .ZN(n3365)
         );
  AOI22_X1 U4342 ( .A1(n3388), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3363) );
  AOI22_X1 U4343 ( .A1(n3785), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4344 ( .A1(n4188), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U4345 ( .A1(n4182), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3360) );
  NAND4_X1 U4346 ( .A1(n3363), .A2(n3362), .A3(n3361), .A4(n3360), .ZN(n3364)
         );
  OR2_X1 U4347 ( .A1(n3450), .A2(n3383), .ZN(n3366) );
  OAI21_X2 U4348 ( .B1(n4342), .B2(STATE2_REG_0__SCAN_IN), .A(n3366), .ZN(
        n3415) );
  NAND2_X1 U4349 ( .A1(n3877), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4350 ( .A1(n3733), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4351 ( .A1(n3790), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4352 ( .A1(n3337), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3371) );
  AOI22_X1 U4353 ( .A1(n4146), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3370) );
  NAND4_X1 U4354 ( .A1(n3373), .A2(n3372), .A3(n3371), .A4(n3370), .ZN(n3380)
         );
  AOI22_X1 U4355 ( .A1(n4188), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4356 ( .A1(n4151), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4357 ( .A1(n3390), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4358 ( .A1(n3015), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3375) );
  NAND4_X1 U4359 ( .A1(n3378), .A2(n3377), .A3(n3376), .A4(n3375), .ZN(n3379)
         );
  OR2_X1 U4360 ( .A1(n3450), .A2(n4085), .ZN(n3381) );
  OAI211_X1 U4361 ( .C1(n3449), .C2(n3383), .A(n3382), .B(n3381), .ZN(n3414)
         );
  AOI22_X1 U4362 ( .A1(n4188), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4363 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n3790), .B1(n4183), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4364 ( .A1(n4151), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3392) );
  AOI22_X1 U4365 ( .A1(n3390), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3391) );
  NAND4_X1 U4366 ( .A1(n3394), .A2(n3393), .A3(n3392), .A4(n3391), .ZN(n3401)
         );
  AOI22_X1 U4367 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n3337), .B1(n3369), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4368 ( .A1(n3354), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4369 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n3733), .B1(n4145), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3397) );
  AOI22_X1 U4370 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n3785), .B1(n4182), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3396) );
  NAND4_X1 U4371 ( .A1(n3399), .A2(n3398), .A3(n3397), .A4(n3396), .ZN(n3400)
         );
  XNOR2_X1 U4372 ( .A(n3547), .B(n4022), .ZN(n3403) );
  INV_X1 U4373 ( .A(n3450), .ZN(n3402) );
  NAND2_X1 U4374 ( .A1(n3403), .A2(n3402), .ZN(n3422) );
  INV_X1 U4375 ( .A(n4022), .ZN(n3406) );
  NAND2_X1 U4376 ( .A1(n3877), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3405) );
  AOI21_X1 U4377 ( .B1(n3005), .B2(n4085), .A(n6474), .ZN(n3404) );
  OR2_X1 U4378 ( .A1(n3450), .A2(n3547), .ZN(n3408) );
  NAND2_X1 U4379 ( .A1(n3415), .A2(n3414), .ZN(n3409) );
  NAND2_X1 U4380 ( .A1(n3410), .A2(n3409), .ZN(n3411) );
  NAND2_X2 U4381 ( .A1(n3412), .A2(n3411), .ZN(n3473) );
  NAND2_X1 U4382 ( .A1(n4481), .A2(n3674), .ZN(n3421) );
  INV_X1 U4383 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n4573) );
  AOI22_X1 U4384 ( .A1(n4207), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n4573), .ZN(n3419) );
  AND2_X1 U4385 ( .A1(n5339), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3435) );
  NAND2_X1 U4386 ( .A1(n3435), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3418) );
  AND2_X1 U4387 ( .A1(n3419), .A2(n3418), .ZN(n3420) );
  NAND2_X1 U4388 ( .A1(n3421), .A2(n3420), .ZN(n4380) );
  INV_X1 U4389 ( .A(n3422), .ZN(n3423) );
  NAND2_X2 U4390 ( .A1(n3426), .A2(n3425), .ZN(n4853) );
  INV_X1 U4391 ( .A(n3202), .ZN(n3427) );
  AOI21_X1 U4392 ( .B1(n4853), .B2(n3427), .A(n4573), .ZN(n4369) );
  INV_X1 U4393 ( .A(n3674), .ZN(n3663) );
  OR2_X1 U4394 ( .A1(n3428), .A2(n3663), .ZN(n3432) );
  AOI22_X1 U4395 ( .A1(n4207), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n4573), .ZN(n3430) );
  NAND2_X1 U4396 ( .A1(n3435), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3429) );
  AND2_X1 U4397 ( .A1(n3430), .A2(n3429), .ZN(n3431) );
  NAND2_X1 U4398 ( .A1(n3432), .A2(n3431), .ZN(n4368) );
  NAND2_X1 U4399 ( .A1(n4369), .A2(n4368), .ZN(n4367) );
  INV_X1 U4400 ( .A(n4368), .ZN(n3433) );
  NAND2_X1 U4401 ( .A1(n3433), .A2(n4202), .ZN(n3434) );
  NAND2_X1 U4402 ( .A1(n4367), .A2(n3434), .ZN(n4379) );
  NAND2_X1 U4403 ( .A1(n4380), .A2(n4379), .ZN(n4382) );
  INV_X1 U4404 ( .A(n3435), .ZN(n3497) );
  OAI21_X1 U4405 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3436), .ZN(n6142) );
  AOI22_X1 U4406 ( .A1(n6142), .A2(n4202), .B1(n4206), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3438) );
  NAND2_X1 U4407 ( .A1(n4207), .A2(EAX_REG_2__SCAN_IN), .ZN(n3437) );
  OAI211_X1 U4408 ( .C1(n3497), .C2(n5336), .A(n3438), .B(n3437), .ZN(n4385)
         );
  NAND2_X1 U4409 ( .A1(n4384), .A2(n4385), .ZN(n3443) );
  INV_X1 U4410 ( .A(n3439), .ZN(n3441) );
  INV_X1 U4411 ( .A(n4382), .ZN(n3440) );
  NAND2_X1 U4412 ( .A1(n3441), .A2(n3440), .ZN(n3442) );
  NAND2_X1 U4413 ( .A1(n3443), .A2(n3442), .ZN(n4383) );
  NAND2_X1 U4414 ( .A1(n3325), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3448) );
  NOR3_X1 U4415 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6441), .A3(n6437), 
        .ZN(n6284) );
  NAND2_X1 U4416 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6284), .ZN(n6282) );
  NAND2_X1 U4417 ( .A1(n6572), .A2(n6282), .ZN(n3445) );
  NAND3_X1 U4418 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4785) );
  INV_X1 U4419 ( .A(n4785), .ZN(n6378) );
  NAND2_X1 U4420 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6378), .ZN(n6364) );
  NAND2_X1 U4421 ( .A1(n3445), .A2(n6364), .ZN(n5128) );
  OAI22_X1 U4422 ( .A1(n6586), .A2(n5128), .B1(n6470), .B2(n6572), .ZN(n3446)
         );
  INV_X1 U4423 ( .A(n3446), .ZN(n3447) );
  NAND2_X1 U4424 ( .A1(n4390), .A2(n6474), .ZN(n3466) );
  AOI22_X1 U4425 ( .A1(n3733), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4426 ( .A1(n3790), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4427 ( .A1(n3337), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4428 ( .A1(n4146), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3452) );
  NAND4_X1 U4429 ( .A1(n3455), .A2(n3454), .A3(n3453), .A4(n3452), .ZN(n3461)
         );
  AOI22_X1 U4430 ( .A1(n4188), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3459) );
  AOI22_X1 U4431 ( .A1(n4151), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3458) );
  AOI22_X1 U4432 ( .A1(n3750), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3457) );
  AOI22_X1 U4433 ( .A1(n4183), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3456) );
  NAND4_X1 U4434 ( .A1(n3459), .A2(n3458), .A3(n3457), .A4(n3456), .ZN(n3460)
         );
  INV_X1 U4435 ( .A(n4044), .ZN(n3463) );
  INV_X1 U4436 ( .A(n3877), .ZN(n3865) );
  INV_X1 U4437 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3462) );
  OAI22_X1 U4438 ( .A1(n3882), .A2(n3463), .B1(n3865), .B2(n3462), .ZN(n3464)
         );
  INV_X1 U4439 ( .A(n3464), .ZN(n3465) );
  XNOR2_X2 U4440 ( .A(n3473), .B(n4479), .ZN(n4042) );
  NAND2_X1 U4441 ( .A1(n4042), .A2(n3674), .ZN(n3472) );
  OAI21_X1 U4442 ( .B1(n3467), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n3494), 
        .ZN(n5344) );
  AOI22_X1 U4443 ( .A1(n5344), .A2(n4202), .B1(n4206), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3469) );
  NAND2_X1 U4444 ( .A1(n3417), .A2(EAX_REG_3__SCAN_IN), .ZN(n3468) );
  OAI211_X1 U4445 ( .C1(n3497), .C2(n4406), .A(n3469), .B(n3468), .ZN(n3470)
         );
  INV_X1 U4446 ( .A(n3470), .ZN(n3471) );
  NAND2_X1 U4447 ( .A1(n4383), .A2(n4389), .ZN(n4388) );
  INV_X1 U4448 ( .A(n4388), .ZN(n3502) );
  INV_X1 U4449 ( .A(n3473), .ZN(n3474) );
  NAND2_X1 U4450 ( .A1(n3474), .A2(n4479), .ZN(n3490) );
  INV_X1 U4451 ( .A(n3490), .ZN(n3488) );
  AOI22_X1 U4452 ( .A1(n3733), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4453 ( .A1(n3388), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3477) );
  AOI22_X1 U4454 ( .A1(n4188), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3476) );
  AOI22_X1 U4455 ( .A1(n3785), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3475) );
  NAND4_X1 U4456 ( .A1(n3478), .A2(n3477), .A3(n3476), .A4(n3475), .ZN(n3484)
         );
  AOI22_X1 U4457 ( .A1(n3750), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4458 ( .A1(n3337), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3481) );
  AOI22_X1 U4459 ( .A1(n4183), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3480) );
  AOI22_X1 U4460 ( .A1(n3790), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3479) );
  NAND4_X1 U4461 ( .A1(n3482), .A2(n3481), .A3(n3480), .A4(n3479), .ZN(n3483)
         );
  NAND2_X1 U4462 ( .A1(n3877), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3485) );
  INV_X1 U4463 ( .A(n3489), .ZN(n3487) );
  NAND2_X1 U4464 ( .A1(n3490), .A2(n3489), .ZN(n3491) );
  INV_X1 U4465 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3493) );
  INV_X1 U4466 ( .A(n3520), .ZN(n3492) );
  AOI21_X1 U4467 ( .B1(n3494), .B2(n3493), .A(n3492), .ZN(n6051) );
  INV_X1 U4468 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4328) );
  NAND2_X1 U4469 ( .A1(n4573), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3496)
         );
  NAND2_X1 U4470 ( .A1(n3417), .A2(EAX_REG_4__SCAN_IN), .ZN(n3495) );
  OAI211_X1 U4471 ( .C1(n3497), .C2(n4328), .A(n3496), .B(n3495), .ZN(n3498)
         );
  NAND2_X1 U4472 ( .A1(n3498), .A2(n3524), .ZN(n3499) );
  OAI21_X1 U4473 ( .B1(n6051), .B2(n3524), .A(n3499), .ZN(n3500) );
  AOI22_X1 U4474 ( .A1(n3733), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3506) );
  AOI22_X1 U4475 ( .A1(n3790), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3505) );
  AOI22_X1 U4476 ( .A1(n3337), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3504) );
  AOI22_X1 U4477 ( .A1(n4146), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3503) );
  NAND4_X1 U4478 ( .A1(n3506), .A2(n3505), .A3(n3504), .A4(n3503), .ZN(n3512)
         );
  AOI22_X1 U4479 ( .A1(n4188), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3510) );
  AOI22_X1 U4480 ( .A1(n4151), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3509) );
  AOI22_X1 U4481 ( .A1(n3750), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4181), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3508) );
  AOI22_X1 U4482 ( .A1(n4183), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3507) );
  NAND4_X1 U4483 ( .A1(n3510), .A2(n3509), .A3(n3508), .A4(n3507), .ZN(n3511)
         );
  INV_X1 U4484 ( .A(n4056), .ZN(n3513) );
  NAND2_X1 U4485 ( .A1(n3877), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3514) );
  NAND2_X1 U4486 ( .A1(n3009), .A2(n3516), .ZN(n3542) );
  INV_X1 U4487 ( .A(n3516), .ZN(n3517) );
  NAND2_X1 U4488 ( .A1(n3518), .A2(n3517), .ZN(n3519) );
  AOI21_X1 U4489 ( .B1(n3520), .B2(n6038), .A(n3525), .ZN(n4558) );
  NAND2_X1 U4490 ( .A1(n3417), .A2(EAX_REG_5__SCAN_IN), .ZN(n3522) );
  NAND2_X1 U4491 ( .A1(n4206), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3521)
         );
  OAI211_X1 U4492 ( .C1(n4558), .C2(n3524), .A(n3522), .B(n3521), .ZN(n3523)
         );
  OAI21_X1 U4493 ( .B1(n3525), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n3549), 
        .ZN(n3526) );
  INV_X1 U4494 ( .A(n3526), .ZN(n6032) );
  AOI22_X1 U4495 ( .A1(n4188), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3530) );
  AOI22_X1 U4496 ( .A1(n3750), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U4497 ( .A1(n3337), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3528) );
  AOI22_X1 U4498 ( .A1(n3790), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3527) );
  NAND4_X1 U4499 ( .A1(n3530), .A2(n3529), .A3(n3528), .A4(n3527), .ZN(n3536)
         );
  AOI22_X1 U4500 ( .A1(n3733), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3534) );
  AOI22_X1 U4501 ( .A1(n3388), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4502 ( .A1(n4181), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3532) );
  AOI22_X1 U4503 ( .A1(n3785), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3531) );
  NAND4_X1 U4504 ( .A1(n3534), .A2(n3533), .A3(n3532), .A4(n3531), .ZN(n3535)
         );
  INV_X1 U4505 ( .A(n4073), .ZN(n3537) );
  NAND2_X1 U4506 ( .A1(n3877), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3538) );
  NAND2_X1 U4507 ( .A1(n3542), .A2(n3543), .ZN(n4063) );
  NAND2_X1 U4508 ( .A1(n4063), .A2(n3674), .ZN(n3541) );
  AOI22_X1 U4509 ( .A1(n4207), .A2(EAX_REG_6__SCAN_IN), .B1(n4206), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3540) );
  OAI211_X1 U4510 ( .C1(n3524), .C2(n6032), .A(n3541), .B(n3540), .ZN(n4453)
         );
  NAND2_X1 U4511 ( .A1(n4450), .A2(n4453), .ZN(n4452) );
  INV_X1 U4512 ( .A(n4452), .ZN(n3554) );
  INV_X1 U4513 ( .A(n3542), .ZN(n3545) );
  INV_X1 U4514 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3546) );
  OAI22_X1 U4515 ( .A1(n3882), .A2(n3547), .B1(n3865), .B2(n3546), .ZN(n3548)
         );
  NAND2_X1 U4516 ( .A1(n4071), .A2(n3674), .ZN(n3553) );
  AOI21_X1 U4517 ( .B1(n3549), .B2(n6023), .A(n3555), .ZN(n5085) );
  AOI22_X1 U4518 ( .A1(n4207), .A2(EAX_REG_7__SCAN_IN), .B1(n4206), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3550) );
  OAI21_X1 U4519 ( .B1(n5085), .B2(n3524), .A(n3550), .ZN(n3551) );
  NAND2_X1 U4520 ( .A1(n3554), .A2(n4911), .ZN(n4912) );
  XOR2_X1 U4521 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3555), .Z(n6013) );
  INV_X1 U4522 ( .A(n6013), .ZN(n5098) );
  AOI22_X1 U4523 ( .A1(n3388), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4524 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n3337), .B1(n3785), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3558) );
  AOI22_X1 U4525 ( .A1(n4188), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4526 ( .A1(n4183), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3556) );
  NAND4_X1 U4527 ( .A1(n3559), .A2(n3558), .A3(n3557), .A4(n3556), .ZN(n3565)
         );
  AOI22_X1 U4528 ( .A1(n3750), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4529 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n3790), .B1(n3369), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4530 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n3354), .B1(n4181), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4531 ( .A1(n3733), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3560) );
  NAND4_X1 U4532 ( .A1(n3563), .A2(n3562), .A3(n3561), .A4(n3560), .ZN(n3564)
         );
  OAI21_X1 U4533 ( .B1(n3565), .B2(n3564), .A(n3674), .ZN(n3568) );
  NAND2_X1 U4534 ( .A1(n3417), .A2(EAX_REG_8__SCAN_IN), .ZN(n3567) );
  NAND2_X1 U4535 ( .A1(n4206), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3566)
         );
  NAND3_X1 U4536 ( .A1(n3568), .A2(n3567), .A3(n3566), .ZN(n3569) );
  AOI21_X1 U4537 ( .B1(n5098), .B2(n4202), .A(n3569), .ZN(n5092) );
  XNOR2_X1 U4538 ( .A(n3572), .B(n5107), .ZN(n5115) );
  AOI22_X1 U4539 ( .A1(n3388), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4540 ( .A1(n3337), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4541 ( .A1(n4188), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4181), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4542 ( .A1(n4146), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3573) );
  NAND4_X1 U4543 ( .A1(n3576), .A2(n3575), .A3(n3574), .A4(n3573), .ZN(n3582)
         );
  AOI22_X1 U4544 ( .A1(n3750), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4151), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4545 ( .A1(n3733), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4546 ( .A1(n3790), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3578) );
  AOI22_X1 U4547 ( .A1(n4183), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3577) );
  NAND4_X1 U4548 ( .A1(n3580), .A2(n3579), .A3(n3578), .A4(n3577), .ZN(n3581)
         );
  OAI21_X1 U4549 ( .B1(n3582), .B2(n3581), .A(n3674), .ZN(n3585) );
  NAND2_X1 U4550 ( .A1(n3417), .A2(EAX_REG_9__SCAN_IN), .ZN(n3584) );
  NAND2_X1 U4551 ( .A1(n4206), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3583)
         );
  NAND3_X1 U4552 ( .A1(n3585), .A2(n3584), .A3(n3583), .ZN(n3586) );
  AOI21_X1 U4553 ( .B1(n5115), .B2(n4202), .A(n3586), .ZN(n5053) );
  XOR2_X1 U4554 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3587), .Z(n6000) );
  AOI22_X1 U4555 ( .A1(n4151), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4556 ( .A1(n3733), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3590) );
  AOI22_X1 U4557 ( .A1(n3388), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4181), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3589) );
  AOI22_X1 U4558 ( .A1(n4183), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3588) );
  NAND4_X1 U4559 ( .A1(n3591), .A2(n3590), .A3(n3589), .A4(n3588), .ZN(n3598)
         );
  AOI22_X1 U4560 ( .A1(n4188), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4561 ( .A1(n3337), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4562 ( .A1(n3354), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4563 ( .A1(n3790), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3593) );
  NAND4_X1 U4564 ( .A1(n3596), .A2(n3595), .A3(n3594), .A4(n3593), .ZN(n3597)
         );
  OR2_X1 U4565 ( .A1(n3598), .A2(n3597), .ZN(n3599) );
  AOI22_X1 U4566 ( .A1(n3674), .A2(n3599), .B1(n4206), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3601) );
  NAND2_X1 U4567 ( .A1(n3417), .A2(EAX_REG_10__SCAN_IN), .ZN(n3600) );
  OAI211_X1 U4568 ( .C1(n6000), .C2(n3524), .A(n3601), .B(n3600), .ZN(n5111)
         );
  AOI22_X1 U4569 ( .A1(n4188), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3605) );
  AOI22_X1 U4570 ( .A1(n3354), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3015), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3604) );
  AOI22_X1 U4571 ( .A1(n3337), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3603) );
  AOI22_X1 U4572 ( .A1(n3750), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4181), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3602) );
  NAND4_X1 U4573 ( .A1(n3605), .A2(n3604), .A3(n3603), .A4(n3602), .ZN(n3611)
         );
  AOI22_X1 U4574 ( .A1(n4151), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4575 ( .A1(n3790), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3608) );
  AOI22_X1 U4576 ( .A1(n3733), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3607) );
  AOI22_X1 U4577 ( .A1(n4146), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3606) );
  NAND4_X1 U4578 ( .A1(n3609), .A2(n3608), .A3(n3607), .A4(n3606), .ZN(n3610)
         );
  NOR2_X1 U4579 ( .A1(n3611), .A2(n3610), .ZN(n3615) );
  XNOR2_X1 U4580 ( .A(n3612), .B(n5170), .ZN(n5259) );
  NAND2_X1 U4581 ( .A1(n5259), .A2(n4202), .ZN(n3614) );
  AOI22_X1 U4582 ( .A1(n4207), .A2(EAX_REG_11__SCAN_IN), .B1(n4206), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3613) );
  OAI211_X1 U4583 ( .C1(n3615), .C2(n3663), .A(n3614), .B(n3613), .ZN(n5122)
         );
  XOR2_X1 U4584 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3616), .Z(n5306) );
  AOI22_X1 U4585 ( .A1(n4151), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4586 ( .A1(n3354), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4587 ( .A1(n3785), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4588 ( .A1(n3790), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3617) );
  NAND4_X1 U4589 ( .A1(n3620), .A2(n3619), .A3(n3618), .A4(n3617), .ZN(n3626)
         );
  AOI22_X1 U4590 ( .A1(n4188), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4591 ( .A1(n3750), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4181), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4592 ( .A1(n3337), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4593 ( .A1(n3733), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3621) );
  NAND4_X1 U4594 ( .A1(n3624), .A2(n3623), .A3(n3622), .A4(n3621), .ZN(n3625)
         );
  OR2_X1 U4595 ( .A1(n3626), .A2(n3625), .ZN(n3627) );
  AOI22_X1 U4596 ( .A1(n3674), .A2(n3627), .B1(n4206), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3629) );
  NAND2_X1 U4597 ( .A1(n3417), .A2(EAX_REG_12__SCAN_IN), .ZN(n3628) );
  OAI211_X1 U4598 ( .C1(n5306), .C2(n3524), .A(n3629), .B(n3628), .ZN(n5184)
         );
  XNOR2_X1 U4599 ( .A(n3630), .B(n3631), .ZN(n5314) );
  NAND2_X1 U4600 ( .A1(n5314), .A2(n4202), .ZN(n3635) );
  INV_X1 U4601 ( .A(n4206), .ZN(n3632) );
  NOR2_X1 U4602 ( .A1(n3632), .A2(n3631), .ZN(n3633) );
  AOI21_X1 U4603 ( .B1(n3417), .B2(EAX_REG_13__SCAN_IN), .A(n3633), .ZN(n3634)
         );
  NAND2_X1 U4604 ( .A1(n3635), .A2(n3634), .ZN(n3647) );
  AOI22_X1 U4605 ( .A1(n3337), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4606 ( .A1(n4151), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3638) );
  AOI22_X1 U4607 ( .A1(n3388), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4608 ( .A1(n3785), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4181), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3636) );
  NAND4_X1 U4609 ( .A1(n3639), .A2(n3638), .A3(n3637), .A4(n3636), .ZN(n3645)
         );
  AOI22_X1 U4610 ( .A1(n3733), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4611 ( .A1(n4188), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4612 ( .A1(n3015), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4613 ( .A1(n3790), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3640) );
  NAND4_X1 U4614 ( .A1(n3643), .A2(n3642), .A3(n3641), .A4(n3640), .ZN(n3644)
         );
  OR2_X1 U4615 ( .A1(n3645), .A2(n3644), .ZN(n3646) );
  AND2_X1 U4616 ( .A1(n3674), .A2(n3646), .ZN(n5267) );
  NAND2_X1 U4617 ( .A1(n5264), .A2(n5267), .ZN(n5265) );
  INV_X1 U4618 ( .A(n3647), .ZN(n3648) );
  NAND2_X1 U4619 ( .A1(n5265), .A2(n5319), .ZN(n3664) );
  AOI22_X1 U4620 ( .A1(n4188), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3652) );
  AOI22_X1 U4621 ( .A1(n3733), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3651) );
  AOI22_X1 U4622 ( .A1(n3337), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3650) );
  AOI22_X1 U4623 ( .A1(n3750), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3649) );
  NAND4_X1 U4624 ( .A1(n3652), .A2(n3651), .A3(n3650), .A4(n3649), .ZN(n3658)
         );
  AOI22_X1 U4625 ( .A1(n3388), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4626 ( .A1(n3790), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3655) );
  AOI22_X1 U4627 ( .A1(n4183), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4181), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4628 ( .A1(n4146), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3653) );
  NAND4_X1 U4629 ( .A1(n3656), .A2(n3655), .A3(n3654), .A4(n3653), .ZN(n3657)
         );
  NOR2_X1 U4630 ( .A1(n3658), .A2(n3657), .ZN(n3662) );
  XNOR2_X1 U4631 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3659), .ZN(n5637)
         );
  AOI22_X1 U4632 ( .A1(n4202), .A2(n5637), .B1(n4206), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3661) );
  NAND2_X1 U4633 ( .A1(n4207), .A2(EAX_REG_14__SCAN_IN), .ZN(n3660) );
  OAI211_X1 U4634 ( .C1(n3663), .C2(n3662), .A(n3661), .B(n3660), .ZN(n5320)
         );
  XNOR2_X1 U4635 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3665), .ZN(n5418)
         );
  INV_X1 U4636 ( .A(n5418), .ZN(n5627) );
  AOI22_X1 U4637 ( .A1(n3790), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4638 ( .A1(n3337), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4639 ( .A1(n4151), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4640 ( .A1(n3733), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3666) );
  NAND4_X1 U4641 ( .A1(n3669), .A2(n3668), .A3(n3667), .A4(n3666), .ZN(n3676)
         );
  AOI22_X1 U4642 ( .A1(n4188), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3673) );
  AOI22_X1 U4643 ( .A1(n3388), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4644 ( .A1(n3015), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4181), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4645 ( .A1(n3354), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3670) );
  NAND4_X1 U4646 ( .A1(n3673), .A2(n3672), .A3(n3671), .A4(n3670), .ZN(n3675)
         );
  OAI21_X1 U4647 ( .B1(n3676), .B2(n3675), .A(n3674), .ZN(n3679) );
  NAND2_X1 U4648 ( .A1(n4207), .A2(EAX_REG_15__SCAN_IN), .ZN(n3678) );
  NAND2_X1 U4649 ( .A1(n4206), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3677)
         );
  NAND3_X1 U4650 ( .A1(n3679), .A2(n3678), .A3(n3677), .ZN(n3680) );
  AOI21_X1 U4651 ( .B1(n5627), .B2(n4202), .A(n3680), .ZN(n5411) );
  XNOR2_X1 U4652 ( .A(n3682), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5992)
         );
  AOI22_X1 U4653 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n3354), .B1(n3733), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4654 ( .A1(n4188), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4655 ( .A1(n3015), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4181), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4656 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n3790), .B1(n4145), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3683) );
  NAND4_X1 U4657 ( .A1(n3686), .A2(n3685), .A3(n3684), .A4(n3683), .ZN(n3692)
         );
  AOI22_X1 U4658 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n3374), .B1(n3016), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4659 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n3337), .B1(n3369), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4660 ( .A1(n3750), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4661 ( .A1(n3785), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3687) );
  NAND4_X1 U4662 ( .A1(n3690), .A2(n3689), .A3(n3688), .A4(n3687), .ZN(n3691)
         );
  NOR2_X1 U4663 ( .A1(n3692), .A2(n3691), .ZN(n3694) );
  AOI22_X1 U4664 ( .A1(n4207), .A2(EAX_REG_16__SCAN_IN), .B1(n4206), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3693) );
  OAI21_X1 U4665 ( .B1(n4173), .B2(n3694), .A(n3693), .ZN(n3695) );
  AOI21_X1 U4666 ( .B1(n5992), .B2(n4202), .A(n3695), .ZN(n5500) );
  NAND2_X1 U4667 ( .A1(n3697), .A2(n3696), .ZN(n5487) );
  AOI22_X1 U4668 ( .A1(n4188), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4669 ( .A1(n3355), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4670 ( .A1(n4151), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4671 ( .A1(n3790), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3698) );
  NAND4_X1 U4672 ( .A1(n3701), .A2(n3700), .A3(n3699), .A4(n3698), .ZN(n3707)
         );
  AOI22_X1 U4673 ( .A1(n3388), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4674 ( .A1(n3337), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4675 ( .A1(n4181), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4676 ( .A1(n3785), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3702) );
  NAND4_X1 U4677 ( .A1(n3705), .A2(n3704), .A3(n3703), .A4(n3702), .ZN(n3706)
         );
  NOR2_X1 U4678 ( .A1(n3707), .A2(n3706), .ZN(n3711) );
  NAND2_X1 U4679 ( .A1(n4573), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3708)
         );
  NAND2_X1 U4680 ( .A1(n3524), .A2(n3708), .ZN(n3709) );
  AOI21_X1 U4681 ( .B1(n3417), .B2(EAX_REG_17__SCAN_IN), .A(n3709), .ZN(n3710)
         );
  OAI21_X1 U4682 ( .B1(n4173), .B2(n3711), .A(n3710), .ZN(n3714) );
  OAI21_X1 U4683 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3712), .A(n3728), 
        .ZN(n5987) );
  OR2_X1 U4684 ( .A1(n3524), .A2(n5987), .ZN(n3713) );
  NAND2_X1 U4685 ( .A1(n3714), .A2(n3713), .ZN(n5488) );
  AOI22_X1 U4686 ( .A1(n3355), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4687 ( .A1(n3790), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4688 ( .A1(n3337), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4689 ( .A1(n4146), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3715) );
  NAND4_X1 U4690 ( .A1(n3718), .A2(n3717), .A3(n3716), .A4(n3715), .ZN(n3724)
         );
  AOI22_X1 U4691 ( .A1(n4188), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3374), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4692 ( .A1(n4151), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4693 ( .A1(n3750), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4181), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4694 ( .A1(n3015), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3719) );
  NAND4_X1 U4695 ( .A1(n3722), .A2(n3721), .A3(n3720), .A4(n3719), .ZN(n3723)
         );
  NOR2_X1 U4696 ( .A1(n3724), .A2(n3723), .ZN(n3727) );
  AOI21_X1 U4697 ( .B1(n3197), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3725) );
  AOI21_X1 U4698 ( .B1(n3417), .B2(EAX_REG_18__SCAN_IN), .A(n3725), .ZN(n3726)
         );
  OAI21_X1 U4699 ( .B1(n4173), .B2(n3727), .A(n3726), .ZN(n3730) );
  XNOR2_X1 U4700 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3728), .ZN(n5612)
         );
  NAND2_X1 U4701 ( .A1(n4202), .A2(n5612), .ZN(n3729) );
  NAND2_X1 U4702 ( .A1(n5399), .A2(n5400), .ZN(n5398) );
  INV_X1 U4703 ( .A(n5398), .ZN(n3749) );
  OR2_X1 U4704 ( .A1(n3731), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3732)
         );
  NAND2_X1 U4705 ( .A1(n3732), .A2(n3764), .ZN(n5909) );
  AOI22_X1 U4706 ( .A1(n3388), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3750), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4707 ( .A1(n4151), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4708 ( .A1(n3733), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4181), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4709 ( .A1(n3337), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3734) );
  NAND4_X1 U4710 ( .A1(n3737), .A2(n3736), .A3(n3735), .A4(n3734), .ZN(n3743)
         );
  AOI22_X1 U4711 ( .A1(n3354), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3015), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4712 ( .A1(n3785), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4713 ( .A1(n4188), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4714 ( .A1(n3790), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3738) );
  NAND4_X1 U4715 ( .A1(n3741), .A2(n3740), .A3(n3739), .A4(n3738), .ZN(n3742)
         );
  NOR2_X1 U4716 ( .A1(n3743), .A2(n3742), .ZN(n3746) );
  INV_X1 U4717 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6730) );
  OAI21_X1 U4718 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6730), .A(n4573), 
        .ZN(n3745) );
  NAND2_X1 U4719 ( .A1(n4207), .A2(EAX_REG_19__SCAN_IN), .ZN(n3744) );
  OAI211_X1 U4720 ( .C1(n4173), .C2(n3746), .A(n3745), .B(n3744), .ZN(n3747)
         );
  OAI21_X1 U4721 ( .B1(n5909), .B2(n3524), .A(n3747), .ZN(n5476) );
  AOI22_X1 U4722 ( .A1(n3750), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3754) );
  AOI22_X1 U4723 ( .A1(n3355), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4724 ( .A1(n4188), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4725 ( .A1(n3369), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3751) );
  NAND4_X1 U4726 ( .A1(n3754), .A2(n3753), .A3(n3752), .A4(n3751), .ZN(n3760)
         );
  AOI22_X1 U4727 ( .A1(n3388), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3758) );
  AOI22_X1 U4728 ( .A1(n3337), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4729 ( .A1(n4181), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4730 ( .A1(n3790), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3755) );
  NAND4_X1 U4731 ( .A1(n3758), .A2(n3757), .A3(n3756), .A4(n3755), .ZN(n3759)
         );
  NOR2_X1 U4732 ( .A1(n3760), .A2(n3759), .ZN(n3763) );
  INV_X1 U4733 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5861) );
  OAI21_X1 U4734 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5861), .A(n3524), .ZN(
        n3761) );
  AOI21_X1 U4735 ( .B1(n3417), .B2(EAX_REG_20__SCAN_IN), .A(n3761), .ZN(n3762)
         );
  OAI21_X1 U4736 ( .B1(n4173), .B2(n3763), .A(n3762), .ZN(n3766) );
  XNOR2_X1 U4737 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n3764), .ZN(n5852)
         );
  NAND2_X1 U4738 ( .A1(n5852), .A2(n4202), .ZN(n3765) );
  NAND2_X1 U4739 ( .A1(n3766), .A2(n3765), .ZN(n5470) );
  AOI22_X1 U4740 ( .A1(n4188), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4741 ( .A1(n3390), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4742 ( .A1(n3790), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4743 ( .A1(n3733), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3767) );
  NAND4_X1 U4744 ( .A1(n3770), .A2(n3769), .A3(n3768), .A4(n3767), .ZN(n3776)
         );
  AOI22_X1 U4745 ( .A1(n3374), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4746 ( .A1(n3337), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4747 ( .A1(n4181), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4748 ( .A1(n3015), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3771) );
  NAND4_X1 U4749 ( .A1(n3774), .A2(n3773), .A3(n3772), .A4(n3771), .ZN(n3775)
         );
  NOR2_X1 U4750 ( .A1(n3776), .A2(n3775), .ZN(n3780) );
  NAND2_X1 U4751 ( .A1(n4573), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3777)
         );
  NAND2_X1 U4752 ( .A1(n3524), .A2(n3777), .ZN(n3778) );
  AOI21_X1 U4753 ( .B1(n3417), .B2(EAX_REG_21__SCAN_IN), .A(n3778), .ZN(n3779)
         );
  OAI21_X1 U4754 ( .B1(n4173), .B2(n3780), .A(n3779), .ZN(n3783) );
  OAI21_X1 U4755 ( .B1(n3781), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n3800), 
        .ZN(n5846) );
  OR2_X1 U4756 ( .A1(n5846), .A2(n3524), .ZN(n3782) );
  NAND2_X1 U4757 ( .A1(n3783), .A2(n3782), .ZN(n5464) );
  AOI22_X1 U4758 ( .A1(n4188), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4759 ( .A1(n3390), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3015), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4760 ( .A1(n3337), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4761 ( .A1(n3733), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3786) );
  NAND4_X1 U4762 ( .A1(n3789), .A2(n3788), .A3(n3787), .A4(n3786), .ZN(n3796)
         );
  AOI22_X1 U4763 ( .A1(n3388), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4764 ( .A1(n3790), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4765 ( .A1(n4181), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4766 ( .A1(n3354), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3791) );
  NAND4_X1 U4767 ( .A1(n3794), .A2(n3793), .A3(n3792), .A4(n3791), .ZN(n3795)
         );
  NOR2_X1 U4768 ( .A1(n3796), .A2(n3795), .ZN(n3799) );
  OAI21_X1 U4769 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5588), .A(n3524), .ZN(
        n3797) );
  AOI21_X1 U4770 ( .B1(n3417), .B2(EAX_REG_22__SCAN_IN), .A(n3797), .ZN(n3798)
         );
  OAI21_X1 U4771 ( .B1(n4173), .B2(n3799), .A(n3798), .ZN(n3802) );
  XNOR2_X1 U4772 ( .A(n3800), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5842)
         );
  NAND2_X1 U4773 ( .A1(n5842), .A2(n4202), .ZN(n3801) );
  XNOR2_X1 U4774 ( .A(n3804), .B(n3803), .ZN(n3805) );
  OR2_X1 U4775 ( .A1(n4173), .A2(n3805), .ZN(n3812) );
  NAND2_X1 U4776 ( .A1(n4124), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3806)
         );
  NAND2_X1 U4777 ( .A1(n3524), .A2(n3806), .ZN(n3807) );
  AOI21_X1 U4778 ( .B1(n3417), .B2(EAX_REG_23__SCAN_IN), .A(n3807), .ZN(n3811)
         );
  OR2_X1 U4779 ( .A1(n3808), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3809)
         );
  NAND2_X1 U4780 ( .A1(n3816), .A2(n3809), .ZN(n5825) );
  NOR2_X1 U4781 ( .A1(n5825), .A2(n3524), .ZN(n3810) );
  AOI21_X1 U4782 ( .B1(n3812), .B2(n3811), .A(n3810), .ZN(n5448) );
  INV_X1 U4783 ( .A(n4173), .ZN(n4197) );
  INV_X1 U4784 ( .A(n3813), .ZN(n3814) );
  XNOR2_X1 U4785 ( .A(n3815), .B(n3814), .ZN(n3820) );
  XNOR2_X1 U4786 ( .A(n3816), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5818)
         );
  NAND2_X1 U4787 ( .A1(n4207), .A2(EAX_REG_24__SCAN_IN), .ZN(n3818) );
  NAND2_X1 U4788 ( .A1(n4206), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3817)
         );
  OAI211_X1 U4789 ( .C1(n5818), .C2(n3524), .A(n3818), .B(n3817), .ZN(n3819)
         );
  AOI21_X1 U4790 ( .B1(n4197), .B2(n3820), .A(n3819), .ZN(n5442) );
  XNOR2_X1 U4791 ( .A(n3822), .B(n3821), .ZN(n3826) );
  NAND2_X1 U4792 ( .A1(n4124), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3823)
         );
  NAND2_X1 U4793 ( .A1(n3524), .A2(n3823), .ZN(n3824) );
  AOI21_X1 U4794 ( .B1(n3417), .B2(EAX_REG_25__SCAN_IN), .A(n3824), .ZN(n3825)
         );
  OAI21_X1 U4795 ( .B1(n3826), .B2(n4173), .A(n3825), .ZN(n3830) );
  OR2_X1 U4796 ( .A1(n3827), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3828)
         );
  NAND2_X1 U4797 ( .A1(n3828), .A2(n3897), .ZN(n5904) );
  NAND2_X1 U4798 ( .A1(n3830), .A2(n3829), .ZN(n5384) );
  INV_X1 U4799 ( .A(n5565), .ZN(n5517) );
  NAND2_X1 U4800 ( .A1(n3088), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3833) );
  NAND2_X1 U4801 ( .A1(n3834), .A2(n3833), .ZN(n3846) );
  INV_X1 U4802 ( .A(n3834), .ZN(n3835) );
  NAND2_X1 U4803 ( .A1(n5336), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3836) );
  INV_X1 U4804 ( .A(n3841), .ZN(n3840) );
  NAND2_X1 U4805 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3841), .ZN(n3842) );
  XNOR2_X1 U4806 ( .A(n3844), .B(n3843), .ZN(n3888) );
  OAI21_X1 U4807 ( .B1(n3882), .B2(n4615), .A(n5338), .ZN(n3856) );
  AOI21_X1 U4808 ( .B1(n3847), .B2(n3846), .A(n3845), .ZN(n3886) );
  OAI21_X1 U4809 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6430), .A(n3847), 
        .ZN(n3849) );
  NOR2_X1 U4810 ( .A1(n3882), .A2(n3849), .ZN(n3852) );
  AND2_X1 U4811 ( .A1(n4615), .A2(n5338), .ZN(n3848) );
  INV_X1 U4812 ( .A(n4111), .ZN(n3850) );
  OAI21_X1 U4813 ( .B1(n3850), .B2(n3849), .A(n3295), .ZN(n3851) );
  NAND2_X1 U4814 ( .A1(n3870), .A2(n3851), .ZN(n3853) );
  OAI211_X1 U4815 ( .C1(n3856), .C2(n3886), .A(n3852), .B(n3853), .ZN(n3855)
         );
  INV_X1 U4816 ( .A(n3853), .ZN(n3854) );
  AOI22_X1 U4817 ( .A1(n3883), .A2(n3855), .B1(n3854), .B2(n3886), .ZN(n3868)
         );
  INV_X1 U4818 ( .A(n3856), .ZN(n3858) );
  INV_X1 U4819 ( .A(n3886), .ZN(n3857) );
  NOR3_X1 U4820 ( .A1(n3858), .A2(n6474), .A3(n3857), .ZN(n3867) );
  OR2_X1 U4821 ( .A1(n3860), .A2(n3859), .ZN(n3862) );
  AND2_X1 U4822 ( .A1(n3862), .A2(n3861), .ZN(n3887) );
  INV_X1 U4823 ( .A(n3887), .ZN(n3863) );
  OAI21_X1 U4824 ( .B1(n3882), .B2(n3863), .A(n3870), .ZN(n3864) );
  NAND2_X1 U4825 ( .A1(n3864), .A2(n3888), .ZN(n3869) );
  OAI21_X1 U4826 ( .B1(n3887), .B2(n3865), .A(n3869), .ZN(n3866) );
  OAI21_X1 U4827 ( .B1(n3868), .B2(n3867), .A(n3866), .ZN(n3875) );
  INV_X1 U4828 ( .A(n3869), .ZN(n3873) );
  INV_X1 U4829 ( .A(n3882), .ZN(n3872) );
  INV_X1 U4830 ( .A(n3870), .ZN(n3871) );
  NAND4_X1 U4831 ( .A1(n3873), .A2(n3887), .A3(n3872), .A4(n3871), .ZN(n3874)
         );
  OAI211_X1 U4832 ( .C1(n3888), .C2(n3883), .A(n3875), .B(n3874), .ZN(n3876)
         );
  NAND3_X1 U4833 ( .A1(n3888), .A2(n3887), .A3(n3886), .ZN(n3890) );
  OAI21_X1 U4834 ( .B1(n3891), .B2(n3890), .A(n3889), .ZN(n6448) );
  NOR2_X1 U4835 ( .A1(n3297), .A2(n3295), .ZN(n3893) );
  NAND2_X1 U4836 ( .A1(n3892), .A2(n3893), .ZN(n6450) );
  NOR2_X1 U4837 ( .A1(n6448), .A2(n6450), .ZN(n5957) );
  NAND2_X1 U4838 ( .A1(n5957), .A2(n4506), .ZN(n4304) );
  NOR2_X1 U4839 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n3894) );
  INV_X1 U4840 ( .A(n3894), .ZN(n6484) );
  NOR3_X1 U4841 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6484), .A3(n4419), .ZN(
        n6479) );
  INV_X1 U4842 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6562) );
  NAND2_X1 U4843 ( .A1(n4419), .A2(n4573), .ZN(n6483) );
  NOR3_X1 U4844 ( .A1(n6474), .A2(n6562), .A3(n6483), .ZN(n6471) );
  AND2_X2 U4845 ( .A1(n4346), .A2(n3894), .ZN(n6133) );
  OR2_X1 U4846 ( .A1(n6471), .A2(n6133), .ZN(n3895) );
  NOR2_X1 U4847 ( .A1(n6479), .A2(n3895), .ZN(n3896) );
  INV_X1 U4848 ( .A(n3897), .ZN(n3898) );
  INV_X1 U4849 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4170) );
  NAND2_X1 U4850 ( .A1(n4162), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4201)
         );
  INV_X1 U4851 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5376) );
  INV_X1 U4852 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3899) );
  NOR2_X1 U4853 ( .A1(n4217), .A2(n4419), .ZN(n3901) );
  NOR2_X1 U4854 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4001) );
  INV_X1 U4855 ( .A(n4001), .ZN(n4002) );
  AND2_X1 U4856 ( .A1(n4989), .A2(n4002), .ZN(n3902) );
  INV_X1 U4857 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6214) );
  NAND2_X1 U4858 ( .A1(n3919), .A2(n6214), .ZN(n3906) );
  INV_X1 U4859 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4990) );
  NAND2_X1 U4860 ( .A1(n4989), .A2(n4990), .ZN(n3905) );
  NAND3_X1 U4861 ( .A1(n4296), .A2(n3906), .A3(n3905), .ZN(n3907) );
  NAND2_X1 U4862 ( .A1(n3919), .A2(EBX_REG_0__SCAN_IN), .ZN(n3909) );
  INV_X1 U4863 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4924) );
  NAND2_X1 U4864 ( .A1(n4296), .A2(n4924), .ZN(n3908) );
  AND2_X1 U4865 ( .A1(n3909), .A2(n3908), .ZN(n4923) );
  OAI21_X1 U4866 ( .B1(n4756), .B2(n5358), .A(n3910), .ZN(n4985) );
  OR2_X1 U4867 ( .A1(n4294), .A2(EBX_REG_2__SCAN_IN), .ZN(n3915) );
  INV_X1 U4868 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3911) );
  NAND2_X1 U4869 ( .A1(n3919), .A2(n3911), .ZN(n3913) );
  INV_X1 U4870 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U4871 ( .A1(n4989), .A2(n6079), .ZN(n3912) );
  NAND3_X1 U4872 ( .A1(n3913), .A2(n4296), .A3(n3912), .ZN(n3914) );
  AND2_X1 U4873 ( .A1(n3915), .A2(n3914), .ZN(n4984) );
  MUX2_X1 U4874 ( .A(n3978), .B(n4296), .S(EBX_REG_3__SCAN_IN), .Z(n3918) );
  OAI21_X1 U4875 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n5359), .A(n3918), 
        .ZN(n4994) );
  MUX2_X1 U4876 ( .A(n4294), .B(n3919), .S(EBX_REG_4__SCAN_IN), .Z(n3921) );
  INV_X1 U4877 ( .A(n3919), .ZN(n3958) );
  NAND2_X1 U4878 ( .A1(n3958), .A2(n5358), .ZN(n3975) );
  NAND2_X1 U4879 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n5358), .ZN(n3920)
         );
  AND3_X1 U4880 ( .A1(n3921), .A2(n3975), .A3(n3920), .ZN(n4538) );
  NOR2_X2 U4881 ( .A1(n4997), .A2(n4538), .ZN(n4537) );
  MUX2_X1 U4882 ( .A(n3978), .B(n4296), .S(EBX_REG_5__SCAN_IN), .Z(n3922) );
  OAI21_X1 U4883 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n5359), .A(n3922), 
        .ZN(n4555) );
  INV_X1 U4884 ( .A(n4555), .ZN(n3923) );
  NAND2_X1 U4885 ( .A1(n4537), .A2(n3923), .ZN(n4919) );
  MUX2_X1 U4886 ( .A(n3978), .B(n4296), .S(EBX_REG_7__SCAN_IN), .Z(n3924) );
  OAI21_X1 U4887 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n5359), .A(n3924), 
        .ZN(n4917) );
  INV_X1 U4888 ( .A(n4917), .ZN(n3929) );
  OR2_X1 U4889 ( .A1(n4294), .A2(EBX_REG_6__SCAN_IN), .ZN(n3928) );
  INV_X1 U4890 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4067) );
  NAND2_X1 U4891 ( .A1(n3919), .A2(n4067), .ZN(n3926) );
  INV_X1 U4892 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U4893 ( .A1(n4989), .A2(n6085), .ZN(n3925) );
  NAND3_X1 U4894 ( .A1(n3926), .A2(n4296), .A3(n3925), .ZN(n3927) );
  NAND2_X1 U4895 ( .A1(n3928), .A2(n3927), .ZN(n4916) );
  OR2_X1 U4896 ( .A1(n4294), .A2(EBX_REG_8__SCAN_IN), .ZN(n3934) );
  INV_X1 U4897 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U4898 ( .A1(n3919), .A2(n5078), .ZN(n3932) );
  INV_X1 U4899 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U4900 ( .A1(n4989), .A2(n6011), .ZN(n3931) );
  NAND3_X1 U4901 ( .A1(n3932), .A2(n4296), .A3(n3931), .ZN(n3933) );
  INV_X1 U4902 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U4903 ( .A1(n4250), .A2(n5058), .ZN(n3937) );
  NAND2_X1 U4904 ( .A1(n4296), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3935)
         );
  OAI211_X1 U4905 ( .C1(n5358), .C2(EBX_REG_9__SCAN_IN), .A(n3919), .B(n3935), 
        .ZN(n3936) );
  MUX2_X1 U4906 ( .A(n4294), .B(n3919), .S(EBX_REG_10__SCAN_IN), .Z(n3939) );
  NAND2_X1 U4907 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n5358), .ZN(n3938) );
  NAND2_X1 U4908 ( .A1(n4296), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3940) );
  OAI211_X1 U4909 ( .C1(n5358), .C2(EBX_REG_11__SCAN_IN), .A(n3919), .B(n3940), 
        .ZN(n3941) );
  OAI21_X1 U4910 ( .B1(n3978), .B2(EBX_REG_11__SCAN_IN), .A(n3941), .ZN(n5124)
         );
  OR2_X1 U4911 ( .A1(n4294), .A2(EBX_REG_12__SCAN_IN), .ZN(n3945) );
  NAND2_X1 U4912 ( .A1(n3919), .A2(n2999), .ZN(n3943) );
  INV_X1 U4913 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5191) );
  NAND2_X1 U4914 ( .A1(n4989), .A2(n5191), .ZN(n3942) );
  NAND3_X1 U4915 ( .A1(n3943), .A2(n4296), .A3(n3942), .ZN(n3944) );
  NAND2_X1 U4916 ( .A1(n3945), .A2(n3944), .ZN(n5185) );
  INV_X1 U4917 ( .A(n5359), .ZN(n3947) );
  INV_X1 U4918 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3946) );
  NAND2_X1 U4919 ( .A1(n3947), .A2(n3946), .ZN(n3949) );
  MUX2_X1 U4920 ( .A(n3978), .B(n4296), .S(EBX_REG_13__SCAN_IN), .Z(n3948) );
  AND2_X1 U4921 ( .A1(n3949), .A2(n3948), .ZN(n5272) );
  MUX2_X1 U4922 ( .A(n4294), .B(n3919), .S(EBX_REG_14__SCAN_IN), .Z(n3951) );
  NAND2_X1 U4923 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5358), .ZN(n3950) );
  MUX2_X1 U4924 ( .A(n3978), .B(n4296), .S(EBX_REG_15__SCAN_IN), .Z(n3952) );
  OAI21_X1 U4925 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n5359), .A(n3952), 
        .ZN(n5414) );
  MUX2_X1 U4926 ( .A(n4294), .B(n3919), .S(EBX_REG_16__SCAN_IN), .Z(n3954) );
  NAND2_X1 U4927 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n5358), .ZN(n3953) );
  NOR2_X2 U4928 ( .A1(n5496), .A2(n5495), .ZN(n5497) );
  INV_X1 U4929 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U4930 ( .A1(n4250), .A2(n5493), .ZN(n3957) );
  NAND2_X1 U4931 ( .A1(n4296), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3955) );
  OAI211_X1 U4932 ( .C1(n5358), .C2(EBX_REG_17__SCAN_IN), .A(n3919), .B(n3955), 
        .ZN(n3956) );
  OR2_X1 U4933 ( .A1(n4294), .A2(EBX_REG_19__SCAN_IN), .ZN(n3963) );
  INV_X1 U4934 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3959) );
  NAND2_X1 U4935 ( .A1(n3919), .A2(n3959), .ZN(n3961) );
  INV_X1 U4936 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U4937 ( .A1(n4989), .A2(n5482), .ZN(n3960) );
  NAND3_X1 U4938 ( .A1(n3961), .A2(n4296), .A3(n3960), .ZN(n3962) );
  AND2_X1 U4939 ( .A1(n3963), .A2(n3962), .ZN(n5478) );
  OR2_X1 U4940 ( .A1(n5359), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3965)
         );
  INV_X1 U4941 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U4942 ( .A1(n4989), .A2(n5475), .ZN(n3964) );
  AND2_X1 U4943 ( .A1(n3965), .A2(n3964), .ZN(n5473) );
  OR2_X1 U4944 ( .A1(n5359), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3966)
         );
  INV_X1 U4945 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U4946 ( .A1(n4989), .A2(n5405), .ZN(n5402) );
  NAND2_X1 U4947 ( .A1(n3966), .A2(n5402), .ZN(n5472) );
  NAND2_X1 U4948 ( .A1(n3904), .A2(EBX_REG_20__SCAN_IN), .ZN(n3968) );
  NAND2_X1 U4949 ( .A1(n5472), .A2(n4296), .ZN(n3967) );
  OAI211_X1 U4950 ( .C1(n5473), .C2(n5472), .A(n3968), .B(n3967), .ZN(n3969)
         );
  INV_X1 U4951 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U4952 ( .A1(n4250), .A2(n5467), .ZN(n3973) );
  NAND2_X1 U4953 ( .A1(n4989), .A2(n5467), .ZN(n3971) );
  NAND2_X1 U4954 ( .A1(n4296), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3970) );
  NAND3_X1 U4955 ( .A1(n3971), .A2(n3919), .A3(n3970), .ZN(n3972) );
  MUX2_X1 U4956 ( .A(n4294), .B(n3919), .S(EBX_REG_22__SCAN_IN), .Z(n3977) );
  NAND2_X1 U4957 ( .A1(n5358), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3974) );
  AND2_X1 U4958 ( .A1(n3975), .A2(n3974), .ZN(n3976) );
  NAND2_X1 U4959 ( .A1(n3977), .A2(n3976), .ZN(n5456) );
  MUX2_X1 U4960 ( .A(n3978), .B(n4296), .S(EBX_REG_23__SCAN_IN), .Z(n3979) );
  OAI21_X1 U4961 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5359), .A(n3979), 
        .ZN(n5451) );
  OR2_X2 U4962 ( .A1(n5450), .A2(n5451), .ZN(n5453) );
  INV_X1 U4963 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U4964 ( .A1(n4250), .A2(n5437), .ZN(n3983) );
  NAND2_X1 U4965 ( .A1(n4989), .A2(n5437), .ZN(n3981) );
  NAND2_X1 U4966 ( .A1(n4296), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3980) );
  NAND3_X1 U4967 ( .A1(n3981), .A2(n3919), .A3(n3980), .ZN(n3982) );
  AND2_X1 U4968 ( .A1(n3983), .A2(n3982), .ZN(n5386) );
  OR2_X1 U4969 ( .A1(n4294), .A2(EBX_REG_24__SCAN_IN), .ZN(n3987) );
  INV_X1 U4970 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5718) );
  NAND2_X1 U4971 ( .A1(n3919), .A2(n5718), .ZN(n3985) );
  INV_X1 U4972 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U4973 ( .A1(n4989), .A2(n5445), .ZN(n3984) );
  NAND3_X1 U4974 ( .A1(n3985), .A2(n4296), .A3(n3984), .ZN(n3986) );
  NAND2_X1 U4975 ( .A1(n3987), .A2(n3986), .ZN(n5443) );
  NAND2_X1 U4976 ( .A1(n5386), .A2(n5443), .ZN(n3988) );
  MUX2_X1 U4977 ( .A(n4294), .B(n3919), .S(EBX_REG_26__SCAN_IN), .Z(n3990) );
  NAND2_X1 U4978 ( .A1(n5358), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3989) );
  NAND2_X1 U4979 ( .A1(n3990), .A2(n3989), .ZN(n3992) );
  AND2_X2 U4980 ( .A1(n5388), .A2(n3992), .ZN(n5693) );
  INV_X1 U4981 ( .A(n5693), .ZN(n3991) );
  OAI21_X1 U4982 ( .B1(n5388), .B2(n3992), .A(n3991), .ZN(n5710) );
  OAI22_X1 U4983 ( .A1(n5517), .A2(n5856), .B1(n6061), .B2(n5710), .ZN(n4013)
         );
  INV_X1 U4984 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U4985 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5836) );
  INV_X1 U4986 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6528) );
  INV_X1 U4987 ( .A(REIP_REG_11__SCAN_IN), .ZN(n3993) );
  INV_X1 U4988 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6518) );
  INV_X1 U4989 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6512) );
  INV_X1 U4990 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6574) );
  INV_X1 U4991 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6508) );
  INV_X1 U4992 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6506) );
  NOR3_X1 U4993 ( .A1(n6574), .A2(n6508), .A3(n6506), .ZN(n6053) );
  NAND2_X1 U4994 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6053), .ZN(n6008) );
  NOR2_X1 U4995 ( .A1(n6512), .A2(n6008), .ZN(n6019) );
  NAND4_X1 U4996 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6019), .A3(
        REIP_REG_7__SCAN_IN), .A4(REIP_REG_6__SCAN_IN), .ZN(n5102) );
  NOR2_X1 U4997 ( .A1(n6518), .A2(n5102), .ZN(n6003) );
  NAND2_X1 U4998 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6003), .ZN(n5174) );
  NAND4_X1 U4999 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .A4(n5269), .ZN(n5429) );
  NAND3_X1 U5000 ( .A1(n5412), .A2(REIP_REG_17__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .ZN(n5863) );
  INV_X1 U5001 ( .A(n5863), .ZN(n3994) );
  NAND4_X1 U5002 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(n3994), .ZN(n5835) );
  INV_X1 U5003 ( .A(n5835), .ZN(n3997) );
  OR2_X1 U5004 ( .A1(n3995), .A2(STATE_REG_0__SCAN_IN), .ZN(n6496) );
  NAND2_X1 U5005 ( .A1(n4615), .A2(n6496), .ZN(n4508) );
  AND3_X1 U5006 ( .A1(n4508), .A2(n4001), .A3(n3295), .ZN(n3996) );
  NAND2_X1 U5007 ( .A1(n3997), .A2(n6054), .ZN(n5847) );
  NAND2_X1 U5008 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5831), .ZN(n5392) );
  INV_X1 U5009 ( .A(n5392), .ZN(n3998) );
  NAND2_X1 U5010 ( .A1(REIP_REG_24__SCAN_IN), .A2(n3998), .ZN(n5385) );
  INV_X1 U5011 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6623) );
  OAI21_X1 U5012 ( .B1(n6542), .B2(n5385), .A(n6623), .ZN(n4000) );
  INV_X1 U5013 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6657) );
  NOR3_X1 U5014 ( .A1(n6657), .A2(n5835), .A3(n5836), .ZN(n5390) );
  NAND3_X1 U5015 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4274) );
  INV_X1 U5016 ( .A(n4274), .ZN(n3999) );
  NAND2_X1 U5017 ( .A1(n6069), .A2(n6068), .ZN(n5864) );
  INV_X1 U5018 ( .A(n5864), .ZN(n5391) );
  AOI21_X1 U5019 ( .B1(n5390), .B2(n3999), .A(n5391), .ZN(n5814) );
  INV_X1 U5020 ( .A(n6496), .ZN(n4502) );
  NAND2_X1 U5021 ( .A1(n4502), .A2(n4001), .ZN(n6466) );
  NAND2_X1 U5022 ( .A1(n3314), .A2(n6466), .ZN(n5366) );
  INV_X1 U5023 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5434) );
  NAND3_X1 U5024 ( .A1(n3295), .A2(n5434), .A3(n4002), .ZN(n4003) );
  NAND2_X1 U5025 ( .A1(n5366), .A2(n4003), .ZN(n4004) );
  AOI22_X1 U5026 ( .A1(EBX_REG_26__SCAN_IN), .A2(n6050), .B1(n5561), .B2(n6071), .ZN(n4006) );
  INV_X1 U5027 ( .A(n4006), .ZN(n4009) );
  OR2_X1 U5028 ( .A1(n4013), .A2(n4012), .ZN(U2801) );
  NAND2_X1 U5029 ( .A1(n4014), .A2(n4082), .ZN(n4018) );
  NAND2_X1 U5030 ( .A1(n4022), .A2(n4023), .ZN(n4033) );
  NAND2_X1 U5031 ( .A1(n4033), .A2(n4034), .ZN(n4043) );
  NAND2_X1 U5032 ( .A1(n4043), .A2(n4044), .ZN(n4055) );
  XNOR2_X1 U5033 ( .A(n4055), .B(n4015), .ZN(n4016) );
  NAND2_X1 U5034 ( .A1(n4016), .A2(n3314), .ZN(n4017) );
  INV_X1 U5035 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4541) );
  INV_X1 U5036 ( .A(n4082), .ZN(n4032) );
  NAND2_X1 U5037 ( .A1(n4580), .A2(n4019), .ZN(n4035) );
  OAI21_X1 U5038 ( .B1(n6592), .B2(n4022), .A(n4035), .ZN(n4020) );
  INV_X1 U5039 ( .A(n4020), .ZN(n4021) );
  OAI21_X1 U5040 ( .B1(n4853), .B2(n4032), .A(n4021), .ZN(n6144) );
  XNOR2_X1 U5041 ( .A(n4029), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4440)
         );
  NAND2_X1 U5042 ( .A1(n4481), .A2(n4082), .ZN(n4028) );
  OAI21_X1 U5043 ( .B1(n4023), .B2(n4022), .A(n4033), .ZN(n4025) );
  INV_X1 U5044 ( .A(n4235), .ZN(n4024) );
  OAI211_X1 U5045 ( .C1(n4025), .C2(n6592), .A(n4024), .B(n5338), .ZN(n4026)
         );
  INV_X1 U5046 ( .A(n4026), .ZN(n4027) );
  NAND2_X1 U5047 ( .A1(n4028), .A2(n4027), .ZN(n4439) );
  NAND2_X1 U5048 ( .A1(n4440), .A2(n4439), .ZN(n4438) );
  INV_X1 U5049 ( .A(n4029), .ZN(n4030) );
  NAND2_X1 U5050 ( .A1(n4030), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4031)
         );
  OAI21_X1 U5051 ( .B1(n4034), .B2(n4033), .A(n4043), .ZN(n4037) );
  INV_X1 U5052 ( .A(n4035), .ZN(n4036) );
  AOI21_X1 U5053 ( .B1(n4037), .B2(n3314), .A(n4036), .ZN(n4038) );
  OAI21_X1 U5054 ( .B1(n6136), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(n6134), 
        .ZN(n4041) );
  NAND2_X1 U5055 ( .A1(n6136), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4040)
         );
  NAND2_X1 U5056 ( .A1(n4041), .A2(n4040), .ZN(n4454) );
  NAND2_X1 U5057 ( .A1(n4042), .A2(n4082), .ZN(n4046) );
  OAI211_X1 U5058 ( .C1(n4044), .C2(n4043), .A(n4055), .B(n3314), .ZN(n4045)
         );
  INV_X1 U5059 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U5060 ( .A1(n4454), .A2(n4455), .ZN(n4049) );
  NAND2_X1 U5061 ( .A1(n4047), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4048)
         );
  NAND2_X1 U5062 ( .A1(n4049), .A2(n4048), .ZN(n4526) );
  NAND2_X1 U5063 ( .A1(n4525), .A2(n4526), .ZN(n4052) );
  NAND2_X1 U5064 ( .A1(n4050), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4051)
         );
  NAND2_X1 U5065 ( .A1(n4053), .A2(n4082), .ZN(n4059) );
  NOR2_X1 U5066 ( .A1(n4055), .A2(n4054), .ZN(n4057) );
  NAND2_X1 U5067 ( .A1(n4057), .A2(n4056), .ZN(n4072) );
  OAI211_X1 U5068 ( .C1(n4057), .C2(n4056), .A(n4072), .B(n3314), .ZN(n4058)
         );
  NAND2_X1 U5069 ( .A1(n4059), .A2(n4058), .ZN(n4060) );
  INV_X1 U5070 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4552) );
  XNOR2_X1 U5071 ( .A(n4060), .B(n4552), .ZN(n4548) );
  NAND2_X1 U5072 ( .A1(n4547), .A2(n4548), .ZN(n4062) );
  NAND2_X1 U5073 ( .A1(n4060), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4061)
         );
  NAND3_X1 U5074 ( .A1(n4081), .A2(n4063), .A3(n4082), .ZN(n4066) );
  XNOR2_X1 U5075 ( .A(n4072), .B(n4073), .ZN(n4064) );
  NAND2_X1 U5076 ( .A1(n4064), .A2(n3314), .ZN(n4065) );
  NAND2_X1 U5077 ( .A1(n4066), .A2(n4065), .ZN(n4068) );
  XNOR2_X1 U5078 ( .A(n4068), .B(n4067), .ZN(n4692) );
  NAND2_X1 U5079 ( .A1(n4691), .A2(n4692), .ZN(n4070) );
  NAND2_X1 U5080 ( .A1(n4068), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4069)
         );
  NAND2_X1 U5081 ( .A1(n4071), .A2(n4082), .ZN(n4077) );
  INV_X1 U5082 ( .A(n4072), .ZN(n4074) );
  NAND2_X1 U5083 ( .A1(n4074), .A2(n4073), .ZN(n4084) );
  XNOR2_X1 U5084 ( .A(n4084), .B(n4085), .ZN(n4075) );
  NAND2_X1 U5085 ( .A1(n4075), .A2(n3314), .ZN(n4076) );
  NAND2_X1 U5086 ( .A1(n4077), .A2(n4076), .ZN(n4078) );
  INV_X1 U5087 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6177) );
  XNOR2_X1 U5088 ( .A(n4078), .B(n6177), .ZN(n5084) );
  NAND2_X1 U5089 ( .A1(n5083), .A2(n5084), .ZN(n4080) );
  NAND2_X1 U5090 ( .A1(n4078), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4079)
         );
  NAND2_X1 U5091 ( .A1(n4080), .A2(n4079), .ZN(n5067) );
  INV_X1 U5092 ( .A(n4084), .ZN(n4086) );
  NAND3_X1 U5093 ( .A1(n4086), .A2(n3314), .A3(n4085), .ZN(n4087) );
  NAND2_X1 U5094 ( .A1(n4090), .A2(n4087), .ZN(n4088) );
  XNOR2_X1 U5095 ( .A(n4088), .B(n5078), .ZN(n5068) );
  NAND2_X1 U5096 ( .A1(n4088), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4089)
         );
  INV_X1 U5097 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U5098 ( .A1(n5618), .A2(n6167), .ZN(n4091) );
  NAND2_X1 U5099 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4093) );
  INV_X1 U5100 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5239) );
  OR2_X1 U5101 ( .A1(n5606), .A2(n5239), .ZN(n5252) );
  INV_X1 U5102 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6153) );
  OR2_X1 U5103 ( .A1(n5606), .A2(n6153), .ZN(n5254) );
  XNOR2_X1 U5104 ( .A(n5618), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5311)
         );
  NAND2_X1 U5105 ( .A1(n5618), .A2(n3946), .ZN(n4094) );
  INV_X1 U5106 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5945) );
  AND2_X1 U5107 ( .A1(n5606), .A2(n5945), .ZN(n5633) );
  INV_X1 U5108 ( .A(n4095), .ZN(n5623) );
  XNOR2_X1 U5109 ( .A(n5618), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5624)
         );
  INV_X1 U5110 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U5111 ( .A1(n5618), .A2(n5794), .ZN(n4096) );
  INV_X1 U5112 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U5113 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U5114 ( .A1(n5606), .A2(n5642), .ZN(n4098) );
  INV_X1 U5115 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5608) );
  INV_X1 U5116 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5921) );
  AND3_X1 U5117 ( .A1(n5608), .A2(n5780), .A3(n5921), .ZN(n4099) );
  NOR2_X1 U5118 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5749) );
  NOR2_X1 U5119 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4101) );
  INV_X1 U5120 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5726) );
  AND4_X1 U5121 ( .A1(n5749), .A2(n4101), .A3(n5718), .A4(n5726), .ZN(n4102)
         );
  NAND2_X1 U5122 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5654) );
  AND2_X1 U5123 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5648) );
  AND2_X1 U5124 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5643) );
  NAND2_X1 U5125 ( .A1(n5648), .A2(n5643), .ZN(n5715) );
  OAI21_X1 U5126 ( .B1(n5654), .B2(n5715), .A(n5618), .ZN(n4103) );
  XNOR2_X1 U5127 ( .A(n5618), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5900)
         );
  INV_X1 U5128 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U5129 ( .A1(n5559), .A2(n3082), .ZN(n5551) );
  NAND2_X1 U5130 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U5131 ( .A1(n5529), .A2(n3086), .ZN(n4107) );
  NOR2_X1 U5132 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5684) );
  INV_X1 U5133 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5540) );
  NAND2_X1 U5134 ( .A1(n5684), .A2(n5540), .ZN(n4104) );
  NOR2_X1 U5135 ( .A1(n5618), .A2(n4104), .ZN(n4221) );
  INV_X1 U5136 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5666) );
  NAND3_X1 U5137 ( .A1(n4221), .A2(n5666), .A3(n5527), .ZN(n4105) );
  NAND2_X1 U5138 ( .A1(n4107), .A2(n4106), .ZN(n4108) );
  XNOR2_X1 U5139 ( .A(n4108), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5663)
         );
  NAND2_X1 U5140 ( .A1(n4344), .A2(n4580), .ZN(n4109) );
  NAND2_X1 U5141 ( .A1(n4110), .A2(n4109), .ZN(n4323) );
  AOI22_X1 U5142 ( .A1(n3374), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4115) );
  AOI22_X1 U5143 ( .A1(n3790), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3015), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4114) );
  AOI22_X1 U5144 ( .A1(n3337), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U5145 ( .A1(n3390), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4112) );
  NAND4_X1 U5146 ( .A1(n4115), .A2(n4114), .A3(n4113), .A4(n4112), .ZN(n4121)
         );
  AOI22_X1 U5147 ( .A1(n3592), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4119) );
  AOI22_X1 U5148 ( .A1(n3354), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U5149 ( .A1(n3355), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4117) );
  AOI22_X1 U5150 ( .A1(n3369), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4116) );
  NAND4_X1 U5151 ( .A1(n4119), .A2(n4118), .A3(n4117), .A4(n4116), .ZN(n4120)
         );
  NOR2_X1 U5152 ( .A1(n4121), .A2(n4120), .ZN(n4144) );
  NAND2_X1 U5153 ( .A1(n4123), .A2(n4122), .ZN(n4143) );
  XNOR2_X1 U5154 ( .A(n4144), .B(n4143), .ZN(n4128) );
  NAND2_X1 U5155 ( .A1(n4124), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4125)
         );
  NAND2_X1 U5156 ( .A1(n3524), .A2(n4125), .ZN(n4126) );
  AOI21_X1 U5157 ( .B1(n3417), .B2(EAX_REG_27__SCAN_IN), .A(n4126), .ZN(n4127)
         );
  OAI21_X1 U5158 ( .B1(n4128), .B2(n4173), .A(n4127), .ZN(n4131) );
  OAI21_X1 U5159 ( .B1(n4129), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n4175), 
        .ZN(n5811) );
  OR2_X1 U5160 ( .A1(n5811), .A2(n3524), .ZN(n4130) );
  AOI22_X1 U5161 ( .A1(n3592), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U5162 ( .A1(n3388), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U5163 ( .A1(n3015), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U5164 ( .A1(n3785), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4133) );
  NAND4_X1 U5165 ( .A1(n4136), .A2(n4135), .A3(n4134), .A4(n4133), .ZN(n4142)
         );
  AOI22_X1 U5166 ( .A1(n3355), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4140) );
  AOI22_X1 U5167 ( .A1(n3337), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4139) );
  AOI22_X1 U5168 ( .A1(n4151), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U5169 ( .A1(n3790), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4182), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4137) );
  NAND4_X1 U5170 ( .A1(n4140), .A2(n4139), .A3(n4138), .A4(n4137), .ZN(n4141)
         );
  NOR2_X1 U5171 ( .A1(n4142), .A2(n4141), .ZN(n4180) );
  NOR2_X1 U5172 ( .A1(n4144), .A2(n4143), .ZN(n4169) );
  AOI22_X1 U5173 ( .A1(n3355), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U5174 ( .A1(n3790), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U5175 ( .A1(n3337), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U5176 ( .A1(n4146), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4147) );
  NAND4_X1 U5177 ( .A1(n4150), .A2(n4149), .A3(n4148), .A4(n4147), .ZN(n4157)
         );
  AOI22_X1 U5178 ( .A1(n3592), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3388), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U5179 ( .A1(n4151), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5180 ( .A1(n3390), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U5181 ( .A1(n4183), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4152) );
  NAND4_X1 U5182 ( .A1(n4155), .A2(n4154), .A3(n4153), .A4(n4152), .ZN(n4156)
         );
  OR2_X1 U5183 ( .A1(n4157), .A2(n4156), .ZN(n4168) );
  NAND2_X1 U5184 ( .A1(n4169), .A2(n4168), .ZN(n4179) );
  XNOR2_X1 U5185 ( .A(n4180), .B(n4179), .ZN(n4161) );
  NAND2_X1 U5186 ( .A1(n4573), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4158)
         );
  NAND2_X1 U5187 ( .A1(n3524), .A2(n4158), .ZN(n4159) );
  AOI21_X1 U5188 ( .B1(n3417), .B2(EAX_REG_29__SCAN_IN), .A(n4159), .ZN(n4160)
         );
  OAI21_X1 U5189 ( .B1(n4161), .B2(n4173), .A(n4160), .ZN(n4167) );
  INV_X1 U5190 ( .A(n4162), .ZN(n4164) );
  INV_X1 U5191 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4163) );
  NAND2_X1 U5192 ( .A1(n4164), .A2(n4163), .ZN(n4165) );
  NAND2_X1 U5193 ( .A1(n4201), .A2(n4165), .ZN(n4287) );
  NAND2_X1 U5194 ( .A1(n4167), .A2(n4166), .ZN(n4225) );
  XNOR2_X1 U5195 ( .A(n4169), .B(n4168), .ZN(n4174) );
  AOI21_X1 U5196 ( .B1(n4170), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4171) );
  AOI21_X1 U5197 ( .B1(n3417), .B2(EAX_REG_28__SCAN_IN), .A(n4171), .ZN(n4172)
         );
  OAI21_X1 U5198 ( .B1(n4174), .B2(n4173), .A(n4172), .ZN(n4177) );
  XNOR2_X1 U5199 ( .A(n4175), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5544)
         );
  NAND2_X1 U5200 ( .A1(n5544), .A2(n4202), .ZN(n4176) );
  NAND2_X1 U5201 ( .A1(n4177), .A2(n4176), .ZN(n4224) );
  NOR2_X1 U5202 ( .A1(n4180), .A2(n4179), .ZN(n4196) );
  AOI22_X1 U5203 ( .A1(n3374), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3390), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4187) );
  AOI22_X1 U5204 ( .A1(n4151), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4186) );
  AOI22_X1 U5205 ( .A1(n4181), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4185) );
  AOI22_X1 U5206 ( .A1(n4183), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4182), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4184) );
  NAND4_X1 U5207 ( .A1(n4187), .A2(n4186), .A3(n4185), .A4(n4184), .ZN(n4194)
         );
  AOI22_X1 U5208 ( .A1(n4188), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4192) );
  AOI22_X1 U5209 ( .A1(n3790), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3785), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4191) );
  AOI22_X1 U5210 ( .A1(n3337), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3369), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4190) );
  AOI22_X1 U5211 ( .A1(n3355), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3185), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4189) );
  NAND4_X1 U5212 ( .A1(n4192), .A2(n4191), .A3(n4190), .A4(n4189), .ZN(n4193)
         );
  NOR2_X1 U5213 ( .A1(n4194), .A2(n4193), .ZN(n4195) );
  XNOR2_X1 U5214 ( .A(n4196), .B(n4195), .ZN(n4198) );
  NAND2_X1 U5215 ( .A1(n4198), .A2(n4197), .ZN(n4205) );
  NAND2_X1 U5216 ( .A1(n4573), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4199)
         );
  NAND2_X1 U5217 ( .A1(n3524), .A2(n4199), .ZN(n4200) );
  AOI21_X1 U5218 ( .B1(n3417), .B2(EAX_REG_30__SCAN_IN), .A(n4200), .ZN(n4204)
         );
  XNOR2_X1 U5219 ( .A(n4201), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5375)
         );
  AND2_X1 U5220 ( .A1(n5375), .A2(n4202), .ZN(n4203) );
  NAND2_X1 U5221 ( .A1(n4234), .A2(n4232), .ZN(n4210) );
  AOI22_X1 U5222 ( .A1(n4207), .A2(EAX_REG_31__SCAN_IN), .B1(n4206), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4208) );
  INV_X1 U5223 ( .A(n4208), .ZN(n4209) );
  XNOR2_X2 U5224 ( .A(n4210), .B(n4209), .ZN(n5509) );
  NAND3_X1 U5225 ( .A1(n6474), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6485) );
  INV_X1 U5226 ( .A(n6485), .ZN(n4211) );
  NOR2_X2 U5227 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6568) );
  INV_X2 U5228 ( .A(n6371), .ZN(n6138) );
  NAND2_X1 U5229 ( .A1(n5509), .A2(n6138), .ZN(n4220) );
  NAND2_X1 U5230 ( .A1(n6587), .A2(n6586), .ZN(n4212) );
  NAND2_X1 U5231 ( .A1(n4212), .A2(n6474), .ZN(n4213) );
  AND2_X2 U5232 ( .A1(n6145), .A2(n4213), .ZN(n6148) );
  NAND2_X1 U5233 ( .A1(n6474), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4215) );
  NAND2_X1 U5234 ( .A1(n6730), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4214) );
  NAND2_X1 U5235 ( .A1(n4215), .A2(n4214), .ZN(n6147) );
  NAND2_X2 U5236 ( .A1(n5610), .A2(n6147), .ZN(n6143) );
  NAND2_X1 U5237 ( .A1(n6133), .A2(REIP_REG_31__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U5238 ( .A1(n6148), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4216)
         );
  OAI211_X1 U5239 ( .C1(n6143), .C2(n4217), .A(n5658), .B(n4216), .ZN(n4218)
         );
  INV_X1 U5240 ( .A(n4218), .ZN(n4219) );
  OAI211_X1 U5241 ( .C1(n5663), .C2(n6145), .A(n4220), .B(n4219), .ZN(U2955)
         );
  XNOR2_X1 U5242 ( .A(n4223), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5681)
         );
  INV_X1 U5243 ( .A(n4224), .ZN(n4270) );
  INV_X1 U5244 ( .A(n4234), .ZN(n4226) );
  NAND2_X1 U5245 ( .A1(n2988), .A2(n6138), .ZN(n4231) );
  AND2_X1 U5246 ( .A1(n6133), .A2(REIP_REG_29__SCAN_IN), .ZN(n5676) );
  AOI21_X1 U5247 ( .B1(n6148), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5676), 
        .ZN(n4228) );
  OAI21_X1 U5248 ( .B1(n6143), .B2(n4287), .A(n4228), .ZN(n4229) );
  INV_X1 U5249 ( .A(n4229), .ZN(n4230) );
  OAI211_X1 U5250 ( .C1(n5681), .C2(n6145), .A(n4231), .B(n4230), .ZN(U2957)
         );
  XNOR2_X1 U5251 ( .A(n4234), .B(n4233), .ZN(n5536) );
  AND2_X1 U5252 ( .A1(n4580), .A2(n4371), .ZN(n4762) );
  AND2_X1 U5253 ( .A1(n4762), .A2(n4511), .ZN(n4317) );
  OAI21_X1 U5254 ( .B1(n4317), .B2(n5359), .A(n4235), .ZN(n4243) );
  NAND2_X1 U5255 ( .A1(n3290), .A2(n3295), .ZN(n4236) );
  NAND2_X1 U5256 ( .A1(n6592), .A2(n4236), .ZN(n4239) );
  NAND2_X1 U5257 ( .A1(n3290), .A2(n3192), .ZN(n4377) );
  OR2_X1 U5258 ( .A1(n4377), .A2(n4237), .ZN(n4238) );
  NAND2_X1 U5259 ( .A1(n4239), .A2(n4238), .ZN(n4314) );
  INV_X1 U5260 ( .A(n5339), .ZN(n4509) );
  NAND2_X1 U5261 ( .A1(n4509), .A2(n4501), .ZN(n4242) );
  NAND2_X1 U5262 ( .A1(n4240), .A2(n3904), .ZN(n4241) );
  NOR2_X1 U5263 ( .A1(n4344), .A2(n4615), .ZN(n4499) );
  NAND2_X1 U5264 ( .A1(n4530), .A2(n4499), .ZN(n4527) );
  NAND3_X1 U5265 ( .A1(n4246), .A2(n3005), .A3(n3296), .ZN(n4372) );
  INV_X1 U5266 ( .A(n4372), .ZN(n4248) );
  NAND3_X1 U5267 ( .A1(n3030), .A2(n4248), .A3(n4989), .ZN(n4249) );
  INV_X1 U5268 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5876) );
  NAND2_X1 U5269 ( .A1(n4250), .A2(n5876), .ZN(n4253) );
  NAND2_X1 U5270 ( .A1(n4296), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4251) );
  OAI211_X1 U5271 ( .C1(n5358), .C2(EBX_REG_27__SCAN_IN), .A(n3919), .B(n4251), 
        .ZN(n4252) );
  AND2_X1 U5272 ( .A1(n4253), .A2(n4252), .ZN(n5692) );
  NAND2_X1 U5273 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n5358), .ZN(n4255) );
  MUX2_X1 U5274 ( .A(n4294), .B(n3919), .S(EBX_REG_28__SCAN_IN), .Z(n4254) );
  AND2_X1 U5275 ( .A1(n4255), .A2(n4254), .ZN(n4276) );
  OR2_X1 U5276 ( .A1(n5359), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4257)
         );
  INV_X1 U5277 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U5278 ( .A1(n4989), .A2(n5435), .ZN(n4256) );
  NAND2_X1 U5279 ( .A1(n4257), .A2(n4256), .ZN(n4299) );
  NAND2_X1 U5280 ( .A1(n5359), .A2(EBX_REG_30__SCAN_IN), .ZN(n4260) );
  NAND2_X1 U5281 ( .A1(n5358), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4259) );
  NAND2_X1 U5282 ( .A1(n4260), .A2(n4259), .ZN(n5356) );
  OAI211_X1 U5283 ( .C1(n4297), .C2(n2986), .A(n5355), .B(n5356), .ZN(n4265)
         );
  NAND2_X1 U5284 ( .A1(n2986), .A2(n3904), .ZN(n4262) );
  INV_X1 U5285 ( .A(n5356), .ZN(n4261) );
  NAND2_X1 U5286 ( .A1(n4262), .A2(n4261), .ZN(n4263) );
  OR2_X1 U5287 ( .A1(n4297), .A2(n4263), .ZN(n4264) );
  INV_X2 U5288 ( .A(n6081), .ZN(n5503) );
  NAND2_X1 U5289 ( .A1(n5485), .A2(EBX_REG_30__SCAN_IN), .ZN(n4266) );
  NOR2_X1 U5290 ( .A1(n4274), .A2(n5392), .ZN(n5813) );
  NAND2_X1 U5291 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5813), .ZN(n4291) );
  OAI22_X1 U5292 ( .A1(n5543), .A2(n5856), .B1(REIP_REG_28__SCAN_IN), .B2(
        n4291), .ZN(n4275) );
  NAND2_X1 U5293 ( .A1(n5695), .A2(n4276), .ZN(n4277) );
  NAND2_X1 U5294 ( .A1(n2986), .A2(n4277), .ZN(n5682) );
  NAND2_X1 U5295 ( .A1(REIP_REG_27__SCAN_IN), .A2(REIP_REG_28__SCAN_IN), .ZN(
        n4278) );
  OAI21_X1 U5296 ( .B1(n5814), .B2(n4278), .A(n5864), .ZN(n5371) );
  INV_X1 U5297 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6662) );
  AOI22_X1 U5298 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n6062), .B1(n5544), 
        .B2(n6071), .ZN(n4279) );
  OAI21_X1 U5299 ( .B1(n5371), .B2(n6662), .A(n4279), .ZN(n4281) );
  AND2_X1 U5300 ( .A1(n6050), .A2(EBX_REG_28__SCAN_IN), .ZN(n4280) );
  INV_X1 U5301 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6741) );
  OAI22_X1 U5302 ( .A1(n4287), .A2(n6047), .B1(n6741), .B2(n5371), .ZN(n4288)
         );
  INV_X1 U5303 ( .A(n4288), .ZN(n4290) );
  AOI22_X1 U5304 ( .A1(EBX_REG_29__SCAN_IN), .A2(n6050), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6062), .ZN(n4289) );
  NAND2_X1 U5305 ( .A1(n5378), .A2(n6741), .ZN(n5370) );
  OR2_X1 U5306 ( .A1(n4294), .A2(EBX_REG_29__SCAN_IN), .ZN(n4298) );
  NOR2_X1 U5307 ( .A1(n2986), .A2(n4298), .ZN(n4295) );
  AOI21_X1 U5308 ( .B1(n4297), .B2(n4296), .A(n4295), .ZN(n5357) );
  OAI211_X1 U5309 ( .C1(n3904), .C2(n4299), .A(n2986), .B(n4298), .ZN(n4300)
         );
  NAND2_X1 U5310 ( .A1(n5357), .A2(n4300), .ZN(n5674) );
  NOR2_X1 U5311 ( .A1(n6587), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4307) );
  AOI21_X1 U5312 ( .B1(n4304), .B2(MEMORYFETCH_REG_SCAN_IN), .A(n4307), .ZN(
        n4305) );
  NAND2_X1 U5313 ( .A1(n4306), .A2(n4305), .ZN(U2788) );
  OR2_X1 U5314 ( .A1(n3314), .A2(n4762), .ZN(n5962) );
  OAI21_X1 U5315 ( .B1(n4307), .B2(READREQUEST_REG_SCAN_IN), .A(n4309), .ZN(
        n4308) );
  OAI21_X1 U5316 ( .B1(n4309), .B2(n5962), .A(n4308), .ZN(U3474) );
  NOR2_X1 U5317 ( .A1(n6450), .A2(n4615), .ZN(n4528) );
  INV_X1 U5318 ( .A(n4528), .ZN(n4351) );
  INV_X1 U5319 ( .A(n4310), .ZN(n4311) );
  OR2_X1 U5320 ( .A1(n4312), .A2(n4311), .ZN(n4520) );
  INV_X1 U5321 ( .A(READY_N), .ZN(n6658) );
  OAI21_X1 U5322 ( .B1(n4989), .B2(n4502), .A(n6658), .ZN(n4313) );
  AOI21_X1 U5323 ( .B1(n4351), .B2(n4520), .A(n4313), .ZN(n4320) );
  INV_X1 U5324 ( .A(n4314), .ZN(n4315) );
  OR2_X1 U5325 ( .A1(n4323), .A2(n4315), .ZN(n4316) );
  NAND2_X1 U5326 ( .A1(n4316), .A2(n6450), .ZN(n4504) );
  INV_X1 U5327 ( .A(n4317), .ZN(n4318) );
  NAND2_X1 U5328 ( .A1(n4504), .A2(n4318), .ZN(n4319) );
  AOI21_X1 U5329 ( .B1(n6453), .B2(n4320), .A(n4319), .ZN(n4321) );
  NAND2_X1 U5330 ( .A1(n4322), .A2(n4321), .ZN(n4327) );
  NOR2_X1 U5331 ( .A1(n4323), .A2(n3298), .ZN(n4517) );
  NAND2_X1 U5332 ( .A1(n6453), .A2(n4517), .ZN(n4326) );
  INV_X1 U5333 ( .A(n4324), .ZN(n4330) );
  NOR2_X1 U5334 ( .A1(READY_N), .A2(n6448), .ZN(n4500) );
  NAND2_X1 U5335 ( .A1(n4330), .A2(n4500), .ZN(n4325) );
  NAND2_X1 U5336 ( .A1(n4326), .A2(n4325), .ZN(n4375) );
  NOR2_X1 U5337 ( .A1(n4327), .A2(n4375), .ZN(n4426) );
  INV_X1 U5338 ( .A(n4426), .ZN(n6435) );
  NAND2_X1 U5339 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4433) );
  OR2_X1 U5340 ( .A1(n6474), .A2(n4433), .ZN(n6559) );
  INV_X1 U5341 ( .A(n6559), .ZN(n4430) );
  AOI22_X1 U5342 ( .A1(n6435), .A2(n4506), .B1(FLUSH_REG_SCAN_IN), .B2(n4430), 
        .ZN(n4332) );
  NAND2_X1 U5343 ( .A1(n6474), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6560) );
  NAND2_X1 U5344 ( .A1(n4332), .A2(n6560), .ZN(n5808) );
  INV_X1 U5345 ( .A(n5008), .ZN(n5135) );
  NOR2_X1 U5346 ( .A1(n3444), .A2(n5135), .ZN(n4329) );
  XNOR2_X1 U5347 ( .A(n4329), .B(n4328), .ZN(n6048) );
  NAND4_X1 U5348 ( .A1(n6048), .A2(n4330), .A3(n6562), .A4(n4419), .ZN(n4331)
         );
  OAI22_X1 U5349 ( .A1(n5808), .A2(n4328), .B1(n4332), .B2(n4331), .ZN(U3455)
         );
  INV_X1 U5350 ( .A(n3428), .ZN(n6315) );
  AND4_X1 U5351 ( .A1(n4324), .A2(n4531), .A3(n4520), .A4(n4373), .ZN(n4334)
         );
  NAND2_X1 U5352 ( .A1(n4530), .A2(n4334), .ZN(n4416) );
  NOR2_X1 U5353 ( .A1(n4344), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4335)
         );
  AOI21_X1 U5354 ( .B1(n6315), .B2(n4416), .A(n4335), .ZN(n6433) );
  INV_X1 U5355 ( .A(n4346), .ZN(n5806) );
  INV_X1 U5356 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6227) );
  AOI22_X1 U5357 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6227), .B1(n4333), .B2(
        n5327), .ZN(n4336) );
  OAI21_X1 U5358 ( .B1(n6433), .B2(n5806), .A(n4336), .ZN(n4337) );
  AND2_X1 U5359 ( .A1(n4528), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6431)
         );
  AOI22_X1 U5360 ( .A1(n5808), .A2(n4337), .B1(n4346), .B2(n6431), .ZN(n4338)
         );
  OAI21_X1 U5361 ( .B1(n4333), .B2(n5808), .A(n4338), .ZN(U3461) );
  INV_X1 U5362 ( .A(n5808), .ZN(n5335) );
  NOR2_X1 U5363 ( .A1(n4340), .A2(n4339), .ZN(n4345) );
  INV_X1 U5364 ( .A(n4345), .ZN(n4348) );
  NOR2_X1 U5365 ( .A1(n4419), .A2(n6227), .ZN(n5333) );
  INV_X1 U5366 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4341) );
  AOI22_X1 U5367 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n4341), .B2(n6214), .ZN(n5332)
         );
  INV_X1 U5368 ( .A(n5332), .ZN(n4347) );
  NAND2_X1 U5369 ( .A1(n4763), .A2(n4416), .ZN(n4343) );
  NAND2_X1 U5370 ( .A1(n4528), .A2(n3088), .ZN(n4410) );
  OAI211_X1 U5371 ( .C1(n4345), .C2(n4344), .A(n4343), .B(n4410), .ZN(n6434)
         );
  AOI222_X1 U5372 ( .A1(n4348), .A2(n5327), .B1(n5333), .B2(n4347), .C1(n6434), 
        .C2(n4346), .ZN(n4350) );
  NAND2_X1 U5373 ( .A1(n5335), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4349) );
  OAI21_X1 U5374 ( .B1(n5335), .B2(n4350), .A(n4349), .ZN(U3460) );
  INV_X1 U5375 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4354) );
  OAI21_X1 U5376 ( .B1(n4351), .B2(n4514), .A(n4445), .ZN(n4352) );
  NAND2_X1 U5377 ( .A1(n6097), .A2(n3295), .ZN(n4475) );
  OR2_X1 U5378 ( .A1(n4433), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6588) );
  AOI22_X1 U5379 ( .A1(n6129), .A2(UWORD_REG_9__SCAN_IN), .B1(n6128), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4353) );
  OAI21_X1 U5380 ( .B1(n4354), .B2(n4475), .A(n4353), .ZN(U2898) );
  INV_X1 U5381 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4356) );
  AOI22_X1 U5382 ( .A1(n6129), .A2(UWORD_REG_10__SCAN_IN), .B1(n6128), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4355) );
  OAI21_X1 U5383 ( .B1(n4356), .B2(n4475), .A(n4355), .ZN(U2897) );
  INV_X1 U5384 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4358) );
  AOI22_X1 U5385 ( .A1(n6129), .A2(UWORD_REG_11__SCAN_IN), .B1(n6128), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4357) );
  OAI21_X1 U5386 ( .B1(n4358), .B2(n4475), .A(n4357), .ZN(U2896) );
  INV_X1 U5387 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4360) );
  AOI22_X1 U5388 ( .A1(n6129), .A2(UWORD_REG_12__SCAN_IN), .B1(n6128), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4359) );
  OAI21_X1 U5389 ( .B1(n4360), .B2(n4475), .A(n4359), .ZN(U2895) );
  INV_X1 U5390 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4362) );
  AOI22_X1 U5391 ( .A1(n6129), .A2(UWORD_REG_13__SCAN_IN), .B1(n6128), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4361) );
  OAI21_X1 U5392 ( .B1(n4362), .B2(n4475), .A(n4361), .ZN(U2894) );
  INV_X1 U5393 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4364) );
  AOI22_X1 U5394 ( .A1(n6129), .A2(UWORD_REG_8__SCAN_IN), .B1(n6128), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4363) );
  OAI21_X1 U5395 ( .B1(n4364), .B2(n4475), .A(n4363), .ZN(U2899) );
  INV_X1 U5396 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4366) );
  AOI22_X1 U5397 ( .A1(n6129), .A2(UWORD_REG_14__SCAN_IN), .B1(n6128), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4365) );
  OAI21_X1 U5398 ( .B1(n4366), .B2(n4475), .A(n4365), .ZN(U2893) );
  OAI21_X1 U5399 ( .B1(n4369), .B2(n4368), .A(n4367), .ZN(n6151) );
  NOR2_X1 U5400 ( .A1(n4373), .A2(n4372), .ZN(n4374) );
  INV_X1 U5401 ( .A(n4377), .ZN(n4378) );
  INV_X1 U5402 ( .A(DATAI_0_), .ZN(n6749) );
  INV_X1 U5403 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6132) );
  OAI222_X1 U5404 ( .A1(n6151), .A2(n5524), .B1(n5299), .B2(n6749), .C1(n5507), 
        .C2(n6132), .ZN(U2891) );
  OR2_X1 U5405 ( .A1(n4380), .A2(n4379), .ZN(n4381) );
  NAND2_X1 U5406 ( .A1(n4382), .A2(n4381), .ZN(n4993) );
  INV_X1 U5407 ( .A(DATAI_1_), .ZN(n4614) );
  INV_X1 U5408 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6127) );
  OAI222_X1 U5409 ( .A1(n4993), .A2(n5524), .B1(n5299), .B2(n4614), .C1(n5507), 
        .C2(n6127), .ZN(U2890) );
  NOR2_X1 U5410 ( .A1(n4384), .A2(n4385), .ZN(n4386) );
  NOR2_X1 U5411 ( .A1(n4383), .A2(n4386), .ZN(n6139) );
  INV_X1 U5412 ( .A(n6139), .ZN(n4387) );
  INV_X1 U5413 ( .A(DATAI_2_), .ZN(n4488) );
  INV_X1 U5414 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6125) );
  OAI222_X1 U5415 ( .A1(n4387), .A2(n5524), .B1(n5299), .B2(n4488), .C1(n5507), 
        .C2(n6125), .ZN(U2889) );
  OAI21_X1 U5416 ( .B1(n4383), .B2(n4389), .A(n4388), .ZN(n5353) );
  INV_X1 U5417 ( .A(DATAI_3_), .ZN(n4584) );
  INV_X1 U5418 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6123) );
  OAI222_X1 U5419 ( .A1(n5353), .A2(n5524), .B1(n5299), .B2(n4584), .C1(n5507), 
        .C2(n6123), .ZN(U2888) );
  INV_X1 U5420 ( .A(n4517), .ZN(n4391) );
  NAND2_X1 U5421 ( .A1(n4527), .A2(n4391), .ZN(n4409) );
  INV_X1 U5422 ( .A(n4393), .ZN(n4399) );
  INV_X1 U5423 ( .A(n4397), .ZN(n4394) );
  OAI211_X1 U5424 ( .C1(n4392), .C2(n4399), .A(n4395), .B(n4394), .ZN(n4396)
         );
  NAND2_X1 U5425 ( .A1(n4409), .A2(n4396), .ZN(n4404) );
  NAND2_X1 U5426 ( .A1(n4397), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4398) );
  NAND2_X1 U5427 ( .A1(n4399), .A2(n4398), .ZN(n4402) );
  OAI21_X1 U5428 ( .B1(n3354), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n4400), 
        .ZN(n5805) );
  NOR2_X1 U5429 ( .A1(n4529), .A2(n5805), .ZN(n4401) );
  AOI21_X1 U5430 ( .B1(n4528), .B2(n4402), .A(n4401), .ZN(n4403) );
  OAI211_X1 U5431 ( .C1(n4406), .C2(n4410), .A(n4404), .B(n4403), .ZN(n4405)
         );
  AOI21_X1 U5432 ( .B1(n3017), .B2(n4416), .A(n4405), .ZN(n5807) );
  MUX2_X1 U5433 ( .A(n4406), .B(n5807), .S(n6435), .Z(n6443) );
  INV_X1 U5434 ( .A(n6443), .ZN(n4420) );
  NAND2_X1 U5435 ( .A1(n4426), .A2(n5336), .ZN(n4418) );
  INV_X1 U5436 ( .A(n4408), .ZN(n6063) );
  XNOR2_X1 U5437 ( .A(n4392), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4414)
         );
  NAND2_X1 U5438 ( .A1(n4409), .A2(n4414), .ZN(n4413) );
  NAND2_X1 U5439 ( .A1(n4528), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4411) );
  MUX2_X1 U5440 ( .A(n4411), .B(n4410), .S(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .Z(n4412) );
  OAI211_X1 U5441 ( .C1(n4414), .C2(n4529), .A(n4413), .B(n4412), .ZN(n4415)
         );
  AOI21_X1 U5442 ( .B1(n6063), .B2(n4416), .A(n4415), .ZN(n5329) );
  NAND2_X1 U5443 ( .A1(n6435), .A2(n5329), .ZN(n4417) );
  NAND3_X1 U5444 ( .A1(n4420), .A2(n6442), .A3(n4419), .ZN(n4424) );
  INV_X1 U5445 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6755) );
  AND2_X1 U5446 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6755), .ZN(n4421) );
  NAND2_X1 U5447 ( .A1(n4422), .A2(n4421), .ZN(n4423) );
  NAND2_X1 U5448 ( .A1(n4424), .A2(n4423), .ZN(n6460) );
  INV_X1 U5449 ( .A(n3095), .ZN(n4425) );
  NAND2_X1 U5450 ( .A1(n6460), .A2(n4425), .ZN(n4435) );
  MUX2_X1 U5451 ( .A(n4426), .B(n6755), .S(STATE2_REG_1__SCAN_IN), .Z(n4429)
         );
  NOR2_X1 U5452 ( .A1(n4324), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4427) );
  AND2_X1 U5453 ( .A1(n6048), .A2(n4427), .ZN(n4428) );
  AOI21_X1 U5454 ( .B1(n4429), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n4428), 
        .ZN(n6458) );
  NAND3_X1 U5455 ( .A1(n4435), .A2(n6458), .A3(n6755), .ZN(n4431) );
  NAND2_X1 U5456 ( .A1(n4431), .A2(n4430), .ZN(n4432) );
  NAND2_X1 U5457 ( .A1(n4432), .A2(n4667), .ZN(n6570) );
  INV_X1 U5458 ( .A(n4433), .ZN(n4434) );
  AND3_X1 U5459 ( .A1(n4435), .A2(n6458), .A3(n4434), .ZN(n6468) );
  NAND2_X1 U5460 ( .A1(n6562), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6567) );
  INV_X1 U5461 ( .A(n6567), .ZN(n5802) );
  OAI22_X1 U5462 ( .A1(n4853), .A2(n6587), .B1(n3428), .B2(n5802), .ZN(n4436)
         );
  OAI21_X1 U5463 ( .B1(n6468), .B2(n4436), .A(n6570), .ZN(n4437) );
  OAI21_X1 U5464 ( .B1(n6570), .B2(n6430), .A(n4437), .ZN(U3465) );
  INV_X1 U5465 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4761) );
  NAND2_X1 U5466 ( .A1(n6133), .A2(REIP_REG_1__SCAN_IN), .ZN(n6207) );
  OAI21_X1 U5467 ( .B1(n5610), .B2(n4761), .A(n6207), .ZN(n4442) );
  OAI21_X1 U5468 ( .B1(n4440), .B2(n4439), .A(n4438), .ZN(n6205) );
  NOR2_X1 U5469 ( .A1(n6205), .A2(n6145), .ZN(n4441) );
  AOI211_X1 U5470 ( .C1(n4761), .C2(n5613), .A(n4442), .B(n4441), .ZN(n4443)
         );
  OAI21_X1 U5471 ( .B1(n6371), .B2(n4993), .A(n4443), .ZN(U2985) );
  INV_X1 U5472 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4447) );
  INV_X2 U5473 ( .A(n4445), .ZN(n4657) );
  OR2_X1 U5474 ( .A1(n4657), .A2(n4444), .ZN(n4625) );
  INV_X1 U5475 ( .A(DATAI_15_), .ZN(n6764) );
  INV_X1 U5476 ( .A(EAX_REG_15__SCAN_IN), .ZN(n4446) );
  OAI222_X1 U5477 ( .A1(n4447), .A2(n4625), .B1(n4607), .B2(n6764), .C1(n4446), 
        .C2(n4445), .ZN(U2954) );
  AND2_X1 U5478 ( .A1(n4448), .A2(n4449), .ZN(n4451) );
  OR2_X1 U5479 ( .A1(n4451), .A2(n4450), .ZN(n4881) );
  INV_X1 U5480 ( .A(DATAI_5_), .ZN(n6770) );
  INV_X1 U5481 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6118) );
  OAI222_X1 U5482 ( .A1(n4881), .A2(n5524), .B1(n5299), .B2(n6770), .C1(n5507), 
        .C2(n6118), .ZN(U2886) );
  OAI21_X1 U5483 ( .B1(n4450), .B2(n4453), .A(n4914), .ZN(n4693) );
  INV_X1 U5484 ( .A(DATAI_6_), .ZN(n4609) );
  INV_X1 U5485 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6116) );
  OAI222_X1 U5486 ( .A1(n4693), .A2(n5524), .B1(n5299), .B2(n4609), .C1(n5507), 
        .C2(n6116), .ZN(U2885) );
  XNOR2_X1 U5487 ( .A(n4454), .B(n4455), .ZN(n6182) );
  INV_X1 U5488 ( .A(n5353), .ZN(n4458) );
  NAND2_X1 U5489 ( .A1(n6148), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4456)
         );
  NAND2_X1 U5490 ( .A1(n6133), .A2(REIP_REG_3__SCAN_IN), .ZN(n6179) );
  OAI211_X1 U5491 ( .C1(n6143), .C2(n5344), .A(n4456), .B(n6179), .ZN(n4457)
         );
  AOI21_X1 U5492 ( .B1(n4458), .B2(n6138), .A(n4457), .ZN(n4459) );
  OAI21_X1 U5493 ( .B1(n6145), .B2(n6182), .A(n4459), .ZN(U2983) );
  INV_X1 U5494 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4461) );
  INV_X2 U5495 ( .A(n6588), .ZN(n6129) );
  AOI22_X1 U5496 ( .A1(n6129), .A2(UWORD_REG_2__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4460) );
  OAI21_X1 U5497 ( .B1(n4461), .B2(n4475), .A(n4460), .ZN(U2905) );
  INV_X1 U5498 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4463) );
  AOI22_X1 U5499 ( .A1(n6129), .A2(UWORD_REG_3__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4462) );
  OAI21_X1 U5500 ( .B1(n4463), .B2(n4475), .A(n4462), .ZN(U2904) );
  INV_X1 U5501 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4465) );
  AOI22_X1 U5502 ( .A1(n6129), .A2(UWORD_REG_6__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4464) );
  OAI21_X1 U5503 ( .B1(n4465), .B2(n4475), .A(n4464), .ZN(U2901) );
  INV_X1 U5504 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4467) );
  AOI22_X1 U5505 ( .A1(n6129), .A2(UWORD_REG_5__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4466) );
  OAI21_X1 U5506 ( .B1(n4467), .B2(n4475), .A(n4466), .ZN(U2902) );
  INV_X1 U5507 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4469) );
  AOI22_X1 U5508 ( .A1(n6129), .A2(UWORD_REG_4__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4468) );
  OAI21_X1 U5509 ( .B1(n4469), .B2(n4475), .A(n4468), .ZN(U2903) );
  INV_X1 U5510 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4471) );
  AOI22_X1 U5511 ( .A1(n6129), .A2(UWORD_REG_7__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4470) );
  OAI21_X1 U5512 ( .B1(n4471), .B2(n4475), .A(n4470), .ZN(U2900) );
  INV_X1 U5513 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4473) );
  AOI22_X1 U5514 ( .A1(n6129), .A2(UWORD_REG_1__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4472) );
  OAI21_X1 U5515 ( .B1(n4473), .B2(n4475), .A(n4472), .ZN(U2906) );
  INV_X1 U5516 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4476) );
  AOI22_X1 U5517 ( .A1(n6129), .A2(UWORD_REG_0__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4474) );
  OAI21_X1 U5518 ( .B1(n4476), .B2(n4475), .A(n4474), .ZN(U2907) );
  INV_X1 U5519 ( .A(n4479), .ZN(n4480) );
  NOR2_X1 U5520 ( .A1(n4482), .A2(n6730), .ZN(n4483) );
  AOI21_X1 U5521 ( .B1(n6281), .B2(n4483), .A(n6587), .ZN(n4495) );
  NOR2_X1 U5522 ( .A1(n4408), .A2(n4763), .ZN(n5136) );
  NAND3_X1 U5523 ( .A1(n5136), .A2(n5135), .A3(n6315), .ZN(n4485) );
  NAND2_X1 U5524 ( .A1(n6437), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4940) );
  OR2_X1 U5525 ( .A1(n4940), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5126)
         );
  NOR2_X1 U5526 ( .A1(n6430), .A2(n5126), .ZN(n4671) );
  INV_X1 U5527 ( .A(n4671), .ZN(n4484) );
  AND2_X1 U5528 ( .A1(n4485), .A2(n4484), .ZN(n4494) );
  INV_X1 U5529 ( .A(n4494), .ZN(n4487) );
  INV_X1 U5530 ( .A(n5126), .ZN(n4486) );
  AOI22_X1 U5531 ( .A1(n4495), .A2(n4487), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4486), .ZN(n4675) );
  NOR2_X2 U5532 ( .A1(n4668), .A2(n4511), .ZN(n6390) );
  INV_X1 U5533 ( .A(DATAI_26_), .ZN(n4490) );
  OR2_X1 U5534 ( .A1(n6371), .A2(n4490), .ZN(n6248) );
  INV_X1 U5535 ( .A(n6281), .ZN(n4491) );
  INV_X1 U5536 ( .A(DATAI_18_), .ZN(n6768) );
  OR2_X1 U5537 ( .A1(n6371), .A2(n6768), .ZN(n6394) );
  OAI22_X1 U5538 ( .A1(n6248), .A2(n5166), .B1(n5047), .B2(n6394), .ZN(n4493)
         );
  AOI21_X1 U5539 ( .B1(n6390), .B2(n4671), .A(n4493), .ZN(n4498) );
  OAI21_X1 U5540 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6562), .A(n5132), 
        .ZN(n4575) );
  AOI22_X1 U5541 ( .A1(n4495), .A2(n4494), .B1(n5126), .B2(n6587), .ZN(n4496)
         );
  NAND2_X1 U5542 ( .A1(n6377), .A2(n4496), .ZN(n4672) );
  NAND2_X1 U5543 ( .A1(n4672), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4497) );
  OAI211_X1 U5544 ( .C1(n4675), .C2(n6336), .A(n4498), .B(n4497), .ZN(U3062)
         );
  INV_X1 U5545 ( .A(n4499), .ZN(n4505) );
  OAI211_X1 U5546 ( .C1(n4615), .C2(n4502), .A(n4501), .B(n4500), .ZN(n4503)
         );
  OAI211_X1 U5547 ( .C1(n6453), .C2(n4505), .A(n4504), .B(n4503), .ZN(n4507)
         );
  NAND2_X1 U5548 ( .A1(n4507), .A2(n4506), .ZN(n4516) );
  NAND2_X1 U5549 ( .A1(n4508), .A2(n6658), .ZN(n4510) );
  OAI211_X1 U5550 ( .C1(n4520), .C2(n4510), .A(n3295), .B(n4509), .ZN(n4512)
         );
  NAND2_X1 U5551 ( .A1(n4512), .A2(n4511), .ZN(n4513) );
  INV_X1 U5552 ( .A(n6457), .ZN(n4518) );
  OR2_X1 U5553 ( .A1(n4518), .A2(n4517), .ZN(n6447) );
  INV_X1 U5554 ( .A(n6447), .ZN(n4523) );
  OAI22_X1 U5555 ( .A1(n4520), .A2(n5358), .B1(n4519), .B2(n3005), .ZN(n4521)
         );
  INV_X1 U5556 ( .A(n4521), .ZN(n4522) );
  NAND3_X1 U5557 ( .A1(n4523), .A2(n4522), .A3(n4324), .ZN(n4524) );
  XNOR2_X1 U5558 ( .A(n4525), .B(n4526), .ZN(n4571) );
  INV_X1 U5559 ( .A(n4527), .ZN(n6454) );
  INV_X1 U5560 ( .A(n5929), .ZN(n6193) );
  AOI21_X1 U5561 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6195) );
  NAND2_X1 U5562 ( .A1(n4536), .A2(n4528), .ZN(n6225) );
  OAI211_X1 U5563 ( .C1(n4531), .C2(n3295), .A(n4530), .B(n4529), .ZN(n4532)
         );
  NAND2_X1 U5564 ( .A1(n4536), .A2(n4532), .ZN(n5930) );
  NAND2_X1 U5565 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5070) );
  INV_X1 U5566 ( .A(n5070), .ZN(n6194) );
  NAND2_X1 U5567 ( .A1(n4533), .A2(n6190), .ZN(n6226) );
  OAI21_X1 U5568 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n5930), .A(n6226), 
        .ZN(n5284) );
  INV_X1 U5569 ( .A(n5284), .ZN(n4534) );
  OAI21_X1 U5570 ( .B1(n5280), .B2(n6194), .A(n4534), .ZN(n6197) );
  AOI21_X1 U5571 ( .B1(n6193), .B2(n6195), .A(n6197), .ZN(n6189) );
  INV_X1 U5572 ( .A(n6189), .ZN(n4545) );
  OAI21_X1 U5573 ( .B1(n4519), .B2(n3284), .A(n6465), .ZN(n4535) );
  INV_X1 U5574 ( .A(n4537), .ZN(n4554) );
  NAND2_X1 U5575 ( .A1(n4997), .A2(n4538), .ZN(n4539) );
  NAND2_X1 U5576 ( .A1(n4554), .A2(n4539), .ZN(n6060) );
  NAND2_X1 U5577 ( .A1(n6133), .A2(REIP_REG_4__SCAN_IN), .ZN(n4567) );
  INV_X1 U5578 ( .A(n6195), .ZN(n4540) );
  OAI21_X1 U5579 ( .B1(n5070), .B2(n6198), .A(n5929), .ZN(n5077) );
  NAND2_X1 U5580 ( .A1(n4540), .A2(n5077), .ZN(n6185) );
  AOI21_X1 U5581 ( .B1(n6188), .B2(n4541), .A(n6185), .ZN(n4542) );
  NAND2_X1 U5582 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4551) );
  NAND2_X1 U5583 ( .A1(n4542), .A2(n4551), .ZN(n4543) );
  OAI211_X1 U5584 ( .C1(n6218), .C2(n6060), .A(n4567), .B(n4543), .ZN(n4544)
         );
  AOI21_X1 U5585 ( .B1(n4545), .B2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4544), 
        .ZN(n4546) );
  OAI21_X1 U5586 ( .B1(n6206), .B2(n4571), .A(n4546), .ZN(U3014) );
  XNOR2_X1 U5587 ( .A(n3008), .B(n4548), .ZN(n4563) );
  INV_X1 U5588 ( .A(n6198), .ZN(n4549) );
  NAND2_X1 U5589 ( .A1(n6194), .A2(n4549), .ZN(n4550) );
  AOI211_X1 U5590 ( .C1(n4550), .C2(n5929), .A(n6195), .B(n4551), .ZN(n4553)
         );
  NOR2_X1 U5591 ( .A1(n4552), .A2(n4551), .ZN(n5069) );
  OAI21_X1 U5592 ( .B1(n5069), .B2(n5782), .A(n6189), .ZN(n4739) );
  OAI21_X1 U5593 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4553), .A(n4739), 
        .ZN(n4557) );
  AOI21_X1 U5594 ( .B1(n4555), .B2(n4554), .A(n3930), .ZN(n6036) );
  AND2_X1 U5595 ( .A1(n6133), .A2(REIP_REG_5__SCAN_IN), .ZN(n4559) );
  AOI21_X1 U5596 ( .B1(n6170), .B2(n6036), .A(n4559), .ZN(n4556) );
  OAI211_X1 U5597 ( .C1(n6206), .C2(n4563), .A(n4557), .B(n4556), .ZN(U3013)
         );
  INV_X1 U5598 ( .A(n4881), .ZN(n6041) );
  INV_X1 U5599 ( .A(n4558), .ZN(n6046) );
  AOI21_X1 U5600 ( .B1(n6148), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4559), 
        .ZN(n4560) );
  OAI21_X1 U5601 ( .B1(n6143), .B2(n6046), .A(n4560), .ZN(n4561) );
  AOI21_X1 U5602 ( .B1(n6041), .B2(n6138), .A(n4561), .ZN(n4562) );
  OAI21_X1 U5603 ( .B1(n6145), .B2(n4563), .A(n4562), .ZN(U2981) );
  INV_X1 U5604 ( .A(n4448), .ZN(n4564) );
  AOI21_X1 U5605 ( .B1(n4565), .B2(n4388), .A(n4564), .ZN(n6052) );
  INV_X1 U5606 ( .A(n6051), .ZN(n4568) );
  NAND2_X1 U5607 ( .A1(n6148), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4566)
         );
  OAI211_X1 U5608 ( .C1(n6143), .C2(n4568), .A(n4567), .B(n4566), .ZN(n4569)
         );
  AOI21_X1 U5609 ( .B1(n6052), .B2(n6138), .A(n4569), .ZN(n4570) );
  OAI21_X1 U5610 ( .B1(n6145), .B2(n4571), .A(n4570), .ZN(U2982) );
  INV_X1 U5611 ( .A(n6052), .ZN(n4926) );
  INV_X1 U5612 ( .A(DATAI_4_), .ZN(n6751) );
  INV_X1 U5613 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6121) );
  OAI222_X1 U5614 ( .A1(n4926), .A2(n5524), .B1(n5299), .B2(n6751), .C1(n5507), 
        .C2(n6121), .ZN(U2887) );
  NAND2_X1 U5615 ( .A1(n4478), .A2(n4479), .ZN(n6370) );
  NAND2_X1 U5616 ( .A1(n4854), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4942) );
  NAND2_X1 U5617 ( .A1(n4942), .A2(n6311), .ZN(n6563) );
  NAND2_X1 U5618 ( .A1(n4482), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5800) );
  INV_X1 U5619 ( .A(n5800), .ZN(n6312) );
  NAND2_X1 U5620 ( .A1(n5801), .A2(n6312), .ZN(n4572) );
  OAI21_X1 U5621 ( .B1(n6563), .B2(n4572), .A(n6568), .ZN(n4578) );
  NAND2_X1 U5622 ( .A1(n4408), .A2(n4763), .ZN(n5201) );
  NOR2_X1 U5623 ( .A1(n3017), .A2(n5201), .ZN(n4702) );
  NOR2_X1 U5624 ( .A1(n6314), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6274)
         );
  AOI21_X1 U5625 ( .B1(n4702), .B2(n6315), .A(n6274), .ZN(n4574) );
  NAND3_X1 U5626 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6572), .A3(n6441), .ZN(n4697) );
  OAI22_X1 U5627 ( .A1(n4578), .A2(n4574), .B1(n4697), .B2(n4573), .ZN(n6276)
         );
  INV_X1 U5628 ( .A(n6276), .ZN(n5005) );
  INV_X1 U5629 ( .A(n4574), .ZN(n4577) );
  AOI21_X1 U5630 ( .B1(n4697), .B2(n6587), .A(n4575), .ZN(n4576) );
  OAI21_X1 U5631 ( .B1(n4578), .B2(n4577), .A(n4576), .ZN(n6277) );
  INV_X1 U5632 ( .A(DATAI_16_), .ZN(n6765) );
  OR2_X1 U5633 ( .A1(n6371), .A2(n6765), .ZN(n6382) );
  NAND2_X1 U5634 ( .A1(n4482), .A2(n4782), .ZN(n6228) );
  INV_X1 U5635 ( .A(n6228), .ZN(n4714) );
  NAND2_X1 U5636 ( .A1(n3078), .A2(n5006), .ZN(n4930) );
  INV_X1 U5637 ( .A(DATAI_24_), .ZN(n4579) );
  OR2_X1 U5638 ( .A1(n6371), .A2(n4579), .ZN(n6242) );
  INV_X1 U5639 ( .A(n6242), .ZN(n6379) );
  NOR2_X2 U5640 ( .A1(n4668), .A2(n4580), .ZN(n6369) );
  AOI22_X1 U5641 ( .A1(n6275), .A2(n6379), .B1(n6369), .B2(n6274), .ZN(n4581)
         );
  OAI21_X1 U5642 ( .B1(n6382), .B2(n6280), .A(n4581), .ZN(n4582) );
  AOI21_X1 U5643 ( .B1(n6277), .B2(INSTQUEUE_REG_3__0__SCAN_IN), .A(n4582), 
        .ZN(n4583) );
  OAI21_X1 U5644 ( .B1(n5005), .B2(n6328), .A(n4583), .ZN(U3044) );
  INV_X1 U5645 ( .A(DATAI_19_), .ZN(n6754) );
  OR2_X1 U5646 ( .A1(n6371), .A2(n6754), .ZN(n6400) );
  INV_X1 U5647 ( .A(DATAI_27_), .ZN(n4585) );
  OR2_X1 U5648 ( .A1(n6371), .A2(n4585), .ZN(n6251) );
  INV_X1 U5649 ( .A(n6251), .ZN(n6397) );
  NOR2_X2 U5650 ( .A1(n4668), .A2(n4586), .ZN(n6396) );
  AOI22_X1 U5651 ( .A1(n6275), .A2(n6397), .B1(n6396), .B2(n6274), .ZN(n4587)
         );
  OAI21_X1 U5652 ( .B1(n6400), .B2(n6280), .A(n4587), .ZN(n4588) );
  AOI21_X1 U5653 ( .B1(n6277), .B2(INSTQUEUE_REG_3__3__SCAN_IN), .A(n4588), 
        .ZN(n4589) );
  OAI21_X1 U5654 ( .B1(n5005), .B2(n6340), .A(n4589), .ZN(U3047) );
  OAI22_X1 U5655 ( .A1(n6242), .A2(n5166), .B1(n5047), .B2(n6382), .ZN(n4590)
         );
  AOI21_X1 U5656 ( .B1(n6369), .B2(n4671), .A(n4590), .ZN(n4592) );
  NAND2_X1 U5657 ( .A1(n4672), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4591) );
  OAI211_X1 U5658 ( .C1(n4675), .C2(n6328), .A(n4592), .B(n4591), .ZN(U3060)
         );
  OAI22_X1 U5659 ( .A1(n6251), .A2(n5166), .B1(n5047), .B2(n6400), .ZN(n4593)
         );
  AOI21_X1 U5660 ( .B1(n6396), .B2(n4671), .A(n4593), .ZN(n4595) );
  NAND2_X1 U5661 ( .A1(n4672), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4594) );
  OAI211_X1 U5662 ( .C1(n4675), .C2(n6340), .A(n4595), .B(n4594), .ZN(U3063)
         );
  AOI22_X1 U5663 ( .A1(n4606), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n4657), .ZN(n4596) );
  NAND2_X1 U5664 ( .A1(n4649), .A2(DATAI_13_), .ZN(n4647) );
  NAND2_X1 U5665 ( .A1(n4596), .A2(n4647), .ZN(U2952) );
  AOI22_X1 U5666 ( .A1(n4606), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n4657), .ZN(n4597) );
  NAND2_X1 U5667 ( .A1(n4649), .A2(DATAI_6_), .ZN(n4630) );
  NAND2_X1 U5668 ( .A1(n4597), .A2(n4630), .ZN(U2930) );
  AOI22_X1 U5669 ( .A1(n4606), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n4657), .ZN(n4598) );
  NAND2_X1 U5670 ( .A1(n4649), .A2(DATAI_3_), .ZN(n4626) );
  NAND2_X1 U5671 ( .A1(n4598), .A2(n4626), .ZN(U2927) );
  AOI22_X1 U5672 ( .A1(n4606), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n4657), .ZN(n4599) );
  INV_X1 U5673 ( .A(DATAI_9_), .ZN(n5090) );
  OR2_X1 U5674 ( .A1(n4607), .A2(n5090), .ZN(n4602) );
  NAND2_X1 U5675 ( .A1(n4599), .A2(n4602), .ZN(U2933) );
  AOI22_X1 U5676 ( .A1(n4606), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n4657), .ZN(n4600) );
  NAND2_X1 U5677 ( .A1(n4649), .A2(DATAI_0_), .ZN(n4639) );
  NAND2_X1 U5678 ( .A1(n4600), .A2(n4639), .ZN(U2924) );
  AOI22_X1 U5679 ( .A1(n4606), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n4657), .ZN(n4601) );
  NAND2_X1 U5680 ( .A1(n4649), .A2(DATAI_10_), .ZN(n4628) );
  NAND2_X1 U5681 ( .A1(n4601), .A2(n4628), .ZN(U2949) );
  AOI22_X1 U5682 ( .A1(n4606), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n4657), .ZN(n4603) );
  NAND2_X1 U5683 ( .A1(n4603), .A2(n4602), .ZN(U2948) );
  AOI22_X1 U5684 ( .A1(n4606), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n4657), .ZN(n4604) );
  NAND2_X1 U5685 ( .A1(n4649), .A2(DATAI_12_), .ZN(n4637) );
  NAND2_X1 U5686 ( .A1(n4604), .A2(n4637), .ZN(U2951) );
  AOI22_X1 U5687 ( .A1(n4606), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n4657), .ZN(n4605) );
  NAND2_X1 U5688 ( .A1(n4649), .A2(DATAI_14_), .ZN(n4641) );
  NAND2_X1 U5689 ( .A1(n4605), .A2(n4641), .ZN(U2953) );
  AOI22_X1 U5690 ( .A1(n4606), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n4657), .ZN(n4608) );
  INV_X1 U5691 ( .A(DATAI_11_), .ZN(n5182) );
  OR2_X1 U5692 ( .A1(n4607), .A2(n5182), .ZN(n4635) );
  NAND2_X1 U5693 ( .A1(n4608), .A2(n4635), .ZN(U2950) );
  NOR2_X2 U5694 ( .A1(n4668), .A2(n3006), .ZN(n6414) );
  INV_X1 U5695 ( .A(DATAI_30_), .ZN(n4610) );
  OR2_X1 U5696 ( .A1(n6371), .A2(n4610), .ZN(n6260) );
  INV_X1 U5697 ( .A(DATAI_22_), .ZN(n6771) );
  OR2_X1 U5698 ( .A1(n6371), .A2(n6771), .ZN(n6418) );
  OAI22_X1 U5699 ( .A1(n6260), .A2(n5166), .B1(n5047), .B2(n6418), .ZN(n4611)
         );
  AOI21_X1 U5700 ( .B1(n6414), .B2(n4671), .A(n4611), .ZN(n4613) );
  NAND2_X1 U5701 ( .A1(n4672), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4612) );
  OAI211_X1 U5702 ( .C1(n4675), .C2(n6352), .A(n4613), .B(n4612), .ZN(U3066)
         );
  NOR2_X2 U5703 ( .A1(n4668), .A2(n4615), .ZN(n6384) );
  INV_X1 U5704 ( .A(DATAI_25_), .ZN(n4616) );
  OR2_X1 U5705 ( .A1(n6371), .A2(n4616), .ZN(n6245) );
  INV_X1 U5706 ( .A(DATAI_17_), .ZN(n6739) );
  OR2_X1 U5707 ( .A1(n6371), .A2(n6739), .ZN(n6388) );
  OAI22_X1 U5708 ( .A1(n6245), .A2(n5166), .B1(n5047), .B2(n6388), .ZN(n4617)
         );
  AOI21_X1 U5709 ( .B1(n6384), .B2(n4671), .A(n4617), .ZN(n4619) );
  NAND2_X1 U5710 ( .A1(n4672), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4618) );
  OAI211_X1 U5711 ( .C1(n4675), .C2(n6332), .A(n4619), .B(n4618), .ZN(U3061)
         );
  NOR2_X2 U5712 ( .A1(n4668), .A2(n3005), .ZN(n6402) );
  INV_X1 U5713 ( .A(DATAI_28_), .ZN(n4621) );
  OR2_X1 U5714 ( .A1(n6371), .A2(n4621), .ZN(n6254) );
  INV_X1 U5715 ( .A(DATAI_20_), .ZN(n6727) );
  OR2_X1 U5716 ( .A1(n6371), .A2(n6727), .ZN(n6406) );
  OAI22_X1 U5717 ( .A1(n6254), .A2(n5166), .B1(n5047), .B2(n6406), .ZN(n4622)
         );
  AOI21_X1 U5718 ( .B1(n6402), .B2(n4671), .A(n4622), .ZN(n4624) );
  NAND2_X1 U5719 ( .A1(n4672), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4623) );
  OAI211_X1 U5720 ( .C1(n4675), .C2(n6344), .A(n4624), .B(n4623), .ZN(U3064)
         );
  AOI22_X1 U5721 ( .A1(n4660), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n4657), .ZN(n4627) );
  NAND2_X1 U5722 ( .A1(n4627), .A2(n4626), .ZN(U2942) );
  AOI22_X1 U5723 ( .A1(n4660), .A2(UWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_26__SCAN_IN), .B2(n4657), .ZN(n4629) );
  NAND2_X1 U5724 ( .A1(n4629), .A2(n4628), .ZN(U2934) );
  AOI22_X1 U5725 ( .A1(n4660), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n4657), .ZN(n4631) );
  NAND2_X1 U5726 ( .A1(n4631), .A2(n4630), .ZN(U2945) );
  AOI22_X1 U5727 ( .A1(n4660), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n4657), .ZN(n4632) );
  NAND2_X1 U5728 ( .A1(n4649), .A2(DATAI_7_), .ZN(n4658) );
  NAND2_X1 U5729 ( .A1(n4632), .A2(n4658), .ZN(U2946) );
  AOI22_X1 U5730 ( .A1(n4660), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n4657), .ZN(n4633) );
  NAND2_X1 U5731 ( .A1(n4649), .A2(DATAI_1_), .ZN(n4651) );
  NAND2_X1 U5732 ( .A1(n4633), .A2(n4651), .ZN(U2940) );
  AOI22_X1 U5733 ( .A1(n4660), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n4657), .ZN(n4634) );
  NAND2_X1 U5734 ( .A1(n4649), .A2(DATAI_2_), .ZN(n4653) );
  NAND2_X1 U5735 ( .A1(n4634), .A2(n4653), .ZN(U2941) );
  AOI22_X1 U5736 ( .A1(n4660), .A2(UWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_27__SCAN_IN), .B2(n4657), .ZN(n4636) );
  NAND2_X1 U5737 ( .A1(n4636), .A2(n4635), .ZN(U2935) );
  AOI22_X1 U5738 ( .A1(n4660), .A2(UWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_28__SCAN_IN), .B2(n4657), .ZN(n4638) );
  NAND2_X1 U5739 ( .A1(n4638), .A2(n4637), .ZN(U2936) );
  AOI22_X1 U5740 ( .A1(n4660), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n4657), .ZN(n4640) );
  NAND2_X1 U5741 ( .A1(n4640), .A2(n4639), .ZN(U2939) );
  AOI22_X1 U5742 ( .A1(n4660), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n4657), .ZN(n4642) );
  NAND2_X1 U5743 ( .A1(n4642), .A2(n4641), .ZN(U2938) );
  AOI22_X1 U5744 ( .A1(n4660), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n4657), .ZN(n4643) );
  NAND2_X1 U5745 ( .A1(n4649), .A2(DATAI_4_), .ZN(n4661) );
  NAND2_X1 U5746 ( .A1(n4643), .A2(n4661), .ZN(U2943) );
  AOI22_X1 U5747 ( .A1(n4660), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n4657), .ZN(n4644) );
  NAND2_X1 U5748 ( .A1(n4649), .A2(DATAI_5_), .ZN(n4645) );
  NAND2_X1 U5749 ( .A1(n4644), .A2(n4645), .ZN(U2944) );
  AOI22_X1 U5750 ( .A1(n4660), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n4657), .ZN(n4646) );
  NAND2_X1 U5751 ( .A1(n4646), .A2(n4645), .ZN(U2929) );
  AOI22_X1 U5752 ( .A1(n4660), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n4657), .ZN(n4648) );
  NAND2_X1 U5753 ( .A1(n4648), .A2(n4647), .ZN(U2937) );
  AOI22_X1 U5754 ( .A1(n4660), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n4657), .ZN(n4650) );
  NAND2_X1 U5755 ( .A1(n4649), .A2(DATAI_8_), .ZN(n4655) );
  NAND2_X1 U5756 ( .A1(n4650), .A2(n4655), .ZN(U2947) );
  AOI22_X1 U5757 ( .A1(n4660), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n4657), .ZN(n4652) );
  NAND2_X1 U5758 ( .A1(n4652), .A2(n4651), .ZN(U2925) );
  AOI22_X1 U5759 ( .A1(n4660), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n4657), .ZN(n4654) );
  NAND2_X1 U5760 ( .A1(n4654), .A2(n4653), .ZN(U2926) );
  AOI22_X1 U5761 ( .A1(n4660), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n4657), .ZN(n4656) );
  NAND2_X1 U5762 ( .A1(n4656), .A2(n4655), .ZN(U2932) );
  AOI22_X1 U5763 ( .A1(n4660), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n4657), .ZN(n4659) );
  NAND2_X1 U5764 ( .A1(n4659), .A2(n4658), .ZN(U2931) );
  AOI22_X1 U5765 ( .A1(n4660), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n4657), .ZN(n4662) );
  NAND2_X1 U5766 ( .A1(n4662), .A2(n4661), .ZN(U2928) );
  INV_X1 U5767 ( .A(DATAI_7_), .ZN(n6617) );
  NOR2_X2 U5768 ( .A1(n4668), .A2(n4246), .ZN(n6422) );
  INV_X1 U5769 ( .A(DATAI_31_), .ZN(n4663) );
  OR2_X1 U5770 ( .A1(n6371), .A2(n4663), .ZN(n6267) );
  INV_X1 U5771 ( .A(DATAI_23_), .ZN(n6748) );
  OR2_X1 U5772 ( .A1(n6371), .A2(n6748), .ZN(n6429) );
  OAI22_X1 U5773 ( .A1(n6267), .A2(n5166), .B1(n5047), .B2(n6429), .ZN(n4664)
         );
  AOI21_X1 U5774 ( .B1(n6422), .B2(n4671), .A(n4664), .ZN(n4666) );
  NAND2_X1 U5775 ( .A1(n4672), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4665) );
  OAI211_X1 U5776 ( .C1(n4675), .C2(n6360), .A(n4666), .B(n4665), .ZN(U3067)
         );
  NOR2_X2 U5777 ( .A1(n4668), .A2(n3282), .ZN(n6408) );
  INV_X1 U5778 ( .A(DATAI_29_), .ZN(n4669) );
  OR2_X1 U5779 ( .A1(n6371), .A2(n4669), .ZN(n6257) );
  INV_X1 U5780 ( .A(DATAI_21_), .ZN(n6665) );
  OR2_X1 U5781 ( .A1(n6371), .A2(n6665), .ZN(n6412) );
  OAI22_X1 U5782 ( .A1(n6257), .A2(n5166), .B1(n5047), .B2(n6412), .ZN(n4670)
         );
  AOI21_X1 U5783 ( .B1(n6408), .B2(n4671), .A(n4670), .ZN(n4674) );
  NAND2_X1 U5784 ( .A1(n4672), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4673) );
  OAI211_X1 U5785 ( .C1(n4675), .C2(n6348), .A(n4674), .B(n4673), .ZN(U3065)
         );
  NAND2_X1 U5786 ( .A1(n3078), .A2(n4676), .ZN(n4684) );
  INV_X1 U5787 ( .A(n4684), .ZN(n4677) );
  NAND2_X1 U5788 ( .A1(n4408), .A2(n4342), .ZN(n4744) );
  INV_X1 U5789 ( .A(n6233), .ZN(n4678) );
  NAND3_X1 U5790 ( .A1(n6572), .A2(n6441), .A3(n6437), .ZN(n6229) );
  NOR2_X1 U5791 ( .A1(n6430), .A2(n6229), .ZN(n4831) );
  AOI21_X1 U5792 ( .B1(n4678), .B2(n6315), .A(n4831), .ZN(n4682) );
  OR2_X1 U5793 ( .A1(n4684), .A2(n6730), .ZN(n4679) );
  AOI22_X1 U5794 ( .A1(n4682), .A2(n4681), .B1(n6587), .B2(n6229), .ZN(n4680)
         );
  NAND2_X1 U5795 ( .A1(n6377), .A2(n4680), .ZN(n4830) );
  INV_X1 U5796 ( .A(n4681), .ZN(n4683) );
  OAI22_X1 U5797 ( .A1(n4683), .A2(n4682), .B1(n4573), .B2(n6229), .ZN(n4829)
         );
  AOI22_X1 U5798 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4830), .B1(n6389), 
        .B2(n4829), .ZN(n4686) );
  NOR2_X2 U5799 ( .A1(n4684), .A2(n4782), .ZN(n6263) );
  INV_X1 U5800 ( .A(n6248), .ZN(n6391) );
  AOI22_X1 U5801 ( .A1(n6263), .A2(n6391), .B1(n6390), .B2(n4831), .ZN(n4685)
         );
  OAI211_X1 U5802 ( .C1(n6394), .C2(n4933), .A(n4686), .B(n4685), .ZN(U3030)
         );
  AOI22_X1 U5803 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4830), .B1(n6368), 
        .B2(n4829), .ZN(n4688) );
  AOI22_X1 U5804 ( .A1(n6263), .A2(n6379), .B1(n6369), .B2(n4831), .ZN(n4687)
         );
  OAI211_X1 U5805 ( .C1(n6382), .C2(n4933), .A(n4688), .B(n4687), .ZN(U3028)
         );
  AOI22_X1 U5806 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4830), .B1(n6395), 
        .B2(n4829), .ZN(n4690) );
  AOI22_X1 U5807 ( .A1(n6263), .A2(n6397), .B1(n6396), .B2(n4831), .ZN(n4689)
         );
  OAI211_X1 U5808 ( .C1(n6400), .C2(n4933), .A(n4690), .B(n4689), .ZN(U3031)
         );
  XNOR2_X1 U5809 ( .A(n2995), .B(n4692), .ZN(n4743) );
  INV_X1 U5810 ( .A(n4693), .ZN(n6083) );
  NAND2_X1 U5811 ( .A1(n6083), .A2(n6138), .ZN(n4696) );
  AND2_X1 U5812 ( .A1(n6133), .A2(REIP_REG_6__SCAN_IN), .ZN(n4740) );
  AND2_X1 U5813 ( .A1(n6148), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4694)
         );
  AOI211_X1 U5814 ( .C1(n5613), .C2(n6032), .A(n4740), .B(n4694), .ZN(n4695)
         );
  OAI211_X1 U5815 ( .C1(n4743), .C2(n6145), .A(n4696), .B(n4695), .ZN(U2980)
         );
  NOR2_X1 U5816 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4697), .ZN(n4929)
         );
  INV_X1 U5817 ( .A(n4929), .ZN(n4701) );
  AND2_X1 U5818 ( .A1(n6568), .A2(n6730), .ZN(n6566) );
  AOI21_X1 U5819 ( .B1(n4933), .B2(n4930), .A(n6566), .ZN(n4698) );
  OAI21_X1 U5820 ( .B1(n4698), .B2(n4702), .A(n6562), .ZN(n4700) );
  AND2_X1 U5821 ( .A1(n4703), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6236) );
  OAI21_X1 U5822 ( .B1(n5205), .B2(n4573), .A(n5132), .ZN(n4784) );
  NOR2_X1 U5823 ( .A1(n6236), .A2(n4784), .ZN(n5210) );
  INV_X1 U5824 ( .A(n5210), .ZN(n4699) );
  INV_X1 U5825 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4709) );
  INV_X1 U5826 ( .A(n4702), .ZN(n4705) );
  NOR2_X1 U5827 ( .A1(n4703), .A2(n4573), .ZN(n5203) );
  NAND3_X1 U5828 ( .A1(n5203), .A2(n5205), .A3(n6572), .ZN(n4704) );
  OAI21_X1 U5829 ( .B1(n4705), .B2(n6587), .A(n4704), .ZN(n4928) );
  AOI22_X1 U5830 ( .A1(n6390), .A2(n4929), .B1(n6389), .B2(n4928), .ZN(n4706)
         );
  OAI21_X1 U5831 ( .B1(n6394), .B2(n4930), .A(n4706), .ZN(n4707) );
  AOI21_X1 U5832 ( .B1(n6391), .B2(n4888), .A(n4707), .ZN(n4708) );
  OAI21_X1 U5833 ( .B1(n4927), .B2(n4709), .A(n4708), .ZN(U3038) );
  INV_X1 U5834 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4713) );
  AOI22_X1 U5835 ( .A1(n6396), .A2(n4929), .B1(n6395), .B2(n4928), .ZN(n4710)
         );
  OAI21_X1 U5836 ( .B1(n6400), .B2(n4930), .A(n4710), .ZN(n4711) );
  AOI21_X1 U5837 ( .B1(n6397), .B2(n4888), .A(n4711), .ZN(n4712) );
  OAI21_X1 U5838 ( .B1(n4927), .B2(n4713), .A(n4712), .ZN(U3039) );
  NOR2_X1 U5839 ( .A1(n6306), .A2(n6587), .ZN(n4715) );
  AOI21_X1 U5840 ( .B1(n4904), .B2(n4715), .A(n6566), .ZN(n4718) );
  INV_X1 U5841 ( .A(n3017), .ZN(n4790) );
  NOR2_X1 U5842 ( .A1(n4790), .A2(n4744), .ZN(n4719) );
  NAND3_X1 U5843 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6441), .A3(n6437), .ZN(n4749) );
  NOR2_X1 U5844 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4749), .ZN(n4901)
         );
  INV_X1 U5845 ( .A(n4901), .ZN(n4716) );
  OAI21_X1 U5846 ( .B1(n3084), .B2(n4573), .A(n5132), .ZN(n4858) );
  AOI211_X1 U5847 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4716), .A(n6236), .B(
        n4858), .ZN(n4717) );
  NAND2_X1 U5848 ( .A1(n4897), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4722) );
  AOI22_X1 U5849 ( .A1(n4719), .A2(n6568), .B1(n5203), .B2(n3084), .ZN(n4898)
         );
  OAI22_X1 U5850 ( .A1(n4899), .A2(n6245), .B1(n4898), .B2(n6332), .ZN(n4720)
         );
  AOI21_X1 U5851 ( .B1(n6384), .B2(n4901), .A(n4720), .ZN(n4721) );
  OAI211_X1 U5852 ( .C1(n6388), .C2(n4904), .A(n4722), .B(n4721), .ZN(U3085)
         );
  NAND2_X1 U5853 ( .A1(n4897), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4725) );
  OAI22_X1 U5854 ( .A1(n4899), .A2(n6248), .B1(n4898), .B2(n6336), .ZN(n4723)
         );
  AOI21_X1 U5855 ( .B1(n6390), .B2(n4901), .A(n4723), .ZN(n4724) );
  OAI211_X1 U5856 ( .C1(n6394), .C2(n4904), .A(n4725), .B(n4724), .ZN(U3086)
         );
  NAND2_X1 U5857 ( .A1(n4897), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4728) );
  OAI22_X1 U5858 ( .A1(n4899), .A2(n6267), .B1(n4898), .B2(n6360), .ZN(n4726)
         );
  AOI21_X1 U5859 ( .B1(n6422), .B2(n4901), .A(n4726), .ZN(n4727) );
  OAI211_X1 U5860 ( .C1(n6429), .C2(n4904), .A(n4728), .B(n4727), .ZN(U3091)
         );
  NAND2_X1 U5861 ( .A1(n4897), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4731) );
  OAI22_X1 U5862 ( .A1(n4899), .A2(n6260), .B1(n4898), .B2(n6352), .ZN(n4729)
         );
  AOI21_X1 U5863 ( .B1(n6414), .B2(n4901), .A(n4729), .ZN(n4730) );
  OAI211_X1 U5864 ( .C1(n6418), .C2(n4904), .A(n4731), .B(n4730), .ZN(U3090)
         );
  NAND2_X1 U5865 ( .A1(n4897), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4734) );
  OAI22_X1 U5866 ( .A1(n4899), .A2(n6254), .B1(n4898), .B2(n6344), .ZN(n4732)
         );
  AOI21_X1 U5867 ( .B1(n6402), .B2(n4901), .A(n4732), .ZN(n4733) );
  OAI211_X1 U5868 ( .C1(n6406), .C2(n4904), .A(n4734), .B(n4733), .ZN(U3088)
         );
  NAND2_X1 U5869 ( .A1(n4897), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4737) );
  OAI22_X1 U5870 ( .A1(n4899), .A2(n6257), .B1(n4898), .B2(n6348), .ZN(n4735)
         );
  AOI21_X1 U5871 ( .B1(n6408), .B2(n4901), .A(n4735), .ZN(n4736) );
  OAI211_X1 U5872 ( .C1(n6412), .C2(n4904), .A(n4737), .B(n4736), .ZN(U3089)
         );
  NOR2_X1 U5873 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6185), .ZN(n4738)
         );
  AOI22_X1 U5874 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4739), .B1(n5069), 
        .B2(n4738), .ZN(n4742) );
  XNOR2_X1 U5875 ( .A(n4919), .B(n4916), .ZN(n6080) );
  AOI21_X1 U5876 ( .B1(n6170), .B2(n6080), .A(n4740), .ZN(n4741) );
  OAI211_X1 U5877 ( .C1(n6206), .C2(n4743), .A(n4742), .B(n4741), .ZN(U3012)
         );
  INV_X1 U5878 ( .A(n4744), .ZN(n4745) );
  NOR2_X1 U5879 ( .A1(n6430), .A2(n4749), .ZN(n4838) );
  AOI21_X1 U5880 ( .B1(n6363), .B2(n4745), .A(n4838), .ZN(n4751) );
  AOI21_X1 U5881 ( .B1(n4746), .B2(STATEBS16_REG_SCAN_IN), .A(n6587), .ZN(
        n4748) );
  AOI22_X1 U5882 ( .A1(n4751), .A2(n4748), .B1(n6587), .B2(n4749), .ZN(n4747)
         );
  NAND2_X1 U5883 ( .A1(n6377), .A2(n4747), .ZN(n4837) );
  INV_X1 U5884 ( .A(n4748), .ZN(n4750) );
  OAI22_X1 U5885 ( .A1(n4751), .A2(n4750), .B1(n4573), .B2(n4749), .ZN(n4836)
         );
  AOI22_X1 U5886 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4837), .B1(n6389), 
        .B2(n4836), .ZN(n4754) );
  INV_X1 U5887 ( .A(n6394), .ZN(n6333) );
  AOI22_X1 U5888 ( .A1(n5236), .A2(n6333), .B1(n4838), .B2(n6390), .ZN(n4753)
         );
  OAI211_X1 U5889 ( .C1(n4904), .C2(n6248), .A(n4754), .B(n4753), .ZN(U3094)
         );
  NAND2_X1 U5890 ( .A1(n6590), .A2(n5958), .ZN(n4755) );
  NAND2_X1 U5891 ( .A1(n4755), .A2(n5856), .ZN(n6067) );
  INV_X1 U5892 ( .A(n6067), .ZN(n5354) );
  OAI22_X1 U5893 ( .A1(n4990), .A2(n6078), .B1(n4756), .B2(n6061), .ZN(n4757)
         );
  AOI21_X1 U5894 ( .B1(n4758), .B2(REIP_REG_1__SCAN_IN), .A(n4757), .ZN(n4759)
         );
  OAI21_X1 U5895 ( .B1(n6039), .B2(n4761), .A(n4759), .ZN(n4760) );
  AOI21_X1 U5896 ( .B1(n6071), .B2(n4761), .A(n4760), .ZN(n4765) );
  AND2_X1 U5897 ( .A1(n6590), .A2(n4762), .ZN(n6064) );
  AOI22_X1 U5898 ( .A1(n6054), .A2(n6574), .B1(n6064), .B2(n4763), .ZN(n4764)
         );
  OAI211_X1 U5899 ( .C1(n5354), .C2(n4993), .A(n4765), .B(n4764), .ZN(U2826)
         );
  AOI22_X1 U5900 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4837), .B1(n6368), 
        .B2(n4836), .ZN(n4767) );
  INV_X1 U5901 ( .A(n6382), .ZN(n6320) );
  AOI22_X1 U5902 ( .A1(n5236), .A2(n6320), .B1(n6369), .B2(n4838), .ZN(n4766)
         );
  OAI211_X1 U5903 ( .C1(n4904), .C2(n6242), .A(n4767), .B(n4766), .ZN(U3092)
         );
  AOI22_X1 U5904 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4837), .B1(n6395), 
        .B2(n4836), .ZN(n4769) );
  INV_X1 U5905 ( .A(n6400), .ZN(n6337) );
  AOI22_X1 U5906 ( .A1(n5236), .A2(n6337), .B1(n4838), .B2(n6396), .ZN(n4768)
         );
  OAI211_X1 U5907 ( .C1(n4904), .C2(n6251), .A(n4769), .B(n4768), .ZN(U3095)
         );
  AOI22_X1 U5908 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4830), .B1(n6383), 
        .B2(n4829), .ZN(n4771) );
  INV_X1 U5909 ( .A(n6245), .ZN(n6385) );
  AOI22_X1 U5910 ( .A1(n6263), .A2(n6385), .B1(n6384), .B2(n4831), .ZN(n4770)
         );
  OAI211_X1 U5911 ( .C1(n6388), .C2(n4933), .A(n4771), .B(n4770), .ZN(U3029)
         );
  AOI22_X1 U5912 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4830), .B1(n6413), 
        .B2(n4829), .ZN(n4773) );
  INV_X1 U5913 ( .A(n6260), .ZN(n6415) );
  AOI22_X1 U5914 ( .A1(n6263), .A2(n6415), .B1(n6414), .B2(n4831), .ZN(n4772)
         );
  OAI211_X1 U5915 ( .C1(n6418), .C2(n4933), .A(n4773), .B(n4772), .ZN(U3034)
         );
  AOI22_X1 U5916 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4830), .B1(n6401), 
        .B2(n4829), .ZN(n4775) );
  INV_X1 U5917 ( .A(n6254), .ZN(n6403) );
  AOI22_X1 U5918 ( .A1(n6263), .A2(n6403), .B1(n6402), .B2(n4831), .ZN(n4774)
         );
  OAI211_X1 U5919 ( .C1(n6406), .C2(n4933), .A(n4775), .B(n4774), .ZN(U3032)
         );
  AOI22_X1 U5920 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4837), .B1(n6401), 
        .B2(n4836), .ZN(n4777) );
  INV_X1 U5921 ( .A(n6406), .ZN(n6341) );
  AOI22_X1 U5922 ( .A1(n5236), .A2(n6341), .B1(n4838), .B2(n6402), .ZN(n4776)
         );
  OAI211_X1 U5923 ( .C1(n4904), .C2(n6254), .A(n4777), .B(n4776), .ZN(U3096)
         );
  AOI22_X1 U5924 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4837), .B1(n6383), 
        .B2(n4836), .ZN(n4779) );
  INV_X1 U5925 ( .A(n6388), .ZN(n6329) );
  AOI22_X1 U5926 ( .A1(n5236), .A2(n6329), .B1(n4838), .B2(n6384), .ZN(n4778)
         );
  OAI211_X1 U5927 ( .C1(n4904), .C2(n6245), .A(n4779), .B(n4778), .ZN(U3093)
         );
  AOI22_X1 U5928 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4837), .B1(n6413), 
        .B2(n4836), .ZN(n4781) );
  INV_X1 U5929 ( .A(n6418), .ZN(n6349) );
  AOI22_X1 U5930 ( .A1(n5236), .A2(n6349), .B1(n4838), .B2(n6414), .ZN(n4780)
         );
  OAI211_X1 U5931 ( .C1(n4904), .C2(n6260), .A(n4781), .B(n4780), .ZN(U3098)
         );
  NOR2_X1 U5932 ( .A1(n4408), .A2(n4342), .ZN(n6362) );
  INV_X1 U5933 ( .A(n6362), .ZN(n5009) );
  NOR2_X2 U5934 ( .A1(n6370), .A2(n5198), .ZN(n6423) );
  OAI21_X1 U5935 ( .B1(n4980), .B2(n6423), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4783) );
  NAND3_X1 U5936 ( .A1(n5009), .A2(n6568), .A3(n4783), .ZN(n4788) );
  NOR2_X1 U5937 ( .A1(n5203), .A2(n4784), .ZN(n5013) );
  NOR2_X1 U5938 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4785), .ZN(n4823)
         );
  INV_X1 U5939 ( .A(n4823), .ZN(n4786) );
  AOI21_X1 U5940 ( .B1(n4786), .B2(STATE2_REG_3__SCAN_IN), .A(n6572), .ZN(
        n4787) );
  INV_X1 U5941 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4794) );
  INV_X1 U5942 ( .A(n6412), .ZN(n6345) );
  NAND2_X1 U5943 ( .A1(n6362), .A2(n6568), .ZN(n5016) );
  NAND3_X1 U5944 ( .A1(n6236), .A2(n5205), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4789) );
  OAI21_X1 U5945 ( .B1(n5016), .B2(n4790), .A(n4789), .ZN(n4819) );
  AOI22_X1 U5946 ( .A1(n6423), .A2(n6345), .B1(n6407), .B2(n4819), .ZN(n4791)
         );
  OAI21_X1 U5947 ( .B1(n4821), .B2(n6257), .A(n4791), .ZN(n4792) );
  AOI21_X1 U5948 ( .B1(n6408), .B2(n4823), .A(n4792), .ZN(n4793) );
  OAI21_X1 U5949 ( .B1(n4826), .B2(n4794), .A(n4793), .ZN(U3137) );
  INV_X1 U5950 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4798) );
  AOI22_X1 U5951 ( .A1(n6423), .A2(n6333), .B1(n6389), .B2(n4819), .ZN(n4795)
         );
  OAI21_X1 U5952 ( .B1(n4821), .B2(n6248), .A(n4795), .ZN(n4796) );
  AOI21_X1 U5953 ( .B1(n6390), .B2(n4823), .A(n4796), .ZN(n4797) );
  OAI21_X1 U5954 ( .B1(n4826), .B2(n4798), .A(n4797), .ZN(U3134) );
  INV_X1 U5955 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4802) );
  AOI22_X1 U5956 ( .A1(n6423), .A2(n6320), .B1(n6368), .B2(n4819), .ZN(n4799)
         );
  OAI21_X1 U5957 ( .B1(n6242), .B2(n4821), .A(n4799), .ZN(n4800) );
  AOI21_X1 U5958 ( .B1(n6369), .B2(n4823), .A(n4800), .ZN(n4801) );
  OAI21_X1 U5959 ( .B1(n4826), .B2(n4802), .A(n4801), .ZN(U3132) );
  INV_X1 U5960 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4806) );
  INV_X1 U5961 ( .A(n6429), .ZN(n6354) );
  AOI22_X1 U5962 ( .A1(n6423), .A2(n6354), .B1(n6420), .B2(n4819), .ZN(n4803)
         );
  OAI21_X1 U5963 ( .B1(n4821), .B2(n6267), .A(n4803), .ZN(n4804) );
  AOI21_X1 U5964 ( .B1(n6422), .B2(n4823), .A(n4804), .ZN(n4805) );
  OAI21_X1 U5965 ( .B1(n4826), .B2(n4806), .A(n4805), .ZN(U3139) );
  INV_X1 U5966 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4810) );
  AOI22_X1 U5967 ( .A1(n6423), .A2(n6337), .B1(n6395), .B2(n4819), .ZN(n4807)
         );
  OAI21_X1 U5968 ( .B1(n4821), .B2(n6251), .A(n4807), .ZN(n4808) );
  AOI21_X1 U5969 ( .B1(n6396), .B2(n4823), .A(n4808), .ZN(n4809) );
  OAI21_X1 U5970 ( .B1(n4826), .B2(n4810), .A(n4809), .ZN(U3135) );
  INV_X1 U5971 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4814) );
  AOI22_X1 U5972 ( .A1(n6423), .A2(n6341), .B1(n6401), .B2(n4819), .ZN(n4811)
         );
  OAI21_X1 U5973 ( .B1(n4821), .B2(n6254), .A(n4811), .ZN(n4812) );
  AOI21_X1 U5974 ( .B1(n6402), .B2(n4823), .A(n4812), .ZN(n4813) );
  OAI21_X1 U5975 ( .B1(n4826), .B2(n4814), .A(n4813), .ZN(U3136) );
  INV_X1 U5976 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4818) );
  AOI22_X1 U5977 ( .A1(n6423), .A2(n6349), .B1(n6413), .B2(n4819), .ZN(n4815)
         );
  OAI21_X1 U5978 ( .B1(n4821), .B2(n6260), .A(n4815), .ZN(n4816) );
  AOI21_X1 U5979 ( .B1(n6414), .B2(n4823), .A(n4816), .ZN(n4817) );
  OAI21_X1 U5980 ( .B1(n4826), .B2(n4818), .A(n4817), .ZN(U3138) );
  INV_X1 U5981 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4825) );
  AOI22_X1 U5982 ( .A1(n6423), .A2(n6329), .B1(n6383), .B2(n4819), .ZN(n4820)
         );
  OAI21_X1 U5983 ( .B1(n4821), .B2(n6245), .A(n4820), .ZN(n4822) );
  AOI21_X1 U5984 ( .B1(n6384), .B2(n4823), .A(n4822), .ZN(n4824) );
  OAI21_X1 U5985 ( .B1(n4826), .B2(n4825), .A(n4824), .ZN(U3133) );
  AOI22_X1 U5986 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4830), .B1(n6407), 
        .B2(n4829), .ZN(n4828) );
  INV_X1 U5987 ( .A(n6257), .ZN(n6409) );
  AOI22_X1 U5988 ( .A1(n6263), .A2(n6409), .B1(n6408), .B2(n4831), .ZN(n4827)
         );
  OAI211_X1 U5989 ( .C1(n6412), .C2(n4933), .A(n4828), .B(n4827), .ZN(U3033)
         );
  AOI22_X1 U5990 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4830), .B1(n6420), 
        .B2(n4829), .ZN(n4833) );
  INV_X1 U5991 ( .A(n6267), .ZN(n6424) );
  AOI22_X1 U5992 ( .A1(n6263), .A2(n6424), .B1(n6422), .B2(n4831), .ZN(n4832)
         );
  OAI211_X1 U5993 ( .C1(n6429), .C2(n4933), .A(n4833), .B(n4832), .ZN(U3035)
         );
  AOI22_X1 U5994 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4837), .B1(n6420), 
        .B2(n4836), .ZN(n4835) );
  AOI22_X1 U5995 ( .A1(n5236), .A2(n6354), .B1(n4838), .B2(n6422), .ZN(n4834)
         );
  OAI211_X1 U5996 ( .C1(n4904), .C2(n6267), .A(n4835), .B(n4834), .ZN(U3099)
         );
  AOI22_X1 U5997 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4837), .B1(n6407), 
        .B2(n4836), .ZN(n4840) );
  AOI22_X1 U5998 ( .A1(n5236), .A2(n6345), .B1(n4838), .B2(n6408), .ZN(n4839)
         );
  OAI211_X1 U5999 ( .C1(n4904), .C2(n6257), .A(n4840), .B(n4839), .ZN(U3097)
         );
  INV_X1 U6000 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4844) );
  AOI22_X1 U6001 ( .A1(n6384), .A2(n4929), .B1(n6383), .B2(n4928), .ZN(n4841)
         );
  OAI21_X1 U6002 ( .B1(n6388), .B2(n4930), .A(n4841), .ZN(n4842) );
  AOI21_X1 U6003 ( .B1(n6385), .B2(n4888), .A(n4842), .ZN(n4843) );
  OAI21_X1 U6004 ( .B1(n4927), .B2(n4844), .A(n4843), .ZN(U3037) );
  INV_X1 U6005 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4848) );
  AOI22_X1 U6006 ( .A1(n6414), .A2(n4929), .B1(n6413), .B2(n4928), .ZN(n4845)
         );
  OAI21_X1 U6007 ( .B1(n6418), .B2(n4930), .A(n4845), .ZN(n4846) );
  AOI21_X1 U6008 ( .B1(n6415), .B2(n4888), .A(n4846), .ZN(n4847) );
  OAI21_X1 U6009 ( .B1(n4927), .B2(n4848), .A(n4847), .ZN(U3042) );
  INV_X1 U6010 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4852) );
  AOI22_X1 U6011 ( .A1(n6402), .A2(n4929), .B1(n6401), .B2(n4928), .ZN(n4849)
         );
  OAI21_X1 U6012 ( .B1(n6406), .B2(n4930), .A(n4849), .ZN(n4850) );
  AOI21_X1 U6013 ( .B1(n6403), .B2(n4888), .A(n4850), .ZN(n4851) );
  OAI21_X1 U6014 ( .B1(n4927), .B2(n4852), .A(n4851), .ZN(U3040) );
  NAND3_X1 U6015 ( .A1(n4978), .A2(n6568), .A3(n6319), .ZN(n4855) );
  INV_X1 U6016 ( .A(n6566), .ZN(n5199) );
  AOI22_X1 U6017 ( .A1(n4855), .A2(n5199), .B1(n5136), .B2(n5008), .ZN(n4857)
         );
  NOR2_X1 U6018 ( .A1(n6572), .A2(n4940), .ZN(n4946) );
  INV_X1 U6019 ( .A(n4946), .ZN(n4938) );
  NOR2_X1 U6020 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4938), .ZN(n4908)
         );
  NOR2_X1 U6021 ( .A1(n4908), .A2(n6562), .ZN(n4856) );
  NAND2_X1 U6022 ( .A1(n4905), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4864)
         );
  INV_X1 U6023 ( .A(n5136), .ZN(n4859) );
  NOR2_X1 U6024 ( .A1(n4859), .A2(n6587), .ZN(n5127) );
  NAND2_X1 U6025 ( .A1(n5127), .A2(n3017), .ZN(n4861) );
  NAND2_X1 U6026 ( .A1(n3084), .A2(n6236), .ZN(n4860) );
  OAI22_X1 U6027 ( .A1(n4978), .A2(n6418), .B1(n4906), .B2(n6352), .ZN(n4862)
         );
  AOI21_X1 U6028 ( .B1(n6414), .B2(n4908), .A(n4862), .ZN(n4863) );
  OAI211_X1 U6029 ( .C1(n6319), .C2(n6260), .A(n4864), .B(n4863), .ZN(U3122)
         );
  NAND2_X1 U6030 ( .A1(n4905), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4867)
         );
  OAI22_X1 U6031 ( .A1(n4978), .A2(n6394), .B1(n4906), .B2(n6336), .ZN(n4865)
         );
  AOI21_X1 U6032 ( .B1(n6390), .B2(n4908), .A(n4865), .ZN(n4866) );
  OAI211_X1 U6033 ( .C1(n6319), .C2(n6248), .A(n4867), .B(n4866), .ZN(U3118)
         );
  NAND2_X1 U6034 ( .A1(n4905), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4870)
         );
  OAI22_X1 U6035 ( .A1(n4978), .A2(n6406), .B1(n4906), .B2(n6344), .ZN(n4868)
         );
  AOI21_X1 U6036 ( .B1(n6402), .B2(n4908), .A(n4868), .ZN(n4869) );
  OAI211_X1 U6037 ( .C1(n6319), .C2(n6254), .A(n4870), .B(n4869), .ZN(U3120)
         );
  NAND2_X1 U6038 ( .A1(n4905), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4873)
         );
  OAI22_X1 U6039 ( .A1(n4978), .A2(n6388), .B1(n4906), .B2(n6332), .ZN(n4871)
         );
  AOI21_X1 U6040 ( .B1(n6384), .B2(n4908), .A(n4871), .ZN(n4872) );
  OAI211_X1 U6041 ( .C1(n6319), .C2(n6245), .A(n4873), .B(n4872), .ZN(U3117)
         );
  NAND2_X1 U6042 ( .A1(n4905), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4876)
         );
  OAI22_X1 U6043 ( .A1(n4978), .A2(n6412), .B1(n4906), .B2(n6348), .ZN(n4874)
         );
  AOI21_X1 U6044 ( .B1(n6408), .B2(n4908), .A(n4874), .ZN(n4875) );
  OAI211_X1 U6045 ( .C1(n6319), .C2(n6257), .A(n4876), .B(n4875), .ZN(U3121)
         );
  NAND2_X1 U6046 ( .A1(n4905), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4879)
         );
  OAI22_X1 U6047 ( .A1(n4978), .A2(n6429), .B1(n4906), .B2(n6360), .ZN(n4877)
         );
  AOI21_X1 U6048 ( .B1(n6422), .B2(n4908), .A(n4877), .ZN(n4878) );
  OAI211_X1 U6049 ( .C1(n6319), .C2(n6267), .A(n4879), .B(n4878), .ZN(U3123)
         );
  AOI22_X1 U6050 ( .A1(n6081), .A2(n6036), .B1(n5485), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4880) );
  OAI21_X1 U6051 ( .B1(n4881), .B2(n5506), .A(n4880), .ZN(U2854) );
  INV_X1 U6052 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4885) );
  AOI22_X1 U6053 ( .A1(n6422), .A2(n4929), .B1(n6420), .B2(n4928), .ZN(n4882)
         );
  OAI21_X1 U6054 ( .B1(n6429), .B2(n4930), .A(n4882), .ZN(n4883) );
  AOI21_X1 U6055 ( .B1(n6424), .B2(n4888), .A(n4883), .ZN(n4884) );
  OAI21_X1 U6056 ( .B1(n4927), .B2(n4885), .A(n4884), .ZN(U3043) );
  INV_X1 U6057 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4890) );
  AOI22_X1 U6058 ( .A1(n6408), .A2(n4929), .B1(n6407), .B2(n4928), .ZN(n4886)
         );
  OAI21_X1 U6059 ( .B1(n6412), .B2(n4930), .A(n4886), .ZN(n4887) );
  AOI21_X1 U6060 ( .B1(n6409), .B2(n4888), .A(n4887), .ZN(n4889) );
  OAI21_X1 U6061 ( .B1(n4927), .B2(n4890), .A(n4889), .ZN(U3041) );
  NAND2_X1 U6062 ( .A1(n4905), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4893)
         );
  OAI22_X1 U6063 ( .A1(n4978), .A2(n6382), .B1(n4906), .B2(n6328), .ZN(n4891)
         );
  AOI21_X1 U6064 ( .B1(n6369), .B2(n4908), .A(n4891), .ZN(n4892) );
  OAI211_X1 U6065 ( .C1(n6319), .C2(n6242), .A(n4893), .B(n4892), .ZN(U3116)
         );
  NAND2_X1 U6066 ( .A1(n4897), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4896) );
  OAI22_X1 U6067 ( .A1(n4899), .A2(n6242), .B1(n4898), .B2(n6328), .ZN(n4894)
         );
  AOI21_X1 U6068 ( .B1(n6369), .B2(n4901), .A(n4894), .ZN(n4895) );
  OAI211_X1 U6069 ( .C1(n6382), .C2(n4904), .A(n4896), .B(n4895), .ZN(U3084)
         );
  NAND2_X1 U6070 ( .A1(n4897), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4903) );
  OAI22_X1 U6071 ( .A1(n4899), .A2(n6251), .B1(n4898), .B2(n6340), .ZN(n4900)
         );
  AOI21_X1 U6072 ( .B1(n6396), .B2(n4901), .A(n4900), .ZN(n4902) );
  OAI211_X1 U6073 ( .C1(n6400), .C2(n4904), .A(n4903), .B(n4902), .ZN(U3087)
         );
  NAND2_X1 U6074 ( .A1(n4905), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4910)
         );
  OAI22_X1 U6075 ( .A1(n4978), .A2(n6400), .B1(n4906), .B2(n6340), .ZN(n4907)
         );
  AOI21_X1 U6076 ( .B1(n6396), .B2(n4908), .A(n4907), .ZN(n4909) );
  OAI211_X1 U6077 ( .C1(n6319), .C2(n6251), .A(n4910), .B(n4909), .ZN(U3119)
         );
  INV_X1 U6078 ( .A(n4911), .ZN(n4915) );
  AOI21_X1 U6079 ( .B1(n4915), .B2(n4914), .A(n3571), .ZN(n6025) );
  INV_X1 U6080 ( .A(n6025), .ZN(n4937) );
  INV_X1 U6081 ( .A(n4916), .ZN(n4918) );
  OAI21_X1 U6082 ( .B1(n4919), .B2(n4918), .A(n4917), .ZN(n4920) );
  AND2_X1 U6083 ( .A1(n4920), .A2(n5074), .ZN(n6169) );
  AOI22_X1 U6084 ( .A1(n6081), .A2(n6169), .B1(EBX_REG_7__SCAN_IN), .B2(n5485), 
        .ZN(n4921) );
  OAI21_X1 U6085 ( .B1(n4937), .B2(n5506), .A(n4921), .ZN(U2852) );
  NOR2_X1 U6086 ( .A1(n5359), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4922)
         );
  OR2_X1 U6087 ( .A1(n4923), .A2(n4922), .ZN(n6217) );
  OAI222_X1 U6088 ( .A1(n6151), .A2(n5506), .B1(n4924), .B2(n5504), .C1(n6217), 
        .C2(n5503), .ZN(U2859) );
  INV_X1 U6089 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4925) );
  OAI222_X1 U6090 ( .A1(n4926), .A2(n5506), .B1(n4925), .B2(n6086), .C1(n5503), 
        .C2(n6060), .ZN(U2855) );
  INV_X1 U6091 ( .A(n4927), .ZN(n4935) );
  AOI22_X1 U6092 ( .A1(n6369), .A2(n4929), .B1(n6368), .B2(n4928), .ZN(n4932)
         );
  OR2_X1 U6093 ( .A1(n4930), .A2(n6382), .ZN(n4931) );
  OAI211_X1 U6094 ( .C1(n4933), .C2(n6242), .A(n4932), .B(n4931), .ZN(n4934)
         );
  AOI21_X1 U6095 ( .B1(n4935), .B2(INSTQUEUE_REG_2__0__SCAN_IN), .A(n4934), 
        .ZN(n4936) );
  INV_X1 U6096 ( .A(n4936), .ZN(U3036) );
  INV_X1 U6097 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6114) );
  OAI222_X1 U6098 ( .A1(n4937), .A2(n5524), .B1(n5299), .B2(n6617), .C1(n5507), 
        .C2(n6114), .ZN(U2884) );
  INV_X1 U6099 ( .A(n6408), .ZN(n4950) );
  NOR2_X1 U6100 ( .A1(n6430), .A2(n4938), .ZN(n4939) );
  INV_X1 U6101 ( .A(n4939), .ZN(n4982) );
  AOI21_X1 U6102 ( .B1(n6363), .B2(n5136), .A(n4939), .ZN(n4943) );
  NAND2_X1 U6103 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4941) );
  OAI22_X1 U6104 ( .A1(n4943), .A2(n6587), .B1(n4941), .B2(n4940), .ZN(n4976)
         );
  NAND2_X1 U6105 ( .A1(n4943), .A2(n4942), .ZN(n4944) );
  OR2_X1 U6106 ( .A1(n6587), .A2(n4944), .ZN(n4945) );
  OAI211_X1 U6107 ( .C1(n6568), .C2(n4946), .A(n4945), .B(n6377), .ZN(n4975)
         );
  AOI22_X1 U6108 ( .A1(n4976), .A2(n6407), .B1(INSTQUEUE_REG_13__5__SCAN_IN), 
        .B2(n4975), .ZN(n4947) );
  OAI21_X1 U6109 ( .B1(n4978), .B2(n6257), .A(n4947), .ZN(n4948) );
  AOI21_X1 U6110 ( .B1(n6345), .B2(n4980), .A(n4948), .ZN(n4949) );
  OAI21_X1 U6111 ( .B1(n4950), .B2(n4982), .A(n4949), .ZN(U3129) );
  INV_X1 U6112 ( .A(n6384), .ZN(n4954) );
  AOI22_X1 U6113 ( .A1(n4976), .A2(n6383), .B1(INSTQUEUE_REG_13__1__SCAN_IN), 
        .B2(n4975), .ZN(n4951) );
  OAI21_X1 U6114 ( .B1(n4978), .B2(n6245), .A(n4951), .ZN(n4952) );
  AOI21_X1 U6115 ( .B1(n6329), .B2(n4980), .A(n4952), .ZN(n4953) );
  OAI21_X1 U6116 ( .B1(n4954), .B2(n4982), .A(n4953), .ZN(U3125) );
  INV_X1 U6117 ( .A(n6422), .ZN(n4958) );
  AOI22_X1 U6118 ( .A1(n4976), .A2(n6420), .B1(INSTQUEUE_REG_13__7__SCAN_IN), 
        .B2(n4975), .ZN(n4955) );
  OAI21_X1 U6119 ( .B1(n4978), .B2(n6267), .A(n4955), .ZN(n4956) );
  AOI21_X1 U6120 ( .B1(n6354), .B2(n4980), .A(n4956), .ZN(n4957) );
  OAI21_X1 U6121 ( .B1(n4958), .B2(n4982), .A(n4957), .ZN(U3131) );
  INV_X1 U6122 ( .A(n6414), .ZN(n4962) );
  AOI22_X1 U6123 ( .A1(n4976), .A2(n6413), .B1(INSTQUEUE_REG_13__6__SCAN_IN), 
        .B2(n4975), .ZN(n4959) );
  OAI21_X1 U6124 ( .B1(n4978), .B2(n6260), .A(n4959), .ZN(n4960) );
  AOI21_X1 U6125 ( .B1(n6349), .B2(n4980), .A(n4960), .ZN(n4961) );
  OAI21_X1 U6126 ( .B1(n4962), .B2(n4982), .A(n4961), .ZN(U3130) );
  INV_X1 U6127 ( .A(n6402), .ZN(n4966) );
  AOI22_X1 U6128 ( .A1(n4976), .A2(n6401), .B1(INSTQUEUE_REG_13__4__SCAN_IN), 
        .B2(n4975), .ZN(n4963) );
  OAI21_X1 U6129 ( .B1(n4978), .B2(n6254), .A(n4963), .ZN(n4964) );
  AOI21_X1 U6130 ( .B1(n6341), .B2(n4980), .A(n4964), .ZN(n4965) );
  OAI21_X1 U6131 ( .B1(n4966), .B2(n4982), .A(n4965), .ZN(U3128) );
  INV_X1 U6132 ( .A(n6396), .ZN(n4970) );
  AOI22_X1 U6133 ( .A1(n4976), .A2(n6395), .B1(INSTQUEUE_REG_13__3__SCAN_IN), 
        .B2(n4975), .ZN(n4967) );
  OAI21_X1 U6134 ( .B1(n4978), .B2(n6251), .A(n4967), .ZN(n4968) );
  AOI21_X1 U6135 ( .B1(n6337), .B2(n4980), .A(n4968), .ZN(n4969) );
  OAI21_X1 U6136 ( .B1(n4970), .B2(n4982), .A(n4969), .ZN(U3127) );
  INV_X1 U6137 ( .A(n6390), .ZN(n4974) );
  AOI22_X1 U6138 ( .A1(n4976), .A2(n6389), .B1(INSTQUEUE_REG_13__2__SCAN_IN), 
        .B2(n4975), .ZN(n4971) );
  OAI21_X1 U6139 ( .B1(n4978), .B2(n6248), .A(n4971), .ZN(n4972) );
  AOI21_X1 U6140 ( .B1(n6333), .B2(n4980), .A(n4972), .ZN(n4973) );
  OAI21_X1 U6141 ( .B1(n4974), .B2(n4982), .A(n4973), .ZN(U3126) );
  INV_X1 U6142 ( .A(n6369), .ZN(n4983) );
  AOI22_X1 U6143 ( .A1(n4976), .A2(n6368), .B1(INSTQUEUE_REG_13__0__SCAN_IN), 
        .B2(n4975), .ZN(n4977) );
  OAI21_X1 U6144 ( .B1(n4978), .B2(n6242), .A(n4977), .ZN(n4979) );
  AOI21_X1 U6145 ( .B1(n6320), .B2(n4980), .A(n4979), .ZN(n4981) );
  OAI21_X1 U6146 ( .B1(n4983), .B2(n4982), .A(n4981), .ZN(U3124) );
  NAND2_X1 U6147 ( .A1(n4985), .A2(n4984), .ZN(n4986) );
  AND2_X1 U6148 ( .A1(n4995), .A2(n4986), .ZN(n6065) );
  INV_X1 U6149 ( .A(n6065), .ZN(n6191) );
  OAI22_X1 U6150 ( .A1(n5503), .A2(n6191), .B1(n6079), .B2(n6086), .ZN(n4987)
         );
  AOI21_X1 U6151 ( .B1(n6139), .B2(n6082), .A(n4987), .ZN(n4988) );
  INV_X1 U6152 ( .A(n4988), .ZN(U2857) );
  XNOR2_X1 U6153 ( .A(n4756), .B(n4989), .ZN(n6208) );
  OAI22_X1 U6154 ( .A1(n5503), .A2(n6208), .B1(n4990), .B2(n6086), .ZN(n4991)
         );
  INV_X1 U6155 ( .A(n4991), .ZN(n4992) );
  OAI21_X1 U6156 ( .B1(n5506), .B2(n4993), .A(n4992), .ZN(U2858) );
  INV_X1 U6157 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4998) );
  NAND2_X1 U6158 ( .A1(n4995), .A2(n4994), .ZN(n4996) );
  NAND2_X1 U6159 ( .A1(n4997), .A2(n4996), .ZN(n6180) );
  OAI222_X1 U6160 ( .A1(n5353), .A2(n5506), .B1(n4998), .B2(n6086), .C1(n6180), 
        .C2(n5503), .ZN(U2856) );
  AOI22_X1 U6161 ( .A1(n6275), .A2(n6409), .B1(n6408), .B2(n6274), .ZN(n4999)
         );
  OAI21_X1 U6162 ( .B1(n6412), .B2(n6280), .A(n4999), .ZN(n5000) );
  AOI21_X1 U6163 ( .B1(n6277), .B2(INSTQUEUE_REG_3__5__SCAN_IN), .A(n5000), 
        .ZN(n5001) );
  OAI21_X1 U6164 ( .B1(n5005), .B2(n6348), .A(n5001), .ZN(U3049) );
  AOI22_X1 U6165 ( .A1(n6275), .A2(n6424), .B1(n6422), .B2(n6274), .ZN(n5002)
         );
  OAI21_X1 U6166 ( .B1(n6429), .B2(n6280), .A(n5002), .ZN(n5003) );
  AOI21_X1 U6167 ( .B1(n6277), .B2(INSTQUEUE_REG_3__7__SCAN_IN), .A(n5003), 
        .ZN(n5004) );
  OAI21_X1 U6168 ( .B1(n5005), .B2(n6360), .A(n5004), .ZN(U3051) );
  INV_X1 U6169 ( .A(n6284), .ZN(n6286) );
  NOR2_X1 U6170 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6286), .ZN(n5049)
         );
  INV_X1 U6171 ( .A(n5049), .ZN(n5012) );
  INV_X1 U6172 ( .A(n6304), .ZN(n5007) );
  AOI21_X1 U6173 ( .B1(n5007), .B2(n5047), .A(n6730), .ZN(n5010) );
  NOR2_X1 U6174 ( .A1(n5009), .A2(n5008), .ZN(n6283) );
  NOR2_X1 U6175 ( .A1(n5010), .A2(n6283), .ZN(n5011) );
  AOI22_X1 U6176 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5012), .B1(n6568), .B2(
        n5011), .ZN(n5014) );
  INV_X1 U6177 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5020) );
  NAND3_X1 U6178 ( .A1(n6236), .A2(n5205), .A3(n6572), .ZN(n5015) );
  OAI21_X1 U6179 ( .B1(n5016), .B2(n3017), .A(n5015), .ZN(n5045) );
  AOI22_X1 U6180 ( .A1(n6304), .A2(n6320), .B1(n6368), .B2(n5045), .ZN(n5017)
         );
  OAI21_X1 U6181 ( .B1(n6242), .B2(n5047), .A(n5017), .ZN(n5018) );
  AOI21_X1 U6182 ( .B1(n6369), .B2(n5049), .A(n5018), .ZN(n5019) );
  OAI21_X1 U6183 ( .B1(n3087), .B2(n5020), .A(n5019), .ZN(U3068) );
  INV_X1 U6184 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5024) );
  AOI22_X1 U6185 ( .A1(n6304), .A2(n6354), .B1(n6420), .B2(n5045), .ZN(n5021)
         );
  OAI21_X1 U6186 ( .B1(n6267), .B2(n5047), .A(n5021), .ZN(n5022) );
  AOI21_X1 U6187 ( .B1(n6422), .B2(n5049), .A(n5022), .ZN(n5023) );
  OAI21_X1 U6188 ( .B1(n3087), .B2(n5024), .A(n5023), .ZN(U3075) );
  INV_X1 U6189 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5028) );
  AOI22_X1 U6190 ( .A1(n6304), .A2(n6329), .B1(n6383), .B2(n5045), .ZN(n5025)
         );
  OAI21_X1 U6191 ( .B1(n6245), .B2(n5047), .A(n5025), .ZN(n5026) );
  AOI21_X1 U6192 ( .B1(n6384), .B2(n5049), .A(n5026), .ZN(n5027) );
  OAI21_X1 U6193 ( .B1(n3087), .B2(n5028), .A(n5027), .ZN(U3069) );
  INV_X1 U6194 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5032) );
  AOI22_X1 U6195 ( .A1(n6304), .A2(n6333), .B1(n6389), .B2(n5045), .ZN(n5029)
         );
  OAI21_X1 U6196 ( .B1(n6248), .B2(n5047), .A(n5029), .ZN(n5030) );
  AOI21_X1 U6197 ( .B1(n6390), .B2(n5049), .A(n5030), .ZN(n5031) );
  OAI21_X1 U6198 ( .B1(n3087), .B2(n5032), .A(n5031), .ZN(U3070) );
  INV_X1 U6199 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5036) );
  AOI22_X1 U6200 ( .A1(n6304), .A2(n6337), .B1(n6395), .B2(n5045), .ZN(n5033)
         );
  OAI21_X1 U6201 ( .B1(n6251), .B2(n5047), .A(n5033), .ZN(n5034) );
  AOI21_X1 U6202 ( .B1(n6396), .B2(n5049), .A(n5034), .ZN(n5035) );
  OAI21_X1 U6203 ( .B1(n3087), .B2(n5036), .A(n5035), .ZN(U3071) );
  INV_X1 U6204 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5040) );
  AOI22_X1 U6205 ( .A1(n6304), .A2(n6341), .B1(n6401), .B2(n5045), .ZN(n5037)
         );
  OAI21_X1 U6206 ( .B1(n6254), .B2(n5047), .A(n5037), .ZN(n5038) );
  AOI21_X1 U6207 ( .B1(n6402), .B2(n5049), .A(n5038), .ZN(n5039) );
  OAI21_X1 U6208 ( .B1(n3087), .B2(n5040), .A(n5039), .ZN(U3072) );
  INV_X1 U6209 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5044) );
  AOI22_X1 U6210 ( .A1(n6304), .A2(n6345), .B1(n6407), .B2(n5045), .ZN(n5041)
         );
  OAI21_X1 U6211 ( .B1(n6257), .B2(n5047), .A(n5041), .ZN(n5042) );
  AOI21_X1 U6212 ( .B1(n6408), .B2(n5049), .A(n5042), .ZN(n5043) );
  OAI21_X1 U6213 ( .B1(n3087), .B2(n5044), .A(n5043), .ZN(U3073) );
  INV_X1 U6214 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5051) );
  AOI22_X1 U6215 ( .A1(n6304), .A2(n6349), .B1(n6413), .B2(n5045), .ZN(n5046)
         );
  OAI21_X1 U6216 ( .B1(n6260), .B2(n5047), .A(n5046), .ZN(n5048) );
  AOI21_X1 U6217 ( .B1(n6414), .B2(n5049), .A(n5048), .ZN(n5050) );
  OAI21_X1 U6218 ( .B1(n3087), .B2(n5051), .A(n5050), .ZN(U3074) );
  AND2_X1 U6219 ( .A1(n5052), .A2(n5053), .ZN(n5055) );
  OR2_X1 U6220 ( .A1(n5055), .A2(n5054), .ZN(n5119) );
  OR2_X1 U6221 ( .A1(n5075), .A2(n5056), .ZN(n5057) );
  AND2_X1 U6222 ( .A1(n5178), .A2(n5057), .ZN(n6162) );
  INV_X1 U6223 ( .A(n6162), .ZN(n5059) );
  OAI22_X1 U6224 ( .A1(n5503), .A2(n5059), .B1(n5058), .B2(n6086), .ZN(n5060)
         );
  INV_X1 U6225 ( .A(n5060), .ZN(n5061) );
  OAI21_X1 U6226 ( .B1(n5119), .B2(n5506), .A(n5061), .ZN(U2850) );
  INV_X1 U6227 ( .A(n6064), .ZN(n5062) );
  OAI22_X1 U6228 ( .A1(n3428), .A2(n5062), .B1(n5354), .B2(n6151), .ZN(n5063)
         );
  AOI21_X1 U6229 ( .B1(REIP_REG_0__SCAN_IN), .B2(n5864), .A(n5063), .ZN(n5066)
         );
  NAND2_X1 U6230 ( .A1(n6039), .A2(n6047), .ZN(n5064) );
  AOI22_X1 U6231 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n5064), .B1(n6050), 
        .B2(EBX_REG_0__SCAN_IN), .ZN(n5065) );
  OAI211_X1 U6232 ( .C1(n6061), .C2(n6217), .A(n5066), .B(n5065), .ZN(U2827)
         );
  XNOR2_X1 U6233 ( .A(n5067), .B(n5068), .ZN(n5101) );
  NAND2_X1 U6234 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5069), .ZN(n5071)
         );
  NOR2_X1 U6235 ( .A1(n5070), .A2(n5071), .ZN(n5283) );
  NOR2_X1 U6236 ( .A1(n6195), .A2(n5071), .ZN(n5287) );
  OAI22_X1 U6237 ( .A1(n5280), .A2(n5283), .B1(n5287), .B2(n5929), .ZN(n5072)
         );
  NOR2_X1 U6238 ( .A1(n5284), .A2(n5072), .ZN(n6178) );
  INV_X1 U6239 ( .A(n6178), .ZN(n5081) );
  AND2_X1 U6240 ( .A1(n5074), .A2(n5073), .ZN(n5076) );
  OR2_X1 U6241 ( .A1(n5076), .A2(n5075), .ZN(n6010) );
  NAND2_X1 U6242 ( .A1(n6133), .A2(REIP_REG_8__SCAN_IN), .ZN(n5097) );
  OAI21_X1 U6243 ( .B1(n6218), .B2(n6010), .A(n5097), .ZN(n5080) );
  NAND2_X1 U6244 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5282) );
  INV_X1 U6245 ( .A(n5282), .ZN(n5247) );
  NAND2_X1 U6246 ( .A1(n5287), .A2(n5077), .ZN(n6173) );
  AOI211_X1 U6247 ( .C1(n6177), .C2(n5078), .A(n5247), .B(n6173), .ZN(n5079)
         );
  AOI211_X1 U6248 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n5081), .A(n5080), 
        .B(n5079), .ZN(n5082) );
  OAI21_X1 U6249 ( .B1(n6206), .B2(n5101), .A(n5082), .ZN(U3010) );
  XOR2_X1 U6250 ( .A(n5084), .B(n5083), .Z(n6175) );
  INV_X1 U6251 ( .A(n6175), .ZN(n5089) );
  INV_X1 U6252 ( .A(n5085), .ZN(n6028) );
  NAND2_X1 U6253 ( .A1(n6133), .A2(REIP_REG_7__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U6254 ( .A1(n6148), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5086)
         );
  OAI211_X1 U6255 ( .C1(n6143), .C2(n6028), .A(n6171), .B(n5086), .ZN(n5087)
         );
  AOI21_X1 U6256 ( .B1(n6025), .B2(n6138), .A(n5087), .ZN(n5088) );
  OAI21_X1 U6257 ( .B1(n5089), .B2(n6145), .A(n5088), .ZN(U2979) );
  INV_X1 U6258 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6110) );
  OAI222_X1 U6259 ( .A1(n5119), .A2(n5524), .B1(n5299), .B2(n5090), .C1(n5507), 
        .C2(n6110), .ZN(U2882) );
  INV_X1 U6260 ( .A(n5052), .ZN(n5091) );
  AOI21_X1 U6261 ( .B1(n5092), .B2(n4912), .A(n5091), .ZN(n6014) );
  OAI22_X1 U6262 ( .A1(n5503), .A2(n6010), .B1(n6011), .B2(n6086), .ZN(n5093)
         );
  AOI21_X1 U6263 ( .B1(n6014), .B2(n6082), .A(n5093), .ZN(n5094) );
  INV_X1 U6264 ( .A(n5094), .ZN(U2851) );
  INV_X1 U6265 ( .A(n6014), .ZN(n5095) );
  INV_X1 U6266 ( .A(DATAI_8_), .ZN(n6619) );
  INV_X1 U6267 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6112) );
  OAI222_X1 U6268 ( .A1(n5095), .A2(n5524), .B1(n5299), .B2(n6619), .C1(n5507), 
        .C2(n6112), .ZN(U2883) );
  NAND2_X1 U6269 ( .A1(n6148), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5096)
         );
  OAI211_X1 U6270 ( .C1(n6143), .C2(n5098), .A(n5097), .B(n5096), .ZN(n5099)
         );
  AOI21_X1 U6271 ( .B1(n6014), .B2(n6138), .A(n5099), .ZN(n5100) );
  OAI21_X1 U6272 ( .B1(n6145), .B2(n5101), .A(n5100), .ZN(U2978) );
  INV_X1 U6273 ( .A(n5102), .ZN(n5103) );
  OAI21_X1 U6274 ( .B1(n6069), .B2(n5103), .A(n6068), .ZN(n6009) );
  NAND2_X1 U6275 ( .A1(n5103), .A2(n6518), .ZN(n5104) );
  NOR2_X1 U6276 ( .A1(n6069), .A2(n5104), .ZN(n6002) );
  INV_X1 U6277 ( .A(n6002), .ZN(n5105) );
  OAI21_X1 U6278 ( .B1(n5115), .B2(n6047), .A(n5105), .ZN(n5109) );
  AOI22_X1 U6279 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6050), .B1(n6066), .B2(n6162), 
        .ZN(n5106) );
  OAI211_X1 U6280 ( .C1(n6039), .C2(n5107), .A(n5106), .B(n6190), .ZN(n5108)
         );
  AOI211_X1 U6281 ( .C1(REIP_REG_9__SCAN_IN), .C2(n6009), .A(n5109), .B(n5108), 
        .ZN(n5110) );
  OAI21_X1 U6282 ( .B1(n5119), .B2(n5856), .A(n5110), .ZN(U2818) );
  INV_X1 U6283 ( .A(n5111), .ZN(n5112) );
  AOI21_X1 U6284 ( .B1(n5112), .B2(n3067), .A(n3018), .ZN(n6001) );
  INV_X1 U6285 ( .A(n6001), .ZN(n5181) );
  INV_X1 U6286 ( .A(DATAI_10_), .ZN(n6673) );
  INV_X1 U6287 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6108) );
  OAI222_X1 U6288 ( .A1(n5181), .A2(n5524), .B1(n5299), .B2(n6673), .C1(n5507), 
        .C2(n6108), .ZN(U2881) );
  XNOR2_X1 U6289 ( .A(n5618), .B(n6167), .ZN(n5114) );
  XNOR2_X1 U6290 ( .A(n5113), .B(n5114), .ZN(n6164) );
  NAND2_X1 U6291 ( .A1(n6164), .A2(n6137), .ZN(n5118) );
  AND2_X1 U6292 ( .A1(n6133), .A2(REIP_REG_9__SCAN_IN), .ZN(n6161) );
  NOR2_X1 U6293 ( .A1(n6143), .A2(n5115), .ZN(n5116) );
  AOI211_X1 U6294 ( .C1(n6148), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6161), 
        .B(n5116), .ZN(n5117) );
  OAI211_X1 U6295 ( .C1(n6371), .C2(n5119), .A(n5118), .B(n5117), .ZN(U2977)
         );
  NOR2_X1 U6296 ( .A1(n3018), .A2(n5122), .ZN(n5123) );
  OR2_X1 U6297 ( .A1(n5121), .A2(n5123), .ZN(n5257) );
  AOI21_X1 U6298 ( .B1(n5124), .B2(n5180), .A(n5186), .ZN(n6154) );
  AOI22_X1 U6299 ( .A1(n6081), .A2(n6154), .B1(n5485), .B2(EBX_REG_11__SCAN_IN), .ZN(n5125) );
  OAI21_X1 U6300 ( .B1(n5257), .B2(n5506), .A(n5125), .ZN(U2848) );
  NOR2_X1 U6301 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5126), .ZN(n5168)
         );
  INV_X1 U6302 ( .A(n5127), .ZN(n5131) );
  INV_X1 U6303 ( .A(n6236), .ZN(n5130) );
  INV_X1 U6304 ( .A(n5128), .ZN(n5129) );
  OR2_X1 U6305 ( .A1(n5205), .A2(n5129), .ZN(n6230) );
  OAI22_X1 U6306 ( .A1(n5131), .A2(n3017), .B1(n5130), .B2(n6230), .ZN(n5164)
         );
  INV_X1 U6307 ( .A(n6230), .ZN(n5133) );
  OAI21_X1 U6308 ( .B1(n5133), .B2(n4573), .A(n5132), .ZN(n6235) );
  NOR2_X1 U6309 ( .A1(n6235), .A2(n5203), .ZN(n5140) );
  NAND2_X1 U6310 ( .A1(n5166), .A2(n6280), .ZN(n5134) );
  NAND2_X1 U6311 ( .A1(n5134), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5138) );
  AOI21_X1 U6312 ( .B1(n5136), .B2(n5135), .A(n6587), .ZN(n5137) );
  NAND2_X1 U6313 ( .A1(n5138), .A2(n5137), .ZN(n5139) );
  AND2_X1 U6314 ( .A1(n5140), .A2(n5139), .ZN(n5141) );
  AOI22_X1 U6315 ( .A1(n5164), .A2(n6368), .B1(INSTQUEUE_REG_4__0__SCAN_IN), 
        .B2(n5163), .ZN(n5142) );
  OAI21_X1 U6316 ( .B1(n5166), .B2(n6382), .A(n5142), .ZN(n5143) );
  AOI21_X1 U6317 ( .B1(n6369), .B2(n5168), .A(n5143), .ZN(n5144) );
  OAI21_X1 U6318 ( .B1(n6242), .B2(n6280), .A(n5144), .ZN(U3052) );
  AOI22_X1 U6319 ( .A1(n5164), .A2(n6413), .B1(INSTQUEUE_REG_4__6__SCAN_IN), 
        .B2(n5163), .ZN(n5145) );
  OAI21_X1 U6320 ( .B1(n5166), .B2(n6418), .A(n5145), .ZN(n5146) );
  AOI21_X1 U6321 ( .B1(n6414), .B2(n5168), .A(n5146), .ZN(n5147) );
  OAI21_X1 U6322 ( .B1(n6260), .B2(n6280), .A(n5147), .ZN(U3058) );
  AOI22_X1 U6323 ( .A1(n5164), .A2(n6383), .B1(INSTQUEUE_REG_4__1__SCAN_IN), 
        .B2(n5163), .ZN(n5148) );
  OAI21_X1 U6324 ( .B1(n5166), .B2(n6388), .A(n5148), .ZN(n5149) );
  AOI21_X1 U6325 ( .B1(n6384), .B2(n5168), .A(n5149), .ZN(n5150) );
  OAI21_X1 U6326 ( .B1(n6245), .B2(n6280), .A(n5150), .ZN(U3053) );
  AOI22_X1 U6327 ( .A1(n5164), .A2(n6401), .B1(INSTQUEUE_REG_4__4__SCAN_IN), 
        .B2(n5163), .ZN(n5151) );
  OAI21_X1 U6328 ( .B1(n5166), .B2(n6406), .A(n5151), .ZN(n5152) );
  AOI21_X1 U6329 ( .B1(n6402), .B2(n5168), .A(n5152), .ZN(n5153) );
  OAI21_X1 U6330 ( .B1(n6254), .B2(n6280), .A(n5153), .ZN(U3056) );
  AOI22_X1 U6331 ( .A1(n5164), .A2(n6395), .B1(INSTQUEUE_REG_4__3__SCAN_IN), 
        .B2(n5163), .ZN(n5154) );
  OAI21_X1 U6332 ( .B1(n5166), .B2(n6400), .A(n5154), .ZN(n5155) );
  AOI21_X1 U6333 ( .B1(n6396), .B2(n5168), .A(n5155), .ZN(n5156) );
  OAI21_X1 U6334 ( .B1(n6251), .B2(n6280), .A(n5156), .ZN(U3055) );
  AOI22_X1 U6335 ( .A1(n5164), .A2(n6389), .B1(INSTQUEUE_REG_4__2__SCAN_IN), 
        .B2(n5163), .ZN(n5157) );
  OAI21_X1 U6336 ( .B1(n5166), .B2(n6394), .A(n5157), .ZN(n5158) );
  AOI21_X1 U6337 ( .B1(n6390), .B2(n5168), .A(n5158), .ZN(n5159) );
  OAI21_X1 U6338 ( .B1(n6248), .B2(n6280), .A(n5159), .ZN(U3054) );
  AOI22_X1 U6339 ( .A1(n5164), .A2(n6420), .B1(INSTQUEUE_REG_4__7__SCAN_IN), 
        .B2(n5163), .ZN(n5160) );
  OAI21_X1 U6340 ( .B1(n5166), .B2(n6429), .A(n5160), .ZN(n5161) );
  AOI21_X1 U6341 ( .B1(n6422), .B2(n5168), .A(n5161), .ZN(n5162) );
  OAI21_X1 U6342 ( .B1(n6267), .B2(n6280), .A(n5162), .ZN(U3059) );
  AOI22_X1 U6343 ( .A1(n5164), .A2(n6407), .B1(INSTQUEUE_REG_4__5__SCAN_IN), 
        .B2(n5163), .ZN(n5165) );
  OAI21_X1 U6344 ( .B1(n5166), .B2(n6412), .A(n5165), .ZN(n5167) );
  AOI21_X1 U6345 ( .B1(n6408), .B2(n5168), .A(n5167), .ZN(n5169) );
  OAI21_X1 U6346 ( .B1(n6257), .B2(n6280), .A(n5169), .ZN(U3057) );
  OAI21_X1 U6347 ( .B1(n6047), .B2(n5259), .A(n6190), .ZN(n5173) );
  INV_X1 U6348 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5171) );
  OAI22_X1 U6349 ( .A1(n5171), .A2(n6078), .B1(n5170), .B2(n6039), .ZN(n5172)
         );
  AOI211_X1 U6350 ( .C1(n6154), .C2(n6066), .A(n5173), .B(n5172), .ZN(n5176)
         );
  NOR2_X1 U6351 ( .A1(n6069), .A2(n5174), .ZN(n5193) );
  NOR2_X1 U6352 ( .A1(n5391), .A2(n5269), .ZN(n5190) );
  OAI21_X1 U6353 ( .B1(n5193), .B2(REIP_REG_11__SCAN_IN), .A(n5190), .ZN(n5175) );
  OAI211_X1 U6354 ( .C1(n5257), .C2(n5856), .A(n5176), .B(n5175), .ZN(U2816)
         );
  NAND2_X1 U6355 ( .A1(n5178), .A2(n5177), .ZN(n5179) );
  NAND2_X1 U6356 ( .A1(n5180), .A2(n5179), .ZN(n5997) );
  INV_X1 U6357 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5998) );
  OAI222_X1 U6358 ( .A1(n5997), .A2(n5503), .B1(n6086), .B2(n5998), .C1(n5181), 
        .C2(n5506), .ZN(U2849) );
  INV_X1 U6359 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6106) );
  OAI222_X1 U6360 ( .A1(n5257), .A2(n5524), .B1(n5299), .B2(n5182), .C1(n5507), 
        .C2(n6106), .ZN(U2880) );
  OAI21_X1 U6361 ( .B1(n5121), .B2(n5184), .A(n2987), .ZN(n5309) );
  NOR2_X1 U6362 ( .A1(n5186), .A2(n5185), .ZN(n5187) );
  OR2_X1 U6363 ( .A1(n3019), .A2(n5187), .ZN(n5293) );
  OAI22_X1 U6364 ( .A1(n5503), .A2(n5293), .B1(n5191), .B2(n6086), .ZN(n5188)
         );
  INV_X1 U6365 ( .A(n5188), .ZN(n5189) );
  OAI21_X1 U6366 ( .B1(n5309), .B2(n5506), .A(n5189), .ZN(U2847) );
  INV_X1 U6367 ( .A(n5190), .ZN(n5195) );
  INV_X1 U6368 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6524) );
  OAI22_X1 U6369 ( .A1(n5191), .A2(n6078), .B1(n6061), .B2(n5293), .ZN(n5192)
         );
  AOI211_X1 U6370 ( .C1(n6062), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6133), 
        .B(n5192), .ZN(n5194) );
  AND2_X1 U6371 ( .A1(n5193), .A2(REIP_REG_11__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6372 ( .A1(n5271), .A2(n6524), .ZN(n5268) );
  OAI211_X1 U6373 ( .C1(n5195), .C2(n6524), .A(n5194), .B(n5268), .ZN(n5196)
         );
  AOI21_X1 U6374 ( .B1(n5306), .B2(n6071), .A(n5196), .ZN(n5197) );
  OAI21_X1 U6375 ( .B1(n5309), .B2(n5856), .A(n5197), .ZN(U2815) );
  NAND2_X1 U6376 ( .A1(n6325), .A2(n6568), .ZN(n5200) );
  OAI21_X1 U6377 ( .B1(n5236), .B2(n5200), .A(n5199), .ZN(n5207) );
  INV_X1 U6378 ( .A(n5201), .ZN(n5202) );
  INV_X1 U6379 ( .A(n5203), .ZN(n6231) );
  NOR2_X1 U6380 ( .A1(n6231), .A2(n6572), .ZN(n5204) );
  NAND3_X1 U6381 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6441), .ZN(n6317) );
  NOR2_X1 U6382 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6317), .ZN(n5233)
         );
  INV_X1 U6383 ( .A(n5233), .ZN(n5208) );
  INV_X1 U6384 ( .A(n6316), .ZN(n5206) );
  AOI22_X1 U6385 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5208), .B1(n5207), .B2(
        n5206), .ZN(n5209) );
  OAI211_X1 U6386 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n4573), .A(n5210), .B(n5209), .ZN(n5232) );
  AOI22_X1 U6387 ( .A1(n6369), .A2(n5233), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5232), .ZN(n5211) );
  OAI21_X1 U6388 ( .B1(n6382), .B2(n6325), .A(n5211), .ZN(n5212) );
  AOI21_X1 U6389 ( .B1(n6379), .B2(n5236), .A(n5212), .ZN(n5213) );
  OAI21_X1 U6390 ( .B1(n5238), .B2(n6328), .A(n5213), .ZN(U3100) );
  AOI22_X1 U6391 ( .A1(n6414), .A2(n5233), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5232), .ZN(n5214) );
  OAI21_X1 U6392 ( .B1(n6418), .B2(n6325), .A(n5214), .ZN(n5215) );
  AOI21_X1 U6393 ( .B1(n5236), .B2(n6415), .A(n5215), .ZN(n5216) );
  OAI21_X1 U6394 ( .B1(n5238), .B2(n6352), .A(n5216), .ZN(U3106) );
  AOI22_X1 U6395 ( .A1(n6384), .A2(n5233), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5232), .ZN(n5217) );
  OAI21_X1 U6396 ( .B1(n6388), .B2(n6325), .A(n5217), .ZN(n5218) );
  AOI21_X1 U6397 ( .B1(n5236), .B2(n6385), .A(n5218), .ZN(n5219) );
  OAI21_X1 U6398 ( .B1(n5238), .B2(n6332), .A(n5219), .ZN(U3101) );
  AOI22_X1 U6399 ( .A1(n6402), .A2(n5233), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5232), .ZN(n5220) );
  OAI21_X1 U6400 ( .B1(n6406), .B2(n6325), .A(n5220), .ZN(n5221) );
  AOI21_X1 U6401 ( .B1(n5236), .B2(n6403), .A(n5221), .ZN(n5222) );
  OAI21_X1 U6402 ( .B1(n5238), .B2(n6344), .A(n5222), .ZN(U3104) );
  AOI22_X1 U6403 ( .A1(n6396), .A2(n5233), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5232), .ZN(n5223) );
  OAI21_X1 U6404 ( .B1(n6400), .B2(n6325), .A(n5223), .ZN(n5224) );
  AOI21_X1 U6405 ( .B1(n5236), .B2(n6397), .A(n5224), .ZN(n5225) );
  OAI21_X1 U6406 ( .B1(n5238), .B2(n6340), .A(n5225), .ZN(U3103) );
  AOI22_X1 U6407 ( .A1(n6390), .A2(n5233), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5232), .ZN(n5226) );
  OAI21_X1 U6408 ( .B1(n6394), .B2(n6325), .A(n5226), .ZN(n5227) );
  AOI21_X1 U6409 ( .B1(n5236), .B2(n6391), .A(n5227), .ZN(n5228) );
  OAI21_X1 U6410 ( .B1(n5238), .B2(n6336), .A(n5228), .ZN(U3102) );
  AOI22_X1 U6411 ( .A1(n6422), .A2(n5233), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5232), .ZN(n5229) );
  OAI21_X1 U6412 ( .B1(n6429), .B2(n6325), .A(n5229), .ZN(n5230) );
  AOI21_X1 U6413 ( .B1(n5236), .B2(n6424), .A(n5230), .ZN(n5231) );
  OAI21_X1 U6414 ( .B1(n5238), .B2(n6360), .A(n5231), .ZN(U3107) );
  AOI22_X1 U6415 ( .A1(n6408), .A2(n5233), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5232), .ZN(n5234) );
  OAI21_X1 U6416 ( .B1(n6412), .B2(n6325), .A(n5234), .ZN(n5235) );
  AOI21_X1 U6417 ( .B1(n5236), .B2(n6409), .A(n5235), .ZN(n5237) );
  OAI21_X1 U6418 ( .B1(n5238), .B2(n6348), .A(n5237), .ZN(U3105) );
  INV_X1 U6419 ( .A(n5252), .ZN(n5240) );
  AND2_X1 U6420 ( .A1(n5606), .A2(n5239), .ZN(n5253) );
  NOR2_X1 U6421 ( .A1(n5240), .A2(n5253), .ZN(n5242) );
  XOR2_X1 U6422 ( .A(n5242), .B(n2991), .Z(n5251) );
  INV_X1 U6423 ( .A(n6000), .ZN(n5244) );
  AOI22_X1 U6424 ( .A1(n6148), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6133), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5243) );
  OAI21_X1 U6425 ( .B1(n6143), .B2(n5244), .A(n5243), .ZN(n5245) );
  AOI21_X1 U6426 ( .B1(n6001), .B2(n6138), .A(n5245), .ZN(n5246) );
  OAI21_X1 U6427 ( .B1(n5251), .B2(n6145), .A(n5246), .ZN(U2976) );
  NOR2_X1 U6428 ( .A1(n5282), .A2(n6173), .ZN(n6163) );
  NAND2_X1 U6429 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5281) );
  OAI211_X1 U6430 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6163), .B(n5281), .ZN(n5250) );
  OAI21_X1 U6431 ( .B1(n5247), .B2(n5782), .A(n6178), .ZN(n6160) );
  INV_X1 U6432 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6521) );
  OAI22_X1 U6433 ( .A1(n6218), .A2(n5997), .B1(n6521), .B2(n6190), .ZN(n5248)
         );
  AOI21_X1 U6434 ( .B1(n6160), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5248), 
        .ZN(n5249) );
  OAI211_X1 U6435 ( .C1(n5251), .C2(n6206), .A(n5250), .B(n5249), .ZN(U3008)
         );
  INV_X1 U6436 ( .A(DATAI_12_), .ZN(n6731) );
  INV_X1 U6437 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6104) );
  OAI222_X1 U6438 ( .A1(n5309), .A2(n5524), .B1(n5299), .B2(n6731), .C1(n5507), 
        .C2(n6104), .ZN(U2879) );
  OAI21_X1 U6439 ( .B1(n2991), .B2(n5253), .A(n5252), .ZN(n5256) );
  OAI21_X1 U6440 ( .B1(n5571), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n5254), 
        .ZN(n5255) );
  XNOR2_X1 U6441 ( .A(n5256), .B(n5255), .ZN(n6155) );
  INV_X1 U6442 ( .A(n6155), .ZN(n5263) );
  INV_X1 U6443 ( .A(n5257), .ZN(n5261) );
  AOI22_X1 U6444 ( .A1(n6148), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n6133), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n5258) );
  OAI21_X1 U6445 ( .B1(n6143), .B2(n5259), .A(n5258), .ZN(n5260) );
  AOI21_X1 U6446 ( .B1(n5261), .B2(n6138), .A(n5260), .ZN(n5262) );
  OAI21_X1 U6447 ( .B1(n5263), .B2(n6145), .A(n5262), .ZN(U2975) );
  OAI21_X1 U6448 ( .B1(n5264), .B2(n5267), .A(n5266), .ZN(n5312) );
  OAI21_X1 U6449 ( .B1(n5391), .B2(n5269), .A(n5268), .ZN(n5276) );
  AOI21_X1 U6450 ( .B1(n6062), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6133), 
        .ZN(n5270) );
  OAI21_X1 U6451 ( .B1(n6047), .B2(n5314), .A(n5270), .ZN(n5275) );
  NAND2_X1 U6452 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5271), .ZN(n5428) );
  OAI21_X1 U6453 ( .B1(n3019), .B2(n5272), .A(n5416), .ZN(n5300) );
  INV_X1 U6454 ( .A(n5300), .ZN(n5949) );
  AOI22_X1 U6455 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6050), .B1(n6066), .B2(n5949), .ZN(n5273) );
  OAI21_X1 U6456 ( .B1(REIP_REG_13__SCAN_IN), .B2(n5428), .A(n5273), .ZN(n5274) );
  AOI211_X1 U6457 ( .C1(n5276), .C2(REIP_REG_13__SCAN_IN), .A(n5275), .B(n5274), .ZN(n5277) );
  OAI21_X1 U6458 ( .B1(n5312), .B2(n5856), .A(n5277), .ZN(U2814) );
  OAI21_X1 U6459 ( .B1(n3026), .B2(n5279), .A(n5278), .ZN(n5302) );
  INV_X1 U6460 ( .A(n5302), .ZN(n5298) );
  INV_X1 U6461 ( .A(n5280), .ZN(n5285) );
  NOR2_X1 U6462 ( .A1(n5282), .A2(n5281), .ZN(n5288) );
  NAND2_X1 U6463 ( .A1(n5283), .A2(n5288), .ZN(n5286) );
  AOI21_X1 U6464 ( .B1(n5285), .B2(n5286), .A(n5284), .ZN(n5935) );
  NOR2_X1 U6465 ( .A1(n6193), .A2(n5747), .ZN(n5291) );
  NAND2_X1 U6466 ( .A1(n5288), .A2(n5287), .ZN(n5292) );
  INV_X1 U6467 ( .A(n5292), .ZN(n5289) );
  OR2_X1 U6468 ( .A1(n5929), .A2(n5289), .ZN(n5933) );
  NAND2_X1 U6469 ( .A1(n5935), .A2(n5933), .ZN(n5290) );
  NOR2_X1 U6470 ( .A1(n6153), .A2(n5290), .ZN(n6159) );
  AOI211_X1 U6471 ( .C1(n5935), .C2(n5291), .A(n6159), .B(n2999), .ZN(n5296)
         );
  NOR2_X1 U6472 ( .A1(n5929), .A2(n5292), .ZN(n5936) );
  NOR3_X1 U6473 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6152), .A3(n6153), 
        .ZN(n5295) );
  NAND2_X1 U6474 ( .A1(n6133), .A2(REIP_REG_12__SCAN_IN), .ZN(n5303) );
  OAI21_X1 U6475 ( .B1(n6218), .B2(n5293), .A(n5303), .ZN(n5294) );
  NOR3_X1 U6476 ( .A1(n5296), .A2(n5295), .A3(n5294), .ZN(n5297) );
  OAI21_X1 U6477 ( .B1(n5298), .B2(n6206), .A(n5297), .ZN(U3006) );
  INV_X1 U6478 ( .A(DATAI_13_), .ZN(n6757) );
  INV_X1 U6479 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6102) );
  OAI222_X1 U6480 ( .A1(n5312), .A2(n5524), .B1(n5299), .B2(n6757), .C1(n6102), 
        .C2(n5507), .ZN(U2878) );
  INV_X1 U6481 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5301) );
  OAI222_X1 U6482 ( .A1(n5312), .A2(n5506), .B1(n5301), .B2(n5504), .C1(n5503), 
        .C2(n5300), .ZN(U2846) );
  NAND2_X1 U6483 ( .A1(n5302), .A2(n6137), .ZN(n5308) );
  INV_X1 U6484 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5304) );
  OAI21_X1 U6485 ( .B1(n5610), .B2(n5304), .A(n5303), .ZN(n5305) );
  AOI21_X1 U6486 ( .B1(n5613), .B2(n5306), .A(n5305), .ZN(n5307) );
  OAI211_X1 U6487 ( .C1(n6371), .C2(n5309), .A(n5308), .B(n5307), .ZN(U2974)
         );
  XNOR2_X1 U6488 ( .A(n5310), .B(n5311), .ZN(n5951) );
  INV_X1 U6489 ( .A(n5951), .ZN(n5318) );
  INV_X1 U6490 ( .A(n5312), .ZN(n5316) );
  AND2_X1 U6491 ( .A1(n6133), .A2(REIP_REG_13__SCAN_IN), .ZN(n5948) );
  AOI21_X1 U6492 ( .B1(n6148), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5948), 
        .ZN(n5313) );
  OAI21_X1 U6493 ( .B1(n6143), .B2(n5314), .A(n5313), .ZN(n5315) );
  AOI21_X1 U6494 ( .B1(n5316), .B2(n6138), .A(n5315), .ZN(n5317) );
  OAI21_X1 U6495 ( .B1(n6145), .B2(n5318), .A(n5317), .ZN(U2973) );
  INV_X1 U6496 ( .A(n5319), .ZN(n5321) );
  NOR2_X1 U6497 ( .A1(n5321), .A2(n5320), .ZN(n5324) );
  INV_X1 U6498 ( .A(n5322), .ZN(n5323) );
  AOI21_X1 U6499 ( .B1(n5324), .B2(n5266), .A(n5323), .ZN(n5639) );
  INV_X1 U6500 ( .A(n5639), .ZN(n5433) );
  XOR2_X1 U6501 ( .A(n5415), .B(n5416), .Z(n5939) );
  AOI22_X1 U6502 ( .A1(n5939), .A2(n6081), .B1(EBX_REG_14__SCAN_IN), .B2(n5485), .ZN(n5325) );
  OAI21_X1 U6503 ( .B1(n5433), .B2(n5506), .A(n5325), .ZN(U2845) );
  AOI22_X1 U6504 ( .A1(n5522), .A2(DATAI_14_), .B1(n6093), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5326) );
  OAI21_X1 U6505 ( .B1(n5433), .B2(n5524), .A(n5326), .ZN(U2877) );
  INV_X1 U6506 ( .A(n4392), .ZN(n5328) );
  AOI21_X1 U6507 ( .B1(n5328), .B2(n5327), .A(n5335), .ZN(n5337) );
  NOR3_X1 U6508 ( .A1(n5328), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6467), 
        .ZN(n5331) );
  NOR2_X1 U6509 ( .A1(n5329), .A2(n5806), .ZN(n5330) );
  AOI211_X1 U6510 ( .C1(n5333), .C2(n5332), .A(n5331), .B(n5330), .ZN(n5334)
         );
  OAI22_X1 U6511 ( .A1(n5337), .A2(n5336), .B1(n5335), .B2(n5334), .ZN(U3459)
         );
  NOR3_X4 U6512 ( .A1(n6093), .A2(n4246), .A3(n5338), .ZN(n6094) );
  AOI22_X1 U6513 ( .A1(n6094), .A2(DATAI_12_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6093), .ZN(n5341) );
  AND2_X1 U6514 ( .A1(n5507), .A2(n5339), .ZN(n6090) );
  NAND2_X1 U6515 ( .A1(n6090), .A2(DATAI_28_), .ZN(n5340) );
  OAI211_X1 U6516 ( .C1(n5543), .C2(n5524), .A(n5341), .B(n5340), .ZN(U2863)
         );
  INV_X1 U6517 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5342) );
  OAI222_X1 U6518 ( .A1(n5506), .A2(n5543), .B1(n6086), .B2(n5342), .C1(n5682), 
        .C2(n5503), .ZN(U2831) );
  OAI21_X1 U6519 ( .B1(n6069), .B2(n6053), .A(n6068), .ZN(n6049) );
  AOI22_X1 U6520 ( .A1(EBX_REG_3__SCAN_IN), .A2(n6050), .B1(n6064), .B2(n3017), 
        .ZN(n5350) );
  INV_X1 U6521 ( .A(n6180), .ZN(n5343) );
  NAND2_X1 U6522 ( .A1(n6066), .A2(n5343), .ZN(n5349) );
  INV_X1 U6523 ( .A(n5344), .ZN(n5345) );
  AOI22_X1 U6524 ( .A1(n6062), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n6071), 
        .B2(n5345), .ZN(n5348) );
  INV_X1 U6525 ( .A(n6053), .ZN(n5346) );
  NAND4_X1 U6526 ( .A1(n6054), .A2(REIP_REG_1__SCAN_IN), .A3(n5346), .A4(
        REIP_REG_2__SCAN_IN), .ZN(n5347) );
  NAND4_X1 U6527 ( .A1(n5350), .A2(n5349), .A3(n5348), .A4(n5347), .ZN(n5351)
         );
  AOI21_X1 U6528 ( .B1(REIP_REG_3__SCAN_IN), .B2(n6049), .A(n5351), .ZN(n5352)
         );
  OAI21_X1 U6529 ( .B1(n5354), .B2(n5353), .A(n5352), .ZN(U2824) );
  INV_X1 U6530 ( .A(n5509), .ZN(n5374) );
  OAI22_X1 U6531 ( .A1(n5359), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n5358), .B2(EBX_REG_31__SCAN_IN), .ZN(n5360) );
  INV_X1 U6532 ( .A(n5362), .ZN(n5367) );
  NAND2_X1 U6533 ( .A1(n6062), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5365)
         );
  INV_X1 U6534 ( .A(REIP_REG_31__SCAN_IN), .ZN(n5363) );
  NAND4_X1 U6535 ( .A1(n5363), .A2(REIP_REG_30__SCAN_IN), .A3(
        REIP_REG_29__SCAN_IN), .A4(n5378), .ZN(n5364) );
  OAI211_X1 U6536 ( .C1(n5367), .C2(n5366), .A(n5365), .B(n5364), .ZN(n5368)
         );
  AOI21_X1 U6537 ( .B1(n5369), .B2(n6066), .A(n5368), .ZN(n5373) );
  NAND3_X1 U6538 ( .A1(n5371), .A2(REIP_REG_30__SCAN_IN), .A3(n5370), .ZN(
        n5379) );
  NAND3_X1 U6539 ( .A1(n5379), .A2(REIP_REG_31__SCAN_IN), .A3(n5864), .ZN(
        n5372) );
  OAI211_X1 U6540 ( .C1(n5374), .C2(n5856), .A(n5373), .B(n5372), .ZN(U2796)
         );
  INV_X1 U6541 ( .A(n5375), .ZN(n5534) );
  OAI22_X1 U6542 ( .A1(n5376), .A2(n6039), .B1(n6047), .B2(n5534), .ZN(n5377)
         );
  AND2_X1 U6543 ( .A1(REIP_REG_29__SCAN_IN), .A2(n5378), .ZN(n5380) );
  OAI21_X1 U6544 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5380), .A(n5379), .ZN(n5381) );
  INV_X1 U6545 ( .A(n3021), .ZN(n5383) );
  OAI22_X1 U6546 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5385), .B1(n5904), .B2(
        n6047), .ZN(n5396) );
  INV_X1 U6547 ( .A(n5453), .ZN(n5387) );
  AOI21_X1 U6548 ( .B1(n5387), .B2(n5443), .A(n5386), .ZN(n5389) );
  OR2_X1 U6549 ( .A1(n5389), .A2(n5388), .ZN(n5914) );
  NOR2_X1 U6550 ( .A1(n5391), .A2(n5390), .ZN(n5830) );
  NOR2_X1 U6551 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5392), .ZN(n5820) );
  OAI21_X1 U6552 ( .B1(n5830), .B2(n5820), .A(REIP_REG_25__SCAN_IN), .ZN(n5394) );
  AOI22_X1 U6553 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6050), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6062), .ZN(n5393) );
  OAI211_X1 U6554 ( .C1(n6061), .C2(n5914), .A(n5394), .B(n5393), .ZN(n5395)
         );
  AOI211_X1 U6555 ( .C1(n5901), .C2(n6033), .A(n5396), .B(n5395), .ZN(n5397)
         );
  INV_X1 U6556 ( .A(n5397), .ZN(U2802) );
  OR2_X1 U6557 ( .A1(n5399), .A2(n5400), .ZN(n5401) );
  NAND2_X1 U6558 ( .A1(n5398), .A2(n5401), .ZN(n5616) );
  MUX2_X1 U6559 ( .A(n5472), .B(n5402), .S(n3904), .Z(n5481) );
  OR2_X1 U6560 ( .A1(n5492), .A2(n5481), .ZN(n5479) );
  INV_X1 U6561 ( .A(n5479), .ZN(n5403) );
  AOI21_X1 U6562 ( .B1(n5492), .B2(n5481), .A(n5403), .ZN(n5924) );
  NAND4_X1 U6563 ( .A1(n5412), .A2(n6054), .A3(REIP_REG_17__SCAN_IN), .A4(
        REIP_REG_16__SCAN_IN), .ZN(n5853) );
  NOR2_X1 U6564 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5853), .ZN(n5862) );
  AOI21_X1 U6565 ( .B1(n6071), .B2(n5612), .A(n5862), .ZN(n5404) );
  OAI21_X1 U6566 ( .B1(n6078), .B2(n5405), .A(n5404), .ZN(n5408) );
  NAND2_X1 U6567 ( .A1(n5864), .A2(n5863), .ZN(n5980) );
  INV_X1 U6568 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6534) );
  NAND2_X1 U6569 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n6062), .ZN(n5406)
         );
  OAI211_X1 U6570 ( .C1(n5980), .C2(n6534), .A(n6190), .B(n5406), .ZN(n5407)
         );
  AOI211_X1 U6571 ( .C1(n5924), .C2(n6066), .A(n5408), .B(n5407), .ZN(n5409)
         );
  OAI21_X1 U6572 ( .B1(n5616), .B2(n5856), .A(n5409), .ZN(U2809) );
  AOI21_X1 U6573 ( .B1(n5411), .B2(n5322), .A(n3697), .ZN(n5629) );
  INV_X1 U6574 ( .A(n5629), .ZN(n5525) );
  INV_X1 U6575 ( .A(n5412), .ZN(n5978) );
  NAND2_X1 U6576 ( .A1(n5864), .A2(n5978), .ZN(n5990) );
  AOI21_X1 U6577 ( .B1(n6528), .B2(n5429), .A(n5990), .ZN(n5422) );
  OAI21_X1 U6578 ( .B1(n6039), .B2(n5413), .A(n6190), .ZN(n5421) );
  OAI21_X1 U6579 ( .B1(n5416), .B2(n5415), .A(n5414), .ZN(n5417) );
  NAND2_X1 U6580 ( .A1(n5417), .A2(n5496), .ZN(n5792) );
  AOI22_X1 U6581 ( .A1(n6050), .A2(EBX_REG_15__SCAN_IN), .B1(n6071), .B2(n5418), .ZN(n5419) );
  OAI21_X1 U6582 ( .B1(n6061), .B2(n5792), .A(n5419), .ZN(n5420) );
  NOR3_X1 U6583 ( .A1(n5422), .A2(n5421), .A3(n5420), .ZN(n5423) );
  OAI21_X1 U6584 ( .B1(n5525), .B2(n5856), .A(n5423), .ZN(U2812) );
  INV_X1 U6585 ( .A(n5637), .ZN(n5427) );
  INV_X1 U6586 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5425) );
  AOI22_X1 U6587 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6050), .B1(n6066), .B2(n5939), .ZN(n5424) );
  OAI211_X1 U6588 ( .C1(n6039), .C2(n5425), .A(n5424), .B(n6190), .ZN(n5426)
         );
  AOI21_X1 U6589 ( .B1(n6071), .B2(n5427), .A(n5426), .ZN(n5432) );
  INV_X1 U6590 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6526) );
  NOR2_X1 U6591 ( .A1(n6526), .A2(n5428), .ZN(n5430) );
  OAI211_X1 U6592 ( .C1(n5430), .C2(REIP_REG_14__SCAN_IN), .A(n5429), .B(n5864), .ZN(n5431) );
  OAI211_X1 U6593 ( .C1(n5433), .C2(n5856), .A(n5432), .B(n5431), .ZN(U2813)
         );
  OAI22_X1 U6594 ( .A1(n5659), .A2(n5503), .B1(n6086), .B2(n5434), .ZN(U2828)
         );
  OAI222_X1 U6595 ( .A1(n5506), .A2(n4286), .B1(n5435), .B2(n5504), .C1(n5674), 
        .C2(n5503), .ZN(U2830) );
  INV_X1 U6596 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5436) );
  OAI222_X1 U6597 ( .A1(n5517), .A2(n5506), .B1(n6086), .B2(n5436), .C1(n5710), 
        .C2(n5503), .ZN(U2833) );
  INV_X1 U6598 ( .A(n5901), .ZN(n5438) );
  OAI222_X1 U6599 ( .A1(n5438), .A2(n5506), .B1(n5437), .B2(n5504), .C1(n5503), 
        .C2(n5914), .ZN(U2834) );
  AOI21_X1 U6600 ( .B1(n5442), .B2(n5440), .A(n5382), .ZN(n5884) );
  INV_X1 U6601 ( .A(n5884), .ZN(n5446) );
  XNOR2_X1 U6602 ( .A(n5453), .B(n5443), .ZN(n5819) );
  INV_X1 U6603 ( .A(n5819), .ZN(n5444) );
  OAI222_X1 U6604 ( .A1(n5506), .A2(n5446), .B1(n5445), .B2(n6086), .C1(n5503), 
        .C2(n5444), .ZN(U2835) );
  OR2_X1 U6605 ( .A1(n5447), .A2(n5448), .ZN(n5449) );
  AND2_X1 U6606 ( .A1(n5440), .A2(n5449), .ZN(n5887) );
  INV_X1 U6607 ( .A(n5887), .ZN(n5455) );
  INV_X1 U6608 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U6609 ( .A1(n5450), .A2(n5451), .ZN(n5452) );
  NAND2_X1 U6610 ( .A1(n5453), .A2(n5452), .ZN(n5828) );
  OAI222_X1 U6611 ( .A1(n5506), .A2(n5455), .B1(n5454), .B2(n6086), .C1(n5828), 
        .C2(n5503), .ZN(U2836) );
  OAI21_X1 U6612 ( .B1(n5457), .B2(n5456), .A(n5450), .ZN(n5838) );
  INV_X1 U6613 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5461) );
  INV_X1 U6614 ( .A(n5447), .ZN(n5459) );
  OAI21_X1 U6615 ( .B1(n5460), .B2(n5458), .A(n5459), .ZN(n5839) );
  OAI222_X1 U6616 ( .A1(n5503), .A2(n5838), .B1(n6086), .B2(n5461), .C1(n5839), 
        .C2(n5506), .ZN(U2837) );
  OR2_X1 U6617 ( .A1(n5462), .A2(n5470), .ZN(n5463) );
  AOI21_X1 U6618 ( .B1(n5464), .B2(n5463), .A(n5458), .ZN(n5890) );
  XNOR2_X1 U6619 ( .A(n5466), .B(n5465), .ZN(n5851) );
  OAI22_X1 U6620 ( .A1(n5851), .A2(n5503), .B1(n5467), .B2(n6086), .ZN(n5468)
         );
  AOI21_X1 U6621 ( .B1(n5890), .B2(n6082), .A(n5468), .ZN(n5469) );
  INV_X1 U6622 ( .A(n5469), .ZN(U2838) );
  XNOR2_X1 U6623 ( .A(n5462), .B(n5470), .ZN(n5893) );
  MUX2_X1 U6624 ( .A(n5472), .B(n4296), .S(n5471), .Z(n5474) );
  XNOR2_X1 U6625 ( .A(n5474), .B(n5473), .ZN(n5858) );
  INV_X1 U6626 ( .A(n5858), .ZN(n5754) );
  OAI222_X1 U6627 ( .A1(n5893), .A2(n5506), .B1(n5475), .B2(n5504), .C1(n5503), 
        .C2(n5754), .ZN(U2839) );
  NAND2_X1 U6628 ( .A1(n5398), .A2(n5476), .ZN(n5477) );
  NAND2_X1 U6629 ( .A1(n5479), .A2(n5478), .ZN(n5480) );
  OAI21_X1 U6630 ( .B1(n5471), .B2(n5481), .A(n5480), .ZN(n5872) );
  OAI22_X1 U6631 ( .A1(n5872), .A2(n5503), .B1(n5482), .B2(n6086), .ZN(n5483)
         );
  AOI21_X1 U6632 ( .B1(n5905), .B2(n6082), .A(n5483), .ZN(n5484) );
  INV_X1 U6633 ( .A(n5484), .ZN(U2840) );
  AOI22_X1 U6634 ( .A1(n5924), .A2(n6081), .B1(EBX_REG_18__SCAN_IN), .B2(n5485), .ZN(n5486) );
  OAI21_X1 U6635 ( .B1(n5616), .B2(n5506), .A(n5486), .ZN(U2841) );
  AND2_X1 U6636 ( .A1(n2989), .A2(n5488), .ZN(n5489) );
  NOR2_X1 U6637 ( .A1(n5399), .A2(n5489), .ZN(n6087) );
  INV_X1 U6638 ( .A(n6087), .ZN(n5494) );
  OR2_X1 U6639 ( .A1(n5497), .A2(n5490), .ZN(n5491) );
  NAND2_X1 U6640 ( .A1(n5492), .A2(n5491), .ZN(n5983) );
  OAI222_X1 U6641 ( .A1(n5494), .A2(n5506), .B1(n5493), .B2(n5504), .C1(n5503), 
        .C2(n5983), .ZN(U2842) );
  AND2_X1 U6642 ( .A1(n5496), .A2(n5495), .ZN(n5498) );
  OR2_X1 U6643 ( .A1(n5498), .A2(n5497), .ZN(n5996) );
  INV_X1 U6644 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5502) );
  INV_X1 U6645 ( .A(n5487), .ZN(n5499) );
  AOI21_X1 U6646 ( .B1(n5500), .B2(n5410), .A(n5499), .ZN(n6092) );
  INV_X1 U6647 ( .A(n6092), .ZN(n5501) );
  OAI222_X1 U6648 ( .A1(n5996), .A2(n5503), .B1(n6086), .B2(n5502), .C1(n5501), 
        .C2(n5506), .ZN(U2843) );
  INV_X1 U6649 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5505) );
  OAI222_X1 U6650 ( .A1(n5525), .A2(n5506), .B1(n5505), .B2(n5504), .C1(n5792), 
        .C2(n5503), .ZN(U2844) );
  AND2_X1 U6651 ( .A1(n5507), .A2(n4246), .ZN(n5508) );
  NAND2_X1 U6652 ( .A1(n5509), .A2(n5508), .ZN(n5511) );
  AOI22_X1 U6653 ( .A1(n6090), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6093), .ZN(n5510) );
  NAND2_X1 U6654 ( .A1(n5511), .A2(n5510), .ZN(U2860) );
  AOI22_X1 U6655 ( .A1(n6090), .A2(DATAI_30_), .B1(n6093), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U6656 ( .A1(n6094), .A2(DATAI_14_), .ZN(n5512) );
  OAI211_X1 U6657 ( .C1(n5514), .C2(n5524), .A(n5513), .B(n5512), .ZN(U2861)
         );
  AOI22_X1 U6658 ( .A1(n6094), .A2(DATAI_10_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6093), .ZN(n5516) );
  NAND2_X1 U6659 ( .A1(n6090), .A2(DATAI_26_), .ZN(n5515) );
  OAI211_X1 U6660 ( .C1(n5517), .C2(n5524), .A(n5516), .B(n5515), .ZN(U2865)
         );
  AOI22_X1 U6661 ( .A1(n6094), .A2(DATAI_6_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n6093), .ZN(n5519) );
  NAND2_X1 U6662 ( .A1(n6090), .A2(DATAI_22_), .ZN(n5518) );
  OAI211_X1 U6663 ( .C1(n5839), .C2(n5524), .A(n5519), .B(n5518), .ZN(U2869)
         );
  AOI22_X1 U6664 ( .A1(n6090), .A2(DATAI_18_), .B1(n6093), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U6665 ( .A1(n6094), .A2(DATAI_2_), .ZN(n5520) );
  OAI211_X1 U6666 ( .C1(n5616), .C2(n5524), .A(n5521), .B(n5520), .ZN(U2873)
         );
  AOI22_X1 U6667 ( .A1(n5522), .A2(DATAI_15_), .B1(n6093), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5523) );
  OAI21_X1 U6668 ( .B1(n5525), .B2(n5524), .A(n5523), .ZN(U2876) );
  INV_X1 U6669 ( .A(n5526), .ZN(n5528) );
  NAND2_X1 U6670 ( .A1(n5528), .A2(n5527), .ZN(n5531) );
  NAND2_X1 U6671 ( .A1(n5529), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U6672 ( .A1(n5531), .A2(n5530), .ZN(n5532) );
  XNOR2_X1 U6673 ( .A(n5532), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5673)
         );
  AND2_X1 U6674 ( .A1(n6133), .A2(REIP_REG_30__SCAN_IN), .ZN(n5665) );
  AOI21_X1 U6675 ( .B1(n6148), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5665), 
        .ZN(n5533) );
  OAI21_X1 U6676 ( .B1(n6143), .B2(n5534), .A(n5533), .ZN(n5535) );
  AOI21_X1 U6677 ( .B1(n5536), .B2(n6138), .A(n5535), .ZN(n5537) );
  OAI21_X1 U6678 ( .B1(n5673), .B2(n6145), .A(n5537), .ZN(U2956) );
  NAND3_X1 U6679 ( .A1(n5559), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5606), .ZN(n5541) );
  NAND2_X1 U6680 ( .A1(n5919), .A2(n5540), .ZN(n5705) );
  OR2_X1 U6681 ( .A1(n5606), .A2(n5705), .ZN(n5538) );
  XNOR2_X1 U6682 ( .A(n5542), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5691)
         );
  INV_X1 U6683 ( .A(n5543), .ZN(n5548) );
  INV_X1 U6684 ( .A(n5544), .ZN(n5546) );
  AND2_X1 U6685 ( .A1(n6133), .A2(REIP_REG_28__SCAN_IN), .ZN(n5686) );
  AOI21_X1 U6686 ( .B1(n6148), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5686), 
        .ZN(n5545) );
  OAI21_X1 U6687 ( .B1(n6143), .B2(n5546), .A(n5545), .ZN(n5547) );
  AOI21_X1 U6688 ( .B1(n5548), .B2(n6138), .A(n5547), .ZN(n5549) );
  OAI21_X1 U6689 ( .B1(n6145), .B2(n5691), .A(n5549), .ZN(U2958) );
  NAND2_X1 U6690 ( .A1(n5551), .A2(n5550), .ZN(n5552) );
  XNOR2_X1 U6691 ( .A(n5552), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5703)
         );
  OR2_X1 U6692 ( .A1(n4132), .A2(n5553), .ZN(n5555) );
  AND2_X1 U6693 ( .A1(n6133), .A2(REIP_REG_27__SCAN_IN), .ZN(n5696) );
  AOI21_X1 U6694 ( .B1(n6148), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5696), 
        .ZN(n5556) );
  OAI21_X1 U6695 ( .B1(n6143), .B2(n5811), .A(n5556), .ZN(n5557) );
  AOI21_X1 U6696 ( .B1(n5879), .B2(n6138), .A(n5557), .ZN(n5558) );
  OAI21_X1 U6697 ( .B1(n5703), .B2(n6145), .A(n5558), .ZN(U2959) );
  XNOR2_X1 U6698 ( .A(n5618), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5560)
         );
  XNOR2_X1 U6699 ( .A(n5559), .B(n5560), .ZN(n5714) );
  INV_X1 U6700 ( .A(n5561), .ZN(n5563) );
  AND2_X1 U6701 ( .A1(n6133), .A2(REIP_REG_26__SCAN_IN), .ZN(n5707) );
  AOI21_X1 U6702 ( .B1(n6148), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5707), 
        .ZN(n5562) );
  OAI21_X1 U6703 ( .B1(n6143), .B2(n5563), .A(n5562), .ZN(n5564) );
  AOI21_X1 U6704 ( .B1(n5565), .B2(n6138), .A(n5564), .ZN(n5566) );
  OAI21_X1 U6705 ( .B1(n6145), .B2(n5714), .A(n5566), .ZN(U2960) );
  NAND2_X1 U6706 ( .A1(n5758), .A2(n3959), .ZN(n5569) );
  AOI21_X1 U6707 ( .B1(n5569), .B2(n5571), .A(n5568), .ZN(n5599) );
  XOR2_X1 U6708 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .B(n5618), .Z(n5600) );
  NOR2_X1 U6709 ( .A1(n2992), .A2(n3080), .ZN(n5592) );
  XNOR2_X1 U6710 ( .A(n5618), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5594)
         );
  INV_X1 U6711 ( .A(n5593), .ZN(n5570) );
  NOR2_X1 U6712 ( .A1(n5618), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5585)
         );
  NAND2_X1 U6713 ( .A1(n5570), .A2(n5585), .ZN(n5579) );
  OAI21_X1 U6714 ( .B1(n5571), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5593), 
        .ZN(n5587) );
  NAND3_X1 U6715 ( .A1(n5606), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5572) );
  XNOR2_X1 U6716 ( .A(n5573), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5722)
         );
  INV_X1 U6717 ( .A(n5818), .ZN(n5575) );
  AND2_X1 U6718 ( .A1(n6133), .A2(REIP_REG_24__SCAN_IN), .ZN(n5720) );
  AOI21_X1 U6719 ( .B1(n6148), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5720), 
        .ZN(n5574) );
  OAI21_X1 U6720 ( .B1(n6143), .B2(n5575), .A(n5574), .ZN(n5576) );
  AOI21_X1 U6721 ( .B1(n5884), .B2(n6138), .A(n5576), .ZN(n5577) );
  OAI21_X1 U6722 ( .B1(n5722), .B2(n6145), .A(n5577), .ZN(U2962) );
  INV_X1 U6723 ( .A(n5578), .ZN(n5580) );
  OAI21_X1 U6724 ( .B1(n5580), .B2(n5715), .A(n5579), .ZN(n5581) );
  XNOR2_X1 U6725 ( .A(n5581), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5729)
         );
  NAND2_X1 U6726 ( .A1(n6133), .A2(REIP_REG_23__SCAN_IN), .ZN(n5723) );
  NAND2_X1 U6727 ( .A1(n6148), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5582)
         );
  OAI211_X1 U6728 ( .C1(n6143), .C2(n5825), .A(n5723), .B(n5582), .ZN(n5583)
         );
  AOI21_X1 U6729 ( .B1(n5887), .B2(n6138), .A(n5583), .ZN(n5584) );
  OAI21_X1 U6730 ( .B1(n5729), .B2(n6145), .A(n5584), .ZN(U2963) );
  AOI21_X1 U6731 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5618), .A(n5585), 
        .ZN(n5586) );
  XNOR2_X1 U6732 ( .A(n5587), .B(n5586), .ZN(n5737) );
  NAND2_X1 U6733 ( .A1(n6133), .A2(REIP_REG_22__SCAN_IN), .ZN(n5731) );
  OAI21_X1 U6734 ( .B1(n5610), .B2(n5588), .A(n5731), .ZN(n5590) );
  NOR2_X1 U6735 ( .A1(n5839), .A2(n6371), .ZN(n5589) );
  AOI211_X1 U6736 ( .C1(n5613), .C2(n5842), .A(n5590), .B(n5589), .ZN(n5591)
         );
  OAI21_X1 U6737 ( .B1(n5737), .B2(n6145), .A(n5591), .ZN(U2964) );
  OAI21_X1 U6738 ( .B1(n5592), .B2(n5594), .A(n5593), .ZN(n5595) );
  INV_X1 U6739 ( .A(n5595), .ZN(n5745) );
  NAND2_X1 U6740 ( .A1(n6133), .A2(REIP_REG_21__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U6741 ( .A1(n6148), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5596)
         );
  OAI211_X1 U6742 ( .C1(n6143), .C2(n5846), .A(n5739), .B(n5596), .ZN(n5597)
         );
  AOI21_X1 U6743 ( .B1(n5890), .B2(n6138), .A(n5597), .ZN(n5598) );
  OAI21_X1 U6744 ( .B1(n5745), .B2(n6145), .A(n5598), .ZN(U2965) );
  AOI21_X1 U6745 ( .B1(n5599), .B2(n5600), .A(n5578), .ZN(n5746) );
  NAND2_X1 U6746 ( .A1(n5746), .A2(n6137), .ZN(n5603) );
  NAND2_X1 U6747 ( .A1(n6133), .A2(REIP_REG_20__SCAN_IN), .ZN(n5753) );
  OAI21_X1 U6748 ( .B1(n5610), .B2(n5861), .A(n5753), .ZN(n5601) );
  AOI21_X1 U6749 ( .B1(n5613), .B2(n5852), .A(n5601), .ZN(n5602) );
  OAI211_X1 U6750 ( .C1(n6371), .C2(n5893), .A(n5603), .B(n5602), .ZN(U2966)
         );
  NAND3_X1 U6751 ( .A1(n5604), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5606), .ZN(n5770) );
  INV_X1 U6752 ( .A(n3059), .ZN(n5607) );
  NOR2_X1 U6753 ( .A1(n5606), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5769)
         );
  NAND3_X1 U6754 ( .A1(n5607), .A2(n5769), .A3(n5921), .ZN(n5772) );
  NAND2_X1 U6755 ( .A1(n5770), .A2(n5772), .ZN(n5609) );
  XNOR2_X1 U6756 ( .A(n5609), .B(n5608), .ZN(n5925) );
  NAND2_X1 U6757 ( .A1(n5925), .A2(n6137), .ZN(n5615) );
  OAI22_X1 U6758 ( .A1(n5610), .A2(n3197), .B1(n6190), .B2(n6534), .ZN(n5611)
         );
  AOI21_X1 U6759 ( .B1(n5613), .B2(n5612), .A(n5611), .ZN(n5614) );
  OAI211_X1 U6760 ( .C1(n6371), .C2(n5616), .A(n5615), .B(n5614), .ZN(U2968)
         );
  XNOR2_X1 U6761 ( .A(n5618), .B(n5780), .ZN(n5619) );
  XNOR2_X1 U6762 ( .A(n5617), .B(n5619), .ZN(n5788) );
  NAND2_X1 U6763 ( .A1(n6133), .A2(REIP_REG_16__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U6764 ( .A1(n6148), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5620)
         );
  OAI211_X1 U6765 ( .C1(n6143), .C2(n5992), .A(n5783), .B(n5620), .ZN(n5621)
         );
  AOI21_X1 U6766 ( .B1(n6092), .B2(n6138), .A(n5621), .ZN(n5622) );
  OAI21_X1 U6767 ( .B1(n6145), .B2(n5788), .A(n5622), .ZN(U2970) );
  OAI21_X1 U6768 ( .B1(n5623), .B2(n5624), .A(n3059), .ZN(n5625) );
  INV_X1 U6769 ( .A(n5625), .ZN(n5797) );
  NAND2_X1 U6770 ( .A1(n6133), .A2(REIP_REG_15__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U6771 ( .A1(n6148), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5626)
         );
  OAI211_X1 U6772 ( .C1(n6143), .C2(n5627), .A(n5790), .B(n5626), .ZN(n5628)
         );
  AOI21_X1 U6773 ( .B1(n5629), .B2(n6138), .A(n5628), .ZN(n5630) );
  OAI21_X1 U6774 ( .B1(n5797), .B2(n6145), .A(n5630), .ZN(U2971) );
  INV_X1 U6775 ( .A(n5632), .ZN(n5634) );
  NOR2_X1 U6776 ( .A1(n5634), .A2(n5633), .ZN(n5635) );
  XNOR2_X1 U6777 ( .A(n3007), .B(n5635), .ZN(n5942) );
  INV_X1 U6778 ( .A(n5942), .ZN(n5641) );
  AND2_X1 U6779 ( .A1(n6133), .A2(REIP_REG_14__SCAN_IN), .ZN(n5938) );
  AOI21_X1 U6780 ( .B1(n6148), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5938), 
        .ZN(n5636) );
  OAI21_X1 U6781 ( .B1(n6143), .B2(n5637), .A(n5636), .ZN(n5638) );
  AOI21_X1 U6782 ( .B1(n5639), .B2(n6138), .A(n5638), .ZN(n5640) );
  OAI21_X1 U6783 ( .B1(n6145), .B2(n5641), .A(n5640), .ZN(U2972) );
  INV_X1 U6784 ( .A(n5656), .ZN(n5683) );
  NAND2_X1 U6785 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5706) );
  NAND3_X1 U6786 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5940) );
  NOR2_X1 U6787 ( .A1(n5945), .A2(n5940), .ZN(n5781) );
  NAND3_X1 U6788 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5781), .ZN(n5646) );
  INV_X1 U6789 ( .A(n5642), .ZN(n5649) );
  NAND2_X1 U6790 ( .A1(n5923), .A2(n5649), .ZN(n5748) );
  INV_X1 U6791 ( .A(n5648), .ZN(n5751) );
  NOR2_X1 U6792 ( .A1(n5748), .A2(n5751), .ZN(n5743) );
  INV_X1 U6793 ( .A(n5643), .ZN(n5644) );
  NAND2_X1 U6794 ( .A1(n5743), .A2(n5644), .ZN(n5732) );
  INV_X1 U6795 ( .A(n5933), .ZN(n5645) );
  OAI21_X1 U6796 ( .B1(n5646), .B2(n5645), .A(n6212), .ZN(n5647) );
  NAND2_X1 U6797 ( .A1(n5935), .A2(n5647), .ZN(n5776) );
  AND2_X1 U6798 ( .A1(n5649), .A2(n5648), .ZN(n5650) );
  NOR2_X1 U6799 ( .A1(n5782), .A2(n5650), .ZN(n5651) );
  NOR2_X1 U6800 ( .A1(n5776), .A2(n5651), .ZN(n5738) );
  NAND2_X1 U6801 ( .A1(n6198), .A2(n5929), .ZN(n5652) );
  NAND2_X1 U6802 ( .A1(n5652), .A2(n5654), .ZN(n5653) );
  AOI21_X1 U6803 ( .B1(n6212), .B2(n5706), .A(n5712), .ZN(n5688) );
  OAI21_X1 U6804 ( .B1(n5782), .B2(n5683), .A(n5688), .ZN(n5678) );
  AOI21_X1 U6805 ( .B1(n6212), .B2(n5527), .A(n5678), .ZN(n5664) );
  OAI21_X1 U6806 ( .B1(n5782), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5664), 
        .ZN(n5661) );
  NOR2_X1 U6807 ( .A1(n5748), .A2(n5715), .ZN(n5727) );
  INV_X1 U6808 ( .A(n5654), .ZN(n5655) );
  NAND2_X1 U6809 ( .A1(n5727), .A2(n5655), .ZN(n5704) );
  NOR2_X1 U6810 ( .A1(n5699), .A2(n5656), .ZN(n5677) );
  NAND4_X1 U6811 ( .A1(n5677), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n4341), .ZN(n5657) );
  OAI211_X1 U6812 ( .C1(n5659), .C2(n6218), .A(n5658), .B(n5657), .ZN(n5660)
         );
  AOI21_X1 U6813 ( .B1(INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5661), .A(n5660), 
        .ZN(n5662) );
  OAI21_X1 U6814 ( .B1(n5663), .B2(n6206), .A(n5662), .ZN(U2987) );
  INV_X1 U6815 ( .A(n5664), .ZN(n5671) );
  INV_X1 U6816 ( .A(n5665), .ZN(n5668) );
  NAND3_X1 U6817 ( .A1(n5677), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5666), .ZN(n5667) );
  OAI211_X1 U6818 ( .C1(n5669), .C2(n6218), .A(n5668), .B(n5667), .ZN(n5670)
         );
  AOI21_X1 U6819 ( .B1(n5671), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5670), 
        .ZN(n5672) );
  OAI21_X1 U6820 ( .B1(n5673), .B2(n6206), .A(n5672), .ZN(U2988) );
  NOR2_X1 U6821 ( .A1(n5674), .A2(n6218), .ZN(n5675) );
  AOI211_X1 U6822 ( .C1(n5677), .C2(n5527), .A(n5676), .B(n5675), .ZN(n5680)
         );
  NAND2_X1 U6823 ( .A1(n5678), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5679) );
  OAI211_X1 U6824 ( .C1(n5681), .C2(n6206), .A(n5680), .B(n5679), .ZN(U2989)
         );
  INV_X1 U6825 ( .A(n5682), .ZN(n5687) );
  NOR3_X1 U6826 ( .A1(n5699), .A2(n5684), .A3(n5683), .ZN(n5685) );
  AOI211_X1 U6827 ( .C1(n6170), .C2(n5687), .A(n5686), .B(n5685), .ZN(n5690)
         );
  INV_X1 U6828 ( .A(n5688), .ZN(n5701) );
  NAND2_X1 U6829 ( .A1(n5701), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5689) );
  OAI211_X1 U6830 ( .C1(n5691), .C2(n6206), .A(n5690), .B(n5689), .ZN(U2990)
         );
  OR2_X1 U6831 ( .A1(n5693), .A2(n5692), .ZN(n5694) );
  NAND2_X1 U6832 ( .A1(n5695), .A2(n5694), .ZN(n5873) );
  INV_X1 U6833 ( .A(n5873), .ZN(n5697) );
  AOI21_X1 U6834 ( .B1(n5697), .B2(n6170), .A(n5696), .ZN(n5698) );
  OAI21_X1 U6835 ( .B1(n5699), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5698), 
        .ZN(n5700) );
  AOI21_X1 U6836 ( .B1(n5701), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5700), 
        .ZN(n5702) );
  OAI21_X1 U6837 ( .B1(n5703), .B2(n6206), .A(n5702), .ZN(U2991) );
  INV_X1 U6838 ( .A(n5704), .ZN(n5913) );
  NAND3_X1 U6839 ( .A1(n5913), .A2(n5706), .A3(n5705), .ZN(n5709) );
  INV_X1 U6840 ( .A(n5707), .ZN(n5708) );
  OAI211_X1 U6841 ( .C1(n6218), .C2(n5710), .A(n5709), .B(n5708), .ZN(n5711)
         );
  AOI21_X1 U6842 ( .B1(n5712), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5711), 
        .ZN(n5713) );
  OAI21_X1 U6843 ( .B1(n5714), .B2(n6206), .A(n5713), .ZN(U2992) );
  INV_X1 U6844 ( .A(n5748), .ZN(n5763) );
  INV_X1 U6845 ( .A(n5715), .ZN(n5716) );
  NAND3_X1 U6846 ( .A1(n5763), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n5716), .ZN(n5717) );
  AOI21_X1 U6847 ( .B1(n5718), .B2(n5717), .A(n5920), .ZN(n5719) );
  AOI211_X1 U6848 ( .C1(n6170), .C2(n5819), .A(n5720), .B(n5719), .ZN(n5721)
         );
  OAI21_X1 U6849 ( .B1(n5722), .B2(n6206), .A(n5721), .ZN(U2994) );
  OAI21_X1 U6850 ( .B1(n5828), .B2(n6218), .A(n5723), .ZN(n5725) );
  NOR2_X1 U6851 ( .A1(n5730), .A2(n5726), .ZN(n5724) );
  AOI211_X1 U6852 ( .C1(n5727), .C2(n5726), .A(n5725), .B(n5724), .ZN(n5728)
         );
  OAI21_X1 U6853 ( .B1(n5729), .B2(n6206), .A(n5728), .ZN(U2995) );
  INV_X1 U6854 ( .A(n5730), .ZN(n5735) );
  OAI21_X1 U6855 ( .B1(n5838), .B2(n6218), .A(n5731), .ZN(n5734) );
  INV_X1 U6856 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5742) );
  NOR2_X1 U6857 ( .A1(n5732), .A2(n5742), .ZN(n5733) );
  AOI211_X1 U6858 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5735), .A(n5734), .B(n5733), .ZN(n5736) );
  OAI21_X1 U6859 ( .B1(n5737), .B2(n6206), .A(n5736), .ZN(U2996) );
  NOR2_X1 U6860 ( .A1(n5738), .A2(n5742), .ZN(n5741) );
  OAI21_X1 U6861 ( .B1(n5851), .B2(n6218), .A(n5739), .ZN(n5740) );
  AOI211_X1 U6862 ( .C1(n5743), .C2(n5742), .A(n5741), .B(n5740), .ZN(n5744)
         );
  OAI21_X1 U6863 ( .B1(n5745), .B2(n6206), .A(n5744), .ZN(U2997) );
  INV_X1 U6864 ( .A(n5746), .ZN(n5757) );
  AOI221_X1 U6865 ( .B1(n6193), .B2(n5921), .C1(n5747), .C2(n5921), .A(n5776), 
        .ZN(n5928) );
  OAI21_X1 U6866 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5782), .A(n5928), 
        .ZN(n5764) );
  NOR2_X1 U6867 ( .A1(n5749), .A2(n5748), .ZN(n5750) );
  NAND2_X1 U6868 ( .A1(n5751), .A2(n5750), .ZN(n5752) );
  OAI211_X1 U6869 ( .C1(n5754), .C2(n6218), .A(n5753), .B(n5752), .ZN(n5755)
         );
  AOI21_X1 U6870 ( .B1(n5764), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5755), 
        .ZN(n5756) );
  OAI21_X1 U6871 ( .B1(n5757), .B2(n6206), .A(n5756), .ZN(U2998) );
  XNOR2_X1 U6872 ( .A(n5618), .B(n3959), .ZN(n5759) );
  XNOR2_X1 U6873 ( .A(n5760), .B(n5759), .ZN(n5906) );
  INV_X1 U6874 ( .A(n5906), .ZN(n5767) );
  INV_X1 U6875 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5761) );
  OAI22_X1 U6876 ( .A1(n5872), .A2(n6218), .B1(n6190), .B2(n5761), .ZN(n5762)
         );
  AOI21_X1 U6877 ( .B1(n5763), .B2(n3959), .A(n5762), .ZN(n5766) );
  NAND2_X1 U6878 ( .A1(n5764), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5765) );
  OAI211_X1 U6879 ( .C1(n5767), .C2(n6206), .A(n5766), .B(n5765), .ZN(U2999)
         );
  INV_X1 U6880 ( .A(n5923), .ZN(n5779) );
  OAI21_X1 U6881 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5618), .A(n5604), 
        .ZN(n5768) );
  OAI21_X1 U6882 ( .B1(n5769), .B2(n5921), .A(n5768), .ZN(n5771) );
  NAND2_X1 U6883 ( .A1(n5771), .A2(n5770), .ZN(n5773) );
  NAND2_X1 U6884 ( .A1(n5773), .A2(n5772), .ZN(n5910) );
  NAND2_X1 U6885 ( .A1(n5910), .A2(n6223), .ZN(n5778) );
  INV_X1 U6886 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5774) );
  OAI22_X1 U6887 ( .A1(n5983), .A2(n6218), .B1(n6190), .B2(n5774), .ZN(n5775)
         );
  AOI21_X1 U6888 ( .B1(n5776), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5775), 
        .ZN(n5777) );
  OAI211_X1 U6889 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5779), .A(n5778), .B(n5777), .ZN(U3001) );
  NOR3_X1 U6890 ( .A1(n6152), .A2(n5940), .A3(n5945), .ZN(n5795) );
  AOI22_X1 U6891 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .B1(n5780), .B2(n5794), .ZN(n5786)
         );
  OAI211_X1 U6892 ( .C1(n5782), .C2(n5781), .A(n5935), .B(n5933), .ZN(n5789)
         );
  NAND2_X1 U6893 ( .A1(n5789), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5784) );
  OAI211_X1 U6894 ( .C1(n6218), .C2(n5996), .A(n5784), .B(n5783), .ZN(n5785)
         );
  AOI21_X1 U6895 ( .B1(n5795), .B2(n5786), .A(n5785), .ZN(n5787) );
  OAI21_X1 U6896 ( .B1(n5788), .B2(n6206), .A(n5787), .ZN(U3002) );
  NAND2_X1 U6897 ( .A1(n5789), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5791) );
  OAI211_X1 U6898 ( .C1(n6218), .C2(n5792), .A(n5791), .B(n5790), .ZN(n5793)
         );
  AOI21_X1 U6899 ( .B1(n5795), .B2(n5794), .A(n5793), .ZN(n5796) );
  OAI21_X1 U6900 ( .B1(n5797), .B2(n6206), .A(n5796), .ZN(U3003) );
  OAI211_X1 U6901 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4482), .A(n5800), .B(
        n6568), .ZN(n5798) );
  OAI21_X1 U6902 ( .B1(n4342), .B2(n5802), .A(n5798), .ZN(n5799) );
  MUX2_X1 U6903 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5799), .S(n6570), 
        .Z(U3464) );
  XNOR2_X1 U6904 ( .A(n5801), .B(n5800), .ZN(n5803) );
  OAI22_X1 U6905 ( .A1(n5803), .A2(n6587), .B1(n4408), .B2(n5802), .ZN(n5804)
         );
  MUX2_X1 U6906 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5804), .S(n6570), 
        .Z(U3463) );
  OAI22_X1 U6907 ( .A1(n5807), .A2(n5806), .B1(n6467), .B2(n5805), .ZN(n5809)
         );
  MUX2_X1 U6908 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5809), .S(n5808), 
        .Z(U3456) );
  AND2_X1 U6909 ( .A1(n6119), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U6910 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6728) );
  AOI22_X1 U6911 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6050), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6062), .ZN(n5810) );
  OAI21_X1 U6912 ( .B1(n5811), .B2(n6047), .A(n5810), .ZN(n5812) );
  AOI221_X1 U6913 ( .B1(n5814), .B2(REIP_REG_27__SCAN_IN), .C1(n5813), .C2(
        n6728), .A(n5812), .ZN(n5817) );
  NOR2_X1 U6914 ( .A1(n5873), .A2(n6061), .ZN(n5815) );
  AOI21_X1 U6915 ( .B1(n5879), .B2(n6033), .A(n5815), .ZN(n5816) );
  NAND2_X1 U6916 ( .A1(n5817), .A2(n5816), .ZN(U2800) );
  AOI22_X1 U6917 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n6062), .B1(n5818), 
        .B2(n6071), .ZN(n5824) );
  AOI22_X1 U6918 ( .A1(EBX_REG_24__SCAN_IN), .A2(n6050), .B1(
        REIP_REG_24__SCAN_IN), .B2(n5830), .ZN(n5823) );
  AOI22_X1 U6919 ( .A1(n5884), .A2(n6033), .B1(n6066), .B2(n5819), .ZN(n5822)
         );
  INV_X1 U6920 ( .A(n5820), .ZN(n5821) );
  NAND4_X1 U6921 ( .A1(n5824), .A2(n5823), .A3(n5822), .A4(n5821), .ZN(U2803)
         );
  INV_X1 U6922 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5826) );
  OAI22_X1 U6923 ( .A1(n5826), .A2(n6039), .B1(n5825), .B2(n6047), .ZN(n5827)
         );
  AOI21_X1 U6924 ( .B1(EBX_REG_23__SCAN_IN), .B2(n6050), .A(n5827), .ZN(n5834)
         );
  NOR2_X1 U6925 ( .A1(n5828), .A2(n6061), .ZN(n5829) );
  AOI21_X1 U6926 ( .B1(n5887), .B2(n6033), .A(n5829), .ZN(n5833) );
  OAI21_X1 U6927 ( .B1(REIP_REG_23__SCAN_IN), .B2(n5831), .A(n5830), .ZN(n5832) );
  NAND3_X1 U6928 ( .A1(n5834), .A2(n5833), .A3(n5832), .ZN(U2804) );
  INV_X1 U6929 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U6930 ( .A1(n5835), .A2(n5864), .ZN(n5854) );
  AOI22_X1 U6931 ( .A1(EBX_REG_22__SCAN_IN), .A2(n6050), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6062), .ZN(n5844) );
  INV_X1 U6932 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6660) );
  INV_X1 U6933 ( .A(n5836), .ZN(n5837) );
  AOI211_X1 U6934 ( .C1(n6539), .C2(n6660), .A(n5837), .B(n5847), .ZN(n5841)
         );
  OAI22_X1 U6935 ( .A1(n5839), .A2(n5856), .B1(n5838), .B2(n6061), .ZN(n5840)
         );
  AOI211_X1 U6936 ( .C1(n6071), .C2(n5842), .A(n5841), .B(n5840), .ZN(n5843)
         );
  OAI211_X1 U6937 ( .C1(n6539), .C2(n5854), .A(n5844), .B(n5843), .ZN(U2805)
         );
  AOI22_X1 U6938 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6050), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6062), .ZN(n5845) );
  OAI21_X1 U6939 ( .B1(n6660), .B2(n5854), .A(n5845), .ZN(n5849) );
  OAI22_X1 U6940 ( .A1(n5847), .A2(REIP_REG_21__SCAN_IN), .B1(n5846), .B2(
        n6047), .ZN(n5848) );
  AOI211_X1 U6941 ( .C1(n5890), .C2(n6033), .A(n5849), .B(n5848), .ZN(n5850)
         );
  OAI21_X1 U6942 ( .B1(n5851), .B2(n6061), .A(n5850), .ZN(U2806) );
  AOI22_X1 U6943 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6050), .B1(n5852), .B2(n6071), .ZN(n5860) );
  NOR2_X1 U6944 ( .A1(n6534), .A2(n5853), .ZN(n5865) );
  AOI21_X1 U6945 ( .B1(REIP_REG_19__SCAN_IN), .B2(n5865), .A(
        REIP_REG_20__SCAN_IN), .ZN(n5855) );
  OAI22_X1 U6946 ( .A1(n5893), .A2(n5856), .B1(n5855), .B2(n5854), .ZN(n5857)
         );
  AOI21_X1 U6947 ( .B1(n6066), .B2(n5858), .A(n5857), .ZN(n5859) );
  OAI211_X1 U6948 ( .C1(n5861), .C2(n6039), .A(n5860), .B(n5859), .ZN(U2807)
         );
  AOI21_X1 U6949 ( .B1(n5864), .B2(n5863), .A(n5862), .ZN(n5869) );
  AOI22_X1 U6950 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n6062), .B1(n5865), 
        .B2(n5761), .ZN(n5868) );
  OAI21_X1 U6951 ( .B1(n6047), .B2(n5909), .A(n6190), .ZN(n5866) );
  AOI21_X1 U6952 ( .B1(n6050), .B2(EBX_REG_19__SCAN_IN), .A(n5866), .ZN(n5867)
         );
  OAI211_X1 U6953 ( .C1(n5869), .C2(n5761), .A(n5868), .B(n5867), .ZN(n5870)
         );
  AOI21_X1 U6954 ( .B1(n5905), .B2(n6033), .A(n5870), .ZN(n5871) );
  OAI21_X1 U6955 ( .B1(n6061), .B2(n5872), .A(n5871), .ZN(U2808) );
  NOR2_X1 U6956 ( .A1(n5873), .A2(n5503), .ZN(n5874) );
  AOI21_X1 U6957 ( .B1(n5879), .B2(n6082), .A(n5874), .ZN(n5875) );
  OAI21_X1 U6958 ( .B1(n6086), .B2(n5876), .A(n5875), .ZN(U2832) );
  AOI22_X1 U6959 ( .A1(n2988), .A2(n6091), .B1(n6090), .B2(DATAI_29_), .ZN(
        n5878) );
  AOI22_X1 U6960 ( .A1(n6094), .A2(DATAI_13_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6093), .ZN(n5877) );
  NAND2_X1 U6961 ( .A1(n5878), .A2(n5877), .ZN(U2862) );
  AOI22_X1 U6962 ( .A1(n5879), .A2(n6091), .B1(n6090), .B2(DATAI_27_), .ZN(
        n5881) );
  AOI22_X1 U6963 ( .A1(n6094), .A2(DATAI_11_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6093), .ZN(n5880) );
  NAND2_X1 U6964 ( .A1(n5881), .A2(n5880), .ZN(U2864) );
  AOI22_X1 U6965 ( .A1(n5901), .A2(n6091), .B1(n6090), .B2(DATAI_25_), .ZN(
        n5883) );
  AOI22_X1 U6966 ( .A1(n6094), .A2(DATAI_9_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6093), .ZN(n5882) );
  NAND2_X1 U6967 ( .A1(n5883), .A2(n5882), .ZN(U2866) );
  AOI22_X1 U6968 ( .A1(n5884), .A2(n6091), .B1(n6090), .B2(DATAI_24_), .ZN(
        n5886) );
  AOI22_X1 U6969 ( .A1(n6094), .A2(DATAI_8_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6093), .ZN(n5885) );
  NAND2_X1 U6970 ( .A1(n5886), .A2(n5885), .ZN(U2867) );
  AOI22_X1 U6971 ( .A1(n5887), .A2(n6091), .B1(n6090), .B2(DATAI_23_), .ZN(
        n5889) );
  AOI22_X1 U6972 ( .A1(n6094), .A2(DATAI_7_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6093), .ZN(n5888) );
  NAND2_X1 U6973 ( .A1(n5889), .A2(n5888), .ZN(U2868) );
  AOI22_X1 U6974 ( .A1(n5890), .A2(n6091), .B1(n6090), .B2(DATAI_21_), .ZN(
        n5892) );
  AOI22_X1 U6975 ( .A1(n6094), .A2(DATAI_5_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n6093), .ZN(n5891) );
  NAND2_X1 U6976 ( .A1(n5892), .A2(n5891), .ZN(U2870) );
  INV_X1 U6977 ( .A(n5893), .ZN(n5894) );
  AOI22_X1 U6978 ( .A1(n5894), .A2(n6091), .B1(n6090), .B2(DATAI_20_), .ZN(
        n5896) );
  AOI22_X1 U6979 ( .A1(n6094), .A2(DATAI_4_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n6093), .ZN(n5895) );
  NAND2_X1 U6980 ( .A1(n5896), .A2(n5895), .ZN(U2871) );
  AOI22_X1 U6981 ( .A1(n5905), .A2(n6091), .B1(n6090), .B2(DATAI_19_), .ZN(
        n5898) );
  AOI22_X1 U6982 ( .A1(n6094), .A2(DATAI_3_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6093), .ZN(n5897) );
  NAND2_X1 U6983 ( .A1(n5898), .A2(n5897), .ZN(U2872) );
  AOI22_X1 U6984 ( .A1(n6133), .A2(REIP_REG_25__SCAN_IN), .B1(n6148), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5903) );
  OAI21_X1 U6985 ( .B1(n5900), .B2(n5899), .A(n3020), .ZN(n5916) );
  AOI22_X1 U6986 ( .A1(n5901), .A2(n6138), .B1(n6137), .B2(n5916), .ZN(n5902)
         );
  OAI211_X1 U6987 ( .C1(n6143), .C2(n5904), .A(n5903), .B(n5902), .ZN(U2961)
         );
  AOI22_X1 U6988 ( .A1(n6133), .A2(REIP_REG_19__SCAN_IN), .B1(n6148), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5908) );
  AOI22_X1 U6989 ( .A1(n5906), .A2(n6137), .B1(n6138), .B2(n5905), .ZN(n5907)
         );
  OAI211_X1 U6990 ( .C1(n6143), .C2(n5909), .A(n5908), .B(n5907), .ZN(U2967)
         );
  AOI22_X1 U6991 ( .A1(n6133), .A2(REIP_REG_17__SCAN_IN), .B1(n6148), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5912) );
  AOI22_X1 U6992 ( .A1(n5910), .A2(n6137), .B1(n6138), .B2(n6087), .ZN(n5911)
         );
  OAI211_X1 U6993 ( .C1(n6143), .C2(n5987), .A(n5912), .B(n5911), .ZN(U2969)
         );
  AOI22_X1 U6994 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6133), .B1(n5913), .B2(
        n5919), .ZN(n5918) );
  INV_X1 U6995 ( .A(n5914), .ZN(n5915) );
  AOI22_X1 U6996 ( .A1(n5916), .A2(n6223), .B1(n6170), .B2(n5915), .ZN(n5917)
         );
  OAI211_X1 U6997 ( .C1(n5920), .C2(n5919), .A(n5918), .B(n5917), .ZN(U2993)
         );
  NOR2_X1 U6998 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5921), .ZN(n5922)
         );
  AOI22_X1 U6999 ( .A1(n6133), .A2(REIP_REG_18__SCAN_IN), .B1(n5923), .B2(
        n5922), .ZN(n5927) );
  AOI22_X1 U7000 ( .A1(n5925), .A2(n6223), .B1(n6170), .B2(n5924), .ZN(n5926)
         );
  OAI211_X1 U7001 ( .C1(n5928), .C2(n5608), .A(n5927), .B(n5926), .ZN(U3000)
         );
  INV_X1 U7002 ( .A(n5930), .ZN(n5937) );
  NAND2_X1 U7003 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5931) );
  NOR2_X1 U7004 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5931), .ZN(n5947)
         );
  INV_X1 U7005 ( .A(n6225), .ZN(n5932) );
  NAND2_X1 U7006 ( .A1(n5930), .A2(n5929), .ZN(n6203) );
  AOI22_X1 U7007 ( .A1(n5932), .A2(n5940), .B1(n5931), .B2(n6203), .ZN(n5934)
         );
  NAND3_X1 U7008 ( .A1(n5935), .A2(n5934), .A3(n5933), .ZN(n5950) );
  AOI221_X1 U7009 ( .B1(n5937), .B2(n5947), .C1(n5936), .C2(n5947), .A(n5950), 
        .ZN(n5946) );
  AOI21_X1 U7010 ( .B1(n5939), .B2(n6170), .A(n5938), .ZN(n5944) );
  NOR2_X1 U7011 ( .A1(n6152), .A2(n5940), .ZN(n5941) );
  AOI22_X1 U7012 ( .A1(n5942), .A2(n6223), .B1(n5941), .B2(n5945), .ZN(n5943)
         );
  OAI211_X1 U7013 ( .C1(n5946), .C2(n5945), .A(n5944), .B(n5943), .ZN(U3004)
         );
  INV_X1 U7014 ( .A(n5947), .ZN(n5954) );
  AOI21_X1 U7015 ( .B1(n6170), .B2(n5949), .A(n5948), .ZN(n5953) );
  AOI22_X1 U7016 ( .A1(n5951), .A2(n6223), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5950), .ZN(n5952) );
  OAI211_X1 U7017 ( .C1(n6152), .C2(n5954), .A(n5953), .B(n5952), .ZN(U3005)
         );
  INV_X1 U7018 ( .A(STATE_REG_1__SCAN_IN), .ZN(n5955) );
  NOR2_X2 U7019 ( .A1(STATE_REG_0__SCAN_IN), .A2(n5955), .ZN(n6786) );
  INV_X1 U7020 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6625) );
  AOI221_X1 U7021 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_0__SCAN_IN), .C1(
        n5955), .C2(STATE_REG_0__SCAN_IN), .A(n6786), .ZN(n6558) );
  OAI21_X1 U7022 ( .B1(n6786), .B2(n6625), .A(n6554), .ZN(U2789) );
  INV_X1 U7023 ( .A(n5956), .ZN(n6446) );
  OAI22_X1 U7024 ( .A1(n6453), .A2(n5958), .B1(n6446), .B2(n5957), .ZN(n5963)
         );
  OAI21_X1 U7025 ( .B1(n5963), .B2(n6477), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5959) );
  OAI21_X1 U7026 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6478), .A(n5959), .ZN(
        U2790) );
  INV_X1 U7027 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6742) );
  NOR2_X1 U7028 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5961) );
  NOR2_X1 U7029 ( .A1(n6786), .A2(n5961), .ZN(n5960) );
  AOI22_X1 U7030 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n6786), .B1(n6742), .B2(
        n5960), .ZN(U2791) );
  OAI21_X1 U7031 ( .B1(BS16_N), .B2(n5961), .A(n6558), .ZN(n6556) );
  OAI21_X1 U7032 ( .B1(n6558), .B2(n6730), .A(n6556), .ZN(U2792) );
  AOI21_X1 U7033 ( .B1(n5962), .B2(n6496), .A(READY_N), .ZN(n6591) );
  NOR2_X1 U7034 ( .A1(n5963), .A2(n6591), .ZN(n6455) );
  NOR2_X1 U7035 ( .A1(n6455), .A2(n6477), .ZN(n6585) );
  OAI21_X1 U7036 ( .B1(n6585), .B2(n6755), .A(n6145), .ZN(U2793) );
  NOR4_X1 U7037 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5967) );
  NOR4_X1 U7038 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n5966) );
  NOR4_X1 U7039 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5965) );
  NOR4_X1 U7040 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5964) );
  NAND4_X1 U7041 ( .A1(n5967), .A2(n5966), .A3(n5965), .A4(n5964), .ZN(n5973)
         );
  NOR4_X1 U7042 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n5971) );
  AOI211_X1 U7043 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_2__SCAN_IN), .B(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n5970) );
  NOR4_X1 U7044 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n5969) );
  NOR4_X1 U7045 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n5968) );
  NAND4_X1 U7046 ( .A1(n5971), .A2(n5970), .A3(n5969), .A4(n5968), .ZN(n5972)
         );
  NOR2_X1 U7047 ( .A1(n5973), .A2(n5972), .ZN(n6581) );
  INV_X1 U7048 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5975) );
  NOR3_X1 U7049 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5976) );
  OAI21_X1 U7050 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5976), .A(n6581), .ZN(n5974)
         );
  OAI21_X1 U7051 ( .B1(n6581), .B2(n5975), .A(n5974), .ZN(U2794) );
  INV_X1 U7052 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6557) );
  AOI21_X1 U7053 ( .B1(n6574), .B2(n6557), .A(n5976), .ZN(n5977) );
  INV_X1 U7054 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6622) );
  INV_X1 U7055 ( .A(n6581), .ZN(n6576) );
  AOI22_X1 U7056 ( .A1(n6581), .A2(n5977), .B1(n6622), .B2(n6576), .ZN(U2795)
         );
  NOR2_X1 U7057 ( .A1(n6069), .A2(n5978), .ZN(n5988) );
  AOI21_X1 U7058 ( .B1(REIP_REG_16__SCAN_IN), .B2(n5988), .A(
        REIP_REG_17__SCAN_IN), .ZN(n5981) );
  INV_X1 U7059 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5979) );
  OAI22_X1 U7060 ( .A1(n5981), .A2(n5980), .B1(n5979), .B2(n6039), .ZN(n5982)
         );
  AOI211_X1 U7061 ( .C1(n6050), .C2(EBX_REG_17__SCAN_IN), .A(n6133), .B(n5982), 
        .ZN(n5986) );
  INV_X1 U7062 ( .A(n5983), .ZN(n5984) );
  AOI22_X1 U7063 ( .A1(n6087), .A2(n6033), .B1(n6066), .B2(n5984), .ZN(n5985)
         );
  OAI211_X1 U7064 ( .C1(n5987), .C2(n6047), .A(n5986), .B(n5985), .ZN(U2810)
         );
  INV_X1 U7065 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6531) );
  AOI22_X1 U7066 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6050), .B1(n5988), .B2(n6531), .ZN(n5989) );
  OAI21_X1 U7067 ( .B1(n6531), .B2(n5990), .A(n5989), .ZN(n5991) );
  AOI211_X1 U7068 ( .C1(n6062), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6133), 
        .B(n5991), .ZN(n5995) );
  INV_X1 U7069 ( .A(n5992), .ZN(n5993) );
  AOI22_X1 U7070 ( .A1(n6092), .A2(n6033), .B1(n5993), .B2(n6071), .ZN(n5994)
         );
  OAI211_X1 U7071 ( .C1(n6061), .C2(n5996), .A(n5995), .B(n5994), .ZN(U2811)
         );
  OAI22_X1 U7072 ( .A1(n5998), .A2(n6078), .B1(n6061), .B2(n5997), .ZN(n5999)
         );
  AOI211_X1 U7073 ( .C1(n6062), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6133), 
        .B(n5999), .ZN(n6007) );
  AOI22_X1 U7074 ( .A1(n6001), .A2(n6033), .B1(n6071), .B2(n6000), .ZN(n6006)
         );
  OAI21_X1 U7075 ( .B1(n6009), .B2(n6002), .A(REIP_REG_10__SCAN_IN), .ZN(n6005) );
  NAND3_X1 U7076 ( .A1(n6054), .A2(n6521), .A3(n6003), .ZN(n6004) );
  NAND4_X1 U7077 ( .A1(n6007), .A2(n6006), .A3(n6005), .A4(n6004), .ZN(U2817)
         );
  INV_X1 U7078 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6516) );
  INV_X1 U7079 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6514) );
  NOR2_X1 U7080 ( .A1(n6516), .A2(n6514), .ZN(n6020) );
  NOR2_X1 U7081 ( .A1(n6069), .A2(n6008), .ZN(n6043) );
  AND2_X1 U7082 ( .A1(n6043), .A2(REIP_REG_5__SCAN_IN), .ZN(n6031) );
  AOI21_X1 U7083 ( .B1(n6020), .B2(n6031), .A(REIP_REG_8__SCAN_IN), .ZN(n6018)
         );
  INV_X1 U7084 ( .A(n6009), .ZN(n6017) );
  OAI22_X1 U7085 ( .A1(n6011), .A2(n6078), .B1(n6061), .B2(n6010), .ZN(n6012)
         );
  AOI211_X1 U7086 ( .C1(n6062), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6133), 
        .B(n6012), .ZN(n6016) );
  AOI22_X1 U7087 ( .A1(n6014), .A2(n6033), .B1(n6071), .B2(n6013), .ZN(n6015)
         );
  OAI211_X1 U7088 ( .C1(n6018), .C2(n6017), .A(n6016), .B(n6015), .ZN(U2819)
         );
  OAI21_X1 U7089 ( .B1(n6069), .B2(n6019), .A(n6068), .ZN(n6042) );
  AOI21_X1 U7090 ( .B1(n6516), .B2(n6514), .A(n6020), .ZN(n6021) );
  AOI22_X1 U7091 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6042), .B1(n6031), .B2(n6021), .ZN(n6027) );
  AOI22_X1 U7092 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6050), .B1(n6066), .B2(n6169), 
        .ZN(n6022) );
  OAI211_X1 U7093 ( .C1(n6039), .C2(n6023), .A(n6190), .B(n6022), .ZN(n6024)
         );
  AOI21_X1 U7094 ( .B1(n6025), .B2(n6033), .A(n6024), .ZN(n6026) );
  OAI211_X1 U7095 ( .C1(n6028), .C2(n6047), .A(n6027), .B(n6026), .ZN(U2820)
         );
  AOI22_X1 U7096 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6062), .B1(n6066), 
        .B2(n6080), .ZN(n6029) );
  OAI211_X1 U7097 ( .C1(n6078), .C2(n6085), .A(n6029), .B(n6190), .ZN(n6030)
         );
  AOI221_X1 U7098 ( .B1(n6042), .B2(REIP_REG_6__SCAN_IN), .C1(n6031), .C2(
        n6514), .A(n6030), .ZN(n6035) );
  AOI22_X1 U7099 ( .A1(n6083), .A2(n6033), .B1(n6071), .B2(n6032), .ZN(n6034)
         );
  NAND2_X1 U7100 ( .A1(n6035), .A2(n6034), .ZN(U2821) );
  AOI22_X1 U7101 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6050), .B1(n6066), .B2(n6036), 
        .ZN(n6037) );
  OAI211_X1 U7102 ( .C1(n6039), .C2(n6038), .A(n6190), .B(n6037), .ZN(n6040)
         );
  AOI21_X1 U7103 ( .B1(n6041), .B2(n6067), .A(n6040), .ZN(n6045) );
  OAI21_X1 U7104 ( .B1(REIP_REG_5__SCAN_IN), .B2(n6043), .A(n6042), .ZN(n6044)
         );
  OAI211_X1 U7105 ( .C1(n6047), .C2(n6046), .A(n6045), .B(n6044), .ZN(U2822)
         );
  AOI22_X1 U7106 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6049), .B1(n6048), .B2(n6064), .ZN(n6059) );
  AOI22_X1 U7107 ( .A1(EBX_REG_4__SCAN_IN), .A2(n6050), .B1(
        PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6062), .ZN(n6057) );
  AOI22_X1 U7108 ( .A1(n6052), .A2(n6067), .B1(n6051), .B2(n6071), .ZN(n6056)
         );
  INV_X1 U7109 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6510) );
  NAND3_X1 U7110 ( .A1(n6054), .A2(n6053), .A3(n6510), .ZN(n6055) );
  AND4_X1 U7111 ( .A1(n6057), .A2(n6056), .A3(n6190), .A4(n6055), .ZN(n6058)
         );
  OAI211_X1 U7112 ( .C1(n6061), .C2(n6060), .A(n6059), .B(n6058), .ZN(U2823)
         );
  AOI222_X1 U7113 ( .A1(n6066), .A2(n6065), .B1(n6064), .B2(n6063), .C1(
        PHYADDRPOINTER_REG_2__SCAN_IN), .C2(n6062), .ZN(n6077) );
  NAND2_X1 U7114 ( .A1(n6139), .A2(n6067), .ZN(n6075) );
  OAI211_X1 U7115 ( .C1(n6069), .C2(REIP_REG_1__SCAN_IN), .A(n6068), .B(
        REIP_REG_2__SCAN_IN), .ZN(n6073) );
  OAI21_X1 U7116 ( .B1(n6069), .B2(n6574), .A(n6506), .ZN(n6072) );
  INV_X1 U7117 ( .A(n6142), .ZN(n6070) );
  AOI22_X1 U7118 ( .A1(n6073), .A2(n6072), .B1(n6071), .B2(n6070), .ZN(n6074)
         );
  AND2_X1 U7119 ( .A1(n6075), .A2(n6074), .ZN(n6076) );
  OAI211_X1 U7120 ( .C1(n6079), .C2(n6078), .A(n6077), .B(n6076), .ZN(U2825)
         );
  AOI22_X1 U7121 ( .A1(n6083), .A2(n6082), .B1(n6081), .B2(n6080), .ZN(n6084)
         );
  OAI21_X1 U7122 ( .B1(n6086), .B2(n6085), .A(n6084), .ZN(U2853) );
  AOI22_X1 U7123 ( .A1(n6087), .A2(n6091), .B1(n6090), .B2(DATAI_17_), .ZN(
        n6089) );
  AOI22_X1 U7124 ( .A1(n6094), .A2(DATAI_1_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n6093), .ZN(n6088) );
  NAND2_X1 U7125 ( .A1(n6089), .A2(n6088), .ZN(U2874) );
  AOI22_X1 U7126 ( .A1(n6092), .A2(n6091), .B1(n6090), .B2(DATAI_16_), .ZN(
        n6096) );
  AOI22_X1 U7127 ( .A1(n6094), .A2(DATAI_0_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n6093), .ZN(n6095) );
  NAND2_X1 U7128 ( .A1(n6096), .A2(n6095), .ZN(U2875) );
  AOI22_X1 U7129 ( .A1(n6129), .A2(LWORD_REG_15__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6098) );
  OAI21_X1 U7130 ( .B1(n4446), .B2(n6131), .A(n6098), .ZN(U2908) );
  INV_X1 U7131 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6100) );
  AOI22_X1 U7132 ( .A1(n6129), .A2(LWORD_REG_14__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6099) );
  OAI21_X1 U7133 ( .B1(n6100), .B2(n6131), .A(n6099), .ZN(U2909) );
  AOI22_X1 U7134 ( .A1(n6129), .A2(LWORD_REG_13__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6101) );
  OAI21_X1 U7135 ( .B1(n6102), .B2(n6131), .A(n6101), .ZN(U2910) );
  AOI22_X1 U7136 ( .A1(n6129), .A2(LWORD_REG_12__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6103) );
  OAI21_X1 U7137 ( .B1(n6104), .B2(n6131), .A(n6103), .ZN(U2911) );
  AOI22_X1 U7138 ( .A1(n6129), .A2(LWORD_REG_11__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6105) );
  OAI21_X1 U7139 ( .B1(n6106), .B2(n6131), .A(n6105), .ZN(U2912) );
  AOI22_X1 U7140 ( .A1(n6129), .A2(LWORD_REG_10__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6107) );
  OAI21_X1 U7141 ( .B1(n6108), .B2(n6131), .A(n6107), .ZN(U2913) );
  AOI22_X1 U7142 ( .A1(n6129), .A2(LWORD_REG_9__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6109) );
  OAI21_X1 U7143 ( .B1(n6110), .B2(n6131), .A(n6109), .ZN(U2914) );
  AOI22_X1 U7144 ( .A1(n6129), .A2(LWORD_REG_8__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6111) );
  OAI21_X1 U7145 ( .B1(n6112), .B2(n6131), .A(n6111), .ZN(U2915) );
  AOI22_X1 U7146 ( .A1(n6129), .A2(LWORD_REG_7__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6113) );
  OAI21_X1 U7147 ( .B1(n6114), .B2(n6131), .A(n6113), .ZN(U2916) );
  AOI22_X1 U7148 ( .A1(n6129), .A2(LWORD_REG_6__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6115) );
  OAI21_X1 U7149 ( .B1(n6116), .B2(n6131), .A(n6115), .ZN(U2917) );
  AOI22_X1 U7150 ( .A1(n6129), .A2(LWORD_REG_5__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6117) );
  OAI21_X1 U7151 ( .B1(n6118), .B2(n6131), .A(n6117), .ZN(U2918) );
  AOI22_X1 U7152 ( .A1(n6129), .A2(LWORD_REG_4__SCAN_IN), .B1(n6119), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6120) );
  OAI21_X1 U7153 ( .B1(n6121), .B2(n6131), .A(n6120), .ZN(U2919) );
  AOI22_X1 U7154 ( .A1(n6129), .A2(LWORD_REG_3__SCAN_IN), .B1(n6128), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6122) );
  OAI21_X1 U7155 ( .B1(n6123), .B2(n6131), .A(n6122), .ZN(U2920) );
  AOI22_X1 U7156 ( .A1(n6129), .A2(LWORD_REG_2__SCAN_IN), .B1(n6128), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6124) );
  OAI21_X1 U7157 ( .B1(n6125), .B2(n6131), .A(n6124), .ZN(U2921) );
  AOI22_X1 U7158 ( .A1(n6129), .A2(LWORD_REG_1__SCAN_IN), .B1(n6128), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6126) );
  OAI21_X1 U7159 ( .B1(n6127), .B2(n6131), .A(n6126), .ZN(U2922) );
  AOI22_X1 U7160 ( .A1(n6129), .A2(LWORD_REG_0__SCAN_IN), .B1(n6128), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6130) );
  OAI21_X1 U7161 ( .B1(n6132), .B2(n6131), .A(n6130), .ZN(U2923) );
  AOI22_X1 U7162 ( .A1(n6133), .A2(REIP_REG_2__SCAN_IN), .B1(n6148), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6141) );
  XNOR2_X1 U7163 ( .A(n6134), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6135)
         );
  XNOR2_X1 U7164 ( .A(n6136), .B(n6135), .ZN(n6196) );
  AOI22_X1 U7165 ( .A1(n6139), .A2(n6138), .B1(n6137), .B2(n6196), .ZN(n6140)
         );
  OAI211_X1 U7166 ( .C1(n6143), .C2(n6142), .A(n6141), .B(n6140), .ZN(U2984)
         );
  OAI21_X1 U7167 ( .B1(n6144), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4029), 
        .ZN(n6215) );
  NAND2_X1 U7168 ( .A1(n6133), .A2(REIP_REG_0__SCAN_IN), .ZN(n6216) );
  OAI21_X1 U7169 ( .B1(n6215), .B2(n6145), .A(n6216), .ZN(n6146) );
  INV_X1 U7170 ( .A(n6146), .ZN(n6150) );
  OAI21_X1 U7171 ( .B1(n6148), .B2(n6147), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6149) );
  OAI211_X1 U7172 ( .C1(n6151), .C2(n6371), .A(n6150), .B(n6149), .ZN(U2986)
         );
  AND2_X1 U7173 ( .A1(n6153), .A2(n6152), .ZN(n6158) );
  AOI22_X1 U7174 ( .A1(n6155), .A2(n6223), .B1(n6170), .B2(n6154), .ZN(n6157)
         );
  NAND2_X1 U7175 ( .A1(n6133), .A2(REIP_REG_11__SCAN_IN), .ZN(n6156) );
  OAI211_X1 U7176 ( .C1(n6159), .C2(n6158), .A(n6157), .B(n6156), .ZN(U3007)
         );
  INV_X1 U7177 ( .A(n6160), .ZN(n6168) );
  AOI21_X1 U7178 ( .B1(n6170), .B2(n6162), .A(n6161), .ZN(n6166) );
  AOI22_X1 U7179 ( .A1(n6164), .A2(n6223), .B1(n6163), .B2(n6167), .ZN(n6165)
         );
  OAI211_X1 U7180 ( .C1(n6168), .C2(n6167), .A(n6166), .B(n6165), .ZN(U3009)
         );
  NAND2_X1 U7181 ( .A1(n6170), .A2(n6169), .ZN(n6172) );
  OAI211_X1 U7182 ( .C1(n6173), .C2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6172), 
        .B(n6171), .ZN(n6174) );
  AOI21_X1 U7183 ( .B1(n6175), .B2(n6223), .A(n6174), .ZN(n6176) );
  OAI21_X1 U7184 ( .B1(n6178), .B2(n6177), .A(n6176), .ZN(U3011) );
  OAI21_X1 U7185 ( .B1(n6218), .B2(n6180), .A(n6179), .ZN(n6181) );
  INV_X1 U7186 ( .A(n6181), .ZN(n6184) );
  OR2_X1 U7187 ( .A1(n6182), .A2(n6206), .ZN(n6183) );
  OAI211_X1 U7188 ( .C1(n6185), .C2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6184), 
        .B(n6183), .ZN(n6186) );
  INV_X1 U7189 ( .A(n6186), .ZN(n6187) );
  OAI21_X1 U7190 ( .B1(n6189), .B2(n6188), .A(n6187), .ZN(U3015) );
  OAI22_X1 U7191 ( .A1(n6218), .A2(n6191), .B1(n6190), .B2(n6506), .ZN(n6192)
         );
  INV_X1 U7192 ( .A(n6192), .ZN(n6202) );
  OAI221_X1 U7193 ( .B1(n6195), .B2(n6194), .C1(n6195), .C2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(n6193), .ZN(n6201) );
  AOI22_X1 U7194 ( .A1(n6197), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6223), 
        .B2(n6196), .ZN(n6200) );
  OR3_X1 U7195 ( .A1(n6214), .A2(n6198), .A3(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6199) );
  NAND4_X1 U7196 ( .A1(n6202), .A2(n6201), .A3(n6200), .A4(n6199), .ZN(U3016)
         );
  NAND2_X1 U7197 ( .A1(n6227), .A2(n6203), .ZN(n6219) );
  NOR2_X1 U7198 ( .A1(n6204), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6211)
         );
  NOR2_X1 U7199 ( .A1(n6206), .A2(n6205), .ZN(n6210) );
  OAI21_X1 U7200 ( .B1(n6218), .B2(n6208), .A(n6207), .ZN(n6209) );
  AOI211_X1 U7201 ( .C1(n6212), .C2(n6211), .A(n6210), .B(n6209), .ZN(n6213)
         );
  OAI221_X1 U7202 ( .B1(n6214), .B2(n6226), .C1(n6214), .C2(n6219), .A(n6213), 
        .ZN(U3017) );
  INV_X1 U7203 ( .A(n6215), .ZN(n6222) );
  OAI21_X1 U7204 ( .B1(n6218), .B2(n6217), .A(n6216), .ZN(n6221) );
  INV_X1 U7205 ( .A(n6219), .ZN(n6220) );
  AOI211_X1 U7206 ( .C1(n6223), .C2(n6222), .A(n6221), .B(n6220), .ZN(n6224)
         );
  OAI221_X1 U7207 ( .B1(n6227), .B2(n6226), .C1(n6227), .C2(n6225), .A(n6224), 
        .ZN(U3018) );
  NOR2_X1 U7208 ( .A1(n6461), .A2(n6570), .ZN(U3019) );
  NOR2_X1 U7209 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6229), .ZN(n6262)
         );
  OAI22_X1 U7210 ( .A1(n6233), .A2(n6587), .B1(n6231), .B2(n6230), .ZN(n6261)
         );
  AOI22_X1 U7211 ( .A1(n6369), .A2(n6262), .B1(n6368), .B2(n6261), .ZN(n6241)
         );
  INV_X1 U7212 ( .A(n6428), .ZN(n6232) );
  OAI21_X1 U7213 ( .B1(n6263), .B2(n6232), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6234) );
  NAND3_X1 U7214 ( .A1(n6234), .A2(n6568), .A3(n6233), .ZN(n6239) );
  INV_X1 U7215 ( .A(n6262), .ZN(n6237) );
  AOI211_X1 U7216 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6237), .A(n6236), .B(
        n6235), .ZN(n6238) );
  NAND2_X1 U7217 ( .A1(n6239), .A2(n6238), .ZN(n6264) );
  AOI22_X1 U7218 ( .A1(n6264), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n6320), 
        .B2(n6263), .ZN(n6240) );
  OAI211_X1 U7219 ( .C1(n6242), .C2(n6428), .A(n6241), .B(n6240), .ZN(U3020)
         );
  AOI22_X1 U7220 ( .A1(n6384), .A2(n6262), .B1(n6383), .B2(n6261), .ZN(n6244)
         );
  AOI22_X1 U7221 ( .A1(n6264), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n6329), 
        .B2(n6263), .ZN(n6243) );
  OAI211_X1 U7222 ( .C1(n6245), .C2(n6428), .A(n6244), .B(n6243), .ZN(U3021)
         );
  AOI22_X1 U7223 ( .A1(n6390), .A2(n6262), .B1(n6389), .B2(n6261), .ZN(n6247)
         );
  AOI22_X1 U7224 ( .A1(n6264), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n6333), 
        .B2(n6263), .ZN(n6246) );
  OAI211_X1 U7225 ( .C1(n6248), .C2(n6428), .A(n6247), .B(n6246), .ZN(U3022)
         );
  AOI22_X1 U7226 ( .A1(n6396), .A2(n6262), .B1(n6395), .B2(n6261), .ZN(n6250)
         );
  AOI22_X1 U7227 ( .A1(n6264), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n6337), 
        .B2(n6263), .ZN(n6249) );
  OAI211_X1 U7228 ( .C1(n6251), .C2(n6428), .A(n6250), .B(n6249), .ZN(U3023)
         );
  AOI22_X1 U7229 ( .A1(n6402), .A2(n6262), .B1(n6401), .B2(n6261), .ZN(n6253)
         );
  AOI22_X1 U7230 ( .A1(n6264), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n6341), 
        .B2(n6263), .ZN(n6252) );
  OAI211_X1 U7231 ( .C1(n6254), .C2(n6428), .A(n6253), .B(n6252), .ZN(U3024)
         );
  AOI22_X1 U7232 ( .A1(n6408), .A2(n6262), .B1(n6407), .B2(n6261), .ZN(n6256)
         );
  AOI22_X1 U7233 ( .A1(n6264), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n6345), 
        .B2(n6263), .ZN(n6255) );
  OAI211_X1 U7234 ( .C1(n6257), .C2(n6428), .A(n6256), .B(n6255), .ZN(U3025)
         );
  AOI22_X1 U7235 ( .A1(n6414), .A2(n6262), .B1(n6413), .B2(n6261), .ZN(n6259)
         );
  AOI22_X1 U7236 ( .A1(n6264), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n6349), 
        .B2(n6263), .ZN(n6258) );
  OAI211_X1 U7237 ( .C1(n6260), .C2(n6428), .A(n6259), .B(n6258), .ZN(U3026)
         );
  AOI22_X1 U7238 ( .A1(n6422), .A2(n6262), .B1(n6420), .B2(n6261), .ZN(n6266)
         );
  AOI22_X1 U7239 ( .A1(n6264), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n6354), 
        .B2(n6263), .ZN(n6265) );
  OAI211_X1 U7240 ( .C1(n6267), .C2(n6428), .A(n6266), .B(n6265), .ZN(U3027)
         );
  AOI22_X1 U7241 ( .A1(n6275), .A2(n6385), .B1(n6384), .B2(n6274), .ZN(n6269)
         );
  AOI22_X1 U7242 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6277), .B1(n6383), 
        .B2(n6276), .ZN(n6268) );
  OAI211_X1 U7243 ( .C1(n6388), .C2(n6280), .A(n6269), .B(n6268), .ZN(U3045)
         );
  AOI22_X1 U7244 ( .A1(n6275), .A2(n6391), .B1(n6390), .B2(n6274), .ZN(n6271)
         );
  AOI22_X1 U7245 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6277), .B1(n6389), 
        .B2(n6276), .ZN(n6270) );
  OAI211_X1 U7246 ( .C1(n6394), .C2(n6280), .A(n6271), .B(n6270), .ZN(U3046)
         );
  AOI22_X1 U7247 ( .A1(n6275), .A2(n6403), .B1(n6402), .B2(n6274), .ZN(n6273)
         );
  AOI22_X1 U7248 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6277), .B1(n6401), 
        .B2(n6276), .ZN(n6272) );
  OAI211_X1 U7249 ( .C1(n6406), .C2(n6280), .A(n6273), .B(n6272), .ZN(U3048)
         );
  AOI22_X1 U7250 ( .A1(n6275), .A2(n6415), .B1(n6414), .B2(n6274), .ZN(n6279)
         );
  AOI22_X1 U7251 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6277), .B1(n6413), 
        .B2(n6276), .ZN(n6278) );
  OAI211_X1 U7252 ( .C1(n6418), .C2(n6280), .A(n6279), .B(n6278), .ZN(U3050)
         );
  NAND2_X1 U7253 ( .A1(n6281), .A2(n6312), .ZN(n6564) );
  AND2_X1 U7254 ( .A1(n6564), .A2(n6568), .ZN(n6288) );
  INV_X1 U7255 ( .A(n6282), .ZN(n6305) );
  AOI21_X1 U7256 ( .B1(n6283), .B2(n6315), .A(n6305), .ZN(n6287) );
  INV_X1 U7257 ( .A(n6287), .ZN(n6285) );
  AOI22_X1 U7258 ( .A1(n6288), .A2(n6285), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6284), .ZN(n6310) );
  AOI22_X1 U7259 ( .A1(n6369), .A2(n6305), .B1(n6306), .B2(n6320), .ZN(n6291)
         );
  AOI22_X1 U7260 ( .A1(n6288), .A2(n6287), .B1(n6286), .B2(n6587), .ZN(n6289)
         );
  NAND2_X1 U7261 ( .A1(n6377), .A2(n6289), .ZN(n6307) );
  AOI22_X1 U7262 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6307), .B1(n6379), 
        .B2(n6304), .ZN(n6290) );
  OAI211_X1 U7263 ( .C1(n6310), .C2(n6328), .A(n6291), .B(n6290), .ZN(U3076)
         );
  AOI22_X1 U7264 ( .A1(n6384), .A2(n6305), .B1(n6306), .B2(n6329), .ZN(n6293)
         );
  AOI22_X1 U7265 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6307), .B1(n6385), 
        .B2(n6304), .ZN(n6292) );
  OAI211_X1 U7266 ( .C1(n6310), .C2(n6332), .A(n6293), .B(n6292), .ZN(U3077)
         );
  AOI22_X1 U7267 ( .A1(n6390), .A2(n6305), .B1(n6304), .B2(n6391), .ZN(n6295)
         );
  AOI22_X1 U7268 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6307), .B1(n6333), 
        .B2(n6306), .ZN(n6294) );
  OAI211_X1 U7269 ( .C1(n6310), .C2(n6336), .A(n6295), .B(n6294), .ZN(U3078)
         );
  AOI22_X1 U7270 ( .A1(n6396), .A2(n6305), .B1(n6306), .B2(n6337), .ZN(n6297)
         );
  AOI22_X1 U7271 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6307), .B1(n6397), 
        .B2(n6304), .ZN(n6296) );
  OAI211_X1 U7272 ( .C1(n6310), .C2(n6340), .A(n6297), .B(n6296), .ZN(U3079)
         );
  AOI22_X1 U7273 ( .A1(n6402), .A2(n6305), .B1(n6304), .B2(n6403), .ZN(n6299)
         );
  AOI22_X1 U7274 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6307), .B1(n6341), 
        .B2(n6306), .ZN(n6298) );
  OAI211_X1 U7275 ( .C1(n6310), .C2(n6344), .A(n6299), .B(n6298), .ZN(U3080)
         );
  AOI22_X1 U7276 ( .A1(n6408), .A2(n6305), .B1(n6304), .B2(n6409), .ZN(n6301)
         );
  AOI22_X1 U7277 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6307), .B1(n6345), 
        .B2(n6306), .ZN(n6300) );
  OAI211_X1 U7278 ( .C1(n6310), .C2(n6348), .A(n6301), .B(n6300), .ZN(U3081)
         );
  AOI22_X1 U7279 ( .A1(n6414), .A2(n6305), .B1(n6304), .B2(n6415), .ZN(n6303)
         );
  AOI22_X1 U7280 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6307), .B1(n6349), 
        .B2(n6306), .ZN(n6302) );
  OAI211_X1 U7281 ( .C1(n6310), .C2(n6352), .A(n6303), .B(n6302), .ZN(U3082)
         );
  AOI22_X1 U7282 ( .A1(n6422), .A2(n6305), .B1(n6304), .B2(n6424), .ZN(n6309)
         );
  AOI22_X1 U7283 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6307), .B1(n6354), 
        .B2(n6306), .ZN(n6308) );
  OAI211_X1 U7284 ( .C1(n6310), .C2(n6360), .A(n6309), .B(n6308), .ZN(U3083)
         );
  INV_X1 U7285 ( .A(n6311), .ZN(n6313) );
  AOI21_X1 U7286 ( .B1(n6313), .B2(n6312), .A(n6587), .ZN(n6322) );
  NOR2_X1 U7287 ( .A1(n6314), .A2(n6572), .ZN(n6353) );
  AOI21_X1 U7288 ( .B1(n6316), .B2(n6315), .A(n6353), .ZN(n6321) );
  INV_X1 U7289 ( .A(n6321), .ZN(n6318) );
  INV_X1 U7290 ( .A(n6317), .ZN(n6324) );
  AOI22_X1 U7291 ( .A1(n6322), .A2(n6318), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6324), .ZN(n6361) );
  AOI22_X1 U7292 ( .A1(n6355), .A2(n6320), .B1(n6369), .B2(n6353), .ZN(n6327)
         );
  NAND2_X1 U7293 ( .A1(n6322), .A2(n6321), .ZN(n6323) );
  OAI211_X1 U7294 ( .C1(n6568), .C2(n6324), .A(n6377), .B(n6323), .ZN(n6357)
         );
  AOI22_X1 U7295 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6357), .B1(n6379), 
        .B2(n6356), .ZN(n6326) );
  OAI211_X1 U7296 ( .C1(n6361), .C2(n6328), .A(n6327), .B(n6326), .ZN(U3108)
         );
  AOI22_X1 U7297 ( .A1(n6355), .A2(n6329), .B1(n6384), .B2(n6353), .ZN(n6331)
         );
  AOI22_X1 U7298 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6357), .B1(n6385), 
        .B2(n6356), .ZN(n6330) );
  OAI211_X1 U7299 ( .C1(n6361), .C2(n6332), .A(n6331), .B(n6330), .ZN(U3109)
         );
  AOI22_X1 U7300 ( .A1(n6355), .A2(n6333), .B1(n6390), .B2(n6353), .ZN(n6335)
         );
  AOI22_X1 U7301 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6357), .B1(n6391), 
        .B2(n6356), .ZN(n6334) );
  OAI211_X1 U7302 ( .C1(n6361), .C2(n6336), .A(n6335), .B(n6334), .ZN(U3110)
         );
  AOI22_X1 U7303 ( .A1(n6356), .A2(n6397), .B1(n6396), .B2(n6353), .ZN(n6339)
         );
  AOI22_X1 U7304 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6357), .B1(n6337), 
        .B2(n6355), .ZN(n6338) );
  OAI211_X1 U7305 ( .C1(n6361), .C2(n6340), .A(n6339), .B(n6338), .ZN(U3111)
         );
  AOI22_X1 U7306 ( .A1(n6356), .A2(n6403), .B1(n6402), .B2(n6353), .ZN(n6343)
         );
  AOI22_X1 U7307 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6357), .B1(n6341), 
        .B2(n6355), .ZN(n6342) );
  OAI211_X1 U7308 ( .C1(n6361), .C2(n6344), .A(n6343), .B(n6342), .ZN(U3112)
         );
  AOI22_X1 U7309 ( .A1(n6355), .A2(n6345), .B1(n6408), .B2(n6353), .ZN(n6347)
         );
  AOI22_X1 U7310 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6357), .B1(n6409), 
        .B2(n6356), .ZN(n6346) );
  OAI211_X1 U7311 ( .C1(n6361), .C2(n6348), .A(n6347), .B(n6346), .ZN(U3113)
         );
  AOI22_X1 U7312 ( .A1(n6355), .A2(n6349), .B1(n6414), .B2(n6353), .ZN(n6351)
         );
  AOI22_X1 U7313 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6357), .B1(n6415), 
        .B2(n6356), .ZN(n6350) );
  OAI211_X1 U7314 ( .C1(n6361), .C2(n6352), .A(n6351), .B(n6350), .ZN(U3114)
         );
  AOI22_X1 U7315 ( .A1(n6355), .A2(n6354), .B1(n6422), .B2(n6353), .ZN(n6359)
         );
  AOI22_X1 U7316 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6357), .B1(n6424), 
        .B2(n6356), .ZN(n6358) );
  OAI211_X1 U7317 ( .C1(n6361), .C2(n6360), .A(n6359), .B(n6358), .ZN(U3115)
         );
  INV_X1 U7318 ( .A(n6364), .ZN(n6421) );
  NAND2_X1 U7319 ( .A1(n6363), .A2(n6362), .ZN(n6365) );
  NAND2_X1 U7320 ( .A1(n6365), .A2(n6364), .ZN(n6373) );
  NAND2_X1 U7321 ( .A1(n6373), .A2(n6568), .ZN(n6367) );
  NAND2_X1 U7322 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6378), .ZN(n6366) );
  NAND2_X1 U7323 ( .A1(n6367), .A2(n6366), .ZN(n6419) );
  AOI22_X1 U7324 ( .A1(n6369), .A2(n6421), .B1(n6368), .B2(n6419), .ZN(n6381)
         );
  INV_X1 U7325 ( .A(n6370), .ZN(n6372) );
  AOI21_X1 U7326 ( .B1(n6372), .B2(n4482), .A(n6371), .ZN(n6375) );
  INV_X1 U7327 ( .A(n6373), .ZN(n6374) );
  OAI21_X1 U7328 ( .B1(n6375), .B2(n6566), .A(n6374), .ZN(n6376) );
  OAI211_X1 U7329 ( .C1(n6378), .C2(n6568), .A(n6377), .B(n6376), .ZN(n6425)
         );
  AOI22_X1 U7330 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6425), .B1(n6379), 
        .B2(n6423), .ZN(n6380) );
  OAI211_X1 U7331 ( .C1(n6382), .C2(n6428), .A(n6381), .B(n6380), .ZN(U3140)
         );
  AOI22_X1 U7332 ( .A1(n6384), .A2(n6421), .B1(n6383), .B2(n6419), .ZN(n6387)
         );
  AOI22_X1 U7333 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n6425), .B1(n6385), 
        .B2(n6423), .ZN(n6386) );
  OAI211_X1 U7334 ( .C1(n6388), .C2(n6428), .A(n6387), .B(n6386), .ZN(U3141)
         );
  AOI22_X1 U7335 ( .A1(n6390), .A2(n6421), .B1(n6389), .B2(n6419), .ZN(n6393)
         );
  AOI22_X1 U7336 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n6425), .B1(n6391), 
        .B2(n6423), .ZN(n6392) );
  OAI211_X1 U7337 ( .C1(n6394), .C2(n6428), .A(n6393), .B(n6392), .ZN(U3142)
         );
  AOI22_X1 U7338 ( .A1(n6396), .A2(n6421), .B1(n6395), .B2(n6419), .ZN(n6399)
         );
  AOI22_X1 U7339 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n6425), .B1(n6397), 
        .B2(n6423), .ZN(n6398) );
  OAI211_X1 U7340 ( .C1(n6400), .C2(n6428), .A(n6399), .B(n6398), .ZN(U3143)
         );
  AOI22_X1 U7341 ( .A1(n6402), .A2(n6421), .B1(n6401), .B2(n6419), .ZN(n6405)
         );
  AOI22_X1 U7342 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n6425), .B1(n6403), 
        .B2(n6423), .ZN(n6404) );
  OAI211_X1 U7343 ( .C1(n6406), .C2(n6428), .A(n6405), .B(n6404), .ZN(U3144)
         );
  AOI22_X1 U7344 ( .A1(n6408), .A2(n6421), .B1(n6407), .B2(n6419), .ZN(n6411)
         );
  AOI22_X1 U7345 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6425), .B1(n6409), 
        .B2(n6423), .ZN(n6410) );
  OAI211_X1 U7346 ( .C1(n6412), .C2(n6428), .A(n6411), .B(n6410), .ZN(U3145)
         );
  AOI22_X1 U7347 ( .A1(n6414), .A2(n6421), .B1(n6413), .B2(n6419), .ZN(n6417)
         );
  AOI22_X1 U7348 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n6425), .B1(n6415), 
        .B2(n6423), .ZN(n6416) );
  OAI211_X1 U7349 ( .C1(n6418), .C2(n6428), .A(n6417), .B(n6416), .ZN(U3146)
         );
  AOI22_X1 U7350 ( .A1(n6422), .A2(n6421), .B1(n6420), .B2(n6419), .ZN(n6427)
         );
  AOI22_X1 U7351 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6425), .B1(n6424), 
        .B2(n6423), .ZN(n6426) );
  OAI211_X1 U7352 ( .C1(n6429), .C2(n6428), .A(n6427), .B(n6426), .ZN(U3147)
         );
  NOR2_X1 U7353 ( .A1(n6431), .A2(n6430), .ZN(n6432) );
  AND2_X1 U7354 ( .A1(n6433), .A2(n6432), .ZN(n6439) );
  INV_X1 U7355 ( .A(n6439), .ZN(n6436) );
  OAI211_X1 U7356 ( .C1(n6437), .C2(n6436), .A(n6435), .B(n6434), .ZN(n6438)
         );
  OAI21_X1 U7357 ( .B1(n6439), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6438), 
        .ZN(n6440) );
  AOI222_X1 U7358 ( .A1(n6442), .A2(n6441), .B1(n6442), .B2(n6440), .C1(n6441), 
        .C2(n6440), .ZN(n6444) );
  AND2_X1 U7359 ( .A1(n6444), .A2(n6443), .ZN(n6445) );
  OAI22_X1 U7360 ( .A1(n6445), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(n6444), .B2(n6443), .ZN(n6462) );
  NOR2_X1 U7361 ( .A1(n6447), .A2(n6446), .ZN(n6451) );
  INV_X1 U7362 ( .A(n6448), .ZN(n6449) );
  OAI22_X1 U7363 ( .A1(n6453), .A2(n6451), .B1(n6450), .B2(n6449), .ZN(n6452)
         );
  AOI21_X1 U7364 ( .B1(n6454), .B2(n6453), .A(n6452), .ZN(n6584) );
  OAI21_X1 U7365 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6455), 
        .ZN(n6456) );
  NAND4_X1 U7366 ( .A1(n6458), .A2(n6584), .A3(n6457), .A4(n6456), .ZN(n6459)
         );
  AOI211_X1 U7367 ( .C1(n6462), .C2(n6461), .A(n6460), .B(n6459), .ZN(n6463)
         );
  INV_X1 U7368 ( .A(n6463), .ZN(n6469) );
  OAI22_X1 U7369 ( .A1(n6469), .A2(n6477), .B1(n6588), .B2(n6658), .ZN(n6464)
         );
  OAI21_X1 U7370 ( .B1(n6466), .B2(n6465), .A(n6464), .ZN(n6561) );
  OAI21_X1 U7371 ( .B1(n6467), .B2(n6483), .A(n6561), .ZN(n6475) );
  OAI21_X1 U7372 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6658), .A(n6561), .ZN(
        n6476) );
  AOI211_X1 U7373 ( .C1(n6470), .C2(n6469), .A(n6468), .B(n6476), .ZN(n6473)
         );
  INV_X1 U7374 ( .A(n6471), .ZN(n6472) );
  OAI221_X1 U7375 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6475), .C1(n6474), .C2(
        n6473), .A(n6472), .ZN(U3148) );
  NAND3_X1 U7376 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6484), .A3(n6476), .ZN(
        n6482) );
  OAI21_X1 U7377 ( .B1(READY_N), .B2(n6478), .A(n6477), .ZN(n6480) );
  AOI21_X1 U7378 ( .B1(n6480), .B2(n6561), .A(n6479), .ZN(n6481) );
  NAND2_X1 U7379 ( .A1(n6482), .A2(n6481), .ZN(U3149) );
  INV_X1 U7380 ( .A(n6483), .ZN(n6593) );
  OAI211_X1 U7381 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6658), .A(n6559), .B(
        n6484), .ZN(n6486) );
  OAI21_X1 U7382 ( .B1(n6593), .B2(n6486), .A(n6485), .ZN(U3150) );
  AND2_X1 U7383 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6554), .ZN(U3151) );
  AND2_X1 U7384 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6554), .ZN(U3152) );
  AND2_X1 U7385 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6554), .ZN(U3153) );
  AND2_X1 U7386 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6554), .ZN(U3154) );
  AND2_X1 U7387 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6554), .ZN(U3155) );
  AND2_X1 U7388 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6554), .ZN(U3156) );
  AND2_X1 U7389 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6554), .ZN(U3157) );
  AND2_X1 U7390 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6554), .ZN(U3158) );
  AND2_X1 U7391 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6554), .ZN(U3159) );
  AND2_X1 U7392 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6554), .ZN(U3160) );
  AND2_X1 U7393 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6554), .ZN(U3161) );
  AND2_X1 U7394 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6554), .ZN(U3162) );
  AND2_X1 U7395 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6554), .ZN(U3163) );
  AND2_X1 U7396 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6554), .ZN(U3164) );
  AND2_X1 U7397 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6554), .ZN(U3165) );
  AND2_X1 U7398 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6554), .ZN(U3166) );
  AND2_X1 U7399 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6554), .ZN(U3167) );
  AND2_X1 U7400 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6554), .ZN(U3168) );
  AND2_X1 U7401 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6554), .ZN(U3169) );
  AND2_X1 U7402 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6554), .ZN(U3170) );
  AND2_X1 U7403 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6554), .ZN(U3171) );
  AND2_X1 U7404 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6554), .ZN(U3172) );
  AND2_X1 U7405 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6554), .ZN(U3173) );
  AND2_X1 U7406 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6554), .ZN(U3174) );
  AND2_X1 U7407 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6554), .ZN(U3175) );
  AND2_X1 U7408 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6554), .ZN(U3176) );
  AND2_X1 U7409 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6554), .ZN(U3177) );
  AND2_X1 U7410 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6554), .ZN(U3178) );
  AND2_X1 U7411 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6554), .ZN(U3179) );
  AND2_X1 U7412 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6554), .ZN(U3180) );
  NAND2_X1 U7413 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6491) );
  NAND2_X1 U7414 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6492) );
  NAND2_X1 U7415 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6498) );
  NAND2_X1 U7416 ( .A1(n6492), .A2(n6498), .ZN(n6488) );
  INV_X1 U7417 ( .A(NA_N), .ZN(n6724) );
  INV_X1 U7418 ( .A(n6489), .ZN(n6487) );
  AOI211_X1 U7419 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6724), .A(
        STATE_REG_0__SCAN_IN), .B(n6487), .ZN(n6503) );
  AOI21_X1 U7420 ( .B1(n6489), .B2(n6488), .A(n6503), .ZN(n6490) );
  OAI221_X1 U7421 ( .B1(n6786), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n6786), 
        .C2(n6491), .A(n6490), .ZN(U3181) );
  INV_X1 U7422 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6499) );
  INV_X1 U7423 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6752) );
  NOR2_X1 U7424 ( .A1(n6499), .A2(n6752), .ZN(n6494) );
  INV_X1 U7425 ( .A(n6491), .ZN(n6493) );
  OAI21_X1 U7426 ( .B1(n6494), .B2(n6493), .A(n6492), .ZN(n6495) );
  NAND3_X1 U7427 ( .A1(n6496), .A2(n6498), .A3(n6495), .ZN(U3182) );
  AOI221_X1 U7428 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6658), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6497) );
  AOI221_X1 U7429 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6497), .C2(HOLD), .A(n6499), .ZN(n6502) );
  OR4_X1 U7430 ( .A1(n6752), .A2(n6499), .A3(n6498), .A4(NA_N), .ZN(n6501) );
  NAND3_X1 U7431 ( .A1(READY_N), .A2(STATE_REG_2__SCAN_IN), .A3(
        STATE_REG_1__SCAN_IN), .ZN(n6500) );
  OAI211_X1 U7432 ( .C1(n6503), .C2(n6502), .A(n6501), .B(n6500), .ZN(U3183)
         );
  NAND2_X1 U7433 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6786), .ZN(n6552) );
  NOR2_X2 U7434 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6598), .ZN(n6550) );
  AOI22_X1 U7435 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6598), .ZN(n6504) );
  OAI21_X1 U7436 ( .B1(n6574), .B2(n6552), .A(n6504), .ZN(U3184) );
  AOI22_X1 U7437 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6598), .ZN(n6505) );
  OAI21_X1 U7438 ( .B1(n6506), .B2(n6552), .A(n6505), .ZN(U3185) );
  AOI22_X1 U7439 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6598), .ZN(n6507) );
  OAI21_X1 U7440 ( .B1(n6508), .B2(n6552), .A(n6507), .ZN(U3186) );
  AOI22_X1 U7441 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6598), .ZN(n6509) );
  OAI21_X1 U7442 ( .B1(n6510), .B2(n6552), .A(n6509), .ZN(U3187) );
  AOI22_X1 U7443 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6598), .ZN(n6511) );
  OAI21_X1 U7444 ( .B1(n6512), .B2(n6552), .A(n6511), .ZN(U3188) );
  AOI22_X1 U7445 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6598), .ZN(n6513) );
  OAI21_X1 U7446 ( .B1(n6514), .B2(n6552), .A(n6513), .ZN(U3189) );
  AOI22_X1 U7447 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6598), .ZN(n6515) );
  OAI21_X1 U7448 ( .B1(n6516), .B2(n6552), .A(n6515), .ZN(U3190) );
  INV_X1 U7449 ( .A(n6552), .ZN(n6547) );
  AOI22_X1 U7450 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6598), .ZN(n6517) );
  OAI21_X1 U7451 ( .B1(n6518), .B2(n6549), .A(n6517), .ZN(U3191) );
  AOI22_X1 U7452 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6598), .ZN(n6519) );
  OAI21_X1 U7453 ( .B1(n6521), .B2(n6549), .A(n6519), .ZN(U3192) );
  AOI22_X1 U7454 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6598), .ZN(n6520) );
  OAI21_X1 U7455 ( .B1(n6521), .B2(n6552), .A(n6520), .ZN(U3193) );
  AOI22_X1 U7456 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6598), .ZN(n6522) );
  OAI21_X1 U7457 ( .B1(n6524), .B2(n6549), .A(n6522), .ZN(U3194) );
  AOI22_X1 U7458 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6598), .ZN(n6523) );
  OAI21_X1 U7459 ( .B1(n6524), .B2(n6552), .A(n6523), .ZN(U3195) );
  AOI22_X1 U7460 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6598), .ZN(n6525) );
  OAI21_X1 U7461 ( .B1(n6526), .B2(n6552), .A(n6525), .ZN(U3196) );
  AOI22_X1 U7462 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6598), .ZN(n6527) );
  OAI21_X1 U7463 ( .B1(n6528), .B2(n6549), .A(n6527), .ZN(U3197) );
  AOI22_X1 U7464 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6598), .ZN(n6529) );
  OAI21_X1 U7465 ( .B1(n6531), .B2(n6549), .A(n6529), .ZN(U3198) );
  AOI22_X1 U7466 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6598), .ZN(n6530) );
  OAI21_X1 U7467 ( .B1(n6531), .B2(n6552), .A(n6530), .ZN(U3199) );
  AOI22_X1 U7468 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6598), .ZN(n6532) );
  OAI21_X1 U7469 ( .B1(n6534), .B2(n6549), .A(n6532), .ZN(U3200) );
  AOI22_X1 U7470 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6598), .ZN(n6533) );
  OAI21_X1 U7471 ( .B1(n6534), .B2(n6552), .A(n6533), .ZN(U3201) );
  AOI22_X1 U7472 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6598), .ZN(n6535) );
  OAI21_X1 U7473 ( .B1(n5761), .B2(n6552), .A(n6535), .ZN(U3202) );
  AOI22_X1 U7474 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6598), .ZN(n6536) );
  OAI21_X1 U7475 ( .B1(n6660), .B2(n6549), .A(n6536), .ZN(U3203) );
  AOI22_X1 U7476 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6598), .ZN(n6537) );
  OAI21_X1 U7477 ( .B1(n6539), .B2(n6549), .A(n6537), .ZN(U3204) );
  AOI22_X1 U7478 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6598), .ZN(n6538) );
  OAI21_X1 U7479 ( .B1(n6539), .B2(n6552), .A(n6538), .ZN(U3205) );
  AOI22_X1 U7480 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6598), .ZN(n6540) );
  OAI21_X1 U7481 ( .B1(n6657), .B2(n6552), .A(n6540), .ZN(U3206) );
  AOI22_X1 U7482 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6598), .ZN(n6541) );
  OAI21_X1 U7483 ( .B1(n6542), .B2(n6549), .A(n6541), .ZN(U3207) );
  AOI22_X1 U7484 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6598), .ZN(n6543) );
  OAI21_X1 U7485 ( .B1(n6623), .B2(n6549), .A(n6543), .ZN(U3208) );
  AOI22_X1 U7486 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6598), .ZN(n6544) );
  OAI21_X1 U7487 ( .B1(n6623), .B2(n6552), .A(n6544), .ZN(U3209) );
  AOI22_X1 U7488 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6598), .ZN(n6545) );
  OAI21_X1 U7489 ( .B1(n6662), .B2(n6549), .A(n6545), .ZN(U3210) );
  AOI22_X1 U7490 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6598), .ZN(n6546) );
  OAI21_X1 U7491 ( .B1(n6741), .B2(n6549), .A(n6546), .ZN(U3211) );
  INV_X1 U7492 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6767) );
  AOI22_X1 U7493 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6547), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6598), .ZN(n6548) );
  OAI21_X1 U7494 ( .B1(n6767), .B2(n6549), .A(n6548), .ZN(U3212) );
  AOI22_X1 U7495 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6598), .ZN(n6551) );
  OAI21_X1 U7496 ( .B1(n6767), .B2(n6552), .A(n6551), .ZN(U3213) );
  MUX2_X1 U7497 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6786), .Z(U3446) );
  MUX2_X1 U7498 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6786), .Z(U3447) );
  MUX2_X1 U7499 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6786), .Z(U3448) );
  INV_X1 U7500 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6555) );
  INV_X1 U7501 ( .A(n6556), .ZN(n6553) );
  AOI21_X1 U7502 ( .B1(n6555), .B2(n6554), .A(n6553), .ZN(U3451) );
  OAI21_X1 U7503 ( .B1(n6558), .B2(n6557), .A(n6556), .ZN(U3452) );
  OAI211_X1 U7504 ( .C1(n6562), .C2(n6561), .A(n6560), .B(n6559), .ZN(U3453)
         );
  INV_X1 U7505 ( .A(n6570), .ZN(n6573) );
  INV_X1 U7506 ( .A(n6563), .ZN(n6565) );
  NAND2_X1 U7507 ( .A1(n6565), .A2(n6564), .ZN(n6569) );
  AOI222_X1 U7508 ( .A1(n6569), .A2(n6568), .B1(n3017), .B2(n6567), .C1(n4042), 
        .C2(n6566), .ZN(n6571) );
  AOI22_X1 U7509 ( .A1(n6573), .A2(n6572), .B1(n6571), .B2(n6570), .ZN(U3462)
         );
  AOI21_X1 U7510 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6575) );
  AOI22_X1 U7511 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6575), .B2(n6574), .ZN(n6578) );
  INV_X1 U7512 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6577) );
  AOI22_X1 U7513 ( .A1(n6581), .A2(n6578), .B1(n6577), .B2(n6576), .ZN(U3468)
         );
  INV_X1 U7514 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6580) );
  OAI21_X1 U7515 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6581), .ZN(n6579) );
  OAI21_X1 U7516 ( .B1(n6581), .B2(n6580), .A(n6579), .ZN(U3469) );
  INV_X1 U7517 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6725) );
  AOI22_X1 U7518 ( .A1(n6786), .A2(READREQUEST_REG_SCAN_IN), .B1(n6725), .B2(
        n6598), .ZN(U3470) );
  INV_X1 U7519 ( .A(MORE_REG_SCAN_IN), .ZN(n6583) );
  INV_X1 U7520 ( .A(n6585), .ZN(n6582) );
  AOI22_X1 U7521 ( .A1(n6585), .A2(n6584), .B1(n6583), .B2(n6582), .ZN(U3471)
         );
  OAI211_X1 U7522 ( .C1(READY_N), .C2(n6588), .A(n6587), .B(n6586), .ZN(n6589)
         );
  NOR2_X1 U7523 ( .A1(n6590), .A2(n6589), .ZN(n6597) );
  OAI211_X1 U7524 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6592), .A(n6591), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6594) );
  AOI21_X1 U7525 ( .B1(n6594), .B2(STATE2_REG_0__SCAN_IN), .A(n6593), .ZN(
        n6596) );
  NAND2_X1 U7526 ( .A1(n6597), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6595) );
  OAI21_X1 U7527 ( .B1(n6597), .B2(n6596), .A(n6595), .ZN(U3472) );
  INV_X1 U7528 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6722) );
  INV_X1 U7529 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6758) );
  AOI22_X1 U7530 ( .A1(n6786), .A2(n6722), .B1(n6758), .B2(n6598), .ZN(U3473)
         );
  OAI22_X1 U7531 ( .A1(REIP_REG_25__SCAN_IN), .A2(keyinput_f57), .B1(DATAI_11_), .B2(keyinput_f20), .ZN(n6599) );
  AOI221_X1 U7532 ( .B1(REIP_REG_25__SCAN_IN), .B2(keyinput_f57), .C1(
        keyinput_f20), .C2(DATAI_11_), .A(n6599), .ZN(n6639) );
  OAI22_X1 U7533 ( .A1(REIP_REG_29__SCAN_IN), .A2(keyinput_f53), .B1(DATAI_29_), .B2(keyinput_f2), .ZN(n6600) );
  AOI221_X1 U7534 ( .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_f53), .C1(
        keyinput_f2), .C2(DATAI_29_), .A(n6600), .ZN(n6638) );
  AOI22_X1 U7535 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(keyinput_f39), .B1(
        DATAI_22_), .B2(keyinput_f9), .ZN(n6601) );
  OAI221_X1 U7536 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_f39), .C1(
        DATAI_22_), .C2(keyinput_f9), .A(n6601), .ZN(n6608) );
  AOI22_X1 U7537 ( .A1(keyinput_f34), .A2(BS16_N), .B1(REIP_REG_27__SCAN_IN), 
        .B2(keyinput_f55), .ZN(n6602) );
  OAI221_X1 U7538 ( .B1(keyinput_f34), .B2(BS16_N), .C1(REIP_REG_27__SCAN_IN), 
        .C2(keyinput_f55), .A(n6602), .ZN(n6607) );
  AOI22_X1 U7539 ( .A1(DATAI_9_), .A2(keyinput_f22), .B1(REIP_REG_20__SCAN_IN), 
        .B2(keyinput_f62), .ZN(n6603) );
  OAI221_X1 U7540 ( .B1(DATAI_9_), .B2(keyinput_f22), .C1(REIP_REG_20__SCAN_IN), .C2(keyinput_f62), .A(n6603), .ZN(n6606) );
  AOI22_X1 U7541 ( .A1(DATAI_19_), .A2(keyinput_f12), .B1(DATAI_14_), .B2(
        keyinput_f17), .ZN(n6604) );
  OAI221_X1 U7542 ( .B1(DATAI_19_), .B2(keyinput_f12), .C1(DATAI_14_), .C2(
        keyinput_f17), .A(n6604), .ZN(n6605) );
  NOR4_X1 U7543 ( .A1(n6608), .A2(n6607), .A3(n6606), .A4(n6605), .ZN(n6611)
         );
  OAI22_X1 U7544 ( .A1(DATAI_16_), .A2(keyinput_f15), .B1(D_C_N_REG_SCAN_IN), 
        .B2(keyinput_f41), .ZN(n6609) );
  AOI221_X1 U7545 ( .B1(DATAI_16_), .B2(keyinput_f15), .C1(keyinput_f41), .C2(
        D_C_N_REG_SCAN_IN), .A(n6609), .ZN(n6610) );
  OAI211_X1 U7546 ( .C1(n6748), .C2(keyinput_f8), .A(n6611), .B(n6610), .ZN(
        n6612) );
  AOI21_X1 U7547 ( .B1(n6748), .B2(keyinput_f8), .A(n6612), .ZN(n6637) );
  XOR2_X1 U7548 ( .A(keyinput_f48), .B(BYTEENABLE_REG_1__SCAN_IN), .Z(n6615)
         );
  AOI22_X1 U7549 ( .A1(n6767), .A2(keyinput_f52), .B1(keyinput_f7), .B2(n4579), 
        .ZN(n6613) );
  OAI221_X1 U7550 ( .B1(n6767), .B2(keyinput_f52), .C1(n4579), .C2(keyinput_f7), .A(n6613), .ZN(n6614) );
  AOI211_X1 U7551 ( .C1(n6617), .C2(keyinput_f24), .A(n6615), .B(n6614), .ZN(
        n6616) );
  OAI21_X1 U7552 ( .B1(n6617), .B2(keyinput_f24), .A(n6616), .ZN(n6635) );
  AOI22_X1 U7553 ( .A1(n6619), .A2(keyinput_f23), .B1(n4663), .B2(keyinput_f0), 
        .ZN(n6618) );
  OAI221_X1 U7554 ( .B1(n6619), .B2(keyinput_f23), .C1(n4663), .C2(keyinput_f0), .A(n6618), .ZN(n6634) );
  AOI22_X1 U7555 ( .A1(n4490), .A2(keyinput_f5), .B1(n4610), .B2(keyinput_f1), 
        .ZN(n6620) );
  OAI221_X1 U7556 ( .B1(n4490), .B2(keyinput_f5), .C1(n4610), .C2(keyinput_f1), 
        .A(n6620), .ZN(n6633) );
  OAI22_X1 U7557 ( .A1(n6623), .A2(keyinput_f56), .B1(n6622), .B2(keyinput_f50), .ZN(n6621) );
  AOI221_X1 U7558 ( .B1(n6623), .B2(keyinput_f56), .C1(keyinput_f50), .C2(
        n6622), .A(n6621), .ZN(n6631) );
  OAI22_X1 U7559 ( .A1(n5761), .A2(keyinput_f63), .B1(n6625), .B2(keyinput_f38), .ZN(n6624) );
  AOI221_X1 U7560 ( .B1(n5761), .B2(keyinput_f63), .C1(keyinput_f38), .C2(
        n6625), .A(n6624), .ZN(n6630) );
  OAI22_X1 U7561 ( .A1(n6758), .A2(keyinput_f40), .B1(n6725), .B2(keyinput_f46), .ZN(n6626) );
  AOI221_X1 U7562 ( .B1(n6758), .B2(keyinput_f40), .C1(keyinput_f46), .C2(
        n6725), .A(n6626), .ZN(n6629) );
  OAI22_X1 U7563 ( .A1(n6757), .A2(keyinput_f18), .B1(n6755), .B2(keyinput_f45), .ZN(n6627) );
  AOI221_X1 U7564 ( .B1(n6757), .B2(keyinput_f18), .C1(keyinput_f45), .C2(
        n6755), .A(n6627), .ZN(n6628) );
  NAND4_X1 U7565 ( .A1(n6631), .A2(n6630), .A3(n6629), .A4(n6628), .ZN(n6632)
         );
  NOR4_X1 U7566 ( .A1(n6635), .A2(n6634), .A3(n6633), .A4(n6632), .ZN(n6636)
         );
  NAND4_X1 U7567 ( .A1(n6639), .A2(n6638), .A3(n6637), .A4(n6636), .ZN(n6684)
         );
  AOI22_X1 U7568 ( .A1(keyinput_f36), .A2(HOLD), .B1(DATAI_6_), .B2(
        keyinput_f25), .ZN(n6640) );
  OAI221_X1 U7569 ( .B1(keyinput_f36), .B2(HOLD), .C1(DATAI_6_), .C2(
        keyinput_f25), .A(n6640), .ZN(n6647) );
  AOI22_X1 U7570 ( .A1(STATEBS16_REG_SCAN_IN), .A2(keyinput_f43), .B1(
        REIP_REG_24__SCAN_IN), .B2(keyinput_f58), .ZN(n6641) );
  OAI221_X1 U7571 ( .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput_f43), .C1(
        REIP_REG_24__SCAN_IN), .C2(keyinput_f58), .A(n6641), .ZN(n6646) );
  AOI22_X1 U7572 ( .A1(DATAI_15_), .A2(keyinput_f16), .B1(DATAI_12_), .B2(
        keyinput_f19), .ZN(n6642) );
  OAI221_X1 U7573 ( .B1(DATAI_15_), .B2(keyinput_f16), .C1(DATAI_12_), .C2(
        keyinput_f19), .A(n6642), .ZN(n6645) );
  AOI22_X1 U7574 ( .A1(DATAI_18_), .A2(keyinput_f13), .B1(DATAI_27_), .B2(
        keyinput_f4), .ZN(n6643) );
  OAI221_X1 U7575 ( .B1(DATAI_18_), .B2(keyinput_f13), .C1(DATAI_27_), .C2(
        keyinput_f4), .A(n6643), .ZN(n6644) );
  NOR4_X1 U7576 ( .A1(n6647), .A2(n6646), .A3(n6645), .A4(n6644), .ZN(n6682)
         );
  AOI22_X1 U7577 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_f32), .B1(
        DATAI_4_), .B2(keyinput_f27), .ZN(n6648) );
  OAI221_X1 U7578 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_f32), .C1(
        DATAI_4_), .C2(keyinput_f27), .A(n6648), .ZN(n6655) );
  AOI22_X1 U7579 ( .A1(DATAI_17_), .A2(keyinput_f14), .B1(DATAI_3_), .B2(
        keyinput_f28), .ZN(n6649) );
  OAI221_X1 U7580 ( .B1(DATAI_17_), .B2(keyinput_f14), .C1(DATAI_3_), .C2(
        keyinput_f28), .A(n6649), .ZN(n6654) );
  AOI22_X1 U7581 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput_f60), .B1(
        REIP_REG_31__SCAN_IN), .B2(keyinput_f51), .ZN(n6650) );
  OAI221_X1 U7582 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_f60), .C1(
        REIP_REG_31__SCAN_IN), .C2(keyinput_f51), .A(n6650), .ZN(n6653) );
  AOI22_X1 U7583 ( .A1(keyinput_f47), .A2(BYTEENABLE_REG_0__SCAN_IN), .B1(
        keyinput_f49), .B2(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6651) );
  OAI221_X1 U7584 ( .B1(keyinput_f47), .B2(BYTEENABLE_REG_0__SCAN_IN), .C1(
        keyinput_f49), .C2(BYTEENABLE_REG_2__SCAN_IN), .A(n6651), .ZN(n6652)
         );
  NOR4_X1 U7585 ( .A1(n6655), .A2(n6654), .A3(n6653), .A4(n6652), .ZN(n6681)
         );
  AOI22_X1 U7586 ( .A1(n6658), .A2(keyinput_f35), .B1(keyinput_f59), .B2(n6657), .ZN(n6656) );
  OAI221_X1 U7587 ( .B1(n6658), .B2(keyinput_f35), .C1(n6657), .C2(
        keyinput_f59), .A(n6656), .ZN(n6669) );
  AOI22_X1 U7588 ( .A1(n6660), .A2(keyinput_f61), .B1(keyinput_f6), .B2(n4616), 
        .ZN(n6659) );
  OAI221_X1 U7589 ( .B1(n6660), .B2(keyinput_f61), .C1(n4616), .C2(keyinput_f6), .A(n6659), .ZN(n6668) );
  INV_X1 U7590 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6663) );
  AOI22_X1 U7591 ( .A1(n6663), .A2(keyinput_f37), .B1(n6662), .B2(keyinput_f54), .ZN(n6661) );
  OAI221_X1 U7592 ( .B1(n6663), .B2(keyinput_f37), .C1(n6662), .C2(
        keyinput_f54), .A(n6661), .ZN(n6667) );
  AOI22_X1 U7593 ( .A1(n6665), .A2(keyinput_f10), .B1(n4621), .B2(keyinput_f3), 
        .ZN(n6664) );
  OAI221_X1 U7594 ( .B1(n6665), .B2(keyinput_f10), .C1(n4621), .C2(keyinput_f3), .A(n6664), .ZN(n6666) );
  NOR4_X1 U7595 ( .A1(n6669), .A2(n6668), .A3(n6667), .A4(n6666), .ZN(n6680)
         );
  AOI22_X1 U7596 ( .A1(keyinput_f33), .A2(NA_N), .B1(DATAI_20_), .B2(
        keyinput_f11), .ZN(n6670) );
  OAI221_X1 U7597 ( .B1(keyinput_f33), .B2(NA_N), .C1(DATAI_20_), .C2(
        keyinput_f11), .A(n6670), .ZN(n6678) );
  AOI22_X1 U7598 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_f42), .B1(
        MORE_REG_SCAN_IN), .B2(keyinput_f44), .ZN(n6671) );
  OAI221_X1 U7599 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_f42), .C1(
        MORE_REG_SCAN_IN), .C2(keyinput_f44), .A(n6671), .ZN(n6677) );
  AOI22_X1 U7600 ( .A1(n6673), .A2(keyinput_f21), .B1(keyinput_f26), .B2(n6770), .ZN(n6672) );
  OAI221_X1 U7601 ( .B1(n6673), .B2(keyinput_f21), .C1(n6770), .C2(
        keyinput_f26), .A(n6672), .ZN(n6676) );
  AOI22_X1 U7602 ( .A1(DATAI_2_), .A2(keyinput_f29), .B1(n6749), .B2(
        keyinput_f31), .ZN(n6674) );
  OAI221_X1 U7603 ( .B1(DATAI_2_), .B2(keyinput_f29), .C1(n6749), .C2(
        keyinput_f31), .A(n6674), .ZN(n6675) );
  NOR4_X1 U7604 ( .A1(n6678), .A2(n6677), .A3(n6676), .A4(n6675), .ZN(n6679)
         );
  NAND4_X1 U7605 ( .A1(n6682), .A2(n6681), .A3(n6680), .A4(n6679), .ZN(n6683)
         );
  OAI22_X1 U7606 ( .A1(n6684), .A2(n6683), .B1(keyinput_f30), .B2(DATAI_1_), 
        .ZN(n6685) );
  AOI21_X1 U7607 ( .B1(keyinput_f30), .B2(DATAI_1_), .A(n6685), .ZN(n6785) );
  AOI22_X1 U7608 ( .A1(ADS_N_REG_SCAN_IN), .A2(keyinput_g38), .B1(
        REIP_REG_25__SCAN_IN), .B2(keyinput_g57), .ZN(n6686) );
  OAI221_X1 U7609 ( .B1(ADS_N_REG_SCAN_IN), .B2(keyinput_g38), .C1(
        REIP_REG_25__SCAN_IN), .C2(keyinput_g57), .A(n6686), .ZN(n6693) );
  AOI22_X1 U7610 ( .A1(DATAI_3_), .A2(keyinput_g28), .B1(DATAI_9_), .B2(
        keyinput_g22), .ZN(n6687) );
  OAI221_X1 U7611 ( .B1(DATAI_3_), .B2(keyinput_g28), .C1(DATAI_9_), .C2(
        keyinput_g22), .A(n6687), .ZN(n6692) );
  AOI22_X1 U7612 ( .A1(DATAI_2_), .A2(keyinput_g29), .B1(DATAI_21_), .B2(
        keyinput_g10), .ZN(n6688) );
  OAI221_X1 U7613 ( .B1(DATAI_2_), .B2(keyinput_g29), .C1(DATAI_21_), .C2(
        keyinput_g10), .A(n6688), .ZN(n6691) );
  AOI22_X1 U7614 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_g50), .B1(
        BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_g49), .ZN(n6689) );
  OAI221_X1 U7615 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_g50), .C1(
        BYTEENABLE_REG_2__SCAN_IN), .C2(keyinput_g49), .A(n6689), .ZN(n6690)
         );
  NOR4_X1 U7616 ( .A1(n6693), .A2(n6692), .A3(n6691), .A4(n6690), .ZN(n6720)
         );
  XOR2_X1 U7617 ( .A(HOLD), .B(keyinput_g36), .Z(n6700) );
  AOI22_X1 U7618 ( .A1(DATAI_24_), .A2(keyinput_g7), .B1(READY_N), .B2(
        keyinput_g35), .ZN(n6694) );
  OAI221_X1 U7619 ( .B1(DATAI_24_), .B2(keyinput_g7), .C1(READY_N), .C2(
        keyinput_g35), .A(n6694), .ZN(n6699) );
  AOI22_X1 U7620 ( .A1(DATAI_6_), .A2(keyinput_g25), .B1(DATAI_25_), .B2(
        keyinput_g6), .ZN(n6695) );
  OAI221_X1 U7621 ( .B1(DATAI_6_), .B2(keyinput_g25), .C1(DATAI_25_), .C2(
        keyinput_g6), .A(n6695), .ZN(n6698) );
  AOI22_X1 U7622 ( .A1(DATAI_8_), .A2(keyinput_g23), .B1(REIP_REG_21__SCAN_IN), 
        .B2(keyinput_g61), .ZN(n6696) );
  OAI221_X1 U7623 ( .B1(DATAI_8_), .B2(keyinput_g23), .C1(REIP_REG_21__SCAN_IN), .C2(keyinput_g61), .A(n6696), .ZN(n6697) );
  NOR4_X1 U7624 ( .A1(n6700), .A2(n6699), .A3(n6698), .A4(n6697), .ZN(n6719)
         );
  AOI22_X1 U7625 ( .A1(READREQUEST_REG_SCAN_IN), .A2(keyinput_g37), .B1(
        REIP_REG_22__SCAN_IN), .B2(keyinput_g60), .ZN(n6701) );
  OAI221_X1 U7626 ( .B1(READREQUEST_REG_SCAN_IN), .B2(keyinput_g37), .C1(
        REIP_REG_22__SCAN_IN), .C2(keyinput_g60), .A(n6701), .ZN(n6708) );
  AOI22_X1 U7627 ( .A1(BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_g47), .B1(
        REIP_REG_28__SCAN_IN), .B2(keyinput_g54), .ZN(n6702) );
  OAI221_X1 U7628 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_g47), .C1(
        REIP_REG_28__SCAN_IN), .C2(keyinput_g54), .A(n6702), .ZN(n6707) );
  AOI22_X1 U7629 ( .A1(DATAI_10_), .A2(keyinput_g21), .B1(REIP_REG_26__SCAN_IN), .B2(keyinput_g56), .ZN(n6703) );
  OAI221_X1 U7630 ( .B1(DATAI_10_), .B2(keyinput_g21), .C1(
        REIP_REG_26__SCAN_IN), .C2(keyinput_g56), .A(n6703), .ZN(n6706) );
  AOI22_X1 U7631 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(keyinput_g39), .B1(
        REIP_REG_19__SCAN_IN), .B2(keyinput_g63), .ZN(n6704) );
  OAI221_X1 U7632 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_g39), .C1(
        REIP_REG_19__SCAN_IN), .C2(keyinput_g63), .A(n6704), .ZN(n6705) );
  NOR4_X1 U7633 ( .A1(n6708), .A2(n6707), .A3(n6706), .A4(n6705), .ZN(n6718)
         );
  AOI22_X1 U7634 ( .A1(DATAI_26_), .A2(keyinput_g5), .B1(REIP_REG_23__SCAN_IN), 
        .B2(keyinput_g59), .ZN(n6709) );
  OAI221_X1 U7635 ( .B1(DATAI_26_), .B2(keyinput_g5), .C1(REIP_REG_23__SCAN_IN), .C2(keyinput_g59), .A(n6709), .ZN(n6716) );
  AOI22_X1 U7636 ( .A1(BS16_N), .A2(keyinput_g34), .B1(REIP_REG_20__SCAN_IN), 
        .B2(keyinput_g62), .ZN(n6710) );
  OAI221_X1 U7637 ( .B1(BS16_N), .B2(keyinput_g34), .C1(REIP_REG_20__SCAN_IN), 
        .C2(keyinput_g62), .A(n6710), .ZN(n6715) );
  AOI22_X1 U7638 ( .A1(MORE_REG_SCAN_IN), .A2(keyinput_g44), .B1(DATAI_30_), 
        .B2(keyinput_g1), .ZN(n6711) );
  OAI221_X1 U7639 ( .B1(MORE_REG_SCAN_IN), .B2(keyinput_g44), .C1(DATAI_30_), 
        .C2(keyinput_g1), .A(n6711), .ZN(n6714) );
  AOI22_X1 U7640 ( .A1(BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_g48), .B1(
        DATAI_28_), .B2(keyinput_g3), .ZN(n6712) );
  OAI221_X1 U7641 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_g48), .C1(
        DATAI_28_), .C2(keyinput_g3), .A(n6712), .ZN(n6713) );
  NOR4_X1 U7642 ( .A1(n6716), .A2(n6715), .A3(n6714), .A4(n6713), .ZN(n6717)
         );
  NAND4_X1 U7643 ( .A1(n6720), .A2(n6719), .A3(n6718), .A4(n6717), .ZN(n6783)
         );
  AOI22_X1 U7644 ( .A1(n4669), .A2(keyinput_g2), .B1(keyinput_g32), .B2(n6722), 
        .ZN(n6721) );
  OAI221_X1 U7645 ( .B1(n4669), .B2(keyinput_g2), .C1(n6722), .C2(keyinput_g32), .A(n6721), .ZN(n6735) );
  AOI22_X1 U7646 ( .A1(n6725), .A2(keyinput_g46), .B1(n6724), .B2(keyinput_g33), .ZN(n6723) );
  OAI221_X1 U7647 ( .B1(n6725), .B2(keyinput_g46), .C1(n6724), .C2(
        keyinput_g33), .A(n6723), .ZN(n6734) );
  AOI22_X1 U7648 ( .A1(n6728), .A2(keyinput_g55), .B1(keyinput_g11), .B2(n6727), .ZN(n6726) );
  OAI221_X1 U7649 ( .B1(n6728), .B2(keyinput_g55), .C1(n6727), .C2(
        keyinput_g11), .A(n6726), .ZN(n6733) );
  AOI22_X1 U7650 ( .A1(n6731), .A2(keyinput_g19), .B1(n6730), .B2(keyinput_g43), .ZN(n6729) );
  OAI221_X1 U7651 ( .B1(n6731), .B2(keyinput_g19), .C1(n6730), .C2(
        keyinput_g43), .A(n6729), .ZN(n6732) );
  NOR4_X1 U7652 ( .A1(n6735), .A2(n6734), .A3(n6733), .A4(n6732), .ZN(n6781)
         );
  AOI22_X1 U7653 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput_g51), .B1(
        REIP_REG_24__SCAN_IN), .B2(keyinput_g58), .ZN(n6736) );
  OAI221_X1 U7654 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_g51), .C1(
        REIP_REG_24__SCAN_IN), .C2(keyinput_g58), .A(n6736), .ZN(n6746) );
  AOI22_X1 U7655 ( .A1(DATAI_7_), .A2(keyinput_g24), .B1(DATAI_11_), .B2(
        keyinput_g20), .ZN(n6737) );
  OAI221_X1 U7656 ( .B1(DATAI_7_), .B2(keyinput_g24), .C1(DATAI_11_), .C2(
        keyinput_g20), .A(n6737), .ZN(n6745) );
  AOI22_X1 U7657 ( .A1(n6739), .A2(keyinput_g14), .B1(n4585), .B2(keyinput_g4), 
        .ZN(n6738) );
  OAI221_X1 U7658 ( .B1(n6739), .B2(keyinput_g14), .C1(n4585), .C2(keyinput_g4), .A(n6738), .ZN(n6744) );
  AOI22_X1 U7659 ( .A1(n6742), .A2(keyinput_g41), .B1(n6741), .B2(keyinput_g53), .ZN(n6740) );
  OAI221_X1 U7660 ( .B1(n6742), .B2(keyinput_g41), .C1(n6741), .C2(
        keyinput_g53), .A(n6740), .ZN(n6743) );
  NOR4_X1 U7661 ( .A1(n6746), .A2(n6745), .A3(n6744), .A4(n6743), .ZN(n6780)
         );
  AOI22_X1 U7662 ( .A1(n6749), .A2(keyinput_g31), .B1(n6748), .B2(keyinput_g8), 
        .ZN(n6747) );
  OAI221_X1 U7663 ( .B1(n6749), .B2(keyinput_g31), .C1(n6748), .C2(keyinput_g8), .A(n6747), .ZN(n6762) );
  AOI22_X1 U7664 ( .A1(n6752), .A2(keyinput_g42), .B1(n6751), .B2(keyinput_g27), .ZN(n6750) );
  OAI221_X1 U7665 ( .B1(n6752), .B2(keyinput_g42), .C1(n6751), .C2(
        keyinput_g27), .A(n6750), .ZN(n6761) );
  AOI22_X1 U7666 ( .A1(n6755), .A2(keyinput_g45), .B1(n6754), .B2(keyinput_g12), .ZN(n6753) );
  OAI221_X1 U7667 ( .B1(n6755), .B2(keyinput_g45), .C1(n6754), .C2(
        keyinput_g12), .A(n6753), .ZN(n6760) );
  AOI22_X1 U7668 ( .A1(n6758), .A2(keyinput_g40), .B1(n6757), .B2(keyinput_g18), .ZN(n6756) );
  OAI221_X1 U7669 ( .B1(n6758), .B2(keyinput_g40), .C1(n6757), .C2(
        keyinput_g18), .A(n6756), .ZN(n6759) );
  NOR4_X1 U7670 ( .A1(n6762), .A2(n6761), .A3(n6760), .A4(n6759), .ZN(n6779)
         );
  AOI22_X1 U7671 ( .A1(n6765), .A2(keyinput_g15), .B1(keyinput_g16), .B2(n6764), .ZN(n6763) );
  OAI221_X1 U7672 ( .B1(n6765), .B2(keyinput_g15), .C1(n6764), .C2(
        keyinput_g16), .A(n6763), .ZN(n6777) );
  AOI22_X1 U7673 ( .A1(n6768), .A2(keyinput_g13), .B1(n6767), .B2(keyinput_g52), .ZN(n6766) );
  OAI221_X1 U7674 ( .B1(n6768), .B2(keyinput_g13), .C1(n6767), .C2(
        keyinput_g52), .A(n6766), .ZN(n6776) );
  AOI22_X1 U7675 ( .A1(n6771), .A2(keyinput_g9), .B1(keyinput_g26), .B2(n6770), 
        .ZN(n6769) );
  OAI221_X1 U7676 ( .B1(n6771), .B2(keyinput_g9), .C1(n6770), .C2(keyinput_g26), .A(n6769), .ZN(n6775) );
  INV_X1 U7677 ( .A(DATAI_14_), .ZN(n6773) );
  AOI22_X1 U7678 ( .A1(n6773), .A2(keyinput_g17), .B1(n4663), .B2(keyinput_g0), 
        .ZN(n6772) );
  OAI221_X1 U7679 ( .B1(n6773), .B2(keyinput_g17), .C1(n4663), .C2(keyinput_g0), .A(n6772), .ZN(n6774) );
  NOR4_X1 U7680 ( .A1(n6777), .A2(n6776), .A3(n6775), .A4(n6774), .ZN(n6778)
         );
  NAND4_X1 U7681 ( .A1(n6781), .A2(n6780), .A3(n6779), .A4(n6778), .ZN(n6782)
         );
  OAI22_X1 U7682 ( .A1(DATAI_1_), .A2(keyinput_g30), .B1(n6783), .B2(n6782), 
        .ZN(n6784) );
  AOI211_X1 U7683 ( .C1(DATAI_1_), .C2(keyinput_g30), .A(n6785), .B(n6784), 
        .ZN(n6788) );
  AOI22_X1 U7684 ( .A1(n6786), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6598), .ZN(n6787) );
  XNOR2_X1 U7685 ( .A(n6788), .B(n6787), .ZN(U3445) );
  AND2_X1 U3572 ( .A1(n3011), .A2(n3012), .ZN(n5631) );
  CLKBUF_X1 U3480 ( .A(n5631), .Z(n3007) );
  CLKBUF_X1 U3575 ( .A(n6128), .Z(n6119) );
endmodule

