

module b21_C_AntiSAT_k_128_4 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049;

  OAI21_X1 U4803 ( .B1(n5449), .B2(n4629), .A(n5453), .ZN(n5471) );
  CLKBUF_X2 U4804 ( .A(n5591), .Z(n5413) );
  INV_X1 U4805 ( .A(n5586), .ZN(n5499) );
  AND3_X1 U4806 ( .A1(n4922), .A2(n4923), .A3(n4921), .ZN(n6920) );
  AND2_X1 U4807 ( .A1(n4851), .A2(n4852), .ZN(n5056) );
  NOR2_X1 U4808 ( .A1(n5607), .A2(n4863), .ZN(n4868) );
  XNOR2_X1 U4809 ( .A(n6296), .B(n6104), .ZN(n8193) );
  INV_X4 U4810 ( .A(n5773), .ZN(n6071) );
  CLKBUF_X1 U4811 ( .A(n6725), .Z(n4300) );
  NAND2_X2 U4812 ( .A1(n5639), .A2(n6565), .ZN(n6574) );
  NAND2_X2 U4813 ( .A1(n6310), .A2(n6783), .ZN(n6769) );
  INV_X1 U4814 ( .A(n5680), .ZN(n8022) );
  NAND2_X1 U4815 ( .A1(n5675), .A2(n8885), .ZN(n5680) );
  XNOR2_X1 U4816 ( .A(n5092), .B(SI_7_), .ZN(n5089) );
  XNOR2_X1 U4817 ( .A(n4968), .B(SI_2_), .ZN(n4966) );
  INV_X1 U4818 ( .A(n6281), .ZN(n6288) );
  INV_X1 U4819 ( .A(n8175), .ZN(n8168) );
  OR2_X1 U4820 ( .A1(n7517), .A2(n7511), .ZN(n7656) );
  NAND2_X1 U4821 ( .A1(n4694), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4693) );
  INV_X2 U4822 ( .A(n5599), .ZN(n4976) );
  NAND4_X1 U4823 ( .A1(n4571), .A2(n4836), .A3(n4569), .A4(n4568), .ZN(n4899)
         );
  AND3_X1 U4824 ( .A1(n5778), .A2(n5777), .A3(n5776), .ZN(n7604) );
  CLKBUF_X3 U4825 ( .A(n5056), .Z(n6344) );
  AOI21_X1 U4827 ( .B1(n9093), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9086), .ZN(
        n9089) );
  AOI21_X1 U4828 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9103), .A(n9100), .ZN(
        n9101) );
  NAND2_X1 U4829 ( .A1(n5490), .A2(n5489), .ZN(n5508) );
  NAND2_X1 U4830 ( .A1(n5914), .A2(n5913), .ZN(n8828) );
  NAND2_X1 U4831 ( .A1(n5692), .A2(n5691), .ZN(n6310) );
  INV_X1 U4832 ( .A(n5679), .ZN(n8890) );
  INV_X1 U4833 ( .A(n9240), .ZN(n9394) );
  XNOR2_X1 U4834 ( .A(n5147), .B(n4824), .ZN(n6660) );
  CLKBUF_X3 U4835 ( .A(n4916), .Z(n4299) );
  NAND4_X1 U4836 ( .A1(n5772), .A2(n5771), .A3(n5770), .A4(n5769), .ZN(n8360)
         );
  INV_X2 U4837 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  AND4_X1 U4838 ( .A1(n4838), .A2(n4875), .A3(n5330), .A4(n4886), .ZN(n4298)
         );
  INV_X4 U4839 ( .A(n5602), .ZN(n5596) );
  OAI211_X1 U4840 ( .C1(n6482), .C2(n6481), .A(n6480), .B(n6479), .ZN(n6484)
         );
  MUX2_X2 U4841 ( .A(n6474), .B(n6473), .S(n6517), .Z(n6482) );
  OAI21_X2 U4842 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        n4696), .ZN(n4695) );
  INV_X2 U4843 ( .A(n5601), .ZN(n5026) );
  AND2_X4 U4844 ( .A1(n6769), .A2(n5700), .ZN(n5880) );
  INV_X2 U4845 ( .A(n6616), .ZN(n5700) );
  XNOR2_X1 U4846 ( .A(n4920), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U4847 ( .A1(n6342), .A2(n6341), .ZN(n9357) );
  OAI21_X1 U4848 ( .B1(n4439), .B2(n4408), .A(n5427), .ZN(n8931) );
  OR2_X1 U4849 ( .A1(n9231), .A2(n9383), .ZN(n9213) );
  NOR3_X1 U4850 ( .A1(n9283), .A2(n9282), .A3(n9281), .ZN(n9280) );
  NAND2_X1 U4851 ( .A1(n5515), .A2(n5514), .ZN(n9389) );
  XNOR2_X1 U4852 ( .A(n5508), .B(n5503), .ZN(n7783) );
  NAND2_X1 U4853 ( .A1(n5973), .A2(n5972), .ZN(n8802) );
  OAI21_X1 U4854 ( .B1(n7913), .B2(n4438), .A(n4304), .ZN(n8041) );
  NAND2_X1 U4855 ( .A1(n5434), .A2(n5433), .ZN(n9409) );
  NAND2_X1 U4856 ( .A1(n5410), .A2(n5409), .ZN(n9414) );
  NAND2_X1 U4857 ( .A1(n5431), .A2(n5430), .ZN(n5449) );
  NAND2_X1 U4858 ( .A1(n5926), .A2(n5925), .ZN(n8824) );
  NAND2_X1 U4859 ( .A1(n5359), .A2(n5358), .ZN(n9423) );
  XNOR2_X1 U4860 ( .A(n5355), .B(n5373), .ZN(n7206) );
  NAND2_X1 U4861 ( .A1(n4404), .A2(n4403), .ZN(n7246) );
  OAI21_X1 U4862 ( .B1(n7540), .B2(n7501), .A(n7500), .ZN(n7788) );
  NAND2_X1 U4863 ( .A1(n4630), .A2(n5326), .ZN(n5371) );
  NAND2_X1 U4864 ( .A1(n5850), .A2(n5849), .ZN(n8108) );
  AND2_X1 U4865 ( .A1(n7657), .A2(n7656), .ZN(n7659) );
  OAI21_X1 U4866 ( .B1(n5299), .B2(n5298), .A(n5297), .ZN(n5325) );
  NOR2_X1 U4867 ( .A1(n8069), .A2(n9671), .ZN(n9702) );
  NAND2_X1 U4868 ( .A1(n5821), .A2(n5820), .ZN(n8855) );
  OAI21_X1 U4869 ( .B1(n5275), .B2(n5274), .A(n5273), .ZN(n5299) );
  NAND2_X2 U4870 ( .A1(n9725), .A2(n7131), .ZN(n9723) );
  INV_X2 U4871 ( .A(n9725), .ZN(n9309) );
  OAI22_X1 U4872 ( .A1(n9808), .A2(n9807), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n9801), .ZN(n9799) );
  NAND2_X2 U4873 ( .A1(n6151), .A2(n6149), .ZN(n6946) );
  XNOR2_X1 U4874 ( .A(n9054), .B(n7214), .ZN(n6889) );
  NOR2_X1 U4875 ( .A1(n6690), .A2(n6689), .ZN(n6688) );
  XNOR2_X1 U4876 ( .A(n5115), .B(n5114), .ZN(n6646) );
  AND3_X1 U4877 ( .A1(n5730), .A2(n5729), .A3(n5728), .ZN(n9952) );
  AND2_X2 U4878 ( .A1(n5586), .A2(n6893), .ZN(n5601) );
  AND2_X2 U4879 ( .A1(n6610), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  AND2_X2 U4880 ( .A1(n4904), .A2(n6890), .ZN(n5586) );
  OR2_X2 U4881 ( .A1(n6891), .A2(n7092), .ZN(n5599) );
  AND4_X1 U4882 ( .A1(n5683), .A2(n5684), .A3(n5681), .A4(n5682), .ZN(n8058)
         );
  OR2_X1 U4883 ( .A1(n9789), .A2(n9788), .ZN(n9791) );
  AND2_X1 U4884 ( .A1(n4867), .A2(n4866), .ZN(n7940) );
  BUF_X2 U4885 ( .A(n5084), .Z(n6317) );
  AND2_X1 U4886 ( .A1(n4426), .A2(n5090), .ZN(n4423) );
  INV_X1 U4887 ( .A(n4852), .ZN(n8024) );
  MUX2_X1 U4888 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4859), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n4862) );
  NAND2_X2 U4889 ( .A1(n8022), .A2(n8890), .ZN(n5963) );
  AND2_X1 U4890 ( .A1(n5679), .A2(n5680), .ZN(n5756) );
  NAND2_X1 U4891 ( .A1(n4903), .A2(n4902), .ZN(n6565) );
  NAND2_X1 U4892 ( .A1(n5690), .A2(n5689), .ZN(n5692) );
  NOR2_X1 U4893 ( .A1(n5612), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4861) );
  MUX2_X1 U4894 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5674), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5675) );
  XNOR2_X1 U4895 ( .A(n4972), .B(SI_3_), .ZN(n4982) );
  NAND2_X1 U4896 ( .A1(n6305), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5694) );
  OR2_X1 U4897 ( .A1(n5676), .A2(n5818), .ZN(n5678) );
  NAND2_X2 U4898 ( .A1(n6617), .A2(P2_U3152), .ZN(n8195) );
  XNOR2_X1 U4899 ( .A(n5013), .B(SI_4_), .ZN(n5010) );
  NOR2_X1 U4900 ( .A1(n4899), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n4847) );
  XNOR2_X1 U4901 ( .A(n5066), .B(SI_6_), .ZN(n5064) );
  NAND2_X2 U4902 ( .A1(n4299), .A2(P1_U3084), .ZN(n9653) );
  AND2_X1 U4903 ( .A1(n4788), .A2(n4787), .ZN(n4786) );
  AND2_X1 U4904 ( .A1(n4984), .A2(n4395), .ZN(n4789) );
  NAND2_X1 U4905 ( .A1(n5672), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5689) );
  AND4_X1 U4906 ( .A1(n5664), .A2(n5663), .A3(n5662), .A4(n5661), .ZN(n5665)
         );
  INV_X1 U4907 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5659) );
  NOR2_X2 U4908 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5657) );
  CLKBUF_X1 U4909 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n9655) );
  INV_X1 U4910 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4886) );
  NOR2_X1 U4911 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n6083) );
  INV_X1 U4912 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5894) );
  OR2_X2 U4913 ( .A1(n8637), .A2(n4511), .ZN(n4510) );
  AND2_X1 U4914 ( .A1(n9174), .A2(n9181), .ZN(n9169) );
  NOR2_X2 U4915 ( .A1(n9373), .A2(n9192), .ZN(n9181) );
  OAI21_X2 U4916 ( .B1(n8559), .B2(n8567), .A(n8481), .ZN(n8540) );
  NOR2_X2 U4917 ( .A1(n8574), .A2(n4538), .ZN(n8559) );
  INV_X1 U4918 ( .A(n5756), .ZN(n4301) );
  INV_X2 U4919 ( .A(n5756), .ZN(n4302) );
  XNOR2_X2 U4920 ( .A(n4985), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9750) );
  NAND2_X1 U4921 ( .A1(n4528), .A2(n4529), .ZN(n7540) );
  INV_X1 U4922 ( .A(n5963), .ZN(n4303) );
  INV_X4 U4923 ( .A(n5963), .ZN(n6018) );
  XNOR2_X2 U4924 ( .A(n5678), .B(n5677), .ZN(n5679) );
  NAND2_X1 U4925 ( .A1(n9005), .A2(n9004), .ZN(n4446) );
  OR2_X1 U4926 ( .A1(n9383), .A2(n9203), .ZN(n9137) );
  OAI21_X1 U4927 ( .B1(n5371), .B2(n5370), .A(n5377), .ZN(n5398) );
  OR2_X1 U4928 ( .A1(n5369), .A2(n5373), .ZN(n5370) );
  AND2_X1 U4929 ( .A1(n5376), .A2(n5375), .ZN(n5377) );
  NOR2_X1 U4930 ( .A1(n4692), .A2(n4425), .ZN(n4424) );
  AND4_X1 U4931 ( .A1(n4324), .A2(n4570), .A3(n4839), .A4(n4840), .ZN(n4569)
         );
  AND2_X1 U4932 ( .A1(n4572), .A2(n4298), .ZN(n4571) );
  INV_X1 U4933 ( .A(n5016), .ZN(n4568) );
  OR2_X1 U4934 ( .A1(n8448), .A2(n6100), .ZN(n6287) );
  NOR2_X1 U4935 ( .A1(n8454), .A2(n4770), .ZN(n4769) );
  INV_X1 U4936 ( .A(n6283), .ZN(n4770) );
  INV_X1 U4937 ( .A(n4429), .ZN(n4428) );
  OAI22_X1 U4938 ( .A1(n9174), .A2(n6521), .B1(n6518), .B2(n6517), .ZN(n4429)
         );
  NAND2_X1 U4939 ( .A1(n9174), .A2(n6518), .ZN(n4430) );
  INV_X1 U4940 ( .A(n8950), .ZN(n9119) );
  AOI21_X1 U4941 ( .B1(n4611), .B2(n4609), .A(n4608), .ZN(n4607) );
  INV_X1 U4942 ( .A(n5249), .ZN(n4608) );
  INV_X1 U4943 ( .A(n4613), .ZN(n4609) );
  OR2_X1 U4944 ( .A1(n8151), .A2(n8150), .ZN(n8152) );
  NAND2_X1 U4945 ( .A1(n7628), .A2(n7629), .ZN(n7635) );
  NAND2_X1 U4946 ( .A1(n8489), .A2(n6279), .ZN(n4682) );
  INV_X1 U4947 ( .A(n7493), .ZN(n7007) );
  AND2_X1 U4948 ( .A1(n6287), .A2(n6285), .ZN(n6137) );
  AND2_X1 U4949 ( .A1(n8448), .A2(n6100), .ZN(n6290) );
  AND2_X1 U4950 ( .A1(n8579), .A2(n6261), .ZN(n4785) );
  AND2_X1 U4951 ( .A1(n6257), .A2(n6252), .ZN(n5989) );
  INV_X1 U4952 ( .A(n4512), .ZN(n4509) );
  NOR2_X1 U4953 ( .A1(n8777), .A2(n8770), .ZN(n8498) );
  INV_X1 U4954 ( .A(n4459), .ZN(n4458) );
  OAI21_X1 U4955 ( .B1(n5596), .B2(n7113), .A(n4410), .ZN(n4977) );
  NAND2_X1 U4956 ( .A1(n5586), .A2(n8978), .ZN(n4410) );
  NAND2_X1 U4957 ( .A1(n4447), .A2(n4446), .ZN(n4444) );
  OR2_X1 U4958 ( .A1(n6920), .A2(n5499), .ZN(n4924) );
  OR2_X1 U4959 ( .A1(n9366), .A2(n6518), .ZN(n6388) );
  OR2_X1 U4960 ( .A1(n9373), .A2(n9197), .ZN(n6509) );
  NAND2_X1 U4961 ( .A1(n9373), .A2(n9197), .ZN(n9160) );
  OR2_X1 U4962 ( .A1(n9379), .A2(n9139), .ZN(n9158) );
  OAI21_X1 U4963 ( .B1(n4563), .B2(n4561), .A(n9132), .ZN(n4560) );
  INV_X1 U4964 ( .A(n4562), .ZN(n4561) );
  NAND2_X1 U4965 ( .A1(n9268), .A2(n9130), .ZN(n4567) );
  OR2_X1 U4966 ( .A1(n9399), .A2(n9131), .ZN(n9153) );
  OR2_X1 U4967 ( .A1(n9409), .A2(n9041), .ZN(n6360) );
  NAND2_X1 U4968 ( .A1(n7816), .A2(n9711), .ZN(n7823) );
  NAND2_X1 U4969 ( .A1(n5576), .A2(n5575), .ZN(n6047) );
  NOR2_X1 U4970 ( .A1(n5016), .A2(n4574), .ZN(n4573) );
  NAND2_X1 U4971 ( .A1(n5325), .A2(n5324), .ZN(n4630) );
  NOR2_X1 U4972 ( .A1(n5226), .A2(n4614), .ZN(n4613) );
  INV_X1 U4973 ( .A(n5196), .ZN(n4614) );
  NAND2_X1 U4974 ( .A1(n4615), .A2(n5148), .ZN(n5170) );
  INV_X1 U4975 ( .A(n5010), .ZN(n5011) );
  NOR2_X1 U4976 ( .A1(n8134), .A2(n4706), .ZN(n4705) );
  INV_X1 U4977 ( .A(n8130), .ZN(n4706) );
  OR2_X1 U4978 ( .A1(n4709), .A2(n8134), .ZN(n4707) );
  AND2_X1 U4979 ( .A1(n8319), .A2(n4710), .ZN(n4709) );
  NAND2_X1 U4980 ( .A1(n8278), .A2(n8130), .ZN(n4710) );
  AOI21_X1 U4982 ( .B1(n4776), .B2(n4777), .A(n4775), .ZN(n4774) );
  INV_X1 U4983 ( .A(n6277), .ZN(n4775) );
  INV_X1 U4984 ( .A(n6019), .ZN(n4776) );
  AND2_X1 U4985 ( .A1(n6031), .A2(n6030), .ZN(n8516) );
  NAND2_X1 U4986 ( .A1(n8541), .A2(n6019), .ZN(n8543) );
  NAND2_X1 U4987 ( .A1(n8586), .A2(n4820), .ZN(n8575) );
  OR2_X1 U4988 ( .A1(n8593), .A2(n8479), .ZN(n4820) );
  NAND2_X1 U4989 ( .A1(n8657), .A2(n8656), .ZN(n4763) );
  OR2_X1 U4990 ( .A1(n8842), .A2(n8458), .ZN(n4527) );
  INV_X1 U4991 ( .A(n4446), .ZN(n4445) );
  AND2_X1 U4992 ( .A1(n6574), .A2(n6617), .ZN(n5021) );
  NOR2_X1 U4993 ( .A1(n7910), .A2(n4791), .ZN(n4790) );
  INV_X1 U4994 ( .A(n5224), .ZN(n4791) );
  NAND2_X1 U4995 ( .A1(n7246), .A2(n5081), .ZN(n5109) );
  AND2_X1 U4996 ( .A1(n9030), .A2(n4461), .ZN(n4459) );
  NAND2_X1 U4997 ( .A1(n5591), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4915) );
  XNOR2_X1 U4998 ( .A(n7922), .B(n7929), .ZN(n7681) );
  OR2_X1 U4999 ( .A1(n4582), .A2(n4353), .ZN(n4580) );
  NOR2_X1 U5000 ( .A1(n6547), .A2(n4584), .ZN(n4582) );
  BUF_X1 U5001 ( .A(n5021), .Z(n6340) );
  NAND2_X1 U5002 ( .A1(n4846), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4848) );
  OAI21_X1 U5003 ( .B1(n4847), .B2(n5122), .A(P1_IR_REG_29__SCAN_IN), .ZN(
        n4849) );
  XNOR2_X1 U5004 ( .A(n4876), .B(n4875), .ZN(n7093) );
  NAND2_X1 U5005 ( .A1(n4466), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4876) );
  INV_X1 U5006 ( .A(n4882), .ZN(n4466) );
  AOI21_X1 U5007 ( .B1(n4885), .B2(n4884), .A(n4883), .ZN(n5383) );
  NOR2_X1 U5008 ( .A1(n5122), .A2(n4838), .ZN(n4884) );
  OR2_X1 U5009 ( .A1(n4882), .A2(n4881), .ZN(n4883) );
  NAND2_X1 U5010 ( .A1(n4880), .A2(n4879), .ZN(n4885) );
  XNOR2_X1 U5011 ( .A(n5038), .B(SI_5_), .ZN(n5036) );
  NAND2_X1 U5012 ( .A1(n5015), .A2(n5014), .ZN(n5037) );
  OAI21_X1 U5013 ( .B1(n4390), .B2(n6196), .A(n6200), .ZN(n4389) );
  AOI21_X1 U5014 ( .B1(n6192), .B2(n6191), .A(n6190), .ZN(n4390) );
  NOR2_X1 U5015 ( .A1(n4419), .A2(n4418), .ZN(n4417) );
  NAND2_X1 U5016 ( .A1(n8008), .A2(n6460), .ZN(n4418) );
  INV_X1 U5017 ( .A(n6455), .ZN(n4419) );
  AND2_X1 U5018 ( .A1(n9339), .A2(n6461), .ZN(n4421) );
  INV_X1 U5019 ( .A(n6462), .ZN(n4422) );
  NAND2_X1 U5020 ( .A1(n4307), .A2(n6460), .ZN(n4420) );
  AND2_X1 U5021 ( .A1(n8247), .A2(n4701), .ZN(n4700) );
  NAND2_X1 U5022 ( .A1(n8301), .A2(n8145), .ZN(n4701) );
  INV_X1 U5023 ( .A(n8145), .ZN(n4698) );
  INV_X1 U5024 ( .A(n5467), .ZN(n4810) );
  AND2_X1 U5025 ( .A1(n9357), .A2(n4617), .ZN(n6415) );
  OR2_X1 U5026 ( .A1(n9357), .A2(n6349), .ZN(n6523) );
  NAND2_X1 U5027 ( .A1(n4628), .A2(n6068), .ZN(n6090) );
  INV_X1 U5028 ( .A(n4611), .ZN(n4610) );
  OR2_X1 U5029 ( .A1(n7620), .A2(n7646), .ZN(n7621) );
  NAND2_X1 U5030 ( .A1(n8156), .A2(n8155), .ZN(n8160) );
  INV_X1 U5031 ( .A(n8288), .ZN(n8156) );
  NAND2_X1 U5032 ( .A1(n4729), .A2(n8116), .ZN(n4728) );
  INV_X1 U5033 ( .A(n8102), .ZN(n4729) );
  NAND2_X1 U5034 ( .A1(n4727), .A2(n8116), .ZN(n4726) );
  INV_X1 U5035 ( .A(n4730), .ZN(n4727) );
  OAI21_X1 U5036 ( .B1(n4392), .B2(n4684), .A(n6276), .ZN(n4391) );
  OAI21_X1 U5037 ( .B1(n4771), .B2(n4768), .A(n4767), .ZN(n4766) );
  NAND2_X1 U5038 ( .A1(n4769), .A2(n6065), .ZN(n4767) );
  AND2_X1 U5039 ( .A1(n6286), .A2(n4772), .ZN(n4771) );
  OR2_X1 U5040 ( .A1(n8776), .A2(n8516), .ZN(n6277) );
  OR2_X1 U5041 ( .A1(n8784), .A2(n8352), .ZN(n6271) );
  NAND2_X1 U5042 ( .A1(n4514), .A2(n8478), .ZN(n4511) );
  INV_X1 U5043 ( .A(n8614), .ZN(n8478) );
  INV_X1 U5044 ( .A(n8628), .ZN(n4755) );
  OR2_X1 U5045 ( .A1(n8802), .A2(n8475), .ZN(n6252) );
  NOR2_X1 U5046 ( .A1(n4494), .A2(n8108), .ZN(n4493) );
  NAND2_X1 U5047 ( .A1(n7990), .A2(n4495), .ZN(n4494) );
  INV_X1 U5048 ( .A(n7895), .ZN(n4525) );
  NAND2_X1 U5049 ( .A1(n6950), .A2(n8554), .ZN(n6956) );
  OR2_X1 U5050 ( .A1(n7794), .A2(n8855), .ZN(n7883) );
  NAND2_X1 U5051 ( .A1(n4740), .A2(n6185), .ZN(n4735) );
  INV_X1 U5052 ( .A(n6169), .ZN(n4743) );
  OAI21_X1 U5053 ( .B1(n7714), .B2(n4741), .A(n6175), .ZN(n4740) );
  NAND2_X1 U5054 ( .A1(n6121), .A2(n6169), .ZN(n4741) );
  NOR2_X1 U5055 ( .A1(n8360), .A2(n7604), .ZN(n6121) );
  OR2_X1 U5056 ( .A1(n7077), .A2(n9952), .ZN(n6117) );
  NAND2_X1 U5057 ( .A1(n7406), .A2(n7311), .ZN(n7428) );
  NAND2_X1 U5058 ( .A1(n8784), .A2(n8352), .ZN(n6272) );
  NOR2_X1 U5059 ( .A1(n4678), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n4677) );
  INV_X1 U5060 ( .A(n4678), .ZN(n4676) );
  NAND2_X1 U5061 ( .A1(n8931), .A2(n8932), .ZN(n5448) );
  XNOR2_X1 U5062 ( .A(n4951), .B(n4976), .ZN(n4952) );
  OR2_X1 U5063 ( .A1(n7908), .A2(n4438), .ZN(n4437) );
  NAND2_X1 U5064 ( .A1(n6316), .A2(n4616), .ZN(n6554) );
  AND2_X1 U5065 ( .A1(n9165), .A2(n6315), .ZN(n4616) );
  AOI21_X1 U5066 ( .B1(n4658), .B2(n6337), .A(n9157), .ZN(n4656) );
  NOR2_X1 U5067 ( .A1(n9227), .A2(n4659), .ZN(n4658) );
  INV_X1 U5068 ( .A(n9155), .ZN(n4659) );
  OR2_X1 U5069 ( .A1(n9389), .A2(n9135), .ZN(n6498) );
  OR2_X1 U5070 ( .A1(n9404), .A2(n9409), .ZN(n4668) );
  NOR2_X1 U5071 ( .A1(n9149), .A2(n4635), .ZN(n4634) );
  INV_X1 U5072 ( .A(n9148), .ZN(n4635) );
  NOR2_X1 U5073 ( .A1(n9146), .A2(n4643), .ZN(n4642) );
  INV_X1 U5074 ( .A(n9331), .ZN(n4590) );
  NAND2_X1 U5075 ( .A1(n4595), .A2(n9331), .ZN(n4592) );
  NOR2_X1 U5076 ( .A1(n9119), .A2(n9439), .ZN(n4675) );
  AND2_X1 U5077 ( .A1(n9119), .A2(n8033), .ZN(n9141) );
  NOR2_X1 U5078 ( .A1(n7829), .A2(n4647), .ZN(n4646) );
  INV_X1 U5079 ( .A(n7827), .ZN(n4647) );
  NOR2_X1 U5080 ( .A1(n4549), .A2(n4305), .ZN(n4548) );
  INV_X1 U5081 ( .A(n4554), .ZN(n4549) );
  AND2_X1 U5082 ( .A1(n4348), .A2(n7474), .ZN(n4600) );
  NOR2_X1 U5083 ( .A1(n7243), .A2(n9023), .ZN(n4673) );
  NAND2_X1 U5084 ( .A1(n7331), .A2(n7329), .ZN(n4602) );
  AOI21_X1 U5085 ( .B1(n7826), .B2(n7825), .A(n7824), .ZN(n9689) );
  NAND2_X1 U5086 ( .A1(n7115), .A2(n7121), .ZN(n7225) );
  NAND2_X1 U5087 ( .A1(n7114), .A2(n7276), .ZN(n7115) );
  INV_X1 U5088 ( .A(n4899), .ZN(n4896) );
  NAND2_X1 U5089 ( .A1(n4627), .A2(n5554), .ZN(n5576) );
  INV_X1 U5090 ( .A(n4622), .ZN(n4621) );
  AOI21_X1 U5091 ( .B1(n4622), .B2(n4624), .A(n4620), .ZN(n4619) );
  AND3_X1 U5092 ( .A1(n4576), .A2(n4324), .A3(n4298), .ZN(n4844) );
  INV_X1 U5093 ( .A(n5450), .ZN(n4629) );
  AND2_X1 U5094 ( .A1(n5326), .A2(n5305), .ZN(n5324) );
  OR2_X1 U5095 ( .A1(n4857), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5253) );
  AND2_X1 U5096 ( .A1(n5251), .A2(n5231), .ZN(n5249) );
  AOI21_X1 U5097 ( .B1(n4613), .B2(n5197), .A(n4612), .ZN(n4611) );
  INV_X1 U5098 ( .A(n5225), .ZN(n4612) );
  AND4_X1 U5099 ( .A1(n4835), .A2(n4834), .A3(n5068), .A4(n4833), .ZN(n4836)
         );
  NAND2_X1 U5100 ( .A1(n5225), .A2(n5204), .ZN(n5226) );
  INV_X1 U5101 ( .A(n5193), .ZN(n5197) );
  NAND2_X1 U5102 ( .A1(n5172), .A2(n5171), .ZN(n5198) );
  NAND2_X1 U5103 ( .A1(n5113), .A2(n5099), .ZN(n5114) );
  OAI21_X1 U5104 ( .B1(n5036), .B2(n4692), .A(n5064), .ZN(n4691) );
  NAND2_X1 U5105 ( .A1(n4688), .A2(n4982), .ZN(n4686) );
  AND2_X1 U5106 ( .A1(n4713), .A2(n8169), .ZN(n4712) );
  AOI21_X1 U5107 ( .B1(n7151), .B2(n7150), .A(n7076), .ZN(n7084) );
  AOI21_X1 U5108 ( .B1(n8279), .B2(n4325), .A(n4703), .ZN(n8225) );
  NOR2_X1 U5109 ( .A1(n4707), .A2(n4704), .ZN(n4703) );
  INV_X1 U5110 ( .A(n8226), .ZN(n4704) );
  INV_X1 U5111 ( .A(n7635), .ZN(n7633) );
  OR2_X1 U5112 ( .A1(n6012), .A2(n8330), .ZN(n6024) );
  OR3_X1 U5113 ( .A1(n7813), .A2(n7950), .A3(n7945), .ZN(n7061) );
  INV_X1 U5114 ( .A(n6957), .ZN(n6947) );
  OR2_X1 U5115 ( .A1(n6832), .A2(n6831), .ZN(n4471) );
  NAND2_X1 U5116 ( .A1(n4471), .A2(n4470), .ZN(n4469) );
  NAND2_X1 U5117 ( .A1(n6804), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4470) );
  AND2_X1 U5118 ( .A1(n4469), .A2(n4468), .ZN(n6854) );
  INV_X1 U5119 ( .A(n6855), .ZN(n4468) );
  NAND2_X1 U5120 ( .A1(n6098), .A2(n6097), .ZN(n8448) );
  NAND2_X1 U5121 ( .A1(n8498), .A2(n8502), .ZN(n8497) );
  NAND2_X1 U5122 ( .A1(n6057), .A2(n6056), .ZN(n8766) );
  AND2_X1 U5123 ( .A1(n6043), .A2(n6042), .ZN(n8488) );
  AND2_X1 U5124 ( .A1(n6064), .A2(n6063), .ZN(n8517) );
  INV_X1 U5125 ( .A(n8507), .ZN(n8514) );
  AND2_X1 U5126 ( .A1(n6278), .A2(n6275), .ZN(n8507) );
  OR2_X1 U5127 ( .A1(n8485), .A2(n8776), .ZN(n8486) );
  INV_X1 U5128 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5939) );
  OR2_X1 U5129 ( .A1(n8788), .A2(n8580), .ZN(n8481) );
  OAI21_X1 U5130 ( .B1(n8613), .B2(n4784), .A(n4781), .ZN(n6009) );
  AOI21_X1 U5131 ( .B1(n4785), .B2(n4783), .A(n4782), .ZN(n4781) );
  INV_X1 U5132 ( .A(n4785), .ZN(n4784) );
  AND2_X1 U5133 ( .A1(n8605), .A2(n4483), .ZN(n8560) );
  NOR2_X1 U5134 ( .A1(n8788), .A2(n4485), .ZN(n4483) );
  XNOR2_X1 U5135 ( .A(n8788), .B(n8580), .ZN(n8567) );
  AND2_X1 U5136 ( .A1(n8566), .A2(n6263), .ZN(n8579) );
  NAND2_X1 U5137 ( .A1(n8615), .A2(n8614), .ZN(n8613) );
  AOI21_X1 U5138 ( .B1(n4514), .B2(n6112), .A(n4334), .ZN(n4512) );
  AND2_X1 U5139 ( .A1(n6252), .A2(n6253), .ZN(n8614) );
  OAI21_X1 U5140 ( .B1(n8688), .B2(n5937), .A(n6228), .ZN(n8657) );
  NOR2_X1 U5141 ( .A1(n8824), .A2(n8468), .ZN(n4537) );
  NOR2_X1 U5142 ( .A1(n8689), .A2(n8690), .ZN(n8688) );
  NOR2_X1 U5143 ( .A1(n8697), .A2(n8464), .ZN(n8682) );
  AND2_X1 U5144 ( .A1(n8832), .A2(n8463), .ZN(n8464) );
  OR2_X1 U5145 ( .A1(n8717), .A2(n8832), .ZN(n8700) );
  OR2_X1 U5146 ( .A1(n7902), .A2(n8355), .ZN(n7872) );
  NAND2_X1 U5147 ( .A1(n4526), .A2(n4525), .ZN(n4524) );
  INV_X1 U5148 ( .A(n7890), .ZN(n4526) );
  OR2_X1 U5149 ( .A1(n8001), .A2(n6959), .ZN(n8728) );
  AND2_X1 U5150 ( .A1(n7720), .A2(n7764), .ZN(n7670) );
  AOI21_X1 U5151 ( .B1(n4530), .B2(n4533), .A(n4335), .ZN(n4529) );
  NAND2_X1 U5152 ( .A1(n8751), .A2(n8750), .ZN(n8749) );
  INV_X1 U5153 ( .A(n8728), .ZN(n8632) );
  INV_X1 U5154 ( .A(n8724), .ZN(n8740) );
  AND2_X1 U5155 ( .A1(n8766), .A2(n8856), .ZN(n8767) );
  NAND2_X1 U5156 ( .A1(n6033), .A2(n6032), .ZN(n8770) );
  OR2_X1 U5157 ( .A1(n8529), .A2(n8776), .ZN(n8777) );
  NAND2_X1 U5158 ( .A1(n5943), .A2(n5942), .ZN(n8818) );
  OR2_X1 U5159 ( .A1(n7303), .A2(n6961), .ZN(n9981) );
  NAND2_X1 U5160 ( .A1(n7061), .A2(n9937), .ZN(n9926) );
  NOR2_X1 U5161 ( .A1(n4794), .A2(n4407), .ZN(n4405) );
  INV_X1 U5162 ( .A(n8940), .ZN(n4457) );
  NOR2_X1 U5163 ( .A1(n4458), .A2(n4455), .ZN(n4454) );
  INV_X1 U5164 ( .A(n4462), .ZN(n4455) );
  NAND2_X1 U5165 ( .A1(n8965), .A2(n4462), .ZN(n4453) );
  NOR2_X1 U5166 ( .A1(n9005), .A2(n9004), .ZN(n4447) );
  AND2_X1 U5167 ( .A1(n4805), .A2(n4803), .ZN(n8902) );
  NOR2_X1 U5168 ( .A1(n4804), .A2(n5486), .ZN(n4803) );
  INV_X1 U5169 ( .A(n4808), .ZN(n4804) );
  NAND2_X1 U5170 ( .A1(n4432), .A2(n4999), .ZN(n8974) );
  NAND2_X1 U5171 ( .A1(n6868), .A2(n4394), .ZN(n4432) );
  OR2_X1 U5172 ( .A1(n5109), .A2(n5110), .ZN(n8920) );
  AOI21_X1 U5173 ( .B1(n9007), .B2(n4317), .A(n4440), .ZN(n4439) );
  NAND2_X1 U5174 ( .A1(n4441), .A2(n5397), .ZN(n4440) );
  NAND2_X1 U5175 ( .A1(n4317), .A2(n4445), .ZN(n4441) );
  NAND2_X1 U5176 ( .A1(n7776), .A2(n5221), .ZN(n4792) );
  NAND2_X1 U5177 ( .A1(n5529), .A2(n5528), .ZN(n4461) );
  NAND2_X1 U5178 ( .A1(n8939), .A2(n8940), .ZN(n4460) );
  AND4_X1 U5179 ( .A1(n5644), .A2(n5643), .A3(n5642), .A4(n5641), .ZN(n6518)
         );
  AND4_X1 U5180 ( .A1(n5569), .A2(n5568), .A3(n5567), .A4(n5566), .ZN(n9139)
         );
  AND4_X1 U5181 ( .A1(n5484), .A2(n5483), .A3(n5482), .A4(n5481), .ZN(n9131)
         );
  AND4_X1 U5182 ( .A1(n5216), .A2(n5215), .A3(n5214), .A4(n5213), .ZN(n9711)
         );
  NAND2_X1 U5183 ( .A1(n6708), .A2(n6587), .ZN(n6690) );
  NOR2_X1 U5184 ( .A1(n7679), .A2(n7680), .ZN(n7922) );
  NAND2_X1 U5185 ( .A1(n6323), .A2(n6322), .ZN(n9366) );
  AND2_X1 U5186 ( .A1(n6388), .A2(n6550), .ZN(n9161) );
  AND2_X1 U5187 ( .A1(n5640), .A2(n5590), .ZN(n9182) );
  NAND2_X1 U5188 ( .A1(n4579), .A2(n4578), .ZN(n9178) );
  NOR2_X1 U5189 ( .A1(n4580), .A2(n9187), .ZN(n4578) );
  AND2_X1 U5190 ( .A1(n4585), .A2(n9137), .ZN(n4584) );
  OR2_X1 U5191 ( .A1(n4586), .A2(n9138), .ZN(n4585) );
  AND2_X1 U5192 ( .A1(n9227), .A2(n6338), .ZN(n4583) );
  AND2_X1 U5193 ( .A1(n9241), .A2(n4658), .ZN(n9225) );
  NAND2_X1 U5194 ( .A1(n9134), .A2(n9133), .ZN(n9222) );
  OR2_X1 U5195 ( .A1(n9394), .A2(n9230), .ZN(n9133) );
  NAND2_X1 U5196 ( .A1(n9394), .A2(n9230), .ZN(n4566) );
  NAND2_X1 U5197 ( .A1(n6498), .A2(n6496), .ZN(n9227) );
  NAND2_X1 U5198 ( .A1(n9243), .A2(n9242), .ZN(n9241) );
  AND2_X1 U5199 ( .A1(n4567), .A2(n9281), .ZN(n4563) );
  NAND2_X1 U5200 ( .A1(n4341), .A2(n4567), .ZN(n4562) );
  AND2_X1 U5201 ( .A1(n9299), .A2(n9312), .ZN(n9282) );
  NAND2_X1 U5202 ( .A1(n6360), .A2(n6475), .ZN(n9281) );
  OR2_X1 U5203 ( .A1(n9414), .A2(n9312), .ZN(n9126) );
  AND2_X1 U5204 ( .A1(n4639), .A2(n4638), .ZN(n4637) );
  NAND2_X1 U5205 ( .A1(n4640), .A2(n9145), .ZN(n4639) );
  INV_X1 U5206 ( .A(n9147), .ZN(n4640) );
  AOI21_X1 U5207 ( .B1(n4595), .B2(n9120), .A(n4312), .ZN(n4593) );
  OR2_X1 U5208 ( .A1(n9439), .A2(n9042), .ZN(n7977) );
  NOR2_X1 U5209 ( .A1(n6458), .A2(n9141), .ZN(n9142) );
  NAND2_X1 U5210 ( .A1(n4649), .A2(n9688), .ZN(n4648) );
  INV_X1 U5211 ( .A(n9689), .ZN(n4649) );
  OR2_X1 U5212 ( .A1(n9704), .A2(n7816), .ZN(n4828) );
  NOR2_X1 U5213 ( .A1(n7817), .A2(n4555), .ZN(n4554) );
  INV_X1 U5214 ( .A(n7748), .ZN(n4555) );
  NAND2_X1 U5215 ( .A1(n7825), .A2(n4556), .ZN(n4552) );
  OR2_X1 U5216 ( .A1(n9701), .A2(n7747), .ZN(n7749) );
  AND4_X1 U5217 ( .A1(n5163), .A2(n5162), .A3(n5161), .A4(n5160), .ZN(n9713)
         );
  AND2_X1 U5218 ( .A1(n7478), .A2(n7480), .ZN(n7334) );
  NAND2_X1 U5219 ( .A1(n7330), .A2(n4601), .ZN(n7475) );
  INV_X1 U5220 ( .A(n4602), .ZN(n4601) );
  AND4_X1 U5221 ( .A1(n5033), .A2(n5032), .A3(n5031), .A4(n5030), .ZN(n7322)
         );
  AND4_X1 U5222 ( .A1(n5063), .A2(n5062), .A3(n5061), .A4(n5060), .ZN(n7336)
         );
  OR2_X1 U5223 ( .A1(n6734), .A2(n6894), .ZN(n9710) );
  OR2_X1 U5224 ( .A1(n7263), .A2(n8978), .ZN(n7280) );
  OAI211_X1 U5225 ( .C1(n4991), .C2(n6633), .A(n4990), .B(n4989), .ZN(n7267)
         );
  OR2_X1 U5226 ( .A1(n4991), .A2(n6618), .ZN(n4923) );
  INV_X1 U5227 ( .A(n9710), .ZN(n9349) );
  INV_X1 U5228 ( .A(n9365), .ZN(n9370) );
  NAND2_X1 U5229 ( .A1(n5585), .A2(n5584), .ZN(n9373) );
  INV_X1 U5230 ( .A(n8978), .ZN(n9847) );
  NAND2_X1 U5231 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4546), .ZN(n4545) );
  INV_X1 U5232 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4546) );
  NOR2_X1 U5233 ( .A1(n4846), .A2(P1_IR_REG_30__SCAN_IN), .ZN(n4544) );
  XNOR2_X1 U5234 ( .A(n5576), .B(n5575), .ZN(n7964) );
  XNOR2_X1 U5235 ( .A(n5553), .B(n5552), .ZN(n7942) );
  NAND2_X1 U5236 ( .A1(n4618), .A2(n4622), .ZN(n5553) );
  NAND2_X1 U5237 ( .A1(n5508), .A2(n4625), .ZN(n4618) );
  NAND2_X1 U5238 ( .A1(n4813), .A2(n4844), .ZN(n4866) );
  INV_X1 U5239 ( .A(n4857), .ZN(n4813) );
  XNOR2_X1 U5240 ( .A(n4890), .B(n4889), .ZN(n5636) );
  XNOR2_X1 U5241 ( .A(n4431), .B(n5226), .ZN(n6698) );
  OAI21_X1 U5242 ( .B1(n5198), .B2(n5197), .A(n5196), .ZN(n4431) );
  INV_X1 U5243 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4397) );
  INV_X1 U5244 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4395) );
  NAND2_X1 U5245 ( .A1(n5866), .A2(n5865), .ZN(n8842) );
  NAND2_X1 U5246 ( .A1(n5983), .A2(n5982), .ZN(n8797) );
  AND2_X1 U5247 ( .A1(n8282), .A2(n8630), .ZN(n8240) );
  NAND2_X1 U5248 ( .A1(n5962), .A2(n5961), .ZN(n8807) );
  NAND2_X1 U5249 ( .A1(n5951), .A2(n5950), .ZN(n8812) );
  INV_X1 U5250 ( .A(n8193), .ZN(n6950) );
  NAND2_X1 U5251 ( .A1(n4382), .A2(n4381), .ZN(n4380) );
  OR2_X1 U5252 ( .A1(n4681), .A2(n4383), .ZN(n4382) );
  NOR2_X1 U5253 ( .A1(n6294), .A2(n6961), .ZN(n4681) );
  AND2_X1 U5254 ( .A1(n6109), .A2(n7702), .ZN(n4745) );
  INV_X1 U5255 ( .A(n8766), .ZN(n8502) );
  OAI211_X1 U5256 ( .C1(n5773), .C2(n6633), .A(n5718), .B(n5717), .ZN(n7445)
         );
  INV_X1 U5257 ( .A(n9033), .ZN(n9008) );
  AND4_X1 U5258 ( .A1(n5439), .A2(n5438), .A3(n5437), .A4(n5436), .ZN(n9041)
         );
  AND2_X1 U5259 ( .A1(n4797), .A2(n4401), .ZN(n4400) );
  OR2_X1 U5260 ( .A1(n5109), .A2(n4399), .ZN(n4398) );
  AND2_X1 U5261 ( .A1(n5145), .A2(n8059), .ZN(n4797) );
  NAND2_X1 U5262 ( .A1(n8059), .A2(n4796), .ZN(n4795) );
  INV_X1 U5263 ( .A(n5146), .ZN(n4796) );
  NAND2_X1 U5264 ( .A1(n4449), .A2(n4448), .ZN(n7694) );
  AND2_X1 U5265 ( .A1(n7695), .A2(n4308), .ZN(n4448) );
  NAND2_X1 U5266 ( .A1(n6526), .A2(n7099), .ZN(n4412) );
  NAND2_X1 U5267 ( .A1(n4414), .A2(n9110), .ZN(n4413) );
  NAND2_X1 U5268 ( .A1(n5209), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4912) );
  NOR2_X1 U5269 ( .A1(n7467), .A2(n7466), .ZN(n7679) );
  OAI21_X1 U5270 ( .B1(n9108), .B2(n9107), .A(n4500), .ZN(n4499) );
  AOI21_X1 U5271 ( .B1(n9109), .B2(n9823), .A(n9825), .ZN(n4500) );
  NAND3_X1 U5272 ( .A1(n5024), .A2(n5023), .A3(n5022), .ZN(n7286) );
  INV_X1 U5273 ( .A(n5636), .ZN(n7538) );
  CLKBUF_X1 U5274 ( .A(n5383), .Z(n9110) );
  OAI21_X1 U5275 ( .B1(n6160), .B2(n6141), .A(n4685), .ZN(n6142) );
  AND2_X1 U5276 ( .A1(n6163), .A2(n6140), .ZN(n4685) );
  NAND3_X1 U5277 ( .A1(n6148), .A2(n6147), .A3(n7430), .ZN(n4386) );
  NAND2_X1 U5278 ( .A1(n4389), .A2(n7876), .ZN(n4388) );
  INV_X1 U5279 ( .A(n6369), .ZN(n6444) );
  NAND2_X1 U5280 ( .A1(n4342), .A2(n4421), .ZN(n4415) );
  NAND2_X1 U5281 ( .A1(n6438), .A2(n6405), .ZN(n6369) );
  NAND2_X1 U5282 ( .A1(n7823), .A2(n7755), .ZN(n6405) );
  OAI21_X1 U5283 ( .B1(n6268), .B2(n6267), .A(n6266), .ZN(n4393) );
  OR2_X1 U5284 ( .A1(n8524), .A2(n6273), .ZN(n4684) );
  OR2_X1 U5285 ( .A1(n8812), .A2(n8250), .ZN(n6241) );
  AND2_X1 U5286 ( .A1(n4787), .A2(n5693), .ZN(n4534) );
  AND2_X1 U5287 ( .A1(n5660), .A2(n5671), .ZN(n4535) );
  INV_X1 U5288 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4787) );
  NAND2_X1 U5289 ( .A1(n5894), .A2(n4679), .ZN(n4678) );
  INV_X1 U5290 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4780) );
  NAND2_X1 U5291 ( .A1(n4814), .A2(n4575), .ZN(n4574) );
  INV_X1 U5292 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4575) );
  AND2_X1 U5293 ( .A1(n4837), .A2(n4815), .ZN(n4814) );
  INV_X1 U5294 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4815) );
  INV_X1 U5295 ( .A(n5552), .ZN(n4620) );
  NAND2_X1 U5296 ( .A1(n5202), .A2(n5201), .ZN(n5225) );
  NAND2_X1 U5297 ( .A1(n5118), .A2(n5117), .ZN(n5148) );
  NAND2_X1 U5298 ( .A1(n5097), .A2(n5096), .ZN(n5113) );
  INV_X1 U5299 ( .A(n4970), .ZN(n4688) );
  NAND2_X1 U5300 ( .A1(n4715), .A2(n4719), .ZN(n4713) );
  AOI21_X1 U5301 ( .B1(n4726), .B2(n4728), .A(n4322), .ZN(n4724) );
  OAI21_X1 U5302 ( .B1(n8302), .B2(n4699), .A(n4697), .ZN(n8151) );
  AOI21_X1 U5303 ( .B1(n4700), .B2(n4698), .A(n4326), .ZN(n4697) );
  INV_X1 U5304 ( .A(n4700), .ZN(n4699) );
  OR2_X1 U5305 ( .A1(n8766), .A2(n8517), .ZN(n6282) );
  INV_X1 U5306 ( .A(n5989), .ZN(n4783) );
  NOR2_X1 U5307 ( .A1(n8797), .A2(n8802), .ZN(n4487) );
  AND2_X1 U5308 ( .A1(n6258), .A2(n6261), .ZN(n6257) );
  OR2_X1 U5309 ( .A1(n5953), .A2(n5952), .ZN(n5965) );
  OR2_X1 U5310 ( .A1(n8818), .A2(n8828), .ZN(n4504) );
  OR2_X1 U5311 ( .A1(n5916), .A2(n5915), .ZN(n5929) );
  NOR2_X1 U5312 ( .A1(n7993), .A2(n4752), .ZN(n4751) );
  INV_X1 U5313 ( .A(n4751), .ZN(n4749) );
  AND2_X1 U5314 ( .A1(n7496), .A2(n4531), .ZN(n4530) );
  NAND2_X1 U5315 ( .A1(n4532), .A2(n7412), .ZN(n4531) );
  INV_X1 U5316 ( .A(n8750), .ZN(n4532) );
  INV_X1 U5317 ( .A(n7412), .ZN(n4533) );
  AND2_X1 U5318 ( .A1(n6141), .A2(n7428), .ZN(n5731) );
  AND2_X1 U5319 ( .A1(n8736), .A2(n6117), .ZN(n6141) );
  OR2_X1 U5320 ( .A1(n8828), .A2(n8272), .ZN(n8669) );
  INV_X1 U5322 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5672) );
  AND2_X1 U5323 ( .A1(n5774), .A2(n4535), .ZN(n4536) );
  INV_X1 U5324 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4891) );
  OR2_X1 U5325 ( .A1(n5794), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5817) );
  INV_X1 U5326 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5057) );
  AND2_X1 U5327 ( .A1(n4998), .A2(n7023), .ZN(n4394) );
  NAND2_X1 U5328 ( .A1(n8994), .A2(n4810), .ZN(n4808) );
  NOR2_X1 U5329 ( .A1(n4809), .A2(n4807), .ZN(n4806) );
  INV_X1 U5330 ( .A(n5447), .ZN(n4807) );
  NOR2_X1 U5331 ( .A1(n8994), .A2(n4810), .ZN(n4809) );
  NAND2_X1 U5332 ( .A1(n6522), .A2(n4332), .ZN(n6529) );
  OAI21_X1 U5333 ( .B1(n6515), .B2(n4430), .A(n4333), .ZN(n6520) );
  AND2_X1 U5334 ( .A1(n6677), .A2(n6583), .ZN(n9767) );
  INV_X1 U5335 ( .A(n4574), .ZN(n4572) );
  NOR2_X1 U5336 ( .A1(n5480), .A2(n8907), .ZN(n5494) );
  NAND2_X1 U5337 ( .A1(n9258), .A2(n4667), .ZN(n4666) );
  INV_X1 U5338 ( .A(n4668), .ZN(n4667) );
  NOR2_X1 U5339 ( .A1(n5435), .A2(n8933), .ZN(n5461) );
  OR2_X1 U5340 ( .A1(n5336), .A2(n5335), .ZN(n5361) );
  AND2_X1 U5341 ( .A1(n5286), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5310) );
  OR2_X1 U5342 ( .A1(n5236), .A2(n5235), .ZN(n5260) );
  NOR2_X1 U5343 ( .A1(n5179), .A2(n5178), .ZN(n5211) );
  OR2_X1 U5344 ( .A1(n5158), .A2(n5157), .ZN(n5179) );
  NOR3_X1 U5345 ( .A1(n9295), .A2(n9394), .A3(n4666), .ZN(n9246) );
  OR2_X1 U5346 ( .A1(n7199), .A2(n7538), .ZN(n6893) );
  AND2_X1 U5347 ( .A1(n7099), .A2(n7538), .ZN(n6891) );
  XNOR2_X1 U5348 ( .A(n6090), .B(n6089), .ZN(n6087) );
  INV_X1 U5349 ( .A(n5506), .ZN(n4626) );
  AOI21_X1 U5350 ( .B1(n5507), .B2(n4625), .A(n4623), .ZN(n4622) );
  INV_X1 U5351 ( .A(n5530), .ZN(n4623) );
  NAND2_X1 U5352 ( .A1(n5488), .A2(n5487), .ZN(n5490) );
  OR2_X1 U5353 ( .A1(n4857), .A2(n4858), .ZN(n5612) );
  NAND2_X1 U5354 ( .A1(n4576), .A2(n4298), .ZN(n4858) );
  OAI21_X1 U5355 ( .B1(n5471), .B2(n5470), .A(n5469), .ZN(n5488) );
  OAI21_X1 U5356 ( .B1(n4874), .B2(n4464), .A(n4463), .ZN(n4887) );
  AOI21_X1 U5357 ( .B1(n4465), .B2(n5122), .A(n5122), .ZN(n4463) );
  INV_X1 U5358 ( .A(n4465), .ZN(n4464) );
  AOI21_X1 U5359 ( .B1(n4873), .B2(P1_IR_REG_31__SCAN_IN), .A(
        P1_IR_REG_20__SCAN_IN), .ZN(n4465) );
  NAND2_X1 U5360 ( .A1(n5403), .A2(n5402), .ZN(n5429) );
  NAND2_X1 U5361 ( .A1(n5401), .A2(n5400), .ZN(n5403) );
  AND2_X1 U5362 ( .A1(n5430), .A2(n5408), .ZN(n5428) );
  NAND2_X1 U5363 ( .A1(n4605), .A2(n4603), .ZN(n5275) );
  AOI21_X1 U5364 ( .B1(n4607), .B2(n4610), .A(n4604), .ZN(n4603) );
  INV_X1 U5365 ( .A(n5251), .ZN(n4604) );
  INV_X1 U5366 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4837) );
  XNOR2_X1 U5367 ( .A(n5194), .B(SI_11_), .ZN(n5193) );
  INV_X1 U5368 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5068) );
  OR2_X1 U5369 ( .A1(n8092), .A2(n8091), .ZN(n4731) );
  NOR2_X1 U5370 ( .A1(n8094), .A2(n4723), .ZN(n4730) );
  INV_X1 U5371 ( .A(n4731), .ZN(n4723) );
  OR2_X1 U5372 ( .A1(n8101), .A2(n8102), .ZN(n4732) );
  OR2_X1 U5373 ( .A1(n5985), .A2(n5984), .ZN(n5993) );
  NAND2_X1 U5374 ( .A1(n7621), .A2(n4331), .ZN(n7629) );
  OR2_X1 U5375 ( .A1(n5884), .A2(n5883), .ZN(n5901) );
  OR2_X1 U5376 ( .A1(n8153), .A2(n4359), .ZN(n8288) );
  OR2_X1 U5377 ( .A1(n5798), .A2(n9586), .ZN(n5826) );
  AND2_X1 U5378 ( .A1(n8327), .A2(n4716), .ZN(n4715) );
  NAND2_X1 U5379 ( .A1(n4718), .A2(n4717), .ZN(n4716) );
  INV_X1 U5380 ( .A(n4720), .ZN(n4717) );
  OR2_X1 U5381 ( .A1(n8164), .A2(n4721), .ZN(n4720) );
  INV_X1 U5382 ( .A(n8255), .ZN(n4721) );
  AOI211_X1 U5383 ( .C1(n8480), .C2(n8291), .A(n8289), .B(n8206), .ZN(n8162)
         );
  OR2_X1 U5384 ( .A1(n8101), .A2(n4728), .ZN(n4725) );
  OAI21_X1 U5385 ( .B1(n4683), .B2(n4682), .A(n4329), .ZN(n6292) );
  INV_X1 U5386 ( .A(n4766), .ZN(n4765) );
  OR2_X1 U5387 ( .A1(n5963), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U5388 ( .A1(n9658), .A2(n9659), .ZN(n9657) );
  AND2_X1 U5389 ( .A1(n9657), .A2(n4480), .ZN(n6776) );
  NAND2_X1 U5390 ( .A1(n6782), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4480) );
  NOR2_X1 U5391 ( .A1(n6776), .A2(n6775), .ZN(n6791) );
  NOR2_X1 U5392 ( .A1(n6854), .A2(n4467), .ZN(n6820) );
  AND2_X1 U5393 ( .A1(n6802), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4467) );
  OR2_X1 U5394 ( .A1(n6843), .A2(n6842), .ZN(n4475) );
  OR2_X1 U5395 ( .A1(n6904), .A2(n6903), .ZN(n4473) );
  NOR2_X1 U5396 ( .A1(n7396), .A2(n4479), .ZN(n7398) );
  AND2_X1 U5397 ( .A1(n7397), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4479) );
  NOR2_X1 U5398 ( .A1(n7399), .A2(n7398), .ZN(n7561) );
  NOR2_X1 U5399 ( .A1(n7561), .A2(n4478), .ZN(n8371) );
  AND2_X1 U5400 ( .A1(n7562), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4478) );
  NAND2_X1 U5401 ( .A1(n8371), .A2(n8372), .ZN(n8370) );
  NOR2_X1 U5402 ( .A1(n8418), .A2(n4378), .ZN(n8422) );
  NAND2_X1 U5403 ( .A1(n8422), .A2(n8421), .ZN(n8430) );
  NOR2_X1 U5404 ( .A1(n8454), .A2(n8497), .ZN(n8453) );
  NAND2_X1 U5405 ( .A1(n6282), .A2(n6283), .ZN(n8492) );
  NAND2_X1 U5406 ( .A1(n6271), .A2(n6272), .ZN(n8546) );
  NOR2_X1 U5407 ( .A1(n8792), .A2(n4539), .ZN(n4538) );
  NAND2_X1 U5408 ( .A1(n8605), .A2(n4487), .ZN(n8588) );
  AOI21_X1 U5409 ( .B1(n4509), .B2(n8478), .A(n8477), .ZN(n4508) );
  NOR2_X1 U5410 ( .A1(n8802), .A2(n8476), .ZN(n8477) );
  INV_X1 U5411 ( .A(n6257), .ZN(n8594) );
  NAND2_X1 U5412 ( .A1(n4761), .A2(n4757), .ZN(n4756) );
  OAI21_X1 U5413 ( .B1(n4758), .B2(n4755), .A(n4757), .ZN(n4754) );
  INV_X1 U5414 ( .A(n6248), .ZN(n4757) );
  AND2_X1 U5415 ( .A1(n8638), .A2(n8627), .ZN(n8605) );
  NAND2_X1 U5416 ( .A1(n8605), .A2(n8612), .ZN(n8606) );
  NOR3_X1 U5417 ( .A1(n8700), .A2(n4502), .A3(n8824), .ZN(n8638) );
  OR2_X1 U5418 ( .A1(n8812), .A2(n4504), .ZN(n4502) );
  NAND2_X1 U5419 ( .A1(n8681), .A2(n8467), .ZN(n8663) );
  NAND2_X1 U5420 ( .A1(n8669), .A2(n6218), .ZN(n8690) );
  NAND2_X1 U5421 ( .A1(n8682), .A2(n8690), .ZN(n8681) );
  OR2_X1 U5422 ( .A1(n8837), .A2(n8273), .ZN(n8705) );
  OR2_X1 U5423 ( .A1(n8837), .A2(n8461), .ZN(n8462) );
  AND2_X1 U5424 ( .A1(n6208), .A2(n6207), .ZN(n8707) );
  NOR2_X1 U5425 ( .A1(n8698), .A2(n8707), .ZN(n8697) );
  NAND2_X1 U5426 ( .A1(n7879), .A2(n4751), .ZN(n4750) );
  INV_X1 U5427 ( .A(n4746), .ZN(n8723) );
  AOI21_X1 U5428 ( .B1(n7879), .B2(n4748), .A(n4747), .ZN(n4746) );
  NOR2_X1 U5429 ( .A1(n8725), .A2(n5877), .ZN(n4747) );
  NOR2_X1 U5430 ( .A1(n8725), .A2(n4749), .ZN(n4748) );
  NAND2_X1 U5431 ( .A1(n4493), .A2(n8722), .ZN(n4492) );
  NAND2_X1 U5432 ( .A1(n8705), .A2(n6214), .ZN(n8725) );
  INV_X1 U5433 ( .A(n4493), .ZN(n4491) );
  INV_X1 U5434 ( .A(n4521), .ZN(n4520) );
  OAI21_X1 U5435 ( .B1(n4525), .B2(n4523), .A(n4337), .ZN(n4521) );
  NOR3_X1 U5436 ( .A1(n7883), .A2(n8108), .A3(n7902), .ZN(n7987) );
  AND2_X1 U5437 ( .A1(n7902), .A2(n8105), .ZN(n7875) );
  NOR2_X1 U5438 ( .A1(n7883), .A2(n7902), .ZN(n7898) );
  OR2_X1 U5439 ( .A1(n8855), .A2(n7897), .ZN(n7891) );
  AND2_X1 U5440 ( .A1(n6198), .A2(n6197), .ZN(n7895) );
  AND2_X1 U5441 ( .A1(n4734), .A2(n4733), .ZN(n7798) );
  NAND2_X1 U5442 ( .A1(n6186), .A2(n6180), .ZN(n4733) );
  AND2_X1 U5443 ( .A1(n6183), .A2(n6186), .ZN(n7664) );
  NAND2_X1 U5444 ( .A1(n4737), .A2(n4739), .ZN(n7516) );
  INV_X1 U5445 ( .A(n4740), .ZN(n4739) );
  NAND2_X1 U5446 ( .A1(n7502), .A2(n4742), .ZN(n4737) );
  NAND2_X1 U5447 ( .A1(n7714), .A2(n7708), .ZN(n7709) );
  AND3_X1 U5448 ( .A1(n8744), .A2(n4316), .A3(n4369), .ZN(n7720) );
  NAND2_X1 U5449 ( .A1(n4738), .A2(n6169), .ZN(n7715) );
  OR2_X1 U5450 ( .A1(n7502), .A2(n6121), .ZN(n4738) );
  NAND2_X1 U5451 ( .A1(n8744), .A2(n4316), .ZN(n7541) );
  AND2_X1 U5452 ( .A1(n8744), .A2(n9960), .ZN(n7542) );
  NAND2_X1 U5453 ( .A1(n6958), .A2(n7445), .ZN(n8736) );
  NOR2_X1 U5454 ( .A1(n8745), .A2(n8752), .ZN(n8744) );
  NAND2_X1 U5455 ( .A1(n6949), .A2(n6948), .ZN(n4517) );
  NOR2_X1 U5456 ( .A1(n8050), .A2(n9938), .ZN(n7350) );
  NAND2_X1 U5457 ( .A1(n8543), .A2(n4777), .ZN(n8528) );
  NAND2_X1 U5458 ( .A1(n8543), .A2(n6272), .ZN(n8525) );
  NAND2_X1 U5459 ( .A1(n5898), .A2(n5897), .ZN(n8832) );
  AND2_X1 U5460 ( .A1(n5809), .A2(n5808), .ZN(n9974) );
  INV_X1 U5461 ( .A(n9981), .ZN(n8857) );
  INV_X1 U5462 ( .A(n8856), .ZN(n9980) );
  NOR2_X1 U5463 ( .A1(n6939), .A2(n7950), .ZN(n9925) );
  OAI21_X2 U5464 ( .B1(n6103), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U5465 ( .A1(n5895), .A2(n5894), .ZN(n5911) );
  AND2_X1 U5466 ( .A1(n5658), .A2(n5657), .ZN(n5726) );
  NOR2_X1 U5467 ( .A1(n5058), .A2(n5057), .ZN(n5082) );
  OR2_X1 U5468 ( .A1(n5501), .A2(n5502), .ZN(n4462) );
  OR2_X1 U5469 ( .A1(n8948), .A2(n8949), .ZN(n8946) );
  OR2_X1 U5470 ( .A1(n4996), .A2(n4995), .ZN(n8972) );
  NAND2_X1 U5471 ( .A1(n5448), .A2(n5447), .ZN(n4811) );
  NAND2_X1 U5472 ( .A1(n4805), .A2(n4808), .ZN(n8993) );
  NOR2_X1 U5473 ( .A1(n5111), .A2(n8921), .ZN(n4399) );
  NAND2_X1 U5474 ( .A1(n5111), .A2(n8921), .ZN(n4401) );
  AND2_X1 U5475 ( .A1(n4956), .A2(n7023), .ZN(n6867) );
  AND2_X1 U5476 ( .A1(n4801), .A2(n8957), .ZN(n4800) );
  NAND2_X1 U5477 ( .A1(n8949), .A2(n5323), .ZN(n4801) );
  NAND2_X1 U5478 ( .A1(n4304), .A2(n4438), .ZN(n4435) );
  OAI21_X1 U5479 ( .B1(n6529), .B2(n6734), .A(n6525), .ZN(n4414) );
  OR2_X1 U5480 ( .A1(n6556), .A2(n6555), .ZN(n6558) );
  AND4_X1 U5481 ( .A1(n4961), .A2(n4960), .A3(n4959), .A4(n4958), .ZN(n7113)
         );
  AND4_X1 U5482 ( .A1(n4981), .A2(n4980), .A3(n4979), .A4(n4978), .ZN(n4993)
         );
  OR2_X1 U5483 ( .A1(n6688), .A2(n6588), .ZN(n4482) );
  NOR2_X1 U5484 ( .A1(n9820), .A2(n9819), .ZN(n9818) );
  NOR2_X1 U5485 ( .A1(n9818), .A2(n4489), .ZN(n9056) );
  AND2_X1 U5486 ( .A1(n9826), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4489) );
  NAND2_X1 U5487 ( .A1(n9056), .A2(n9057), .ZN(n9055) );
  AOI21_X1 U5488 ( .B1(n7465), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7464), .ZN(
        n7678) );
  NAND2_X1 U5489 ( .A1(n4655), .A2(n4654), .ZN(n9199) );
  AOI21_X1 U5490 ( .B1(n4656), .B2(n4657), .A(n6353), .ZN(n4654) );
  INV_X1 U5491 ( .A(n4658), .ZN(n4657) );
  OR2_X1 U5492 ( .A1(n4561), .A2(n4323), .ZN(n4557) );
  INV_X1 U5493 ( .A(n4560), .ZN(n4559) );
  NOR2_X1 U5494 ( .A1(n9295), .A2(n4666), .ZN(n9254) );
  NOR2_X1 U5495 ( .A1(n9295), .A2(n4668), .ZN(n9273) );
  NAND2_X1 U5496 ( .A1(n4634), .A2(n4632), .ZN(n4631) );
  NAND2_X1 U5497 ( .A1(n4319), .A2(n9346), .ZN(n4633) );
  OR2_X1 U5498 ( .A1(n9314), .A2(n9414), .ZN(n9295) );
  NOR2_X1 U5499 ( .A1(n5361), .A2(n5360), .ZN(n5386) );
  AND2_X1 U5500 ( .A1(n4591), .A2(n4588), .ZN(n9308) );
  INV_X1 U5501 ( .A(n4589), .ZN(n4588) );
  OAI21_X1 U5502 ( .B1(n4593), .B2(n4590), .A(n4336), .ZN(n4589) );
  AND2_X1 U5503 ( .A1(n8013), .A2(n4350), .ZN(n9323) );
  AND2_X1 U5504 ( .A1(n8013), .A2(n4311), .ZN(n9341) );
  NAND2_X1 U5505 ( .A1(n8013), .A2(n4675), .ZN(n9342) );
  AND2_X1 U5506 ( .A1(n5309), .A2(n5308), .ZN(n8950) );
  NAND2_X1 U5507 ( .A1(n9680), .A2(n7827), .ZN(n4645) );
  NAND2_X1 U5508 ( .A1(n8007), .A2(n8008), .ZN(n8006) );
  AND4_X1 U5509 ( .A1(n5265), .A2(n5264), .A3(n5263), .A4(n5262), .ZN(n9690)
         );
  AND2_X1 U5510 ( .A1(n9682), .A2(n7973), .ZN(n8013) );
  INV_X1 U5511 ( .A(n4551), .ZN(n4550) );
  OAI21_X1 U5512 ( .B1(n4552), .B2(n4305), .A(n7819), .ZN(n4551) );
  NOR2_X1 U5513 ( .A1(n4828), .A2(n9697), .ZN(n9682) );
  OAI211_X1 U5514 ( .C1(n7330), .C2(n4599), .A(n4598), .B(n7476), .ZN(n7744)
         );
  INV_X1 U5515 ( .A(n4600), .ZN(n4599) );
  NAND2_X1 U5516 ( .A1(n4602), .A2(n4600), .ZN(n4598) );
  AND2_X1 U5517 ( .A1(n4306), .A2(n4671), .ZN(n4670) );
  AOI21_X1 U5518 ( .B1(n4653), .B2(n7478), .A(n4652), .ZN(n4651) );
  INV_X1 U5519 ( .A(n7480), .ZN(n4652) );
  NAND2_X1 U5520 ( .A1(n7228), .A2(n4306), .ZN(n8071) );
  NAND2_X1 U5521 ( .A1(n7228), .A2(n4673), .ZN(n7339) );
  AND4_X1 U5522 ( .A1(n5088), .A2(n5087), .A3(n5086), .A4(n5085), .ZN(n8076)
         );
  AND2_X1 U5523 ( .A1(n7225), .A2(n7124), .ZN(n7126) );
  AND2_X1 U5524 ( .A1(n7124), .A2(n7123), .ZN(n7125) );
  AND2_X1 U5525 ( .A1(n7228), .A2(n7230), .ZN(n7229) );
  AND4_X1 U5526 ( .A1(n5008), .A2(n5007), .A3(n5006), .A4(n5005), .ZN(n7220)
         );
  INV_X1 U5527 ( .A(n7267), .ZN(n7264) );
  AND2_X1 U5528 ( .A1(n6921), .A2(n7214), .ZN(n7265) );
  AND2_X1 U5529 ( .A1(n6915), .A2(n6883), .ZN(n6884) );
  NOR2_X1 U5530 ( .A1(n6325), .A2(n7238), .ZN(n6917) );
  AND2_X1 U5531 ( .A1(n6325), .A2(n6885), .ZN(n4540) );
  AND2_X1 U5532 ( .A1(n6920), .A2(n7238), .ZN(n6921) );
  NAND2_X1 U5533 ( .A1(n6316), .A2(n6315), .ZN(n9360) );
  AND2_X1 U5534 ( .A1(n4664), .A2(n4663), .ZN(n9376) );
  AOI22_X1 U5535 ( .A1(n9188), .A2(n9349), .B1(n9347), .B2(n9211), .ZN(n4663)
         );
  NAND2_X1 U5536 ( .A1(n9189), .A2(n9352), .ZN(n4664) );
  XNOR2_X1 U5537 ( .A(n6095), .B(n6094), .ZN(n8884) );
  XNOR2_X1 U5538 ( .A(n6087), .B(SI_30_), .ZN(n8888) );
  XNOR2_X1 U5539 ( .A(n6067), .B(n6066), .ZN(n8021) );
  AND2_X1 U5540 ( .A1(n6049), .A2(n6048), .ZN(n6067) );
  XNOR2_X1 U5541 ( .A(n5583), .B(n5582), .ZN(n8000) );
  NAND2_X1 U5542 ( .A1(n6047), .A2(n6045), .ZN(n5583) );
  OR2_X1 U5543 ( .A1(n4901), .A2(n4845), .ZN(n4902) );
  NAND2_X1 U5544 ( .A1(n5354), .A2(n5372), .ZN(n5355) );
  NOR2_X1 U5545 ( .A1(n5253), .A2(n4877), .ZN(n5306) );
  NAND2_X1 U5546 ( .A1(n5205), .A2(n4837), .ZN(n4857) );
  NAND2_X1 U5547 ( .A1(n4606), .A2(n4611), .ZN(n5250) );
  NAND2_X1 U5548 ( .A1(n5198), .A2(n4613), .ZN(n4606) );
  AND2_X1 U5549 ( .A1(n5018), .A2(n4836), .ZN(n5205) );
  OR2_X1 U5550 ( .A1(n5100), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5121) );
  AND2_X1 U5551 ( .A1(n4427), .A2(n4426), .ZN(n5091) );
  NAND2_X1 U5552 ( .A1(n4505), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4985) );
  INV_X1 U5553 ( .A(n4945), .ZN(n4505) );
  XNOR2_X1 U5554 ( .A(n4940), .B(n4919), .ZN(n4939) );
  NAND2_X1 U5555 ( .A1(n6021), .A2(n6020), .ZN(n8776) );
  INV_X1 U5556 ( .A(n8461), .ZN(n8273) );
  NAND2_X1 U5557 ( .A1(n4732), .A2(n4731), .ZN(n8093) );
  OAI21_X1 U5558 ( .B1(n7072), .B2(n7071), .A(n7070), .ZN(n7151) );
  NAND2_X1 U5559 ( .A1(n4702), .A2(n4707), .ZN(n8227) );
  NAND2_X1 U5560 ( .A1(n8279), .A2(n4705), .ZN(n4702) );
  AND2_X1 U5561 ( .A1(n7017), .A2(n7016), .ZN(n8053) );
  INV_X1 U5562 ( .A(n8354), .ZN(n7994) );
  INV_X1 U5563 ( .A(n8163), .ZN(n8258) );
  NAND2_X1 U5564 ( .A1(n7939), .A2(n6071), .ZN(n5999) );
  INV_X1 U5565 ( .A(n7415), .ZN(n9960) );
  NAND2_X1 U5566 ( .A1(n8058), .A2(n9938), .ZN(n7346) );
  AND2_X1 U5567 ( .A1(n7004), .A2(n6998), .ZN(n8282) );
  NAND2_X1 U5568 ( .A1(n4708), .A2(n8130), .ZN(n8320) );
  OR2_X1 U5569 ( .A1(n8279), .A2(n8278), .ZN(n4708) );
  AOI21_X1 U5570 ( .B1(n7372), .B2(n7371), .A(n4816), .ZN(n7373) );
  INV_X1 U5571 ( .A(n8240), .ZN(n8342) );
  NAND2_X1 U5572 ( .A1(n4714), .A2(n4718), .ZN(n8328) );
  NAND2_X1 U5573 ( .A1(n8163), .A2(n4720), .ZN(n4714) );
  INV_X1 U5574 ( .A(n8349), .ZN(n8325) );
  AND2_X1 U5575 ( .A1(n6024), .A2(n6013), .ZN(n8551) );
  INV_X1 U5576 ( .A(n8336), .ZN(n8346) );
  OR2_X1 U5577 ( .A1(n7061), .A2(n6571), .ZN(n8353) );
  NAND4_X1 U5578 ( .A1(n5787), .A2(n5786), .A3(n5785), .A4(n5784), .ZN(n8359)
         );
  OR2_X1 U5579 ( .A1(n5754), .A2(n5783), .ZN(n5784) );
  OR2_X1 U5580 ( .A1(n4302), .A2(n5782), .ZN(n5785) );
  OR2_X1 U5581 ( .A1(n5754), .A2(n5767), .ZN(n5770) );
  NAND4_X1 U5582 ( .A1(n5739), .A2(n5738), .A3(n5737), .A4(n5736), .ZN(n8362)
         );
  NAND4_X1 U5583 ( .A1(n5724), .A2(n5723), .A3(n5722), .A4(n5721), .ZN(n7077)
         );
  OR2_X1 U5584 ( .A1(n4302), .A2(n5720), .ZN(n5722) );
  OR2_X1 U5585 ( .A1(n5754), .A2(n8743), .ZN(n5721) );
  INV_X1 U5586 ( .A(n6958), .ZN(n8363) );
  XNOR2_X1 U5587 ( .A(n5701), .B(P2_IR_REG_1__SCAN_IN), .ZN(n7047) );
  INV_X1 U5588 ( .A(n4471), .ZN(n6830) );
  INV_X1 U5589 ( .A(n4469), .ZN(n6856) );
  INV_X1 U5590 ( .A(n4475), .ZN(n6901) );
  AND2_X1 U5591 ( .A1(n4475), .A2(n4474), .ZN(n6904) );
  NAND2_X1 U5592 ( .A1(n6906), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4474) );
  INV_X1 U5593 ( .A(n4473), .ZN(n7173) );
  AND2_X1 U5594 ( .A1(n4473), .A2(n4472), .ZN(n7176) );
  NAND2_X1 U5595 ( .A1(n7178), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4472) );
  AND2_X1 U5596 ( .A1(n5878), .A2(n5864), .ZN(n7955) );
  XNOR2_X1 U5597 ( .A(n4476), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U5598 ( .A1(n8430), .A2(n4477), .ZN(n4476) );
  OR2_X1 U5599 ( .A1(n8432), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4477) );
  AOI21_X1 U5600 ( .B1(n8512), .B2(n8519), .A(n8518), .ZN(n8773) );
  INV_X1 U5601 ( .A(n8770), .ZN(n8511) );
  NAND2_X1 U5602 ( .A1(n6011), .A2(n6010), .ZN(n8784) );
  NAND2_X1 U5603 ( .A1(n7942), .A2(n6071), .ZN(n6011) );
  AND2_X1 U5604 ( .A1(n5941), .A2(n6105), .ZN(n8554) );
  AND2_X1 U5605 ( .A1(n8597), .A2(n6261), .ZN(n8578) );
  NAND2_X1 U5606 ( .A1(n4507), .A2(n4512), .ZN(n8604) );
  OR2_X1 U5607 ( .A1(n8637), .A2(n4513), .ZN(n4507) );
  INV_X1 U5608 ( .A(n4753), .ZN(n8629) );
  OAI21_X1 U5609 ( .B1(n8657), .B2(n4762), .A(n4759), .ZN(n4753) );
  AND2_X1 U5610 ( .A1(n4515), .A2(n4516), .ZN(n8623) );
  NAND2_X1 U5611 ( .A1(n8637), .A2(n8643), .ZN(n4515) );
  AND2_X1 U5612 ( .A1(n4763), .A2(n4761), .ZN(n8642) );
  NAND2_X1 U5613 ( .A1(n4524), .A2(n4522), .ZN(n7986) );
  NAND2_X1 U5614 ( .A1(n4524), .A2(n7872), .ZN(n7873) );
  OR2_X1 U5615 ( .A1(n7543), .A2(n9981), .ZN(n8530) );
  NAND2_X2 U5616 ( .A1(n5791), .A2(n5790), .ZN(n8239) );
  NAND2_X1 U5617 ( .A1(n8749), .A2(n7412), .ZN(n7497) );
  INV_X1 U5618 ( .A(n8553), .ZN(n8746) );
  OAI211_X1 U5619 ( .C1(n5773), .C2(n6631), .A(n5709), .B(n5708), .ZN(n7311)
         );
  OR2_X1 U5620 ( .A1(n9926), .A2(n7296), .ZN(n8553) );
  INV_X1 U5621 ( .A(n8721), .ZN(n8753) );
  INV_X1 U5622 ( .A(n8530), .ZN(n8748) );
  OR2_X1 U5623 ( .A1(n8765), .A2(n9981), .ZN(n4506) );
  AND2_X1 U5624 ( .A1(n7057), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9937) );
  XNOR2_X1 U5625 ( .A(n6085), .B(n5667), .ZN(n7493) );
  INV_X1 U5626 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6106) );
  INV_X1 U5627 ( .A(n8554), .ZN(n8440) );
  INV_X1 U5628 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6637) );
  INV_X1 U5629 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6620) );
  AND2_X1 U5630 ( .A1(n4402), .A2(n7245), .ZN(n4403) );
  NAND2_X1 U5631 ( .A1(n8974), .A2(n4405), .ZN(n4404) );
  AND4_X1 U5632 ( .A1(n5595), .A2(n5594), .A3(n5593), .A4(n5592), .ZN(n9197)
         );
  AND2_X1 U5633 ( .A1(n4456), .A2(n4355), .ZN(n4452) );
  AOI21_X1 U5634 ( .B1(n4457), .B2(n4459), .A(n4364), .ZN(n4456) );
  NAND2_X1 U5635 ( .A1(n5562), .A2(n5561), .ZN(n9379) );
  NAND2_X1 U5636 ( .A1(n7528), .A2(n5146), .ZN(n8061) );
  AOI21_X1 U5637 ( .B1(n9007), .B2(n4443), .A(n4445), .ZN(n4442) );
  INV_X1 U5638 ( .A(n4447), .ZN(n4443) );
  NAND2_X1 U5639 ( .A1(n9029), .A2(n4812), .ZN(n5632) );
  NOR2_X1 U5640 ( .A1(n5574), .A2(n4364), .ZN(n4812) );
  NAND2_X1 U5641 ( .A1(n4802), .A2(n6865), .ZN(n6756) );
  INV_X1 U5642 ( .A(n8986), .ZN(n4408) );
  NAND2_X1 U5643 ( .A1(n8946), .A2(n5323), .ZN(n8958) );
  NAND2_X1 U5644 ( .A1(n4975), .A2(n4974), .ZN(n8978) );
  AND2_X1 U5645 ( .A1(n4965), .A2(n4964), .ZN(n4975) );
  NAND2_X1 U5646 ( .A1(n5009), .A2(n5725), .ZN(n4974) );
  NAND2_X1 U5647 ( .A1(n8919), .A2(n8921), .ZN(n5112) );
  INV_X1 U5648 ( .A(n4439), .ZN(n8985) );
  NAND2_X1 U5649 ( .A1(n4792), .A2(n5224), .ZN(n7909) );
  NAND2_X1 U5650 ( .A1(n4811), .A2(n5467), .ZN(n8996) );
  NAND2_X1 U5651 ( .A1(n5460), .A2(n5459), .ZN(n9404) );
  INV_X1 U5652 ( .A(n6757), .ZN(n4933) );
  NAND2_X1 U5653 ( .A1(n4460), .A2(n4459), .ZN(n9029) );
  NAND2_X1 U5654 ( .A1(n5539), .A2(n5538), .ZN(n9383) );
  NAND2_X1 U5655 ( .A1(n7942), .A2(n5009), .ZN(n5539) );
  INV_X1 U5656 ( .A(n7336), .ZN(n9049) );
  INV_X1 U5657 ( .A(n7322), .ZN(n9050) );
  INV_X1 U5658 ( .A(n7220), .ZN(n9051) );
  AND2_X1 U5659 ( .A1(n9785), .A2(n9784), .ZN(n9787) );
  INV_X1 U5660 ( .A(n4482), .ZN(n9801) );
  NOR2_X1 U5661 ( .A1(n4482), .A2(n4481), .ZN(n9808) );
  NAND2_X1 U5662 ( .A1(n9055), .A2(n4488), .ZN(n6985) );
  OR2_X1 U5663 ( .A1(n6982), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4488) );
  XNOR2_X1 U5664 ( .A(n7678), .B(n7677), .ZN(n7467) );
  NOR2_X1 U5665 ( .A1(n7924), .A2(n7923), .ZN(n7927) );
  OR2_X1 U5666 ( .A1(n9376), .A2(n9309), .ZN(n4662) );
  AND2_X1 U5667 ( .A1(n4579), .A2(n4577), .ZN(n9180) );
  INV_X1 U5668 ( .A(n4580), .ZN(n4577) );
  NAND2_X1 U5669 ( .A1(n4581), .A2(n4584), .ZN(n9191) );
  NAND2_X1 U5670 ( .A1(n9241), .A2(n9155), .ZN(n9226) );
  NAND2_X1 U5671 ( .A1(n4558), .A2(n4562), .ZN(n9253) );
  NAND2_X1 U5672 ( .A1(n9279), .A2(n4563), .ZN(n4558) );
  INV_X1 U5673 ( .A(n9404), .ZN(n9268) );
  NAND2_X1 U5674 ( .A1(n9279), .A2(n9281), .ZN(n4565) );
  NAND2_X1 U5675 ( .A1(n4636), .A2(n9148), .ZN(n9301) );
  NAND2_X1 U5676 ( .A1(n4637), .A2(n4641), .ZN(n4636) );
  INV_X1 U5677 ( .A(n9414), .ZN(n9299) );
  NAND2_X1 U5678 ( .A1(n4641), .A2(n4639), .ZN(n9311) );
  NAND2_X1 U5679 ( .A1(n5385), .A2(n5384), .ZN(n9419) );
  NAND2_X1 U5680 ( .A1(n4587), .A2(n4593), .ZN(n9322) );
  OR2_X1 U5681 ( .A1(n7979), .A2(n4594), .ZN(n4587) );
  AND2_X1 U5682 ( .A1(n4597), .A2(n4596), .ZN(n9340) );
  NAND2_X1 U5683 ( .A1(n4648), .A2(n7827), .ZN(n7828) );
  NAND2_X1 U5684 ( .A1(n4553), .A2(n4552), .ZN(n9681) );
  NAND2_X1 U5685 ( .A1(n7749), .A2(n4554), .ZN(n4553) );
  NAND2_X1 U5686 ( .A1(n7749), .A2(n7748), .ZN(n7818) );
  NAND2_X1 U5687 ( .A1(n5208), .A2(n5207), .ZN(n7816) );
  NAND2_X1 U5688 ( .A1(n5156), .A2(n5155), .ZN(n9671) );
  NAND2_X1 U5689 ( .A1(n7475), .A2(n7474), .ZN(n8068) );
  NAND2_X1 U5690 ( .A1(n7333), .A2(n7332), .ZN(n7479) );
  AND2_X1 U5691 ( .A1(n9725), .A2(n7200), .ZN(n9706) );
  INV_X1 U5692 ( .A(n9911), .ZN(n9909) );
  AND2_X1 U5693 ( .A1(n9370), .A2(n9369), .ZN(n9371) );
  OAI22_X1 U5694 ( .A1(n5122), .A2(n4544), .B1(P1_IR_REG_31__SCAN_IN), .B2(
        P1_IR_REG_30__SCAN_IN), .ZN(n4543) );
  XNOR2_X1 U5695 ( .A(n4409), .B(P1_IR_REG_26__SCAN_IN), .ZN(n7943) );
  NAND2_X1 U5696 ( .A1(n4866), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4409) );
  MUX2_X1 U5697 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4865), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n4867) );
  NAND2_X1 U5698 ( .A1(n4690), .A2(n5040), .ZN(n5065) );
  NAND2_X1 U5699 ( .A1(n5037), .A2(n5036), .ZN(n4690) );
  INV_X1 U5700 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6626) );
  AND2_X1 U5701 ( .A1(n5020), .A2(n5019), .ZN(n9783) );
  NAND2_X1 U5702 ( .A1(n4689), .A2(n4970), .ZN(n4983) );
  NAND2_X1 U5703 ( .A1(n4380), .A2(n7702), .ZN(n4680) );
  AND2_X1 U5704 ( .A1(n4449), .A2(n4308), .ZN(n7696) );
  NAND2_X1 U5705 ( .A1(n4411), .A2(n6564), .ZN(n6569) );
  OAI21_X1 U5706 ( .B1(n9111), .B2(n9110), .A(n4497), .ZN(P1_U3260) );
  AOI21_X1 U5707 ( .B1(n4499), .B2(n9110), .A(n4498), .ZN(n4497) );
  OAI21_X1 U5708 ( .B1(n9773), .B2(n4696), .A(n9112), .ZN(n4498) );
  NAND2_X1 U5709 ( .A1(n4665), .A2(n4660), .ZN(P1_U3263) );
  OR2_X1 U5710 ( .A1(n9377), .A2(n9356), .ZN(n4665) );
  AND2_X1 U5711 ( .A1(n4662), .A2(n4661), .ZN(n4660) );
  AOI21_X1 U5712 ( .B1(n9374), .B2(n9706), .A(n9190), .ZN(n4661) );
  NAND2_X1 U5713 ( .A1(n6112), .A2(n6237), .ZN(n4762) );
  INV_X1 U5714 ( .A(n7406), .ZN(n7009) );
  NAND2_X1 U5715 ( .A1(n6574), .A2(n4299), .ZN(n4991) );
  INV_X2 U5716 ( .A(n4991), .ZN(n5009) );
  AND2_X1 U5717 ( .A1(n4437), .A2(n8042), .ZN(n4304) );
  NAND2_X1 U5718 ( .A1(n4320), .A2(n5003), .ZN(n4794) );
  AND2_X1 U5719 ( .A1(n9697), .A2(n9043), .ZN(n4305) );
  NAND2_X1 U5720 ( .A1(n6199), .A2(n7872), .ZN(n4523) );
  INV_X1 U5721 ( .A(n4762), .ZN(n4761) );
  INV_X2 U5722 ( .A(n4301), .ZN(n5695) );
  AND2_X1 U5723 ( .A1(n4673), .A2(n4672), .ZN(n4306) );
  AND2_X1 U5724 ( .A1(n6457), .A2(n6517), .ZN(n4307) );
  AND2_X1 U5725 ( .A1(n4379), .A2(n4795), .ZN(n4308) );
  AND2_X1 U5726 ( .A1(n4340), .A2(n4536), .ZN(n4309) );
  AND2_X1 U5727 ( .A1(n8996), .A2(n8994), .ZN(n4310) );
  INV_X1 U5728 ( .A(n7243), .ZN(n7328) );
  INV_X1 U5729 ( .A(n6112), .ZN(n8643) );
  AND2_X1 U5730 ( .A1(n6241), .A2(n6246), .ZN(n6112) );
  AND2_X1 U5731 ( .A1(n5285), .A2(n5284), .ZN(n8016) );
  INV_X1 U5732 ( .A(n8016), .ZN(n9439) );
  NAND2_X1 U5733 ( .A1(n5999), .A2(n5998), .ZN(n8788) );
  AND2_X1 U5734 ( .A1(n8812), .A2(n8631), .ZN(n8474) );
  AND2_X1 U5735 ( .A1(n4675), .A2(n4674), .ZN(n4311) );
  INV_X1 U5736 ( .A(n4759), .ZN(n4758) );
  AOI21_X1 U5737 ( .B1(n4761), .B2(n4760), .A(n6236), .ZN(n4759) );
  NOR2_X1 U5738 ( .A1(n4674), .A2(n9121), .ZN(n4312) );
  AND2_X1 U5739 ( .A1(n6283), .A2(n6086), .ZN(n4313) );
  AND2_X1 U5740 ( .A1(n4744), .A2(n6314), .ZN(n4314) );
  OR2_X1 U5741 ( .A1(n9445), .A2(n9690), .ZN(n7969) );
  AND2_X1 U5742 ( .A1(n4435), .A2(n5293), .ZN(n4315) );
  AND2_X1 U5743 ( .A1(n9965), .A2(n9960), .ZN(n4316) );
  NAND2_X1 U5744 ( .A1(n4798), .A2(n5145), .ZN(n7528) );
  AND2_X2 U5745 ( .A1(n4852), .A2(n9651), .ZN(n5084) );
  NAND4_X1 U5746 ( .A1(n4856), .A2(n4855), .A3(n4854), .A4(n4853), .ZN(n6325)
         );
  INV_X2 U5747 ( .A(n6574), .ZN(n4988) );
  NOR2_X1 U5748 ( .A1(n5673), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n5676) );
  NOR2_X1 U5749 ( .A1(n5016), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5018) );
  NAND2_X1 U5750 ( .A1(n7655), .A2(n7665), .ZN(n6177) );
  INV_X1 U5751 ( .A(n5269), .ZN(n4438) );
  NAND2_X1 U5752 ( .A1(n8597), .A2(n4785), .ZN(n8565) );
  OR2_X1 U5753 ( .A1(n8842), .A2(n8727), .ZN(n5877) );
  INV_X1 U5754 ( .A(n6616), .ZN(n4916) );
  AND2_X1 U5755 ( .A1(n4444), .A2(n8914), .ZN(n4317) );
  AND2_X1 U5756 ( .A1(n9404), .A2(n9286), .ZN(n4318) );
  AND2_X1 U5757 ( .A1(n5774), .A2(n5660), .ZN(n5788) );
  AND2_X1 U5758 ( .A1(n4634), .A2(n4642), .ZN(n4319) );
  NAND2_X1 U5759 ( .A1(n5052), .A2(n7320), .ZN(n4320) );
  XNOR2_X1 U5760 ( .A(n8776), .B(n8516), .ZN(n8524) );
  INV_X1 U5761 ( .A(n8524), .ZN(n4779) );
  AND2_X1 U5762 ( .A1(n7908), .A2(n4438), .ZN(n4321) );
  INV_X1 U5763 ( .A(n8058), .ZN(n6945) );
  INV_X1 U5764 ( .A(n4719), .ZN(n4718) );
  NOR2_X1 U5765 ( .A1(n8256), .A2(n8255), .ZN(n4719) );
  INV_X1 U5766 ( .A(n7332), .ZN(n4653) );
  AND4_X1 U5767 ( .A1(n5713), .A2(n5712), .A3(n5711), .A4(n5710), .ZN(n6958)
         );
  NAND2_X1 U5768 ( .A1(n5334), .A2(n5333), .ZN(n9428) );
  INV_X1 U5769 ( .A(n9428), .ZN(n4674) );
  NAND2_X1 U5770 ( .A1(n9158), .A2(n6506), .ZN(n9200) );
  AND2_X1 U5771 ( .A1(n8265), .A2(n8117), .ZN(n4322) );
  NAND2_X1 U5772 ( .A1(n9651), .A2(n8024), .ZN(n5210) );
  INV_X2 U5773 ( .A(n5210), .ZN(n5591) );
  NAND2_X1 U5774 ( .A1(n8613), .A2(n5989), .ZN(n8597) );
  INV_X1 U5775 ( .A(n8656), .ZN(n4760) );
  NAND3_X1 U5776 ( .A1(n4945), .A2(n4789), .A3(n4832), .ZN(n5016) );
  AND2_X1 U5777 ( .A1(n9399), .A2(n9271), .ZN(n4323) );
  AND3_X1 U5778 ( .A1(n4843), .A2(n4860), .A3(n4842), .ZN(n4324) );
  AND2_X1 U5779 ( .A1(n4705), .A2(n8226), .ZN(n4325) );
  NAND2_X1 U5780 ( .A1(n5991), .A2(n5990), .ZN(n8792) );
  INV_X1 U5781 ( .A(n8792), .ZN(n4486) );
  NAND2_X1 U5782 ( .A1(n4789), .A2(n4945), .ZN(n4962) );
  AND2_X1 U5783 ( .A1(n8148), .A2(n8147), .ZN(n4326) );
  XOR2_X1 U5784 ( .A(n8492), .B(n8491), .Z(n4327) );
  AND2_X1 U5785 ( .A1(n8950), .A2(n9348), .ZN(n6458) );
  INV_X1 U5786 ( .A(n9023), .ZN(n7230) );
  NOR2_X1 U5787 ( .A1(n8627), .A2(n8645), .ZN(n4328) );
  AND3_X1 U5788 ( .A1(n6286), .A2(n6284), .A3(n6285), .ZN(n4329) );
  NAND2_X1 U5789 ( .A1(n5067), .A2(SI_6_), .ZN(n4330) );
  NAND2_X1 U5790 ( .A1(n6509), .A2(n9160), .ZN(n9179) );
  NAND2_X1 U5791 ( .A1(n7644), .A2(n7626), .ZN(n4331) );
  AND2_X1 U5792 ( .A1(n6524), .A2(n6523), .ZN(n4332) );
  AND2_X1 U5793 ( .A1(n6516), .A2(n4428), .ZN(n4333) );
  INV_X1 U5794 ( .A(n7817), .ZN(n4556) );
  AND2_X1 U5795 ( .A1(n8627), .A2(n8645), .ZN(n4334) );
  AND2_X1 U5796 ( .A1(n7498), .A2(n9960), .ZN(n4335) );
  INV_X1 U5797 ( .A(n5040), .ZN(n4692) );
  NAND2_X1 U5798 ( .A1(n9423), .A2(n9350), .ZN(n4336) );
  INV_X1 U5799 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4679) );
  INV_X1 U5800 ( .A(n4485), .ZN(n4484) );
  NAND2_X1 U5801 ( .A1(n4487), .A2(n4486), .ZN(n4485) );
  OR2_X1 U5802 ( .A1(n8848), .A2(n7994), .ZN(n4337) );
  NAND3_X1 U5803 ( .A1(n4844), .A2(n4836), .A3(n4573), .ZN(n4338) );
  INV_X1 U5804 ( .A(n4595), .ZN(n4594) );
  AOI21_X1 U5805 ( .B1(n9142), .B2(n4596), .A(n9122), .ZN(n4595) );
  OR2_X1 U5806 ( .A1(n4811), .A2(n5467), .ZN(n4339) );
  INV_X1 U5807 ( .A(n4514), .ZN(n4513) );
  NOR2_X1 U5808 ( .A1(n4328), .A2(n8474), .ZN(n4514) );
  AND2_X1 U5809 ( .A1(n6202), .A2(n6201), .ZN(n7876) );
  AND4_X1 U5810 ( .A1(n5707), .A2(n5706), .A3(n5705), .A4(n5704), .ZN(n7406)
         );
  AND2_X1 U5811 ( .A1(n4788), .A2(n4534), .ZN(n4340) );
  INV_X1 U5812 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5122) );
  INV_X1 U5813 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4875) );
  AND2_X1 U5814 ( .A1(n5479), .A2(n5478), .ZN(n9258) );
  INV_X1 U5815 ( .A(n9258), .ZN(n9399) );
  OR2_X1 U5816 ( .A1(n9129), .A2(n4318), .ZN(n4341) );
  NAND2_X1 U5817 ( .A1(n4420), .A2(n4422), .ZN(n4342) );
  AND2_X1 U5818 ( .A1(n4565), .A2(n4564), .ZN(n4343) );
  AND2_X1 U5819 ( .A1(n4846), .A2(P1_IR_REG_30__SCAN_IN), .ZN(n4344) );
  NOR2_X1 U5820 ( .A1(n8768), .A2(n8767), .ZN(n4345) );
  AND2_X1 U5821 ( .A1(n9383), .A2(n9203), .ZN(n9138) );
  AND2_X1 U5822 ( .A1(n6177), .A2(n6186), .ZN(n4346) );
  AND2_X1 U5823 ( .A1(n8459), .A2(n6203), .ZN(n4347) );
  NAND2_X1 U5824 ( .A1(n9886), .A2(n9047), .ZN(n4348) );
  AND2_X1 U5825 ( .A1(n4583), .A2(n9200), .ZN(n4349) );
  AND2_X1 U5826 ( .A1(n9328), .A2(n4311), .ZN(n4350) );
  OR2_X1 U5827 ( .A1(n4769), .A2(n4313), .ZN(n4351) );
  AND2_X1 U5828 ( .A1(n6530), .A2(n7453), .ZN(n4352) );
  AND2_X1 U5829 ( .A1(n9196), .A2(n9139), .ZN(n4353) );
  AND2_X1 U5830 ( .A1(n4460), .A2(n4461), .ZN(n4354) );
  OR2_X1 U5831 ( .A1(n8770), .A2(n8488), .ZN(n6278) );
  OR2_X1 U5832 ( .A1(n4458), .A2(n4453), .ZN(n4355) );
  AND2_X1 U5833 ( .A1(n4535), .A2(n5672), .ZN(n4356) );
  OR2_X1 U5834 ( .A1(n4304), .A2(n4321), .ZN(n4357) );
  INV_X1 U5835 ( .A(n4523), .ZN(n4522) );
  INV_X1 U5836 ( .A(n4778), .ZN(n4777) );
  NAND2_X1 U5837 ( .A1(n4779), .A2(n6272), .ZN(n4778) );
  NAND2_X1 U5838 ( .A1(n4973), .A2(SI_3_), .ZN(n4358) );
  INV_X1 U5839 ( .A(n6108), .ZN(n8174) );
  XOR2_X1 U5840 ( .A(n8797), .B(n8175), .Z(n4359) );
  AND2_X1 U5841 ( .A1(n4725), .A2(n4726), .ZN(n4360) );
  AND2_X1 U5842 ( .A1(n8013), .A2(n8016), .ZN(n4361) );
  NAND2_X1 U5843 ( .A1(n6073), .A2(n6072), .ZN(n8454) );
  INV_X1 U5844 ( .A(n8454), .ZN(n4773) );
  INV_X1 U5845 ( .A(n8108), .ZN(n8848) );
  OR2_X1 U5846 ( .A1(n7979), .A2(n9142), .ZN(n4597) );
  INV_X1 U5847 ( .A(n4442), .ZN(n8913) );
  AND4_X1 U5848 ( .A1(n5241), .A2(n5240), .A3(n5239), .A4(n5238), .ZN(n8040)
         );
  NAND2_X1 U5849 ( .A1(n5895), .A2(n4676), .ZN(n4362) );
  OR2_X1 U5850 ( .A1(n8792), .A2(n8480), .ZN(n8566) );
  INV_X1 U5851 ( .A(n8566), .ZN(n4782) );
  INV_X1 U5852 ( .A(n4501), .ZN(n8652) );
  NOR3_X1 U5853 ( .A1(n8700), .A2(n8824), .A3(n4504), .ZN(n4501) );
  INV_X1 U5854 ( .A(n4503), .ZN(n8664) );
  NOR3_X1 U5855 ( .A1(n8700), .A2(n8824), .A3(n8828), .ZN(n4503) );
  NAND2_X1 U5856 ( .A1(n4763), .A2(n6237), .ZN(n4363) );
  AND2_X1 U5857 ( .A1(n5551), .A2(n5550), .ZN(n4364) );
  INV_X1 U5858 ( .A(n4625), .ZN(n4624) );
  NOR2_X1 U5859 ( .A1(n5531), .A2(n4626), .ZN(n4625) );
  NAND2_X1 U5860 ( .A1(n8605), .A2(n4484), .ZN(n4365) );
  AND3_X1 U5861 ( .A1(n5997), .A2(n5996), .A3(n5995), .ZN(n8480) );
  INV_X1 U5862 ( .A(n8480), .ZN(n4539) );
  INV_X1 U5863 ( .A(n9120), .ZN(n4596) );
  AND2_X1 U5864 ( .A1(n9119), .A2(n9348), .ZN(n9120) );
  INV_X1 U5865 ( .A(n9729), .ZN(n9697) );
  AND2_X1 U5866 ( .A1(n5234), .A2(n5233), .ZN(n9729) );
  INV_X1 U5867 ( .A(n4669), .ZN(n9288) );
  NOR2_X1 U5868 ( .A1(n9295), .A2(n9409), .ZN(n4669) );
  AND2_X1 U5869 ( .A1(n4732), .A2(n4730), .ZN(n4366) );
  AND2_X1 U5870 ( .A1(n5493), .A2(n5492), .ZN(n9240) );
  AND2_X1 U5871 ( .A1(n5258), .A2(n5257), .ZN(n7973) );
  INV_X1 U5872 ( .A(n7973), .ZN(n9445) );
  AND2_X1 U5873 ( .A1(n4648), .A2(n4646), .ZN(n4367) );
  AND2_X1 U5874 ( .A1(n4750), .A2(n5877), .ZN(n4368) );
  AND2_X1 U5875 ( .A1(n7604), .A2(n9969), .ZN(n4369) );
  INV_X1 U5876 ( .A(n9136), .ZN(n4586) );
  NOR2_X1 U5877 ( .A1(n9389), .A2(n9244), .ZN(n9136) );
  INV_X1 U5878 ( .A(n8474), .ZN(n4516) );
  NAND2_X1 U5879 ( .A1(n6867), .A2(n4433), .ZN(n6868) );
  NAND2_X1 U5880 ( .A1(n6396), .A2(n6395), .ZN(n6531) );
  NAND2_X1 U5881 ( .A1(n5837), .A2(n5836), .ZN(n7902) );
  INV_X1 U5882 ( .A(n7902), .ZN(n4495) );
  AND2_X1 U5883 ( .A1(n8974), .A2(n5003), .ZN(n7317) );
  AND3_X1 U5884 ( .A1(n8744), .A2(n4316), .A3(n7604), .ZN(n4370) );
  AND2_X1 U5885 ( .A1(n4406), .A2(n5055), .ZN(n4371) );
  INV_X1 U5886 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4396) );
  NAND2_X1 U5887 ( .A1(n4519), .A2(n4520), .ZN(n8460) );
  NAND2_X1 U5888 ( .A1(n5882), .A2(n5881), .ZN(n8837) );
  NAND2_X1 U5889 ( .A1(n7139), .A2(n7138), .ZN(n7333) );
  NAND2_X1 U5890 ( .A1(n5788), .A2(n4788), .ZN(n6307) );
  NAND2_X1 U5891 ( .A1(n5788), .A2(n4786), .ZN(n4372) );
  NOR2_X1 U5892 ( .A1(n7278), .A2(n7279), .ZN(n4373) );
  INV_X1 U5893 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6104) );
  INV_X1 U5894 ( .A(n4450), .ZN(n4798) );
  NAND2_X1 U5895 ( .A1(n5112), .A2(n8920), .ZN(n4450) );
  NOR2_X1 U5896 ( .A1(n7714), .A2(n4743), .ZN(n4742) );
  NOR2_X1 U5897 ( .A1(n7883), .A2(n4492), .ZN(n4490) );
  NAND2_X1 U5898 ( .A1(n8090), .A2(n8087), .ZN(n4374) );
  INV_X1 U5899 ( .A(n4496), .ZN(n8718) );
  NOR2_X1 U5900 ( .A1(n7883), .A2(n4491), .ZN(n4496) );
  AND3_X1 U5901 ( .A1(n4736), .A2(n4735), .A3(n6177), .ZN(n4375) );
  AND2_X1 U5902 ( .A1(n7330), .A2(n7329), .ZN(n4376) );
  AND2_X1 U5903 ( .A1(n6066), .A2(n6048), .ZN(n4377) );
  NAND2_X1 U5904 ( .A1(n4786), .A2(n4536), .ZN(n6305) );
  INV_X1 U5905 ( .A(n4794), .ZN(n4793) );
  XNOR2_X1 U5906 ( .A(n4898), .B(n4897), .ZN(n5639) );
  INV_X1 U5907 ( .A(n8926), .ZN(n4672) );
  NAND2_X1 U5908 ( .A1(n5128), .A2(n5127), .ZN(n9886) );
  INV_X1 U5909 ( .A(n9886), .ZN(n4671) );
  AND2_X1 U5910 ( .A1(n8972), .A2(n4997), .ZN(n7021) );
  AND4_X1 U5911 ( .A1(n5699), .A2(n5698), .A3(n5697), .A4(n5696), .ZN(n6957)
         );
  AND2_X1 U5912 ( .A1(n8419), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4378) );
  NAND2_X1 U5913 ( .A1(n5169), .A2(n5168), .ZN(n4379) );
  INV_X1 U5914 ( .A(n6086), .ZN(n4768) );
  NOR2_X1 U5915 ( .A1(n7057), .A2(P2_U3152), .ZN(n7702) );
  NAND2_X1 U5916 ( .A1(n7303), .A2(n6956), .ZN(n7005) );
  INV_X1 U5917 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4696) );
  INV_X1 U5918 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n4481) );
  NAND2_X1 U5919 ( .A1(n7493), .A2(n8193), .ZN(n7303) );
  NAND2_X1 U5920 ( .A1(n4681), .A2(n7006), .ZN(n4381) );
  INV_X1 U5921 ( .A(n6295), .ZN(n4383) );
  NAND2_X1 U5922 ( .A1(n4384), .A2(n6162), .ZN(n6167) );
  NAND2_X1 U5923 ( .A1(n4385), .A2(n6154), .ZN(n4384) );
  NAND2_X1 U5924 ( .A1(n4387), .A2(n4386), .ZN(n4385) );
  NAND2_X1 U5925 ( .A1(n6142), .A2(n6288), .ZN(n4387) );
  NAND2_X1 U5926 ( .A1(n4388), .A2(n4347), .ZN(n6217) );
  AND2_X2 U5927 ( .A1(n5788), .A2(n5665), .ZN(n5895) );
  NOR2_X2 U5928 ( .A1(n5743), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5774) );
  AOI21_X1 U5929 ( .B1(n4391), .B2(n6278), .A(n6280), .ZN(n4683) );
  AOI21_X1 U5930 ( .B1(n4393), .B2(n6271), .A(n6270), .ZN(n4392) );
  NAND2_X1 U5931 ( .A1(n4994), .A2(n8976), .ZN(n4998) );
  XNOR2_X1 U5932 ( .A(n5000), .B(n5001), .ZN(n8976) );
  AND2_X2 U5933 ( .A1(n4397), .A2(n4396), .ZN(n4945) );
  NAND2_X1 U5934 ( .A1(n4398), .A2(n4400), .ZN(n4449) );
  NAND2_X1 U5935 ( .A1(n5109), .A2(n5110), .ZN(n8919) );
  OR2_X1 U5936 ( .A1(n5055), .A2(n4407), .ZN(n4402) );
  NAND2_X1 U5937 ( .A1(n8974), .A2(n4793), .ZN(n4406) );
  INV_X1 U5938 ( .A(n7244), .ZN(n4407) );
  OAI21_X2 U5939 ( .B1(n8964), .B2(n8965), .A(n4462), .ZN(n8939) );
  NAND2_X2 U5940 ( .A1(n4792), .A2(n4790), .ZN(n7913) );
  NAND3_X1 U5941 ( .A1(n4352), .A2(n4413), .A3(n4412), .ZN(n4411) );
  NAND3_X1 U5942 ( .A1(n4416), .A2(n6464), .A3(n4415), .ZN(n6470) );
  NAND3_X1 U5943 ( .A1(n6456), .A2(n4421), .A3(n4417), .ZN(n4416) );
  NAND2_X1 U5944 ( .A1(n4427), .A2(n4423), .ZN(n5094) );
  NAND2_X1 U5945 ( .A1(n4691), .A2(n4330), .ZN(n4426) );
  NAND2_X1 U5946 ( .A1(n4424), .A2(n5015), .ZN(n4427) );
  NAND2_X1 U5947 ( .A1(n4330), .A2(n5014), .ZN(n4425) );
  NAND2_X1 U5948 ( .A1(n6754), .A2(n6865), .ZN(n4433) );
  NAND2_X1 U5949 ( .A1(n7913), .A2(n4321), .ZN(n8045) );
  NAND2_X1 U5950 ( .A1(n4434), .A2(n4315), .ZN(n8027) );
  NAND2_X1 U5951 ( .A1(n7913), .A2(n4357), .ZN(n4434) );
  NAND2_X1 U5952 ( .A1(n4436), .A2(n5269), .ZN(n8043) );
  NAND2_X1 U5953 ( .A1(n7913), .A2(n7908), .ZN(n4436) );
  NAND2_X1 U5954 ( .A1(n4451), .A2(n4452), .ZN(n8895) );
  NAND2_X1 U5955 ( .A1(n8964), .A2(n4454), .ZN(n4451) );
  NOR2_X1 U5956 ( .A1(n4874), .A2(n4873), .ZN(n4882) );
  INV_X1 U5957 ( .A(n4490), .ZN(n8717) );
  NOR2_X1 U5958 ( .A1(n8700), .A2(n8828), .ZN(n8684) );
  NAND3_X1 U5959 ( .A1(n4506), .A2(n8769), .A3(n4345), .ZN(n8866) );
  AND2_X2 U5960 ( .A1(n4510), .A2(n4508), .ZN(n8587) );
  OAI21_X1 U5961 ( .B1(n4517), .B2(n7409), .A(n7408), .ZN(n7425) );
  XNOR2_X1 U5962 ( .A(n4517), .B(n6113), .ZN(n7316) );
  NAND2_X1 U5963 ( .A1(n4518), .A2(n4527), .ZN(n8715) );
  NAND3_X1 U5964 ( .A1(n4519), .A2(n7993), .A3(n4520), .ZN(n4518) );
  NAND2_X1 U5965 ( .A1(n7890), .A2(n4522), .ZN(n4519) );
  NAND2_X1 U5966 ( .A1(n8751), .A2(n4530), .ZN(n4528) );
  NAND4_X1 U5967 ( .A1(n4788), .A2(n5774), .A3(n4534), .A4(n4356), .ZN(n5673)
         );
  AOI21_X2 U5968 ( .B1(n8663), .B2(n8470), .A(n4537), .ZN(n8651) );
  NOR2_X2 U5969 ( .A1(n8575), .A2(n8579), .ZN(n8574) );
  OR2_X1 U5970 ( .A1(n7788), .A2(n7787), .ZN(n7869) );
  AOI22_X1 U5971 ( .A1(n8508), .A2(n8514), .B1(n8488), .B2(n8511), .ZN(n8490)
         );
  NAND2_X1 U5972 ( .A1(n8715), .A2(n8725), .ZN(n8714) );
  NOR2_X1 U5973 ( .A1(n7799), .A2(n7867), .ZN(n7868) );
  NAND2_X2 U5974 ( .A1(n6175), .A2(n6174), .ZN(n7714) );
  NAND2_X1 U5975 ( .A1(n7709), .A2(n7509), .ZN(n7511) );
  NAND2_X1 U5976 ( .A1(n8473), .A2(n4819), .ZN(n8637) );
  NAND2_X1 U5977 ( .A1(n7792), .A2(n7791), .ZN(n7866) );
  INV_X1 U5978 ( .A(n8359), .ZN(n7593) );
  NAND2_X1 U5979 ( .A1(n7593), .A2(n8239), .ZN(n6175) );
  OR2_X2 U5980 ( .A1(n7512), .A2(n7517), .ZN(n7786) );
  NAND2_X2 U5981 ( .A1(n5094), .A2(n5093), .ZN(n5115) );
  NAND2_X1 U5982 ( .A1(n4891), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4694) );
  NAND2_X1 U5983 ( .A1(n8714), .A2(n8462), .ZN(n8698) );
  NAND2_X1 U5984 ( .A1(n4540), .A2(n6916), .ZN(n6915) );
  OAI21_X1 U5985 ( .B1(n4540), .B2(n6916), .A(n6915), .ZN(n7097) );
  OR2_X1 U5986 ( .A1(n4847), .A2(n4545), .ZN(n4542) );
  NAND2_X1 U5987 ( .A1(n4847), .A2(n4846), .ZN(n9645) );
  NAND3_X1 U5988 ( .A1(n4542), .A2(n4541), .A3(n4543), .ZN(n9651) );
  NAND2_X1 U5989 ( .A1(n4847), .A2(n4344), .ZN(n4541) );
  NAND2_X1 U5990 ( .A1(n7749), .A2(n4548), .ZN(n4547) );
  NAND2_X1 U5991 ( .A1(n4547), .A2(n4550), .ZN(n7972) );
  OAI22_X1 U5992 ( .A1(n9279), .A2(n4557), .B1(n4559), .B2(n4323), .ZN(n9239)
         );
  NAND2_X1 U5993 ( .A1(n9239), .A2(n4566), .ZN(n9134) );
  INV_X1 U5994 ( .A(n9129), .ZN(n4564) );
  AND3_X1 U5995 ( .A1(n4839), .A2(n4840), .A3(n4841), .ZN(n4576) );
  AND2_X1 U5996 ( .A1(n4841), .A2(n4845), .ZN(n4570) );
  NAND2_X1 U5997 ( .A1(n9222), .A2(n4349), .ZN(n4579) );
  NAND2_X1 U5998 ( .A1(n9222), .A2(n4583), .ZN(n4581) );
  AOI21_X1 U5999 ( .B1(n9222), .B2(n9227), .A(n9136), .ZN(n9207) );
  OR2_X1 U6000 ( .A1(n7979), .A2(n4592), .ZN(n4591) );
  NAND2_X1 U6001 ( .A1(n5198), .A2(n4607), .ZN(n4605) );
  NAND2_X1 U6002 ( .A1(n5147), .A2(n4824), .ZN(n4615) );
  OAI21_X2 U6003 ( .B1(n5115), .B2(n5114), .A(n5113), .ZN(n5147) );
  NAND2_X1 U6004 ( .A1(n6554), .A2(n8113), .ZN(n4617) );
  OAI21_X1 U6005 ( .B1(n5508), .B2(n5507), .A(n5506), .ZN(n5532) );
  OAI21_X1 U6006 ( .B1(n5508), .B2(n4621), .A(n4619), .ZN(n4627) );
  NAND2_X1 U6007 ( .A1(n6049), .A2(n4377), .ZN(n4628) );
  MUX2_X1 U6008 ( .A(n6626), .B(n6623), .S(n6616), .Z(n5038) );
  MUX2_X1 U6009 ( .A(n5432), .B(n7495), .S(n6617), .Z(n5451) );
  INV_X1 U6010 ( .A(n9310), .ZN(n4638) );
  NAND2_X1 U6011 ( .A1(n4633), .A2(n4631), .ZN(n9283) );
  INV_X1 U6012 ( .A(n4637), .ZN(n4632) );
  NAND2_X1 U6013 ( .A1(n9346), .A2(n4642), .ZN(n4641) );
  NAND2_X1 U6014 ( .A1(n9346), .A2(n9144), .ZN(n9330) );
  INV_X1 U6015 ( .A(n9144), .ZN(n4643) );
  AOI21_X1 U6016 ( .B1(n4646), .B2(n9689), .A(n4644), .ZN(n8007) );
  OAI21_X1 U6017 ( .B1(n7829), .B2(n4645), .A(n7969), .ZN(n4644) );
  NAND2_X1 U6018 ( .A1(n4650), .A2(n4651), .ZN(n8075) );
  NAND3_X1 U6019 ( .A1(n7139), .A2(n7138), .A3(n7478), .ZN(n4650) );
  NAND2_X1 U6020 ( .A1(n9243), .A2(n4656), .ZN(n4655) );
  NAND2_X1 U6021 ( .A1(n4670), .A2(n7228), .ZN(n8069) );
  NAND2_X1 U6022 ( .A1(n5895), .A2(n4677), .ZN(n6082) );
  INV_X1 U6023 ( .A(n6082), .ZN(n6084) );
  NAND2_X1 U6024 ( .A1(n4680), .A2(n4314), .ZN(P2_U3244) );
  MUX2_X1 U6025 ( .A(n6139), .B(n6138), .S(n6281), .Z(n6160) );
  NOR2_X2 U6026 ( .A1(n7005), .A2(n8440), .ZN(n6281) );
  NAND2_X1 U6027 ( .A1(n4967), .A2(n4966), .ZN(n4689) );
  NAND3_X1 U6028 ( .A1(n4687), .A2(n4686), .A3(n4358), .ZN(n5012) );
  NAND3_X1 U6029 ( .A1(n4967), .A2(n4982), .A3(n4966), .ZN(n4687) );
  NAND2_X2 U6030 ( .A1(n4695), .A2(n4693), .ZN(n6616) );
  OAI21_X1 U6031 ( .B1(n8302), .B2(n8301), .A(n8145), .ZN(n8248) );
  NAND2_X1 U6032 ( .A1(n8163), .A2(n4715), .ZN(n4711) );
  OAI21_X1 U6033 ( .B1(n8163), .B2(n4719), .A(n4715), .ZN(n8326) );
  NAND2_X1 U6034 ( .A1(n4711), .A2(n4712), .ZN(n8183) );
  NAND2_X1 U6035 ( .A1(n4722), .A2(n4724), .ZN(n8121) );
  NAND2_X1 U6036 ( .A1(n8101), .A2(n4726), .ZN(n4722) );
  NAND3_X1 U6037 ( .A1(n4736), .A2(n4735), .A3(n4346), .ZN(n4734) );
  NAND3_X1 U6038 ( .A1(n4742), .A2(n7502), .A3(n6185), .ZN(n4736) );
  NAND2_X1 U6039 ( .A1(n6110), .A2(n4745), .ZN(n4744) );
  NAND2_X1 U6040 ( .A1(n7879), .A2(n6201), .ZN(n7992) );
  INV_X1 U6041 ( .A(n4750), .ZN(n7991) );
  INV_X1 U6042 ( .A(n6201), .ZN(n4752) );
  OAI21_X1 U6043 ( .B1(n8657), .B2(n4756), .A(n4754), .ZN(n8615) );
  NAND2_X1 U6044 ( .A1(n4764), .A2(n4765), .ZN(n6101) );
  NAND2_X1 U6045 ( .A1(n8491), .A2(n4351), .ZN(n4764) );
  NAND2_X1 U6046 ( .A1(n6065), .A2(n6283), .ZN(n4772) );
  OAI21_X1 U6047 ( .B1(n8541), .B2(n4778), .A(n4774), .ZN(n8513) );
  NAND3_X1 U6048 ( .A1(n5658), .A2(n5657), .A3(n5659), .ZN(n5741) );
  NAND4_X1 U6049 ( .A1(n4780), .A2(n5658), .A3(n5657), .A4(n5659), .ZN(n5743)
         );
  AND2_X2 U6050 ( .A1(n5670), .A2(n5665), .ZN(n4788) );
  NAND2_X1 U6051 ( .A1(n4799), .A2(n4800), .ZN(n5350) );
  NAND2_X1 U6052 ( .A1(n8948), .A2(n5323), .ZN(n4799) );
  NAND3_X1 U6053 ( .A1(n4802), .A2(n6865), .A3(n4933), .ZN(n6754) );
  NAND2_X1 U6054 ( .A1(n4927), .A2(n4928), .ZN(n6865) );
  NAND2_X1 U6055 ( .A1(n4930), .A2(n4929), .ZN(n4802) );
  NAND2_X1 U6056 ( .A1(n5448), .A2(n4806), .ZN(n4805) );
  INV_X1 U6057 ( .A(n5632), .ZN(n5633) );
  NAND2_X1 U6058 ( .A1(n4899), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4898) );
  NAND2_X1 U6059 ( .A1(n9246), .A2(n9223), .ZN(n9231) );
  XNOR2_X1 U6060 ( .A(n5532), .B(n5531), .ZN(n7939) );
  XNOR2_X1 U6061 ( .A(n4486), .B(n8175), .ZN(n8291) );
  NAND2_X1 U6062 ( .A1(n4918), .A2(n5687), .ZN(n4940) );
  AND2_X1 U6063 ( .A1(n8855), .A2(n7897), .ZN(n6193) );
  NOR2_X1 U6064 ( .A1(n4896), .A2(n4900), .ZN(n4903) );
  NAND2_X1 U6065 ( .A1(n4829), .A2(n4998), .ZN(n4999) );
  AOI21_X1 U6066 ( .B1(n6325), .B2(n5601), .A(n4906), .ZN(n6764) );
  XNOR2_X1 U6067 ( .A(n4977), .B(n4976), .ZN(n5000) );
  AND2_X1 U6068 ( .A1(n7370), .A2(n7369), .ZN(n4816) );
  NAND2_X1 U6069 ( .A1(n7297), .A2(n8553), .ZN(n8667) );
  INV_X1 U6070 ( .A(n5021), .ZN(n5034) );
  AND2_X1 U6071 ( .A1(n9445), .A2(n7974), .ZN(n4817) );
  OR2_X1 U6072 ( .A1(n9445), .A2(n7974), .ZN(n4818) );
  OR2_X1 U6073 ( .A1(n8655), .A2(n8644), .ZN(n4819) );
  OR2_X1 U6074 ( .A1(n9184), .A2(n9197), .ZN(n4821) );
  AND2_X1 U6075 ( .A1(n5631), .A2(n4825), .ZN(n4822) );
  AND3_X1 U6076 ( .A1(n5981), .A2(n5980), .A3(n5979), .ZN(n8475) );
  AND2_X1 U6077 ( .A1(n5171), .A2(n5153), .ZN(n4823) );
  AND2_X1 U6078 ( .A1(n5148), .A2(n5120), .ZN(n4824) );
  INV_X1 U6079 ( .A(n9690), .ZN(n7974) );
  AND4_X1 U6080 ( .A1(n5522), .A2(n5521), .A3(n5520), .A4(n5519), .ZN(n9135)
         );
  AND2_X1 U6081 ( .A1(n8893), .A2(n5630), .ZN(n4825) );
  AND2_X1 U6082 ( .A1(n8894), .A2(n8893), .ZN(n4826) );
  OR2_X1 U6083 ( .A1(n7976), .A2(n8016), .ZN(n4827) );
  NAND2_X1 U6084 ( .A1(n7021), .A2(n8976), .ZN(n4829) );
  INV_X1 U6085 ( .A(n8828), .ZN(n8466) );
  INV_X1 U6086 ( .A(n9389), .ZN(n9223) );
  NOR2_X1 U6087 ( .A1(n5310), .A2(n5287), .ZN(n4830) );
  OAI21_X1 U6088 ( .B1(n7419), .B2(n6116), .A(n6140), .ZN(n7544) );
  AND3_X1 U6089 ( .A1(n4936), .A2(n4935), .A3(n4934), .ZN(n4831) );
  AND2_X1 U6090 ( .A1(n6153), .A2(n6157), .ZN(n6154) );
  INV_X1 U6091 ( .A(n7707), .ZN(n6165) );
  NOR2_X1 U6092 ( .A1(n6171), .A2(n7714), .ZN(n6172) );
  AND2_X1 U6093 ( .A1(n6233), .A2(n6232), .ZN(n6234) );
  NOR2_X1 U6094 ( .A1(n6242), .A2(n6248), .ZN(n6243) );
  INV_X1 U6095 ( .A(n6156), .ZN(n5732) );
  INV_X1 U6096 ( .A(n8450), .ZN(n6100) );
  AOI21_X1 U6097 ( .B1(n6141), .B2(n6114), .A(n5732), .ZN(n5733) );
  INV_X1 U6098 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U6099 ( .A1(n9054), .A2(n5602), .ZN(n4950) );
  INV_X1 U6100 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4832) );
  NAND2_X1 U6101 ( .A1(n8291), .A2(n8157), .ZN(n8155) );
  AND2_X1 U6102 ( .A1(n6143), .A2(n6149), .ZN(n6953) );
  INV_X1 U6103 ( .A(n6177), .ZN(n6182) );
  OAI22_X1 U6104 ( .A1(n4993), .A2(n5596), .B1(n7264), .B2(n5499), .ZN(n4992)
         );
  NAND2_X1 U6105 ( .A1(n8158), .A2(n8290), .ZN(n8159) );
  AND2_X1 U6106 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5747) );
  INV_X1 U6107 ( .A(n7514), .ZN(n7517) );
  NOR2_X1 U6108 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4900) );
  NOR2_X1 U6109 ( .A1(n5260), .A2(n5259), .ZN(n5286) );
  NAND2_X1 U6110 ( .A1(n9051), .A2(n9853), .ZN(n6421) );
  INV_X1 U6111 ( .A(n7940), .ZN(n5608) );
  AND2_X1 U6112 ( .A1(n5122), .A2(n4838), .ZN(n4881) );
  OR2_X1 U6113 ( .A1(n5373), .A2(n5372), .ZN(n5376) );
  INV_X1 U6114 ( .A(n5089), .ZN(n5090) );
  INV_X1 U6115 ( .A(n5929), .ZN(n5927) );
  NAND2_X1 U6116 ( .A1(n8160), .A2(n8159), .ZN(n8161) );
  OR2_X1 U6117 ( .A1(n5977), .A2(n8313), .ZN(n5985) );
  OR2_X1 U6118 ( .A1(n5851), .A2(n7567), .ZN(n5869) );
  INV_X1 U6119 ( .A(n8475), .ZN(n8476) );
  OR2_X1 U6120 ( .A1(n7786), .A2(n7790), .ZN(n7787) );
  OAI21_X1 U6121 ( .B1(n8723), .B2(n5909), .A(n6207), .ZN(n8689) );
  OR2_X1 U6122 ( .A1(n5773), .A2(n6629), .ZN(n5730) );
  AOI22_X1 U6123 ( .A1(n6885), .A2(n5586), .B1(n4907), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n4908) );
  NAND2_X1 U6124 ( .A1(n5411), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5435) );
  OR2_X1 U6125 ( .A1(n5130), .A2(n5129), .ZN(n5158) );
  AND2_X1 U6126 ( .A1(n5589), .A2(n5565), .ZN(n9194) );
  AND3_X1 U6127 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5029) );
  AND2_X1 U6128 ( .A1(n9366), .A2(n9887), .ZN(n9367) );
  INV_X1 U6129 ( .A(n9179), .ZN(n9187) );
  AOI21_X1 U6130 ( .B1(n9143), .B2(n9142), .A(n9141), .ZN(n9346) );
  OR2_X1 U6131 ( .A1(n6090), .A2(n6089), .ZN(n6091) );
  NAND2_X1 U6132 ( .A1(n5151), .A2(n5150), .ZN(n5171) );
  INV_X1 U6133 ( .A(n8361), .ZN(n7384) );
  NAND2_X1 U6134 ( .A1(n7964), .A2(n6071), .ZN(n6021) );
  NAND2_X1 U6135 ( .A1(n5927), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5953) );
  OR2_X1 U6136 ( .A1(n5780), .A2(n5779), .ZN(n5798) );
  INV_X1 U6137 ( .A(n8345), .ZN(n8314) );
  NAND2_X1 U6138 ( .A1(n5695), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5711) );
  INV_X1 U6139 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9586) );
  INV_X1 U6140 ( .A(n8492), .ZN(n8489) );
  NAND2_X1 U6141 ( .A1(n8447), .A2(n8352), .ZN(n8483) );
  AND2_X1 U6142 ( .A1(n6232), .A2(n6237), .ZN(n8656) );
  INV_X1 U6143 ( .A(n8458), .ZN(n8727) );
  AND2_X1 U6144 ( .A1(n7001), .A2(n8001), .ZN(n8630) );
  AND2_X1 U6145 ( .A1(n6956), .A2(n6955), .ZN(n8724) );
  AND2_X1 U6146 ( .A1(n9939), .A2(n6997), .ZN(n8856) );
  AND2_X1 U6147 ( .A1(n6163), .A2(n6157), .ZN(n7546) );
  AND2_X1 U6148 ( .A1(n7945), .A2(n6938), .ZN(n6939) );
  OR2_X1 U6149 ( .A1(n5034), .A2(n6626), .ZN(n5022) );
  AND2_X1 U6150 ( .A1(n5386), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5411) );
  INV_X1 U6151 ( .A(n9366), .ZN(n9174) );
  AND2_X1 U6152 ( .A1(n9409), .A2(n9302), .ZN(n9129) );
  NOR2_X1 U6153 ( .A1(n9368), .A2(n9367), .ZN(n9369) );
  AND2_X1 U6154 ( .A1(n6459), .A2(n7970), .ZN(n8008) );
  AOI21_X1 U6155 ( .B1(n7126), .B2(n7224), .A(n7125), .ZN(n7127) );
  INV_X1 U6156 ( .A(n9887), .ZN(n9852) );
  AND2_X1 U6157 ( .A1(n8282), .A2(n8632), .ZN(n8345) );
  INV_X1 U6158 ( .A(n9917), .ZN(n9912) );
  AND2_X1 U6159 ( .A1(n6774), .A2(n6773), .ZN(n9914) );
  AND2_X1 U6160 ( .A1(n7986), .A2(n7874), .ZN(n8847) );
  NOR2_X1 U6161 ( .A1(n9933), .A2(n6944), .ZN(n7292) );
  OR3_X1 U6162 ( .A1(n6950), .A2(n6961), .A3(n8440), .ZN(n8854) );
  INV_X1 U6163 ( .A(n9985), .ZN(n8861) );
  AND2_X1 U6164 ( .A1(n6943), .A2(n6942), .ZN(n6967) );
  AND2_X1 U6165 ( .A1(n9024), .A2(n9887), .ZN(n9038) );
  AND4_X1 U6166 ( .A1(n5498), .A2(n5497), .A3(n5496), .A4(n5495), .ZN(n9259)
         );
  AND4_X1 U6167 ( .A1(n5291), .A2(n5290), .A3(n5289), .A4(n5288), .ZN(n7976)
         );
  AND2_X1 U6168 ( .A1(n6338), .A2(n9137), .ZN(n9210) );
  AND2_X1 U6169 ( .A1(n9329), .A2(n9144), .ZN(n9339) );
  AND2_X1 U6170 ( .A1(n6895), .A2(n6894), .ZN(n9347) );
  OR2_X1 U6171 ( .A1(n5649), .A2(n9837), .ZN(n9685) );
  AND2_X1 U6172 ( .A1(n5650), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9033) );
  INV_X1 U6173 ( .A(n9873), .ZN(n9892) );
  AND2_X1 U6174 ( .A1(n6517), .A2(n7093), .ZN(n9884) );
  INV_X1 U6175 ( .A(n6611), .ZN(n6980) );
  INV_X1 U6176 ( .A(n8446), .ZN(n9920) );
  INV_X1 U6177 ( .A(n8333), .ZN(n8341) );
  NAND2_X1 U6178 ( .A1(n7004), .A2(n7003), .ZN(n8349) );
  INV_X1 U6179 ( .A(n8516), .ZN(n8485) );
  INV_X1 U6180 ( .A(n8448), .ZN(n8760) );
  XNOR2_X1 U6181 ( .A(n8508), .B(n8507), .ZN(n8774) );
  INV_X1 U6182 ( .A(n8667), .ZN(n8686) );
  INV_X1 U6183 ( .A(n10001), .ZN(n9999) );
  INV_X1 U6184 ( .A(n9988), .ZN(n9987) );
  INV_X1 U6185 ( .A(n9931), .ZN(n9934) );
  XNOR2_X1 U6186 ( .A(n6303), .B(n6302), .ZN(n7813) );
  INV_X1 U6187 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9501) );
  INV_X1 U6188 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6623) );
  XNOR2_X1 U6189 ( .A(n8895), .B(n4826), .ZN(n8901) );
  NOR2_X1 U6190 ( .A1(n5635), .A2(n5653), .ZN(n5654) );
  OR2_X1 U6191 ( .A1(n5637), .A2(n5629), .ZN(n9012) );
  INV_X1 U6192 ( .A(n9259), .ZN(n9230) );
  XOR2_X1 U6193 ( .A(n9169), .B(n9360), .Z(n9363) );
  NAND2_X1 U6194 ( .A1(n7130), .A2(n9685), .ZN(n9725) );
  OR2_X1 U6195 ( .A1(n9831), .A2(n9837), .ZN(n9835) );
  INV_X1 U6196 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U6197 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4835) );
  NOR2_X1 U6198 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4834) );
  INV_X1 U6199 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4833) );
  INV_X1 U6200 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4838) );
  INV_X1 U6201 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5330) );
  NOR2_X1 U6202 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4841) );
  NOR2_X1 U6203 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4840) );
  NOR2_X1 U6204 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n4839) );
  INV_X1 U6205 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4843) );
  INV_X1 U6206 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4860) );
  INV_X1 U6207 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4842) );
  INV_X1 U6208 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4845) );
  INV_X1 U6209 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4897) );
  INV_X1 U6210 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4846) );
  NAND2_X1 U6211 ( .A1(n4849), .A2(n4848), .ZN(n4850) );
  NAND2_X1 U6212 ( .A1(n4850), .A2(n9645), .ZN(n4852) );
  NAND2_X1 U6213 ( .A1(n5591), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4856) );
  INV_X1 U6214 ( .A(n9651), .ZN(n4851) );
  AND2_X2 U6215 ( .A1(n4851), .A2(n8024), .ZN(n5209) );
  NAND2_X1 U6216 ( .A1(n5209), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4855) );
  NAND2_X1 U6217 ( .A1(n5056), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n4854) );
  NAND2_X1 U6218 ( .A1(n5084), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4853) );
  INV_X1 U6219 ( .A(n4861), .ZN(n5614) );
  NAND2_X1 U6220 ( .A1(n5614), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4859) );
  NAND2_X1 U6221 ( .A1(n4861), .A2(n4860), .ZN(n4864) );
  NAND2_X1 U6222 ( .A1(n4862), .A2(n4864), .ZN(n5607) );
  INV_X1 U6223 ( .A(n7943), .ZN(n4863) );
  NAND2_X1 U6224 ( .A1(n4864), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4865) );
  NAND2_X2 U6225 ( .A1(n4868), .A2(n7940), .ZN(n4904) );
  INV_X1 U6226 ( .A(n5205), .ZN(n4874) );
  NOR2_X1 U6227 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4872) );
  NOR2_X1 U6228 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4871) );
  NOR2_X1 U6229 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n4870) );
  NOR2_X1 U6230 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4869) );
  NAND4_X1 U6231 ( .A1(n4872), .A2(n4871), .A3(n4870), .A4(n4869), .ZN(n4873)
         );
  XNOR2_X1 U6232 ( .A(n4887), .B(n4886), .ZN(n5628) );
  INV_X1 U6233 ( .A(n5628), .ZN(n7472) );
  NAND2_X1 U6234 ( .A1(n7472), .A2(n7093), .ZN(n6890) );
  INV_X1 U6235 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5282) );
  INV_X1 U6236 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6237 ( .A1(n5282), .A2(n5254), .ZN(n4877) );
  INV_X1 U6238 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4878) );
  NAND2_X1 U6239 ( .A1(n5306), .A2(n4878), .ZN(n5329) );
  INV_X1 U6240 ( .A(n5329), .ZN(n4880) );
  NOR2_X1 U6241 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n4879) );
  INV_X1 U6242 ( .A(n5383), .ZN(n7099) );
  NAND2_X1 U6243 ( .A1(n7099), .A2(n7093), .ZN(n7199) );
  NAND2_X1 U6244 ( .A1(n4887), .A2(n4886), .ZN(n4888) );
  NAND2_X1 U6245 ( .A1(n4888), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4890) );
  INV_X1 U6246 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4889) );
  INV_X1 U6247 ( .A(n4299), .ZN(n6617) );
  INV_X1 U6248 ( .A(SI_0_), .ZN(n4893) );
  INV_X1 U6249 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4892) );
  OAI21_X1 U6250 ( .B1(n6617), .B2(n4893), .A(n4892), .ZN(n4895) );
  AND2_X1 U6251 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4894) );
  NAND2_X1 U6252 ( .A1(n4916), .A2(n4894), .ZN(n4918) );
  AND2_X1 U6253 ( .A1(n4895), .A2(n4918), .ZN(n9656) );
  NAND2_X1 U6254 ( .A1(n4338), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4901) );
  MUX2_X1 U6255 ( .A(n9655), .B(n9656), .S(n6574), .Z(n6885) );
  INV_X1 U6256 ( .A(n6890), .ZN(n7092) );
  AND2_X4 U6257 ( .A1(n7092), .A2(n4904), .ZN(n5602) );
  NAND2_X1 U6258 ( .A1(n6885), .A2(n5602), .ZN(n4905) );
  OAI21_X1 U6259 ( .B1(n4396), .B2(n4904), .A(n4905), .ZN(n4906) );
  NAND2_X1 U6260 ( .A1(n6325), .A2(n5602), .ZN(n4909) );
  INV_X1 U6261 ( .A(n4904), .ZN(n4907) );
  NAND2_X1 U6262 ( .A1(n4909), .A2(n4908), .ZN(n6763) );
  NAND2_X1 U6263 ( .A1(n6764), .A2(n6763), .ZN(n6762) );
  INV_X1 U6264 ( .A(n6763), .ZN(n4910) );
  NAND2_X1 U6265 ( .A1(n4910), .A2(n5599), .ZN(n4911) );
  NAND2_X1 U6266 ( .A1(n6762), .A2(n4911), .ZN(n4927) );
  NAND2_X1 U6267 ( .A1(n5056), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4914) );
  NAND2_X1 U6268 ( .A1(n5084), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4913) );
  NAND4_X4 U6269 ( .A1(n4915), .A2(n4914), .A3(n4913), .A4(n4912), .ZN(n6326)
         );
  NAND2_X1 U6270 ( .A1(n6326), .A2(n5602), .ZN(n4925) );
  AND2_X1 U6271 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4917) );
  NAND2_X1 U6272 ( .A1(n6616), .A2(n4917), .ZN(n5687) );
  INV_X1 U6273 ( .A(SI_1_), .ZN(n4919) );
  INV_X2 U6274 ( .A(n6616), .ZN(n5327) );
  MUX2_X1 U6275 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5327), .Z(n4938) );
  XNOR2_X1 U6276 ( .A(n4939), .B(n4938), .ZN(n6618) );
  NAND2_X1 U6277 ( .A1(n5021), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4922) );
  NAND2_X1 U6278 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n9655), .ZN(n4920) );
  NAND2_X1 U6279 ( .A1(n4988), .A2(n4300), .ZN(n4921) );
  NAND2_X1 U6280 ( .A1(n4925), .A2(n4924), .ZN(n4926) );
  XNOR2_X1 U6281 ( .A(n4926), .B(n4976), .ZN(n4928) );
  INV_X1 U6282 ( .A(n4927), .ZN(n4930) );
  INV_X1 U6283 ( .A(n4928), .ZN(n4929) );
  NAND2_X1 U6284 ( .A1(n6326), .A2(n5601), .ZN(n4932) );
  OR2_X1 U6285 ( .A1(n6920), .A2(n5596), .ZN(n4931) );
  NAND2_X1 U6286 ( .A1(n4932), .A2(n4931), .ZN(n6757) );
  NAND2_X1 U6287 ( .A1(n5056), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n4937) );
  NAND2_X1 U6288 ( .A1(n5591), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n4936) );
  NAND2_X1 U6289 ( .A1(n5209), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4935) );
  NAND2_X1 U6290 ( .A1(n5084), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4934) );
  NAND2_X2 U6291 ( .A1(n4937), .A2(n4831), .ZN(n9054) );
  NAND2_X1 U6292 ( .A1(n4939), .A2(n4938), .ZN(n4942) );
  NAND2_X1 U6293 ( .A1(n4940), .A2(SI_1_), .ZN(n4941) );
  NAND2_X1 U6294 ( .A1(n4942), .A2(n4941), .ZN(n4967) );
  INV_X1 U6295 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6621) );
  INV_X1 U6296 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4943) );
  MUX2_X1 U6297 ( .A(n6621), .B(n4943), .S(n5327), .Z(n4968) );
  XNOR2_X1 U6298 ( .A(n4967), .B(n4966), .ZN(n6631) );
  INV_X1 U6299 ( .A(n6631), .ZN(n4944) );
  NAND2_X1 U6300 ( .A1(n5009), .A2(n4944), .ZN(n4948) );
  NAND2_X1 U6301 ( .A1(n5021), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4947) );
  NAND2_X1 U6302 ( .A1(n4988), .A2(n9750), .ZN(n4946) );
  AND3_X2 U6303 ( .A1(n4948), .A2(n4947), .A3(n4946), .ZN(n7214) );
  OR2_X1 U6304 ( .A1(n7214), .A2(n5499), .ZN(n4949) );
  NAND2_X1 U6305 ( .A1(n4950), .A2(n4949), .ZN(n4951) );
  INV_X1 U6306 ( .A(n7214), .ZN(n6872) );
  AOI22_X1 U6307 ( .A1(n9054), .A2(n5601), .B1(n6872), .B2(n5602), .ZN(n4953)
         );
  NAND2_X1 U6308 ( .A1(n4952), .A2(n4953), .ZN(n7023) );
  INV_X1 U6309 ( .A(n4952), .ZN(n4955) );
  INV_X1 U6310 ( .A(n4953), .ZN(n4954) );
  NAND2_X1 U6311 ( .A1(n4955), .A2(n4954), .ZN(n4956) );
  NAND2_X1 U6312 ( .A1(n5056), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n4961) );
  NAND2_X1 U6313 ( .A1(n5084), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4960) );
  INV_X1 U6314 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n4957) );
  XNOR2_X1 U6315 ( .A(n4957), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n8981) );
  NAND2_X1 U6316 ( .A1(n5413), .A2(n8981), .ZN(n4959) );
  NAND2_X1 U6317 ( .A1(n5209), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n4958) );
  NAND2_X1 U6318 ( .A1(n5021), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4965) );
  NAND2_X1 U6319 ( .A1(n4962), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4963) );
  XNOR2_X1 U6320 ( .A(n4963), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9769) );
  NAND2_X1 U6321 ( .A1(n4988), .A2(n9769), .ZN(n4964) );
  INV_X1 U6322 ( .A(n4968), .ZN(n4969) );
  NAND2_X1 U6323 ( .A1(n4969), .A2(SI_2_), .ZN(n4970) );
  INV_X1 U6324 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n4971) );
  MUX2_X1 U6325 ( .A(n6620), .B(n4971), .S(n5327), .Z(n4972) );
  INV_X1 U6326 ( .A(n4972), .ZN(n4973) );
  MUX2_X1 U6327 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n4299), .Z(n5013) );
  XNOR2_X1 U6328 ( .A(n5012), .B(n5010), .ZN(n5725) );
  INV_X1 U6329 ( .A(n5725), .ZN(n6629) );
  OAI22_X1 U6330 ( .A1(n7113), .A2(n5026), .B1(n9847), .B2(n5596), .ZN(n5001)
         );
  NAND2_X1 U6331 ( .A1(n5056), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n4981) );
  NAND2_X1 U6332 ( .A1(n5084), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4980) );
  NAND2_X1 U6333 ( .A1(n5209), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4979) );
  INV_X1 U6334 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7029) );
  NAND2_X1 U6335 ( .A1(n5591), .A2(n7029), .ZN(n4978) );
  XNOR2_X1 U6336 ( .A(n4983), .B(n4982), .ZN(n6633) );
  NAND2_X1 U6337 ( .A1(n5021), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4990) );
  INV_X1 U6338 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4984) );
  NAND2_X1 U6339 ( .A1(n4985), .A2(n4984), .ZN(n4986) );
  NAND2_X1 U6340 ( .A1(n4986), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4987) );
  XNOR2_X2 U6341 ( .A(n4987), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U6342 ( .A1(n4988), .A2(n6673), .ZN(n4989) );
  XNOR2_X1 U6343 ( .A(n4992), .B(n5599), .ZN(n4996) );
  OAI22_X1 U6344 ( .A1(n4993), .A2(n5026), .B1(n7264), .B2(n5596), .ZN(n4995)
         );
  INV_X1 U6345 ( .A(n8972), .ZN(n4994) );
  NAND2_X1 U6346 ( .A1(n4996), .A2(n4995), .ZN(n4997) );
  INV_X1 U6347 ( .A(n5000), .ZN(n5002) );
  OR2_X1 U6348 ( .A1(n5002), .A2(n5001), .ZN(n5003) );
  NAND2_X1 U6349 ( .A1(n5056), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5008) );
  NAND2_X1 U6350 ( .A1(n6317), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5007) );
  AOI21_X1 U6351 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5004) );
  NOR2_X1 U6352 ( .A1(n5004), .A2(n5029), .ZN(n7283) );
  NAND2_X1 U6353 ( .A1(n5413), .A2(n7283), .ZN(n5006) );
  INV_X1 U6354 ( .A(n5209), .ZN(n6321) );
  NAND2_X1 U6355 ( .A1(n5209), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5005) );
  NAND2_X1 U6356 ( .A1(n5012), .A2(n5011), .ZN(n5015) );
  NAND2_X1 U6357 ( .A1(n5013), .A2(SI_4_), .ZN(n5014) );
  XNOR2_X1 U6358 ( .A(n5037), .B(n5036), .ZN(n6625) );
  OR2_X1 U6359 ( .A1(n4991), .A2(n6625), .ZN(n5024) );
  NAND2_X1 U6360 ( .A1(n5016), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5017) );
  MUX2_X1 U6361 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5017), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5020) );
  INV_X1 U6362 ( .A(n5018), .ZN(n5019) );
  NAND2_X1 U6363 ( .A1(n4988), .A2(n9783), .ZN(n5023) );
  INV_X1 U6364 ( .A(n7286), .ZN(n9853) );
  OAI22_X1 U6365 ( .A1(n7220), .A2(n5596), .B1(n9853), .B2(n5499), .ZN(n5025)
         );
  XNOR2_X1 U6366 ( .A(n5025), .B(n4976), .ZN(n5052) );
  OR2_X1 U6367 ( .A1(n7220), .A2(n5026), .ZN(n5028) );
  NAND2_X1 U6368 ( .A1(n7286), .A2(n5602), .ZN(n5027) );
  NAND2_X1 U6369 ( .A1(n5028), .A2(n5027), .ZN(n5053) );
  INV_X1 U6370 ( .A(n5053), .ZN(n7320) );
  NAND2_X1 U6371 ( .A1(n5209), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5033) );
  NAND2_X1 U6372 ( .A1(n6344), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5032) );
  NAND2_X1 U6373 ( .A1(n5029), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5058) );
  OAI21_X1 U6374 ( .B1(n5029), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5058), .ZN(
        n7231) );
  INV_X1 U6375 ( .A(n7231), .ZN(n9021) );
  NAND2_X1 U6376 ( .A1(n5413), .A2(n9021), .ZN(n5031) );
  NAND2_X1 U6377 ( .A1(n6317), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5030) );
  OR2_X1 U6378 ( .A1(n5018), .A2(n5122), .ZN(n5035) );
  XNOR2_X1 U6379 ( .A(n5035), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6634) );
  AOI22_X1 U6380 ( .A1(n5021), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n4988), .B2(
        n6634), .ZN(n5043) );
  INV_X1 U6381 ( .A(n5038), .ZN(n5039) );
  NAND2_X1 U6382 ( .A1(n5039), .A2(SI_5_), .ZN(n5040) );
  INV_X1 U6383 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5041) );
  MUX2_X1 U6384 ( .A(n6637), .B(n5041), .S(n4299), .Z(n5066) );
  XNOR2_X1 U6385 ( .A(n5065), .B(n5064), .ZN(n6636) );
  OR2_X1 U6386 ( .A1(n6636), .A2(n4991), .ZN(n5042) );
  NAND2_X1 U6387 ( .A1(n5043), .A2(n5042), .ZN(n9023) );
  OAI22_X1 U6388 ( .A1(n7322), .A2(n5596), .B1(n7230), .B2(n5499), .ZN(n5044)
         );
  XNOR2_X1 U6389 ( .A(n5044), .B(n4976), .ZN(n5048) );
  OR2_X1 U6390 ( .A1(n7322), .A2(n5026), .ZN(n5046) );
  NAND2_X1 U6391 ( .A1(n9023), .A2(n5602), .ZN(n5045) );
  NAND2_X1 U6392 ( .A1(n5046), .A2(n5045), .ZN(n5049) );
  INV_X1 U6393 ( .A(n5049), .ZN(n5047) );
  NAND2_X1 U6394 ( .A1(n5048), .A2(n5047), .ZN(n7244) );
  INV_X1 U6395 ( .A(n5048), .ZN(n5050) );
  NAND2_X1 U6396 ( .A1(n5050), .A2(n5049), .ZN(n5051) );
  NAND2_X1 U6397 ( .A1(n7244), .A2(n5051), .ZN(n9016) );
  INV_X1 U6398 ( .A(n5052), .ZN(n7318) );
  AND2_X1 U6399 ( .A1(n7318), .A2(n5053), .ZN(n5054) );
  NOR2_X1 U6400 ( .A1(n9016), .A2(n5054), .ZN(n5055) );
  NAND2_X1 U6401 ( .A1(n6343), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5063) );
  NAND2_X1 U6402 ( .A1(n5056), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5062) );
  AND2_X1 U6403 ( .A1(n5058), .A2(n5057), .ZN(n5059) );
  NOR2_X1 U6404 ( .A1(n5082), .A2(n5059), .ZN(n7132) );
  NAND2_X1 U6405 ( .A1(n5413), .A2(n7132), .ZN(n5061) );
  NAND2_X1 U6406 ( .A1(n5084), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5060) );
  INV_X1 U6407 ( .A(n5066), .ZN(n5067) );
  MUX2_X1 U6408 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5700), .Z(n5092) );
  XNOR2_X1 U6409 ( .A(n5091), .B(n5089), .ZN(n6642) );
  NAND2_X1 U6410 ( .A1(n6642), .A2(n5009), .ZN(n5071) );
  NAND2_X1 U6411 ( .A1(n5018), .A2(n5068), .ZN(n5100) );
  NAND2_X1 U6412 ( .A1(n5100), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5069) );
  XNOR2_X1 U6413 ( .A(n5069), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6691) );
  AOI22_X1 U6414 ( .A1(n5021), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n4988), .B2(
        n6691), .ZN(n5070) );
  NAND2_X1 U6415 ( .A1(n5071), .A2(n5070), .ZN(n7243) );
  NAND2_X1 U6416 ( .A1(n7243), .A2(n5586), .ZN(n5072) );
  OAI21_X1 U6417 ( .B1(n7336), .B2(n5596), .A(n5072), .ZN(n5073) );
  XNOR2_X1 U6418 ( .A(n5073), .B(n4976), .ZN(n5077) );
  OR2_X1 U6419 ( .A1(n7336), .A2(n5026), .ZN(n5075) );
  NAND2_X1 U6420 ( .A1(n7243), .A2(n5602), .ZN(n5074) );
  NAND2_X1 U6421 ( .A1(n5075), .A2(n5074), .ZN(n5078) );
  INV_X1 U6422 ( .A(n5078), .ZN(n5076) );
  NAND2_X1 U6423 ( .A1(n5077), .A2(n5076), .ZN(n5081) );
  INV_X1 U6424 ( .A(n5077), .ZN(n5079) );
  NAND2_X1 U6425 ( .A1(n5079), .A2(n5078), .ZN(n5080) );
  AND2_X1 U6426 ( .A1(n5081), .A2(n5080), .ZN(n7245) );
  NAND2_X1 U6427 ( .A1(n6343), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5088) );
  NAND2_X1 U6428 ( .A1(n5056), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5087) );
  NAND2_X1 U6429 ( .A1(n5082), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5130) );
  OR2_X1 U6430 ( .A1(n5082), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5083) );
  AND2_X1 U6431 ( .A1(n5130), .A2(n5083), .ZN(n8925) );
  NAND2_X1 U6432 ( .A1(n5413), .A2(n8925), .ZN(n5086) );
  NAND2_X1 U6433 ( .A1(n5084), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5085) );
  OR2_X1 U6434 ( .A1(n8076), .A2(n5026), .ZN(n5105) );
  NAND2_X1 U6435 ( .A1(n5092), .A2(SI_7_), .ZN(n5093) );
  INV_X1 U6436 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5095) );
  MUX2_X1 U6437 ( .A(n9501), .B(n5095), .S(n4299), .Z(n5097) );
  INV_X1 U6438 ( .A(SI_8_), .ZN(n5096) );
  INV_X1 U6439 ( .A(n5097), .ZN(n5098) );
  NAND2_X1 U6440 ( .A1(n5098), .A2(SI_8_), .ZN(n5099) );
  NAND2_X1 U6441 ( .A1(n6646), .A2(n5009), .ZN(n5103) );
  NAND2_X1 U6442 ( .A1(n5121), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5101) );
  XNOR2_X1 U6443 ( .A(n5101), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9807) );
  AOI22_X1 U6444 ( .A1(n5021), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n4988), .B2(
        n9807), .ZN(n5102) );
  NAND2_X1 U6445 ( .A1(n5103), .A2(n5102), .ZN(n8926) );
  NAND2_X1 U6446 ( .A1(n8926), .A2(n5602), .ZN(n5104) );
  AND2_X1 U6447 ( .A1(n5105), .A2(n5104), .ZN(n5110) );
  NAND2_X1 U6448 ( .A1(n8926), .A2(n5586), .ZN(n5107) );
  OR2_X1 U6449 ( .A1(n8076), .A2(n5596), .ZN(n5106) );
  NAND2_X1 U6450 ( .A1(n5107), .A2(n5106), .ZN(n5108) );
  XNOR2_X1 U6451 ( .A(n5108), .B(n5599), .ZN(n8921) );
  INV_X1 U6452 ( .A(n5110), .ZN(n5111) );
  INV_X1 U6453 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6663) );
  INV_X1 U6454 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5116) );
  MUX2_X1 U6455 ( .A(n6663), .B(n5116), .S(n4299), .Z(n5118) );
  INV_X1 U6456 ( .A(SI_9_), .ZN(n5117) );
  INV_X1 U6457 ( .A(n5118), .ZN(n5119) );
  NAND2_X1 U6458 ( .A1(n5119), .A2(SI_9_), .ZN(n5120) );
  NAND2_X1 U6459 ( .A1(n6660), .A2(n5009), .ZN(n5128) );
  NOR2_X1 U6460 ( .A1(n5121), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5125) );
  OR2_X1 U6461 ( .A1(n5125), .A2(n5122), .ZN(n5123) );
  INV_X1 U6462 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5124) );
  MUX2_X1 U6463 ( .A(n5123), .B(P1_IR_REG_31__SCAN_IN), .S(n5124), .Z(n5126)
         );
  NAND2_X1 U6464 ( .A1(n5125), .A2(n5124), .ZN(n5174) );
  NAND2_X1 U6465 ( .A1(n5126), .A2(n5174), .ZN(n6611) );
  AOI22_X1 U6466 ( .A1(n5021), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n4988), .B2(
        n6980), .ZN(n5127) );
  NAND2_X1 U6467 ( .A1(n9886), .A2(n5586), .ZN(n5137) );
  INV_X1 U6468 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U6469 ( .A1(n5130), .A2(n5129), .ZN(n5131) );
  AND2_X1 U6470 ( .A1(n5158), .A2(n5131), .ZN(n8072) );
  NAND2_X1 U6471 ( .A1(n5413), .A2(n8072), .ZN(n5135) );
  NAND2_X1 U6472 ( .A1(n5056), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5134) );
  NAND2_X1 U6473 ( .A1(n6317), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5133) );
  NAND2_X1 U6474 ( .A1(n6343), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5132) );
  NAND4_X1 U6475 ( .A1(n5135), .A2(n5134), .A3(n5133), .A4(n5132), .ZN(n9047)
         );
  NAND2_X1 U6476 ( .A1(n9047), .A2(n5602), .ZN(n5136) );
  NAND2_X1 U6477 ( .A1(n5137), .A2(n5136), .ZN(n5138) );
  XNOR2_X1 U6478 ( .A(n5138), .B(n4976), .ZN(n5140) );
  AND2_X1 U6479 ( .A1(n9047), .A2(n5601), .ZN(n5139) );
  AOI21_X1 U6480 ( .B1(n9886), .B2(n5602), .A(n5139), .ZN(n5141) );
  NAND2_X1 U6481 ( .A1(n5140), .A2(n5141), .ZN(n5146) );
  INV_X1 U6482 ( .A(n5140), .ZN(n5143) );
  INV_X1 U6483 ( .A(n5141), .ZN(n5142) );
  NAND2_X1 U6484 ( .A1(n5143), .A2(n5142), .ZN(n5144) );
  NAND2_X1 U6485 ( .A1(n5146), .A2(n5144), .ZN(n7530) );
  INV_X1 U6486 ( .A(n7530), .ZN(n5145) );
  INV_X1 U6487 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6682) );
  INV_X1 U6488 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5149) );
  MUX2_X1 U6489 ( .A(n6682), .B(n5149), .S(n5700), .Z(n5151) );
  INV_X1 U6490 ( .A(SI_10_), .ZN(n5150) );
  INV_X1 U6491 ( .A(n5151), .ZN(n5152) );
  NAND2_X1 U6492 ( .A1(n5152), .A2(SI_10_), .ZN(n5153) );
  XNOR2_X1 U6493 ( .A(n5170), .B(n4823), .ZN(n6664) );
  NAND2_X1 U6494 ( .A1(n6664), .A2(n5009), .ZN(n5156) );
  NAND2_X1 U6495 ( .A1(n5174), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5154) );
  XNOR2_X1 U6496 ( .A(n5154), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9826) );
  AOI22_X1 U6497 ( .A1(n6340), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n4988), .B2(
        n9826), .ZN(n5155) );
  NAND2_X1 U6498 ( .A1(n9671), .A2(n5586), .ZN(n5165) );
  NAND2_X1 U6499 ( .A1(n6344), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5163) );
  NAND2_X1 U6500 ( .A1(n6317), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5162) );
  INV_X1 U6501 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U6502 ( .A1(n5158), .A2(n5157), .ZN(n5159) );
  AND2_X1 U6503 ( .A1(n5179), .A2(n5159), .ZN(n8062) );
  NAND2_X1 U6504 ( .A1(n5413), .A2(n8062), .ZN(n5161) );
  NAND2_X1 U6505 ( .A1(n5209), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5160) );
  OR2_X1 U6506 ( .A1(n9713), .A2(n5596), .ZN(n5164) );
  NAND2_X1 U6507 ( .A1(n5165), .A2(n5164), .ZN(n5166) );
  XNOR2_X1 U6508 ( .A(n5166), .B(n4976), .ZN(n5169) );
  NOR2_X1 U6509 ( .A1(n9713), .A2(n5026), .ZN(n5167) );
  AOI21_X1 U6510 ( .B1(n9671), .B2(n5602), .A(n5167), .ZN(n5168) );
  OR2_X1 U6511 ( .A1(n5169), .A2(n5168), .ZN(n8059) );
  NAND2_X1 U6512 ( .A1(n5170), .A2(n4823), .ZN(n5172) );
  INV_X1 U6513 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6684) );
  INV_X1 U6514 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5173) );
  MUX2_X1 U6515 ( .A(n6684), .B(n5173), .S(n5700), .Z(n5194) );
  XNOR2_X1 U6516 ( .A(n5198), .B(n5193), .ZN(n6666) );
  NAND2_X1 U6517 ( .A1(n6666), .A2(n5009), .ZN(n5177) );
  OAI21_X1 U6518 ( .B1(n5174), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5175) );
  XNOR2_X1 U6519 ( .A(n5175), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6982) );
  AOI22_X1 U6520 ( .A1(n6340), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n4988), .B2(
        n6982), .ZN(n5176) );
  NAND2_X1 U6521 ( .A1(n5177), .A2(n5176), .ZN(n7753) );
  NAND2_X1 U6522 ( .A1(n7753), .A2(n5586), .ZN(n5186) );
  NAND2_X1 U6523 ( .A1(n5209), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U6524 ( .A1(n6344), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5183) );
  INV_X1 U6525 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5178) );
  AND2_X1 U6526 ( .A1(n5179), .A2(n5178), .ZN(n5180) );
  NOR2_X1 U6527 ( .A1(n5211), .A2(n5180), .ZN(n9721) );
  NAND2_X1 U6528 ( .A1(n5413), .A2(n9721), .ZN(n5182) );
  NAND2_X1 U6529 ( .A1(n6317), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5181) );
  NAND4_X1 U6530 ( .A1(n5184), .A2(n5183), .A3(n5182), .A4(n5181), .ZN(n9045)
         );
  NAND2_X1 U6531 ( .A1(n9045), .A2(n5602), .ZN(n5185) );
  NAND2_X1 U6532 ( .A1(n5186), .A2(n5185), .ZN(n5187) );
  XNOR2_X1 U6533 ( .A(n5187), .B(n5599), .ZN(n5191) );
  AND2_X1 U6534 ( .A1(n9045), .A2(n5601), .ZN(n5188) );
  AOI21_X1 U6535 ( .B1(n7753), .B2(n5602), .A(n5188), .ZN(n5189) );
  XNOR2_X1 U6536 ( .A(n5191), .B(n5189), .ZN(n7695) );
  INV_X1 U6537 ( .A(n5189), .ZN(n5190) );
  NAND2_X1 U6538 ( .A1(n5191), .A2(n5190), .ZN(n5192) );
  NAND2_X1 U6539 ( .A1(n7694), .A2(n5192), .ZN(n7776) );
  INV_X1 U6540 ( .A(n5194), .ZN(n5195) );
  NAND2_X1 U6541 ( .A1(n5195), .A2(SI_11_), .ZN(n5196) );
  INV_X1 U6542 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5200) );
  INV_X1 U6543 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5199) );
  MUX2_X1 U6544 ( .A(n5200), .B(n5199), .S(n5700), .Z(n5202) );
  INV_X1 U6545 ( .A(SI_12_), .ZN(n5201) );
  INV_X1 U6546 ( .A(n5202), .ZN(n5203) );
  NAND2_X1 U6547 ( .A1(n5203), .A2(SI_12_), .ZN(n5204) );
  NAND2_X1 U6548 ( .A1(n6698), .A2(n5009), .ZN(n5208) );
  OR2_X1 U6549 ( .A1(n5205), .A2(n5122), .ZN(n5206) );
  XNOR2_X1 U6550 ( .A(n5206), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7166) );
  AOI22_X1 U6551 ( .A1(n6340), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n4988), .B2(
        n7166), .ZN(n5207) );
  NAND2_X1 U6552 ( .A1(n7816), .A2(n5586), .ZN(n5218) );
  NAND2_X1 U6553 ( .A1(n5209), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U6554 ( .A1(n6344), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5215) );
  OR2_X1 U6555 ( .A1(n5211), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5212) );
  NAND2_X1 U6556 ( .A1(n5211), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5236) );
  AND2_X1 U6557 ( .A1(n5212), .A2(n5236), .ZN(n7777) );
  NAND2_X1 U6558 ( .A1(n5591), .A2(n7777), .ZN(n5214) );
  NAND2_X1 U6559 ( .A1(n6317), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5213) );
  OR2_X1 U6560 ( .A1(n9711), .A2(n5596), .ZN(n5217) );
  NAND2_X1 U6561 ( .A1(n5218), .A2(n5217), .ZN(n5219) );
  XNOR2_X1 U6562 ( .A(n5219), .B(n4976), .ZN(n7774) );
  NOR2_X1 U6563 ( .A1(n9711), .A2(n5026), .ZN(n5220) );
  AOI21_X1 U6564 ( .B1(n7816), .B2(n5602), .A(n5220), .ZN(n5222) );
  NAND2_X1 U6565 ( .A1(n7774), .A2(n5222), .ZN(n5221) );
  INV_X1 U6566 ( .A(n7774), .ZN(n5223) );
  INV_X1 U6567 ( .A(n5222), .ZN(n7773) );
  NAND2_X1 U6568 ( .A1(n5223), .A2(n7773), .ZN(n5224) );
  INV_X1 U6569 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6751) );
  INV_X1 U6570 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5227) );
  MUX2_X1 U6571 ( .A(n6751), .B(n5227), .S(n5700), .Z(n5229) );
  INV_X1 U6572 ( .A(SI_13_), .ZN(n5228) );
  NAND2_X1 U6573 ( .A1(n5229), .A2(n5228), .ZN(n5251) );
  INV_X1 U6574 ( .A(n5229), .ZN(n5230) );
  NAND2_X1 U6575 ( .A1(n5230), .A2(SI_13_), .ZN(n5231) );
  XNOR2_X1 U6576 ( .A(n5250), .B(n5249), .ZN(n6744) );
  NAND2_X1 U6577 ( .A1(n6744), .A2(n5009), .ZN(n5234) );
  NAND2_X1 U6578 ( .A1(n4857), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5232) );
  XNOR2_X1 U6579 ( .A(n5232), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7465) );
  AOI22_X1 U6580 ( .A1(n6340), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n4988), .B2(
        n7465), .ZN(n5233) );
  NAND2_X1 U6581 ( .A1(n6344), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U6582 ( .A1(n6343), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5240) );
  INV_X1 U6583 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U6584 ( .A1(n5236), .A2(n5235), .ZN(n5237) );
  AND2_X1 U6585 ( .A1(n5260), .A2(n5237), .ZN(n7916) );
  NAND2_X1 U6586 ( .A1(n5413), .A2(n7916), .ZN(n5239) );
  NAND2_X1 U6587 ( .A1(n5084), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5238) );
  OAI22_X1 U6588 ( .A1(n9729), .A2(n5499), .B1(n8040), .B2(n5596), .ZN(n5242)
         );
  XNOR2_X1 U6589 ( .A(n5242), .B(n5599), .ZN(n5245) );
  OR2_X1 U6590 ( .A1(n9729), .A2(n5596), .ZN(n5244) );
  OR2_X1 U6591 ( .A1(n8040), .A2(n5026), .ZN(n5243) );
  NAND2_X1 U6592 ( .A1(n5244), .A2(n5243), .ZN(n5246) );
  AND2_X1 U6593 ( .A1(n5245), .A2(n5246), .ZN(n7910) );
  INV_X1 U6594 ( .A(n5245), .ZN(n5248) );
  INV_X1 U6595 ( .A(n5246), .ZN(n5247) );
  NAND2_X1 U6596 ( .A1(n5248), .A2(n5247), .ZN(n7908) );
  INV_X1 U6597 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6753) );
  INV_X1 U6598 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5252) );
  MUX2_X1 U6599 ( .A(n6753), .B(n5252), .S(n5700), .Z(n5271) );
  XNOR2_X1 U6600 ( .A(n5271), .B(SI_14_), .ZN(n5270) );
  XNOR2_X1 U6601 ( .A(n5275), .B(n5270), .ZN(n6746) );
  NAND2_X1 U6602 ( .A1(n6746), .A2(n5009), .ZN(n5258) );
  NAND2_X1 U6603 ( .A1(n5253), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5255) );
  NAND2_X1 U6604 ( .A1(n5255), .A2(n5254), .ZN(n5281) );
  OR2_X1 U6605 ( .A1(n5255), .A2(n5254), .ZN(n5256) );
  AND2_X1 U6606 ( .A1(n5281), .A2(n5256), .ZN(n7686) );
  AOI22_X1 U6607 ( .A1(n6340), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n4988), .B2(
        n7686), .ZN(n5257) );
  NAND2_X1 U6608 ( .A1(n6344), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U6609 ( .A1(n6343), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5264) );
  INV_X1 U6610 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5259) );
  AND2_X1 U6611 ( .A1(n5260), .A2(n5259), .ZN(n5261) );
  NOR2_X1 U6612 ( .A1(n5286), .A2(n5261), .ZN(n8037) );
  NAND2_X1 U6613 ( .A1(n5591), .A2(n8037), .ZN(n5263) );
  NAND2_X1 U6614 ( .A1(n6317), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5262) );
  OAI22_X1 U6615 ( .A1(n7973), .A2(n5499), .B1(n9690), .B2(n5596), .ZN(n5266)
         );
  XNOR2_X1 U6616 ( .A(n5266), .B(n4976), .ZN(n5269) );
  OR2_X1 U6617 ( .A1(n7973), .A2(n5596), .ZN(n5268) );
  OR2_X1 U6618 ( .A1(n9690), .A2(n5026), .ZN(n5267) );
  NAND2_X1 U6619 ( .A1(n5268), .A2(n5267), .ZN(n8042) );
  INV_X1 U6620 ( .A(n5270), .ZN(n5274) );
  INV_X1 U6621 ( .A(n5271), .ZN(n5272) );
  NAND2_X1 U6622 ( .A1(n5272), .A2(SI_14_), .ZN(n5273) );
  INV_X1 U6623 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6991) );
  INV_X1 U6624 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n5276) );
  MUX2_X1 U6625 ( .A(n6991), .B(n5276), .S(n5700), .Z(n5278) );
  INV_X1 U6626 ( .A(SI_15_), .ZN(n5277) );
  NAND2_X1 U6627 ( .A1(n5278), .A2(n5277), .ZN(n5297) );
  INV_X1 U6628 ( .A(n5278), .ZN(n5279) );
  NAND2_X1 U6629 ( .A1(n5279), .A2(SI_15_), .ZN(n5280) );
  NAND2_X1 U6630 ( .A1(n5297), .A2(n5280), .ZN(n5298) );
  XNOR2_X1 U6631 ( .A(n5299), .B(n5298), .ZN(n6876) );
  NAND2_X1 U6632 ( .A1(n6876), .A2(n5009), .ZN(n5285) );
  NAND2_X1 U6633 ( .A1(n5281), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5283) );
  XNOR2_X1 U6634 ( .A(n5283), .B(n5282), .ZN(n7929) );
  INV_X1 U6635 ( .A(n7929), .ZN(n7690) );
  AOI22_X1 U6636 ( .A1(n6340), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n4988), .B2(
        n7690), .ZN(n5284) );
  NAND2_X1 U6637 ( .A1(n6344), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6638 ( .A1(n6317), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5290) );
  NOR2_X1 U6639 ( .A1(n5286), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5287) );
  NAND2_X1 U6640 ( .A1(n5413), .A2(n4830), .ZN(n5289) );
  NAND2_X1 U6641 ( .A1(n6343), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5288) );
  OAI22_X1 U6642 ( .A1(n8016), .A2(n5499), .B1(n7976), .B2(n5596), .ZN(n5292)
         );
  XNOR2_X1 U6643 ( .A(n5292), .B(n4976), .ZN(n5293) );
  OAI22_X1 U6644 ( .A1(n8016), .A2(n5596), .B1(n7976), .B2(n5026), .ZN(n8030)
         );
  NAND2_X1 U6645 ( .A1(n8027), .A2(n8030), .ZN(n5296) );
  NAND2_X1 U6646 ( .A1(n8041), .A2(n8045), .ZN(n5295) );
  INV_X1 U6647 ( .A(n5293), .ZN(n5294) );
  NAND2_X1 U6648 ( .A1(n5295), .A2(n5294), .ZN(n8028) );
  NAND2_X1 U6649 ( .A1(n5296), .A2(n8028), .ZN(n8948) );
  INV_X1 U6650 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5301) );
  INV_X1 U6651 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5300) );
  MUX2_X1 U6652 ( .A(n5301), .B(n5300), .S(n5327), .Z(n5303) );
  INV_X1 U6653 ( .A(SI_16_), .ZN(n5302) );
  NAND2_X1 U6654 ( .A1(n5303), .A2(n5302), .ZN(n5326) );
  INV_X1 U6655 ( .A(n5303), .ZN(n5304) );
  NAND2_X1 U6656 ( .A1(n5304), .A2(SI_16_), .ZN(n5305) );
  XNOR2_X1 U6657 ( .A(n5325), .B(n5324), .ZN(n6926) );
  NAND2_X1 U6658 ( .A1(n6926), .A2(n5009), .ZN(n5309) );
  OR2_X1 U6659 ( .A1(n5306), .A2(n5122), .ZN(n5307) );
  XNOR2_X1 U6660 ( .A(n5307), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9078) );
  AOI22_X1 U6661 ( .A1(n6340), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n4988), .B2(
        n9078), .ZN(n5308) );
  NAND2_X1 U6662 ( .A1(n6343), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6663 ( .A1(n6344), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6664 ( .A1(n5310), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5336) );
  OR2_X1 U6665 ( .A1(n5310), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5311) );
  AND2_X1 U6666 ( .A1(n5336), .A2(n5311), .ZN(n8951) );
  NAND2_X1 U6667 ( .A1(n5591), .A2(n8951), .ZN(n5313) );
  NAND2_X1 U6668 ( .A1(n6317), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5312) );
  NAND4_X1 U6669 ( .A1(n5315), .A2(n5314), .A3(n5313), .A4(n5312), .ZN(n9348)
         );
  INV_X1 U6670 ( .A(n9348), .ZN(n8033) );
  OAI22_X1 U6671 ( .A1(n8950), .A2(n5499), .B1(n8033), .B2(n5596), .ZN(n5316)
         );
  XNOR2_X1 U6672 ( .A(n5316), .B(n5599), .ZN(n5319) );
  OR2_X1 U6673 ( .A1(n8950), .A2(n5596), .ZN(n5318) );
  NAND2_X1 U6674 ( .A1(n9348), .A2(n5601), .ZN(n5317) );
  NAND2_X1 U6675 ( .A1(n5318), .A2(n5317), .ZN(n5320) );
  XNOR2_X1 U6676 ( .A(n5319), .B(n5320), .ZN(n8949) );
  INV_X1 U6677 ( .A(n5319), .ZN(n5322) );
  INV_X1 U6678 ( .A(n5320), .ZN(n5321) );
  NAND2_X1 U6679 ( .A1(n5322), .A2(n5321), .ZN(n5323) );
  INV_X1 U6680 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9602) );
  INV_X1 U6681 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5328) );
  MUX2_X1 U6682 ( .A(n9602), .B(n5328), .S(n5327), .Z(n5352) );
  XNOR2_X1 U6683 ( .A(n5352), .B(SI_17_), .ZN(n5351) );
  XNOR2_X1 U6684 ( .A(n5371), .B(n5351), .ZN(n7103) );
  NAND2_X1 U6685 ( .A1(n7103), .A2(n5009), .ZN(n5334) );
  NAND2_X1 U6686 ( .A1(n5329), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6687 ( .A1(n5331), .A2(n5330), .ZN(n5356) );
  OR2_X1 U6688 ( .A1(n5331), .A2(n5330), .ZN(n5332) );
  AND2_X1 U6689 ( .A1(n5356), .A2(n5332), .ZN(n9093) );
  AOI22_X1 U6690 ( .A1(n6340), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n4988), .B2(
        n9093), .ZN(n5333) );
  NAND2_X1 U6691 ( .A1(n9428), .A2(n5586), .ZN(n5343) );
  NAND2_X1 U6692 ( .A1(n6343), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U6693 ( .A1(n6344), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5340) );
  INV_X1 U6694 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U6695 ( .A1(n5336), .A2(n5335), .ZN(n5337) );
  AND2_X1 U6696 ( .A1(n5361), .A2(n5337), .ZN(n9343) );
  NAND2_X1 U6697 ( .A1(n5413), .A2(n9343), .ZN(n5339) );
  NAND2_X1 U6698 ( .A1(n6317), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5338) );
  NAND4_X1 U6699 ( .A1(n5341), .A2(n5340), .A3(n5339), .A4(n5338), .ZN(n9333)
         );
  NAND2_X1 U6700 ( .A1(n9333), .A2(n5602), .ZN(n5342) );
  NAND2_X1 U6701 ( .A1(n5343), .A2(n5342), .ZN(n5344) );
  XNOR2_X1 U6702 ( .A(n5344), .B(n5599), .ZN(n5346) );
  AND2_X1 U6703 ( .A1(n9333), .A2(n5601), .ZN(n5345) );
  AOI21_X1 U6704 ( .B1(n9428), .B2(n5602), .A(n5345), .ZN(n5347) );
  XNOR2_X1 U6705 ( .A(n5346), .B(n5347), .ZN(n8957) );
  INV_X1 U6706 ( .A(n5346), .ZN(n5348) );
  NAND2_X1 U6707 ( .A1(n5348), .A2(n5347), .ZN(n5349) );
  NAND2_X1 U6708 ( .A1(n5350), .A2(n5349), .ZN(n9007) );
  INV_X1 U6709 ( .A(n5351), .ZN(n5369) );
  OR2_X1 U6710 ( .A1(n5371), .A2(n5369), .ZN(n5354) );
  INV_X1 U6711 ( .A(n5352), .ZN(n5353) );
  NAND2_X1 U6712 ( .A1(n5353), .A2(SI_17_), .ZN(n5372) );
  MUX2_X1 U6713 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5700), .Z(n5374) );
  XNOR2_X1 U6714 ( .A(n5374), .B(SI_18_), .ZN(n5373) );
  NAND2_X1 U6715 ( .A1(n7206), .A2(n5009), .ZN(n5359) );
  NAND2_X1 U6716 ( .A1(n5356), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5357) );
  XNOR2_X1 U6717 ( .A(n5357), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9103) );
  AOI22_X1 U6718 ( .A1(n6340), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9103), .B2(
        n4988), .ZN(n5358) );
  NAND2_X1 U6719 ( .A1(n9423), .A2(n5586), .ZN(n5366) );
  INV_X1 U6720 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5360) );
  AND2_X1 U6721 ( .A1(n5361), .A2(n5360), .ZN(n5362) );
  OR2_X1 U6722 ( .A1(n5362), .A2(n5386), .ZN(n9325) );
  AOI22_X1 U6723 ( .A1(n6317), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n6344), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U6724 ( .A1(n6343), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5363) );
  OAI211_X1 U6725 ( .C1(n9325), .C2(n5210), .A(n5364), .B(n5363), .ZN(n9350)
         );
  NAND2_X1 U6726 ( .A1(n9350), .A2(n5602), .ZN(n5365) );
  NAND2_X1 U6727 ( .A1(n5366), .A2(n5365), .ZN(n5367) );
  XNOR2_X1 U6728 ( .A(n5367), .B(n4976), .ZN(n9005) );
  AND2_X1 U6729 ( .A1(n9350), .A2(n5601), .ZN(n5368) );
  AOI21_X1 U6730 ( .B1(n9423), .B2(n5602), .A(n5368), .ZN(n9004) );
  NAND2_X1 U6731 ( .A1(n5374), .A2(SI_18_), .ZN(n5375) );
  INV_X1 U6732 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7345) );
  INV_X1 U6733 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n5378) );
  MUX2_X1 U6734 ( .A(n7345), .B(n5378), .S(n5700), .Z(n5380) );
  INV_X1 U6735 ( .A(SI_19_), .ZN(n5379) );
  NAND2_X1 U6736 ( .A1(n5380), .A2(n5379), .ZN(n5402) );
  INV_X1 U6737 ( .A(n5380), .ZN(n5381) );
  NAND2_X1 U6738 ( .A1(n5381), .A2(SI_19_), .ZN(n5382) );
  NAND2_X1 U6739 ( .A1(n5402), .A2(n5382), .ZN(n5399) );
  XNOR2_X1 U6740 ( .A(n5398), .B(n5399), .ZN(n7290) );
  NAND2_X1 U6741 ( .A1(n7290), .A2(n5009), .ZN(n5385) );
  AOI22_X1 U6742 ( .A1(n6340), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9110), .B2(
        n4988), .ZN(n5384) );
  NAND2_X1 U6743 ( .A1(n9419), .A2(n5586), .ZN(n5391) );
  NOR2_X1 U6744 ( .A1(n5386), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5387) );
  OR2_X1 U6745 ( .A1(n5411), .A2(n5387), .ZN(n9318) );
  AOI22_X1 U6746 ( .A1(n6343), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n6344), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U6747 ( .A1(n6317), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5388) );
  OAI211_X1 U6748 ( .C1(n9318), .C2(n5210), .A(n5389), .B(n5388), .ZN(n9334)
         );
  NAND2_X1 U6749 ( .A1(n9334), .A2(n5602), .ZN(n5390) );
  NAND2_X1 U6750 ( .A1(n5391), .A2(n5390), .ZN(n5392) );
  XNOR2_X1 U6751 ( .A(n5392), .B(n5599), .ZN(n5394) );
  AND2_X1 U6752 ( .A1(n9334), .A2(n5601), .ZN(n5393) );
  AOI21_X1 U6753 ( .B1(n9419), .B2(n5602), .A(n5393), .ZN(n5395) );
  XNOR2_X1 U6754 ( .A(n5394), .B(n5395), .ZN(n8914) );
  INV_X1 U6755 ( .A(n5394), .ZN(n5396) );
  NAND2_X1 U6756 ( .A1(n5396), .A2(n5395), .ZN(n5397) );
  INV_X1 U6757 ( .A(n5398), .ZN(n5401) );
  INV_X1 U6758 ( .A(n5399), .ZN(n5400) );
  INV_X1 U6759 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7457) );
  INV_X1 U6760 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n5404) );
  MUX2_X1 U6761 ( .A(n7457), .B(n5404), .S(n5700), .Z(n5406) );
  INV_X1 U6762 ( .A(SI_20_), .ZN(n5405) );
  NAND2_X1 U6763 ( .A1(n5406), .A2(n5405), .ZN(n5430) );
  INV_X1 U6764 ( .A(n5406), .ZN(n5407) );
  NAND2_X1 U6765 ( .A1(n5407), .A2(SI_20_), .ZN(n5408) );
  XNOR2_X1 U6766 ( .A(n5429), .B(n5428), .ZN(n7452) );
  NAND2_X1 U6767 ( .A1(n7452), .A2(n5009), .ZN(n5410) );
  NAND2_X1 U6768 ( .A1(n6340), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5409) );
  NAND2_X1 U6769 ( .A1(n9414), .A2(n5586), .ZN(n5421) );
  OR2_X1 U6770 ( .A1(n5411), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5412) );
  AND2_X1 U6771 ( .A1(n5412), .A2(n5435), .ZN(n9297) );
  NAND2_X1 U6772 ( .A1(n9297), .A2(n5413), .ZN(n5419) );
  INV_X1 U6773 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U6774 ( .A1(n6344), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U6775 ( .A1(n6317), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5414) );
  OAI211_X1 U6776 ( .C1(n6321), .C2(n5416), .A(n5415), .B(n5414), .ZN(n5417)
         );
  INV_X1 U6777 ( .A(n5417), .ZN(n5418) );
  NAND2_X1 U6778 ( .A1(n5419), .A2(n5418), .ZN(n9312) );
  NAND2_X1 U6779 ( .A1(n9312), .A2(n5602), .ZN(n5420) );
  NAND2_X1 U6780 ( .A1(n5421), .A2(n5420), .ZN(n5422) );
  XNOR2_X1 U6781 ( .A(n5422), .B(n5599), .ZN(n5424) );
  AND2_X1 U6782 ( .A1(n9312), .A2(n5601), .ZN(n5423) );
  AOI21_X1 U6783 ( .B1(n9414), .B2(n5602), .A(n5423), .ZN(n5425) );
  XNOR2_X1 U6784 ( .A(n5424), .B(n5425), .ZN(n8986) );
  INV_X1 U6785 ( .A(n5424), .ZN(n5426) );
  NAND2_X1 U6786 ( .A1(n5426), .A2(n5425), .ZN(n5427) );
  NAND2_X1 U6787 ( .A1(n5429), .A2(n5428), .ZN(n5431) );
  INV_X1 U6788 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7495) );
  INV_X1 U6789 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n5432) );
  XNOR2_X1 U6790 ( .A(n5451), .B(SI_21_), .ZN(n5450) );
  XNOR2_X1 U6791 ( .A(n5449), .B(n5450), .ZN(n7471) );
  NAND2_X1 U6792 ( .A1(n7471), .A2(n5009), .ZN(n5434) );
  NAND2_X1 U6793 ( .A1(n6340), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U6794 ( .A1(n9409), .A2(n5586), .ZN(n5441) );
  NAND2_X1 U6795 ( .A1(n6343), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U6796 ( .A1(n6344), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5438) );
  INV_X1 U6797 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8933) );
  AOI21_X1 U6798 ( .B1(n8933), .B2(n5435), .A(n5461), .ZN(n9289) );
  NAND2_X1 U6799 ( .A1(n5591), .A2(n9289), .ZN(n5437) );
  NAND2_X1 U6800 ( .A1(n6317), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5436) );
  OR2_X1 U6801 ( .A1(n9041), .A2(n5596), .ZN(n5440) );
  NAND2_X1 U6802 ( .A1(n5441), .A2(n5440), .ZN(n5442) );
  XNOR2_X1 U6803 ( .A(n5442), .B(n5599), .ZN(n5444) );
  NOR2_X1 U6804 ( .A1(n9041), .A2(n5026), .ZN(n5443) );
  AOI21_X1 U6805 ( .B1(n9409), .B2(n5602), .A(n5443), .ZN(n5445) );
  XNOR2_X1 U6806 ( .A(n5444), .B(n5445), .ZN(n8932) );
  INV_X1 U6807 ( .A(n5444), .ZN(n5446) );
  NAND2_X1 U6808 ( .A1(n5446), .A2(n5445), .ZN(n5447) );
  INV_X1 U6809 ( .A(n5451), .ZN(n5452) );
  NAND2_X1 U6810 ( .A1(n5452), .A2(SI_21_), .ZN(n5453) );
  INV_X1 U6811 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8196) );
  INV_X1 U6812 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n5454) );
  MUX2_X1 U6813 ( .A(n8196), .B(n5454), .S(n5700), .Z(n5456) );
  INV_X1 U6814 ( .A(SI_22_), .ZN(n5455) );
  NAND2_X1 U6815 ( .A1(n5456), .A2(n5455), .ZN(n5469) );
  INV_X1 U6816 ( .A(n5456), .ZN(n5457) );
  NAND2_X1 U6817 ( .A1(n5457), .A2(SI_22_), .ZN(n5458) );
  NAND2_X1 U6818 ( .A1(n5469), .A2(n5458), .ZN(n5470) );
  XNOR2_X1 U6819 ( .A(n5471), .B(n5470), .ZN(n7537) );
  NAND2_X1 U6820 ( .A1(n7537), .A2(n5009), .ZN(n5460) );
  NAND2_X1 U6821 ( .A1(n6340), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U6822 ( .A1(n6343), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U6823 ( .A1(n6344), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U6824 ( .A1(n5461), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5480) );
  OAI21_X1 U6825 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n5461), .A(n5480), .ZN(
        n8999) );
  INV_X1 U6826 ( .A(n8999), .ZN(n9274) );
  NAND2_X1 U6827 ( .A1(n5413), .A2(n9274), .ZN(n5463) );
  NAND2_X1 U6828 ( .A1(n6317), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5462) );
  NAND4_X1 U6829 ( .A1(n5465), .A2(n5464), .A3(n5463), .A4(n5462), .ZN(n9286)
         );
  AND2_X1 U6830 ( .A1(n9286), .A2(n5601), .ZN(n5466) );
  AOI21_X1 U6831 ( .B1(n9404), .B2(n5602), .A(n5466), .ZN(n5467) );
  INV_X1 U6832 ( .A(n9286), .ZN(n9130) );
  OAI22_X1 U6833 ( .A1(n9268), .A2(n5499), .B1(n9130), .B2(n5596), .ZN(n5468)
         );
  XNOR2_X1 U6834 ( .A(n5468), .B(n5599), .ZN(n8994) );
  INV_X1 U6835 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5473) );
  INV_X1 U6836 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5472) );
  MUX2_X1 U6837 ( .A(n5473), .B(n5472), .S(n5700), .Z(n5475) );
  INV_X1 U6838 ( .A(SI_23_), .ZN(n5474) );
  NAND2_X1 U6839 ( .A1(n5475), .A2(n5474), .ZN(n5489) );
  INV_X1 U6840 ( .A(n5475), .ZN(n5476) );
  NAND2_X1 U6841 ( .A1(n5476), .A2(SI_23_), .ZN(n5477) );
  AND2_X1 U6842 ( .A1(n5489), .A2(n5477), .ZN(n5487) );
  XNOR2_X1 U6843 ( .A(n5488), .B(n5487), .ZN(n7701) );
  NAND2_X1 U6844 ( .A1(n7701), .A2(n5009), .ZN(n5479) );
  NAND2_X1 U6845 ( .A1(n6340), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U6846 ( .A1(n6343), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U6847 ( .A1(n6344), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5483) );
  INV_X1 U6848 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8907) );
  AOI21_X1 U6849 ( .B1(n8907), .B2(n5480), .A(n5494), .ZN(n9256) );
  NAND2_X1 U6850 ( .A1(n5591), .A2(n9256), .ZN(n5482) );
  NAND2_X1 U6851 ( .A1(n6317), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5481) );
  OAI22_X1 U6852 ( .A1(n9258), .A2(n5499), .B1(n9131), .B2(n5596), .ZN(n5485)
         );
  XNOR2_X1 U6853 ( .A(n5485), .B(n5599), .ZN(n5486) );
  INV_X1 U6854 ( .A(n9131), .ZN(n9271) );
  AOI22_X1 U6855 ( .A1(n9399), .A2(n5602), .B1(n5601), .B2(n9271), .ZN(n8905)
         );
  NAND2_X1 U6856 ( .A1(n8993), .A2(n5486), .ZN(n8903) );
  OAI21_X2 U6857 ( .B1(n8902), .B2(n8905), .A(n8903), .ZN(n8964) );
  INV_X1 U6858 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7811) );
  INV_X1 U6859 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n5491) );
  MUX2_X1 U6860 ( .A(n7811), .B(n5491), .S(n5700), .Z(n5504) );
  XNOR2_X1 U6861 ( .A(n5504), .B(SI_24_), .ZN(n5503) );
  NAND2_X1 U6862 ( .A1(n7783), .A2(n5009), .ZN(n5493) );
  NAND2_X1 U6863 ( .A1(n6340), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U6864 ( .A1(n6344), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U6865 ( .A1(n6317), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U6866 ( .A1(n5494), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5516) );
  OAI21_X1 U6867 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n5494), .A(n5516), .ZN(
        n8967) );
  INV_X1 U6868 ( .A(n8967), .ZN(n9248) );
  NAND2_X1 U6869 ( .A1(n5413), .A2(n9248), .ZN(n5496) );
  NAND2_X1 U6870 ( .A1(n6343), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5495) );
  OAI22_X1 U6871 ( .A1(n9240), .A2(n5499), .B1(n9259), .B2(n5596), .ZN(n5500)
         );
  XNOR2_X1 U6872 ( .A(n5500), .B(n5599), .ZN(n5501) );
  OAI22_X1 U6873 ( .A1(n9240), .A2(n5596), .B1(n9259), .B2(n5026), .ZN(n5502)
         );
  XNOR2_X1 U6874 ( .A(n5501), .B(n5502), .ZN(n8965) );
  INV_X1 U6875 ( .A(n5503), .ZN(n5507) );
  INV_X1 U6876 ( .A(n5504), .ZN(n5505) );
  NAND2_X1 U6877 ( .A1(n5505), .A2(SI_24_), .ZN(n5506) );
  INV_X1 U6878 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7947) );
  INV_X1 U6879 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n5509) );
  MUX2_X1 U6880 ( .A(n7947), .B(n5509), .S(n5700), .Z(n5511) );
  INV_X1 U6881 ( .A(SI_25_), .ZN(n5510) );
  NAND2_X1 U6882 ( .A1(n5511), .A2(n5510), .ZN(n5530) );
  INV_X1 U6883 ( .A(n5511), .ZN(n5512) );
  NAND2_X1 U6884 ( .A1(n5512), .A2(SI_25_), .ZN(n5513) );
  NAND2_X1 U6885 ( .A1(n5530), .A2(n5513), .ZN(n5531) );
  NAND2_X1 U6886 ( .A1(n7939), .A2(n5009), .ZN(n5515) );
  NAND2_X1 U6887 ( .A1(n6340), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U6888 ( .A1(n6344), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U6889 ( .A1(n5084), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5521) );
  INV_X1 U6890 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9583) );
  NAND2_X1 U6891 ( .A1(n9583), .A2(n5516), .ZN(n5518) );
  INV_X1 U6892 ( .A(n5516), .ZN(n5517) );
  NAND2_X1 U6893 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n5517), .ZN(n5541) );
  AND2_X1 U6894 ( .A1(n5518), .A2(n5541), .ZN(n9234) );
  NAND2_X1 U6895 ( .A1(n5591), .A2(n9234), .ZN(n5520) );
  NAND2_X1 U6896 ( .A1(n6343), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5519) );
  OAI22_X1 U6897 ( .A1(n9223), .A2(n5596), .B1(n9135), .B2(n5026), .ZN(n5527)
         );
  NAND2_X1 U6898 ( .A1(n9389), .A2(n5586), .ZN(n5524) );
  OR2_X1 U6899 ( .A1(n9135), .A2(n5596), .ZN(n5523) );
  NAND2_X1 U6900 ( .A1(n5524), .A2(n5523), .ZN(n5525) );
  XNOR2_X1 U6901 ( .A(n5525), .B(n5599), .ZN(n5526) );
  XOR2_X1 U6902 ( .A(n5527), .B(n5526), .Z(n8940) );
  INV_X1 U6903 ( .A(n5526), .ZN(n5529) );
  INV_X1 U6904 ( .A(n5527), .ZN(n5528) );
  INV_X1 U6905 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7948) );
  INV_X1 U6906 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5533) );
  MUX2_X1 U6907 ( .A(n7948), .B(n5533), .S(n4299), .Z(n5535) );
  INV_X1 U6908 ( .A(SI_26_), .ZN(n5534) );
  NAND2_X1 U6909 ( .A1(n5535), .A2(n5534), .ZN(n5554) );
  INV_X1 U6910 ( .A(n5535), .ZN(n5536) );
  NAND2_X1 U6911 ( .A1(n5536), .A2(SI_26_), .ZN(n5537) );
  AND2_X1 U6912 ( .A1(n5554), .A2(n5537), .ZN(n5552) );
  NAND2_X1 U6913 ( .A1(n6340), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U6914 ( .A1(n6343), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U6915 ( .A1(n6344), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5545) );
  INV_X1 U6916 ( .A(n5541), .ZN(n5540) );
  NAND2_X1 U6917 ( .A1(n5540), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5564) );
  INV_X1 U6918 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9031) );
  NAND2_X1 U6919 ( .A1(n5541), .A2(n9031), .ZN(n5542) );
  AND2_X1 U6920 ( .A1(n5564), .A2(n5542), .ZN(n9215) );
  NAND2_X1 U6921 ( .A1(n5591), .A2(n9215), .ZN(n5544) );
  NAND2_X1 U6922 ( .A1(n6317), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5543) );
  NAND4_X1 U6923 ( .A1(n5546), .A2(n5545), .A3(n5544), .A4(n5543), .ZN(n9203)
         );
  AOI22_X1 U6924 ( .A1(n9383), .A2(n5602), .B1(n5601), .B2(n9203), .ZN(n5549)
         );
  AOI22_X1 U6925 ( .A1(n9383), .A2(n5586), .B1(n5602), .B2(n9203), .ZN(n5547)
         );
  XNOR2_X1 U6926 ( .A(n5547), .B(n5599), .ZN(n5548) );
  XOR2_X1 U6927 ( .A(n5549), .B(n5548), .Z(n9030) );
  INV_X1 U6928 ( .A(n5548), .ZN(n5551) );
  INV_X1 U6929 ( .A(n5549), .ZN(n5550) );
  INV_X1 U6930 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5556) );
  INV_X1 U6931 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5555) );
  MUX2_X1 U6932 ( .A(n5556), .B(n5555), .S(n5700), .Z(n5558) );
  INV_X1 U6933 ( .A(SI_27_), .ZN(n5557) );
  NAND2_X1 U6934 ( .A1(n5558), .A2(n5557), .ZN(n6045) );
  INV_X1 U6935 ( .A(n5558), .ZN(n5559) );
  NAND2_X1 U6936 ( .A1(n5559), .A2(SI_27_), .ZN(n5560) );
  AND2_X1 U6937 ( .A1(n6045), .A2(n5560), .ZN(n5575) );
  NAND2_X1 U6938 ( .A1(n7964), .A2(n5009), .ZN(n5562) );
  NAND2_X1 U6939 ( .A1(n6340), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U6940 ( .A1(n9379), .A2(n5586), .ZN(n5571) );
  NAND2_X1 U6941 ( .A1(n6344), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U6942 ( .A1(n5084), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5568) );
  INV_X1 U6943 ( .A(n5564), .ZN(n5563) );
  NAND2_X1 U6944 ( .A1(n5563), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5589) );
  INV_X1 U6945 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8896) );
  NAND2_X1 U6946 ( .A1(n5564), .A2(n8896), .ZN(n5565) );
  NAND2_X1 U6947 ( .A1(n5413), .A2(n9194), .ZN(n5567) );
  NAND2_X1 U6948 ( .A1(n6343), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5566) );
  OR2_X1 U6949 ( .A1(n9139), .A2(n5596), .ZN(n5570) );
  NAND2_X1 U6950 ( .A1(n5571), .A2(n5570), .ZN(n5572) );
  XNOR2_X1 U6951 ( .A(n5572), .B(n4976), .ZN(n5606) );
  NOR2_X1 U6952 ( .A1(n9139), .A2(n5026), .ZN(n5573) );
  AOI21_X1 U6953 ( .B1(n9379), .B2(n5602), .A(n5573), .ZN(n5605) );
  OR2_X1 U6954 ( .A1(n5606), .A2(n5605), .ZN(n8894) );
  INV_X1 U6955 ( .A(n8894), .ZN(n5574) );
  INV_X1 U6956 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5578) );
  INV_X1 U6957 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5577) );
  MUX2_X1 U6958 ( .A(n5578), .B(n5577), .S(n5700), .Z(n5580) );
  INV_X1 U6959 ( .A(SI_28_), .ZN(n5579) );
  NAND2_X1 U6960 ( .A1(n5580), .A2(n5579), .ZN(n6044) );
  INV_X1 U6961 ( .A(n5580), .ZN(n5581) );
  NAND2_X1 U6962 ( .A1(n5581), .A2(SI_28_), .ZN(n6048) );
  AND2_X1 U6963 ( .A1(n6044), .A2(n6048), .ZN(n5582) );
  NAND2_X1 U6964 ( .A1(n8000), .A2(n5009), .ZN(n5585) );
  NAND2_X1 U6965 ( .A1(n6340), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U6966 ( .A1(n9373), .A2(n5586), .ZN(n5598) );
  NAND2_X1 U6967 ( .A1(n6343), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U6968 ( .A1(n6344), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5594) );
  INV_X1 U6969 ( .A(n5589), .ZN(n5587) );
  NAND2_X1 U6970 ( .A1(n5587), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n5640) );
  INV_X1 U6971 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U6972 ( .A1(n5589), .A2(n5588), .ZN(n5590) );
  NAND2_X1 U6973 ( .A1(n5591), .A2(n9182), .ZN(n5593) );
  NAND2_X1 U6974 ( .A1(n5084), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5592) );
  OR2_X1 U6975 ( .A1(n9197), .A2(n5596), .ZN(n5597) );
  NAND2_X1 U6976 ( .A1(n5598), .A2(n5597), .ZN(n5600) );
  XNOR2_X1 U6977 ( .A(n5600), .B(n5599), .ZN(n5604) );
  INV_X1 U6978 ( .A(n9197), .ZN(n9166) );
  AOI22_X1 U6979 ( .A1(n9373), .A2(n5602), .B1(n5601), .B2(n9166), .ZN(n5603)
         );
  XNOR2_X1 U6980 ( .A(n5604), .B(n5603), .ZN(n5634) );
  INV_X1 U6981 ( .A(n5634), .ZN(n5631) );
  NAND2_X1 U6982 ( .A1(n5606), .A2(n5605), .ZN(n8893) );
  NAND3_X1 U6983 ( .A1(n5608), .A2(P1_B_REG_SCAN_IN), .A3(n5607), .ZN(n5611)
         );
  OAI21_X1 U6984 ( .B1(n5607), .B2(P1_B_REG_SCAN_IN), .A(n7943), .ZN(n5609) );
  INV_X1 U6985 ( .A(n5609), .ZN(n5610) );
  NAND2_X1 U6986 ( .A1(n5611), .A2(n5610), .ZN(n9830) );
  OAI22_X1 U6987 ( .A1(n9830), .A2(P1_D_REG_1__SCAN_IN), .B1(n7940), .B2(n7943), .ZN(n7089) );
  NAND2_X1 U6988 ( .A1(n5612), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5613) );
  MUX2_X1 U6989 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5613), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n5615) );
  NAND2_X1 U6990 ( .A1(n5615), .A2(n5614), .ZN(n6572) );
  AND2_X1 U6991 ( .A1(n6572), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5616) );
  NAND2_X1 U6992 ( .A1(n4904), .A2(n5616), .ZN(n9837) );
  NOR2_X1 U6993 ( .A1(n7089), .A2(n9837), .ZN(n9836) );
  INV_X1 U6994 ( .A(n5607), .ZN(n7784) );
  OAI22_X1 U6995 ( .A1(n9830), .A2(P1_D_REG_0__SCAN_IN), .B1(n7943), .B2(n7784), .ZN(n6739) );
  NOR4_X1 U6996 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5625) );
  NOR4_X1 U6997 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5624) );
  OR4_X1 U6998 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5622) );
  NOR4_X1 U6999 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5620) );
  NOR4_X1 U7000 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n5619) );
  NOR4_X1 U7001 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5618) );
  NOR4_X1 U7002 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5617) );
  NAND4_X1 U7003 ( .A1(n5620), .A2(n5619), .A3(n5618), .A4(n5617), .ZN(n5621)
         );
  NOR4_X1 U7004 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5622), .A4(n5621), .ZN(n5623) );
  AND3_X1 U7005 ( .A1(n5625), .A2(n5624), .A3(n5623), .ZN(n5626) );
  NOR2_X1 U7006 ( .A1(n9830), .A2(n5626), .ZN(n6738) );
  OR2_X1 U7007 ( .A1(n6739), .A2(n6738), .ZN(n5646) );
  INV_X1 U7008 ( .A(n5646), .ZN(n5627) );
  AND2_X1 U7009 ( .A1(n9836), .A2(n5627), .ZN(n5638) );
  INV_X1 U7010 ( .A(n5638), .ZN(n5637) );
  NAND2_X1 U7011 ( .A1(n5636), .A2(n5628), .ZN(n7198) );
  INV_X1 U7012 ( .A(n7198), .ZN(n6737) );
  AND2_X2 U7013 ( .A1(n7199), .A2(n6737), .ZN(n9887) );
  AND2_X1 U7014 ( .A1(n7472), .A2(n7538), .ZN(n6895) );
  OR2_X1 U7015 ( .A1(n9887), .A2(n6895), .ZN(n5629) );
  INV_X1 U7016 ( .A(n9012), .ZN(n5630) );
  NAND2_X1 U7017 ( .A1(n5632), .A2(n4822), .ZN(n5656) );
  NAND3_X1 U7018 ( .A1(n5633), .A2(n5630), .A3(n5634), .ZN(n5655) );
  NOR3_X1 U7019 ( .A1(n5631), .A2(n9012), .A3(n8893), .ZN(n5635) );
  INV_X1 U7020 ( .A(n9373), .ZN(n9184) );
  AND2_X1 U7021 ( .A1(n9110), .A2(n5636), .ZN(n6517) );
  NAND2_X1 U7022 ( .A1(n9884), .A2(n5628), .ZN(n5649) );
  NAND2_X1 U7023 ( .A1(n5637), .A2(n9685), .ZN(n9024) );
  INV_X1 U7024 ( .A(n9038), .ZN(n7921) );
  AND2_X1 U7025 ( .A1(n6891), .A2(n7092), .ZN(n6732) );
  AND2_X1 U7026 ( .A1(n5638), .A2(n6732), .ZN(n5645) );
  NAND2_X1 U7027 ( .A1(n5645), .A2(n5639), .ZN(n9035) );
  INV_X1 U7028 ( .A(n9035), .ZN(n9022) );
  NAND2_X1 U7029 ( .A1(n6343), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U7030 ( .A1(n6344), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5643) );
  INV_X1 U7031 ( .A(n5640), .ZN(n9171) );
  NAND2_X1 U7032 ( .A1(n5413), .A2(n9171), .ZN(n5642) );
  NAND2_X1 U7033 ( .A1(n6317), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5641) );
  INV_X1 U7034 ( .A(n6518), .ZN(n9188) );
  AOI22_X1 U7035 ( .A1(n9022), .A2(n9188), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n5652) );
  INV_X1 U7036 ( .A(n5639), .ZN(n6894) );
  NAND2_X1 U7037 ( .A1(n5645), .A2(n6894), .ZN(n9032) );
  INV_X1 U7038 ( .A(n9032), .ZN(n9020) );
  INV_X1 U7039 ( .A(n9139), .ZN(n9211) );
  NAND2_X1 U7040 ( .A1(n5649), .A2(n5646), .ZN(n5648) );
  NAND2_X1 U7041 ( .A1(n7199), .A2(n6895), .ZN(n6758) );
  AND3_X1 U7042 ( .A1(n6758), .A2(n4904), .A3(n6572), .ZN(n5647) );
  NAND2_X1 U7043 ( .A1(n5648), .A2(n5647), .ZN(n6878) );
  AND2_X1 U7044 ( .A1(n5649), .A2(n7089), .ZN(n6741) );
  OR2_X1 U7045 ( .A1(n6878), .A2(n6741), .ZN(n5650) );
  AOI22_X1 U7046 ( .A1(n9020), .A2(n9211), .B1(n9182), .B2(n9033), .ZN(n5651)
         );
  OAI211_X1 U7047 ( .C1(n9184), .C2(n7921), .A(n5652), .B(n5651), .ZN(n5653)
         );
  NAND3_X1 U7048 ( .A1(n5656), .A2(n5655), .A3(n5654), .ZN(P1_U3218) );
  NOR2_X2 U7049 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5658) );
  NOR2_X1 U7050 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5664) );
  NOR2_X1 U7051 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5663) );
  NOR2_X1 U7052 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5662) );
  NOR2_X1 U7053 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5661) );
  NOR2_X1 U7054 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5666) );
  INV_X1 U7055 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6298) );
  NAND3_X1 U7056 ( .A1(n6083), .A2(n5666), .A3(n6298), .ZN(n5669) );
  INV_X1 U7057 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5938) );
  INV_X1 U7058 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5667) );
  NAND4_X1 U7059 ( .A1(n5938), .A2(n4679), .A3(n5894), .A4(n5667), .ZN(n5668)
         );
  NOR2_X1 U7060 ( .A1(n5669), .A2(n5668), .ZN(n5670) );
  INV_X1 U7061 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5671) );
  INV_X1 U7062 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5693) );
  INV_X1 U7063 ( .A(n5676), .ZN(n8885) );
  NAND2_X1 U7064 ( .A1(n5691), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5674) );
  INV_X1 U7065 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U7066 ( .A1(n6018), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5684) );
  AND2_X4 U7067 ( .A1(n5679), .A2(n8022), .ZN(n6077) );
  NAND2_X1 U7068 ( .A1(n6077), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U7069 ( .A1(n5695), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5682) );
  NAND2_X4 U7070 ( .A1(n8890), .A2(n5680), .ZN(n5754) );
  INV_X1 U7071 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7046) );
  OR2_X1 U7072 ( .A1(n5754), .A2(n7046), .ZN(n5681) );
  NAND2_X1 U7073 ( .A1(n6617), .A2(SI_0_), .ZN(n5686) );
  INV_X1 U7074 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7075 ( .A1(n5686), .A2(n5685), .ZN(n5688) );
  AND2_X1 U7076 ( .A1(n5688), .A2(n5687), .ZN(n8892) );
  OAI21_X1 U7077 ( .B1(n4309), .B2(n5818), .A(P2_IR_REG_28__SCAN_IN), .ZN(
        n5690) );
  XNOR2_X2 U7078 ( .A(n5694), .B(n5693), .ZN(n6783) );
  MUX2_X1 U7079 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8892), .S(n6769), .Z(n9938) );
  NAND2_X1 U7080 ( .A1(n6077), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U7081 ( .A1(n5695), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5698) );
  NAND2_X1 U7082 ( .A1(n4303), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5697) );
  INV_X1 U7083 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7048) );
  OR2_X1 U7084 ( .A1(n5754), .A2(n7048), .ZN(n5696) );
  NAND2_X1 U7086 ( .A1(n5880), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5703) );
  INV_X4 U7087 ( .A(n6769), .ZN(n5740) );
  NAND2_X1 U7088 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5701) );
  NAND2_X1 U7089 ( .A1(n5740), .A2(n7047), .ZN(n5702) );
  OAI211_X2 U7090 ( .C1(n5773), .C2(n6618), .A(n5703), .B(n5702), .ZN(n8050)
         );
  NAND2_X1 U7091 ( .A1(n6957), .A2(n8050), .ZN(n6151) );
  NAND2_X1 U7092 ( .A1(n7346), .A2(n6151), .ZN(n6143) );
  INV_X1 U7093 ( .A(n8050), .ZN(n9945) );
  NAND2_X1 U7094 ( .A1(n6947), .A2(n9945), .ZN(n6149) );
  NAND2_X1 U7095 ( .A1(n5695), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5707) );
  INV_X1 U7096 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7312) );
  OR2_X1 U7097 ( .A1(n5754), .A2(n7312), .ZN(n5706) );
  NAND2_X1 U7098 ( .A1(n6018), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U7099 ( .A1(n6077), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U7100 ( .A1(n5880), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5709) );
  OAI21_X1 U7101 ( .B1(P2_IR_REG_1__SCAN_IN), .B2(P2_IR_REG_0__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5714) );
  XNOR2_X1 U7102 ( .A(n5714), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6782) );
  NAND2_X1 U7103 ( .A1(n5740), .A2(n6782), .ZN(n5708) );
  INV_X1 U7104 ( .A(n7311), .ZN(n7407) );
  NAND2_X1 U7105 ( .A1(n7009), .A2(n7407), .ZN(n6144) );
  NAND2_X1 U7106 ( .A1(n6144), .A2(n7428), .ZN(n6113) );
  NAND2_X1 U7107 ( .A1(n6953), .A2(n7409), .ZN(n6954) );
  INV_X1 U7108 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6779) );
  OR2_X1 U7109 ( .A1(n5754), .A2(n6779), .ZN(n5713) );
  NAND2_X1 U7110 ( .A1(n6077), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U7111 ( .A1(n5880), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5718) );
  INV_X1 U7112 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9559) );
  NAND2_X1 U7113 ( .A1(n5714), .A2(n9559), .ZN(n5715) );
  NAND2_X1 U7114 ( .A1(n5715), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5716) );
  XNOR2_X1 U7115 ( .A(n5716), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6806) );
  NAND2_X1 U7116 ( .A1(n5740), .A2(n6806), .ZN(n5717) );
  INV_X1 U7117 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7153) );
  INV_X1 U7118 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6829) );
  NAND2_X1 U7119 ( .A1(n7153), .A2(n6829), .ZN(n5719) );
  NAND2_X1 U7120 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5751) );
  AND2_X1 U7121 ( .A1(n5719), .A2(n5751), .ZN(n8747) );
  NAND2_X1 U7122 ( .A1(n6018), .A2(n8747), .ZN(n5724) );
  NAND2_X1 U7123 ( .A1(n6077), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5723) );
  INV_X1 U7124 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5720) );
  INV_X1 U7125 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U7126 ( .A1(n5880), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5729) );
  INV_X1 U7127 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5818) );
  OR2_X1 U7128 ( .A1(n5726), .A2(n5818), .ZN(n5727) );
  XNOR2_X1 U7129 ( .A(n5727), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U7130 ( .A1(n5740), .A2(n6804), .ZN(n5728) );
  NAND2_X1 U7131 ( .A1(n6954), .A2(n5731), .ZN(n5734) );
  INV_X1 U7132 ( .A(n7445), .ZN(n7410) );
  NAND2_X1 U7133 ( .A1(n8363), .A2(n7410), .ZN(n6155) );
  NAND2_X1 U7134 ( .A1(n6155), .A2(n8736), .ZN(n6114) );
  NAND2_X1 U7135 ( .A1(n7077), .A2(n9952), .ZN(n6156) );
  NAND2_X1 U7136 ( .A1(n5734), .A2(n5733), .ZN(n7419) );
  XNOR2_X1 U7137 ( .A(n5751), .B(P2_REG3_REG_5__SCAN_IN), .ZN(n7414) );
  NAND2_X1 U7138 ( .A1(n6018), .A2(n7414), .ZN(n5739) );
  NAND2_X1 U7139 ( .A1(n6077), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5738) );
  INV_X1 U7140 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5735) );
  OR2_X1 U7141 ( .A1(n4302), .A2(n5735), .ZN(n5737) );
  INV_X1 U7142 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7422) );
  OR2_X1 U7143 ( .A1(n5754), .A2(n7422), .ZN(n5736) );
  NAND2_X1 U7144 ( .A1(n5880), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U7145 ( .A1(n5741), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5742) );
  MUX2_X1 U7146 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5742), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5744) );
  AND2_X1 U7147 ( .A1(n5744), .A2(n5743), .ZN(n6802) );
  NAND2_X1 U7148 ( .A1(n5740), .A2(n6802), .ZN(n5745) );
  OAI211_X1 U7149 ( .C1(n5773), .C2(n6625), .A(n5746), .B(n5745), .ZN(n7415)
         );
  AND2_X1 U7150 ( .A1(n8362), .A2(n9960), .ZN(n6116) );
  INV_X1 U7151 ( .A(n8362), .ZN(n7498) );
  NAND2_X1 U7152 ( .A1(n7498), .A2(n7415), .ZN(n6140) );
  INV_X1 U7153 ( .A(n5751), .ZN(n5748) );
  NAND2_X1 U7154 ( .A1(n5748), .A2(n5747), .ZN(n5765) );
  INV_X1 U7155 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5750) );
  INV_X1 U7156 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5749) );
  OAI21_X1 U7157 ( .B1(n5751), .B2(n5750), .A(n5749), .ZN(n5752) );
  AND2_X1 U7158 ( .A1(n5765), .A2(n5752), .ZN(n7375) );
  NAND2_X1 U7159 ( .A1(n6018), .A2(n7375), .ZN(n5760) );
  NAND2_X1 U7160 ( .A1(n6077), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5759) );
  INV_X1 U7161 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5753) );
  OR2_X1 U7162 ( .A1(n5754), .A2(n5753), .ZN(n5758) );
  INV_X1 U7163 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5755) );
  OR2_X1 U7164 ( .A1(n4302), .A2(n5755), .ZN(n5757) );
  NAND4_X1 U7165 ( .A1(n5760), .A2(n5759), .A3(n5758), .A4(n5757), .ZN(n8361)
         );
  NAND2_X1 U7166 ( .A1(n5880), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U7167 ( .A1(n5743), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5761) );
  XNOR2_X1 U7168 ( .A(n5761), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6800) );
  NAND2_X1 U7169 ( .A1(n5740), .A2(n6800), .ZN(n5762) );
  OAI211_X1 U7170 ( .C1(n5773), .C2(n6636), .A(n5763), .B(n5762), .ZN(n7499)
         );
  NAND2_X1 U7171 ( .A1(n7384), .A2(n7499), .ZN(n6163) );
  INV_X1 U7172 ( .A(n7499), .ZN(n9965) );
  NAND2_X1 U7173 ( .A1(n8361), .A2(n9965), .ZN(n6157) );
  NAND2_X1 U7174 ( .A1(n7544), .A2(n7546), .ZN(n7545) );
  NAND2_X1 U7175 ( .A1(n7545), .A2(n6163), .ZN(n7502) );
  INV_X1 U7176 ( .A(n5765), .ZN(n5764) );
  NAND2_X1 U7177 ( .A1(n5764), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5780) );
  INV_X1 U7178 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7383) );
  NAND2_X1 U7179 ( .A1(n5765), .A2(n7383), .ZN(n5766) );
  AND2_X1 U7180 ( .A1(n5780), .A2(n5766), .ZN(n7602) );
  NAND2_X1 U7181 ( .A1(n6018), .A2(n7602), .ZN(n5772) );
  NAND2_X1 U7182 ( .A1(n6077), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5771) );
  INV_X1 U7183 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5767) );
  INV_X1 U7184 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5768) );
  OR2_X1 U7185 ( .A1(n4302), .A2(n5768), .ZN(n5769) );
  NAND2_X1 U7186 ( .A1(n6642), .A2(n6071), .ZN(n5778) );
  OR2_X1 U7187 ( .A1(n5774), .A2(n5818), .ZN(n5775) );
  XNOR2_X1 U7188 ( .A(n5775), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6845) );
  NAND2_X1 U7189 ( .A1(n5740), .A2(n6845), .ZN(n5777) );
  NAND2_X1 U7190 ( .A1(n5880), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n5776) );
  NAND2_X1 U7191 ( .A1(n8360), .A2(n7604), .ZN(n6169) );
  INV_X1 U7192 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U7193 ( .A1(n5780), .A2(n5779), .ZN(n5781) );
  AND2_X1 U7194 ( .A1(n5798), .A2(n5781), .ZN(n8242) );
  NAND2_X1 U7195 ( .A1(n6018), .A2(n8242), .ZN(n5787) );
  NAND2_X1 U7196 ( .A1(n6077), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5786) );
  INV_X1 U7197 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5782) );
  INV_X1 U7198 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U7199 ( .A1(n6646), .A2(n6071), .ZN(n5791) );
  OR2_X1 U7200 ( .A1(n5788), .A2(n5818), .ZN(n5789) );
  XNOR2_X1 U7201 ( .A(n5789), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6906) );
  AOI22_X1 U7202 ( .A1(n5880), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5740), .B2(
        n6906), .ZN(n5790) );
  INV_X1 U7203 ( .A(n8239), .ZN(n9969) );
  NAND2_X1 U7204 ( .A1(n9969), .A2(n8359), .ZN(n6174) );
  NAND2_X1 U7205 ( .A1(n6660), .A2(n6071), .ZN(n5797) );
  INV_X1 U7206 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U7207 ( .A1(n5788), .A2(n5792), .ZN(n5794) );
  NAND2_X1 U7208 ( .A1(n5794), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5793) );
  MUX2_X1 U7209 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5793), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n5795) );
  AND2_X1 U7210 ( .A1(n5795), .A2(n5817), .ZN(n7178) );
  AOI22_X1 U7211 ( .A1(n5880), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5740), .B2(
        n7178), .ZN(n5796) );
  AND2_X2 U7212 ( .A1(n5797), .A2(n5796), .ZN(n7764) );
  NAND2_X1 U7213 ( .A1(n6077), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5806) );
  NAND2_X1 U7214 ( .A1(n5798), .A2(n9586), .ZN(n5799) );
  NAND2_X1 U7215 ( .A1(n5826), .A2(n5799), .ZN(n7597) );
  INV_X1 U7216 ( .A(n7597), .ZN(n5800) );
  NAND2_X1 U7217 ( .A1(n6018), .A2(n5800), .ZN(n5805) );
  INV_X1 U7218 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5801) );
  OR2_X1 U7219 ( .A1(n4302), .A2(n5801), .ZN(n5804) );
  INV_X1 U7220 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5802) );
  OR2_X1 U7221 ( .A1(n5754), .A2(n5802), .ZN(n5803) );
  NAND4_X1 U7222 ( .A1(n5806), .A2(n5805), .A3(n5804), .A4(n5803), .ZN(n8358)
         );
  NAND2_X1 U7223 ( .A1(n7764), .A2(n8358), .ZN(n6185) );
  INV_X1 U7224 ( .A(n7764), .ZN(n7655) );
  INV_X1 U7225 ( .A(n8358), .ZN(n7665) );
  NAND2_X1 U7226 ( .A1(n6664), .A2(n6071), .ZN(n5809) );
  NAND2_X1 U7227 ( .A1(n5817), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5807) );
  XNOR2_X1 U7228 ( .A(n5807), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7397) );
  AOI22_X1 U7229 ( .A1(n6096), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5740), .B2(
        n7397), .ZN(n5808) );
  NAND2_X1 U7230 ( .A1(n6077), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5815) );
  XNOR2_X1 U7231 ( .A(n5826), .B(P2_REG3_REG_10__SCAN_IN), .ZN(n8220) );
  NAND2_X1 U7232 ( .A1(n6018), .A2(n8220), .ZN(n5814) );
  INV_X1 U7233 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5810) );
  OR2_X1 U7234 ( .A1(n4302), .A2(n5810), .ZN(n5813) );
  INV_X1 U7235 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5811) );
  OR2_X1 U7236 ( .A1(n5754), .A2(n5811), .ZN(n5812) );
  NAND4_X1 U7237 ( .A1(n5815), .A2(n5814), .A3(n5813), .A4(n5812), .ZN(n8357)
         );
  AND2_X1 U7238 ( .A1(n9974), .A2(n8357), .ZN(n6180) );
  INV_X1 U7239 ( .A(n9974), .ZN(n8218) );
  INV_X1 U7240 ( .A(n8357), .ZN(n5816) );
  NAND2_X1 U7241 ( .A1(n8218), .A2(n5816), .ZN(n6186) );
  NAND2_X1 U7242 ( .A1(n6666), .A2(n6071), .ZN(n5821) );
  NOR2_X1 U7243 ( .A1(n5817), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5834) );
  OR2_X1 U7244 ( .A1(n5834), .A2(n5818), .ZN(n5819) );
  XNOR2_X1 U7245 ( .A(n5819), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7562) );
  AOI22_X1 U7246 ( .A1(n6096), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5740), .B2(
        n7562), .ZN(n5820) );
  INV_X1 U7247 ( .A(n5826), .ZN(n5823) );
  AND2_X1 U7248 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n5822) );
  NAND2_X1 U7249 ( .A1(n5823), .A2(n5822), .ZN(n5839) );
  INV_X1 U7250 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5825) );
  INV_X1 U7251 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5824) );
  OAI21_X1 U7252 ( .B1(n5826), .B2(n5825), .A(n5824), .ZN(n5827) );
  AND2_X1 U7253 ( .A1(n5839), .A2(n5827), .ZN(n7795) );
  NAND2_X1 U7254 ( .A1(n6018), .A2(n7795), .ZN(n5832) );
  NAND2_X1 U7255 ( .A1(n6077), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5831) );
  INV_X1 U7256 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5828) );
  OR2_X1 U7257 ( .A1(n4302), .A2(n5828), .ZN(n5830) );
  INV_X1 U7258 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7391) );
  OR2_X1 U7259 ( .A1(n5754), .A2(n7391), .ZN(n5829) );
  NAND4_X1 U7260 ( .A1(n5832), .A2(n5831), .A3(n5830), .A4(n5829), .ZN(n8356)
         );
  INV_X1 U7261 ( .A(n8356), .ZN(n7897) );
  NOR2_X1 U7262 ( .A1(n7798), .A2(n6193), .ZN(n7893) );
  NAND2_X1 U7263 ( .A1(n6698), .A2(n6071), .ZN(n5837) );
  INV_X1 U7264 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U7265 ( .A1(n5834), .A2(n5833), .ZN(n5847) );
  NAND2_X1 U7266 ( .A1(n5847), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5835) );
  XNOR2_X1 U7267 ( .A(n5835), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8369) );
  AOI22_X1 U7268 ( .A1(n6096), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5740), .B2(
        n8369), .ZN(n5836) );
  NAND2_X1 U7269 ( .A1(n6077), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5846) );
  INV_X1 U7270 ( .A(n5839), .ZN(n5838) );
  NAND2_X1 U7271 ( .A1(n5838), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5851) );
  INV_X1 U7272 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9503) );
  NAND2_X1 U7273 ( .A1(n5839), .A2(n9503), .ZN(n5840) );
  AND2_X1 U7274 ( .A1(n5851), .A2(n5840), .ZN(n7901) );
  NAND2_X1 U7275 ( .A1(n6018), .A2(n7901), .ZN(n5845) );
  INV_X1 U7276 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5841) );
  OR2_X1 U7277 ( .A1(n4302), .A2(n5841), .ZN(n5844) );
  INV_X1 U7278 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5842) );
  OR2_X1 U7279 ( .A1(n5754), .A2(n5842), .ZN(n5843) );
  NAND4_X1 U7280 ( .A1(n5846), .A2(n5845), .A3(n5844), .A4(n5843), .ZN(n8355)
         );
  INV_X1 U7281 ( .A(n8355), .ZN(n8105) );
  OR2_X1 U7282 ( .A1(n7902), .A2(n8105), .ZN(n6198) );
  NAND2_X1 U7283 ( .A1(n6198), .A2(n7891), .ZN(n6195) );
  NOR2_X1 U7284 ( .A1(n7893), .A2(n6195), .ZN(n7877) );
  NAND2_X1 U7285 ( .A1(n6744), .A2(n6071), .ZN(n5850) );
  OR2_X1 U7286 ( .A1(n5847), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5848) );
  NAND2_X1 U7287 ( .A1(n5848), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5860) );
  XNOR2_X1 U7288 ( .A(n5860), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7734) );
  AOI22_X1 U7289 ( .A1(n6096), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5740), .B2(
        n7734), .ZN(n5849) );
  INV_X1 U7290 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7567) );
  NAND2_X1 U7291 ( .A1(n5851), .A2(n7567), .ZN(n5852) );
  AND2_X1 U7292 ( .A1(n5869), .A2(n5852), .ZN(n8103) );
  NAND2_X1 U7293 ( .A1(n6018), .A2(n8103), .ZN(n5858) );
  NAND2_X1 U7294 ( .A1(n6077), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5857) );
  INV_X1 U7295 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n5853) );
  OR2_X1 U7296 ( .A1(n4302), .A2(n5853), .ZN(n5856) );
  INV_X1 U7297 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5854) );
  OR2_X1 U7298 ( .A1(n5754), .A2(n5854), .ZN(n5855) );
  NAND4_X1 U7299 ( .A1(n5858), .A2(n5857), .A3(n5856), .A4(n5855), .ZN(n8354)
         );
  OR2_X1 U7300 ( .A1(n8108), .A2(n7994), .ZN(n6202) );
  NAND2_X1 U7301 ( .A1(n8108), .A2(n7994), .ZN(n6201) );
  OAI21_X1 U7302 ( .B1(n7877), .B2(n7875), .A(n7876), .ZN(n7879) );
  NAND2_X1 U7303 ( .A1(n6746), .A2(n6071), .ZN(n5866) );
  INV_X1 U7304 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U7305 ( .A1(n5860), .A2(n5859), .ZN(n5861) );
  NAND2_X1 U7306 ( .A1(n5861), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5863) );
  INV_X1 U7307 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U7308 ( .A1(n5863), .A2(n5862), .ZN(n5878) );
  OR2_X1 U7309 ( .A1(n5863), .A2(n5862), .ZN(n5864) );
  AOI22_X1 U7310 ( .A1(n6096), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5740), .B2(
        n7955), .ZN(n5865) );
  INV_X1 U7311 ( .A(n5869), .ZN(n5867) );
  NAND2_X1 U7312 ( .A1(n5867), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5884) );
  INV_X1 U7313 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7314 ( .A1(n5869), .A2(n5868), .ZN(n5870) );
  AND2_X1 U7315 ( .A1(n5884), .A2(n5870), .ZN(n8095) );
  NAND2_X1 U7316 ( .A1(n6018), .A2(n8095), .ZN(n5876) );
  NAND2_X1 U7317 ( .A1(n6077), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5875) );
  INV_X1 U7318 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n5871) );
  OR2_X1 U7319 ( .A1(n4302), .A2(n5871), .ZN(n5874) );
  INV_X1 U7320 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5872) );
  OR2_X1 U7321 ( .A1(n5754), .A2(n5872), .ZN(n5873) );
  NAND4_X1 U7322 ( .A1(n5876), .A2(n5875), .A3(n5874), .A4(n5873), .ZN(n8458)
         );
  NAND2_X1 U7323 ( .A1(n8842), .A2(n8727), .ZN(n6204) );
  NAND2_X1 U7324 ( .A1(n5877), .A2(n6204), .ZN(n7993) );
  INV_X1 U7325 ( .A(n5877), .ZN(n6213) );
  NAND2_X1 U7326 ( .A1(n6876), .A2(n6071), .ZN(n5882) );
  NAND2_X1 U7327 ( .A1(n5878), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5879) );
  XNOR2_X1 U7328 ( .A(n5879), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8390) );
  AOI22_X1 U7329 ( .A1(n8390), .A2(n5740), .B1(n5880), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U7330 ( .A1(n6077), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5891) );
  INV_X1 U7331 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5883) );
  NAND2_X1 U7332 ( .A1(n5884), .A2(n5883), .ZN(n5885) );
  AND2_X1 U7333 ( .A1(n5901), .A2(n5885), .ZN(n8719) );
  NAND2_X1 U7334 ( .A1(n6018), .A2(n8719), .ZN(n5890) );
  INV_X1 U7335 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n5886) );
  OR2_X1 U7336 ( .A1(n4302), .A2(n5886), .ZN(n5889) );
  INV_X1 U7337 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n5887) );
  OR2_X1 U7338 ( .A1(n5754), .A2(n5887), .ZN(n5888) );
  NAND4_X1 U7339 ( .A1(n5891), .A2(n5890), .A3(n5889), .A4(n5888), .ZN(n8461)
         );
  NAND2_X1 U7340 ( .A1(n8837), .A2(n8273), .ZN(n6214) );
  NAND2_X1 U7341 ( .A1(n6926), .A2(n6071), .ZN(n5898) );
  NOR2_X1 U7342 ( .A1(n5895), .A2(n5818), .ZN(n5892) );
  MUX2_X1 U7343 ( .A(n5818), .B(n5892), .S(P2_IR_REG_16__SCAN_IN), .Z(n5893)
         );
  INV_X1 U7344 ( .A(n5893), .ZN(n5896) );
  AND2_X1 U7345 ( .A1(n5896), .A2(n5911), .ZN(n8407) );
  AOI22_X1 U7346 ( .A1(n6096), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5740), .B2(
        n8407), .ZN(n5897) );
  INV_X1 U7347 ( .A(n5901), .ZN(n5899) );
  NAND2_X1 U7348 ( .A1(n5899), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5916) );
  INV_X1 U7349 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U7350 ( .A1(n5901), .A2(n5900), .ZN(n5902) );
  AND2_X1 U7351 ( .A1(n5916), .A2(n5902), .ZN(n8702) );
  NAND2_X1 U7352 ( .A1(n6018), .A2(n8702), .ZN(n5908) );
  NAND2_X1 U7353 ( .A1(n6077), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5907) );
  INV_X1 U7354 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n5903) );
  OR2_X1 U7355 ( .A1(n4302), .A2(n5903), .ZN(n5906) );
  INV_X1 U7356 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5904) );
  OR2_X1 U7357 ( .A1(n5754), .A2(n5904), .ZN(n5905) );
  NAND4_X1 U7358 ( .A1(n5908), .A2(n5907), .A3(n5906), .A4(n5905), .ZN(n8463)
         );
  INV_X1 U7359 ( .A(n8463), .ZN(n8729) );
  OR2_X1 U7360 ( .A1(n8832), .A2(n8729), .ZN(n6208) );
  NAND2_X1 U7361 ( .A1(n8832), .A2(n8729), .ZN(n6207) );
  NAND2_X1 U7362 ( .A1(n8707), .A2(n8705), .ZN(n5909) );
  NAND2_X1 U7363 ( .A1(n7103), .A2(n6071), .ZN(n5914) );
  NAND2_X1 U7364 ( .A1(n5911), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5910) );
  MUX2_X1 U7365 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5910), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5912) );
  AND2_X1 U7366 ( .A1(n5912), .A2(n4362), .ZN(n8419) );
  AOI22_X1 U7367 ( .A1(n6096), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5740), .B2(
        n8419), .ZN(n5913) );
  INV_X1 U7368 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U7369 ( .A1(n5916), .A2(n5915), .ZN(n5917) );
  AND2_X1 U7370 ( .A1(n5929), .A2(n5917), .ZN(n8685) );
  NAND2_X1 U7371 ( .A1(n6018), .A2(n8685), .ZN(n5923) );
  NAND2_X1 U7372 ( .A1(n6077), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5922) );
  INV_X1 U7373 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n5918) );
  OR2_X1 U7374 ( .A1(n5754), .A2(n5918), .ZN(n5921) );
  INV_X1 U7375 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n5919) );
  OR2_X1 U7376 ( .A1(n4302), .A2(n5919), .ZN(n5920) );
  NAND4_X1 U7377 ( .A1(n5923), .A2(n5922), .A3(n5921), .A4(n5920), .ZN(n8465)
         );
  INV_X1 U7378 ( .A(n8465), .ZN(n8272) );
  NAND2_X1 U7379 ( .A1(n8828), .A2(n8272), .ZN(n6218) );
  NAND2_X1 U7380 ( .A1(n7206), .A2(n6071), .ZN(n5926) );
  NAND2_X1 U7381 ( .A1(n4362), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5924) );
  XNOR2_X1 U7382 ( .A(n5924), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8432) );
  AOI22_X1 U7383 ( .A1(n6096), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5740), .B2(
        n8432), .ZN(n5925) );
  INV_X1 U7384 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7385 ( .A1(n5929), .A2(n5928), .ZN(n5930) );
  AND2_X1 U7386 ( .A1(n5953), .A2(n5930), .ZN(n8675) );
  NAND2_X1 U7387 ( .A1(n6018), .A2(n8675), .ZN(n5935) );
  NAND2_X1 U7388 ( .A1(n6077), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5934) );
  INV_X1 U7389 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8666) );
  OR2_X1 U7390 ( .A1(n5754), .A2(n8666), .ZN(n5933) );
  INV_X1 U7391 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n5931) );
  OR2_X1 U7392 ( .A1(n4302), .A2(n5931), .ZN(n5932) );
  NAND4_X1 U7393 ( .A1(n5935), .A2(n5934), .A3(n5933), .A4(n5932), .ZN(n8468)
         );
  INV_X1 U7394 ( .A(n8468), .ZN(n8469) );
  NOR2_X1 U7395 ( .A1(n8824), .A2(n8469), .ZN(n6231) );
  AND2_X1 U7396 ( .A1(n8824), .A2(n8469), .ZN(n5936) );
  NOR2_X1 U7397 ( .A1(n6231), .A2(n5936), .ZN(n8672) );
  NAND2_X1 U7398 ( .A1(n8672), .A2(n8669), .ZN(n5937) );
  INV_X1 U7399 ( .A(n5936), .ZN(n6228) );
  NAND2_X1 U7400 ( .A1(n7290), .A2(n6071), .ZN(n5943) );
  NAND2_X1 U7401 ( .A1(n6082), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U7402 ( .A1(n5940), .A2(n5939), .ZN(n6105) );
  OR2_X1 U7403 ( .A1(n5940), .A2(n5939), .ZN(n5941) );
  AOI22_X1 U7404 ( .A1(n6096), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5740), .B2(
        n8554), .ZN(n5942) );
  XNOR2_X1 U7405 ( .A(n5953), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U7406 ( .A1(n4303), .A2(n8653), .ZN(n5949) );
  NAND2_X1 U7407 ( .A1(n6077), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5948) );
  INV_X1 U7408 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5944) );
  OR2_X1 U7409 ( .A1(n5754), .A2(n5944), .ZN(n5947) );
  INV_X1 U7410 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n5945) );
  OR2_X1 U7411 ( .A1(n4302), .A2(n5945), .ZN(n5946) );
  NAND4_X1 U7412 ( .A1(n5949), .A2(n5948), .A3(n5947), .A4(n5946), .ZN(n8471)
         );
  INV_X1 U7413 ( .A(n8471), .ZN(n8644) );
  OR2_X1 U7414 ( .A1(n8818), .A2(n8644), .ZN(n6232) );
  NAND2_X1 U7415 ( .A1(n8818), .A2(n8644), .ZN(n6237) );
  NAND2_X1 U7416 ( .A1(n7452), .A2(n6071), .ZN(n5951) );
  NAND2_X1 U7417 ( .A1(n5880), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5950) );
  INV_X1 U7418 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8231) );
  INV_X1 U7419 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8303) );
  OAI21_X1 U7420 ( .B1(n5953), .B2(n8231), .A(n8303), .ZN(n5954) );
  NAND2_X1 U7421 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .ZN(n5952) );
  AND2_X1 U7422 ( .A1(n5954), .A2(n5965), .ZN(n8639) );
  NAND2_X1 U7423 ( .A1(n4303), .A2(n8639), .ZN(n5960) );
  NAND2_X1 U7424 ( .A1(n6077), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5959) );
  INV_X1 U7425 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5955) );
  OR2_X1 U7426 ( .A1(n5754), .A2(n5955), .ZN(n5958) );
  INV_X1 U7427 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n5956) );
  OR2_X1 U7428 ( .A1(n4302), .A2(n5956), .ZN(n5957) );
  NAND4_X1 U7429 ( .A1(n5960), .A2(n5959), .A3(n5958), .A4(n5957), .ZN(n8631)
         );
  INV_X1 U7430 ( .A(n8631), .ZN(n8250) );
  NAND2_X1 U7431 ( .A1(n8812), .A2(n8250), .ZN(n6246) );
  INV_X1 U7432 ( .A(n6241), .ZN(n6236) );
  NAND2_X1 U7433 ( .A1(n7471), .A2(n6071), .ZN(n5962) );
  NAND2_X1 U7434 ( .A1(n5880), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5961) );
  INV_X1 U7435 ( .A(n5965), .ZN(n5964) );
  NAND2_X1 U7436 ( .A1(n5964), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5977) );
  INV_X1 U7437 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8249) );
  NAND2_X1 U7438 ( .A1(n5965), .A2(n8249), .ZN(n5966) );
  NAND2_X1 U7439 ( .A1(n5977), .A2(n5966), .ZN(n8624) );
  OR2_X1 U7440 ( .A1(n5963), .A2(n8624), .ZN(n5971) );
  NAND2_X1 U7441 ( .A1(n5695), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U7442 ( .A1(n6077), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5969) );
  INV_X1 U7443 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n5967) );
  OR2_X1 U7444 ( .A1(n5754), .A2(n5967), .ZN(n5968) );
  NAND4_X1 U7445 ( .A1(n5971), .A2(n5970), .A3(n5969), .A4(n5968), .ZN(n8616)
         );
  XNOR2_X1 U7446 ( .A(n8807), .B(n8616), .ZN(n8628) );
  INV_X1 U7447 ( .A(n8616), .ZN(n8645) );
  AND2_X1 U7448 ( .A1(n8807), .A2(n8645), .ZN(n6248) );
  NAND2_X1 U7449 ( .A1(n7537), .A2(n6071), .ZN(n5973) );
  NAND2_X1 U7450 ( .A1(n5880), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5972) );
  INV_X1 U7451 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9491) );
  OR2_X1 U7452 ( .A1(n4302), .A2(n9491), .ZN(n5976) );
  INV_X1 U7453 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5974) );
  OR2_X1 U7454 ( .A1(n5754), .A2(n5974), .ZN(n5975) );
  AND2_X1 U7455 ( .A1(n5976), .A2(n5975), .ZN(n5981) );
  INV_X1 U7456 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8313) );
  NAND2_X1 U7457 ( .A1(n5977), .A2(n8313), .ZN(n5978) );
  NAND2_X1 U7458 ( .A1(n5985), .A2(n5978), .ZN(n8609) );
  OR2_X1 U7459 ( .A1(n8609), .A2(n5963), .ZN(n5980) );
  NAND2_X1 U7460 ( .A1(n6077), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U7461 ( .A1(n8802), .A2(n8475), .ZN(n6253) );
  NAND2_X1 U7462 ( .A1(n7701), .A2(n6071), .ZN(n5983) );
  NAND2_X1 U7463 ( .A1(n5880), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5982) );
  INV_X1 U7464 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7465 ( .A1(n5985), .A2(n5984), .ZN(n5986) );
  NAND2_X1 U7466 ( .A1(n5993), .A2(n5986), .ZN(n8590) );
  INV_X1 U7467 ( .A(n5754), .ZN(n6074) );
  AOI22_X1 U7468 ( .A1(n6074), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n5695), .B2(
        P2_REG0_REG_23__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U7469 ( .A1(n6077), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5987) );
  OAI211_X1 U7470 ( .C1(n8590), .C2(n5963), .A(n5988), .B(n5987), .ZN(n8617)
         );
  INV_X1 U7471 ( .A(n8617), .ZN(n8479) );
  OR2_X1 U7472 ( .A1(n8797), .A2(n8479), .ZN(n6258) );
  NAND2_X1 U7473 ( .A1(n8797), .A2(n8479), .ZN(n6261) );
  NAND2_X1 U7474 ( .A1(n7783), .A2(n6071), .ZN(n5991) );
  NAND2_X1 U7475 ( .A1(n5880), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5990) );
  INV_X1 U7476 ( .A(n5993), .ZN(n5992) );
  NAND2_X1 U7477 ( .A1(n5992), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6001) );
  INV_X1 U7478 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8294) );
  NAND2_X1 U7479 ( .A1(n5993), .A2(n8294), .ZN(n5994) );
  AND2_X1 U7480 ( .A1(n6001), .A2(n5994), .ZN(n8576) );
  NAND2_X1 U7481 ( .A1(n8576), .A2(n6018), .ZN(n5997) );
  AOI22_X1 U7482 ( .A1(n6074), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n5695), .B2(
        P2_REG0_REG_24__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7483 ( .A1(n6077), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7484 ( .A1(n8792), .A2(n8480), .ZN(n6263) );
  NAND2_X1 U7485 ( .A1(n5880), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5998) );
  INV_X1 U7486 ( .A(n6001), .ZN(n6000) );
  NAND2_X1 U7487 ( .A1(n6000), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6012) );
  INV_X1 U7488 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9526) );
  NAND2_X1 U7489 ( .A1(n6001), .A2(n9526), .ZN(n6002) );
  NAND2_X1 U7490 ( .A1(n6012), .A2(n6002), .ZN(n8561) );
  OR2_X1 U7491 ( .A1(n8561), .A2(n5963), .ZN(n6008) );
  INV_X1 U7492 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6005) );
  INV_X1 U7493 ( .A(n6077), .ZN(n6060) );
  NAND2_X1 U7494 ( .A1(n6074), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U7495 ( .A1(n5695), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6003) );
  OAI211_X1 U7496 ( .C1(n6005), .C2(n6060), .A(n6004), .B(n6003), .ZN(n6006)
         );
  INV_X1 U7497 ( .A(n6006), .ZN(n6007) );
  NAND2_X1 U7498 ( .A1(n6008), .A2(n6007), .ZN(n8580) );
  NAND2_X1 U7499 ( .A1(n6009), .A2(n8567), .ZN(n8541) );
  NAND2_X1 U7500 ( .A1(n5880), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6010) );
  INV_X1 U7501 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8330) );
  NAND2_X1 U7502 ( .A1(n6012), .A2(n8330), .ZN(n6013) );
  INV_X1 U7503 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7504 ( .A1(n6074), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7505 ( .A1(n5695), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6014) );
  OAI211_X1 U7506 ( .C1(n6016), .C2(n6060), .A(n6015), .B(n6014), .ZN(n6017)
         );
  AOI21_X1 U7507 ( .B1(n8551), .B2(n4303), .A(n6017), .ZN(n8352) );
  INV_X1 U7508 ( .A(n8580), .ZN(n8295) );
  NOR2_X1 U7509 ( .A1(n8788), .A2(n8295), .ZN(n6269) );
  NOR2_X1 U7510 ( .A1(n8546), .A2(n6269), .ZN(n6019) );
  NAND2_X1 U7511 ( .A1(n5880), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6020) );
  INV_X1 U7512 ( .A(n6024), .ZN(n6022) );
  NAND2_X1 U7513 ( .A1(n6022), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6036) );
  INV_X1 U7514 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7515 ( .A1(n6024), .A2(n6023), .ZN(n6025) );
  NAND2_X1 U7516 ( .A1(n6036), .A2(n6025), .ZN(n8532) );
  OR2_X1 U7517 ( .A1(n8532), .A2(n5963), .ZN(n6031) );
  INV_X1 U7518 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U7519 ( .A1(n6077), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U7520 ( .A1(n6074), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6026) );
  OAI211_X1 U7521 ( .C1(n4302), .C2(n6028), .A(n6027), .B(n6026), .ZN(n6029)
         );
  INV_X1 U7522 ( .A(n6029), .ZN(n6030) );
  NAND2_X1 U7523 ( .A1(n8000), .A2(n6071), .ZN(n6033) );
  NAND2_X1 U7524 ( .A1(n5880), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6032) );
  INV_X1 U7525 ( .A(n6036), .ZN(n6034) );
  NAND2_X1 U7526 ( .A1(n6034), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8499) );
  INV_X1 U7527 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7528 ( .A1(n6036), .A2(n6035), .ZN(n6037) );
  NAND2_X1 U7529 ( .A1(n8499), .A2(n6037), .ZN(n8188) );
  OR2_X1 U7530 ( .A1(n8188), .A2(n5963), .ZN(n6043) );
  INV_X1 U7531 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7532 ( .A1(n6074), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7533 ( .A1(n5695), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6038) );
  OAI211_X1 U7534 ( .C1(n6040), .C2(n6060), .A(n6039), .B(n6038), .ZN(n6041)
         );
  INV_X1 U7535 ( .A(n6041), .ZN(n6042) );
  NAND2_X1 U7536 ( .A1(n8770), .A2(n8488), .ZN(n6275) );
  NAND2_X1 U7537 ( .A1(n8513), .A2(n8507), .ZN(n8512) );
  NAND2_X1 U7538 ( .A1(n8512), .A2(n6278), .ZN(n8491) );
  AND2_X1 U7539 ( .A1(n6045), .A2(n6044), .ZN(n6046) );
  NAND2_X1 U7540 ( .A1(n6047), .A2(n6046), .ZN(n6049) );
  INV_X1 U7541 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n6051) );
  INV_X1 U7542 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n6050) );
  MUX2_X1 U7543 ( .A(n6051), .B(n6050), .S(n5327), .Z(n6053) );
  INV_X1 U7544 ( .A(SI_29_), .ZN(n6052) );
  NAND2_X1 U7545 ( .A1(n6053), .A2(n6052), .ZN(n6068) );
  INV_X1 U7546 ( .A(n6053), .ZN(n6054) );
  NAND2_X1 U7547 ( .A1(n6054), .A2(SI_29_), .ZN(n6055) );
  AND2_X1 U7548 ( .A1(n6068), .A2(n6055), .ZN(n6066) );
  NAND2_X1 U7549 ( .A1(n8021), .A2(n6071), .ZN(n6057) );
  NAND2_X1 U7550 ( .A1(n6096), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6056) );
  OR2_X1 U7551 ( .A1(n8499), .A2(n5963), .ZN(n6064) );
  INV_X1 U7552 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7553 ( .A1(n5695), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7554 ( .A1(n6074), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6058) );
  OAI211_X1 U7555 ( .C1(n6061), .C2(n6060), .A(n6059), .B(n6058), .ZN(n6062)
         );
  INV_X1 U7556 ( .A(n6062), .ZN(n6063) );
  INV_X1 U7557 ( .A(n6282), .ZN(n6065) );
  NAND2_X1 U7558 ( .A1(n8766), .A2(n8517), .ZN(n6283) );
  INV_X1 U7559 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n6070) );
  INV_X1 U7560 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n6069) );
  MUX2_X1 U7561 ( .A(n6070), .B(n6069), .S(n6617), .Z(n6089) );
  NAND2_X1 U7562 ( .A1(n8888), .A2(n6071), .ZN(n6073) );
  NAND2_X1 U7563 ( .A1(n6096), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6072) );
  INV_X1 U7564 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9591) );
  NAND2_X1 U7565 ( .A1(n6074), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7566 ( .A1(n6077), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6075) );
  OAI211_X1 U7567 ( .C1(n4302), .C2(n9591), .A(n6076), .B(n6075), .ZN(n8493)
         );
  INV_X1 U7568 ( .A(n8493), .ZN(n6099) );
  OR2_X1 U7569 ( .A1(n8454), .A2(n6099), .ZN(n6286) );
  INV_X1 U7570 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7571 ( .A1(n6077), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6080) );
  INV_X1 U7572 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6078) );
  OR2_X1 U7573 ( .A1(n4302), .A2(n6078), .ZN(n6079) );
  OAI211_X1 U7574 ( .C1(n5754), .C2(n6081), .A(n6080), .B(n6079), .ZN(n8450)
         );
  NAND2_X1 U7575 ( .A1(n6084), .A2(n6083), .ZN(n6103) );
  NAND2_X1 U7576 ( .A1(n6103), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6085) );
  OR2_X1 U7577 ( .A1(n8450), .A2(n7493), .ZN(n6086) );
  INV_X1 U7578 ( .A(n6087), .ZN(n6088) );
  NAND2_X1 U7579 ( .A1(n6088), .A2(SI_30_), .ZN(n6092) );
  NAND2_X1 U7580 ( .A1(n6092), .A2(n6091), .ZN(n6095) );
  MUX2_X1 U7581 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n6617), .Z(n6093) );
  XNOR2_X1 U7582 ( .A(n6093), .B(SI_31_), .ZN(n6094) );
  NAND2_X1 U7583 ( .A1(n8884), .A2(n6071), .ZN(n6098) );
  NAND2_X1 U7584 ( .A1(n6096), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7585 ( .A1(n8454), .A2(n6099), .ZN(n6285) );
  AOI21_X1 U7586 ( .B1(n6101), .B2(n6137), .A(n6290), .ZN(n6102) );
  XNOR2_X1 U7587 ( .A(n6102), .B(n8440), .ZN(n6110) );
  NAND2_X1 U7588 ( .A1(n6105), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6107) );
  XNOR2_X1 U7589 ( .A(n6107), .B(n6106), .ZN(n7455) );
  NAND2_X1 U7590 ( .A1(n7455), .A2(n8440), .ZN(n6997) );
  OR2_X1 U7591 ( .A1(n7303), .A2(n6997), .ZN(n6108) );
  INV_X1 U7592 ( .A(n7455), .ZN(n6961) );
  NAND2_X1 U7593 ( .A1(n6961), .A2(n7007), .ZN(n6955) );
  NAND2_X1 U7594 ( .A1(n6108), .A2(n6955), .ZN(n6109) );
  INV_X1 U7595 ( .A(n6137), .ZN(n6132) );
  INV_X1 U7596 ( .A(n6290), .ZN(n6111) );
  NAND2_X1 U7597 ( .A1(n6111), .A2(n6286), .ZN(n6135) );
  INV_X1 U7598 ( .A(n8690), .ZN(n6210) );
  INV_X1 U7599 ( .A(n7876), .ZN(n6199) );
  INV_X1 U7600 ( .A(n7875), .ZN(n6197) );
  INV_X1 U7601 ( .A(n6113), .ZN(n7409) );
  INV_X1 U7602 ( .A(n6114), .ZN(n7430) );
  INV_X1 U7603 ( .A(n9938), .ZN(n6115) );
  NAND2_X1 U7604 ( .A1(n6945), .A2(n6115), .ZN(n7033) );
  AND2_X1 U7605 ( .A1(n7346), .A2(n7033), .ZN(n7307) );
  AND4_X1 U7606 ( .A1(n7409), .A2(n6961), .A3(n7430), .A4(n7307), .ZN(n6120)
         );
  INV_X1 U7607 ( .A(n6116), .ZN(n6158) );
  NAND2_X1 U7608 ( .A1(n6140), .A2(n6158), .ZN(n7496) );
  INV_X1 U7609 ( .A(n7496), .ZN(n6119) );
  NAND2_X1 U7610 ( .A1(n6117), .A2(n6156), .ZN(n8750) );
  NOR2_X1 U7611 ( .A1(n6946), .A2(n8750), .ZN(n6118) );
  NAND4_X1 U7612 ( .A1(n6120), .A2(n6119), .A3(n7546), .A4(n6118), .ZN(n6122)
         );
  NAND2_X1 U7613 ( .A1(n6185), .A2(n6177), .ZN(n7514) );
  INV_X1 U7614 ( .A(n6121), .ZN(n6168) );
  AND2_X2 U7615 ( .A1(n6168), .A2(n6169), .ZN(n7707) );
  NOR4_X1 U7616 ( .A1(n6122), .A2(n7514), .A3(n6165), .A4(n7714), .ZN(n6124)
         );
  INV_X1 U7617 ( .A(n6193), .ZN(n6123) );
  NAND2_X1 U7618 ( .A1(n7891), .A2(n6123), .ZN(n7865) );
  INV_X1 U7619 ( .A(n7865), .ZN(n7799) );
  INV_X1 U7620 ( .A(n6180), .ZN(n6183) );
  NAND4_X1 U7621 ( .A1(n7895), .A2(n6124), .A3(n7799), .A4(n7664), .ZN(n6125)
         );
  NOR4_X1 U7622 ( .A1(n8725), .A2(n7993), .A3(n6199), .A4(n6125), .ZN(n6126)
         );
  NAND4_X1 U7623 ( .A1(n8672), .A2(n6210), .A3(n8707), .A4(n6126), .ZN(n6127)
         );
  NOR4_X1 U7624 ( .A1(n8478), .A2(n8643), .A3(n4760), .A4(n6127), .ZN(n6128)
         );
  NAND4_X1 U7625 ( .A1(n8579), .A2(n6257), .A3(n6128), .A4(n8628), .ZN(n6129)
         );
  NOR2_X1 U7626 ( .A1(n8546), .A2(n6129), .ZN(n6130) );
  NAND4_X1 U7627 ( .A1(n8507), .A2(n6130), .A3(n8567), .A4(n4779), .ZN(n6131)
         );
  NOR4_X1 U7628 ( .A1(n6132), .A2(n6135), .A3(n8492), .A4(n6131), .ZN(n6133)
         );
  XNOR2_X1 U7629 ( .A(n6133), .B(n8554), .ZN(n6134) );
  OAI22_X1 U7630 ( .A1(n6134), .A2(n7007), .B1(n6961), .B2(n6956), .ZN(n6295)
         );
  INV_X1 U7631 ( .A(n6135), .ZN(n6136) );
  MUX2_X1 U7632 ( .A(n6137), .B(n6136), .S(n6288), .Z(n6293) );
  NAND2_X1 U7633 ( .A1(n6158), .A2(n6156), .ZN(n6139) );
  NAND2_X1 U7634 ( .A1(n6117), .A2(n6140), .ZN(n6138) );
  INV_X1 U7635 ( .A(n6160), .ZN(n6148) );
  AND2_X1 U7636 ( .A1(n7033), .A2(n7007), .ZN(n6145) );
  OAI211_X1 U7637 ( .C1(n6143), .C2(n6145), .A(n6144), .B(n6149), .ZN(n6146)
         );
  NAND3_X1 U7638 ( .A1(n6146), .A2(n7428), .A3(n6288), .ZN(n6147) );
  NAND2_X1 U7639 ( .A1(n6149), .A2(n7033), .ZN(n6150) );
  NAND3_X1 U7640 ( .A1(n7428), .A2(n6151), .A3(n6150), .ZN(n6152) );
  NAND3_X1 U7641 ( .A1(n6152), .A2(n6281), .A3(n6144), .ZN(n6153) );
  AND2_X1 U7642 ( .A1(n6156), .A2(n6155), .ZN(n6159) );
  OAI211_X1 U7643 ( .C1(n6160), .C2(n6159), .A(n6158), .B(n6157), .ZN(n6161)
         );
  NAND2_X1 U7644 ( .A1(n6161), .A2(n6281), .ZN(n6162) );
  NOR2_X1 U7645 ( .A1(n6163), .A2(n6288), .ZN(n6164) );
  NOR2_X1 U7646 ( .A1(n6165), .A2(n6164), .ZN(n6166) );
  NAND2_X1 U7647 ( .A1(n6167), .A2(n6166), .ZN(n6173) );
  MUX2_X1 U7648 ( .A(n6169), .B(n6168), .S(n6288), .Z(n6170) );
  INV_X1 U7649 ( .A(n6170), .ZN(n6171) );
  NAND2_X1 U7650 ( .A1(n6173), .A2(n6172), .ZN(n6178) );
  MUX2_X1 U7651 ( .A(n6175), .B(n6174), .S(n6288), .Z(n6176) );
  NAND3_X1 U7652 ( .A1(n6178), .A2(n6177), .A3(n6176), .ZN(n6192) );
  NAND2_X1 U7653 ( .A1(n6186), .A2(n6288), .ZN(n6184) );
  INV_X1 U7654 ( .A(n6185), .ZN(n6179) );
  OR3_X1 U7655 ( .A1(n6180), .A2(n6179), .A3(n6288), .ZN(n6181) );
  OAI21_X1 U7656 ( .B1(n6182), .B2(n6184), .A(n6181), .ZN(n6191) );
  OAI211_X1 U7657 ( .C1(n6185), .C2(n6184), .A(n6183), .B(n7891), .ZN(n6189)
         );
  INV_X1 U7658 ( .A(n6186), .ZN(n6187) );
  OR2_X1 U7659 ( .A1(n6193), .A2(n6187), .ZN(n6188) );
  MUX2_X1 U7660 ( .A(n6189), .B(n6188), .S(n6281), .Z(n6190) );
  OR2_X1 U7661 ( .A1(n7875), .A2(n6193), .ZN(n6194) );
  MUX2_X1 U7662 ( .A(n6195), .B(n6194), .S(n6288), .Z(n6196) );
  MUX2_X1 U7663 ( .A(n6198), .B(n6197), .S(n6281), .Z(n6200) );
  INV_X1 U7664 ( .A(n7993), .ZN(n8459) );
  MUX2_X1 U7665 ( .A(n6202), .B(n6201), .S(n6281), .Z(n6203) );
  INV_X1 U7666 ( .A(n8725), .ZN(n6205) );
  NAND3_X1 U7667 ( .A1(n6217), .A2(n6205), .A3(n6204), .ZN(n6206) );
  NAND2_X1 U7668 ( .A1(n6206), .A2(n8705), .ZN(n6211) );
  MUX2_X1 U7669 ( .A(n6208), .B(n6207), .S(n6288), .Z(n6209) );
  NAND2_X1 U7670 ( .A1(n6210), .A2(n6209), .ZN(n6219) );
  INV_X1 U7671 ( .A(n6219), .ZN(n6225) );
  NAND2_X1 U7672 ( .A1(n6211), .A2(n6225), .ZN(n6212) );
  NAND2_X1 U7673 ( .A1(n6212), .A2(n8669), .ZN(n6222) );
  NOR2_X1 U7674 ( .A1(n8725), .A2(n6213), .ZN(n6216) );
  INV_X1 U7675 ( .A(n6214), .ZN(n6215) );
  AOI21_X1 U7676 ( .B1(n6217), .B2(n6216), .A(n6215), .ZN(n6220) );
  OAI211_X1 U7677 ( .C1(n6220), .C2(n6219), .A(n6218), .B(n6228), .ZN(n6221)
         );
  MUX2_X1 U7678 ( .A(n6222), .B(n6221), .S(n6281), .Z(n6223) );
  INV_X1 U7679 ( .A(n6223), .ZN(n6227) );
  INV_X1 U7680 ( .A(n8707), .ZN(n6224) );
  AOI21_X1 U7681 ( .B1(n6225), .B2(n6224), .A(n6231), .ZN(n6226) );
  NAND2_X1 U7682 ( .A1(n6227), .A2(n6226), .ZN(n6235) );
  NAND2_X1 U7683 ( .A1(n6235), .A2(n6228), .ZN(n6230) );
  NAND2_X1 U7684 ( .A1(n6246), .A2(n6237), .ZN(n6229) );
  AOI21_X1 U7685 ( .B1(n6230), .B2(n6232), .A(n6229), .ZN(n6240) );
  INV_X1 U7686 ( .A(n6231), .ZN(n6233) );
  NAND2_X1 U7687 ( .A1(n6235), .A2(n6234), .ZN(n6238) );
  AOI21_X1 U7688 ( .B1(n6238), .B2(n6237), .A(n6236), .ZN(n6239) );
  MUX2_X1 U7689 ( .A(n6240), .B(n6239), .S(n6281), .Z(n6251) );
  OR2_X1 U7690 ( .A1(n8807), .A2(n8645), .ZN(n6249) );
  NAND2_X1 U7691 ( .A1(n6249), .A2(n6241), .ZN(n6244) );
  INV_X1 U7692 ( .A(n6253), .ZN(n6242) );
  OAI21_X1 U7693 ( .B1(n6251), .B2(n6244), .A(n6243), .ZN(n6245) );
  NAND2_X1 U7694 ( .A1(n6245), .A2(n6252), .ZN(n6256) );
  INV_X1 U7695 ( .A(n6246), .ZN(n6247) );
  OR2_X1 U7696 ( .A1(n6248), .A2(n6247), .ZN(n6250) );
  OAI21_X1 U7697 ( .B1(n6251), .B2(n6250), .A(n6249), .ZN(n6254) );
  INV_X1 U7698 ( .A(n6252), .ZN(n8595) );
  AOI21_X1 U7699 ( .B1(n6254), .B2(n6253), .A(n8595), .ZN(n6255) );
  MUX2_X1 U7700 ( .A(n6256), .B(n6255), .S(n6281), .Z(n6260) );
  AND2_X1 U7701 ( .A1(n8579), .A2(n6258), .ZN(n6259) );
  OAI22_X1 U7702 ( .A1(n6260), .A2(n8594), .B1(n6259), .B2(n6288), .ZN(n6264)
         );
  AOI21_X1 U7703 ( .B1(n6263), .B2(n6261), .A(n6281), .ZN(n6262) );
  AOI21_X1 U7704 ( .B1(n6264), .B2(n6263), .A(n6262), .ZN(n6268) );
  OAI21_X1 U7705 ( .B1(n6281), .B2(n8566), .A(n8567), .ZN(n6267) );
  AND2_X1 U7706 ( .A1(n8788), .A2(n8295), .ZN(n6265) );
  OAI21_X1 U7707 ( .B1(n8546), .B2(n6265), .A(n6288), .ZN(n6266) );
  INV_X1 U7708 ( .A(n6269), .ZN(n8542) );
  AOI21_X1 U7709 ( .B1(n6271), .B2(n8542), .A(n6288), .ZN(n6270) );
  NOR2_X1 U7710 ( .A1(n6272), .A2(n6288), .ZN(n6273) );
  NAND3_X1 U7711 ( .A1(n8776), .A2(n8516), .A3(n6288), .ZN(n6274) );
  AND2_X1 U7712 ( .A1(n6275), .A2(n6274), .ZN(n6276) );
  AOI21_X1 U7713 ( .B1(n6278), .B2(n6277), .A(n6288), .ZN(n6280) );
  NAND3_X1 U7714 ( .A1(n8770), .A2(n8488), .A3(n6281), .ZN(n6279) );
  MUX2_X1 U7715 ( .A(n6283), .B(n6282), .S(n6281), .Z(n6284) );
  INV_X1 U7716 ( .A(n6287), .ZN(n6289) );
  MUX2_X1 U7717 ( .A(n6290), .B(n6289), .S(n6288), .Z(n6291) );
  AOI21_X1 U7718 ( .B1(n6293), .B2(n6292), .A(n6291), .ZN(n6294) );
  NAND2_X1 U7719 ( .A1(n6296), .A2(n6104), .ZN(n6297) );
  NAND2_X1 U7720 ( .A1(n6297), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U7721 ( .A1(n6299), .A2(n6298), .ZN(n6301) );
  OR2_X1 U7722 ( .A1(n6299), .A2(n6298), .ZN(n6300) );
  NAND2_X1 U7723 ( .A1(n6301), .A2(n6300), .ZN(n7057) );
  INV_X1 U7724 ( .A(n7702), .ZN(n6767) );
  NAND2_X1 U7725 ( .A1(n6301), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6303) );
  INV_X1 U7726 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U7727 ( .A1(n4372), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6304) );
  MUX2_X1 U7728 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6304), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6306) );
  NAND2_X1 U7729 ( .A1(n6306), .A2(n6305), .ZN(n7950) );
  NAND2_X1 U7730 ( .A1(n6307), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6308) );
  MUX2_X1 U7731 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6308), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6309) );
  NAND2_X1 U7732 ( .A1(n6309), .A2(n4372), .ZN(n7945) );
  INV_X1 U7733 ( .A(n9926), .ZN(n6312) );
  INV_X1 U7734 ( .A(n6783), .ZN(n8449) );
  INV_X1 U7735 ( .A(n6997), .ZN(n6311) );
  AND2_X1 U7736 ( .A1(n6950), .A2(n7007), .ZN(n7001) );
  INV_X1 U7737 ( .A(n6310), .ZN(n8001) );
  NAND4_X1 U7738 ( .A1(n6312), .A2(n8449), .A3(n6311), .A4(n8630), .ZN(n6313)
         );
  OAI211_X1 U7739 ( .C1(n6950), .C2(n6767), .A(n6313), .B(P2_B_REG_SCAN_IN), 
        .ZN(n6314) );
  NAND2_X1 U7740 ( .A1(n8888), .A2(n5009), .ZN(n6316) );
  NAND2_X1 U7741 ( .A1(n6340), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6315) );
  INV_X1 U7742 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U7743 ( .A1(n6317), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U7744 ( .A1(n6344), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6318) );
  OAI211_X1 U7745 ( .C1(n6321), .C2(n6320), .A(n6319), .B(n6318), .ZN(n9165)
         );
  INV_X1 U7746 ( .A(n9165), .ZN(n6350) );
  NAND2_X1 U7747 ( .A1(n8021), .A2(n5009), .ZN(n6323) );
  NAND2_X1 U7748 ( .A1(n6340), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6322) );
  NAND2_X1 U7749 ( .A1(n9366), .A2(n6518), .ZN(n6550) );
  NAND2_X1 U7750 ( .A1(n9389), .A2(n9135), .ZN(n6496) );
  XNOR2_X1 U7751 ( .A(n9394), .B(n9230), .ZN(n9242) );
  INV_X1 U7752 ( .A(n9242), .ZN(n6337) );
  NAND2_X1 U7753 ( .A1(n9399), .A2(n9131), .ZN(n6382) );
  NAND2_X1 U7754 ( .A1(n9153), .A2(n6382), .ZN(n9262) );
  NAND2_X1 U7755 ( .A1(n9409), .A2(n9041), .ZN(n6475) );
  INV_X1 U7756 ( .A(n9281), .ZN(n6335) );
  AND2_X1 U7757 ( .A1(n9268), .A2(n9286), .ZN(n9152) );
  NAND2_X1 U7758 ( .A1(n9404), .A2(n9130), .ZN(n9151) );
  INV_X1 U7759 ( .A(n9151), .ZN(n6324) );
  NOR2_X1 U7760 ( .A1(n9152), .A2(n6324), .ZN(n9270) );
  INV_X1 U7761 ( .A(n9312), .ZN(n9128) );
  AND2_X1 U7762 ( .A1(n9414), .A2(n9128), .ZN(n9149) );
  NOR2_X1 U7763 ( .A1(n9282), .A2(n9149), .ZN(n9300) );
  INV_X1 U7764 ( .A(n9334), .ZN(n9124) );
  OR2_X1 U7765 ( .A1(n9419), .A2(n9124), .ZN(n6469) );
  NAND2_X1 U7766 ( .A1(n9419), .A2(n9124), .ZN(n9148) );
  NAND2_X1 U7767 ( .A1(n6469), .A2(n9148), .ZN(n9310) );
  INV_X1 U7768 ( .A(n9350), .ZN(n8960) );
  OR2_X1 U7769 ( .A1(n9423), .A2(n8960), .ZN(n6468) );
  NAND2_X1 U7770 ( .A1(n9423), .A2(n8960), .ZN(n9145) );
  NAND2_X1 U7771 ( .A1(n6468), .A2(n9145), .ZN(n9331) );
  INV_X1 U7772 ( .A(n9333), .ZN(n9121) );
  OR2_X1 U7773 ( .A1(n9428), .A2(n9121), .ZN(n9329) );
  NAND2_X1 U7774 ( .A1(n9428), .A2(n9121), .ZN(n9144) );
  INV_X1 U7775 ( .A(n9339), .ZN(n9345) );
  OR2_X1 U7776 ( .A1(n9439), .A2(n7976), .ZN(n6459) );
  NAND2_X1 U7777 ( .A1(n9439), .A2(n7976), .ZN(n7970) );
  NAND2_X1 U7778 ( .A1(n9445), .A2(n9690), .ZN(n6451) );
  NAND2_X1 U7779 ( .A1(n7969), .A2(n6451), .ZN(n7829) );
  INV_X1 U7780 ( .A(n9045), .ZN(n8064) );
  XNOR2_X1 U7781 ( .A(n7753), .B(n8064), .ZN(n9708) );
  OR2_X1 U7782 ( .A1(n7816), .A2(n9711), .ZN(n6438) );
  NAND2_X1 U7783 ( .A1(n6438), .A2(n7823), .ZN(n7822) );
  INV_X1 U7784 ( .A(n6885), .ZN(n7238) );
  AND2_X1 U7785 ( .A1(n6325), .A2(n7238), .ZN(n6532) );
  NOR2_X1 U7786 ( .A1(n6917), .A2(n6532), .ZN(n6733) );
  XNOR2_X2 U7787 ( .A(n6326), .B(n6920), .ZN(n6916) );
  INV_X1 U7788 ( .A(n6916), .ZN(n6918) );
  INV_X1 U7789 ( .A(n6889), .ZN(n6397) );
  NAND2_X1 U7790 ( .A1(n4993), .A2(n7267), .ZN(n6537) );
  NAND4_X1 U7791 ( .A1(n6733), .A2(n6918), .A3(n6397), .A4(n6537), .ZN(n6329)
         );
  NAND2_X1 U7792 ( .A1(n7322), .A2(n9023), .ZN(n6425) );
  NAND2_X1 U7793 ( .A1(n7220), .A2(n7286), .ZN(n6422) );
  NAND2_X1 U7794 ( .A1(n6425), .A2(n6422), .ZN(n6400) );
  NAND2_X1 U7795 ( .A1(n7113), .A2(n8978), .ZN(n7120) );
  INV_X1 U7796 ( .A(n7120), .ZN(n6419) );
  OR2_X1 U7797 ( .A1(n6400), .A2(n6419), .ZN(n6539) );
  NAND2_X1 U7798 ( .A1(n9050), .A2(n7230), .ZN(n6426) );
  NAND2_X1 U7799 ( .A1(n6426), .A2(n6421), .ZN(n6327) );
  NAND2_X1 U7800 ( .A1(n6425), .A2(n6327), .ZN(n7136) );
  INV_X1 U7801 ( .A(n7113), .ZN(n9052) );
  NAND2_X1 U7802 ( .A1(n9052), .A2(n9847), .ZN(n7135) );
  INV_X1 U7803 ( .A(n4993), .ZN(n9053) );
  NAND2_X1 U7804 ( .A1(n9053), .A2(n7264), .ZN(n6417) );
  AND2_X1 U7805 ( .A1(n7135), .A2(n6417), .ZN(n6328) );
  NAND2_X1 U7806 ( .A1(n7136), .A2(n6328), .ZN(n6393) );
  NAND2_X1 U7807 ( .A1(n7336), .A2(n7243), .ZN(n7332) );
  NAND2_X1 U7808 ( .A1(n7328), .A2(n9049), .ZN(n6427) );
  NAND2_X1 U7809 ( .A1(n7332), .A2(n6427), .ZN(n7141) );
  NOR4_X1 U7810 ( .A1(n6329), .A2(n6539), .A3(n6393), .A4(n7141), .ZN(n6330)
         );
  OR2_X1 U7811 ( .A1(n9671), .A2(n9713), .ZN(n6437) );
  NAND2_X1 U7812 ( .A1(n9671), .A2(n9713), .ZN(n6432) );
  NAND2_X1 U7813 ( .A1(n6437), .A2(n6432), .ZN(n7743) );
  INV_X1 U7814 ( .A(n7743), .ZN(n7477) );
  INV_X1 U7815 ( .A(n9047), .ZN(n7337) );
  OR2_X1 U7816 ( .A1(n9886), .A2(n7337), .ZN(n7482) );
  NAND2_X1 U7817 ( .A1(n9886), .A2(n7337), .ZN(n7481) );
  AND2_X1 U7818 ( .A1(n7482), .A2(n7481), .ZN(n8074) );
  OR2_X1 U7819 ( .A1(n8076), .A2(n8926), .ZN(n7478) );
  NAND2_X1 U7820 ( .A1(n8926), .A2(n8076), .ZN(n7480) );
  NAND4_X1 U7821 ( .A1(n6330), .A2(n7477), .A3(n8074), .A4(n7334), .ZN(n6331)
         );
  NOR4_X1 U7822 ( .A1(n7829), .A2(n9708), .A3(n7822), .A4(n6331), .ZN(n6332)
         );
  XNOR2_X1 U7823 ( .A(n9697), .B(n8040), .ZN(n9680) );
  INV_X1 U7824 ( .A(n9680), .ZN(n9688) );
  NAND4_X1 U7825 ( .A1(n8008), .A2(n9142), .A3(n6332), .A4(n9688), .ZN(n6333)
         );
  NOR4_X1 U7826 ( .A1(n9310), .A2(n9331), .A3(n9345), .A4(n6333), .ZN(n6334)
         );
  NAND4_X1 U7827 ( .A1(n6335), .A2(n9270), .A3(n9300), .A4(n6334), .ZN(n6336)
         );
  OR4_X1 U7828 ( .A1(n9227), .A2(n6337), .A3(n9262), .A4(n6336), .ZN(n6339) );
  INV_X1 U7829 ( .A(n9138), .ZN(n6338) );
  NAND2_X1 U7830 ( .A1(n9379), .A2(n9139), .ZN(n6506) );
  NOR4_X1 U7831 ( .A1(n6339), .A2(n9210), .A3(n9200), .A4(n9179), .ZN(n6348)
         );
  NAND2_X1 U7832 ( .A1(n8884), .A2(n5009), .ZN(n6342) );
  NAND2_X1 U7833 ( .A1(n6340), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n6341) );
  NAND2_X1 U7834 ( .A1(n6343), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6347) );
  NAND2_X1 U7835 ( .A1(n5084), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U7836 ( .A1(n6344), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6345) );
  NAND3_X1 U7837 ( .A1(n6347), .A2(n6346), .A3(n6345), .ZN(n8113) );
  INV_X1 U7838 ( .A(n8113), .ZN(n6349) );
  NAND2_X1 U7839 ( .A1(n9357), .A2(n6349), .ZN(n6557) );
  NAND4_X1 U7840 ( .A1(n6554), .A2(n9161), .A3(n6348), .A4(n6557), .ZN(n6352)
         );
  NAND2_X1 U7841 ( .A1(n9360), .A2(n6350), .ZN(n6351) );
  NAND2_X1 U7842 ( .A1(n6523), .A2(n6351), .ZN(n6556) );
  OAI21_X1 U7843 ( .B1(n6352), .B2(n6556), .A(n5628), .ZN(n6525) );
  INV_X1 U7844 ( .A(n6525), .ZN(n6414) );
  INV_X1 U7845 ( .A(n6415), .ZN(n6519) );
  INV_X1 U7846 ( .A(n9203), .ZN(n9224) );
  NAND2_X1 U7847 ( .A1(n9383), .A2(n9224), .ZN(n9156) );
  INV_X1 U7848 ( .A(n9156), .ZN(n6353) );
  NAND2_X1 U7849 ( .A1(n9158), .A2(n6353), .ZN(n6354) );
  AND2_X1 U7850 ( .A1(n6354), .A2(n6506), .ZN(n6355) );
  NAND2_X1 U7851 ( .A1(n6355), .A2(n9160), .ZN(n6546) );
  OR2_X1 U7852 ( .A1(n9383), .A2(n9224), .ZN(n6356) );
  NAND2_X1 U7853 ( .A1(n6356), .A2(n6498), .ZN(n9157) );
  NAND2_X1 U7854 ( .A1(n9240), .A2(n9230), .ZN(n6383) );
  AND2_X1 U7855 ( .A1(n6383), .A2(n9153), .ZN(n6483) );
  INV_X1 U7856 ( .A(n6483), .ZN(n6381) );
  INV_X1 U7857 ( .A(n6360), .ZN(n6357) );
  OR2_X1 U7858 ( .A1(n9152), .A2(n6357), .ZN(n6481) );
  AND2_X1 U7859 ( .A1(n6468), .A2(n9329), .ZN(n9147) );
  AND2_X1 U7860 ( .A1(n9148), .A2(n9145), .ZN(n6465) );
  INV_X1 U7861 ( .A(n6465), .ZN(n6359) );
  INV_X1 U7862 ( .A(n6469), .ZN(n6358) );
  NOR2_X1 U7863 ( .A1(n9282), .A2(n6358), .ZN(n6466) );
  OAI21_X1 U7864 ( .B1(n9147), .B2(n6359), .A(n6466), .ZN(n6364) );
  INV_X1 U7865 ( .A(n9152), .ZN(n6363) );
  NAND2_X1 U7866 ( .A1(n6360), .A2(n9149), .ZN(n6361) );
  AND2_X1 U7867 ( .A1(n6361), .A2(n6475), .ZN(n6362) );
  NAND2_X1 U7868 ( .A1(n9151), .A2(n6362), .ZN(n6365) );
  NAND2_X1 U7869 ( .A1(n6363), .A2(n6365), .ZN(n6479) );
  OAI21_X1 U7870 ( .B1(n6481), .B2(n6364), .A(n6479), .ZN(n6379) );
  INV_X1 U7871 ( .A(n6365), .ZN(n6391) );
  AND2_X1 U7872 ( .A1(n9145), .A2(n9144), .ZN(n6463) );
  INV_X1 U7873 ( .A(n6463), .ZN(n6407) );
  INV_X1 U7874 ( .A(n7970), .ZN(n6366) );
  OR2_X1 U7875 ( .A1(n9141), .A2(n6366), .ZN(n6457) );
  INV_X1 U7876 ( .A(n6457), .ZN(n6390) );
  NAND2_X1 U7877 ( .A1(n7753), .A2(n8064), .ZN(n7755) );
  INV_X1 U7878 ( .A(n6437), .ZN(n6367) );
  NAND2_X1 U7879 ( .A1(n7482), .A2(n7478), .ZN(n6435) );
  NAND2_X1 U7880 ( .A1(n6432), .A2(n7481), .ZN(n6439) );
  NAND2_X1 U7881 ( .A1(n6439), .A2(n6437), .ZN(n7751) );
  OAI21_X1 U7882 ( .B1(n6367), .B2(n6435), .A(n7751), .ZN(n6368) );
  NOR2_X1 U7883 ( .A1(n6405), .A2(n6368), .ZN(n6373) );
  OAI21_X1 U7884 ( .B1(n7822), .B2(n9708), .A(n6369), .ZN(n6370) );
  INV_X1 U7885 ( .A(n8040), .ZN(n9043) );
  NAND2_X1 U7886 ( .A1(n9729), .A2(n9043), .ZN(n6450) );
  AND2_X1 U7887 ( .A1(n6370), .A2(n6450), .ZN(n6443) );
  INV_X1 U7888 ( .A(n6443), .ZN(n6372) );
  NAND2_X1 U7889 ( .A1(n9697), .A2(n8040), .ZN(n7827) );
  NAND2_X1 U7890 ( .A1(n6451), .A2(n7827), .ZN(n6449) );
  INV_X1 U7891 ( .A(n6449), .ZN(n6371) );
  OAI21_X1 U7892 ( .B1(n6373), .B2(n6372), .A(n6371), .ZN(n6374) );
  NAND3_X1 U7893 ( .A1(n6374), .A2(n6459), .A3(n7969), .ZN(n6375) );
  AOI21_X1 U7894 ( .B1(n6390), .B2(n6375), .A(n6458), .ZN(n6376) );
  NOR2_X1 U7895 ( .A1(n6407), .A2(n6376), .ZN(n6377) );
  NAND3_X1 U7896 ( .A1(n6391), .A2(n6377), .A3(n9148), .ZN(n6378) );
  NAND2_X1 U7897 ( .A1(n6379), .A2(n6378), .ZN(n6380) );
  NOR2_X1 U7898 ( .A1(n6381), .A2(n6380), .ZN(n6386) );
  NAND2_X1 U7899 ( .A1(n9394), .A2(n9259), .ZN(n9155) );
  AND2_X1 U7900 ( .A1(n9155), .A2(n6382), .ZN(n6480) );
  INV_X1 U7901 ( .A(n6480), .ZN(n6384) );
  NAND2_X1 U7902 ( .A1(n6384), .A2(n6383), .ZN(n6385) );
  NAND2_X1 U7903 ( .A1(n6496), .A2(n6385), .ZN(n6488) );
  NOR2_X1 U7904 ( .A1(n6386), .A2(n6488), .ZN(n6387) );
  NOR2_X1 U7905 ( .A1(n9157), .A2(n6387), .ZN(n6389) );
  OAI211_X1 U7906 ( .C1(n6546), .C2(n6389), .A(n6388), .B(n6509), .ZN(n6551)
         );
  NAND3_X1 U7907 ( .A1(n6391), .A2(n6390), .A3(n9148), .ZN(n6392) );
  OR3_X1 U7908 ( .A1(n6546), .A2(n6488), .A3(n6392), .ZN(n6549) );
  INV_X1 U7909 ( .A(n6427), .ZN(n6545) );
  INV_X1 U7910 ( .A(n6393), .ZN(n6541) );
  NAND2_X1 U7911 ( .A1(n6918), .A2(n6917), .ZN(n6396) );
  INV_X1 U7912 ( .A(n6326), .ZN(n6394) );
  INV_X1 U7913 ( .A(n6920), .ZN(n7094) );
  NAND2_X1 U7914 ( .A1(n6394), .A2(n7094), .ZN(n6395) );
  NAND2_X1 U7915 ( .A1(n6531), .A2(n6397), .ZN(n6398) );
  INV_X1 U7916 ( .A(n9054), .ZN(n7116) );
  NAND2_X1 U7917 ( .A1(n7116), .A2(n6872), .ZN(n6536) );
  NAND2_X1 U7918 ( .A1(n6398), .A2(n6536), .ZN(n7256) );
  INV_X1 U7919 ( .A(n6537), .ZN(n6399) );
  OAI211_X1 U7920 ( .C1(n6419), .C2(n6399), .A(n6421), .B(n7135), .ZN(n6402)
         );
  INV_X1 U7921 ( .A(n6400), .ZN(n6401) );
  NAND2_X1 U7922 ( .A1(n6402), .A2(n6401), .ZN(n6403) );
  AOI22_X1 U7923 ( .A1(n6541), .A2(n7256), .B1(n6403), .B2(n6426), .ZN(n6408)
         );
  NAND3_X1 U7924 ( .A1(n7751), .A2(n7480), .A3(n7332), .ZN(n6404) );
  OR3_X1 U7925 ( .A1(n6449), .A2(n6405), .A3(n6404), .ZN(n6406) );
  NOR2_X1 U7926 ( .A1(n6407), .A2(n6406), .ZN(n6543) );
  OAI21_X1 U7927 ( .B1(n6545), .B2(n6408), .A(n6543), .ZN(n6409) );
  OAI22_X1 U7928 ( .A1(n6549), .A2(n6409), .B1(n9158), .B2(n6546), .ZN(n6411)
         );
  NAND2_X1 U7929 ( .A1(n8113), .A2(n9165), .ZN(n6410) );
  NAND2_X1 U7930 ( .A1(n9360), .A2(n6410), .ZN(n6516) );
  OAI211_X1 U7931 ( .C1(n6551), .C2(n6411), .A(n6516), .B(n6550), .ZN(n6412)
         );
  INV_X1 U7932 ( .A(n6523), .ZN(n6527) );
  AOI211_X1 U7933 ( .C1(n6519), .C2(n6412), .A(n5628), .B(n6527), .ZN(n6413)
         );
  NOR2_X1 U7934 ( .A1(n6414), .A2(n6413), .ZN(n6526) );
  INV_X1 U7935 ( .A(n6517), .ZN(n6521) );
  NAND2_X1 U7936 ( .A1(n6557), .A2(n6521), .ZN(n6514) );
  NOR2_X1 U7937 ( .A1(n6415), .A2(n9174), .ZN(n6416) );
  MUX2_X1 U7938 ( .A(n6416), .B(n9188), .S(n6517), .Z(n6512) );
  NAND2_X1 U7939 ( .A1(n6537), .A2(n6417), .ZN(n7261) );
  INV_X1 U7940 ( .A(n7261), .ZN(n7255) );
  NAND2_X1 U7941 ( .A1(n7256), .A2(n7255), .ZN(n6418) );
  NAND2_X1 U7942 ( .A1(n6418), .A2(n6537), .ZN(n7187) );
  OR2_X1 U7943 ( .A1(n7187), .A2(n6419), .ZN(n6420) );
  AND2_X1 U7944 ( .A1(n6420), .A2(n7135), .ZN(n7274) );
  NAND2_X1 U7945 ( .A1(n6421), .A2(n6422), .ZN(n7114) );
  INV_X1 U7946 ( .A(n7114), .ZN(n7279) );
  NAND2_X1 U7947 ( .A1(n7274), .A2(n7279), .ZN(n7273) );
  NAND2_X1 U7948 ( .A1(n7273), .A2(n6422), .ZN(n7219) );
  NAND2_X1 U7949 ( .A1(n7219), .A2(n6426), .ZN(n6424) );
  AND2_X1 U7950 ( .A1(n7332), .A2(n6425), .ZN(n6423) );
  AOI21_X1 U7951 ( .B1(n6424), .B2(n6423), .A(n6545), .ZN(n6430) );
  AND2_X1 U7952 ( .A1(n6425), .A2(n6426), .ZN(n7123) );
  INV_X1 U7953 ( .A(n7123), .ZN(n7226) );
  OR2_X1 U7954 ( .A1(n7219), .A2(n7226), .ZN(n7222) );
  AND2_X1 U7955 ( .A1(n6427), .A2(n6426), .ZN(n6428) );
  AOI21_X1 U7956 ( .B1(n7222), .B2(n6428), .A(n4653), .ZN(n6429) );
  MUX2_X1 U7957 ( .A(n6430), .B(n6429), .S(n6517), .Z(n6436) );
  NAND2_X1 U7958 ( .A1(n7481), .A2(n7480), .ZN(n6431) );
  AOI21_X1 U7959 ( .B1(n6436), .B2(n7478), .A(n6431), .ZN(n6434) );
  AND2_X1 U7960 ( .A1(n6437), .A2(n7482), .ZN(n7750) );
  INV_X1 U7961 ( .A(n7750), .ZN(n6433) );
  OAI211_X1 U7962 ( .C1(n6434), .C2(n6433), .A(n7823), .B(n6432), .ZN(n6442)
         );
  AOI21_X1 U7963 ( .B1(n6436), .B2(n7480), .A(n6435), .ZN(n6440) );
  OAI211_X1 U7964 ( .C1(n6440), .C2(n6439), .A(n6438), .B(n6437), .ZN(n6441)
         );
  MUX2_X1 U7965 ( .A(n6442), .B(n6441), .S(n6517), .Z(n6448) );
  AND2_X1 U7966 ( .A1(n6443), .A2(n7969), .ZN(n6446) );
  NOR2_X1 U7967 ( .A1(n6449), .A2(n6444), .ZN(n6445) );
  MUX2_X1 U7968 ( .A(n6446), .B(n6445), .S(n6517), .Z(n6447) );
  OAI21_X1 U7969 ( .B1(n6448), .B2(n9708), .A(n6447), .ZN(n6456) );
  NAND2_X1 U7970 ( .A1(n6449), .A2(n7969), .ZN(n6454) );
  NAND2_X1 U7971 ( .A1(n7969), .A2(n6450), .ZN(n6452) );
  NAND2_X1 U7972 ( .A1(n6452), .A2(n6451), .ZN(n6453) );
  MUX2_X1 U7973 ( .A(n6454), .B(n6453), .S(n6517), .Z(n6455) );
  INV_X1 U7974 ( .A(n6458), .ZN(n6460) );
  AOI21_X1 U7975 ( .B1(n6460), .B2(n6459), .A(n6517), .ZN(n6462) );
  NAND2_X1 U7976 ( .A1(n9141), .A2(n6521), .ZN(n6461) );
  MUX2_X1 U7977 ( .A(n9147), .B(n6463), .S(n6517), .Z(n6464) );
  NAND2_X1 U7978 ( .A1(n6470), .A2(n6465), .ZN(n6467) );
  NAND2_X1 U7979 ( .A1(n6467), .A2(n6466), .ZN(n6474) );
  NAND3_X1 U7980 ( .A1(n6470), .A2(n6469), .A3(n6468), .ZN(n6472) );
  INV_X1 U7981 ( .A(n9149), .ZN(n6471) );
  NAND3_X1 U7982 ( .A1(n6472), .A2(n6471), .A3(n9148), .ZN(n6473) );
  INV_X1 U7983 ( .A(n9282), .ZN(n6476) );
  INV_X1 U7984 ( .A(n6475), .ZN(n9150) );
  AOI21_X1 U7985 ( .B1(n6482), .B2(n6476), .A(n9150), .ZN(n6477) );
  OAI21_X1 U7986 ( .B1(n6477), .B2(n6481), .A(n9151), .ZN(n6478) );
  NAND2_X1 U7987 ( .A1(n6478), .A2(n6483), .ZN(n6487) );
  NAND2_X1 U7988 ( .A1(n6484), .A2(n6483), .ZN(n6485) );
  INV_X1 U7989 ( .A(n6498), .ZN(n9208) );
  AOI21_X1 U7990 ( .B1(n6485), .B2(n9155), .A(n9208), .ZN(n6486) );
  MUX2_X1 U7991 ( .A(n6487), .B(n6486), .S(n6521), .Z(n6490) );
  NAND2_X1 U7992 ( .A1(n6488), .A2(n6517), .ZN(n6489) );
  NAND2_X1 U7993 ( .A1(n6490), .A2(n6489), .ZN(n6503) );
  NAND2_X1 U7994 ( .A1(n9383), .A2(n6498), .ZN(n6491) );
  NAND2_X1 U7995 ( .A1(n6506), .A2(n6491), .ZN(n6494) );
  NAND2_X1 U7996 ( .A1(n6496), .A2(n9203), .ZN(n6492) );
  NAND2_X1 U7997 ( .A1(n9158), .A2(n6492), .ZN(n6493) );
  MUX2_X1 U7998 ( .A(n6494), .B(n6493), .S(n6521), .Z(n6495) );
  OAI21_X1 U7999 ( .B1(n6503), .B2(n9200), .A(n6495), .ZN(n6505) );
  NOR2_X1 U8000 ( .A1(n6496), .A2(n9203), .ZN(n6497) );
  NOR2_X1 U8001 ( .A1(n6497), .A2(n9383), .ZN(n6501) );
  NAND2_X1 U8002 ( .A1(n6498), .A2(n9224), .ZN(n6499) );
  NAND2_X1 U8003 ( .A1(n9156), .A2(n6499), .ZN(n6500) );
  MUX2_X1 U8004 ( .A(n6501), .B(n6500), .S(n6517), .Z(n6502) );
  OAI21_X1 U8005 ( .B1(n6503), .B2(n9137), .A(n6502), .ZN(n6504) );
  NAND2_X1 U8006 ( .A1(n6505), .A2(n6504), .ZN(n6508) );
  MUX2_X1 U8007 ( .A(n6506), .B(n9158), .S(n6517), .Z(n6507) );
  NAND3_X1 U8008 ( .A1(n6508), .A2(n9187), .A3(n6507), .ZN(n6511) );
  MUX2_X1 U8009 ( .A(n9160), .B(n6509), .S(n6521), .Z(n6510) );
  AND2_X2 U8010 ( .A1(n6511), .A2(n6510), .ZN(n6515) );
  NAND2_X1 U8011 ( .A1(n6512), .A2(n6515), .ZN(n6513) );
  MUX2_X1 U8012 ( .A(n6514), .B(n6513), .S(n6516), .Z(n6524) );
  MUX2_X1 U8013 ( .A(n6521), .B(n6520), .S(n6519), .Z(n6522) );
  INV_X1 U8014 ( .A(n6895), .ZN(n6734) );
  NOR3_X1 U8015 ( .A1(n6527), .A2(n7538), .A3(n5628), .ZN(n6528) );
  NAND2_X1 U8016 ( .A1(n6529), .A2(n6528), .ZN(n6530) );
  AOI21_X1 U8017 ( .B1(n6326), .B2(n6920), .A(n5628), .ZN(n6534) );
  INV_X1 U8018 ( .A(n6532), .ZN(n6533) );
  AND2_X1 U8019 ( .A1(n6534), .A2(n6533), .ZN(n6535) );
  OAI22_X1 U8020 ( .A1(n6531), .A2(n6535), .B1(n7116), .B2(n6872), .ZN(n6538)
         );
  NAND3_X1 U8021 ( .A1(n6538), .A2(n6537), .A3(n6536), .ZN(n6542) );
  NAND2_X1 U8022 ( .A1(n6539), .A2(n7136), .ZN(n7140) );
  INV_X1 U8023 ( .A(n7140), .ZN(n6540) );
  AOI21_X1 U8024 ( .B1(n6542), .B2(n6541), .A(n6540), .ZN(n6544) );
  OAI21_X1 U8025 ( .B1(n6545), .B2(n6544), .A(n6543), .ZN(n6548) );
  INV_X1 U8026 ( .A(n9200), .ZN(n6547) );
  OAI22_X1 U8027 ( .A1(n6549), .A2(n6548), .B1(n6547), .B2(n6546), .ZN(n6552)
         );
  OAI21_X1 U8028 ( .B1(n6552), .B2(n6551), .A(n6550), .ZN(n6553) );
  AND2_X1 U8029 ( .A1(n6554), .A2(n6553), .ZN(n6555) );
  NAND2_X1 U8030 ( .A1(n6558), .A2(n6557), .ZN(n6562) );
  NAND2_X1 U8031 ( .A1(n9110), .A2(n7093), .ZN(n6561) );
  INV_X1 U8032 ( .A(n7199), .ZN(n6559) );
  NAND2_X1 U8033 ( .A1(n6562), .A2(n6559), .ZN(n6560) );
  NOR2_X1 U8034 ( .A1(n6572), .A2(P1_U3084), .ZN(n7704) );
  OAI211_X1 U8035 ( .C1(n6562), .C2(n6561), .A(n6560), .B(n7704), .ZN(n6563)
         );
  INV_X1 U8036 ( .A(n6563), .ZN(n6564) );
  INV_X1 U8037 ( .A(n7704), .ZN(n6567) );
  INV_X1 U8038 ( .A(n9837), .ZN(n6641) );
  INV_X1 U8039 ( .A(n6565), .ZN(n6650) );
  NAND4_X1 U8040 ( .A1(n6732), .A2(n6641), .A3(n6894), .A4(n6650), .ZN(n6566)
         );
  OAI211_X1 U8041 ( .C1(n7538), .C2(n6567), .A(n6566), .B(P1_B_REG_SCAN_IN), 
        .ZN(n6568) );
  NAND2_X1 U8042 ( .A1(n6569), .A2(n6568), .ZN(P1_U3240) );
  INV_X1 U8043 ( .A(n6572), .ZN(n6570) );
  NOR2_X1 U8044 ( .A1(n4904), .A2(n6570), .ZN(n6610) );
  INV_X1 U8045 ( .A(n9937), .ZN(n6571) );
  INV_X2 U8046 ( .A(n8353), .ZN(P2_U3966) );
  NAND2_X1 U8047 ( .A1(n4904), .A2(n6734), .ZN(n6573) );
  NAND2_X1 U8048 ( .A1(n6573), .A2(n6572), .ZN(n6608) );
  NAND2_X1 U8049 ( .A1(n6608), .A2(n6574), .ZN(n6655) );
  NAND2_X1 U8050 ( .A1(n6655), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AND2_X1 U8051 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7533) );
  NOR2_X1 U8052 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6691), .ZN(n6588) );
  INV_X1 U8053 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7146) );
  MUX2_X1 U8054 ( .A(n7146), .B(P1_REG2_REG_7__SCAN_IN), .S(n6691), .Z(n6689)
         );
  NAND2_X1 U8055 ( .A1(n6634), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6587) );
  NOR2_X1 U8056 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9783), .ZN(n6585) );
  INV_X1 U8057 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6575) );
  MUX2_X1 U8058 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6575), .S(n9750), .Z(n6579)
         );
  INV_X1 U8059 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6576) );
  MUX2_X1 U8060 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6576), .S(n6725), .Z(n6577)
         );
  AND2_X1 U8061 ( .A1(n9655), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6724) );
  NAND2_X1 U8062 ( .A1(n6577), .A2(n6724), .ZN(n6726) );
  NAND2_X1 U8063 ( .A1(n4300), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6578) );
  NAND2_X1 U8064 ( .A1(n6726), .A2(n6578), .ZN(n9751) );
  NAND2_X1 U8065 ( .A1(n6579), .A2(n9751), .ZN(n9755) );
  NAND2_X1 U8066 ( .A1(n9750), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6674) );
  NAND2_X1 U8067 ( .A1(n9755), .A2(n6674), .ZN(n6582) );
  INV_X1 U8068 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6580) );
  MUX2_X1 U8069 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6580), .S(n6673), .Z(n6581)
         );
  NAND2_X1 U8070 ( .A1(n6582), .A2(n6581), .ZN(n6677) );
  NAND2_X1 U8071 ( .A1(n6673), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6583) );
  INV_X1 U8072 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6584) );
  MUX2_X1 U8073 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6584), .S(n9769), .Z(n9766)
         );
  NAND2_X1 U8074 ( .A1(n9767), .A2(n9766), .ZN(n9765) );
  OAI21_X1 U8075 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9769), .A(n9765), .ZN(
        n9785) );
  INV_X1 U8076 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7284) );
  MUX2_X1 U8077 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7284), .S(n9783), .Z(n9784)
         );
  NOR2_X1 U8078 ( .A1(n6585), .A2(n9787), .ZN(n6710) );
  INV_X1 U8079 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6586) );
  MUX2_X1 U8080 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6586), .S(n6634), .Z(n6709)
         );
  NAND2_X1 U8081 ( .A1(n6710), .A2(n6709), .ZN(n6708) );
  NAND2_X1 U8082 ( .A1(n6980), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6589) );
  OAI21_X1 U8083 ( .B1(n6980), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6589), .ZN(
        n6590) );
  NOR2_X1 U8084 ( .A1(n9799), .A2(n6590), .ZN(n6979) );
  NOR2_X1 U8085 ( .A1(n6565), .A2(P1_U3084), .ZN(n7965) );
  NAND2_X1 U8086 ( .A1(n6608), .A2(n7965), .ZN(n9107) );
  INV_X1 U8087 ( .A(n9107), .ZN(n9806) );
  AND2_X1 U8088 ( .A1(n9806), .A2(n6894), .ZN(n9798) );
  INV_X1 U8089 ( .A(n9798), .ZN(n9817) );
  AOI211_X1 U8090 ( .C1(n9799), .C2(n6590), .A(n6979), .B(n9817), .ZN(n6614)
         );
  NOR2_X1 U8091 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6691), .ZN(n6602) );
  NOR2_X1 U8092 ( .A1(n6634), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6600) );
  NAND2_X1 U8093 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9783), .ZN(n6599) );
  INV_X1 U8094 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6591) );
  MUX2_X1 U8095 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6591), .S(n9750), .Z(n9760)
         );
  INV_X1 U8096 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6592) );
  MUX2_X1 U8097 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6592), .S(n4300), .Z(n6593)
         );
  AND2_X1 U8098 ( .A1(n9655), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6720) );
  NAND2_X1 U8099 ( .A1(n6593), .A2(n6720), .ZN(n6718) );
  NAND2_X1 U8100 ( .A1(n4300), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6594) );
  NAND2_X1 U8101 ( .A1(n6718), .A2(n6594), .ZN(n9761) );
  NAND2_X1 U8102 ( .A1(n9760), .A2(n9761), .ZN(n9759) );
  NAND2_X1 U8103 ( .A1(n9750), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U8104 ( .A1(n9759), .A2(n6669), .ZN(n6597) );
  INV_X1 U8105 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6595) );
  MUX2_X1 U8106 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6595), .S(n6673), .Z(n6596)
         );
  NAND2_X1 U8107 ( .A1(n6597), .A2(n6596), .ZN(n6671) );
  NAND2_X1 U8108 ( .A1(n6673), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6598) );
  AND2_X1 U8109 ( .A1(n6671), .A2(n6598), .ZN(n9776) );
  INV_X1 U8110 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9899) );
  MUX2_X1 U8111 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9899), .S(n9769), .Z(n9777)
         );
  NAND2_X1 U8112 ( .A1(n9776), .A2(n9777), .ZN(n9775) );
  OAI21_X1 U8113 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9769), .A(n9775), .ZN(
        n9789) );
  INV_X1 U8114 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9901) );
  MUX2_X1 U8115 ( .A(n9901), .B(P1_REG1_REG_5__SCAN_IN), .S(n9783), .Z(n9788)
         );
  NAND2_X1 U8116 ( .A1(n6599), .A2(n9791), .ZN(n6704) );
  INV_X1 U8117 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9903) );
  INV_X1 U8118 ( .A(n6634), .ZN(n6706) );
  AOI22_X1 U8119 ( .A1(n6634), .A2(n9903), .B1(P1_REG1_REG_6__SCAN_IN), .B2(
        n6706), .ZN(n6703) );
  NOR2_X1 U8120 ( .A1(n6704), .A2(n6703), .ZN(n6702) );
  NOR2_X1 U8121 ( .A1(n6600), .A2(n6702), .ZN(n6687) );
  INV_X1 U8122 ( .A(n6691), .ZN(n6601) );
  INV_X1 U8123 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9905) );
  AOI22_X1 U8124 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6601), .B1(n6691), .B2(
        n9905), .ZN(n6686) );
  NOR2_X1 U8125 ( .A1(n6687), .A2(n6686), .ZN(n6685) );
  NOR2_X1 U8126 ( .A1(n6602), .A2(n6685), .ZN(n9805) );
  INV_X1 U8127 ( .A(n9805), .ZN(n6603) );
  INV_X1 U8128 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9907) );
  NOR2_X1 U8129 ( .A1(n6603), .A2(n9907), .ZN(n6604) );
  OAI22_X1 U8130 ( .A1(n6604), .A2(n9807), .B1(P1_REG1_REG_8__SCAN_IN), .B2(
        n9805), .ZN(n9803) );
  INV_X1 U8131 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6605) );
  MUX2_X1 U8132 ( .A(n6605), .B(P1_REG1_REG_9__SCAN_IN), .S(n6611), .Z(n6606)
         );
  NAND2_X1 U8133 ( .A1(n9803), .A2(n6606), .ZN(n6972) );
  OAI21_X1 U8134 ( .B1(n9803), .B2(n6606), .A(n6972), .ZN(n6609) );
  OR2_X1 U8135 ( .A1(n5639), .A2(P1_U3084), .ZN(n8004) );
  NOR2_X1 U8136 ( .A1(n8004), .A2(n6650), .ZN(n6607) );
  AND2_X1 U8137 ( .A1(n6608), .A2(n6607), .ZN(n9823) );
  AND2_X1 U8138 ( .A1(n6609), .A2(n9823), .ZN(n6613) );
  AND2_X1 U8139 ( .A1(n9806), .A2(n5639), .ZN(n9825) );
  INV_X1 U8140 ( .A(n9825), .ZN(n9060) );
  OR2_X1 U8141 ( .A1(P1_U3083), .A2(n6610), .ZN(n9773) );
  INV_X1 U8142 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10041) );
  OAI22_X1 U8143 ( .A1(n9060), .A2(n6611), .B1(n9773), .B2(n10041), .ZN(n6612)
         );
  OR4_X1 U8144 ( .A1(n7533), .A2(n6614), .A3(n6613), .A4(n6612), .ZN(P1_U3250)
         );
  NOR2_X1 U8145 ( .A1(n5327), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9647) );
  INV_X1 U8146 ( .A(n9647), .ZN(n6627) );
  INV_X1 U8147 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6615) );
  INV_X1 U8148 ( .A(n4300), .ZN(n6723) );
  OAI222_X1 U8149 ( .A1(n6627), .A2(n6615), .B1(n9653), .B2(n6618), .C1(
        P1_U3084), .C2(n6723), .ZN(P1_U3352) );
  NOR2_X1 U8150 ( .A1(n6616), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8889) );
  INV_X1 U8151 ( .A(n8889), .ZN(n8197) );
  INV_X1 U8152 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6619) );
  INV_X1 U8153 ( .A(n7047), .ZN(n6781) );
  OAI222_X1 U8154 ( .A1(n8197), .A2(n6619), .B1(n8195), .B2(n6618), .C1(
        P2_U3152), .C2(n6781), .ZN(P2_U3357) );
  INV_X1 U8155 ( .A(n6806), .ZN(n6790) );
  OAI222_X1 U8156 ( .A1(n8197), .A2(n6620), .B1(n8195), .B2(n6633), .C1(
        P2_U3152), .C2(n6790), .ZN(P2_U3355) );
  INV_X1 U8157 ( .A(n6782), .ZN(n9661) );
  OAI222_X1 U8158 ( .A1(n8197), .A2(n6621), .B1(n8195), .B2(n6631), .C1(
        P2_U3152), .C2(n9661), .ZN(P2_U3356) );
  INV_X1 U8159 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6622) );
  INV_X1 U8160 ( .A(n6804), .ZN(n6839) );
  OAI222_X1 U8161 ( .A1(n8197), .A2(n6622), .B1(n8195), .B2(n6629), .C1(
        P2_U3152), .C2(n6839), .ZN(P2_U3354) );
  INV_X1 U8162 ( .A(n6802), .ZN(n6864) );
  OAI222_X1 U8163 ( .A1(n8197), .A2(n6623), .B1(n8195), .B2(n6625), .C1(
        P2_U3152), .C2(n6864), .ZN(P2_U3353) );
  INV_X1 U8164 ( .A(n9783), .ZN(n6624) );
  OAI222_X1 U8165 ( .A1(n6627), .A2(n6626), .B1(n9653), .B2(n6625), .C1(
        P1_U3084), .C2(n6624), .ZN(P1_U3348) );
  INV_X1 U8166 ( .A(n6627), .ZN(n9650) );
  AOI22_X1 U8167 ( .A1(n9650), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9769), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6628) );
  OAI21_X1 U8168 ( .B1(n6629), .B2(n9653), .A(n6628), .ZN(P1_U3349) );
  AOI22_X1 U8169 ( .A1(n9650), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n9750), .ZN(n6630) );
  OAI21_X1 U8170 ( .B1(n6631), .B2(n9653), .A(n6630), .ZN(P1_U3351) );
  AOI22_X1 U8171 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n9650), .B1(n6673), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6632) );
  OAI21_X1 U8172 ( .B1(n6633), .B2(n9653), .A(n6632), .ZN(P1_U3350) );
  AOI22_X1 U8173 ( .A1(n6634), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9647), .ZN(n6635) );
  OAI21_X1 U8174 ( .B1(n6636), .B2(n9653), .A(n6635), .ZN(P1_U3347) );
  INV_X1 U8175 ( .A(n6800), .ZN(n6828) );
  OAI222_X1 U8176 ( .A1(n8197), .A2(n6637), .B1(n8195), .B2(n6636), .C1(
        P2_U3152), .C2(n6828), .ZN(P2_U3352) );
  INV_X1 U8177 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6640) );
  INV_X1 U8178 ( .A(n6739), .ZN(n6638) );
  NAND2_X1 U8179 ( .A1(n6638), .A2(n6641), .ZN(n6639) );
  OAI21_X1 U8180 ( .B1(n6641), .B2(n6640), .A(n6639), .ZN(P1_U3440) );
  INV_X1 U8181 ( .A(n6642), .ZN(n6644) );
  AOI22_X1 U8182 ( .A1(n6691), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9647), .ZN(n6643) );
  OAI21_X1 U8183 ( .B1(n6644), .B2(n9653), .A(n6643), .ZN(P1_U3346) );
  INV_X1 U8184 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6645) );
  INV_X1 U8185 ( .A(n6845), .ZN(n6817) );
  OAI222_X1 U8186 ( .A1(n8197), .A2(n6645), .B1(n8195), .B2(n6644), .C1(
        P2_U3152), .C2(n6817), .ZN(P2_U3351) );
  INV_X1 U8187 ( .A(n6646), .ZN(n6648) );
  AOI22_X1 U8188 ( .A1(n9807), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9647), .ZN(n6647) );
  OAI21_X1 U8189 ( .B1(n6648), .B2(n9653), .A(n6647), .ZN(P1_U3345) );
  INV_X1 U8190 ( .A(n6906), .ZN(n6853) );
  OAI222_X1 U8191 ( .A1(n8197), .A2(n9501), .B1(n8195), .B2(n6648), .C1(
        P2_U3152), .C2(n6853), .ZN(P2_U3350) );
  INV_X1 U8192 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6659) );
  INV_X1 U8193 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6649) );
  NAND2_X1 U8194 ( .A1(n6650), .A2(n6649), .ZN(n6651) );
  NAND2_X1 U8195 ( .A1(n6894), .A2(n6651), .ZN(n6653) );
  INV_X1 U8196 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6880) );
  AOI21_X1 U8197 ( .B1(n6565), .B2(n6880), .A(n9655), .ZN(n6652) );
  NAND2_X1 U8198 ( .A1(n6653), .A2(n4396), .ZN(n9748) );
  OAI211_X1 U8199 ( .C1(n6653), .C2(n6652), .A(n9748), .B(P1_STATE_REG_SCAN_IN), .ZN(n6654) );
  INV_X1 U8200 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7237) );
  OAI22_X1 U8201 ( .A1(n6655), .A2(n6654), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7237), .ZN(n6656) );
  INV_X1 U8202 ( .A(n6656), .ZN(n6658) );
  NAND3_X1 U8203 ( .A1(n9823), .A2(n9655), .A3(n6880), .ZN(n6657) );
  OAI211_X1 U8204 ( .C1(n9773), .C2(n6659), .A(n6658), .B(n6657), .ZN(P1_U3241) );
  INV_X1 U8205 ( .A(n6660), .ZN(n6662) );
  AOI22_X1 U8206 ( .A1(n6980), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9647), .ZN(n6661) );
  OAI21_X1 U8207 ( .B1(n6662), .B2(n9653), .A(n6661), .ZN(P1_U3344) );
  INV_X1 U8208 ( .A(n7178), .ZN(n6914) );
  OAI222_X1 U8209 ( .A1(n8197), .A2(n6663), .B1(n8195), .B2(n6662), .C1(n6914), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8210 ( .A(n6664), .ZN(n6681) );
  AOI22_X1 U8211 ( .A1(n9826), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9647), .ZN(n6665) );
  OAI21_X1 U8212 ( .B1(n6681), .B2(n9653), .A(n6665), .ZN(P1_U3343) );
  INV_X1 U8213 ( .A(n6666), .ZN(n6683) );
  AOI22_X1 U8214 ( .A1(n6982), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9650), .ZN(n6667) );
  OAI21_X1 U8215 ( .B1(n6683), .B2(n9653), .A(n6667), .ZN(P1_U3342) );
  INV_X1 U8216 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6680) );
  AND2_X1 U8217 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7028) );
  MUX2_X1 U8218 ( .A(n6595), .B(P1_REG1_REG_3__SCAN_IN), .S(n6673), .Z(n6668)
         );
  NAND3_X1 U8219 ( .A1(n9759), .A2(n6669), .A3(n6668), .ZN(n6670) );
  AND3_X1 U8220 ( .A1(n9823), .A2(n6671), .A3(n6670), .ZN(n6672) );
  AOI211_X1 U8221 ( .C1(n9825), .C2(n6673), .A(n7028), .B(n6672), .ZN(n6679)
         );
  MUX2_X1 U8222 ( .A(n6580), .B(P1_REG2_REG_3__SCAN_IN), .S(n6673), .Z(n6675)
         );
  NAND3_X1 U8223 ( .A1(n6675), .A2(n9755), .A3(n6674), .ZN(n6676) );
  NAND3_X1 U8224 ( .A1(n9798), .A2(n6677), .A3(n6676), .ZN(n6678) );
  OAI211_X1 U8225 ( .C1(n6680), .C2(n9773), .A(n6679), .B(n6678), .ZN(P1_U3244) );
  INV_X1 U8226 ( .A(n7397), .ZN(n7186) );
  OAI222_X1 U8227 ( .A1(n8197), .A2(n6682), .B1(n8195), .B2(n6681), .C1(n7186), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8228 ( .A(n7562), .ZN(n7555) );
  OAI222_X1 U8229 ( .A1(n8197), .A2(n6684), .B1(n8195), .B2(n6683), .C1(n7555), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  AOI21_X1 U8230 ( .B1(n6687), .B2(n6686), .A(n6685), .ZN(n6697) );
  INV_X1 U8231 ( .A(n9823), .ZN(n9072) );
  AOI21_X1 U8232 ( .B1(n6690), .B2(n6689), .A(n6688), .ZN(n6694) );
  AND2_X1 U8233 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7251) );
  AOI21_X1 U8234 ( .B1(n9825), .B2(n6691), .A(n7251), .ZN(n6693) );
  INV_X1 U8235 ( .A(n9773), .ZN(n9827) );
  NAND2_X1 U8236 ( .A1(n9827), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n6692) );
  OAI211_X1 U8237 ( .C1(n6694), .C2(n9817), .A(n6693), .B(n6692), .ZN(n6695)
         );
  INV_X1 U8238 ( .A(n6695), .ZN(n6696) );
  OAI21_X1 U8239 ( .B1(n6697), .B2(n9072), .A(n6696), .ZN(P1_U3248) );
  INV_X1 U8240 ( .A(n6698), .ZN(n6701) );
  AOI22_X1 U8241 ( .A1(n8369), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n8889), .ZN(n6699) );
  OAI21_X1 U8242 ( .B1(n6701), .B2(n8195), .A(n6699), .ZN(P2_U3346) );
  AOI22_X1 U8243 ( .A1(n7166), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9650), .ZN(n6700) );
  OAI21_X1 U8244 ( .B1(n6701), .B2(n9653), .A(n6700), .ZN(P1_U3341) );
  AOI21_X1 U8245 ( .B1(n6704), .B2(n6703), .A(n6702), .ZN(n6713) );
  INV_X1 U8246 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6705) );
  NOR2_X1 U8247 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6705), .ZN(n9019) );
  NOR2_X1 U8248 ( .A1(n9060), .A2(n6706), .ZN(n6707) );
  AOI211_X1 U8249 ( .C1(n9827), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n9019), .B(
        n6707), .ZN(n6712) );
  OAI211_X1 U8250 ( .C1(n6710), .C2(n6709), .A(n9798), .B(n6708), .ZN(n6711)
         );
  OAI211_X1 U8251 ( .C1(n6713), .C2(n9072), .A(n6712), .B(n6711), .ZN(P1_U3247) );
  NAND2_X1 U8252 ( .A1(n9926), .A2(n6767), .ZN(n6714) );
  NAND2_X1 U8253 ( .A1(n6714), .A2(n5740), .ZN(n6716) );
  INV_X1 U8254 ( .A(n7001), .ZN(n6959) );
  OR2_X1 U8255 ( .A1(n9926), .A2(n6959), .ZN(n6715) );
  AND2_X1 U8256 ( .A1(n6716), .A2(n6715), .ZN(n8446) );
  NOR2_X1 U8257 ( .A1(n9920), .A2(P2_U3966), .ZN(P2_U3151) );
  NAND2_X1 U8258 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(P1_U3084), .ZN(n6722) );
  MUX2_X1 U8259 ( .A(n6592), .B(P1_REG1_REG_1__SCAN_IN), .S(n4300), .Z(n6717)
         );
  INV_X1 U8260 ( .A(n6717), .ZN(n6719) );
  OAI211_X1 U8261 ( .C1(n6720), .C2(n6719), .A(n9823), .B(n6718), .ZN(n6721)
         );
  OAI211_X1 U8262 ( .C1(n9060), .C2(n6723), .A(n6722), .B(n6721), .ZN(n6730)
         );
  INV_X1 U8263 ( .A(n6724), .ZN(n9747) );
  MUX2_X1 U8264 ( .A(n6576), .B(P1_REG2_REG_1__SCAN_IN), .S(n4300), .Z(n6728)
         );
  INV_X1 U8265 ( .A(n6726), .ZN(n6727) );
  AOI211_X1 U8266 ( .C1(n9747), .C2(n6728), .A(n6727), .B(n9817), .ZN(n6729)
         );
  AOI211_X1 U8267 ( .C1(P1_ADDR_REG_1__SCAN_IN), .C2(n9827), .A(n6730), .B(
        n6729), .ZN(n6731) );
  INV_X1 U8268 ( .A(n6731), .ZN(P1_U3242) );
  OR3_X1 U8269 ( .A1(n6733), .A2(n6732), .A3(n6737), .ZN(n6736) );
  NAND2_X1 U8270 ( .A1(n6326), .A2(n9349), .ZN(n6735) );
  NAND2_X1 U8271 ( .A1(n6736), .A2(n6735), .ZN(n7241) );
  AOI21_X1 U8272 ( .B1(n6885), .B2(n6737), .A(n7241), .ZN(n6882) );
  NOR2_X1 U8273 ( .A1(n6738), .A2(n9837), .ZN(n6740) );
  AND3_X1 U8274 ( .A1(n6740), .A2(n6739), .A3(n6758), .ZN(n7091) );
  AND2_X2 U8275 ( .A1(n6741), .A2(n7091), .ZN(n9897) );
  INV_X1 U8276 ( .A(n9897), .ZN(n9895) );
  INV_X1 U8277 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6742) );
  OR2_X1 U8278 ( .A1(n9897), .A2(n6742), .ZN(n6743) );
  OAI21_X1 U8279 ( .B1(n6882), .B2(n9895), .A(n6743), .ZN(P1_U3454) );
  INV_X1 U8280 ( .A(n6744), .ZN(n6750) );
  AOI22_X1 U8281 ( .A1(n7465), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9650), .ZN(n6745) );
  OAI21_X1 U8282 ( .B1(n6750), .B2(n9653), .A(n6745), .ZN(P1_U3340) );
  INV_X1 U8283 ( .A(n6746), .ZN(n6752) );
  AOI22_X1 U8284 ( .A1(n7686), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9647), .ZN(n6747) );
  OAI21_X1 U8285 ( .B1(n6752), .B2(n9653), .A(n6747), .ZN(P1_U3339) );
  INV_X1 U8286 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6749) );
  NAND2_X1 U8287 ( .A1(n8113), .A2(P1_U4006), .ZN(n6748) );
  OAI21_X1 U8288 ( .B1(P1_U4006), .B2(n6749), .A(n6748), .ZN(P1_U3586) );
  INV_X1 U8289 ( .A(n7734), .ZN(n7559) );
  OAI222_X1 U8290 ( .A1(n8197), .A2(n6751), .B1(n8195), .B2(n6750), .C1(n7559), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8291 ( .A(n7955), .ZN(n7731) );
  OAI222_X1 U8292 ( .A1(n8197), .A2(n6753), .B1(n8195), .B2(n6752), .C1(n7731), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8293 ( .A(n6754), .ZN(n6755) );
  AOI21_X1 U8294 ( .B1(n6757), .B2(n6756), .A(n6755), .ZN(n6761) );
  AOI22_X1 U8295 ( .A1(n9020), .A2(n6325), .B1(n9022), .B2(n9054), .ZN(n6760)
         );
  NAND2_X1 U8296 ( .A1(n9024), .A2(n6758), .ZN(n6871) );
  AOI22_X1 U8297 ( .A1(n9038), .A2(n7094), .B1(n6871), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6759) );
  OAI211_X1 U8298 ( .C1(n6761), .C2(n9012), .A(n6760), .B(n6759), .ZN(P1_U3220) );
  AOI22_X1 U8299 ( .A1(n9022), .A2(n6326), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n6871), .ZN(n6766) );
  OAI21_X1 U8300 ( .B1(n6764), .B2(n6763), .A(n6762), .ZN(n9746) );
  NAND2_X1 U8301 ( .A1(n9746), .A2(n5630), .ZN(n6765) );
  OAI211_X1 U8302 ( .C1(n7921), .C2(n7238), .A(n6766), .B(n6765), .ZN(P1_U3230) );
  OR2_X1 U8303 ( .A1(n9926), .A2(n7001), .ZN(n6768) );
  OAI211_X1 U8304 ( .C1(P2_U3152), .C2(n7061), .A(n6768), .B(n6767), .ZN(n6774) );
  NAND2_X1 U8305 ( .A1(n6774), .A2(n6769), .ZN(n6770) );
  NAND2_X1 U8306 ( .A1(n6770), .A2(n8353), .ZN(n6785) );
  NAND2_X1 U8307 ( .A1(n6785), .A2(n6310), .ZN(n9915) );
  NOR2_X1 U8308 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7153), .ZN(n6778) );
  INV_X1 U8309 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6965) );
  MUX2_X1 U8310 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6965), .S(n6782), .Z(n9659)
         );
  INV_X1 U8311 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9990) );
  XNOR2_X1 U8312 ( .A(n7047), .B(n9990), .ZN(n7042) );
  AND2_X1 U8313 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n7041) );
  NAND2_X1 U8314 ( .A1(n7042), .A2(n7041), .ZN(n7040) );
  NAND2_X1 U8315 ( .A1(n7047), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6771) );
  NAND2_X1 U8316 ( .A1(n7040), .A2(n6771), .ZN(n9658) );
  NAND2_X1 U8317 ( .A1(n6806), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6772) );
  OAI21_X1 U8318 ( .B1(n6806), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6772), .ZN(
        n6775) );
  AND2_X1 U8319 ( .A1(n6769), .A2(n6783), .ZN(n6773) );
  INV_X1 U8320 ( .A(n9914), .ZN(n7952) );
  AOI211_X1 U8321 ( .C1(n6776), .C2(n6775), .A(n6791), .B(n7952), .ZN(n6777)
         );
  AOI211_X1 U8322 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n9920), .A(n6778), .B(
        n6777), .ZN(n6789) );
  MUX2_X1 U8323 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6779), .S(n6806), .Z(n6787)
         );
  MUX2_X1 U8324 ( .A(n7048), .B(P2_REG2_REG_1__SCAN_IN), .S(n7047), .Z(n6780)
         );
  INV_X1 U8325 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9923) );
  OR3_X1 U8326 ( .A1(n6780), .A2(n7046), .A3(n9923), .ZN(n7049) );
  OAI21_X1 U8327 ( .B1(n7048), .B2(n6781), .A(n7049), .ZN(n9665) );
  MUX2_X1 U8328 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n7312), .S(n6782), .Z(n9664)
         );
  NAND2_X1 U8329 ( .A1(n9665), .A2(n9664), .ZN(n9663) );
  OAI21_X1 U8330 ( .B1(n7312), .B2(n9661), .A(n9663), .ZN(n6786) );
  NOR2_X1 U8331 ( .A1(n6310), .A2(n6783), .ZN(n6784) );
  NAND2_X1 U8332 ( .A1(n6785), .A2(n6784), .ZN(n9917) );
  NAND2_X1 U8333 ( .A1(n6787), .A2(n6786), .ZN(n6807) );
  OAI211_X1 U8334 ( .C1(n6787), .C2(n6786), .A(n9912), .B(n6807), .ZN(n6788)
         );
  OAI211_X1 U8335 ( .C1(n9915), .C2(n6790), .A(n6789), .B(n6788), .ZN(P2_U3248) );
  NOR2_X1 U8336 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7383), .ZN(n6799) );
  AOI21_X1 U8337 ( .B1(n6806), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6791), .ZN(
        n6832) );
  NAND2_X1 U8338 ( .A1(n6804), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6792) );
  OAI21_X1 U8339 ( .B1(n6804), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6792), .ZN(
        n6831) );
  NAND2_X1 U8340 ( .A1(n6802), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6793) );
  OAI21_X1 U8341 ( .B1(n6802), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6793), .ZN(
        n6855) );
  INV_X1 U8342 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6794) );
  MUX2_X1 U8343 ( .A(n6794), .B(P2_REG1_REG_6__SCAN_IN), .S(n6800), .Z(n6819)
         );
  NOR2_X1 U8344 ( .A1(n6820), .A2(n6819), .ZN(n6818) );
  AOI21_X1 U8345 ( .B1(n6800), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6818), .ZN(
        n6797) );
  INV_X1 U8346 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6795) );
  MUX2_X1 U8347 ( .A(n6795), .B(P2_REG1_REG_7__SCAN_IN), .S(n6845), .Z(n6796)
         );
  NOR2_X1 U8348 ( .A1(n6797), .A2(n6796), .ZN(n6840) );
  AOI211_X1 U8349 ( .C1(n6797), .C2(n6796), .A(n6840), .B(n7952), .ZN(n6798)
         );
  AOI211_X1 U8350 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n9920), .A(n6799), .B(
        n6798), .ZN(n6816) );
  NAND2_X1 U8351 ( .A1(n6800), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6811) );
  MUX2_X1 U8352 ( .A(n5753), .B(P2_REG2_REG_6__SCAN_IN), .S(n6800), .Z(n6801)
         );
  INV_X1 U8353 ( .A(n6801), .ZN(n6824) );
  NAND2_X1 U8354 ( .A1(n6802), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6810) );
  MUX2_X1 U8355 ( .A(n7422), .B(P2_REG2_REG_5__SCAN_IN), .S(n6802), .Z(n6803)
         );
  INV_X1 U8356 ( .A(n6803), .ZN(n6860) );
  NAND2_X1 U8357 ( .A1(n6804), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6809) );
  MUX2_X1 U8358 ( .A(n8743), .B(P2_REG2_REG_4__SCAN_IN), .S(n6804), .Z(n6805)
         );
  INV_X1 U8359 ( .A(n6805), .ZN(n6835) );
  NAND2_X1 U8360 ( .A1(n6806), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U8361 ( .A1(n6808), .A2(n6807), .ZN(n6836) );
  NAND2_X1 U8362 ( .A1(n6835), .A2(n6836), .ZN(n6834) );
  NAND2_X1 U8363 ( .A1(n6809), .A2(n6834), .ZN(n6861) );
  NAND2_X1 U8364 ( .A1(n6860), .A2(n6861), .ZN(n6859) );
  NAND2_X1 U8365 ( .A1(n6810), .A2(n6859), .ZN(n6825) );
  NAND2_X1 U8366 ( .A1(n6824), .A2(n6825), .ZN(n6823) );
  NAND2_X1 U8367 ( .A1(n6811), .A2(n6823), .ZN(n6814) );
  MUX2_X1 U8368 ( .A(n5767), .B(P2_REG2_REG_7__SCAN_IN), .S(n6845), .Z(n6812)
         );
  INV_X1 U8369 ( .A(n6812), .ZN(n6813) );
  NAND2_X1 U8370 ( .A1(n6813), .A2(n6814), .ZN(n6846) );
  OAI211_X1 U8371 ( .C1(n6814), .C2(n6813), .A(n9912), .B(n6846), .ZN(n6815)
         );
  OAI211_X1 U8372 ( .C1(n9915), .C2(n6817), .A(n6816), .B(n6815), .ZN(P2_U3252) );
  NAND2_X1 U8373 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7377) );
  INV_X1 U8374 ( .A(n7377), .ZN(n6822) );
  AOI211_X1 U8375 ( .C1(n6820), .C2(n6819), .A(n6818), .B(n7952), .ZN(n6821)
         );
  AOI211_X1 U8376 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n9920), .A(n6822), .B(
        n6821), .ZN(n6827) );
  OAI211_X1 U8377 ( .C1(n6825), .C2(n6824), .A(n9912), .B(n6823), .ZN(n6826)
         );
  OAI211_X1 U8378 ( .C1(n9915), .C2(n6828), .A(n6827), .B(n6826), .ZN(P2_U3251) );
  NOR2_X1 U8379 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6829), .ZN(n7065) );
  AOI211_X1 U8380 ( .C1(n6832), .C2(n6831), .A(n6830), .B(n7952), .ZN(n6833)
         );
  AOI211_X1 U8381 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n9920), .A(n7065), .B(
        n6833), .ZN(n6838) );
  OAI211_X1 U8382 ( .C1(n6836), .C2(n6835), .A(n9912), .B(n6834), .ZN(n6837)
         );
  OAI211_X1 U8383 ( .C1(n9915), .C2(n6839), .A(n6838), .B(n6837), .ZN(P2_U3249) );
  AND2_X1 U8384 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n8241) );
  AOI21_X1 U8385 ( .B1(n6845), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6840), .ZN(
        n6843) );
  INV_X1 U8386 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6841) );
  MUX2_X1 U8387 ( .A(n6841), .B(P2_REG1_REG_8__SCAN_IN), .S(n6906), .Z(n6842)
         );
  AOI211_X1 U8388 ( .C1(n6843), .C2(n6842), .A(n6901), .B(n7952), .ZN(n6844)
         );
  AOI211_X1 U8389 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n9920), .A(n8241), .B(
        n6844), .ZN(n6852) );
  NAND2_X1 U8390 ( .A1(n6845), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6847) );
  NAND2_X1 U8391 ( .A1(n6847), .A2(n6846), .ZN(n6850) );
  MUX2_X1 U8392 ( .A(n5783), .B(P2_REG2_REG_8__SCAN_IN), .S(n6906), .Z(n6848)
         );
  INV_X1 U8393 ( .A(n6848), .ZN(n6849) );
  NAND2_X1 U8394 ( .A1(n6849), .A2(n6850), .ZN(n6907) );
  OAI211_X1 U8395 ( .C1(n6850), .C2(n6849), .A(n9912), .B(n6907), .ZN(n6851)
         );
  OAI211_X1 U8396 ( .C1(n9915), .C2(n6853), .A(n6852), .B(n6851), .ZN(P2_U3253) );
  NOR2_X1 U8397 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5750), .ZN(n6858) );
  AOI211_X1 U8398 ( .C1(n6856), .C2(n6855), .A(n6854), .B(n7952), .ZN(n6857)
         );
  AOI211_X1 U8399 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n9920), .A(n6858), .B(
        n6857), .ZN(n6863) );
  OAI211_X1 U8400 ( .C1(n6861), .C2(n6860), .A(n9912), .B(n6859), .ZN(n6862)
         );
  OAI211_X1 U8401 ( .C1(n9915), .C2(n6864), .A(n6863), .B(n6862), .ZN(P2_U3250) );
  INV_X1 U8402 ( .A(n6865), .ZN(n6866) );
  NOR2_X1 U8403 ( .A1(n6867), .A2(n6866), .ZN(n6870) );
  INV_X1 U8404 ( .A(n6868), .ZN(n6869) );
  AOI21_X1 U8405 ( .B1(n6870), .B2(n6754), .A(n6869), .ZN(n6875) );
  AOI22_X1 U8406 ( .A1(n9020), .A2(n6326), .B1(n9022), .B2(n9053), .ZN(n6874)
         );
  AOI22_X1 U8407 ( .A1(n9038), .A2(n6872), .B1(n6871), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n6873) );
  OAI211_X1 U8408 ( .C1(n6875), .C2(n9012), .A(n6874), .B(n6873), .ZN(P1_U3235) );
  INV_X1 U8409 ( .A(n6876), .ZN(n6990) );
  AOI22_X1 U8410 ( .A1(n7690), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n9650), .ZN(n6877) );
  OAI21_X1 U8411 ( .B1(n6990), .B2(n9653), .A(n6877), .ZN(P1_U3338) );
  INV_X1 U8412 ( .A(n6878), .ZN(n6879) );
  AND2_X2 U8413 ( .A1(n9033), .A2(n6879), .ZN(n9911) );
  NAND2_X1 U8414 ( .A1(n9909), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6881) );
  OAI21_X1 U8415 ( .B1(n6882), .B2(n9909), .A(n6881), .ZN(P1_U3523) );
  NAND2_X1 U8416 ( .A1(n6326), .A2(n7094), .ZN(n6883) );
  NAND2_X1 U8417 ( .A1(n6884), .A2(n6889), .ZN(n7118) );
  OAI21_X1 U8418 ( .B1(n6884), .B2(n6889), .A(n7118), .ZN(n7216) );
  NOR2_X1 U8419 ( .A1(n6921), .A2(n7214), .ZN(n6886) );
  OR2_X1 U8420 ( .A1(n7265), .A2(n6886), .ZN(n7210) );
  INV_X1 U8421 ( .A(n7093), .ZN(n7453) );
  OR2_X1 U8422 ( .A1(n7198), .A2(n7453), .ZN(n9854) );
  OAI22_X1 U8423 ( .A1(n7210), .A2(n9854), .B1(n7214), .B2(n9852), .ZN(n6899)
         );
  NAND2_X1 U8424 ( .A1(n9110), .A2(n7538), .ZN(n6888) );
  NAND2_X1 U8425 ( .A1(n7472), .A2(n7453), .ZN(n6887) );
  AND2_X1 U8426 ( .A1(n6888), .A2(n6887), .ZN(n9716) );
  XNOR2_X1 U8427 ( .A(n6531), .B(n6889), .ZN(n6898) );
  NAND2_X1 U8428 ( .A1(n6891), .A2(n6890), .ZN(n6892) );
  OAI21_X1 U8429 ( .B1(n6893), .B2(n5628), .A(n6892), .ZN(n9719) );
  NAND2_X1 U8430 ( .A1(n7216), .A2(n9719), .ZN(n6897) );
  AOI22_X1 U8431 ( .A1(n9053), .A2(n9349), .B1(n9347), .B2(n6326), .ZN(n6896)
         );
  OAI211_X1 U8432 ( .C1(n9716), .C2(n6898), .A(n6897), .B(n6896), .ZN(n7208)
         );
  AOI211_X1 U8433 ( .C1(n9884), .C2(n7216), .A(n6899), .B(n7208), .ZN(n7054)
         );
  NAND2_X1 U8434 ( .A1(n9909), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6900) );
  OAI21_X1 U8435 ( .B1(n7054), .B2(n9909), .A(n6900), .ZN(P1_U3525) );
  NOR2_X1 U8436 ( .A1(n9586), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7594) );
  INV_X1 U8437 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6902) );
  MUX2_X1 U8438 ( .A(n6902), .B(P2_REG1_REG_9__SCAN_IN), .S(n7178), .Z(n6903)
         );
  AOI211_X1 U8439 ( .C1(n6904), .C2(n6903), .A(n7173), .B(n7952), .ZN(n6905)
         );
  AOI211_X1 U8440 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n9920), .A(n7594), .B(
        n6905), .ZN(n6913) );
  NAND2_X1 U8441 ( .A1(n6906), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6908) );
  NAND2_X1 U8442 ( .A1(n6908), .A2(n6907), .ZN(n6911) );
  MUX2_X1 U8443 ( .A(n5802), .B(P2_REG2_REG_9__SCAN_IN), .S(n7178), .Z(n6909)
         );
  INV_X1 U8444 ( .A(n6909), .ZN(n6910) );
  NAND2_X1 U8445 ( .A1(n6910), .A2(n6911), .ZN(n7179) );
  OAI211_X1 U8446 ( .C1(n6911), .C2(n6910), .A(n9912), .B(n7179), .ZN(n6912)
         );
  OAI211_X1 U8447 ( .C1(n9915), .C2(n6914), .A(n6913), .B(n6912), .ZN(P2_U3254) );
  INV_X1 U8448 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6925) );
  OR2_X1 U8449 ( .A1(n9719), .A2(n9884), .ZN(n9873) );
  INV_X1 U8450 ( .A(n9716), .ZN(n9352) );
  XNOR2_X1 U8451 ( .A(n6918), .B(n6917), .ZN(n6919) );
  AOI222_X1 U8452 ( .A1(n9352), .A2(n6919), .B1(n9054), .B2(n9349), .C1(n6325), 
        .C2(n9347), .ZN(n7096) );
  INV_X1 U8453 ( .A(n9854), .ZN(n9888) );
  OAI21_X1 U8454 ( .B1(n6920), .B2(n7238), .A(n9888), .ZN(n6922) );
  NOR2_X1 U8455 ( .A1(n6922), .A2(n6921), .ZN(n7100) );
  AOI21_X1 U8456 ( .B1(n9887), .B2(n7094), .A(n7100), .ZN(n6923) );
  OAI211_X1 U8457 ( .C1(n9892), .C2(n7097), .A(n7096), .B(n6923), .ZN(n7111)
         );
  NAND2_X1 U8458 ( .A1(n7111), .A2(n9897), .ZN(n6924) );
  OAI21_X1 U8459 ( .B1(n9897), .B2(n6925), .A(n6924), .ZN(P1_U3457) );
  INV_X1 U8460 ( .A(n6926), .ZN(n6929) );
  AOI22_X1 U8461 ( .A1(n9078), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9650), .ZN(n6927) );
  OAI21_X1 U8462 ( .B1(n6929), .B2(n9653), .A(n6927), .ZN(P1_U3337) );
  AOI22_X1 U8463 ( .A1(n8407), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8889), .ZN(n6928) );
  OAI21_X1 U8464 ( .B1(n6929), .B2(n8195), .A(n6928), .ZN(P2_U3342) );
  NOR4_X1 U8465 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6933) );
  NOR4_X1 U8466 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6932) );
  NOR4_X1 U8467 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6931) );
  NOR4_X1 U8468 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6930) );
  NAND4_X1 U8469 ( .A1(n6933), .A2(n6932), .A3(n6931), .A4(n6930), .ZN(n6941)
         );
  NOR2_X1 U8470 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .ZN(
        n6937) );
  NOR4_X1 U8471 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n6936) );
  NOR4_X1 U8472 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6935) );
  NOR4_X1 U8473 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6934) );
  NAND4_X1 U8474 ( .A1(n6937), .A2(n6936), .A3(n6935), .A4(n6934), .ZN(n6940)
         );
  XNOR2_X1 U8475 ( .A(n7813), .B(P2_B_REG_SCAN_IN), .ZN(n6938) );
  OAI21_X1 U8476 ( .B1(n6941), .B2(n6940), .A(n9925), .ZN(n6992) );
  AND2_X1 U8477 ( .A1(n7001), .A2(n6997), .ZN(n7059) );
  NOR2_X1 U8478 ( .A1(n9926), .A2(n7059), .ZN(n6995) );
  NAND2_X1 U8479 ( .A1(n6992), .A2(n6995), .ZN(n7293) );
  NOR2_X1 U8480 ( .A1(n8854), .A2(n7007), .ZN(n6994) );
  NOR2_X1 U8481 ( .A1(n7293), .A2(n6994), .ZN(n6943) );
  INV_X1 U8482 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9935) );
  AND2_X1 U8483 ( .A1(n7945), .A2(n7950), .ZN(n9936) );
  AOI21_X1 U8484 ( .B1(n9925), .B2(n9935), .A(n9936), .ZN(n7294) );
  INV_X1 U8485 ( .A(n7294), .ZN(n6942) );
  AND2_X1 U8486 ( .A1(n7813), .A2(n7950), .ZN(n9933) );
  INV_X1 U8487 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9932) );
  AND2_X1 U8488 ( .A1(n9925), .A2(n9932), .ZN(n6944) );
  AND2_X2 U8489 ( .A1(n6967), .A2(n7292), .ZN(n10001) );
  NAND2_X1 U8490 ( .A1(n6945), .A2(n9938), .ZN(n7357) );
  NAND2_X1 U8491 ( .A1(n6946), .A2(n7357), .ZN(n7356) );
  NAND2_X1 U8492 ( .A1(n7356), .A2(n8050), .ZN(n6949) );
  INV_X1 U8493 ( .A(n7357), .ZN(n7011) );
  CLKBUF_X1 U8494 ( .A(n6947), .Z(n8364) );
  NAND2_X1 U8495 ( .A1(n7011), .A2(n8364), .ZN(n6948) );
  MUX2_X1 U8496 ( .A(n6950), .B(n6959), .S(n7455), .Z(n6952) );
  AND2_X1 U8497 ( .A1(n7303), .A2(n8440), .ZN(n6951) );
  NAND2_X1 U8498 ( .A1(n6952), .A2(n6951), .ZN(n7719) );
  NAND2_X1 U8499 ( .A1(n7719), .A2(n8854), .ZN(n9985) );
  OAI21_X1 U8500 ( .B1(n6953), .B2(n7409), .A(n6954), .ZN(n6960) );
  INV_X1 U8501 ( .A(n8630), .ZN(n8726) );
  OAI22_X1 U8502 ( .A1(n6957), .A2(n8726), .B1(n6958), .B2(n8728), .ZN(n6999)
         );
  AOI21_X1 U8503 ( .B1(n6960), .B2(n8740), .A(n6999), .ZN(n7313) );
  INV_X1 U8504 ( .A(n7303), .ZN(n9939) );
  NAND2_X1 U8505 ( .A1(n7350), .A2(n7407), .ZN(n7436) );
  OAI211_X1 U8506 ( .C1(n7350), .C2(n7407), .A(n8857), .B(n7436), .ZN(n7309)
         );
  INV_X1 U8507 ( .A(n7309), .ZN(n6962) );
  AOI21_X1 U8508 ( .B1(n8856), .B2(n7311), .A(n6962), .ZN(n6963) );
  OAI211_X1 U8509 ( .C1(n7316), .C2(n8861), .A(n7313), .B(n6963), .ZN(n6968)
         );
  NAND2_X1 U8510 ( .A1(n10001), .A2(n6968), .ZN(n6964) );
  OAI21_X1 U8511 ( .B1(n10001), .B2(n6965), .A(n6964), .ZN(P2_U3522) );
  INV_X1 U8512 ( .A(n7292), .ZN(n6966) );
  AND2_X2 U8513 ( .A1(n6967), .A2(n6966), .ZN(n9988) );
  INV_X1 U8514 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6970) );
  NAND2_X1 U8515 ( .A1(n9988), .A2(n6968), .ZN(n6969) );
  OAI21_X1 U8516 ( .B1(n9988), .B2(n6970), .A(n6969), .ZN(P2_U3457) );
  INV_X1 U8517 ( .A(n6982), .ZN(n9059) );
  INV_X1 U8518 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9741) );
  AOI22_X1 U8519 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n6982), .B1(n9059), .B2(
        n9741), .ZN(n9065) );
  INV_X1 U8520 ( .A(n9826), .ZN(n6971) );
  INV_X1 U8521 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9678) );
  AOI22_X1 U8522 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n9826), .B1(n6971), .B2(
        n9678), .ZN(n9815) );
  OAI21_X1 U8523 ( .B1(n6980), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6972), .ZN(
        n9814) );
  NAND2_X1 U8524 ( .A1(n9815), .A2(n9814), .ZN(n9813) );
  OAI21_X1 U8525 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n9826), .A(n9813), .ZN(
        n9064) );
  NAND2_X1 U8526 ( .A1(n9065), .A2(n9064), .ZN(n9063) );
  OAI21_X1 U8527 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6982), .A(n9063), .ZN(
        n6975) );
  INV_X1 U8528 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6973) );
  MUX2_X1 U8529 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6973), .S(n7166), .Z(n6974)
         );
  NAND2_X1 U8530 ( .A1(n6974), .A2(n6975), .ZN(n7159) );
  OAI21_X1 U8531 ( .B1(n6975), .B2(n6974), .A(n7159), .ZN(n6988) );
  INV_X1 U8532 ( .A(n7166), .ZN(n6977) );
  NAND2_X1 U8533 ( .A1(n9827), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6976) );
  NAND2_X1 U8534 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n7778) );
  OAI211_X1 U8535 ( .C1(n9060), .C2(n6977), .A(n6976), .B(n7778), .ZN(n6987)
         );
  INV_X1 U8536 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6978) );
  AOI22_X1 U8537 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6982), .B1(n9059), .B2(
        n6978), .ZN(n9057) );
  AOI21_X1 U8538 ( .B1(n6980), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6979), .ZN(
        n9820) );
  NAND2_X1 U8539 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n9826), .ZN(n6981) );
  OAI21_X1 U8540 ( .B1(n9826), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6981), .ZN(
        n9819) );
  INV_X1 U8541 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6983) );
  MUX2_X1 U8542 ( .A(n6983), .B(P1_REG2_REG_12__SCAN_IN), .S(n7166), .Z(n6984)
         );
  NOR2_X1 U8543 ( .A1(n6984), .A2(n6985), .ZN(n7165) );
  AOI211_X1 U8544 ( .C1(n6985), .C2(n6984), .A(n7165), .B(n9817), .ZN(n6986)
         );
  AOI211_X1 U8545 ( .C1(n9823), .C2(n6988), .A(n6987), .B(n6986), .ZN(n6989)
         );
  INV_X1 U8546 ( .A(n6989), .ZN(P1_U3253) );
  INV_X1 U8547 ( .A(n8390), .ZN(n8379) );
  OAI222_X1 U8548 ( .A1(n8197), .A2(n6991), .B1(n8195), .B2(n6990), .C1(
        P2_U3152), .C2(n8379), .ZN(P2_U3343) );
  AND2_X1 U8549 ( .A1(n6992), .A2(n7292), .ZN(n6993) );
  NAND2_X1 U8550 ( .A1(n7294), .A2(n6993), .ZN(n6996) );
  INV_X1 U8551 ( .A(n6994), .ZN(n7296) );
  NAND2_X1 U8552 ( .A1(n6996), .A2(n7296), .ZN(n7063) );
  AND2_X1 U8553 ( .A1(n7063), .A2(n6995), .ZN(n7039) );
  INV_X1 U8554 ( .A(n7039), .ZN(n8055) );
  INV_X1 U8555 ( .A(n6996), .ZN(n7004) );
  NOR2_X1 U8556 ( .A1(n9926), .A2(n6997), .ZN(n6998) );
  AOI22_X1 U8557 ( .A1(n8055), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n8282), .B2(
        n6999), .ZN(n7020) );
  NOR2_X1 U8558 ( .A1(n9926), .A2(n9980), .ZN(n7000) );
  NAND2_X1 U8559 ( .A1(n7063), .A2(n7000), .ZN(n8336) );
  OR2_X1 U8560 ( .A1(n8856), .A2(n7001), .ZN(n7002) );
  NOR2_X1 U8561 ( .A1(n9926), .A2(n7002), .ZN(n7003) );
  INV_X1 U8562 ( .A(n7005), .ZN(n7006) );
  NAND2_X1 U8563 ( .A1(n7006), .A2(n7493), .ZN(n7008) );
  NAND2_X1 U8564 ( .A1(n7455), .A2(n7007), .ZN(n7298) );
  NAND2_X4 U8565 ( .A1(n7008), .A2(n7298), .ZN(n8175) );
  XNOR2_X1 U8566 ( .A(n7407), .B(n8175), .ZN(n7067) );
  INV_X2 U8567 ( .A(n8174), .ZN(n8154) );
  NAND2_X1 U8568 ( .A1(n7009), .A2(n8154), .ZN(n7066) );
  XNOR2_X1 U8569 ( .A(n7067), .B(n7066), .ZN(n7071) );
  NOR2_X1 U8570 ( .A1(n8175), .A2(n9938), .ZN(n7010) );
  AOI21_X1 U8571 ( .B1(n7011), .B2(n6108), .A(n7010), .ZN(n8052) );
  XNOR2_X1 U8572 ( .A(n9945), .B(n8175), .ZN(n7013) );
  NAND2_X1 U8573 ( .A1(n8364), .A2(n6108), .ZN(n7012) );
  NAND2_X1 U8574 ( .A1(n7013), .A2(n7012), .ZN(n7017) );
  INV_X1 U8575 ( .A(n7012), .ZN(n7015) );
  INV_X1 U8576 ( .A(n7013), .ZN(n7014) );
  NAND2_X1 U8577 ( .A1(n7015), .A2(n7014), .ZN(n7016) );
  NAND2_X1 U8578 ( .A1(n8052), .A2(n8053), .ZN(n8051) );
  NAND2_X1 U8579 ( .A1(n8051), .A2(n7017), .ZN(n7072) );
  XOR2_X1 U8580 ( .A(n7071), .B(n7072), .Z(n7018) );
  AOI22_X1 U8581 ( .A1(n8346), .A2(n7311), .B1(n8325), .B2(n7018), .ZN(n7019)
         );
  NAND2_X1 U8582 ( .A1(n7020), .A2(n7019), .ZN(P2_U3239) );
  INV_X1 U8583 ( .A(n7023), .ZN(n7022) );
  NOR2_X1 U8584 ( .A1(n7021), .A2(n7022), .ZN(n7026) );
  NAND2_X1 U8585 ( .A1(n6868), .A2(n7023), .ZN(n7024) );
  NAND2_X1 U8586 ( .A1(n7024), .A2(n7021), .ZN(n8973) );
  INV_X1 U8587 ( .A(n8973), .ZN(n7025) );
  AOI21_X1 U8588 ( .B1(n7026), .B2(n6868), .A(n7025), .ZN(n7032) );
  INV_X1 U8589 ( .A(n9024), .ZN(n7254) );
  NAND2_X1 U8590 ( .A1(n7267), .A2(n9887), .ZN(n9839) );
  NOR2_X1 U8591 ( .A1(n7254), .A2(n9839), .ZN(n7027) );
  AOI211_X1 U8592 ( .C1(n9020), .C2(n9054), .A(n7028), .B(n7027), .ZN(n7031)
         );
  AOI22_X1 U8593 ( .A1(n9022), .A2(n9052), .B1(n9033), .B2(n7029), .ZN(n7030)
         );
  OAI211_X1 U8594 ( .C1(n7032), .C2(n9012), .A(n7031), .B(n7030), .ZN(P1_U3216) );
  INV_X1 U8595 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7300) );
  AOI22_X1 U8596 ( .A1(n8345), .A2(n8364), .B1(n8346), .B2(n9938), .ZN(n7038)
         );
  INV_X1 U8597 ( .A(n7346), .ZN(n7036) );
  INV_X1 U8598 ( .A(n7033), .ZN(n7034) );
  MUX2_X1 U8599 ( .A(n7034), .B(n9938), .S(n8174), .Z(n7035) );
  OAI21_X1 U8600 ( .B1(n7036), .B2(n7035), .A(n8325), .ZN(n7037) );
  OAI211_X1 U8601 ( .C1(n7039), .C2(n7300), .A(n7038), .B(n7037), .ZN(P2_U3234) );
  INV_X1 U8602 ( .A(n9915), .ZN(n8388) );
  INV_X1 U8603 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7353) );
  OAI211_X1 U8604 ( .C1(n7042), .C2(n7041), .A(n9914), .B(n7040), .ZN(n7044)
         );
  NAND2_X1 U8605 ( .A1(n9920), .A2(P2_ADDR_REG_1__SCAN_IN), .ZN(n7043) );
  OAI211_X1 U8606 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7353), .A(n7044), .B(n7043), .ZN(n7045) );
  AOI21_X1 U8607 ( .B1(n7047), .B2(n8388), .A(n7045), .ZN(n7053) );
  NOR2_X1 U8608 ( .A1(n9923), .A2(n7046), .ZN(n7051) );
  MUX2_X1 U8609 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n7048), .S(n7047), .Z(n7050)
         );
  OAI211_X1 U8610 ( .C1(n7051), .C2(n7050), .A(n9912), .B(n7049), .ZN(n7052)
         );
  NAND2_X1 U8611 ( .A1(n7053), .A2(n7052), .ZN(P2_U3246) );
  INV_X1 U8612 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7056) );
  OR2_X1 U8613 ( .A1(n7054), .A2(n9895), .ZN(n7055) );
  OAI21_X1 U8614 ( .B1(n9897), .B2(n7056), .A(n7055), .ZN(P1_U3460) );
  INV_X1 U8615 ( .A(n7057), .ZN(n7058) );
  NOR2_X1 U8616 ( .A1(n7059), .A2(n7058), .ZN(n7060) );
  AND2_X1 U8617 ( .A1(n7061), .A2(n7060), .ZN(n7062) );
  AOI21_X2 U8618 ( .B1(n7063), .B2(n7062), .A(P2_U3152), .ZN(n8333) );
  INV_X1 U8619 ( .A(n8747), .ZN(n7088) );
  OAI22_X1 U8620 ( .A1(n6958), .A2(n8726), .B1(n7498), .B2(n8728), .ZN(n8739)
         );
  NOR2_X1 U8621 ( .A1(n8336), .A2(n9952), .ZN(n7064) );
  AOI211_X1 U8622 ( .C1(n8282), .C2(n8739), .A(n7065), .B(n7064), .ZN(n7087)
         );
  INV_X1 U8623 ( .A(n7066), .ZN(n7069) );
  INV_X1 U8624 ( .A(n7067), .ZN(n7068) );
  NAND2_X1 U8625 ( .A1(n7069), .A2(n7068), .ZN(n7070) );
  XNOR2_X1 U8626 ( .A(n8175), .B(n7445), .ZN(n7073) );
  NAND2_X1 U8627 ( .A1(n8363), .A2(n8154), .ZN(n7074) );
  XNOR2_X1 U8628 ( .A(n7073), .B(n7074), .ZN(n7150) );
  INV_X1 U8629 ( .A(n7073), .ZN(n7075) );
  NOR2_X1 U8630 ( .A1(n7075), .A2(n7074), .ZN(n7076) );
  XNOR2_X1 U8631 ( .A(n8168), .B(n9952), .ZN(n7081) );
  INV_X1 U8632 ( .A(n7081), .ZN(n7079) );
  AND2_X1 U8633 ( .A1(n7077), .A2(n6108), .ZN(n7080) );
  INV_X1 U8634 ( .A(n7080), .ZN(n7078) );
  NAND2_X1 U8635 ( .A1(n7079), .A2(n7078), .ZN(n7105) );
  NAND2_X1 U8636 ( .A1(n7081), .A2(n7080), .ZN(n7082) );
  AND2_X1 U8637 ( .A1(n7105), .A2(n7082), .ZN(n7083) );
  NAND2_X1 U8638 ( .A1(n7084), .A2(n7083), .ZN(n7106) );
  OAI21_X1 U8639 ( .B1(n7084), .B2(n7083), .A(n7106), .ZN(n7085) );
  NAND2_X1 U8640 ( .A1(n7085), .A2(n8325), .ZN(n7086) );
  OAI211_X1 U8641 ( .C1(n8341), .C2(n7088), .A(n7087), .B(n7086), .ZN(P2_U3232) );
  INV_X1 U8642 ( .A(n7089), .ZN(n7090) );
  NAND2_X1 U8643 ( .A1(n7091), .A2(n7090), .ZN(n7130) );
  AND2_X1 U8644 ( .A1(n9110), .A2(n7092), .ZN(n7196) );
  NOR2_X1 U8645 ( .A1(n9719), .A2(n7196), .ZN(n7128) );
  INV_X1 U8646 ( .A(n9685), .ZN(n9720) );
  NOR2_X1 U8647 ( .A1(n7198), .A2(n7093), .ZN(n7131) );
  AOI22_X1 U8648 ( .A1(n9720), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n7131), .B2(
        n7094), .ZN(n7095) );
  OAI211_X1 U8649 ( .C1(n7128), .C2(n7097), .A(n7096), .B(n7095), .ZN(n7098)
         );
  NAND2_X1 U8650 ( .A1(n7098), .A2(n9725), .ZN(n7102) );
  AND2_X1 U8651 ( .A1(n9725), .A2(n7099), .ZN(n9306) );
  NAND2_X1 U8652 ( .A1(n9306), .A2(n7100), .ZN(n7101) );
  OAI211_X1 U8653 ( .C1(n6576), .C2(n9725), .A(n7102), .B(n7101), .ZN(P1_U3290) );
  INV_X1 U8654 ( .A(n7103), .ZN(n7157) );
  AOI22_X1 U8655 ( .A1(n9093), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9650), .ZN(n7104) );
  OAI21_X1 U8656 ( .B1(n7157), .B2(n9653), .A(n7104), .ZN(P1_U3336) );
  NAND2_X1 U8657 ( .A1(n7106), .A2(n7105), .ZN(n7365) );
  XNOR2_X1 U8658 ( .A(n9960), .B(n8175), .ZN(n7368) );
  NAND2_X1 U8659 ( .A1(n8362), .A2(n8154), .ZN(n7367) );
  XNOR2_X1 U8660 ( .A(n7368), .B(n7367), .ZN(n7366) );
  XNOR2_X1 U8661 ( .A(n7365), .B(n7366), .ZN(n7110) );
  INV_X1 U8662 ( .A(n7077), .ZN(n7431) );
  OAI22_X1 U8663 ( .A1(n7431), .A2(n8726), .B1(n7384), .B2(n8728), .ZN(n7420)
         );
  AOI22_X1 U8664 ( .A1(n8282), .A2(n7420), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n7107) );
  OAI21_X1 U8665 ( .B1(n9960), .B2(n8336), .A(n7107), .ZN(n7108) );
  AOI21_X1 U8666 ( .B1(n7414), .B2(n8333), .A(n7108), .ZN(n7109) );
  OAI21_X1 U8667 ( .B1(n7110), .B2(n8349), .A(n7109), .ZN(P2_U3229) );
  NAND2_X1 U8668 ( .A1(n7111), .A2(n9911), .ZN(n7112) );
  OAI21_X1 U8669 ( .B1(n9911), .B2(n6592), .A(n7112), .ZN(P1_U3524) );
  NAND2_X1 U8670 ( .A1(n7113), .A2(n9847), .ZN(n7276) );
  NAND2_X1 U8671 ( .A1(n9051), .A2(n7286), .ZN(n7121) );
  NAND2_X1 U8672 ( .A1(n7322), .A2(n7230), .ZN(n7124) );
  NAND2_X1 U8673 ( .A1(n7116), .A2(n7214), .ZN(n7117) );
  NAND2_X1 U8674 ( .A1(n7118), .A2(n7117), .ZN(n7262) );
  NAND2_X1 U8675 ( .A1(n7262), .A2(n7261), .ZN(n7260) );
  NAND2_X1 U8676 ( .A1(n4993), .A2(n7264), .ZN(n7119) );
  NAND2_X1 U8677 ( .A1(n7260), .A2(n7119), .ZN(n7188) );
  NAND2_X1 U8678 ( .A1(n7120), .A2(n7135), .ZN(n7189) );
  AND2_X1 U8679 ( .A1(n7189), .A2(n7121), .ZN(n7122) );
  NAND2_X1 U8680 ( .A1(n7188), .A2(n7122), .ZN(n7224) );
  NAND2_X1 U8681 ( .A1(n7127), .A2(n7141), .ZN(n7330) );
  OAI21_X1 U8682 ( .B1(n7127), .B2(n7141), .A(n7330), .ZN(n9874) );
  INV_X1 U8683 ( .A(n9874), .ZN(n7149) );
  INV_X1 U8684 ( .A(n7128), .ZN(n7129) );
  NAND2_X1 U8685 ( .A1(n9725), .A2(n7129), .ZN(n9356) );
  NAND2_X1 U8686 ( .A1(n7265), .A2(n7264), .ZN(n7263) );
  NOR2_X2 U8687 ( .A1(n7280), .A2(n7286), .ZN(n7228) );
  OAI211_X1 U8688 ( .C1(n7229), .C2(n7328), .A(n9888), .B(n7339), .ZN(n9869)
         );
  INV_X1 U8689 ( .A(n9869), .ZN(n7134) );
  NOR2_X1 U8690 ( .A1(n7130), .A2(n9110), .ZN(n7982) );
  INV_X1 U8691 ( .A(n7132), .ZN(n7249) );
  OAI22_X1 U8692 ( .A1(n9723), .A2(n7328), .B1(n9685), .B2(n7249), .ZN(n7133)
         );
  AOI21_X1 U8693 ( .B1(n7134), .B2(n7982), .A(n7133), .ZN(n7148) );
  AND2_X1 U8694 ( .A1(n7136), .A2(n7135), .ZN(n7137) );
  NAND2_X1 U8695 ( .A1(n7187), .A2(n7137), .ZN(n7142) );
  NAND2_X1 U8696 ( .A1(n7142), .A2(n7140), .ZN(n7139) );
  INV_X1 U8697 ( .A(n7141), .ZN(n7138) );
  NAND3_X1 U8698 ( .A1(n7142), .A2(n7141), .A3(n7140), .ZN(n7143) );
  NAND2_X1 U8699 ( .A1(n7333), .A2(n7143), .ZN(n7145) );
  INV_X1 U8700 ( .A(n9347), .ZN(n9712) );
  OAI22_X1 U8701 ( .A1(n7322), .A2(n9712), .B1(n8076), .B2(n9710), .ZN(n7144)
         );
  AOI21_X1 U8702 ( .B1(n7145), .B2(n9352), .A(n7144), .ZN(n9871) );
  MUX2_X1 U8703 ( .A(n7146), .B(n9871), .S(n9725), .Z(n7147) );
  OAI211_X1 U8704 ( .C1(n7149), .C2(n9356), .A(n7148), .B(n7147), .ZN(P1_U3284) );
  XNOR2_X1 U8705 ( .A(n7151), .B(n7150), .ZN(n7156) );
  OAI22_X1 U8706 ( .A1(n8314), .A2(n7431), .B1(n7410), .B2(n8336), .ZN(n7152)
         );
  AOI21_X1 U8707 ( .B1(n8240), .B2(n7009), .A(n7152), .ZN(n7155) );
  MUX2_X1 U8708 ( .A(P2_STATE_REG_SCAN_IN), .B(n8341), .S(n7153), .Z(n7154) );
  OAI211_X1 U8709 ( .C1(n8349), .C2(n7156), .A(n7155), .B(n7154), .ZN(P2_U3220) );
  INV_X1 U8710 ( .A(n8419), .ZN(n8405) );
  OAI222_X1 U8711 ( .A1(n8197), .A2(n9602), .B1(n8195), .B2(n7157), .C1(n8405), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8712 ( .A(n7465), .ZN(n7164) );
  NAND2_X1 U8713 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7915) );
  INV_X1 U8714 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7158) );
  MUX2_X1 U8715 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7158), .S(n7465), .Z(n7161)
         );
  OAI21_X1 U8716 ( .B1(n7166), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7159), .ZN(
        n7160) );
  NAND2_X1 U8717 ( .A1(n7161), .A2(n7160), .ZN(n7459) );
  OAI21_X1 U8718 ( .B1(n7161), .B2(n7160), .A(n7459), .ZN(n7162) );
  NAND2_X1 U8719 ( .A1(n9823), .A2(n7162), .ZN(n7163) );
  OAI211_X1 U8720 ( .C1(n9060), .C2(n7164), .A(n7915), .B(n7163), .ZN(n7171)
         );
  AOI21_X1 U8721 ( .B1(n7166), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7165), .ZN(
        n7169) );
  NAND2_X1 U8722 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7465), .ZN(n7167) );
  OAI21_X1 U8723 ( .B1(n7465), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7167), .ZN(
        n7168) );
  NOR2_X1 U8724 ( .A1(n7169), .A2(n7168), .ZN(n7464) );
  AOI211_X1 U8725 ( .C1(n7169), .C2(n7168), .A(n7464), .B(n9817), .ZN(n7170)
         );
  AOI211_X1 U8726 ( .C1(P1_ADDR_REG_13__SCAN_IN), .C2(n9827), .A(n7171), .B(
        n7170), .ZN(n7172) );
  INV_X1 U8727 ( .A(n7172), .ZN(P1_U3254) );
  AND2_X1 U8728 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n8219) );
  INV_X1 U8729 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7174) );
  MUX2_X1 U8730 ( .A(n7174), .B(P2_REG1_REG_10__SCAN_IN), .S(n7397), .Z(n7175)
         );
  NOR2_X1 U8731 ( .A1(n7176), .A2(n7175), .ZN(n7396) );
  AOI211_X1 U8732 ( .C1(n7176), .C2(n7175), .A(n7396), .B(n7952), .ZN(n7177)
         );
  AOI211_X1 U8733 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n9920), .A(n8219), .B(
        n7177), .ZN(n7185) );
  NAND2_X1 U8734 ( .A1(n7178), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7180) );
  NAND2_X1 U8735 ( .A1(n7180), .A2(n7179), .ZN(n7183) );
  MUX2_X1 U8736 ( .A(n5811), .B(P2_REG2_REG_10__SCAN_IN), .S(n7397), .Z(n7181)
         );
  INV_X1 U8737 ( .A(n7181), .ZN(n7182) );
  NAND2_X1 U8738 ( .A1(n7182), .A2(n7183), .ZN(n7389) );
  OAI211_X1 U8739 ( .C1(n7183), .C2(n7182), .A(n9912), .B(n7389), .ZN(n7184)
         );
  OAI211_X1 U8740 ( .C1(n9915), .C2(n7186), .A(n7185), .B(n7184), .ZN(P2_U3255) );
  XNOR2_X1 U8741 ( .A(n7187), .B(n7189), .ZN(n7194) );
  NAND2_X1 U8742 ( .A1(n7188), .A2(n7189), .ZN(n7277) );
  OR2_X1 U8743 ( .A1(n7188), .A2(n7189), .ZN(n7190) );
  NAND2_X1 U8744 ( .A1(n7277), .A2(n7190), .ZN(n9850) );
  NAND2_X1 U8745 ( .A1(n9850), .A2(n9719), .ZN(n7193) );
  OAI22_X1 U8746 ( .A1(n4993), .A2(n9712), .B1(n7220), .B2(n9710), .ZN(n7191)
         );
  INV_X1 U8747 ( .A(n7191), .ZN(n7192) );
  OAI211_X1 U8748 ( .C1(n9716), .C2(n7194), .A(n7193), .B(n7192), .ZN(n9848)
         );
  MUX2_X1 U8749 ( .A(n9848), .B(P1_REG2_REG_4__SCAN_IN), .S(n9309), .Z(n7195)
         );
  INV_X1 U8750 ( .A(n7195), .ZN(n7205) );
  NAND2_X1 U8751 ( .A1(n9725), .A2(n7196), .ZN(n8017) );
  INV_X1 U8752 ( .A(n8017), .ZN(n9707) );
  NAND2_X1 U8753 ( .A1(n7263), .A2(n8978), .ZN(n7197) );
  AND2_X1 U8754 ( .A1(n7280), .A2(n7197), .ZN(n9845) );
  NOR2_X1 U8755 ( .A1(n7199), .A2(n7198), .ZN(n7200) );
  NAND2_X1 U8756 ( .A1(n9845), .A2(n9706), .ZN(n7202) );
  NAND2_X1 U8757 ( .A1(n9720), .A2(n8981), .ZN(n7201) );
  OAI211_X1 U8758 ( .C1(n9847), .C2(n9723), .A(n7202), .B(n7201), .ZN(n7203)
         );
  AOI21_X1 U8759 ( .B1(n9850), .B2(n9707), .A(n7203), .ZN(n7204) );
  NAND2_X1 U8760 ( .A1(n7205), .A2(n7204), .ZN(P1_U3287) );
  INV_X1 U8761 ( .A(n7206), .ZN(n7236) );
  AOI22_X1 U8762 ( .A1(n9103), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9650), .ZN(n7207) );
  OAI21_X1 U8763 ( .B1(n7236), .B2(n9653), .A(n7207), .ZN(P1_U3335) );
  MUX2_X1 U8764 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n7208), .S(n9725), .Z(n7209)
         );
  INV_X1 U8765 ( .A(n7209), .ZN(n7218) );
  INV_X1 U8766 ( .A(n7210), .ZN(n7211) );
  NAND2_X1 U8767 ( .A1(n9706), .A2(n7211), .ZN(n7213) );
  NAND2_X1 U8768 ( .A1(n9720), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7212) );
  OAI211_X1 U8769 ( .C1(n7214), .C2(n9723), .A(n7213), .B(n7212), .ZN(n7215)
         );
  AOI21_X1 U8770 ( .B1(n7216), .B2(n9707), .A(n7215), .ZN(n7217) );
  NAND2_X1 U8771 ( .A1(n7218), .A2(n7217), .ZN(P1_U3289) );
  AOI21_X1 U8772 ( .B1(n7219), .B2(n7226), .A(n9716), .ZN(n7223) );
  OAI22_X1 U8773 ( .A1(n7220), .A2(n9712), .B1(n7336), .B2(n9710), .ZN(n7221)
         );
  AOI21_X1 U8774 ( .B1(n7223), .B2(n7222), .A(n7221), .ZN(n9864) );
  AND2_X1 U8775 ( .A1(n7225), .A2(n7224), .ZN(n7227) );
  XNOR2_X1 U8776 ( .A(n7227), .B(n7226), .ZN(n9865) );
  INV_X1 U8777 ( .A(n9865), .ZN(n9867) );
  INV_X1 U8778 ( .A(n9356), .ZN(n7270) );
  NAND2_X1 U8779 ( .A1(n9867), .A2(n7270), .ZN(n7235) );
  INV_X1 U8780 ( .A(n7228), .ZN(n7281) );
  AOI21_X1 U8781 ( .B1(n9023), .B2(n7281), .A(n7229), .ZN(n9862) );
  NOR2_X1 U8782 ( .A1(n9723), .A2(n7230), .ZN(n7233) );
  OAI22_X1 U8783 ( .A1(n9725), .A2(n6586), .B1(n7231), .B2(n9685), .ZN(n7232)
         );
  AOI211_X1 U8784 ( .C1(n9862), .C2(n9706), .A(n7233), .B(n7232), .ZN(n7234)
         );
  OAI211_X1 U8785 ( .C1(n9309), .C2(n9864), .A(n7235), .B(n7234), .ZN(P1_U3285) );
  INV_X1 U8786 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n9488) );
  INV_X1 U8787 ( .A(n8432), .ZN(n8425) );
  OAI222_X1 U8788 ( .A1(n8197), .A2(n9488), .B1(n8195), .B2(n7236), .C1(
        P2_U3152), .C2(n8425), .ZN(P2_U3340) );
  OAI22_X1 U8789 ( .A1(n9725), .A2(n6649), .B1(n7237), .B2(n9685), .ZN(n7240)
         );
  INV_X1 U8790 ( .A(n9706), .ZN(n9118) );
  AOI21_X1 U8791 ( .B1(n9118), .B2(n9723), .A(n7238), .ZN(n7239) );
  AOI211_X1 U8792 ( .C1(n9725), .C2(n7241), .A(n7240), .B(n7239), .ZN(n7242)
         );
  INV_X1 U8793 ( .A(n7242), .ZN(P1_U3291) );
  NAND2_X1 U8794 ( .A1(n7243), .A2(n9887), .ZN(n9870) );
  NOR3_X1 U8795 ( .A1(n4371), .A2(n4407), .A3(n7245), .ZN(n7248) );
  INV_X1 U8796 ( .A(n7246), .ZN(n7247) );
  OAI21_X1 U8797 ( .B1(n7248), .B2(n7247), .A(n5630), .ZN(n7253) );
  OAI22_X1 U8798 ( .A1(n9008), .A2(n7249), .B1(n9035), .B2(n8076), .ZN(n7250)
         );
  AOI211_X1 U8799 ( .C1(n9020), .C2(n9050), .A(n7251), .B(n7250), .ZN(n7252)
         );
  OAI211_X1 U8800 ( .C1(n7254), .C2(n9870), .A(n7253), .B(n7252), .ZN(P1_U3211) );
  XNOR2_X1 U8801 ( .A(n7256), .B(n7255), .ZN(n7257) );
  NAND2_X1 U8802 ( .A1(n7257), .A2(n9352), .ZN(n7259) );
  AOI22_X1 U8803 ( .A1(n9052), .A2(n9349), .B1(n9347), .B2(n9054), .ZN(n7258)
         );
  NAND2_X1 U8804 ( .A1(n7259), .A2(n7258), .ZN(n9841) );
  INV_X1 U8805 ( .A(n9841), .ZN(n7272) );
  OAI21_X1 U8806 ( .B1(n7262), .B2(n7261), .A(n7260), .ZN(n9843) );
  OAI21_X1 U8807 ( .B1(n7265), .B2(n7264), .A(n7263), .ZN(n9840) );
  INV_X1 U8808 ( .A(n9723), .ZN(n9698) );
  OAI22_X1 U8809 ( .A1(n9725), .A2(n6580), .B1(n9685), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n7266) );
  AOI21_X1 U8810 ( .B1(n9698), .B2(n7267), .A(n7266), .ZN(n7268) );
  OAI21_X1 U8811 ( .B1(n9118), .B2(n9840), .A(n7268), .ZN(n7269) );
  AOI21_X1 U8812 ( .B1(n9843), .B2(n7270), .A(n7269), .ZN(n7271) );
  OAI21_X1 U8813 ( .B1(n7272), .B2(n9309), .A(n7271), .ZN(P1_U3288) );
  OAI21_X1 U8814 ( .B1(n7279), .B2(n7274), .A(n7273), .ZN(n7275) );
  AOI222_X1 U8815 ( .A1(n9352), .A2(n7275), .B1(n9050), .B2(n9349), .C1(n9052), 
        .C2(n9347), .ZN(n9856) );
  NAND2_X1 U8816 ( .A1(n7277), .A2(n7276), .ZN(n7278) );
  AOI21_X1 U8817 ( .B1(n7279), .B2(n7278), .A(n4373), .ZN(n9859) );
  INV_X1 U8818 ( .A(n7280), .ZN(n7282) );
  OAI21_X1 U8819 ( .B1(n9853), .B2(n7282), .A(n7281), .ZN(n9855) );
  INV_X1 U8820 ( .A(n7283), .ZN(n7323) );
  OAI22_X1 U8821 ( .A1(n9725), .A2(n7284), .B1(n7323), .B2(n9685), .ZN(n7285)
         );
  AOI21_X1 U8822 ( .B1(n9698), .B2(n7286), .A(n7285), .ZN(n7287) );
  OAI21_X1 U8823 ( .B1(n9855), .B2(n9118), .A(n7287), .ZN(n7288) );
  AOI21_X1 U8824 ( .B1(n9859), .B2(n7270), .A(n7288), .ZN(n7289) );
  OAI21_X1 U8825 ( .B1(n9856), .B2(n9309), .A(n7289), .ZN(P1_U3286) );
  INV_X1 U8826 ( .A(n7290), .ZN(n7344) );
  AOI22_X1 U8827 ( .A1(n9110), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n9650), .ZN(n7291) );
  OAI21_X1 U8828 ( .B1(n7344), .B2(n9653), .A(n7291), .ZN(P1_U3334) );
  NOR2_X1 U8829 ( .A1(n7293), .A2(n7292), .ZN(n7295) );
  AND2_X1 U8830 ( .A1(n7295), .A2(n7294), .ZN(n7302) );
  INV_X1 U8831 ( .A(n7302), .ZN(n7297) );
  OR2_X1 U8832 ( .A1(n7298), .A2(n8440), .ZN(n7443) );
  NAND2_X1 U8833 ( .A1(n7719), .A2(n7443), .ZN(n7299) );
  NAND2_X1 U8834 ( .A1(n8667), .A2(n7299), .ZN(n8735) );
  INV_X1 U8835 ( .A(n7307), .ZN(n9940) );
  AOI22_X1 U8836 ( .A1(n9940), .A2(n8740), .B1(n8632), .B2(n8364), .ZN(n9942)
         );
  OAI22_X1 U8837 ( .A1(n8742), .A2(n9942), .B1(n7300), .B2(n8553), .ZN(n7301)
         );
  AOI21_X1 U8838 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n8686), .A(n7301), .ZN(
        n7306) );
  NAND2_X1 U8839 ( .A1(n7302), .A2(n8440), .ZN(n7543) );
  NOR2_X1 U8840 ( .A1(n7303), .A2(n7455), .ZN(n7304) );
  NAND2_X1 U8841 ( .A1(n8667), .A2(n7304), .ZN(n8721) );
  OAI21_X1 U8842 ( .B1(n8748), .B2(n8753), .A(n9938), .ZN(n7305) );
  OAI211_X1 U8843 ( .C1(n7307), .C2(n8735), .A(n7306), .B(n7305), .ZN(P2_U3296) );
  INV_X1 U8844 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7308) );
  OAI22_X1 U8845 ( .A1(n7543), .A2(n7309), .B1(n7308), .B2(n8553), .ZN(n7310)
         );
  AOI21_X1 U8846 ( .B1(n8753), .B2(n7311), .A(n7310), .ZN(n7315) );
  MUX2_X1 U8847 ( .A(n7313), .B(n7312), .S(n8686), .Z(n7314) );
  OAI211_X1 U8848 ( .C1(n8735), .C2(n7316), .A(n7315), .B(n7314), .ZN(P2_U3294) );
  NOR2_X1 U8849 ( .A1(n7317), .A2(n7318), .ZN(n9014) );
  AOI21_X1 U8850 ( .B1(n7317), .B2(n7318), .A(n9014), .ZN(n7319) );
  NAND2_X1 U8851 ( .A1(n7319), .A2(n7320), .ZN(n9017) );
  OAI21_X1 U8852 ( .B1(n7320), .B2(n7319), .A(n9017), .ZN(n7321) );
  NAND2_X1 U8853 ( .A1(n7321), .A2(n5630), .ZN(n7327) );
  NAND2_X1 U8854 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9794) );
  INV_X1 U8855 ( .A(n9794), .ZN(n7325) );
  OAI22_X1 U8856 ( .A1(n9008), .A2(n7323), .B1(n9035), .B2(n7322), .ZN(n7324)
         );
  AOI211_X1 U8857 ( .C1(n9020), .C2(n9052), .A(n7325), .B(n7324), .ZN(n7326)
         );
  OAI211_X1 U8858 ( .C1(n9853), .C2(n7921), .A(n7327), .B(n7326), .ZN(P1_U3225) );
  NAND2_X1 U8859 ( .A1(n7336), .A2(n7328), .ZN(n7329) );
  INV_X1 U8860 ( .A(n7334), .ZN(n7331) );
  OAI21_X1 U8861 ( .B1(n4376), .B2(n7331), .A(n7475), .ZN(n9880) );
  XOR2_X1 U8862 ( .A(n7334), .B(n7479), .Z(n7335) );
  OAI222_X1 U8863 ( .A1(n9710), .A2(n7337), .B1(n9712), .B2(n7336), .C1(n7335), 
        .C2(n9716), .ZN(n9876) );
  INV_X1 U8864 ( .A(n8071), .ZN(n7338) );
  AOI21_X1 U8865 ( .B1(n8926), .B2(n7339), .A(n7338), .ZN(n9878) );
  NAND2_X1 U8866 ( .A1(n9878), .A2(n9706), .ZN(n7341) );
  AOI22_X1 U8867 ( .A1(n9309), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n8925), .B2(
        n9720), .ZN(n7340) );
  OAI211_X1 U8868 ( .C1(n4672), .C2(n9723), .A(n7341), .B(n7340), .ZN(n7342)
         );
  AOI21_X1 U8869 ( .B1(n9876), .B2(n9725), .A(n7342), .ZN(n7343) );
  OAI21_X1 U8870 ( .B1(n9880), .B2(n9356), .A(n7343), .ZN(P1_U3283) );
  OAI222_X1 U8871 ( .A1(n8197), .A2(n7345), .B1(n8195), .B2(n7344), .C1(
        P2_U3152), .C2(n8440), .ZN(P2_U3339) );
  INV_X2 U8872 ( .A(n8667), .ZN(n8742) );
  XNOR2_X1 U8873 ( .A(n7346), .B(n6946), .ZN(n7347) );
  NAND2_X1 U8874 ( .A1(n7347), .A2(n8740), .ZN(n7349) );
  AOI22_X1 U8875 ( .A1(n8630), .A2(n6945), .B1(n7009), .B2(n8632), .ZN(n7348)
         );
  AND2_X1 U8876 ( .A1(n7349), .A2(n7348), .ZN(n9946) );
  NOR2_X1 U8877 ( .A1(n8686), .A2(n9946), .ZN(n7355) );
  INV_X1 U8878 ( .A(n7350), .ZN(n7352) );
  AOI21_X1 U8879 ( .B1(n8050), .B2(n9938), .A(n9981), .ZN(n7351) );
  NAND2_X1 U8880 ( .A1(n7352), .A2(n7351), .ZN(n9944) );
  OAI22_X1 U8881 ( .A1(n7543), .A2(n9944), .B1(n7353), .B2(n8553), .ZN(n7354)
         );
  AOI211_X1 U8882 ( .C1(n8742), .C2(P2_REG2_REG_1__SCAN_IN), .A(n7355), .B(
        n7354), .ZN(n7359) );
  INV_X1 U8883 ( .A(n8735), .ZN(n8754) );
  OAI21_X1 U8884 ( .B1(n6946), .B2(n7357), .A(n7356), .ZN(n9949) );
  AOI22_X1 U8885 ( .A1(n8754), .A2(n9949), .B1(n8753), .B2(n8050), .ZN(n7358)
         );
  NAND2_X1 U8886 ( .A1(n7359), .A2(n7358), .ZN(P2_U3295) );
  XNOR2_X1 U8887 ( .A(n9965), .B(n8175), .ZN(n7361) );
  NAND2_X1 U8888 ( .A1(n8361), .A2(n8154), .ZN(n7360) );
  NAND2_X1 U8889 ( .A1(n7361), .A2(n7360), .ZN(n7574) );
  INV_X1 U8890 ( .A(n7360), .ZN(n7363) );
  INV_X1 U8891 ( .A(n7361), .ZN(n7362) );
  NAND2_X1 U8892 ( .A1(n7363), .A2(n7362), .ZN(n7364) );
  AND2_X1 U8893 ( .A1(n7574), .A2(n7364), .ZN(n7374) );
  INV_X1 U8894 ( .A(n7365), .ZN(n7372) );
  INV_X1 U8895 ( .A(n7366), .ZN(n7371) );
  INV_X1 U8896 ( .A(n7367), .ZN(n7370) );
  INV_X1 U8897 ( .A(n7368), .ZN(n7369) );
  NAND2_X1 U8898 ( .A1(n7373), .A2(n7374), .ZN(n7577) );
  OAI21_X1 U8899 ( .B1(n7374), .B2(n7373), .A(n7577), .ZN(n7380) );
  OAI22_X1 U8900 ( .A1(n8342), .A2(n7498), .B1(n9965), .B2(n8336), .ZN(n7379)
         );
  INV_X1 U8901 ( .A(n7375), .ZN(n7548) );
  NAND2_X1 U8902 ( .A1(n8345), .A2(n8360), .ZN(n7376) );
  OAI211_X1 U8903 ( .C1(n8341), .C2(n7548), .A(n7377), .B(n7376), .ZN(n7378)
         );
  AOI211_X1 U8904 ( .C1(n7380), .C2(n8325), .A(n7379), .B(n7378), .ZN(n7381)
         );
  INV_X1 U8905 ( .A(n7381), .ZN(P2_U3241) );
  NAND2_X1 U8906 ( .A1(n7577), .A2(n7574), .ZN(n7382) );
  XNOR2_X1 U8907 ( .A(n7604), .B(n8175), .ZN(n7578) );
  NAND2_X1 U8908 ( .A1(n8360), .A2(n8154), .ZN(n7579) );
  XNOR2_X1 U8909 ( .A(n7578), .B(n7579), .ZN(n7573) );
  XNOR2_X1 U8910 ( .A(n7382), .B(n7573), .ZN(n7388) );
  OAI22_X1 U8911 ( .A1(n8336), .A2(n7604), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7383), .ZN(n7386) );
  OAI22_X1 U8912 ( .A1(n7384), .A2(n8342), .B1(n8314), .B2(n7593), .ZN(n7385)
         );
  AOI211_X1 U8913 ( .C1(n7602), .C2(n8333), .A(n7386), .B(n7385), .ZN(n7387)
         );
  OAI21_X1 U8914 ( .B1(n7388), .B2(n8349), .A(n7387), .ZN(P2_U3215) );
  NAND2_X1 U8915 ( .A1(n7397), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7390) );
  NAND2_X1 U8916 ( .A1(n7390), .A2(n7389), .ZN(n7393) );
  MUX2_X1 U8917 ( .A(n7391), .B(P2_REG2_REG_11__SCAN_IN), .S(n7562), .Z(n7392)
         );
  NOR2_X1 U8918 ( .A1(n7393), .A2(n7392), .ZN(n7554) );
  AOI21_X1 U8919 ( .B1(n7393), .B2(n7392), .A(n7554), .ZN(n7405) );
  AND2_X1 U8920 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7394) );
  AOI21_X1 U8921 ( .B1(n9920), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7394), .ZN(
        n7402) );
  INV_X1 U8922 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7395) );
  MUX2_X1 U8923 ( .A(n7395), .B(P2_REG1_REG_11__SCAN_IN), .S(n7562), .Z(n7399)
         );
  AOI21_X1 U8924 ( .B1(n7399), .B2(n7398), .A(n7561), .ZN(n7400) );
  NAND2_X1 U8925 ( .A1(n9914), .A2(n7400), .ZN(n7401) );
  OAI211_X1 U8926 ( .C1(n9915), .C2(n7555), .A(n7402), .B(n7401), .ZN(n7403)
         );
  INV_X1 U8927 ( .A(n7403), .ZN(n7404) );
  OAI21_X1 U8928 ( .B1(n7405), .B2(n9917), .A(n7404), .ZN(P2_U3256) );
  NAND2_X1 U8929 ( .A1(n7406), .A2(n7407), .ZN(n7408) );
  NAND2_X1 U8930 ( .A1(n7425), .A2(n6114), .ZN(n7427) );
  NAND2_X1 U8931 ( .A1(n6958), .A2(n7410), .ZN(n7411) );
  NAND2_X1 U8932 ( .A1(n7427), .A2(n7411), .ZN(n8751) );
  NAND2_X1 U8933 ( .A1(n7431), .A2(n9952), .ZN(n7412) );
  XNOR2_X1 U8934 ( .A(n7497), .B(n7496), .ZN(n9962) );
  NOR2_X1 U8935 ( .A1(n8686), .A2(n8554), .ZN(n8695) );
  INV_X1 U8936 ( .A(n8695), .ZN(n7417) );
  OR2_X1 U8937 ( .A1(n7436), .A2(n7445), .ZN(n8745) );
  INV_X1 U8938 ( .A(n9952), .ZN(n8752) );
  INV_X1 U8939 ( .A(n7542), .ZN(n7413) );
  OAI211_X1 U8940 ( .C1(n9960), .C2(n8744), .A(n7413), .B(n8857), .ZN(n9958)
         );
  AOI22_X1 U8941 ( .A1(n8753), .A2(n7415), .B1(n8746), .B2(n7414), .ZN(n7416)
         );
  OAI21_X1 U8942 ( .B1(n7417), .B2(n9958), .A(n7416), .ZN(n7418) );
  AOI21_X1 U8943 ( .B1(n8754), .B2(n9962), .A(n7418), .ZN(n7424) );
  XNOR2_X1 U8944 ( .A(n7419), .B(n7496), .ZN(n7421) );
  AOI21_X1 U8945 ( .B1(n7421), .B2(n8740), .A(n7420), .ZN(n9959) );
  MUX2_X1 U8946 ( .A(n9959), .B(n7422), .S(n8742), .Z(n7423) );
  NAND2_X1 U8947 ( .A1(n7424), .A2(n7423), .ZN(P2_U3291) );
  INV_X1 U8948 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7439) );
  OR2_X1 U8949 ( .A1(n7425), .A2(n6114), .ZN(n7426) );
  AND2_X1 U8950 ( .A1(n7427), .A2(n7426), .ZN(n7451) );
  NAND2_X1 U8951 ( .A1(n6954), .A2(n7428), .ZN(n7429) );
  NAND2_X1 U8952 ( .A1(n7429), .A2(n7430), .ZN(n8737) );
  OAI21_X1 U8953 ( .B1(n7430), .B2(n7429), .A(n8737), .ZN(n7434) );
  OAI22_X1 U8954 ( .A1(n7406), .A2(n8726), .B1(n7431), .B2(n8728), .ZN(n7433)
         );
  NOR2_X1 U8955 ( .A1(n7451), .A2(n7719), .ZN(n7432) );
  AOI211_X1 U8956 ( .C1(n8740), .C2(n7434), .A(n7433), .B(n7432), .ZN(n7444)
         );
  INV_X1 U8957 ( .A(n8745), .ZN(n7435) );
  AOI211_X1 U8958 ( .C1(n7445), .C2(n7436), .A(n9981), .B(n7435), .ZN(n7448)
         );
  AOI21_X1 U8959 ( .B1(n8856), .B2(n7445), .A(n7448), .ZN(n7437) );
  OAI211_X1 U8960 ( .C1(n7451), .C2(n8854), .A(n7444), .B(n7437), .ZN(n7440)
         );
  NAND2_X1 U8961 ( .A1(n7440), .A2(n10001), .ZN(n7438) );
  OAI21_X1 U8962 ( .B1(n10001), .B2(n7439), .A(n7438), .ZN(P2_U3523) );
  INV_X1 U8963 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7442) );
  NAND2_X1 U8964 ( .A1(n7440), .A2(n9988), .ZN(n7441) );
  OAI21_X1 U8965 ( .B1(n9988), .B2(n7442), .A(n7441), .ZN(P2_U3460) );
  NOR2_X1 U8966 ( .A1(n8686), .A2(n7443), .ZN(n7888) );
  INV_X1 U8967 ( .A(n7888), .ZN(n7726) );
  INV_X1 U8968 ( .A(n7444), .ZN(n7446) );
  AOI22_X1 U8969 ( .A1(n7446), .A2(n8667), .B1(n8753), .B2(n7445), .ZN(n7450)
         );
  INV_X1 U8970 ( .A(n7543), .ZN(n8679) );
  OAI22_X1 U8971 ( .A1(n8667), .A2(n6779), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8553), .ZN(n7447) );
  AOI21_X1 U8972 ( .B1(n8679), .B2(n7448), .A(n7447), .ZN(n7449) );
  OAI211_X1 U8973 ( .C1(n7451), .C2(n7726), .A(n7450), .B(n7449), .ZN(P2_U3293) );
  INV_X1 U8974 ( .A(n7452), .ZN(n7456) );
  AOI22_X1 U8975 ( .A1(n7453), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n9650), .ZN(n7454) );
  OAI21_X1 U8976 ( .B1(n7456), .B2(n9653), .A(n7454), .ZN(P1_U3333) );
  OAI222_X1 U8977 ( .A1(n8197), .A2(n7457), .B1(n8195), .B2(n7456), .C1(n7455), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  INV_X1 U8978 ( .A(n7686), .ZN(n7677) );
  NAND2_X1 U8979 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8038) );
  INV_X1 U8980 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7458) );
  MUX2_X1 U8981 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n7458), .S(n7686), .Z(n7461)
         );
  OAI21_X1 U8982 ( .B1(n7465), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7459), .ZN(
        n7460) );
  NAND2_X1 U8983 ( .A1(n7461), .A2(n7460), .ZN(n7685) );
  OAI21_X1 U8984 ( .B1(n7461), .B2(n7460), .A(n7685), .ZN(n7462) );
  NAND2_X1 U8985 ( .A1(n9823), .A2(n7462), .ZN(n7463) );
  OAI211_X1 U8986 ( .C1(n9060), .C2(n7677), .A(n8038), .B(n7463), .ZN(n7469)
         );
  INV_X1 U8987 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7466) );
  AOI211_X1 U8988 ( .C1(n7467), .C2(n7466), .A(n7679), .B(n9817), .ZN(n7468)
         );
  AOI211_X1 U8989 ( .C1(P1_ADDR_REG_14__SCAN_IN), .C2(n9827), .A(n7469), .B(
        n7468), .ZN(n7470) );
  INV_X1 U8990 ( .A(n7470), .ZN(P1_U3255) );
  INV_X1 U8991 ( .A(n7471), .ZN(n7494) );
  AOI22_X1 U8992 ( .A1(n7472), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n9650), .ZN(n7473) );
  OAI21_X1 U8993 ( .B1(n7494), .B2(n9653), .A(n7473), .ZN(P1_U3332) );
  INV_X1 U8994 ( .A(n8076), .ZN(n9048) );
  NAND2_X1 U8995 ( .A1(n8926), .A2(n9048), .ZN(n7474) );
  OR2_X1 U8996 ( .A1(n9886), .A2(n9047), .ZN(n7476) );
  XNOR2_X1 U8997 ( .A(n7744), .B(n7477), .ZN(n9674) );
  INV_X1 U8998 ( .A(n7481), .ZN(n7483) );
  OAI21_X1 U8999 ( .B1(n8075), .B2(n7483), .A(n7482), .ZN(n7484) );
  XNOR2_X1 U9000 ( .A(n7484), .B(n7743), .ZN(n7485) );
  NAND2_X1 U9001 ( .A1(n7485), .A2(n9352), .ZN(n7487) );
  AOI22_X1 U9002 ( .A1(n9347), .A2(n9047), .B1(n9045), .B2(n9349), .ZN(n7486)
         );
  NAND2_X1 U9003 ( .A1(n7487), .A2(n7486), .ZN(n9669) );
  INV_X1 U9004 ( .A(n9671), .ZN(n7490) );
  AOI211_X1 U9005 ( .C1(n9671), .C2(n8069), .A(n9854), .B(n9702), .ZN(n9670)
         );
  NAND2_X1 U9006 ( .A1(n9670), .A2(n7982), .ZN(n7489) );
  AOI22_X1 U9007 ( .A1(n9309), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n8062), .B2(
        n9720), .ZN(n7488) );
  OAI211_X1 U9008 ( .C1(n7490), .C2(n9723), .A(n7489), .B(n7488), .ZN(n7491)
         );
  AOI21_X1 U9009 ( .B1(n9725), .B2(n9669), .A(n7491), .ZN(n7492) );
  OAI21_X1 U9010 ( .B1(n9674), .B2(n9356), .A(n7492), .ZN(P1_U3281) );
  OAI222_X1 U9011 ( .A1(n8197), .A2(n7495), .B1(n8195), .B2(n7494), .C1(n7493), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  NOR2_X1 U9012 ( .A1(n8361), .A2(n7499), .ZN(n7501) );
  NAND2_X1 U9013 ( .A1(n8361), .A2(n7499), .ZN(n7500) );
  XNOR2_X1 U9014 ( .A(n7788), .B(n6165), .ZN(n7610) );
  XNOR2_X1 U9015 ( .A(n7502), .B(n7707), .ZN(n7503) );
  AOI222_X1 U9016 ( .A1(n8740), .A2(n7503), .B1(n8359), .B2(n8632), .C1(n8361), 
        .C2(n8630), .ZN(n7605) );
  INV_X1 U9017 ( .A(n7604), .ZN(n7504) );
  AOI21_X1 U9018 ( .B1(n7504), .B2(n7541), .A(n4370), .ZN(n7608) );
  AOI22_X1 U9019 ( .A1(n7608), .A2(n8857), .B1(n8856), .B2(n7504), .ZN(n7505)
         );
  OAI211_X1 U9020 ( .C1(n8861), .C2(n7610), .A(n7605), .B(n7505), .ZN(n8863)
         );
  NAND2_X1 U9021 ( .A1(n8863), .A2(n9988), .ZN(n7506) );
  OAI21_X1 U9022 ( .B1(n9988), .B2(n5768), .A(n7506), .ZN(P2_U3472) );
  AND2_X1 U9023 ( .A1(n8359), .A2(n8239), .ZN(n7508) );
  OR2_X2 U9024 ( .A1(n7707), .A2(n7508), .ZN(n7512) );
  OR2_X1 U9025 ( .A1(n7788), .A2(n7512), .ZN(n7510) );
  INV_X1 U9026 ( .A(n8360), .ZN(n7507) );
  NAND2_X1 U9027 ( .A1(n7507), .A2(n7604), .ZN(n7708) );
  INV_X1 U9028 ( .A(n7508), .ZN(n7509) );
  NAND2_X1 U9029 ( .A1(n7510), .A2(n7511), .ZN(n7515) );
  OR2_X1 U9030 ( .A1(n7788), .A2(n7786), .ZN(n7660) );
  AND2_X1 U9031 ( .A1(n7656), .A2(n7660), .ZN(n7513) );
  OAI21_X1 U9032 ( .B1(n7515), .B2(n7514), .A(n7513), .ZN(n7767) );
  INV_X1 U9033 ( .A(n7719), .ZN(n7882) );
  XNOR2_X1 U9034 ( .A(n7516), .B(n7517), .ZN(n7518) );
  NAND2_X1 U9035 ( .A1(n7518), .A2(n8740), .ZN(n7520) );
  AOI22_X1 U9036 ( .A1(n8630), .A2(n8359), .B1(n8357), .B2(n8632), .ZN(n7519)
         );
  NAND2_X1 U9037 ( .A1(n7520), .A2(n7519), .ZN(n7521) );
  AOI21_X1 U9038 ( .B1(n7767), .B2(n7882), .A(n7521), .ZN(n7769) );
  NOR2_X1 U9039 ( .A1(n7720), .A2(n7764), .ZN(n7522) );
  OR2_X1 U9040 ( .A1(n7670), .A2(n7522), .ZN(n7765) );
  NAND2_X1 U9041 ( .A1(n8742), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7523) );
  OAI21_X1 U9042 ( .B1(n8553), .B2(n7597), .A(n7523), .ZN(n7524) );
  AOI21_X1 U9043 ( .B1(n8753), .B2(n7655), .A(n7524), .ZN(n7525) );
  OAI21_X1 U9044 ( .B1(n8530), .B2(n7765), .A(n7525), .ZN(n7526) );
  AOI21_X1 U9045 ( .B1(n7767), .B2(n7888), .A(n7526), .ZN(n7527) );
  OAI21_X1 U9046 ( .B1(n7769), .B2(n8742), .A(n7527), .ZN(P2_U3287) );
  INV_X1 U9047 ( .A(n7528), .ZN(n7529) );
  AOI21_X1 U9048 ( .B1(n7530), .B2(n4450), .A(n7529), .ZN(n7536) );
  INV_X1 U9049 ( .A(n8072), .ZN(n7531) );
  OAI22_X1 U9050 ( .A1(n9008), .A2(n7531), .B1(n9035), .B2(n9713), .ZN(n7532)
         );
  AOI211_X1 U9051 ( .C1(n9020), .C2(n9048), .A(n7533), .B(n7532), .ZN(n7535)
         );
  NAND2_X1 U9052 ( .A1(n9038), .A2(n9886), .ZN(n7534) );
  OAI211_X1 U9053 ( .C1(n7536), .C2(n9012), .A(n7535), .B(n7534), .ZN(P1_U3229) );
  INV_X1 U9054 ( .A(n7537), .ZN(n8194) );
  AOI22_X1 U9055 ( .A1(n7538), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n9650), .ZN(n7539) );
  OAI21_X1 U9056 ( .B1(n8194), .B2(n9653), .A(n7539), .ZN(P1_U3331) );
  XOR2_X1 U9057 ( .A(n7546), .B(n7540), .Z(n9967) );
  OAI211_X1 U9058 ( .C1(n7542), .C2(n9965), .A(n8857), .B(n7541), .ZN(n9963)
         );
  OAI22_X1 U9059 ( .A1(n8721), .A2(n9965), .B1(n7543), .B2(n9963), .ZN(n7551)
         );
  OAI21_X1 U9060 ( .B1(n7546), .B2(n7544), .A(n7545), .ZN(n7547) );
  AOI222_X1 U9061 ( .A1(n8740), .A2(n7547), .B1(n8360), .B2(n8632), .C1(n8362), 
        .C2(n8630), .ZN(n9964) );
  OAI21_X1 U9062 ( .B1(n7548), .B2(n8553), .A(n9964), .ZN(n7549) );
  MUX2_X1 U9063 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7549), .S(n8667), .Z(n7550)
         );
  AOI211_X1 U9064 ( .C1(n8754), .C2(n9967), .A(n7551), .B(n7550), .ZN(n7552)
         );
  INV_X1 U9065 ( .A(n7552), .ZN(P2_U3290) );
  NAND2_X1 U9066 ( .A1(n8369), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7556) );
  MUX2_X1 U9067 ( .A(n5842), .B(P2_REG2_REG_12__SCAN_IN), .S(n8369), .Z(n7553)
         );
  INV_X1 U9068 ( .A(n7553), .ZN(n8366) );
  AOI21_X1 U9069 ( .B1(n7555), .B2(n7391), .A(n7554), .ZN(n8367) );
  NAND2_X1 U9070 ( .A1(n8366), .A2(n8367), .ZN(n8365) );
  NAND2_X1 U9071 ( .A1(n7556), .A2(n8365), .ZN(n7558) );
  AOI22_X1 U9072 ( .A1(n7734), .A2(n5854), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7559), .ZN(n7557) );
  NOR2_X1 U9073 ( .A1(n7558), .A2(n7557), .ZN(n7727) );
  AOI21_X1 U9074 ( .B1(n7558), .B2(n7557), .A(n7727), .ZN(n7572) );
  INV_X1 U9075 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7560) );
  AOI22_X1 U9076 ( .A1(n7734), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n7560), .B2(
        n7559), .ZN(n7565) );
  INV_X1 U9077 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7563) );
  MUX2_X1 U9078 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7563), .S(n8369), .Z(n8372)
         );
  OAI21_X1 U9079 ( .B1(n8369), .B2(P2_REG1_REG_12__SCAN_IN), .A(n8370), .ZN(
        n7564) );
  NAND2_X1 U9080 ( .A1(n7565), .A2(n7564), .ZN(n7733) );
  OAI21_X1 U9081 ( .B1(n7565), .B2(n7564), .A(n7733), .ZN(n7566) );
  NAND2_X1 U9082 ( .A1(n7566), .A2(n9914), .ZN(n7571) );
  INV_X1 U9083 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7568) );
  OAI22_X1 U9084 ( .A1(n8446), .A2(n7568), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7567), .ZN(n7569) );
  AOI21_X1 U9085 ( .B1(n8388), .B2(n7734), .A(n7569), .ZN(n7570) );
  OAI211_X1 U9086 ( .C1(n7572), .C2(n9917), .A(n7571), .B(n7570), .ZN(P2_U3258) );
  INV_X1 U9087 ( .A(n7573), .ZN(n7575) );
  AND2_X1 U9088 ( .A1(n7575), .A2(n7574), .ZN(n7576) );
  NAND2_X1 U9089 ( .A1(n7577), .A2(n7576), .ZN(n7583) );
  INV_X1 U9090 ( .A(n7578), .ZN(n7581) );
  INV_X1 U9091 ( .A(n7579), .ZN(n7580) );
  NAND2_X1 U9092 ( .A1(n7581), .A2(n7580), .ZN(n7582) );
  NAND2_X1 U9093 ( .A1(n7583), .A2(n7582), .ZN(n8237) );
  XNOR2_X1 U9094 ( .A(n8239), .B(n8175), .ZN(n7586) );
  NAND2_X1 U9095 ( .A1(n8359), .A2(n8154), .ZN(n7584) );
  XNOR2_X1 U9096 ( .A(n7586), .B(n7584), .ZN(n8236) );
  INV_X1 U9097 ( .A(n7584), .ZN(n7585) );
  AND2_X1 U9098 ( .A1(n7586), .A2(n7585), .ZN(n7587) );
  AOI21_X2 U9099 ( .B1(n8237), .B2(n8236), .A(n7587), .ZN(n7632) );
  XNOR2_X1 U9100 ( .A(n7764), .B(n8175), .ZN(n7588) );
  NAND2_X1 U9101 ( .A1(n8358), .A2(n8154), .ZN(n7589) );
  NAND2_X1 U9102 ( .A1(n7588), .A2(n7589), .ZN(n8213) );
  INV_X1 U9103 ( .A(n7588), .ZN(n7591) );
  INV_X1 U9104 ( .A(n7589), .ZN(n7590) );
  NAND2_X1 U9105 ( .A1(n7591), .A2(n7590), .ZN(n7592) );
  AND2_X1 U9106 ( .A1(n8213), .A2(n7592), .ZN(n7630) );
  NAND2_X1 U9107 ( .A1(n7632), .A2(n7630), .ZN(n8214) );
  OAI21_X1 U9108 ( .B1(n7632), .B2(n7630), .A(n8214), .ZN(n7600) );
  OAI22_X1 U9109 ( .A1(n8342), .A2(n7593), .B1(n7764), .B2(n8336), .ZN(n7599)
         );
  INV_X1 U9110 ( .A(n7594), .ZN(n7596) );
  NAND2_X1 U9111 ( .A1(n8345), .A2(n8357), .ZN(n7595) );
  OAI211_X1 U9112 ( .C1(n8341), .C2(n7597), .A(n7596), .B(n7595), .ZN(n7598)
         );
  AOI211_X1 U9113 ( .C1(n7600), .C2(n8325), .A(n7599), .B(n7598), .ZN(n7601)
         );
  INV_X1 U9114 ( .A(n7601), .ZN(P2_U3233) );
  AOI22_X1 U9115 ( .A1(n8742), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n7602), .B2(
        n8746), .ZN(n7603) );
  OAI21_X1 U9116 ( .B1(n7604), .B2(n8721), .A(n7603), .ZN(n7607) );
  NOR2_X1 U9117 ( .A1(n7605), .A2(n8686), .ZN(n7606) );
  AOI211_X1 U9118 ( .C1(n7608), .C2(n8748), .A(n7607), .B(n7606), .ZN(n7609)
         );
  OAI21_X1 U9119 ( .B1(n8735), .B2(n7610), .A(n7609), .ZN(P2_U3289) );
  XNOR2_X1 U9120 ( .A(n7902), .B(n8168), .ZN(n7611) );
  NAND2_X1 U9121 ( .A1(n8355), .A2(n8154), .ZN(n7612) );
  NAND2_X1 U9122 ( .A1(n7611), .A2(n7612), .ZN(n8088) );
  INV_X1 U9123 ( .A(n7611), .ZN(n7614) );
  INV_X1 U9124 ( .A(n7612), .ZN(n7613) );
  NAND2_X1 U9125 ( .A1(n7614), .A2(n7613), .ZN(n7615) );
  NAND2_X1 U9126 ( .A1(n8088), .A2(n7615), .ZN(n7637) );
  XNOR2_X1 U9127 ( .A(n9974), .B(n8175), .ZN(n7622) );
  NAND2_X1 U9128 ( .A1(n8357), .A2(n8154), .ZN(n7623) );
  XNOR2_X1 U9129 ( .A(n7622), .B(n7623), .ZN(n8216) );
  INV_X1 U9130 ( .A(n8216), .ZN(n7616) );
  AND2_X1 U9131 ( .A1(n7616), .A2(n8213), .ZN(n7643) );
  XNOR2_X1 U9132 ( .A(n8855), .B(n8175), .ZN(n7619) );
  NAND2_X1 U9133 ( .A1(n8356), .A2(n8154), .ZN(n7618) );
  INV_X1 U9134 ( .A(n7618), .ZN(n7617) );
  NAND2_X1 U9135 ( .A1(n7619), .A2(n7617), .ZN(n7626) );
  INV_X1 U9136 ( .A(n7626), .ZN(n7620) );
  XNOR2_X1 U9137 ( .A(n7619), .B(n7618), .ZN(n7646) );
  AND2_X1 U9138 ( .A1(n7643), .A2(n7621), .ZN(n7634) );
  NAND2_X1 U9139 ( .A1(n8214), .A2(n7634), .ZN(n7627) );
  INV_X1 U9140 ( .A(n7622), .ZN(n7625) );
  INV_X1 U9141 ( .A(n7623), .ZN(n7624) );
  NAND2_X1 U9142 ( .A1(n7625), .A2(n7624), .ZN(n7644) );
  NAND2_X1 U9143 ( .A1(n7627), .A2(n7629), .ZN(n7636) );
  INV_X1 U9144 ( .A(n7637), .ZN(n7628) );
  AND2_X1 U9145 ( .A1(n7630), .A2(n7633), .ZN(n7631) );
  NAND2_X1 U9146 ( .A1(n7632), .A2(n7631), .ZN(n8090) );
  OR2_X1 U9147 ( .A1(n7635), .A2(n7634), .ZN(n8087) );
  AOI21_X1 U9148 ( .B1(n7637), .B2(n7636), .A(n4374), .ZN(n7642) );
  AOI22_X1 U9149 ( .A1(n8240), .A2(n8356), .B1(n8333), .B2(n7901), .ZN(n7639)
         );
  NOR2_X1 U9150 ( .A1(n9503), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8368) );
  INV_X1 U9151 ( .A(n8368), .ZN(n7638) );
  OAI211_X1 U9152 ( .C1(n7994), .C2(n8314), .A(n7639), .B(n7638), .ZN(n7640)
         );
  AOI21_X1 U9153 ( .B1(n8346), .B2(n7902), .A(n7640), .ZN(n7641) );
  OAI21_X1 U9154 ( .B1(n7642), .B2(n8349), .A(n7641), .ZN(P2_U3226) );
  NAND2_X1 U9155 ( .A1(n8214), .A2(n7643), .ZN(n7645) );
  NAND2_X1 U9156 ( .A1(n7645), .A2(n7644), .ZN(n7647) );
  XNOR2_X1 U9157 ( .A(n7647), .B(n7646), .ZN(n7654) );
  INV_X1 U9158 ( .A(n7795), .ZN(n7651) );
  NAND2_X1 U9159 ( .A1(n8355), .A2(n8632), .ZN(n7649) );
  NAND2_X1 U9160 ( .A1(n8357), .A2(n8630), .ZN(n7648) );
  NAND2_X1 U9161 ( .A1(n7649), .A2(n7648), .ZN(n7800) );
  AOI22_X1 U9162 ( .A1(n8282), .A2(n7800), .B1(P2_REG3_REG_11__SCAN_IN), .B2(
        P2_U3152), .ZN(n7650) );
  OAI21_X1 U9163 ( .B1(n8341), .B2(n7651), .A(n7650), .ZN(n7652) );
  AOI21_X1 U9164 ( .B1(n8346), .B2(n8855), .A(n7652), .ZN(n7653) );
  OAI21_X1 U9165 ( .B1(n7654), .B2(n8349), .A(n7653), .ZN(P2_U3238) );
  INV_X1 U9166 ( .A(n7664), .ZN(n7658) );
  OR2_X1 U9167 ( .A1(n8358), .A2(n7655), .ZN(n7657) );
  AND2_X2 U9168 ( .A1(n7658), .A2(n7659), .ZN(n7789) );
  NAND2_X1 U9169 ( .A1(n7660), .A2(n7789), .ZN(n7663) );
  NAND2_X1 U9170 ( .A1(n7660), .A2(n7659), .ZN(n7661) );
  NAND2_X1 U9171 ( .A1(n7661), .A2(n7664), .ZN(n7662) );
  NAND2_X1 U9172 ( .A1(n7663), .A2(n7662), .ZN(n7669) );
  XOR2_X1 U9173 ( .A(n4375), .B(n7664), .Z(n7667) );
  OAI22_X1 U9174 ( .A1(n7665), .A2(n8726), .B1(n7897), .B2(n8728), .ZN(n7666)
         );
  AOI21_X1 U9175 ( .B1(n7667), .B2(n8740), .A(n7666), .ZN(n7668) );
  OAI21_X1 U9176 ( .B1(n7669), .B2(n7719), .A(n7668), .ZN(n9976) );
  INV_X1 U9177 ( .A(n9976), .ZN(n7676) );
  INV_X1 U9178 ( .A(n7669), .ZN(n9978) );
  NAND2_X1 U9179 ( .A1(n7670), .A2(n9974), .ZN(n7794) );
  OR2_X1 U9180 ( .A1(n7670), .A2(n9974), .ZN(n7671) );
  NAND2_X1 U9181 ( .A1(n7794), .A2(n7671), .ZN(n9975) );
  AOI22_X1 U9182 ( .A1(n8742), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n8220), .B2(
        n8746), .ZN(n7673) );
  NAND2_X1 U9183 ( .A1(n8753), .A2(n8218), .ZN(n7672) );
  OAI211_X1 U9184 ( .C1(n9975), .C2(n8530), .A(n7673), .B(n7672), .ZN(n7674)
         );
  AOI21_X1 U9185 ( .B1(n9978), .B2(n7888), .A(n7674), .ZN(n7675) );
  OAI21_X1 U9186 ( .B1(n7676), .B2(n8742), .A(n7675), .ZN(P2_U3286) );
  INV_X1 U9187 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7693) );
  NOR2_X1 U9188 ( .A1(n7678), .A2(n7677), .ZN(n7680) );
  INV_X1 U9189 ( .A(n7681), .ZN(n7684) );
  INV_X1 U9190 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7682) );
  NOR2_X1 U9191 ( .A1(n7682), .A2(n7681), .ZN(n7923) );
  INV_X1 U9192 ( .A(n7923), .ZN(n7683) );
  OAI211_X1 U9193 ( .C1(n7684), .C2(P1_REG2_REG_15__SCAN_IN), .A(n9798), .B(
        n7683), .ZN(n7692) );
  NAND2_X1 U9194 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8031) );
  INV_X1 U9195 ( .A(n8031), .ZN(n7689) );
  OAI21_X1 U9196 ( .B1(n7686), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7685), .ZN(
        n7928) );
  XNOR2_X1 U9197 ( .A(n7929), .B(n7928), .ZN(n7687) );
  INV_X1 U9198 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9601) );
  NOR2_X1 U9199 ( .A1(n9601), .A2(n7687), .ZN(n7930) );
  AOI211_X1 U9200 ( .C1(n7687), .C2(n9601), .A(n7930), .B(n9072), .ZN(n7688)
         );
  AOI211_X1 U9201 ( .C1(n9825), .C2(n7690), .A(n7689), .B(n7688), .ZN(n7691)
         );
  OAI211_X1 U9202 ( .C1(n9773), .C2(n7693), .A(n7692), .B(n7691), .ZN(P1_U3256) );
  INV_X1 U9203 ( .A(n7753), .ZN(n9735) );
  OAI211_X1 U9204 ( .C1(n7696), .C2(n7695), .A(n7694), .B(n5630), .ZN(n7700)
         );
  INV_X1 U9205 ( .A(n9711), .ZN(n9044) );
  AND2_X1 U9206 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3084), .ZN(n9062) );
  INV_X1 U9207 ( .A(n9721), .ZN(n7697) );
  OAI22_X1 U9208 ( .A1(n9008), .A2(n7697), .B1(n9032), .B2(n9713), .ZN(n7698)
         );
  AOI211_X1 U9209 ( .C1(n9022), .C2(n9044), .A(n9062), .B(n7698), .ZN(n7699)
         );
  OAI211_X1 U9210 ( .C1(n9735), .C2(n7921), .A(n7700), .B(n7699), .ZN(P1_U3234) );
  INV_X1 U9211 ( .A(n7701), .ZN(n7706) );
  AOI21_X1 U9212 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8889), .A(n7702), .ZN(
        n7703) );
  OAI21_X1 U9213 ( .B1(n7706), .B2(n8195), .A(n7703), .ZN(P2_U3335) );
  AOI21_X1 U9214 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9650), .A(n7704), .ZN(
        n7705) );
  OAI21_X1 U9215 ( .B1(n7706), .B2(n9653), .A(n7705), .ZN(P1_U3330) );
  OR2_X1 U9216 ( .A1(n7788), .A2(n7707), .ZN(n7711) );
  AND2_X1 U9217 ( .A1(n7711), .A2(n7708), .ZN(n7713) );
  INV_X1 U9218 ( .A(n7709), .ZN(n7710) );
  NAND2_X1 U9219 ( .A1(n7711), .A2(n7710), .ZN(n7712) );
  OAI21_X1 U9220 ( .B1(n7713), .B2(n7714), .A(n7712), .ZN(n9968) );
  AOI22_X1 U9221 ( .A1(n8630), .A2(n8360), .B1(n8358), .B2(n8632), .ZN(n7718)
         );
  XNOR2_X1 U9222 ( .A(n7715), .B(n7714), .ZN(n7716) );
  NAND2_X1 U9223 ( .A1(n7716), .A2(n8740), .ZN(n7717) );
  OAI211_X1 U9224 ( .C1(n9968), .C2(n7719), .A(n7718), .B(n7717), .ZN(n9971)
         );
  NAND2_X1 U9225 ( .A1(n9971), .A2(n8667), .ZN(n7725) );
  INV_X1 U9226 ( .A(n7720), .ZN(n7721) );
  OAI21_X1 U9227 ( .B1(n9969), .B2(n4370), .A(n7721), .ZN(n9970) );
  AOI22_X1 U9228 ( .A1(n8742), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n8242), .B2(
        n8746), .ZN(n7722) );
  OAI21_X1 U9229 ( .B1(n9970), .B2(n8530), .A(n7722), .ZN(n7723) );
  AOI21_X1 U9230 ( .B1(n8753), .B2(n8239), .A(n7723), .ZN(n7724) );
  OAI211_X1 U9231 ( .C1(n9968), .C2(n7726), .A(n7725), .B(n7724), .ZN(P2_U3288) );
  NOR2_X1 U9232 ( .A1(n7734), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7728) );
  NOR2_X1 U9233 ( .A1(n7728), .A2(n7727), .ZN(n7730) );
  AOI22_X1 U9234 ( .A1(n7955), .A2(n5872), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7731), .ZN(n7729) );
  NOR2_X1 U9235 ( .A1(n7730), .A2(n7729), .ZN(n7956) );
  AOI21_X1 U9236 ( .B1(n7730), .B2(n7729), .A(n7956), .ZN(n7742) );
  INV_X1 U9237 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7732) );
  AOI22_X1 U9238 ( .A1(n7955), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n7732), .B2(
        n7731), .ZN(n7736) );
  OAI21_X1 U9239 ( .B1(n7734), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7733), .ZN(
        n7735) );
  NAND2_X1 U9240 ( .A1(n7736), .A2(n7735), .ZN(n7951) );
  OAI21_X1 U9241 ( .B1(n7736), .B2(n7735), .A(n7951), .ZN(n7737) );
  NAND2_X1 U9242 ( .A1(n7737), .A2(n9914), .ZN(n7741) );
  INV_X1 U9243 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U9244 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8096) );
  OAI21_X1 U9245 ( .B1(n8446), .B2(n7738), .A(n8096), .ZN(n7739) );
  AOI21_X1 U9246 ( .B1(n8388), .B2(n7955), .A(n7739), .ZN(n7740) );
  OAI211_X1 U9247 ( .C1(n7742), .C2(n9917), .A(n7741), .B(n7740), .ZN(P2_U3259) );
  NAND2_X1 U9248 ( .A1(n7744), .A2(n7743), .ZN(n7746) );
  INV_X1 U9249 ( .A(n9713), .ZN(n9046) );
  OR2_X1 U9250 ( .A1(n9671), .A2(n9046), .ZN(n7745) );
  NAND2_X1 U9251 ( .A1(n7746), .A2(n7745), .ZN(n9701) );
  NOR2_X1 U9252 ( .A1(n7753), .A2(n9045), .ZN(n7747) );
  NAND2_X1 U9253 ( .A1(n7753), .A2(n9045), .ZN(n7748) );
  XNOR2_X1 U9254 ( .A(n7818), .B(n7822), .ZN(n7808) );
  NAND2_X1 U9255 ( .A1(n8075), .A2(n7750), .ZN(n7752) );
  NAND2_X1 U9256 ( .A1(n7752), .A2(n7751), .ZN(n9709) );
  OR2_X1 U9257 ( .A1(n7753), .A2(n8064), .ZN(n7754) );
  NAND2_X1 U9258 ( .A1(n9709), .A2(n7754), .ZN(n7756) );
  NAND2_X1 U9259 ( .A1(n7756), .A2(n7755), .ZN(n7826) );
  XNOR2_X1 U9260 ( .A(n7826), .B(n7822), .ZN(n7757) );
  OAI222_X1 U9261 ( .A1(n9710), .A2(n8040), .B1(n9712), .B2(n8064), .C1(n7757), 
        .C2(n9716), .ZN(n7805) );
  INV_X1 U9262 ( .A(n7816), .ZN(n7761) );
  NAND2_X1 U9263 ( .A1(n9702), .A2(n9735), .ZN(n9704) );
  INV_X1 U9264 ( .A(n4828), .ZN(n7758) );
  AOI211_X1 U9265 ( .C1(n7816), .C2(n9704), .A(n9854), .B(n7758), .ZN(n7806)
         );
  NAND2_X1 U9266 ( .A1(n7806), .A2(n7982), .ZN(n7760) );
  AOI22_X1 U9267 ( .A1(n9309), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7777), .B2(
        n9720), .ZN(n7759) );
  OAI211_X1 U9268 ( .C1(n7761), .C2(n9723), .A(n7760), .B(n7759), .ZN(n7762)
         );
  AOI21_X1 U9269 ( .B1(n9725), .B2(n7805), .A(n7762), .ZN(n7763) );
  OAI21_X1 U9270 ( .B1(n7808), .B2(n9356), .A(n7763), .ZN(P1_U3279) );
  INV_X1 U9271 ( .A(n8854), .ZN(n9979) );
  OAI22_X1 U9272 ( .A1(n7765), .A2(n9981), .B1(n7764), .B2(n9980), .ZN(n7766)
         );
  AOI21_X1 U9273 ( .B1(n7767), .B2(n9979), .A(n7766), .ZN(n7768) );
  AND2_X1 U9274 ( .A1(n7769), .A2(n7768), .ZN(n7771) );
  MUX2_X1 U9275 ( .A(n5801), .B(n7771), .S(n9988), .Z(n7770) );
  INV_X1 U9276 ( .A(n7770), .ZN(P2_U3478) );
  MUX2_X1 U9277 ( .A(n6902), .B(n7771), .S(n10001), .Z(n7772) );
  INV_X1 U9278 ( .A(n7772), .ZN(P2_U3529) );
  XNOR2_X1 U9279 ( .A(n7774), .B(n7773), .ZN(n7775) );
  XNOR2_X1 U9280 ( .A(n7776), .B(n7775), .ZN(n7782) );
  AOI22_X1 U9281 ( .A1(n9020), .A2(n9045), .B1(n9033), .B2(n7777), .ZN(n7779)
         );
  OAI211_X1 U9282 ( .C1(n8040), .C2(n9035), .A(n7779), .B(n7778), .ZN(n7780)
         );
  AOI21_X1 U9283 ( .B1(n7816), .B2(n9038), .A(n7780), .ZN(n7781) );
  OAI21_X1 U9284 ( .B1(n7782), .B2(n9012), .A(n7781), .ZN(P1_U3222) );
  INV_X1 U9285 ( .A(n7783), .ZN(n7812) );
  AOI22_X1 U9286 ( .A1(n7784), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n9647), .ZN(n7785) );
  OAI21_X1 U9287 ( .B1(n7812), .B2(n9653), .A(n7785), .ZN(P1_U3329) );
  AND2_X1 U9288 ( .A1(n8218), .A2(n8357), .ZN(n7790) );
  INV_X1 U9289 ( .A(n7789), .ZN(n7792) );
  INV_X1 U9290 ( .A(n7790), .ZN(n7791) );
  AND2_X1 U9291 ( .A1(n7869), .A2(n7866), .ZN(n7793) );
  XNOR2_X1 U9292 ( .A(n7793), .B(n7865), .ZN(n8862) );
  INV_X1 U9293 ( .A(n7883), .ZN(n7900) );
  AOI21_X1 U9294 ( .B1(n8855), .B2(n7794), .A(n7900), .ZN(n8858) );
  INV_X1 U9295 ( .A(n8855), .ZN(n7797) );
  AOI22_X1 U9296 ( .A1(n8742), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7795), .B2(
        n8746), .ZN(n7796) );
  OAI21_X1 U9297 ( .B1(n7797), .B2(n8721), .A(n7796), .ZN(n7803) );
  XNOR2_X1 U9298 ( .A(n7798), .B(n7799), .ZN(n7801) );
  AOI21_X1 U9299 ( .B1(n7801), .B2(n8740), .A(n7800), .ZN(n8860) );
  NOR2_X1 U9300 ( .A1(n8860), .A2(n8742), .ZN(n7802) );
  AOI211_X1 U9301 ( .C1(n8858), .C2(n8748), .A(n7803), .B(n7802), .ZN(n7804)
         );
  OAI21_X1 U9302 ( .B1(n8735), .B2(n8862), .A(n7804), .ZN(P2_U3285) );
  INV_X1 U9303 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7810) );
  AOI211_X1 U9304 ( .C1(n9887), .C2(n7816), .A(n7806), .B(n7805), .ZN(n7807)
         );
  OAI21_X1 U9305 ( .B1(n7808), .B2(n9892), .A(n7807), .ZN(n7814) );
  NAND2_X1 U9306 ( .A1(n7814), .A2(n9897), .ZN(n7809) );
  OAI21_X1 U9307 ( .B1(n9897), .B2(n7810), .A(n7809), .ZN(P1_U3490) );
  OAI222_X1 U9308 ( .A1(P2_U3152), .A2(n7813), .B1(n8195), .B2(n7812), .C1(
        n7811), .C2(n8197), .ZN(P2_U3334) );
  NAND2_X1 U9309 ( .A1(n7814), .A2(n9911), .ZN(n7815) );
  OAI21_X1 U9310 ( .B1(n9911), .B2(n6973), .A(n7815), .ZN(P1_U3535) );
  AND2_X1 U9311 ( .A1(n7816), .A2(n9044), .ZN(n7817) );
  NAND2_X1 U9312 ( .A1(n9729), .A2(n8040), .ZN(n7819) );
  XOR2_X1 U9313 ( .A(n7972), .B(n7829), .Z(n9448) );
  INV_X1 U9314 ( .A(n9682), .ZN(n7820) );
  AOI211_X1 U9315 ( .C1(n9445), .C2(n7820), .A(n9854), .B(n8013), .ZN(n9444)
         );
  AOI22_X1 U9316 ( .A1(n9309), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8037), .B2(
        n9720), .ZN(n7821) );
  OAI21_X1 U9317 ( .B1(n7973), .B2(n9723), .A(n7821), .ZN(n7833) );
  INV_X1 U9318 ( .A(n7822), .ZN(n7825) );
  INV_X1 U9319 ( .A(n7823), .ZN(n7824) );
  AOI211_X1 U9320 ( .C1(n7829), .C2(n7828), .A(n9716), .B(n4367), .ZN(n7831)
         );
  OAI22_X1 U9321 ( .A1(n8040), .A2(n9712), .B1(n7976), .B2(n9710), .ZN(n7830)
         );
  NOR2_X1 U9322 ( .A1(n7831), .A2(n7830), .ZN(n9447) );
  NOR2_X1 U9323 ( .A1(n9447), .A2(n9309), .ZN(n7832) );
  AOI211_X1 U9324 ( .C1(n7982), .C2(n9444), .A(n7833), .B(n7832), .ZN(n7834)
         );
  OAI21_X1 U9325 ( .B1(n9448), .B2(n9356), .A(n7834), .ZN(P1_U3277) );
  INV_X1 U9326 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10037) );
  NOR2_X1 U9327 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7835) );
  AOI21_X1 U9328 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7835), .ZN(n10009) );
  NOR2_X1 U9329 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7836) );
  AOI21_X1 U9330 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7836), .ZN(n10012) );
  NOR2_X1 U9331 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7837) );
  AOI21_X1 U9332 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7837), .ZN(n10015) );
  NOR2_X1 U9333 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7838) );
  AOI21_X1 U9334 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7838), .ZN(n10018) );
  NOR2_X1 U9335 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7839) );
  AOI21_X1 U9336 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7839), .ZN(n10021) );
  NOR2_X1 U9337 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7845) );
  XNOR2_X1 U9338 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10049) );
  NAND2_X1 U9339 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7843) );
  XOR2_X1 U9340 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10047) );
  NAND2_X1 U9341 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7841) );
  XOR2_X1 U9342 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10045) );
  AOI21_X1 U9343 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10002) );
  INV_X1 U9344 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10006) );
  NAND3_X1 U9345 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10004) );
  OAI21_X1 U9346 ( .B1(n10002), .B2(n10006), .A(n10004), .ZN(n10044) );
  NAND2_X1 U9347 ( .A1(n10045), .A2(n10044), .ZN(n7840) );
  NAND2_X1 U9348 ( .A1(n7841), .A2(n7840), .ZN(n10046) );
  NAND2_X1 U9349 ( .A1(n10047), .A2(n10046), .ZN(n7842) );
  NAND2_X1 U9350 ( .A1(n7843), .A2(n7842), .ZN(n10048) );
  NOR2_X1 U9351 ( .A1(n10049), .A2(n10048), .ZN(n7844) );
  NOR2_X1 U9352 ( .A1(n7845), .A2(n7844), .ZN(n7846) );
  NOR2_X1 U9353 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7846), .ZN(n10033) );
  AND2_X1 U9354 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7846), .ZN(n10032) );
  NOR2_X1 U9355 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10032), .ZN(n7847) );
  NOR2_X1 U9356 ( .A1(n10033), .A2(n7847), .ZN(n7848) );
  NAND2_X1 U9357 ( .A1(n7848), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7850) );
  XOR2_X1 U9358 ( .A(n7848), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10031) );
  NAND2_X1 U9359 ( .A1(n10031), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7849) );
  NAND2_X1 U9360 ( .A1(n7850), .A2(n7849), .ZN(n7851) );
  NAND2_X1 U9361 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7851), .ZN(n7853) );
  XOR2_X1 U9362 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7851), .Z(n10043) );
  NAND2_X1 U9363 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10043), .ZN(n7852) );
  NAND2_X1 U9364 ( .A1(n7853), .A2(n7852), .ZN(n7854) );
  NAND2_X1 U9365 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7854), .ZN(n7856) );
  XOR2_X1 U9366 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7854), .Z(n10042) );
  NAND2_X1 U9367 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10042), .ZN(n7855) );
  NAND2_X1 U9368 ( .A1(n7856), .A2(n7855), .ZN(n7857) );
  AND2_X1 U9369 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7857), .ZN(n7858) );
  XNOR2_X1 U9370 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7857), .ZN(n10040) );
  NOR2_X1 U9371 ( .A1(n10041), .A2(n10040), .ZN(n10039) );
  NOR2_X1 U9372 ( .A1(n7858), .A2(n10039), .ZN(n10030) );
  NAND2_X1 U9373 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7859) );
  OAI21_X1 U9374 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7859), .ZN(n10029) );
  NOR2_X1 U9375 ( .A1(n10030), .A2(n10029), .ZN(n10028) );
  AOI21_X1 U9376 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10028), .ZN(n10027) );
  NAND2_X1 U9377 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7860) );
  OAI21_X1 U9378 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7860), .ZN(n10026) );
  NOR2_X1 U9379 ( .A1(n10027), .A2(n10026), .ZN(n10025) );
  AOI21_X1 U9380 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10025), .ZN(n10024) );
  NOR2_X1 U9381 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7861) );
  AOI21_X1 U9382 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7861), .ZN(n10023) );
  NAND2_X1 U9383 ( .A1(n10024), .A2(n10023), .ZN(n10022) );
  OAI21_X1 U9384 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10022), .ZN(n10020) );
  NAND2_X1 U9385 ( .A1(n10021), .A2(n10020), .ZN(n10019) );
  OAI21_X1 U9386 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10019), .ZN(n10017) );
  NAND2_X1 U9387 ( .A1(n10018), .A2(n10017), .ZN(n10016) );
  OAI21_X1 U9388 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10016), .ZN(n10014) );
  NAND2_X1 U9389 ( .A1(n10015), .A2(n10014), .ZN(n10013) );
  OAI21_X1 U9390 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10013), .ZN(n10011) );
  NAND2_X1 U9391 ( .A1(n10012), .A2(n10011), .ZN(n10010) );
  OAI21_X1 U9392 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10010), .ZN(n10008) );
  NAND2_X1 U9393 ( .A1(n10009), .A2(n10008), .ZN(n10007) );
  OAI21_X1 U9394 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10007), .ZN(n10036) );
  NOR2_X1 U9395 ( .A1(n10037), .A2(n10036), .ZN(n7862) );
  NAND2_X1 U9396 ( .A1(n10037), .A2(n10036), .ZN(n10035) );
  OAI21_X1 U9397 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7862), .A(n10035), .ZN(
        n7864) );
  INV_X1 U9398 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8445) );
  XNOR2_X1 U9399 ( .A(n8445), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7863) );
  XNOR2_X1 U9400 ( .A(n7864), .B(n7863), .ZN(ADD_1071_U4) );
  INV_X1 U9401 ( .A(n7866), .ZN(n7867) );
  NAND2_X1 U9402 ( .A1(n7869), .A2(n7868), .ZN(n7871) );
  NAND2_X1 U9403 ( .A1(n8855), .A2(n8356), .ZN(n7870) );
  NAND2_X1 U9404 ( .A1(n7871), .A2(n7870), .ZN(n7890) );
  NAND2_X1 U9405 ( .A1(n7873), .A2(n7876), .ZN(n7874) );
  OAI22_X1 U9406 ( .A1(n8105), .A2(n8726), .B1(n8727), .B2(n8728), .ZN(n7881)
         );
  OR3_X1 U9407 ( .A1(n7877), .A2(n7876), .A3(n7875), .ZN(n7878) );
  AOI21_X1 U9408 ( .B1(n7879), .B2(n7878), .A(n8724), .ZN(n7880) );
  AOI211_X1 U9409 ( .C1(n8847), .C2(n7882), .A(n7881), .B(n7880), .ZN(n8852)
         );
  NOR2_X1 U9410 ( .A1(n7898), .A2(n8848), .ZN(n7884) );
  OR2_X1 U9411 ( .A1(n7987), .A2(n7884), .ZN(n8849) );
  AOI22_X1 U9412 ( .A1(n8742), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8103), .B2(
        n8746), .ZN(n7886) );
  NAND2_X1 U9413 ( .A1(n8753), .A2(n8108), .ZN(n7885) );
  OAI211_X1 U9414 ( .C1(n8849), .C2(n8530), .A(n7886), .B(n7885), .ZN(n7887)
         );
  AOI21_X1 U9415 ( .B1(n8847), .B2(n7888), .A(n7887), .ZN(n7889) );
  OAI21_X1 U9416 ( .B1(n8852), .B2(n8686), .A(n7889), .ZN(P2_U3283) );
  XNOR2_X1 U9417 ( .A(n7890), .B(n7895), .ZN(n9986) );
  INV_X1 U9418 ( .A(n9986), .ZN(n7907) );
  INV_X1 U9419 ( .A(n7891), .ZN(n7892) );
  NOR2_X1 U9420 ( .A1(n7893), .A2(n7892), .ZN(n7894) );
  XOR2_X1 U9421 ( .A(n7895), .B(n7894), .Z(n7896) );
  OAI222_X1 U9422 ( .A1(n8728), .A2(n7994), .B1(n8726), .B2(n7897), .C1(n8724), 
        .C2(n7896), .ZN(n9983) );
  INV_X1 U9423 ( .A(n7898), .ZN(n7899) );
  OAI21_X1 U9424 ( .B1(n4495), .B2(n7900), .A(n7899), .ZN(n9982) );
  AOI22_X1 U9425 ( .A1(n8742), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7901), .B2(
        n8746), .ZN(n7904) );
  NAND2_X1 U9426 ( .A1(n8753), .A2(n7902), .ZN(n7903) );
  OAI211_X1 U9427 ( .C1(n9982), .C2(n8530), .A(n7904), .B(n7903), .ZN(n7905)
         );
  AOI21_X1 U9428 ( .B1(n9983), .B2(n8667), .A(n7905), .ZN(n7906) );
  OAI21_X1 U9429 ( .B1(n8735), .B2(n7907), .A(n7906), .ZN(P2_U3284) );
  INV_X1 U9430 ( .A(n7908), .ZN(n7912) );
  OAI21_X1 U9431 ( .B1(n7912), .B2(n7910), .A(n7909), .ZN(n7911) );
  OAI21_X1 U9432 ( .B1(n7913), .B2(n7912), .A(n7911), .ZN(n7914) );
  NAND2_X1 U9433 ( .A1(n7914), .A2(n5630), .ZN(n7920) );
  INV_X1 U9434 ( .A(n7915), .ZN(n7918) );
  INV_X1 U9435 ( .A(n7916), .ZN(n9686) );
  OAI22_X1 U9436 ( .A1(n9008), .A2(n9686), .B1(n9035), .B2(n9690), .ZN(n7917)
         );
  AOI211_X1 U9437 ( .C1(n9020), .C2(n9044), .A(n7918), .B(n7917), .ZN(n7919)
         );
  OAI211_X1 U9438 ( .C1(n9729), .C2(n7921), .A(n7920), .B(n7919), .ZN(P1_U3232) );
  NOR2_X1 U9439 ( .A1(n7922), .A2(n7929), .ZN(n7924) );
  NAND2_X1 U9440 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9078), .ZN(n7925) );
  OAI21_X1 U9441 ( .B1(n9078), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7925), .ZN(
        n7926) );
  NOR2_X1 U9442 ( .A1(n7927), .A2(n7926), .ZN(n9077) );
  AOI211_X1 U9443 ( .C1(n7927), .C2(n7926), .A(n9077), .B(n9817), .ZN(n7938)
         );
  NOR2_X1 U9444 ( .A1(n7929), .A2(n7928), .ZN(n7931) );
  NOR2_X1 U9445 ( .A1(n7931), .A2(n7930), .ZN(n7933) );
  XNOR2_X1 U9446 ( .A(n9078), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7932) );
  NOR2_X1 U9447 ( .A1(n7933), .A2(n7932), .ZN(n9071) );
  AOI211_X1 U9448 ( .C1(n7933), .C2(n7932), .A(n9071), .B(n9072), .ZN(n7937)
         );
  INV_X1 U9449 ( .A(n9078), .ZN(n7935) );
  NAND2_X1 U9450 ( .A1(n9827), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7934) );
  NAND2_X1 U9451 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8952) );
  OAI211_X1 U9452 ( .C1(n9060), .C2(n7935), .A(n7934), .B(n8952), .ZN(n7936)
         );
  OR3_X1 U9453 ( .A1(n7938), .A2(n7937), .A3(n7936), .ZN(P1_U3257) );
  INV_X1 U9454 ( .A(n7939), .ZN(n7946) );
  AOI22_X1 U9455 ( .A1(n7940), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n9647), .ZN(n7941) );
  OAI21_X1 U9456 ( .B1(n7946), .B2(n9653), .A(n7941), .ZN(P1_U3328) );
  INV_X1 U9457 ( .A(n7942), .ZN(n7949) );
  AOI22_X1 U9458 ( .A1(n7943), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n9650), .ZN(n7944) );
  OAI21_X1 U9459 ( .B1(n7949), .B2(n9653), .A(n7944), .ZN(P1_U3327) );
  OAI222_X1 U9460 ( .A1(n8197), .A2(n7947), .B1(n8195), .B2(n7946), .C1(
        P2_U3152), .C2(n7945), .ZN(P2_U3333) );
  OAI222_X1 U9461 ( .A1(P2_U3152), .A2(n7950), .B1(n8195), .B2(n7949), .C1(
        n7948), .C2(n8197), .ZN(P2_U3332) );
  OAI21_X1 U9462 ( .B1(n7955), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7951), .ZN(
        n8378) );
  XNOR2_X1 U9463 ( .A(n8378), .B(n8379), .ZN(n7954) );
  INV_X1 U9464 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7953) );
  NOR2_X1 U9465 ( .A1(n7953), .A2(n7954), .ZN(n8380) );
  AOI211_X1 U9466 ( .C1(n7954), .C2(n7953), .A(n8380), .B(n7952), .ZN(n7963)
         );
  NOR2_X1 U9467 ( .A1(n7955), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7957) );
  NOR2_X1 U9468 ( .A1(n7957), .A2(n7956), .ZN(n8389) );
  XNOR2_X1 U9469 ( .A(n8389), .B(n8390), .ZN(n7958) );
  NOR2_X1 U9470 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7958), .ZN(n8391) );
  AOI21_X1 U9471 ( .B1(n7958), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8391), .ZN(
        n7959) );
  NOR2_X1 U9472 ( .A1(n7959), .A2(n9917), .ZN(n7962) );
  NOR2_X1 U9473 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5883), .ZN(n8344) );
  AOI21_X1 U9474 ( .B1(n9920), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8344), .ZN(
        n7960) );
  OAI21_X1 U9475 ( .B1(n9915), .B2(n8379), .A(n7960), .ZN(n7961) );
  OR3_X1 U9476 ( .A1(n7963), .A2(n7962), .A3(n7961), .ZN(P2_U3260) );
  INV_X1 U9477 ( .A(n7964), .ZN(n7968) );
  AOI21_X1 U9478 ( .B1(n9647), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7965), .ZN(
        n7966) );
  OAI21_X1 U9479 ( .B1(n7968), .B2(n9653), .A(n7966), .ZN(P1_U3326) );
  AOI22_X1 U9480 ( .A1(n8449), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n8889), .ZN(n7967) );
  OAI21_X1 U9481 ( .B1(n7968), .B2(n8195), .A(n7967), .ZN(P2_U3331) );
  NAND2_X1 U9482 ( .A1(n8006), .A2(n7970), .ZN(n9143) );
  XNOR2_X1 U9483 ( .A(n9143), .B(n9142), .ZN(n7971) );
  INV_X1 U9484 ( .A(n7976), .ZN(n9042) );
  AOI222_X1 U9485 ( .A1(n9352), .A2(n7971), .B1(n9333), .B2(n9349), .C1(n9042), 
        .C2(n9347), .ZN(n9437) );
  INV_X1 U9486 ( .A(n7972), .ZN(n7975) );
  AOI21_X1 U9487 ( .B1(n7975), .B2(n4818), .A(n4817), .ZN(n8009) );
  NAND2_X1 U9488 ( .A1(n8009), .A2(n4827), .ZN(n7978) );
  NAND2_X1 U9489 ( .A1(n7978), .A2(n7977), .ZN(n7979) );
  NAND2_X1 U9490 ( .A1(n7979), .A2(n9142), .ZN(n9433) );
  NAND3_X1 U9491 ( .A1(n4597), .A2(n7270), .A3(n9433), .ZN(n7985) );
  OAI211_X1 U9492 ( .C1(n4361), .C2(n8950), .A(n9888), .B(n9342), .ZN(n9435)
         );
  INV_X1 U9493 ( .A(n9435), .ZN(n7983) );
  AOI22_X1 U9494 ( .A1(n9309), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n8951), .B2(
        n9720), .ZN(n7980) );
  OAI21_X1 U9495 ( .B1(n8950), .B2(n9723), .A(n7980), .ZN(n7981) );
  AOI21_X1 U9496 ( .B1(n7983), .B2(n7982), .A(n7981), .ZN(n7984) );
  OAI211_X1 U9497 ( .C1(n9309), .C2(n9437), .A(n7985), .B(n7984), .ZN(P1_U3275) );
  XNOR2_X1 U9498 ( .A(n8460), .B(n7993), .ZN(n8846) );
  INV_X1 U9499 ( .A(n7987), .ZN(n7988) );
  INV_X1 U9500 ( .A(n8842), .ZN(n7990) );
  AOI21_X1 U9501 ( .B1(n8842), .B2(n7988), .A(n4496), .ZN(n8843) );
  AOI22_X1 U9502 ( .A1(n8742), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8095), .B2(
        n8746), .ZN(n7989) );
  OAI21_X1 U9503 ( .B1(n7990), .B2(n8721), .A(n7989), .ZN(n7998) );
  AOI211_X1 U9504 ( .C1(n7993), .C2(n7992), .A(n8724), .B(n7991), .ZN(n7996)
         );
  OAI22_X1 U9505 ( .A1(n7994), .A2(n8726), .B1(n8273), .B2(n8728), .ZN(n7995)
         );
  NOR2_X1 U9506 ( .A1(n7996), .A2(n7995), .ZN(n8845) );
  NOR2_X1 U9507 ( .A1(n8845), .A2(n8686), .ZN(n7997) );
  AOI211_X1 U9508 ( .C1(n8843), .C2(n8748), .A(n7998), .B(n7997), .ZN(n7999)
         );
  OAI21_X1 U9509 ( .B1(n8735), .B2(n8846), .A(n7999), .ZN(P2_U3282) );
  INV_X1 U9510 ( .A(n8000), .ZN(n8005) );
  AOI22_X1 U9511 ( .A1(n8001), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n8889), .ZN(n8002) );
  OAI21_X1 U9512 ( .B1(n8005), .B2(n8195), .A(n8002), .ZN(P2_U3330) );
  NAND2_X1 U9513 ( .A1(n9650), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8003) );
  OAI211_X1 U9514 ( .C1(n8005), .C2(n9653), .A(n8004), .B(n8003), .ZN(P1_U3325) );
  OAI21_X1 U9515 ( .B1(n8008), .B2(n8007), .A(n8006), .ZN(n8012) );
  OAI22_X1 U9516 ( .A1(n8033), .A2(n9710), .B1(n9690), .B2(n9712), .ZN(n8011)
         );
  XNOR2_X1 U9517 ( .A(n8009), .B(n8008), .ZN(n9443) );
  INV_X1 U9518 ( .A(n9719), .ZN(n9881) );
  NOR2_X1 U9519 ( .A1(n9443), .A2(n9881), .ZN(n8010) );
  AOI211_X1 U9520 ( .C1(n9352), .C2(n8012), .A(n8011), .B(n8010), .ZN(n9442)
         );
  INV_X1 U9521 ( .A(n8013), .ZN(n8014) );
  AOI21_X1 U9522 ( .B1(n9439), .B2(n8014), .A(n4361), .ZN(n9440) );
  AOI22_X1 U9523 ( .A1(n9309), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n4830), .B2(
        n9720), .ZN(n8015) );
  OAI21_X1 U9524 ( .B1(n8016), .B2(n9723), .A(n8015), .ZN(n8019) );
  NOR2_X1 U9525 ( .A1(n9443), .A2(n8017), .ZN(n8018) );
  AOI211_X1 U9526 ( .C1(n9440), .C2(n9706), .A(n8019), .B(n8018), .ZN(n8020)
         );
  OAI21_X1 U9527 ( .B1(n9442), .B2(n9309), .A(n8020), .ZN(P1_U3276) );
  INV_X1 U9528 ( .A(n8021), .ZN(n8026) );
  AOI22_X1 U9529 ( .A1(n8022), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n8889), .ZN(n8023) );
  OAI21_X1 U9530 ( .B1(n8026), .B2(n8195), .A(n8023), .ZN(P2_U3329) );
  AOI22_X1 U9531 ( .A1(n8024), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9650), .ZN(n8025) );
  OAI21_X1 U9532 ( .B1(n8026), .B2(n9653), .A(n8025), .ZN(P1_U3324) );
  NAND2_X1 U9533 ( .A1(n8028), .A2(n8027), .ZN(n8029) );
  XOR2_X1 U9534 ( .A(n8030), .B(n8029), .Z(n8036) );
  AOI22_X1 U9535 ( .A1(n9020), .A2(n7974), .B1(n4830), .B2(n9033), .ZN(n8032)
         );
  OAI211_X1 U9536 ( .C1(n8033), .C2(n9035), .A(n8032), .B(n8031), .ZN(n8034)
         );
  AOI21_X1 U9537 ( .B1(n9439), .B2(n9038), .A(n8034), .ZN(n8035) );
  OAI21_X1 U9538 ( .B1(n8036), .B2(n9012), .A(n8035), .ZN(P1_U3239) );
  AOI22_X1 U9539 ( .A1(n9022), .A2(n9042), .B1(n9033), .B2(n8037), .ZN(n8039)
         );
  OAI211_X1 U9540 ( .C1(n8040), .C2(n9032), .A(n8039), .B(n8038), .ZN(n8048)
         );
  INV_X1 U9541 ( .A(n8041), .ZN(n8046) );
  AOI21_X1 U9542 ( .B1(n8045), .B2(n8043), .A(n8042), .ZN(n8044) );
  AOI211_X1 U9543 ( .C1(n8046), .C2(n8045), .A(n9012), .B(n8044), .ZN(n8047)
         );
  AOI211_X1 U9544 ( .C1(n9038), .C2(n9445), .A(n8048), .B(n8047), .ZN(n8049)
         );
  INV_X1 U9545 ( .A(n8049), .ZN(P1_U3213) );
  AOI22_X1 U9546 ( .A1(n8345), .A2(n7009), .B1(n8346), .B2(n8050), .ZN(n8057)
         );
  OAI21_X1 U9547 ( .B1(n8053), .B2(n8052), .A(n8051), .ZN(n8054) );
  AOI22_X1 U9548 ( .A1(n8055), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n8325), .B2(
        n8054), .ZN(n8056) );
  OAI211_X1 U9549 ( .C1(n8342), .C2(n8058), .A(n8057), .B(n8056), .ZN(P2_U3224) );
  NAND2_X1 U9550 ( .A1(n4379), .A2(n8059), .ZN(n8060) );
  XNOR2_X1 U9551 ( .A(n8061), .B(n8060), .ZN(n8067) );
  AOI22_X1 U9552 ( .A1(n9020), .A2(n9047), .B1(n8062), .B2(n9033), .ZN(n8063)
         );
  NAND2_X1 U9553 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3084), .ZN(n9816) );
  OAI211_X1 U9554 ( .C1(n8064), .C2(n9035), .A(n8063), .B(n9816), .ZN(n8065)
         );
  AOI21_X1 U9555 ( .B1(n9038), .B2(n9671), .A(n8065), .ZN(n8066) );
  OAI21_X1 U9556 ( .B1(n8067), .B2(n9012), .A(n8066), .ZN(P1_U3215) );
  XOR2_X1 U9557 ( .A(n8074), .B(n8068), .Z(n9893) );
  INV_X1 U9558 ( .A(n8069), .ZN(n8070) );
  AOI21_X1 U9559 ( .B1(n9886), .B2(n8071), .A(n8070), .ZN(n9889) );
  AOI22_X1 U9560 ( .A1(n9309), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n8072), .B2(
        n9720), .ZN(n8073) );
  OAI21_X1 U9561 ( .B1(n4671), .B2(n9723), .A(n8073), .ZN(n8080) );
  XNOR2_X1 U9562 ( .A(n8075), .B(n8074), .ZN(n8078) );
  OAI22_X1 U9563 ( .A1(n8076), .A2(n9712), .B1(n9713), .B2(n9710), .ZN(n8077)
         );
  AOI21_X1 U9564 ( .B1(n8078), .B2(n9352), .A(n8077), .ZN(n9891) );
  NOR2_X1 U9565 ( .A1(n9891), .A2(n9309), .ZN(n8079) );
  AOI211_X1 U9566 ( .C1(n9889), .C2(n9706), .A(n8080), .B(n8079), .ZN(n8081)
         );
  OAI21_X1 U9567 ( .B1(n9893), .B2(n9356), .A(n8081), .ZN(P1_U3282) );
  XNOR2_X1 U9568 ( .A(n8842), .B(n8168), .ZN(n8082) );
  NAND2_X1 U9569 ( .A1(n8458), .A2(n8154), .ZN(n8083) );
  NAND2_X1 U9570 ( .A1(n8082), .A2(n8083), .ZN(n8116) );
  INV_X1 U9571 ( .A(n8082), .ZN(n8085) );
  INV_X1 U9572 ( .A(n8083), .ZN(n8084) );
  NAND2_X1 U9573 ( .A1(n8085), .A2(n8084), .ZN(n8086) );
  NAND2_X1 U9574 ( .A1(n8116), .A2(n8086), .ZN(n8094) );
  AND2_X1 U9575 ( .A1(n8088), .A2(n8087), .ZN(n8089) );
  NAND2_X1 U9576 ( .A1(n8090), .A2(n8089), .ZN(n8101) );
  XNOR2_X1 U9577 ( .A(n8108), .B(n8168), .ZN(n8092) );
  NAND2_X1 U9578 ( .A1(n8354), .A2(n8154), .ZN(n8091) );
  XNOR2_X1 U9579 ( .A(n8092), .B(n8091), .ZN(n8102) );
  AOI21_X1 U9580 ( .B1(n8094), .B2(n8093), .A(n4366), .ZN(n8100) );
  AOI22_X1 U9581 ( .A1(n8240), .A2(n8354), .B1(n8333), .B2(n8095), .ZN(n8097)
         );
  OAI211_X1 U9582 ( .C1(n8273), .C2(n8314), .A(n8097), .B(n8096), .ZN(n8098)
         );
  AOI21_X1 U9583 ( .B1(n8346), .B2(n8842), .A(n8098), .ZN(n8099) );
  OAI21_X1 U9584 ( .B1(n8100), .B2(n8349), .A(n8099), .ZN(P2_U3217) );
  XNOR2_X1 U9585 ( .A(n8101), .B(n8102), .ZN(n8110) );
  OAI22_X1 U9586 ( .A1(n8314), .A2(n8727), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7567), .ZN(n8107) );
  INV_X1 U9587 ( .A(n8103), .ZN(n8104) );
  OAI22_X1 U9588 ( .A1(n8342), .A2(n8105), .B1(n8341), .B2(n8104), .ZN(n8106)
         );
  AOI211_X1 U9589 ( .C1(n8346), .C2(n8108), .A(n8107), .B(n8106), .ZN(n8109)
         );
  OAI21_X1 U9590 ( .B1(n8110), .B2(n8349), .A(n8109), .ZN(P2_U3236) );
  INV_X1 U9591 ( .A(n9423), .ZN(n9328) );
  INV_X1 U9592 ( .A(n9419), .ZN(n9123) );
  NAND2_X1 U9593 ( .A1(n9323), .A2(n9123), .ZN(n9314) );
  OR2_X2 U9594 ( .A1(n9213), .A2(n9379), .ZN(n9192) );
  INV_X1 U9595 ( .A(P1_B_REG_SCAN_IN), .ZN(n8111) );
  NOR2_X1 U9596 ( .A1(n6565), .A2(n8111), .ZN(n8112) );
  NOR2_X1 U9597 ( .A1(n9710), .A2(n8112), .ZN(n9164) );
  NAND2_X1 U9598 ( .A1(n8113), .A2(n9164), .ZN(n9362) );
  NOR2_X1 U9599 ( .A1(n9309), .A2(n9362), .ZN(n9115) );
  INV_X1 U9600 ( .A(n9360), .ZN(n9113) );
  NOR2_X1 U9601 ( .A1(n9113), .A2(n9723), .ZN(n8114) );
  AOI211_X1 U9602 ( .C1(n9309), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9115), .B(
        n8114), .ZN(n8115) );
  OAI21_X1 U9603 ( .B1(n9363), .B2(n9118), .A(n8115), .ZN(P1_U3262) );
  NAND2_X1 U9604 ( .A1(n8617), .A2(n8154), .ZN(n8289) );
  XNOR2_X1 U9605 ( .A(n8837), .B(n8168), .ZN(n8265) );
  NAND2_X1 U9606 ( .A1(n8461), .A2(n8154), .ZN(n8117) );
  XNOR2_X1 U9607 ( .A(n8832), .B(n8175), .ZN(n8122) );
  NAND2_X1 U9608 ( .A1(n8463), .A2(n8154), .ZN(n8123) );
  XNOR2_X1 U9609 ( .A(n8122), .B(n8123), .ZN(n8267) );
  INV_X1 U9610 ( .A(n8265), .ZN(n8118) );
  INV_X1 U9611 ( .A(n8117), .ZN(n8339) );
  NAND2_X1 U9612 ( .A1(n8118), .A2(n8339), .ZN(n8119) );
  AND2_X1 U9613 ( .A1(n8267), .A2(n8119), .ZN(n8120) );
  NAND2_X1 U9614 ( .A1(n8121), .A2(n8120), .ZN(n8269) );
  INV_X1 U9615 ( .A(n8122), .ZN(n8124) );
  NAND2_X1 U9616 ( .A1(n8124), .A2(n8123), .ZN(n8125) );
  NAND2_X1 U9617 ( .A1(n8269), .A2(n8125), .ZN(n8279) );
  XNOR2_X1 U9618 ( .A(n8828), .B(n8168), .ZN(n8126) );
  NAND2_X1 U9619 ( .A1(n8465), .A2(n8154), .ZN(n8127) );
  XNOR2_X1 U9620 ( .A(n8126), .B(n8127), .ZN(n8278) );
  INV_X1 U9621 ( .A(n8126), .ZN(n8129) );
  INV_X1 U9622 ( .A(n8127), .ZN(n8128) );
  NAND2_X1 U9623 ( .A1(n8129), .A2(n8128), .ZN(n8130) );
  XNOR2_X1 U9624 ( .A(n8824), .B(n8175), .ZN(n8133) );
  NAND2_X1 U9625 ( .A1(n8468), .A2(n8154), .ZN(n8131) );
  XNOR2_X1 U9626 ( .A(n8133), .B(n8131), .ZN(n8319) );
  INV_X1 U9627 ( .A(n8131), .ZN(n8132) );
  AND2_X1 U9628 ( .A1(n8133), .A2(n8132), .ZN(n8134) );
  XNOR2_X1 U9629 ( .A(n8818), .B(n8168), .ZN(n8135) );
  NAND2_X1 U9630 ( .A1(n8471), .A2(n8154), .ZN(n8136) );
  NAND2_X1 U9631 ( .A1(n8135), .A2(n8136), .ZN(n8140) );
  INV_X1 U9632 ( .A(n8135), .ZN(n8138) );
  INV_X1 U9633 ( .A(n8136), .ZN(n8137) );
  NAND2_X1 U9634 ( .A1(n8138), .A2(n8137), .ZN(n8139) );
  AND2_X1 U9635 ( .A1(n8140), .A2(n8139), .ZN(n8226) );
  NAND2_X1 U9636 ( .A1(n8225), .A2(n8140), .ZN(n8302) );
  XNOR2_X1 U9637 ( .A(n8812), .B(n8168), .ZN(n8141) );
  NAND2_X1 U9638 ( .A1(n8631), .A2(n8154), .ZN(n8142) );
  XNOR2_X1 U9639 ( .A(n8141), .B(n8142), .ZN(n8301) );
  INV_X1 U9640 ( .A(n8141), .ZN(n8144) );
  INV_X1 U9641 ( .A(n8142), .ZN(n8143) );
  NAND2_X1 U9642 ( .A1(n8144), .A2(n8143), .ZN(n8145) );
  XNOR2_X1 U9643 ( .A(n8807), .B(n8175), .ZN(n8148) );
  NAND2_X1 U9644 ( .A1(n8616), .A2(n8154), .ZN(n8146) );
  XNOR2_X1 U9645 ( .A(n8148), .B(n8146), .ZN(n8247) );
  INV_X1 U9646 ( .A(n8146), .ZN(n8147) );
  XNOR2_X1 U9647 ( .A(n8802), .B(n8168), .ZN(n8149) );
  XNOR2_X1 U9648 ( .A(n8151), .B(n8149), .ZN(n8311) );
  NAND2_X1 U9649 ( .A1(n8476), .A2(n8154), .ZN(n8310) );
  NAND2_X1 U9650 ( .A1(n8311), .A2(n8310), .ZN(n8309) );
  INV_X1 U9651 ( .A(n8149), .ZN(n8150) );
  NAND2_X1 U9652 ( .A1(n8309), .A2(n8152), .ZN(n8153) );
  XNOR2_X1 U9653 ( .A(n8153), .B(n4359), .ZN(n8206) );
  NAND2_X1 U9654 ( .A1(n4539), .A2(n8154), .ZN(n8157) );
  INV_X1 U9655 ( .A(n8291), .ZN(n8158) );
  INV_X1 U9656 ( .A(n8157), .ZN(n8290) );
  OR2_X2 U9657 ( .A1(n8162), .A2(n8161), .ZN(n8163) );
  XNOR2_X1 U9658 ( .A(n8788), .B(n8175), .ZN(n8164) );
  NAND2_X1 U9659 ( .A1(n8580), .A2(n8154), .ZN(n8255) );
  INV_X1 U9660 ( .A(n8164), .ZN(n8256) );
  XNOR2_X1 U9661 ( .A(n8784), .B(n8168), .ZN(n8166) );
  OR2_X1 U9662 ( .A1(n8352), .A2(n8174), .ZN(n8165) );
  NOR2_X1 U9663 ( .A1(n8166), .A2(n8165), .ZN(n8167) );
  AOI21_X1 U9664 ( .B1(n8166), .B2(n8165), .A(n8167), .ZN(n8327) );
  INV_X1 U9665 ( .A(n8167), .ZN(n8198) );
  XNOR2_X1 U9666 ( .A(n8776), .B(n8168), .ZN(n8173) );
  NAND2_X1 U9667 ( .A1(n8485), .A2(n8154), .ZN(n8172) );
  NOR2_X1 U9668 ( .A1(n8173), .A2(n8172), .ZN(n8171) );
  INV_X1 U9669 ( .A(n8171), .ZN(n8170) );
  AND2_X1 U9670 ( .A1(n8198), .A2(n8170), .ZN(n8169) );
  AOI21_X1 U9671 ( .B1(n8173), .B2(n8172), .A(n8171), .ZN(n8200) );
  OR2_X1 U9672 ( .A1(n8171), .A2(n8200), .ZN(n8181) );
  AND2_X1 U9673 ( .A1(n8183), .A2(n8181), .ZN(n8187) );
  NOR2_X1 U9674 ( .A1(n8511), .A2(n8856), .ZN(n8179) );
  INV_X1 U9675 ( .A(n8179), .ZN(n8177) );
  NOR2_X1 U9676 ( .A1(n8488), .A2(n8174), .ZN(n8176) );
  XNOR2_X1 U9677 ( .A(n8176), .B(n8175), .ZN(n8178) );
  MUX2_X1 U9678 ( .A(n8770), .B(n8177), .S(n8178), .Z(n8186) );
  MUX2_X1 U9679 ( .A(n8179), .B(n8511), .S(n8178), .Z(n8180) );
  AND2_X1 U9680 ( .A1(n8181), .A2(n8180), .ZN(n8182) );
  NAND2_X1 U9681 ( .A1(n8183), .A2(n8182), .ZN(n8185) );
  OAI21_X1 U9682 ( .B1(n8511), .B2(n8336), .A(n8349), .ZN(n8184) );
  OAI211_X1 U9683 ( .C1(n8187), .C2(n8186), .A(n8185), .B(n8184), .ZN(n8192)
         );
  INV_X1 U9684 ( .A(n8517), .ZN(n8351) );
  INV_X1 U9685 ( .A(n8188), .ZN(n8509) );
  AOI22_X1 U9686 ( .A1(n8345), .A2(n8351), .B1(n8333), .B2(n8509), .ZN(n8190)
         );
  AOI22_X1 U9687 ( .A1(n8240), .A2(n8485), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8189) );
  AND2_X1 U9688 ( .A1(n8190), .A2(n8189), .ZN(n8191) );
  NAND2_X1 U9689 ( .A1(n8192), .A2(n8191), .ZN(P2_U3222) );
  OAI222_X1 U9690 ( .A1(n8197), .A2(n8196), .B1(n8195), .B2(n8194), .C1(
        P2_U3152), .C2(n8193), .ZN(P2_U3336) );
  NAND2_X1 U9691 ( .A1(n8326), .A2(n8198), .ZN(n8201) );
  NAND2_X1 U9692 ( .A1(n8201), .A2(n8200), .ZN(n8199) );
  OAI211_X1 U9693 ( .C1(n8201), .C2(n8200), .A(n8199), .B(n8325), .ZN(n8205)
         );
  OAI22_X1 U9694 ( .A1(n8488), .A2(n8728), .B1(n8352), .B2(n8726), .ZN(n8526)
         );
  AOI22_X1 U9695 ( .A1(n8526), .A2(n8282), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8202) );
  OAI21_X1 U9696 ( .B1(n8532), .B2(n8341), .A(n8202), .ZN(n8203) );
  AOI21_X1 U9697 ( .B1(n8776), .B2(n8346), .A(n8203), .ZN(n8204) );
  NAND2_X1 U9698 ( .A1(n8205), .A2(n8204), .ZN(P2_U3216) );
  XNOR2_X1 U9699 ( .A(n8206), .B(n8289), .ZN(n8212) );
  OR2_X1 U9700 ( .A1(n8480), .A2(n8728), .ZN(n8208) );
  NAND2_X1 U9701 ( .A1(n8476), .A2(n8630), .ZN(n8207) );
  NAND2_X1 U9702 ( .A1(n8208), .A2(n8207), .ZN(n8599) );
  AOI22_X1 U9703 ( .A1(n8282), .A2(n8599), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8209) );
  OAI21_X1 U9704 ( .B1(n8341), .B2(n8590), .A(n8209), .ZN(n8210) );
  AOI21_X1 U9705 ( .B1(n8797), .B2(n8346), .A(n8210), .ZN(n8211) );
  OAI21_X1 U9706 ( .B1(n8212), .B2(n8349), .A(n8211), .ZN(P2_U3218) );
  NAND2_X1 U9707 ( .A1(n8214), .A2(n8213), .ZN(n8215) );
  XOR2_X1 U9708 ( .A(n8216), .B(n8215), .Z(n8217) );
  NAND2_X1 U9709 ( .A1(n8217), .A2(n8325), .ZN(n8224) );
  AOI22_X1 U9710 ( .A1(n8240), .A2(n8358), .B1(n8346), .B2(n8218), .ZN(n8223)
         );
  AOI21_X1 U9711 ( .B1(n8345), .B2(n8356), .A(n8219), .ZN(n8222) );
  NAND2_X1 U9712 ( .A1(n8333), .A2(n8220), .ZN(n8221) );
  NAND4_X1 U9713 ( .A1(n8224), .A2(n8223), .A3(n8222), .A4(n8221), .ZN(
        P2_U3219) );
  INV_X1 U9714 ( .A(n8818), .ZN(n8655) );
  OAI21_X1 U9715 ( .B1(n8227), .B2(n8226), .A(n8225), .ZN(n8228) );
  NAND2_X1 U9716 ( .A1(n8228), .A2(n8325), .ZN(n8235) );
  INV_X1 U9717 ( .A(n8282), .ZN(n8331) );
  NAND2_X1 U9718 ( .A1(n8468), .A2(n8630), .ZN(n8230) );
  NAND2_X1 U9719 ( .A1(n8631), .A2(n8632), .ZN(n8229) );
  NAND2_X1 U9720 ( .A1(n8230), .A2(n8229), .ZN(n8658) );
  INV_X1 U9721 ( .A(n8658), .ZN(n8232) );
  OAI22_X1 U9722 ( .A1(n8331), .A2(n8232), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8231), .ZN(n8233) );
  AOI21_X1 U9723 ( .B1(n8653), .B2(n8333), .A(n8233), .ZN(n8234) );
  OAI211_X1 U9724 ( .C1(n8655), .C2(n8336), .A(n8235), .B(n8234), .ZN(P2_U3221) );
  XOR2_X1 U9725 ( .A(n8237), .B(n8236), .Z(n8238) );
  NAND2_X1 U9726 ( .A1(n8238), .A2(n8325), .ZN(n8246) );
  AOI22_X1 U9727 ( .A1(n8240), .A2(n8360), .B1(n8346), .B2(n8239), .ZN(n8245)
         );
  AOI21_X1 U9728 ( .B1(n8345), .B2(n8358), .A(n8241), .ZN(n8244) );
  NAND2_X1 U9729 ( .A1(n8333), .A2(n8242), .ZN(n8243) );
  NAND4_X1 U9730 ( .A1(n8246), .A2(n8245), .A3(n8244), .A4(n8243), .ZN(
        P2_U3223) );
  XNOR2_X1 U9731 ( .A(n8248), .B(n8247), .ZN(n8254) );
  OAI22_X1 U9732 ( .A1(n8314), .A2(n8475), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8249), .ZN(n8252) );
  OAI22_X1 U9733 ( .A1(n8342), .A2(n8250), .B1(n8341), .B2(n8624), .ZN(n8251)
         );
  AOI211_X1 U9734 ( .C1(n8807), .C2(n8346), .A(n8252), .B(n8251), .ZN(n8253)
         );
  OAI21_X1 U9735 ( .B1(n8254), .B2(n8349), .A(n8253), .ZN(P2_U3225) );
  XNOR2_X1 U9736 ( .A(n8256), .B(n8255), .ZN(n8257) );
  XNOR2_X1 U9737 ( .A(n8258), .B(n8257), .ZN(n8264) );
  OR2_X1 U9738 ( .A1(n8352), .A2(n8728), .ZN(n8260) );
  OR2_X1 U9739 ( .A1(n8480), .A2(n8726), .ZN(n8259) );
  NAND2_X1 U9740 ( .A1(n8260), .A2(n8259), .ZN(n8569) );
  AOI22_X1 U9741 ( .A1(n8282), .A2(n8569), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8261) );
  OAI21_X1 U9742 ( .B1(n8341), .B2(n8561), .A(n8261), .ZN(n8262) );
  AOI21_X1 U9743 ( .B1(n8788), .B2(n8346), .A(n8262), .ZN(n8263) );
  OAI21_X1 U9744 ( .B1(n8264), .B2(n8349), .A(n8263), .ZN(P2_U3227) );
  INV_X1 U9745 ( .A(n8832), .ZN(n8704) );
  NAND2_X1 U9746 ( .A1(n4360), .A2(n8265), .ZN(n8266) );
  OAI21_X1 U9747 ( .B1(n4360), .B2(n8265), .A(n8266), .ZN(n8338) );
  NOR2_X1 U9748 ( .A1(n8338), .A2(n8339), .ZN(n8337) );
  INV_X1 U9749 ( .A(n8266), .ZN(n8268) );
  NOR3_X1 U9750 ( .A1(n8337), .A2(n8268), .A3(n8267), .ZN(n8271) );
  INV_X1 U9751 ( .A(n8269), .ZN(n8270) );
  OAI21_X1 U9752 ( .B1(n8271), .B2(n8270), .A(n8325), .ZN(n8277) );
  OAI22_X1 U9753 ( .A1(n8273), .A2(n8726), .B1(n8272), .B2(n8728), .ZN(n8709)
         );
  INV_X1 U9754 ( .A(n8709), .ZN(n8274) );
  NAND2_X1 U9755 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8385) );
  OAI21_X1 U9756 ( .B1(n8331), .B2(n8274), .A(n8385), .ZN(n8275) );
  AOI21_X1 U9757 ( .B1(n8702), .B2(n8333), .A(n8275), .ZN(n8276) );
  OAI211_X1 U9758 ( .C1(n8704), .C2(n8336), .A(n8277), .B(n8276), .ZN(P2_U3228) );
  XNOR2_X1 U9759 ( .A(n8279), .B(n8278), .ZN(n8287) );
  INV_X1 U9760 ( .A(n8685), .ZN(n8284) );
  NAND2_X1 U9761 ( .A1(n8463), .A2(n8630), .ZN(n8281) );
  NAND2_X1 U9762 ( .A1(n8468), .A2(n8632), .ZN(n8280) );
  NAND2_X1 U9763 ( .A1(n8281), .A2(n8280), .ZN(n8691) );
  AOI22_X1 U9764 ( .A1(n8282), .A2(n8691), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n8283) );
  OAI21_X1 U9765 ( .B1(n8341), .B2(n8284), .A(n8283), .ZN(n8285) );
  AOI21_X1 U9766 ( .B1(n8828), .B2(n8346), .A(n8285), .ZN(n8286) );
  OAI21_X1 U9767 ( .B1(n8287), .B2(n8349), .A(n8286), .ZN(P2_U3230) );
  OAI21_X1 U9768 ( .B1(n8206), .B2(n8289), .A(n8288), .ZN(n8293) );
  XNOR2_X1 U9769 ( .A(n8291), .B(n8290), .ZN(n8292) );
  XNOR2_X1 U9770 ( .A(n8293), .B(n8292), .ZN(n8300) );
  OAI22_X1 U9771 ( .A1(n8314), .A2(n8295), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8294), .ZN(n8298) );
  INV_X1 U9772 ( .A(n8576), .ZN(n8296) );
  OAI22_X1 U9773 ( .A1(n8342), .A2(n8479), .B1(n8341), .B2(n8296), .ZN(n8297)
         );
  AOI211_X1 U9774 ( .C1(n8792), .C2(n8346), .A(n8298), .B(n8297), .ZN(n8299)
         );
  OAI21_X1 U9775 ( .B1(n8300), .B2(n8349), .A(n8299), .ZN(P2_U3231) );
  XNOR2_X1 U9776 ( .A(n8302), .B(n8301), .ZN(n8308) );
  OAI22_X1 U9777 ( .A1(n8314), .A2(n8645), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8303), .ZN(n8306) );
  INV_X1 U9778 ( .A(n8639), .ZN(n8304) );
  OAI22_X1 U9779 ( .A1(n8342), .A2(n8644), .B1(n8341), .B2(n8304), .ZN(n8305)
         );
  AOI211_X1 U9780 ( .C1(n8812), .C2(n8346), .A(n8306), .B(n8305), .ZN(n8307)
         );
  OAI21_X1 U9781 ( .B1(n8308), .B2(n8349), .A(n8307), .ZN(P2_U3235) );
  OAI21_X1 U9782 ( .B1(n8311), .B2(n8310), .A(n8309), .ZN(n8312) );
  NAND2_X1 U9783 ( .A1(n8312), .A2(n8325), .ZN(n8318) );
  OAI22_X1 U9784 ( .A1(n8314), .A2(n8479), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8313), .ZN(n8316) );
  OAI22_X1 U9785 ( .A1(n8342), .A2(n8645), .B1(n8341), .B2(n8609), .ZN(n8315)
         );
  AOI211_X1 U9786 ( .C1(n8802), .C2(n8346), .A(n8316), .B(n8315), .ZN(n8317)
         );
  NAND2_X1 U9787 ( .A1(n8318), .A2(n8317), .ZN(P2_U3237) );
  XNOR2_X1 U9788 ( .A(n8320), .B(n8319), .ZN(n8324) );
  AOI22_X1 U9789 ( .A1(n8630), .A2(n8465), .B1(n8471), .B2(n8632), .ZN(n8673)
         );
  NAND2_X1 U9790 ( .A1(n8333), .A2(n8675), .ZN(n8321) );
  NAND2_X1 U9791 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8424) );
  OAI211_X1 U9792 ( .C1(n8331), .C2(n8673), .A(n8321), .B(n8424), .ZN(n8322)
         );
  AOI21_X1 U9793 ( .B1(n8824), .B2(n8346), .A(n8322), .ZN(n8323) );
  OAI21_X1 U9794 ( .B1(n8324), .B2(n8349), .A(n8323), .ZN(P2_U3240) );
  INV_X1 U9795 ( .A(n8784), .ZN(n8447) );
  OAI211_X1 U9796 ( .C1(n8328), .C2(n8327), .A(n8326), .B(n8325), .ZN(n8335)
         );
  AND2_X1 U9797 ( .A1(n8580), .A2(n8630), .ZN(n8329) );
  AOI21_X1 U9798 ( .B1(n8485), .B2(n8632), .A(n8329), .ZN(n8547) );
  OAI22_X1 U9799 ( .A1(n8547), .A2(n8331), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8330), .ZN(n8332) );
  AOI21_X1 U9800 ( .B1(n8551), .B2(n8333), .A(n8332), .ZN(n8334) );
  OAI211_X1 U9801 ( .C1(n8447), .C2(n8336), .A(n8335), .B(n8334), .ZN(P2_U3242) );
  AOI21_X1 U9802 ( .B1(n8339), .B2(n8338), .A(n8337), .ZN(n8350) );
  INV_X1 U9803 ( .A(n8719), .ZN(n8340) );
  OAI22_X1 U9804 ( .A1(n8342), .A2(n8727), .B1(n8341), .B2(n8340), .ZN(n8343)
         );
  AOI211_X1 U9805 ( .C1(n8345), .C2(n8463), .A(n8344), .B(n8343), .ZN(n8348)
         );
  NAND2_X1 U9806 ( .A1(n8837), .A2(n8346), .ZN(n8347) );
  OAI211_X1 U9807 ( .C1(n8350), .C2(n8349), .A(n8348), .B(n8347), .ZN(P2_U3243) );
  MUX2_X1 U9808 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8450), .S(P2_U3966), .Z(
        P2_U3583) );
  MUX2_X1 U9809 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8493), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9810 ( .A(n8351), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8353), .Z(
        P2_U3581) );
  INV_X1 U9811 ( .A(n8488), .ZN(n8495) );
  MUX2_X1 U9812 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8495), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U9813 ( .A(n8485), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8353), .Z(
        P2_U3579) );
  INV_X1 U9814 ( .A(n8352), .ZN(n8482) );
  MUX2_X1 U9815 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8482), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U9816 ( .A(n8580), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8353), .Z(
        P2_U3577) );
  MUX2_X1 U9817 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n4539), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U9818 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8617), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U9819 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8476), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9820 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8616), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9821 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8631), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9822 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8471), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9823 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8468), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9824 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8465), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9825 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8463), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9826 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8461), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9827 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8458), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9828 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8354), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9829 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8355), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9830 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8356), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9831 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8357), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9832 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8358), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9833 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8359), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9834 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8360), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9835 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8361), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9836 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8362), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9837 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n7077), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9838 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8363), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U9839 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n7009), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U9840 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8364), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U9841 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6945), .S(P2_U3966), .Z(
        P2_U3552) );
  OAI211_X1 U9842 ( .C1(n8367), .C2(n8366), .A(n9912), .B(n8365), .ZN(n8377)
         );
  AOI21_X1 U9843 ( .B1(n9920), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8368), .ZN(
        n8376) );
  NAND2_X1 U9844 ( .A1(n8388), .A2(n8369), .ZN(n8375) );
  OAI21_X1 U9845 ( .B1(n8372), .B2(n8371), .A(n8370), .ZN(n8373) );
  NAND2_X1 U9846 ( .A1(n9914), .A2(n8373), .ZN(n8374) );
  NAND4_X1 U9847 ( .A1(n8377), .A2(n8376), .A3(n8375), .A4(n8374), .ZN(
        P2_U3257) );
  NOR2_X1 U9848 ( .A1(n8379), .A2(n8378), .ZN(n8381) );
  NOR2_X1 U9849 ( .A1(n8381), .A2(n8380), .ZN(n8383) );
  XOR2_X1 U9850 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8407), .Z(n8382) );
  NAND2_X1 U9851 ( .A1(n8382), .A2(n8383), .ZN(n8406) );
  OAI21_X1 U9852 ( .B1(n8383), .B2(n8382), .A(n8406), .ZN(n8384) );
  NAND2_X1 U9853 ( .A1(n8384), .A2(n9914), .ZN(n8398) );
  INV_X1 U9854 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8386) );
  OAI21_X1 U9855 ( .B1(n8446), .B2(n8386), .A(n8385), .ZN(n8387) );
  AOI21_X1 U9856 ( .B1(n8388), .B2(n8407), .A(n8387), .ZN(n8397) );
  NOR2_X1 U9857 ( .A1(n8390), .A2(n8389), .ZN(n8392) );
  NOR2_X1 U9858 ( .A1(n8392), .A2(n8391), .ZN(n8395) );
  MUX2_X1 U9859 ( .A(n5904), .B(P2_REG2_REG_16__SCAN_IN), .S(n8407), .Z(n8393)
         );
  INV_X1 U9860 ( .A(n8393), .ZN(n8394) );
  NAND2_X1 U9861 ( .A1(n8394), .A2(n8395), .ZN(n8399) );
  OAI211_X1 U9862 ( .C1(n8395), .C2(n8394), .A(n9912), .B(n8399), .ZN(n8396)
         );
  NAND3_X1 U9863 ( .A1(n8398), .A2(n8397), .A3(n8396), .ZN(P2_U3261) );
  NAND2_X1 U9864 ( .A1(n8407), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8400) );
  NAND2_X1 U9865 ( .A1(n8400), .A2(n8399), .ZN(n8403) );
  MUX2_X1 U9866 ( .A(n5918), .B(P2_REG2_REG_17__SCAN_IN), .S(n8419), .Z(n8401)
         );
  INV_X1 U9867 ( .A(n8401), .ZN(n8402) );
  NAND2_X1 U9868 ( .A1(n8402), .A2(n8403), .ZN(n8415) );
  OAI211_X1 U9869 ( .C1(n8403), .C2(n8402), .A(n9912), .B(n8415), .ZN(n8414)
         );
  AND2_X1 U9870 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8404) );
  AOI21_X1 U9871 ( .B1(n9920), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8404), .ZN(
        n8413) );
  OR2_X1 U9872 ( .A1(n9915), .A2(n8405), .ZN(n8412) );
  OAI21_X1 U9873 ( .B1(n8407), .B2(P2_REG1_REG_16__SCAN_IN), .A(n8406), .ZN(
        n8409) );
  XNOR2_X1 U9874 ( .A(n8419), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8408) );
  NOR2_X1 U9875 ( .A1(n8408), .A2(n8409), .ZN(n8418) );
  AOI21_X1 U9876 ( .B1(n8409), .B2(n8408), .A(n8418), .ZN(n8410) );
  NAND2_X1 U9877 ( .A1(n9914), .A2(n8410), .ZN(n8411) );
  NAND4_X1 U9878 ( .A1(n8414), .A2(n8413), .A3(n8412), .A4(n8411), .ZN(
        P2_U3262) );
  NAND2_X1 U9879 ( .A1(n8419), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8416) );
  NAND2_X1 U9880 ( .A1(n8416), .A2(n8415), .ZN(n8431) );
  XNOR2_X1 U9881 ( .A(n8432), .B(n8431), .ZN(n8417) );
  NOR2_X1 U9882 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8417), .ZN(n8433) );
  AOI21_X1 U9883 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8417), .A(n8433), .ZN(
        n8429) );
  INV_X1 U9884 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8420) );
  AOI22_X1 U9885 ( .A1(n8432), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n8420), .B2(
        n8425), .ZN(n8421) );
  OAI21_X1 U9886 ( .B1(n8422), .B2(n8421), .A(n8430), .ZN(n8427) );
  NAND2_X1 U9887 ( .A1(n9920), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n8423) );
  OAI211_X1 U9888 ( .C1(n9915), .C2(n8425), .A(n8424), .B(n8423), .ZN(n8426)
         );
  AOI21_X1 U9889 ( .B1(n8427), .B2(n9914), .A(n8426), .ZN(n8428) );
  OAI21_X1 U9890 ( .B1(n8429), .B2(n9917), .A(n8428), .ZN(P2_U3263) );
  INV_X1 U9891 ( .A(n8439), .ZN(n8437) );
  NOR2_X1 U9892 ( .A1(n8432), .A2(n8431), .ZN(n8434) );
  NOR2_X1 U9893 ( .A1(n8434), .A2(n8433), .ZN(n8435) );
  XOR2_X1 U9894 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8435), .Z(n8438) );
  OAI21_X1 U9895 ( .B1(n8438), .B2(n9917), .A(n9915), .ZN(n8436) );
  AOI21_X1 U9896 ( .B1(n8437), .B2(n9914), .A(n8436), .ZN(n8442) );
  AOI22_X1 U9897 ( .A1(n8439), .A2(n9914), .B1(n8438), .B2(n9912), .ZN(n8441)
         );
  MUX2_X1 U9898 ( .A(n8442), .B(n8441), .S(n8440), .Z(n8444) );
  NAND2_X1 U9899 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8443) );
  OAI211_X1 U9900 ( .C1(n8446), .C2(n8445), .A(n8444), .B(n8443), .ZN(P2_U3264) );
  INV_X1 U9901 ( .A(n8824), .ZN(n8668) );
  INV_X1 U9902 ( .A(n8807), .ZN(n8627) );
  INV_X1 U9903 ( .A(n8802), .ZN(n8612) );
  INV_X1 U9904 ( .A(n8788), .ZN(n8564) );
  NAND2_X1 U9905 ( .A1(n8560), .A2(n8447), .ZN(n8529) );
  XNOR2_X1 U9906 ( .A(n8453), .B(n8448), .ZN(n8758) );
  NAND2_X1 U9907 ( .A1(n8758), .A2(n8748), .ZN(n8452) );
  AOI21_X1 U9908 ( .B1(n8449), .B2(P2_B_REG_SCAN_IN), .A(n8728), .ZN(n8494) );
  NAND2_X1 U9909 ( .A1(n8494), .A2(n8450), .ZN(n8762) );
  NOR2_X1 U9910 ( .A1(n8686), .A2(n8762), .ZN(n8455) );
  AOI21_X1 U9911 ( .B1(n8742), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8455), .ZN(
        n8451) );
  OAI211_X1 U9912 ( .C1(n8760), .C2(n8721), .A(n8452), .B(n8451), .ZN(P2_U3265) );
  AOI21_X1 U9913 ( .B1(n8497), .B2(n8454), .A(n8453), .ZN(n8761) );
  NAND2_X1 U9914 ( .A1(n8761), .A2(n8748), .ZN(n8457) );
  AOI21_X1 U9915 ( .B1(n8742), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8455), .ZN(
        n8456) );
  OAI211_X1 U9916 ( .C1(n4773), .C2(n8721), .A(n8457), .B(n8456), .ZN(P2_U3266) );
  NAND2_X1 U9917 ( .A1(n8466), .A2(n8272), .ZN(n8467) );
  NAND2_X1 U9918 ( .A1(n8824), .A2(n8468), .ZN(n8470) );
  OR2_X1 U9919 ( .A1(n8818), .A2(n8471), .ZN(n8472) );
  NAND2_X1 U9920 ( .A1(n8651), .A2(n8472), .ZN(n8473) );
  NAND2_X1 U9921 ( .A1(n8587), .A2(n8594), .ZN(n8586) );
  INV_X1 U9922 ( .A(n8797), .ZN(n8593) );
  NAND2_X1 U9923 ( .A1(n8540), .A2(n8546), .ZN(n8484) );
  NAND2_X1 U9924 ( .A1(n8484), .A2(n8483), .ZN(n8523) );
  NAND2_X1 U9925 ( .A1(n8523), .A2(n8524), .ZN(n8487) );
  NAND2_X1 U9926 ( .A1(n8487), .A2(n8486), .ZN(n8508) );
  XNOR2_X1 U9927 ( .A(n8490), .B(n8489), .ZN(n8764) );
  INV_X1 U9928 ( .A(n8764), .ZN(n8506) );
  AOI22_X1 U9929 ( .A1(n8495), .A2(n8630), .B1(n8494), .B2(n8493), .ZN(n8496)
         );
  OAI21_X1 U9930 ( .B1(n4327), .B2(n8724), .A(n8496), .ZN(n8768) );
  OAI21_X1 U9931 ( .B1(n8498), .B2(n8502), .A(n8497), .ZN(n8765) );
  NOR2_X1 U9932 ( .A1(n8765), .A2(n8530), .ZN(n8504) );
  INV_X1 U9933 ( .A(n8499), .ZN(n8500) );
  AOI22_X1 U9934 ( .A1(n8742), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8500), .B2(
        n8746), .ZN(n8501) );
  OAI21_X1 U9935 ( .B1(n8502), .B2(n8721), .A(n8501), .ZN(n8503) );
  AOI211_X1 U9936 ( .C1(n8768), .C2(n8667), .A(n8504), .B(n8503), .ZN(n8505)
         );
  OAI21_X1 U9937 ( .B1(n8506), .B2(n8735), .A(n8505), .ZN(P2_U3267) );
  XNOR2_X1 U9938 ( .A(n8511), .B(n8777), .ZN(n8771) );
  AOI22_X1 U9939 ( .A1(n8742), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8509), .B2(
        n8746), .ZN(n8510) );
  OAI21_X1 U9940 ( .B1(n8511), .B2(n8721), .A(n8510), .ZN(n8521) );
  INV_X1 U9941 ( .A(n8513), .ZN(n8515) );
  AOI21_X1 U9942 ( .B1(n8515), .B2(n8514), .A(n8724), .ZN(n8519) );
  OAI22_X1 U9943 ( .A1(n8517), .A2(n8728), .B1(n8516), .B2(n8726), .ZN(n8518)
         );
  NOR2_X1 U9944 ( .A1(n8773), .A2(n8686), .ZN(n8520) );
  AOI211_X1 U9945 ( .C1(n8748), .C2(n8771), .A(n8521), .B(n8520), .ZN(n8522)
         );
  OAI21_X1 U9946 ( .B1(n8774), .B2(n8735), .A(n8522), .ZN(P2_U3268) );
  XNOR2_X1 U9947 ( .A(n8523), .B(n4779), .ZN(n8781) );
  AOI21_X1 U9948 ( .B1(n8525), .B2(n8524), .A(n8724), .ZN(n8527) );
  AOI21_X1 U9949 ( .B1(n8528), .B2(n8527), .A(n8526), .ZN(n8780) );
  INV_X1 U9950 ( .A(n8780), .ZN(n8538) );
  INV_X1 U9951 ( .A(n8529), .ZN(n8549) );
  INV_X1 U9952 ( .A(n8776), .ZN(n8535) );
  NOR2_X1 U9953 ( .A1(n8549), .A2(n8535), .ZN(n8775) );
  INV_X1 U9954 ( .A(n8777), .ZN(n8531) );
  NOR3_X1 U9955 ( .A1(n8775), .A2(n8531), .A3(n8530), .ZN(n8537) );
  INV_X1 U9956 ( .A(n8532), .ZN(n8533) );
  AOI22_X1 U9957 ( .A1(n8742), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8533), .B2(
        n8746), .ZN(n8534) );
  OAI21_X1 U9958 ( .B1(n8535), .B2(n8721), .A(n8534), .ZN(n8536) );
  AOI211_X1 U9959 ( .C1(n8538), .C2(n8667), .A(n8537), .B(n8536), .ZN(n8539)
         );
  OAI21_X1 U9960 ( .B1(n8781), .B2(n8735), .A(n8539), .ZN(P2_U3269) );
  XOR2_X1 U9961 ( .A(n8540), .B(n8546), .Z(n8786) );
  AOI22_X1 U9962 ( .A1(n8784), .A2(n8753), .B1(n8742), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8558) );
  NAND2_X1 U9963 ( .A1(n8541), .A2(n8542), .ZN(n8545) );
  INV_X1 U9964 ( .A(n8543), .ZN(n8544) );
  AOI21_X1 U9965 ( .B1(n8546), .B2(n8545), .A(n8544), .ZN(n8548) );
  OAI21_X1 U9966 ( .B1(n8548), .B2(n8724), .A(n8547), .ZN(n8782) );
  INV_X1 U9967 ( .A(n8560), .ZN(n8550) );
  AOI211_X1 U9968 ( .C1(n8784), .C2(n8550), .A(n9981), .B(n8549), .ZN(n8783)
         );
  INV_X1 U9969 ( .A(n8783), .ZN(n8555) );
  INV_X1 U9970 ( .A(n8551), .ZN(n8552) );
  OAI22_X1 U9971 ( .A1(n8555), .A2(n8554), .B1(n8553), .B2(n8552), .ZN(n8556)
         );
  OAI21_X1 U9972 ( .B1(n8782), .B2(n8556), .A(n8667), .ZN(n8557) );
  OAI211_X1 U9973 ( .C1(n8786), .C2(n8735), .A(n8558), .B(n8557), .ZN(P2_U3270) );
  XOR2_X1 U9974 ( .A(n8559), .B(n8567), .Z(n8791) );
  AOI211_X1 U9975 ( .C1(n8788), .C2(n4365), .A(n9981), .B(n8560), .ZN(n8787)
         );
  INV_X1 U9976 ( .A(n8561), .ZN(n8562) );
  AOI22_X1 U9977 ( .A1(n8742), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8562), .B2(
        n8746), .ZN(n8563) );
  OAI21_X1 U9978 ( .B1(n8564), .B2(n8721), .A(n8563), .ZN(n8572) );
  NOR2_X1 U9979 ( .A1(n8567), .A2(n4782), .ZN(n8568) );
  AOI21_X1 U9980 ( .B1(n8565), .B2(n8568), .A(n8724), .ZN(n8570) );
  AOI21_X1 U9981 ( .B1(n8541), .B2(n8570), .A(n8569), .ZN(n8790) );
  NOR2_X1 U9982 ( .A1(n8790), .A2(n8686), .ZN(n8571) );
  AOI211_X1 U9983 ( .C1(n8787), .C2(n8695), .A(n8572), .B(n8571), .ZN(n8573)
         );
  OAI21_X1 U9984 ( .B1(n8791), .B2(n8735), .A(n8573), .ZN(P2_U3271) );
  AOI21_X1 U9985 ( .B1(n8579), .B2(n8575), .A(n8574), .ZN(n8796) );
  XNOR2_X1 U9986 ( .A(n8588), .B(n4486), .ZN(n8793) );
  AOI22_X1 U9987 ( .A1(n8742), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8576), .B2(
        n8746), .ZN(n8577) );
  OAI21_X1 U9988 ( .B1(n4486), .B2(n8721), .A(n8577), .ZN(n8584) );
  OAI211_X1 U9989 ( .C1(n8579), .C2(n8578), .A(n8565), .B(n8740), .ZN(n8582)
         );
  AOI22_X1 U9990 ( .A1(n8580), .A2(n8632), .B1(n8630), .B2(n8617), .ZN(n8581)
         );
  AND2_X1 U9991 ( .A1(n8582), .A2(n8581), .ZN(n8795) );
  NOR2_X1 U9992 ( .A1(n8795), .A2(n8742), .ZN(n8583) );
  AOI211_X1 U9993 ( .C1(n8793), .C2(n8748), .A(n8584), .B(n8583), .ZN(n8585)
         );
  OAI21_X1 U9994 ( .B1(n8796), .B2(n8735), .A(n8585), .ZN(P2_U3272) );
  OAI21_X1 U9995 ( .B1(n8587), .B2(n8594), .A(n8586), .ZN(n8801) );
  INV_X1 U9996 ( .A(n8588), .ZN(n8589) );
  AOI21_X1 U9997 ( .B1(n8797), .B2(n8606), .A(n8589), .ZN(n8798) );
  INV_X1 U9998 ( .A(n8590), .ZN(n8591) );
  AOI22_X1 U9999 ( .A1(n8742), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8591), .B2(
        n8746), .ZN(n8592) );
  OAI21_X1 U10000 ( .B1(n8593), .B2(n8721), .A(n8592), .ZN(n8602) );
  INV_X1 U10001 ( .A(n8613), .ZN(n8596) );
  OAI21_X1 U10002 ( .B1(n8596), .B2(n8595), .A(n8594), .ZN(n8598) );
  AOI21_X1 U10003 ( .B1(n8598), .B2(n8597), .A(n8724), .ZN(n8600) );
  NOR2_X1 U10004 ( .A1(n8600), .A2(n8599), .ZN(n8800) );
  NOR2_X1 U10005 ( .A1(n8800), .A2(n8686), .ZN(n8601) );
  AOI211_X1 U10006 ( .C1(n8798), .C2(n8748), .A(n8602), .B(n8601), .ZN(n8603)
         );
  OAI21_X1 U10007 ( .B1(n8735), .B2(n8801), .A(n8603), .ZN(P2_U3273) );
  XNOR2_X1 U10008 ( .A(n8604), .B(n8614), .ZN(n8806) );
  INV_X1 U10009 ( .A(n8605), .ZN(n8608) );
  INV_X1 U10010 ( .A(n8606), .ZN(n8607) );
  AOI21_X1 U10011 ( .B1(n8802), .B2(n8608), .A(n8607), .ZN(n8803) );
  INV_X1 U10012 ( .A(n8609), .ZN(n8610) );
  AOI22_X1 U10013 ( .A1(n8686), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8610), .B2(
        n8746), .ZN(n8611) );
  OAI21_X1 U10014 ( .B1(n8612), .B2(n8721), .A(n8611), .ZN(n8621) );
  OAI211_X1 U10015 ( .C1(n8615), .C2(n8614), .A(n8613), .B(n8740), .ZN(n8619)
         );
  AOI22_X1 U10016 ( .A1(n8617), .A2(n8632), .B1(n8630), .B2(n8616), .ZN(n8618)
         );
  AND2_X1 U10017 ( .A1(n8619), .A2(n8618), .ZN(n8805) );
  NOR2_X1 U10018 ( .A1(n8805), .A2(n8686), .ZN(n8620) );
  AOI211_X1 U10019 ( .C1(n8803), .C2(n8748), .A(n8621), .B(n8620), .ZN(n8622)
         );
  OAI21_X1 U10020 ( .B1(n8806), .B2(n8735), .A(n8622), .ZN(P2_U3274) );
  XNOR2_X1 U10021 ( .A(n8623), .B(n8628), .ZN(n8811) );
  XNOR2_X1 U10022 ( .A(n8638), .B(n8807), .ZN(n8808) );
  INV_X1 U10023 ( .A(n8624), .ZN(n8625) );
  AOI22_X1 U10024 ( .A1(n8686), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8625), .B2(
        n8746), .ZN(n8626) );
  OAI21_X1 U10025 ( .B1(n8627), .B2(n8721), .A(n8626), .ZN(n8635) );
  XNOR2_X1 U10026 ( .A(n8629), .B(n8628), .ZN(n8633) );
  AOI222_X1 U10027 ( .A1(n8740), .A2(n8633), .B1(n8476), .B2(n8632), .C1(n8631), .C2(n8630), .ZN(n8810) );
  NOR2_X1 U10028 ( .A1(n8810), .A2(n8742), .ZN(n8634) );
  AOI211_X1 U10029 ( .C1(n8808), .C2(n8748), .A(n8635), .B(n8634), .ZN(n8636)
         );
  OAI21_X1 U10030 ( .B1(n8811), .B2(n8735), .A(n8636), .ZN(P2_U3275) );
  XNOR2_X1 U10031 ( .A(n8637), .B(n8643), .ZN(n8816) );
  AOI21_X1 U10032 ( .B1(n8812), .B2(n8652), .A(n8638), .ZN(n8813) );
  INV_X1 U10033 ( .A(n8812), .ZN(n8641) );
  AOI22_X1 U10034 ( .A1(n8686), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8639), .B2(
        n8746), .ZN(n8640) );
  OAI21_X1 U10035 ( .B1(n8641), .B2(n8721), .A(n8640), .ZN(n8649) );
  AOI211_X1 U10036 ( .C1(n8643), .C2(n4363), .A(n8724), .B(n8642), .ZN(n8647)
         );
  OAI22_X1 U10037 ( .A1(n8645), .A2(n8728), .B1(n8644), .B2(n8726), .ZN(n8646)
         );
  NOR2_X1 U10038 ( .A1(n8647), .A2(n8646), .ZN(n8815) );
  NOR2_X1 U10039 ( .A1(n8815), .A2(n8686), .ZN(n8648) );
  AOI211_X1 U10040 ( .C1(n8813), .C2(n8748), .A(n8649), .B(n8648), .ZN(n8650)
         );
  OAI21_X1 U10041 ( .B1(n8735), .B2(n8816), .A(n8650), .ZN(P2_U3276) );
  XNOR2_X1 U10042 ( .A(n8651), .B(n4760), .ZN(n8821) );
  AOI211_X1 U10043 ( .C1(n8818), .C2(n8664), .A(n9981), .B(n4501), .ZN(n8817)
         );
  AOI22_X1 U10044 ( .A1(n8686), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8653), .B2(
        n8746), .ZN(n8654) );
  OAI21_X1 U10045 ( .B1(n8655), .B2(n8721), .A(n8654), .ZN(n8661) );
  XNOR2_X1 U10046 ( .A(n8657), .B(n8656), .ZN(n8659) );
  AOI21_X1 U10047 ( .B1(n8659), .B2(n8740), .A(n8658), .ZN(n8820) );
  NOR2_X1 U10048 ( .A1(n8820), .A2(n8742), .ZN(n8660) );
  AOI211_X1 U10049 ( .C1(n8817), .C2(n8695), .A(n8661), .B(n8660), .ZN(n8662)
         );
  OAI21_X1 U10050 ( .B1(n8821), .B2(n8735), .A(n8662), .ZN(P2_U3277) );
  XNOR2_X1 U10051 ( .A(n8663), .B(n8672), .ZN(n8826) );
  INV_X1 U10052 ( .A(n8684), .ZN(n8665) );
  AOI211_X1 U10053 ( .C1(n8824), .C2(n8665), .A(n9981), .B(n4503), .ZN(n8823)
         );
  OAI22_X1 U10054 ( .A1(n8668), .A2(n8721), .B1(n8667), .B2(n8666), .ZN(n8678)
         );
  INV_X1 U10055 ( .A(n8669), .ZN(n8670) );
  NOR2_X1 U10056 ( .A1(n8688), .A2(n8670), .ZN(n8671) );
  XOR2_X1 U10057 ( .A(n8672), .B(n8671), .Z(n8674) );
  OAI21_X1 U10058 ( .B1(n8674), .B2(n8724), .A(n8673), .ZN(n8822) );
  AOI21_X1 U10059 ( .B1(n8675), .B2(n8746), .A(n8822), .ZN(n8676) );
  NOR2_X1 U10060 ( .A1(n8676), .A2(n8686), .ZN(n8677) );
  AOI211_X1 U10061 ( .C1(n8823), .C2(n8679), .A(n8678), .B(n8677), .ZN(n8680)
         );
  OAI21_X1 U10062 ( .B1(n8826), .B2(n8735), .A(n8680), .ZN(P2_U3278) );
  OAI21_X1 U10063 ( .B1(n8682), .B2(n8690), .A(n8681), .ZN(n8683) );
  INV_X1 U10064 ( .A(n8683), .ZN(n8831) );
  AOI211_X1 U10065 ( .C1(n8828), .C2(n8700), .A(n9981), .B(n8684), .ZN(n8827)
         );
  AOI22_X1 U10066 ( .A1(n8686), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8685), .B2(
        n8746), .ZN(n8687) );
  OAI21_X1 U10067 ( .B1(n8466), .B2(n8721), .A(n8687), .ZN(n8694) );
  AOI211_X1 U10068 ( .C1(n8690), .C2(n8689), .A(n8724), .B(n8688), .ZN(n8692)
         );
  NOR2_X1 U10069 ( .A1(n8692), .A2(n8691), .ZN(n8830) );
  NOR2_X1 U10070 ( .A1(n8830), .A2(n8742), .ZN(n8693) );
  AOI211_X1 U10071 ( .C1(n8827), .C2(n8695), .A(n8694), .B(n8693), .ZN(n8696)
         );
  OAI21_X1 U10072 ( .B1(n8735), .B2(n8831), .A(n8696), .ZN(P2_U3279) );
  AOI21_X1 U10073 ( .B1(n8707), .B2(n8698), .A(n8697), .ZN(n8699) );
  INV_X1 U10074 ( .A(n8699), .ZN(n8836) );
  INV_X1 U10075 ( .A(n8700), .ZN(n8701) );
  AOI21_X1 U10076 ( .B1(n8832), .B2(n8717), .A(n8701), .ZN(n8833) );
  AOI22_X1 U10077 ( .A1(n8742), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8702), .B2(
        n8746), .ZN(n8703) );
  OAI21_X1 U10078 ( .B1(n8704), .B2(n8721), .A(n8703), .ZN(n8712) );
  INV_X1 U10079 ( .A(n8705), .ZN(n8706) );
  NOR2_X1 U10080 ( .A1(n8723), .A2(n8706), .ZN(n8708) );
  XNOR2_X1 U10081 ( .A(n8708), .B(n8707), .ZN(n8710) );
  AOI21_X1 U10082 ( .B1(n8710), .B2(n8740), .A(n8709), .ZN(n8835) );
  NOR2_X1 U10083 ( .A1(n8835), .A2(n8742), .ZN(n8711) );
  AOI211_X1 U10084 ( .C1(n8833), .C2(n8748), .A(n8712), .B(n8711), .ZN(n8713)
         );
  OAI21_X1 U10085 ( .B1(n8735), .B2(n8836), .A(n8713), .ZN(P2_U3280) );
  OAI21_X1 U10086 ( .B1(n8715), .B2(n8725), .A(n8714), .ZN(n8716) );
  INV_X1 U10087 ( .A(n8716), .ZN(n8841) );
  AOI21_X1 U10088 ( .B1(n8837), .B2(n8718), .A(n4490), .ZN(n8838) );
  INV_X1 U10089 ( .A(n8837), .ZN(n8722) );
  AOI22_X1 U10090 ( .A1(n8742), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8719), .B2(
        n8746), .ZN(n8720) );
  OAI21_X1 U10091 ( .B1(n8722), .B2(n8721), .A(n8720), .ZN(n8733) );
  AOI211_X1 U10092 ( .C1(n4368), .C2(n8725), .A(n8724), .B(n8723), .ZN(n8731)
         );
  OAI22_X1 U10093 ( .A1(n8729), .A2(n8728), .B1(n8727), .B2(n8726), .ZN(n8730)
         );
  NOR2_X1 U10094 ( .A1(n8731), .A2(n8730), .ZN(n8840) );
  NOR2_X1 U10095 ( .A1(n8840), .A2(n8742), .ZN(n8732) );
  AOI211_X1 U10096 ( .C1(n8838), .C2(n8748), .A(n8733), .B(n8732), .ZN(n8734)
         );
  OAI21_X1 U10097 ( .B1(n8841), .B2(n8735), .A(n8734), .ZN(P2_U3281) );
  NAND2_X1 U10098 ( .A1(n8737), .A2(n8736), .ZN(n8738) );
  XOR2_X1 U10099 ( .A(n8750), .B(n8738), .Z(n8741) );
  AOI21_X1 U10100 ( .B1(n8741), .B2(n8740), .A(n8739), .ZN(n9954) );
  MUX2_X1 U10101 ( .A(n9954), .B(n8743), .S(n8742), .Z(n8757) );
  AOI21_X1 U10102 ( .B1(n8752), .B2(n8745), .A(n8744), .ZN(n9951) );
  AOI22_X1 U10103 ( .A1(n8748), .A2(n9951), .B1(n8747), .B2(n8746), .ZN(n8756)
         );
  OAI21_X1 U10104 ( .B1(n8751), .B2(n8750), .A(n8749), .ZN(n9957) );
  AOI22_X1 U10105 ( .A1(n9957), .A2(n8754), .B1(n8753), .B2(n8752), .ZN(n8755)
         );
  NAND3_X1 U10106 ( .A1(n8757), .A2(n8756), .A3(n8755), .ZN(P2_U3292) );
  NAND2_X1 U10107 ( .A1(n8758), .A2(n8857), .ZN(n8759) );
  OAI211_X1 U10108 ( .C1(n8760), .C2(n9980), .A(n8759), .B(n8762), .ZN(n8864)
         );
  MUX2_X1 U10109 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8864), .S(n10001), .Z(
        P2_U3551) );
  NAND2_X1 U10110 ( .A1(n8761), .A2(n8857), .ZN(n8763) );
  OAI211_X1 U10111 ( .C1(n4773), .C2(n9980), .A(n8763), .B(n8762), .ZN(n8865)
         );
  MUX2_X1 U10112 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8865), .S(n10001), .Z(
        P2_U3550) );
  NAND2_X1 U10113 ( .A1(n8764), .A2(n9985), .ZN(n8769) );
  MUX2_X1 U10114 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8866), .S(n10001), .Z(
        P2_U3549) );
  AOI22_X1 U10115 ( .A1(n8771), .A2(n8857), .B1(n8856), .B2(n8770), .ZN(n8772)
         );
  OAI211_X1 U10116 ( .C1(n8774), .C2(n8861), .A(n8773), .B(n8772), .ZN(n8867)
         );
  MUX2_X1 U10117 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8867), .S(n10001), .Z(
        P2_U3548) );
  NOR2_X1 U10118 ( .A1(n8775), .A2(n9981), .ZN(n8778) );
  AOI22_X1 U10119 ( .A1(n8778), .A2(n8777), .B1(n8856), .B2(n8776), .ZN(n8779)
         );
  OAI211_X1 U10120 ( .C1(n8781), .C2(n8861), .A(n8780), .B(n8779), .ZN(n8868)
         );
  MUX2_X1 U10121 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8868), .S(n10001), .Z(
        P2_U3547) );
  AOI211_X1 U10122 ( .C1(n8856), .C2(n8784), .A(n8783), .B(n8782), .ZN(n8785)
         );
  OAI21_X1 U10123 ( .B1(n8786), .B2(n8861), .A(n8785), .ZN(n8869) );
  MUX2_X1 U10124 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8869), .S(n10001), .Z(
        P2_U3546) );
  AOI21_X1 U10125 ( .B1(n8856), .B2(n8788), .A(n8787), .ZN(n8789) );
  OAI211_X1 U10126 ( .C1(n8791), .C2(n8861), .A(n8790), .B(n8789), .ZN(n8870)
         );
  MUX2_X1 U10127 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8870), .S(n10001), .Z(
        P2_U3545) );
  AOI22_X1 U10128 ( .A1(n8793), .A2(n8857), .B1(n8856), .B2(n8792), .ZN(n8794)
         );
  OAI211_X1 U10129 ( .C1(n8796), .C2(n8861), .A(n8795), .B(n8794), .ZN(n8871)
         );
  MUX2_X1 U10130 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8871), .S(n10001), .Z(
        P2_U3544) );
  AOI22_X1 U10131 ( .A1(n8798), .A2(n8857), .B1(n8856), .B2(n8797), .ZN(n8799)
         );
  OAI211_X1 U10132 ( .C1(n8861), .C2(n8801), .A(n8800), .B(n8799), .ZN(n8872)
         );
  MUX2_X1 U10133 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8872), .S(n10001), .Z(
        P2_U3543) );
  AOI22_X1 U10134 ( .A1(n8803), .A2(n8857), .B1(n8856), .B2(n8802), .ZN(n8804)
         );
  OAI211_X1 U10135 ( .C1(n8806), .C2(n8861), .A(n8805), .B(n8804), .ZN(n8873)
         );
  MUX2_X1 U10136 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8873), .S(n10001), .Z(
        P2_U3542) );
  AOI22_X1 U10137 ( .A1(n8808), .A2(n8857), .B1(n8856), .B2(n8807), .ZN(n8809)
         );
  OAI211_X1 U10138 ( .C1(n8861), .C2(n8811), .A(n8810), .B(n8809), .ZN(n8874)
         );
  MUX2_X1 U10139 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8874), .S(n10001), .Z(
        P2_U3541) );
  AOI22_X1 U10140 ( .A1(n8813), .A2(n8857), .B1(n8856), .B2(n8812), .ZN(n8814)
         );
  OAI211_X1 U10141 ( .C1(n8861), .C2(n8816), .A(n8815), .B(n8814), .ZN(n8875)
         );
  MUX2_X1 U10142 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8875), .S(n10001), .Z(
        P2_U3540) );
  AOI21_X1 U10143 ( .B1(n8856), .B2(n8818), .A(n8817), .ZN(n8819) );
  OAI211_X1 U10144 ( .C1(n8821), .C2(n8861), .A(n8820), .B(n8819), .ZN(n8876)
         );
  MUX2_X1 U10145 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8876), .S(n10001), .Z(
        P2_U3539) );
  AOI211_X1 U10146 ( .C1(n8856), .C2(n8824), .A(n8823), .B(n8822), .ZN(n8825)
         );
  OAI21_X1 U10147 ( .B1(n8861), .B2(n8826), .A(n8825), .ZN(n8877) );
  MUX2_X1 U10148 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8877), .S(n10001), .Z(
        P2_U3538) );
  AOI21_X1 U10149 ( .B1(n8856), .B2(n8828), .A(n8827), .ZN(n8829) );
  OAI211_X1 U10150 ( .C1(n8861), .C2(n8831), .A(n8830), .B(n8829), .ZN(n8878)
         );
  MUX2_X1 U10151 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8878), .S(n10001), .Z(
        P2_U3537) );
  AOI22_X1 U10152 ( .A1(n8833), .A2(n8857), .B1(n8856), .B2(n8832), .ZN(n8834)
         );
  OAI211_X1 U10153 ( .C1(n8836), .C2(n8861), .A(n8835), .B(n8834), .ZN(n8879)
         );
  MUX2_X1 U10154 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8879), .S(n10001), .Z(
        P2_U3536) );
  AOI22_X1 U10155 ( .A1(n8838), .A2(n8857), .B1(n8856), .B2(n8837), .ZN(n8839)
         );
  OAI211_X1 U10156 ( .C1(n8861), .C2(n8841), .A(n8840), .B(n8839), .ZN(n8880)
         );
  MUX2_X1 U10157 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8880), .S(n10001), .Z(
        P2_U3535) );
  AOI22_X1 U10158 ( .A1(n8843), .A2(n8857), .B1(n8856), .B2(n8842), .ZN(n8844)
         );
  OAI211_X1 U10159 ( .C1(n8861), .C2(n8846), .A(n8845), .B(n8844), .ZN(n8881)
         );
  MUX2_X1 U10160 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8881), .S(n10001), .Z(
        P2_U3534) );
  INV_X1 U10161 ( .A(n8847), .ZN(n8853) );
  OAI22_X1 U10162 ( .A1(n8849), .A2(n9981), .B1(n8848), .B2(n9980), .ZN(n8850)
         );
  INV_X1 U10163 ( .A(n8850), .ZN(n8851) );
  OAI211_X1 U10164 ( .C1(n8854), .C2(n8853), .A(n8852), .B(n8851), .ZN(n8882)
         );
  MUX2_X1 U10165 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8882), .S(n10001), .Z(
        P2_U3533) );
  AOI22_X1 U10166 ( .A1(n8858), .A2(n8857), .B1(n8856), .B2(n8855), .ZN(n8859)
         );
  OAI211_X1 U10167 ( .C1(n8862), .C2(n8861), .A(n8860), .B(n8859), .ZN(n8883)
         );
  MUX2_X1 U10168 ( .A(n8883), .B(P2_REG1_REG_11__SCAN_IN), .S(n9999), .Z(
        P2_U3531) );
  MUX2_X1 U10169 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n8863), .S(n10001), .Z(
        P2_U3527) );
  MUX2_X1 U10170 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8864), .S(n9988), .Z(
        P2_U3519) );
  MUX2_X1 U10171 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8865), .S(n9988), .Z(
        P2_U3518) );
  MUX2_X1 U10172 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8866), .S(n9988), .Z(
        P2_U3517) );
  MUX2_X1 U10173 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8867), .S(n9988), .Z(
        P2_U3516) );
  MUX2_X1 U10174 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8868), .S(n9988), .Z(
        P2_U3515) );
  MUX2_X1 U10175 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8869), .S(n9988), .Z(
        P2_U3514) );
  MUX2_X1 U10176 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8870), .S(n9988), .Z(
        P2_U3513) );
  MUX2_X1 U10177 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8871), .S(n9988), .Z(
        P2_U3512) );
  MUX2_X1 U10178 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8872), .S(n9988), .Z(
        P2_U3511) );
  MUX2_X1 U10179 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8873), .S(n9988), .Z(
        P2_U3510) );
  MUX2_X1 U10180 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8874), .S(n9988), .Z(
        P2_U3509) );
  MUX2_X1 U10181 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8875), .S(n9988), .Z(
        P2_U3508) );
  MUX2_X1 U10182 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8876), .S(n9988), .Z(
        P2_U3507) );
  MUX2_X1 U10183 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8877), .S(n9988), .Z(
        P2_U3505) );
  MUX2_X1 U10184 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8878), .S(n9988), .Z(
        P2_U3502) );
  MUX2_X1 U10185 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8879), .S(n9988), .Z(
        P2_U3499) );
  MUX2_X1 U10186 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8880), .S(n9988), .Z(
        P2_U3496) );
  MUX2_X1 U10187 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8881), .S(n9988), .Z(
        P2_U3493) );
  MUX2_X1 U10188 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8882), .S(n9988), .Z(
        P2_U3490) );
  MUX2_X1 U10189 ( .A(n8883), .B(P2_REG0_REG_11__SCAN_IN), .S(n9987), .Z(
        P2_U3484) );
  INV_X1 U10190 ( .A(n8884), .ZN(n9649) );
  NOR4_X1 U10191 ( .A1(n8885), .A2(P2_IR_REG_30__SCAN_IN), .A3(n5818), .A4(
        P2_U3152), .ZN(n8886) );
  AOI21_X1 U10192 ( .B1(n8889), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8886), .ZN(
        n8887) );
  OAI21_X1 U10193 ( .B1(n9649), .B2(n8195), .A(n8887), .ZN(P2_U3327) );
  INV_X1 U10194 ( .A(n8888), .ZN(n9654) );
  AOI22_X1 U10195 ( .A1(n8890), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8889), .ZN(n8891) );
  OAI21_X1 U10196 ( .B1(n9654), .B2(n8195), .A(n8891), .ZN(P2_U3328) );
  MUX2_X1 U10197 ( .A(n8892), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  OAI22_X1 U10198 ( .A1(n9032), .A2(n9224), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8896), .ZN(n8899) );
  INV_X1 U10199 ( .A(n9194), .ZN(n8897) );
  OAI22_X1 U10200 ( .A1(n9008), .A2(n8897), .B1(n9035), .B2(n9197), .ZN(n8898)
         );
  AOI211_X1 U10201 ( .C1(n9379), .C2(n9038), .A(n8899), .B(n8898), .ZN(n8900)
         );
  OAI21_X1 U10202 ( .B1(n8901), .B2(n9012), .A(n8900), .ZN(P1_U3212) );
  INV_X1 U10203 ( .A(n8902), .ZN(n8904) );
  NAND2_X1 U10204 ( .A1(n8904), .A2(n8903), .ZN(n8906) );
  XNOR2_X1 U10205 ( .A(n8906), .B(n8905), .ZN(n8912) );
  OAI22_X1 U10206 ( .A1(n9032), .A2(n9130), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8907), .ZN(n8910) );
  INV_X1 U10207 ( .A(n9256), .ZN(n8908) );
  OAI22_X1 U10208 ( .A1(n9008), .A2(n8908), .B1(n9035), .B2(n9259), .ZN(n8909)
         );
  AOI211_X1 U10209 ( .C1(n9399), .C2(n9038), .A(n8910), .B(n8909), .ZN(n8911)
         );
  OAI21_X1 U10210 ( .B1(n8912), .B2(n9012), .A(n8911), .ZN(P1_U3214) );
  XOR2_X1 U10211 ( .A(n8913), .B(n8914), .Z(n8918) );
  NAND2_X1 U10212 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9112) );
  OAI21_X1 U10213 ( .B1(n9128), .B2(n9035), .A(n9112), .ZN(n8916) );
  OAI22_X1 U10214 ( .A1(n9008), .A2(n9318), .B1(n9032), .B2(n8960), .ZN(n8915)
         );
  AOI211_X1 U10215 ( .C1(n9419), .C2(n9038), .A(n8916), .B(n8915), .ZN(n8917)
         );
  OAI21_X1 U10216 ( .B1(n8918), .B2(n9012), .A(n8917), .ZN(P1_U3217) );
  NAND2_X1 U10217 ( .A1(n8920), .A2(n8919), .ZN(n8922) );
  XNOR2_X1 U10218 ( .A(n8922), .B(n8921), .ZN(n8923) );
  NAND2_X1 U10219 ( .A1(n8923), .A2(n5630), .ZN(n8930) );
  INV_X1 U10220 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8924) );
  NOR2_X1 U10221 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8924), .ZN(n9797) );
  AOI21_X1 U10222 ( .B1(n9020), .B2(n9049), .A(n9797), .ZN(n8929) );
  AOI22_X1 U10223 ( .A1(n9022), .A2(n9047), .B1(n9033), .B2(n8925), .ZN(n8928)
         );
  AND2_X1 U10224 ( .A1(n8926), .A2(n9887), .ZN(n9877) );
  NAND2_X1 U10225 ( .A1(n9877), .A2(n9024), .ZN(n8927) );
  NAND4_X1 U10226 ( .A1(n8930), .A2(n8929), .A3(n8928), .A4(n8927), .ZN(
        P1_U3219) );
  XOR2_X1 U10227 ( .A(n8931), .B(n8932), .Z(n8938) );
  OAI22_X1 U10228 ( .A1(n9035), .A2(n9130), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8933), .ZN(n8936) );
  INV_X1 U10229 ( .A(n9289), .ZN(n8934) );
  OAI22_X1 U10230 ( .A1(n8934), .A2(n9008), .B1(n9128), .B2(n9032), .ZN(n8935)
         );
  AOI211_X1 U10231 ( .C1(n9409), .C2(n9038), .A(n8936), .B(n8935), .ZN(n8937)
         );
  OAI21_X1 U10232 ( .B1(n8938), .B2(n9012), .A(n8937), .ZN(P1_U3221) );
  XOR2_X1 U10233 ( .A(n8940), .B(n8939), .Z(n8945) );
  OAI22_X1 U10234 ( .A1(n9035), .A2(n9224), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9583), .ZN(n8943) );
  INV_X1 U10235 ( .A(n9234), .ZN(n8941) );
  OAI22_X1 U10236 ( .A1(n9008), .A2(n8941), .B1(n9032), .B2(n9259), .ZN(n8942)
         );
  AOI211_X1 U10237 ( .C1(n9389), .C2(n9038), .A(n8943), .B(n8942), .ZN(n8944)
         );
  OAI21_X1 U10238 ( .B1(n8945), .B2(n9012), .A(n8944), .ZN(P1_U3223) );
  INV_X1 U10239 ( .A(n8946), .ZN(n8947) );
  AOI21_X1 U10240 ( .B1(n8949), .B2(n8948), .A(n8947), .ZN(n8956) );
  NOR2_X1 U10241 ( .A1(n8950), .A2(n9852), .ZN(n9434) );
  AOI22_X1 U10242 ( .A1(n9020), .A2(n9042), .B1(n8951), .B2(n9033), .ZN(n8953)
         );
  OAI211_X1 U10243 ( .C1(n9121), .C2(n9035), .A(n8953), .B(n8952), .ZN(n8954)
         );
  AOI21_X1 U10244 ( .B1(n9434), .B2(n9024), .A(n8954), .ZN(n8955) );
  OAI21_X1 U10245 ( .B1(n8956), .B2(n9012), .A(n8955), .ZN(P1_U3224) );
  XOR2_X1 U10246 ( .A(n8958), .B(n8957), .Z(n8963) );
  AOI22_X1 U10247 ( .A1(n9020), .A2(n9348), .B1(n9343), .B2(n9033), .ZN(n8959)
         );
  NAND2_X1 U10248 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9070) );
  OAI211_X1 U10249 ( .C1(n8960), .C2(n9035), .A(n8959), .B(n9070), .ZN(n8961)
         );
  AOI21_X1 U10250 ( .B1(n9428), .B2(n9038), .A(n8961), .ZN(n8962) );
  OAI21_X1 U10251 ( .B1(n8963), .B2(n9012), .A(n8962), .ZN(P1_U3226) );
  XOR2_X1 U10252 ( .A(n8965), .B(n8964), .Z(n8971) );
  INV_X1 U10253 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8966) );
  OAI22_X1 U10254 ( .A1(n9035), .A2(n9135), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8966), .ZN(n8969) );
  OAI22_X1 U10255 ( .A1(n9008), .A2(n8967), .B1(n9032), .B2(n9131), .ZN(n8968)
         );
  AOI211_X1 U10256 ( .C1(n9394), .C2(n9038), .A(n8969), .B(n8968), .ZN(n8970)
         );
  OAI21_X1 U10257 ( .B1(n8971), .B2(n9012), .A(n8970), .ZN(P1_U3227) );
  NAND2_X1 U10258 ( .A1(n8973), .A2(n8972), .ZN(n8975) );
  OAI21_X1 U10259 ( .B1(n8976), .B2(n8975), .A(n8974), .ZN(n8977) );
  NAND2_X1 U10260 ( .A1(n8977), .A2(n5630), .ZN(n8984) );
  AOI22_X1 U10261 ( .A1(n9022), .A2(n9051), .B1(n9038), .B2(n8978), .ZN(n8983)
         );
  NAND2_X1 U10262 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9781) );
  INV_X1 U10263 ( .A(n9781), .ZN(n8980) );
  NOR2_X1 U10264 ( .A1(n9032), .A2(n4993), .ZN(n8979) );
  AOI211_X1 U10265 ( .C1(n9033), .C2(n8981), .A(n8980), .B(n8979), .ZN(n8982)
         );
  NAND3_X1 U10266 ( .A1(n8984), .A2(n8983), .A3(n8982), .ZN(P1_U3228) );
  XOR2_X1 U10267 ( .A(n8985), .B(n8986), .Z(n8992) );
  INV_X1 U10268 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8987) );
  OAI22_X1 U10269 ( .A1(n9035), .A2(n9041), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8987), .ZN(n8990) );
  INV_X1 U10270 ( .A(n9297), .ZN(n8988) );
  OAI22_X1 U10271 ( .A1(n8988), .A2(n9008), .B1(n9032), .B2(n9124), .ZN(n8989)
         );
  AOI211_X1 U10272 ( .C1(n9414), .C2(n9038), .A(n8990), .B(n8989), .ZN(n8991)
         );
  OAI21_X1 U10273 ( .B1(n8992), .B2(n9012), .A(n8991), .ZN(P1_U3231) );
  INV_X1 U10274 ( .A(n8993), .ZN(n8997) );
  NAND2_X1 U10275 ( .A1(n4310), .A2(n4339), .ZN(n8995) );
  AOI22_X1 U10276 ( .A1(n8997), .A2(n8996), .B1(n8995), .B2(n8994), .ZN(n9003)
         );
  INV_X1 U10277 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8998) );
  OAI22_X1 U10278 ( .A1(n9032), .A2(n9041), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8998), .ZN(n9001) );
  OAI22_X1 U10279 ( .A1(n9008), .A2(n8999), .B1(n9035), .B2(n9131), .ZN(n9000)
         );
  AOI211_X1 U10280 ( .C1(n9404), .C2(n9038), .A(n9001), .B(n9000), .ZN(n9002)
         );
  OAI21_X1 U10281 ( .B1(n9003), .B2(n9012), .A(n9002), .ZN(P1_U3233) );
  XNOR2_X1 U10282 ( .A(n9005), .B(n9004), .ZN(n9006) );
  XNOR2_X1 U10283 ( .A(n9007), .B(n9006), .ZN(n9013) );
  NAND2_X1 U10284 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9085) );
  OAI21_X1 U10285 ( .B1(n9035), .B2(n9124), .A(n9085), .ZN(n9010) );
  OAI22_X1 U10286 ( .A1(n9008), .A2(n9325), .B1(n9032), .B2(n9121), .ZN(n9009)
         );
  AOI211_X1 U10287 ( .C1(n9423), .C2(n9038), .A(n9010), .B(n9009), .ZN(n9011)
         );
  OAI21_X1 U10288 ( .B1(n9013), .B2(n9012), .A(n9011), .ZN(P1_U3236) );
  INV_X1 U10289 ( .A(n9014), .ZN(n9015) );
  AND3_X1 U10290 ( .A1(n9017), .A2(n9016), .A3(n9015), .ZN(n9018) );
  OAI21_X1 U10291 ( .B1(n9018), .B2(n4371), .A(n5630), .ZN(n9028) );
  AOI21_X1 U10292 ( .B1(n9020), .B2(n9051), .A(n9019), .ZN(n9027) );
  AOI22_X1 U10293 ( .A1(n9022), .A2(n9049), .B1(n9033), .B2(n9021), .ZN(n9026)
         );
  AND2_X1 U10294 ( .A1(n9023), .A2(n9887), .ZN(n9861) );
  NAND2_X1 U10295 ( .A1(n9024), .A2(n9861), .ZN(n9025) );
  NAND4_X1 U10296 ( .A1(n9028), .A2(n9027), .A3(n9026), .A4(n9025), .ZN(
        P1_U3237) );
  OAI211_X1 U10297 ( .C1(n4354), .C2(n9030), .A(n9029), .B(n5630), .ZN(n9040)
         );
  OAI22_X1 U10298 ( .A1(n9032), .A2(n9135), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9031), .ZN(n9037) );
  NAND2_X1 U10299 ( .A1(n9033), .A2(n9215), .ZN(n9034) );
  OAI21_X1 U10300 ( .B1(n9035), .B2(n9139), .A(n9034), .ZN(n9036) );
  AOI211_X1 U10301 ( .C1(n9383), .C2(n9038), .A(n9037), .B(n9036), .ZN(n9039)
         );
  NAND2_X1 U10302 ( .A1(n9040), .A2(n9039), .ZN(P1_U3238) );
  MUX2_X1 U10303 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9165), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10304 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9188), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10305 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9166), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10306 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9211), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10307 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9203), .S(P1_U4006), .Z(
        P1_U3581) );
  INV_X1 U10308 ( .A(n9135), .ZN(n9244) );
  MUX2_X1 U10309 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9244), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10310 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9230), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10311 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9271), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10312 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9286), .S(P1_U4006), .Z(
        P1_U3577) );
  INV_X1 U10313 ( .A(n9041), .ZN(n9302) );
  MUX2_X1 U10314 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9302), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10315 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9312), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10316 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9334), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10317 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9350), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10318 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9333), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10319 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9348), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10320 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9042), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10321 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n7974), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10322 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9043), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10323 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9044), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10324 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9045), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10325 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9046), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10326 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9047), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10327 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9048), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10328 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9049), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10329 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9050), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10330 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9051), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10331 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9052), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10332 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9053), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10333 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9054), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10334 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6326), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10335 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6325), .S(P1_U4006), .Z(
        P1_U3555) );
  OAI21_X1 U10336 ( .B1(n9057), .B2(n9056), .A(n9055), .ZN(n9058) );
  NAND2_X1 U10337 ( .A1(n9058), .A2(n9798), .ZN(n9069) );
  NOR2_X1 U10338 ( .A1(n9060), .A2(n9059), .ZN(n9061) );
  AOI211_X1 U10339 ( .C1(P1_ADDR_REG_11__SCAN_IN), .C2(n9827), .A(n9062), .B(
        n9061), .ZN(n9068) );
  OAI21_X1 U10340 ( .B1(n9065), .B2(n9064), .A(n9063), .ZN(n9066) );
  NAND2_X1 U10341 ( .A1(n9066), .A2(n9823), .ZN(n9067) );
  NAND3_X1 U10342 ( .A1(n9069), .A2(n9068), .A3(n9067), .ZN(P1_U3252) );
  INV_X1 U10343 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9084) );
  INV_X1 U10344 ( .A(n9070), .ZN(n9076) );
  AOI21_X1 U10345 ( .B1(n9078), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9071), .ZN(
        n9074) );
  XNOR2_X1 U10346 ( .A(n9093), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9073) );
  NOR2_X1 U10347 ( .A1(n9074), .A2(n9073), .ZN(n9092) );
  AOI211_X1 U10348 ( .C1(n9074), .C2(n9073), .A(n9092), .B(n9072), .ZN(n9075)
         );
  AOI211_X1 U10349 ( .C1(n9825), .C2(n9093), .A(n9076), .B(n9075), .ZN(n9083)
         );
  AOI21_X1 U10350 ( .B1(n9078), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9077), .ZN(
        n9080) );
  XNOR2_X1 U10351 ( .A(n9093), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n9079) );
  NOR2_X1 U10352 ( .A1(n9080), .A2(n9079), .ZN(n9086) );
  AOI211_X1 U10353 ( .C1(n9080), .C2(n9079), .A(n9086), .B(n9817), .ZN(n9081)
         );
  INV_X1 U10354 ( .A(n9081), .ZN(n9082) );
  OAI211_X1 U10355 ( .C1(n9084), .C2(n9773), .A(n9083), .B(n9082), .ZN(
        P1_U3258) );
  INV_X1 U10356 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9099) );
  INV_X1 U10357 ( .A(n9085), .ZN(n9091) );
  NAND2_X1 U10358 ( .A1(n9103), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9087) );
  OAI21_X1 U10359 ( .B1(n9103), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9087), .ZN(
        n9088) );
  NOR2_X1 U10360 ( .A1(n9089), .A2(n9088), .ZN(n9100) );
  AOI211_X1 U10361 ( .C1(n9089), .C2(n9088), .A(n9100), .B(n9817), .ZN(n9090)
         );
  AOI211_X1 U10362 ( .C1(n9103), .C2(n9825), .A(n9091), .B(n9090), .ZN(n9098)
         );
  XOR2_X1 U10363 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9103), .Z(n9095) );
  AOI21_X1 U10364 ( .B1(n9093), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9092), .ZN(
        n9094) );
  NAND2_X1 U10365 ( .A1(n9095), .A2(n9094), .ZN(n9102) );
  OAI21_X1 U10366 ( .B1(n9095), .B2(n9094), .A(n9102), .ZN(n9096) );
  NAND2_X1 U10367 ( .A1(n9096), .A2(n9823), .ZN(n9097) );
  OAI211_X1 U10368 ( .C1(n9773), .C2(n9099), .A(n9098), .B(n9097), .ZN(
        P1_U3259) );
  XNOR2_X1 U10369 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9101), .ZN(n9108) );
  OAI21_X1 U10370 ( .B1(n9103), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9102), .ZN(
        n9105) );
  INV_X1 U10371 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9104) );
  XOR2_X1 U10372 ( .A(n9105), .B(n9104), .Z(n9106) );
  AOI22_X1 U10373 ( .A1(n9108), .A2(n9798), .B1(n9823), .B2(n9106), .ZN(n9111)
         );
  INV_X1 U10374 ( .A(n9106), .ZN(n9109) );
  NAND2_X1 U10375 ( .A1(n9113), .A2(n9169), .ZN(n9114) );
  XNOR2_X1 U10376 ( .A(n9114), .B(n9357), .ZN(n9359) );
  AOI21_X1 U10377 ( .B1(n9309), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9115), .ZN(
        n9117) );
  NAND2_X1 U10378 ( .A1(n9357), .A2(n9698), .ZN(n9116) );
  OAI211_X1 U10379 ( .C1(n9359), .C2(n9118), .A(n9117), .B(n9116), .ZN(
        P1_U3261) );
  NOR2_X1 U10380 ( .A1(n9428), .A2(n9333), .ZN(n9122) );
  NAND2_X1 U10381 ( .A1(n9419), .A2(n9334), .ZN(n9125) );
  AOI22_X1 U10382 ( .A1(n9308), .A2(n9125), .B1(n9124), .B2(n9123), .ZN(n9294)
         );
  NAND2_X1 U10383 ( .A1(n9294), .A2(n9126), .ZN(n9127) );
  OAI21_X1 U10384 ( .B1(n9128), .B2(n9299), .A(n9127), .ZN(n9279) );
  NAND2_X1 U10385 ( .A1(n9258), .A2(n9131), .ZN(n9132) );
  INV_X1 U10386 ( .A(n9379), .ZN(n9196) );
  NAND2_X1 U10387 ( .A1(n9178), .A2(n4821), .ZN(n9140) );
  XNOR2_X1 U10388 ( .A(n9140), .B(n9161), .ZN(n9364) );
  INV_X1 U10389 ( .A(n9364), .ZN(n9177) );
  INV_X1 U10390 ( .A(n9145), .ZN(n9146) );
  NOR2_X1 U10391 ( .A1(n9280), .A2(n9150), .ZN(n9269) );
  OAI21_X1 U10392 ( .B1(n9269), .B2(n9152), .A(n9151), .ZN(n9261) );
  NOR2_X1 U10393 ( .A1(n9261), .A2(n9262), .ZN(n9260) );
  INV_X1 U10394 ( .A(n9153), .ZN(n9154) );
  NOR2_X1 U10395 ( .A1(n9260), .A2(n9154), .ZN(n9243) );
  NOR2_X1 U10396 ( .A1(n9199), .A2(n9200), .ZN(n9198) );
  INV_X1 U10397 ( .A(n9158), .ZN(n9159) );
  NOR2_X1 U10398 ( .A1(n9198), .A2(n9159), .ZN(n9186) );
  NAND2_X1 U10399 ( .A1(n9186), .A2(n9187), .ZN(n9185) );
  NAND2_X1 U10400 ( .A1(n9185), .A2(n9160), .ZN(n9163) );
  INV_X1 U10401 ( .A(n9161), .ZN(n9162) );
  XNOR2_X1 U10402 ( .A(n9163), .B(n9162), .ZN(n9168) );
  AOI22_X1 U10403 ( .A1(n9166), .A2(n9347), .B1(n9165), .B2(n9164), .ZN(n9167)
         );
  OAI21_X1 U10404 ( .B1(n9168), .B2(n9716), .A(n9167), .ZN(n9365) );
  INV_X1 U10405 ( .A(n9181), .ZN(n9170) );
  AOI211_X1 U10406 ( .C1(n9366), .C2(n9170), .A(n9854), .B(n9169), .ZN(n9368)
         );
  NAND2_X1 U10407 ( .A1(n9368), .A2(n9306), .ZN(n9173) );
  AOI22_X1 U10408 ( .A1(n9309), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9171), .B2(
        n9720), .ZN(n9172) );
  OAI211_X1 U10409 ( .C1(n9174), .C2(n9723), .A(n9173), .B(n9172), .ZN(n9175)
         );
  AOI21_X1 U10410 ( .B1(n9365), .B2(n9725), .A(n9175), .ZN(n9176) );
  OAI21_X1 U10411 ( .B1(n9177), .B2(n9356), .A(n9176), .ZN(P1_U3355) );
  OAI21_X1 U10412 ( .B1(n9180), .B2(n9179), .A(n9178), .ZN(n9377) );
  AOI21_X1 U10413 ( .B1(n9373), .B2(n9192), .A(n9181), .ZN(n9374) );
  AOI22_X1 U10414 ( .A1(n9309), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9182), .B2(
        n9720), .ZN(n9183) );
  OAI21_X1 U10415 ( .B1(n9184), .B2(n9723), .A(n9183), .ZN(n9190) );
  OAI21_X1 U10416 ( .B1(n9187), .B2(n9186), .A(n9185), .ZN(n9189) );
  XOR2_X1 U10417 ( .A(n9191), .B(n9200), .Z(n9382) );
  INV_X1 U10418 ( .A(n9192), .ZN(n9193) );
  AOI211_X1 U10419 ( .C1(n9379), .C2(n9213), .A(n9854), .B(n9193), .ZN(n9378)
         );
  AOI22_X1 U10420 ( .A1(n9309), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9194), .B2(
        n9720), .ZN(n9195) );
  OAI21_X1 U10421 ( .B1(n9196), .B2(n9723), .A(n9195), .ZN(n9205) );
  NOR2_X1 U10422 ( .A1(n9197), .A2(n9710), .ZN(n9202) );
  AOI211_X1 U10423 ( .C1(n9200), .C2(n9199), .A(n9716), .B(n9198), .ZN(n9201)
         );
  AOI211_X1 U10424 ( .C1(n9347), .C2(n9203), .A(n9202), .B(n9201), .ZN(n9381)
         );
  NOR2_X1 U10425 ( .A1(n9381), .A2(n9309), .ZN(n9204) );
  AOI211_X1 U10426 ( .C1(n9306), .C2(n9378), .A(n9205), .B(n9204), .ZN(n9206)
         );
  OAI21_X1 U10427 ( .B1(n9382), .B2(n9356), .A(n9206), .ZN(P1_U3264) );
  XNOR2_X1 U10428 ( .A(n9207), .B(n9210), .ZN(n9387) );
  NOR2_X1 U10429 ( .A1(n9225), .A2(n9208), .ZN(n9209) );
  XOR2_X1 U10430 ( .A(n9210), .B(n9209), .Z(n9212) );
  AOI222_X1 U10431 ( .A1(n9352), .A2(n9212), .B1(n9211), .B2(n9349), .C1(n9244), .C2(n9347), .ZN(n9386) );
  INV_X1 U10432 ( .A(n9386), .ZN(n9220) );
  INV_X1 U10433 ( .A(n9383), .ZN(n9218) );
  INV_X1 U10434 ( .A(n9213), .ZN(n9214) );
  AOI21_X1 U10435 ( .B1(n9383), .B2(n9231), .A(n9214), .ZN(n9384) );
  NAND2_X1 U10436 ( .A1(n9384), .A2(n9706), .ZN(n9217) );
  AOI22_X1 U10437 ( .A1(n9309), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9215), .B2(
        n9720), .ZN(n9216) );
  OAI211_X1 U10438 ( .C1(n9218), .C2(n9723), .A(n9217), .B(n9216), .ZN(n9219)
         );
  AOI21_X1 U10439 ( .B1(n9220), .B2(n9725), .A(n9219), .ZN(n9221) );
  OAI21_X1 U10440 ( .B1(n9387), .B2(n9356), .A(n9221), .ZN(P1_U3265) );
  XOR2_X1 U10441 ( .A(n9227), .B(n9222), .Z(n9392) );
  NOR2_X1 U10442 ( .A1(n9223), .A2(n9723), .ZN(n9237) );
  NOR2_X1 U10443 ( .A1(n9224), .A2(n9710), .ZN(n9229) );
  AOI211_X1 U10444 ( .C1(n9227), .C2(n9226), .A(n9716), .B(n9225), .ZN(n9228)
         );
  AOI211_X1 U10445 ( .C1(n9347), .C2(n9230), .A(n9229), .B(n9228), .ZN(n9391)
         );
  INV_X1 U10446 ( .A(n9246), .ZN(n9233) );
  INV_X1 U10447 ( .A(n9231), .ZN(n9232) );
  AOI211_X1 U10448 ( .C1(n9389), .C2(n9233), .A(n9854), .B(n9232), .ZN(n9388)
         );
  AOI22_X1 U10449 ( .A1(n9388), .A2(n7099), .B1(n9720), .B2(n9234), .ZN(n9235)
         );
  AOI21_X1 U10450 ( .B1(n9391), .B2(n9235), .A(n9309), .ZN(n9236) );
  AOI211_X1 U10451 ( .C1(n9309), .C2(P1_REG2_REG_25__SCAN_IN), .A(n9237), .B(
        n9236), .ZN(n9238) );
  OAI21_X1 U10452 ( .B1(n9392), .B2(n9356), .A(n9238), .ZN(P1_U3266) );
  XNOR2_X1 U10453 ( .A(n9239), .B(n9242), .ZN(n9397) );
  NOR2_X1 U10454 ( .A1(n9240), .A2(n9723), .ZN(n9251) );
  OAI21_X1 U10455 ( .B1(n9243), .B2(n9242), .A(n9241), .ZN(n9245) );
  AOI222_X1 U10456 ( .A1(n9352), .A2(n9245), .B1(n9244), .B2(n9349), .C1(n9271), .C2(n9347), .ZN(n9396) );
  INV_X1 U10457 ( .A(n9254), .ZN(n9247) );
  AOI211_X1 U10458 ( .C1(n9394), .C2(n9247), .A(n9854), .B(n9246), .ZN(n9393)
         );
  AOI22_X1 U10459 ( .A1(n9393), .A2(n7099), .B1(n9720), .B2(n9248), .ZN(n9249)
         );
  AOI21_X1 U10460 ( .B1(n9396), .B2(n9249), .A(n9309), .ZN(n9250) );
  AOI211_X1 U10461 ( .C1(n9309), .C2(P1_REG2_REG_24__SCAN_IN), .A(n9251), .B(
        n9250), .ZN(n9252) );
  OAI21_X1 U10462 ( .B1(n9397), .B2(n9356), .A(n9252), .ZN(P1_U3267) );
  XNOR2_X1 U10463 ( .A(n9253), .B(n9262), .ZN(n9402) );
  INV_X1 U10464 ( .A(n9273), .ZN(n9255) );
  AOI211_X1 U10465 ( .C1(n9399), .C2(n9255), .A(n9854), .B(n9254), .ZN(n9398)
         );
  AOI22_X1 U10466 ( .A1(n9309), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9256), .B2(
        n9720), .ZN(n9257) );
  OAI21_X1 U10467 ( .B1(n9258), .B2(n9723), .A(n9257), .ZN(n9266) );
  NOR2_X1 U10468 ( .A1(n9259), .A2(n9710), .ZN(n9264) );
  AOI211_X1 U10469 ( .C1(n9262), .C2(n9261), .A(n9716), .B(n9260), .ZN(n9263)
         );
  AOI211_X1 U10470 ( .C1(n9347), .C2(n9286), .A(n9264), .B(n9263), .ZN(n9401)
         );
  NOR2_X1 U10471 ( .A1(n9401), .A2(n9309), .ZN(n9265) );
  AOI211_X1 U10472 ( .C1(n9398), .C2(n9306), .A(n9266), .B(n9265), .ZN(n9267)
         );
  OAI21_X1 U10473 ( .B1(n9402), .B2(n9356), .A(n9267), .ZN(P1_U3268) );
  XNOR2_X1 U10474 ( .A(n4343), .B(n9270), .ZN(n9407) );
  NOR2_X1 U10475 ( .A1(n9268), .A2(n9723), .ZN(n9277) );
  XOR2_X1 U10476 ( .A(n9270), .B(n9269), .Z(n9272) );
  AOI222_X1 U10477 ( .A1(n9352), .A2(n9272), .B1(n9271), .B2(n9349), .C1(n9302), .C2(n9347), .ZN(n9406) );
  AOI211_X1 U10478 ( .C1(n9404), .C2(n9288), .A(n9854), .B(n9273), .ZN(n9403)
         );
  AOI22_X1 U10479 ( .A1(n9403), .A2(n7099), .B1(n9720), .B2(n9274), .ZN(n9275)
         );
  AOI21_X1 U10480 ( .B1(n9406), .B2(n9275), .A(n9309), .ZN(n9276) );
  AOI211_X1 U10481 ( .C1(n9309), .C2(P1_REG2_REG_22__SCAN_IN), .A(n9277), .B(
        n9276), .ZN(n9278) );
  OAI21_X1 U10482 ( .B1(n9407), .B2(n9356), .A(n9278), .ZN(P1_U3269) );
  XNOR2_X1 U10483 ( .A(n9279), .B(n9281), .ZN(n9412) );
  AOI22_X1 U10484 ( .A1(n9409), .A2(n9698), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9309), .ZN(n9293) );
  INV_X1 U10485 ( .A(n9280), .ZN(n9285) );
  OAI21_X1 U10486 ( .B1(n9283), .B2(n9282), .A(n9281), .ZN(n9284) );
  NAND2_X1 U10487 ( .A1(n9285), .A2(n9284), .ZN(n9287) );
  AOI222_X1 U10488 ( .A1(n9352), .A2(n9287), .B1(n9286), .B2(n9349), .C1(n9312), .C2(n9347), .ZN(n9411) );
  AOI211_X1 U10489 ( .C1(n9409), .C2(n9295), .A(n9854), .B(n4669), .ZN(n9408)
         );
  AOI22_X1 U10490 ( .A1(n9408), .A2(n7099), .B1(n9720), .B2(n9289), .ZN(n9290)
         );
  AOI21_X1 U10491 ( .B1(n9411), .B2(n9290), .A(n9309), .ZN(n9291) );
  INV_X1 U10492 ( .A(n9291), .ZN(n9292) );
  OAI211_X1 U10493 ( .C1(n9412), .C2(n9356), .A(n9293), .B(n9292), .ZN(
        P1_U3270) );
  XOR2_X1 U10494 ( .A(n9294), .B(n9300), .Z(n9417) );
  INV_X1 U10495 ( .A(n9295), .ZN(n9296) );
  AOI211_X1 U10496 ( .C1(n9414), .C2(n9314), .A(n9854), .B(n9296), .ZN(n9413)
         );
  AOI22_X1 U10497 ( .A1(n9309), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9297), .B2(
        n9720), .ZN(n9298) );
  OAI21_X1 U10498 ( .B1(n9299), .B2(n9723), .A(n9298), .ZN(n9305) );
  XNOR2_X1 U10499 ( .A(n9301), .B(n9300), .ZN(n9303) );
  AOI222_X1 U10500 ( .A1(n9352), .A2(n9303), .B1(n9302), .B2(n9349), .C1(n9334), .C2(n9347), .ZN(n9416) );
  NOR2_X1 U10501 ( .A1(n9416), .A2(n9309), .ZN(n9304) );
  AOI211_X1 U10502 ( .C1(n9413), .C2(n9306), .A(n9305), .B(n9304), .ZN(n9307)
         );
  OAI21_X1 U10503 ( .B1(n9417), .B2(n9356), .A(n9307), .ZN(P1_U3271) );
  XOR2_X1 U10504 ( .A(n9308), .B(n9310), .Z(n9422) );
  AOI22_X1 U10505 ( .A1(n9419), .A2(n9698), .B1(P1_REG2_REG_19__SCAN_IN), .B2(
        n9309), .ZN(n9321) );
  XNOR2_X1 U10506 ( .A(n9311), .B(n9310), .ZN(n9313) );
  AOI222_X1 U10507 ( .A1(n9352), .A2(n9313), .B1(n9312), .B2(n9349), .C1(n9350), .C2(n9347), .ZN(n9421) );
  INV_X1 U10508 ( .A(n9323), .ZN(n9316) );
  INV_X1 U10509 ( .A(n9314), .ZN(n9315) );
  AOI211_X1 U10510 ( .C1(n9419), .C2(n9316), .A(n9854), .B(n9315), .ZN(n9418)
         );
  NAND2_X1 U10511 ( .A1(n9418), .A2(n7099), .ZN(n9317) );
  OAI211_X1 U10512 ( .C1(n9685), .C2(n9318), .A(n9421), .B(n9317), .ZN(n9319)
         );
  NAND2_X1 U10513 ( .A1(n9319), .A2(n9725), .ZN(n9320) );
  OAI211_X1 U10514 ( .C1(n9422), .C2(n9356), .A(n9321), .B(n9320), .ZN(
        P1_U3272) );
  XNOR2_X1 U10515 ( .A(n9322), .B(n9331), .ZN(n9427) );
  INV_X1 U10516 ( .A(n9341), .ZN(n9324) );
  AOI21_X1 U10517 ( .B1(n9423), .B2(n9324), .A(n9323), .ZN(n9424) );
  INV_X1 U10518 ( .A(n9325), .ZN(n9326) );
  AOI22_X1 U10519 ( .A1(n9309), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9326), .B2(
        n9720), .ZN(n9327) );
  OAI21_X1 U10520 ( .B1(n9328), .B2(n9723), .A(n9327), .ZN(n9337) );
  NAND2_X1 U10521 ( .A1(n9330), .A2(n9329), .ZN(n9332) );
  XNOR2_X1 U10522 ( .A(n9332), .B(n9331), .ZN(n9335) );
  AOI222_X1 U10523 ( .A1(n9352), .A2(n9335), .B1(n9334), .B2(n9349), .C1(n9333), .C2(n9347), .ZN(n9426) );
  NOR2_X1 U10524 ( .A1(n9426), .A2(n9309), .ZN(n9336) );
  AOI211_X1 U10525 ( .C1(n9424), .C2(n9706), .A(n9337), .B(n9336), .ZN(n9338)
         );
  OAI21_X1 U10526 ( .B1(n9427), .B2(n9356), .A(n9338), .ZN(P1_U3273) );
  XNOR2_X1 U10527 ( .A(n9340), .B(n9339), .ZN(n9432) );
  AOI21_X1 U10528 ( .B1(n9428), .B2(n9342), .A(n9341), .ZN(n9429) );
  AOI22_X1 U10529 ( .A1(n9309), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9343), .B2(
        n9720), .ZN(n9344) );
  OAI21_X1 U10530 ( .B1(n4674), .B2(n9723), .A(n9344), .ZN(n9354) );
  XNOR2_X1 U10531 ( .A(n9346), .B(n9345), .ZN(n9351) );
  AOI222_X1 U10532 ( .A1(n9352), .A2(n9351), .B1(n9350), .B2(n9349), .C1(n9348), .C2(n9347), .ZN(n9431) );
  NOR2_X1 U10533 ( .A1(n9431), .A2(n9309), .ZN(n9353) );
  AOI211_X1 U10534 ( .C1(n9429), .C2(n9706), .A(n9354), .B(n9353), .ZN(n9355)
         );
  OAI21_X1 U10535 ( .B1(n9432), .B2(n9356), .A(n9355), .ZN(P1_U3274) );
  NAND2_X1 U10536 ( .A1(n9357), .A2(n9887), .ZN(n9358) );
  OAI211_X1 U10537 ( .C1(n9359), .C2(n9854), .A(n9358), .B(n9362), .ZN(n9449)
         );
  MUX2_X1 U10538 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9449), .S(n9911), .Z(
        P1_U3554) );
  NAND2_X1 U10539 ( .A1(n9360), .A2(n9887), .ZN(n9361) );
  OAI211_X1 U10540 ( .C1(n9363), .C2(n9854), .A(n9362), .B(n9361), .ZN(n9450)
         );
  MUX2_X1 U10541 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9450), .S(n9911), .Z(
        P1_U3553) );
  NAND2_X1 U10542 ( .A1(n9364), .A2(n9873), .ZN(n9372) );
  NAND2_X1 U10543 ( .A1(n9372), .A2(n9371), .ZN(n9629) );
  MUX2_X1 U10544 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9629), .S(n9911), .Z(
        P1_U3552) );
  AOI22_X1 U10545 ( .A1(n9374), .A2(n9888), .B1(n9887), .B2(n9373), .ZN(n9375)
         );
  OAI211_X1 U10546 ( .C1(n9377), .C2(n9892), .A(n9376), .B(n9375), .ZN(n9630)
         );
  MUX2_X1 U10547 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9630), .S(n9911), .Z(
        P1_U3551) );
  AOI21_X1 U10548 ( .B1(n9887), .B2(n9379), .A(n9378), .ZN(n9380) );
  OAI211_X1 U10549 ( .C1(n9382), .C2(n9892), .A(n9381), .B(n9380), .ZN(n9631)
         );
  MUX2_X1 U10550 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9631), .S(n9911), .Z(
        P1_U3550) );
  AOI22_X1 U10551 ( .A1(n9384), .A2(n9888), .B1(n9887), .B2(n9383), .ZN(n9385)
         );
  OAI211_X1 U10552 ( .C1(n9387), .C2(n9892), .A(n9386), .B(n9385), .ZN(n9632)
         );
  MUX2_X1 U10553 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9632), .S(n9911), .Z(
        P1_U3549) );
  AOI21_X1 U10554 ( .B1(n9887), .B2(n9389), .A(n9388), .ZN(n9390) );
  OAI211_X1 U10555 ( .C1(n9392), .C2(n9892), .A(n9391), .B(n9390), .ZN(n9633)
         );
  MUX2_X1 U10556 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9633), .S(n9911), .Z(
        P1_U3548) );
  AOI21_X1 U10557 ( .B1(n9887), .B2(n9394), .A(n9393), .ZN(n9395) );
  OAI211_X1 U10558 ( .C1(n9397), .C2(n9892), .A(n9396), .B(n9395), .ZN(n9634)
         );
  MUX2_X1 U10559 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9634), .S(n9911), .Z(
        P1_U3547) );
  AOI21_X1 U10560 ( .B1(n9887), .B2(n9399), .A(n9398), .ZN(n9400) );
  OAI211_X1 U10561 ( .C1(n9402), .C2(n9892), .A(n9401), .B(n9400), .ZN(n9635)
         );
  MUX2_X1 U10562 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9635), .S(n9911), .Z(
        P1_U3546) );
  AOI21_X1 U10563 ( .B1(n9887), .B2(n9404), .A(n9403), .ZN(n9405) );
  OAI211_X1 U10564 ( .C1(n9407), .C2(n9892), .A(n9406), .B(n9405), .ZN(n9636)
         );
  MUX2_X1 U10565 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9636), .S(n9911), .Z(
        P1_U3545) );
  AOI21_X1 U10566 ( .B1(n9887), .B2(n9409), .A(n9408), .ZN(n9410) );
  OAI211_X1 U10567 ( .C1(n9412), .C2(n9892), .A(n9411), .B(n9410), .ZN(n9637)
         );
  MUX2_X1 U10568 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9637), .S(n9911), .Z(
        P1_U3544) );
  AOI21_X1 U10569 ( .B1(n9887), .B2(n9414), .A(n9413), .ZN(n9415) );
  OAI211_X1 U10570 ( .C1(n9417), .C2(n9892), .A(n9416), .B(n9415), .ZN(n9638)
         );
  MUX2_X1 U10571 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9638), .S(n9911), .Z(
        P1_U3543) );
  AOI21_X1 U10572 ( .B1(n9887), .B2(n9419), .A(n9418), .ZN(n9420) );
  OAI211_X1 U10573 ( .C1(n9422), .C2(n9892), .A(n9421), .B(n9420), .ZN(n9639)
         );
  MUX2_X1 U10574 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9639), .S(n9911), .Z(
        P1_U3542) );
  AOI22_X1 U10575 ( .A1(n9424), .A2(n9888), .B1(n9887), .B2(n9423), .ZN(n9425)
         );
  OAI211_X1 U10576 ( .C1(n9427), .C2(n9892), .A(n9426), .B(n9425), .ZN(n9640)
         );
  MUX2_X1 U10577 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9640), .S(n9911), .Z(
        P1_U3541) );
  AOI22_X1 U10578 ( .A1(n9429), .A2(n9888), .B1(n9887), .B2(n9428), .ZN(n9430)
         );
  OAI211_X1 U10579 ( .C1(n9432), .C2(n9892), .A(n9431), .B(n9430), .ZN(n9641)
         );
  MUX2_X1 U10580 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9641), .S(n9911), .Z(
        P1_U3540) );
  NAND3_X1 U10581 ( .A1(n4597), .A2(n9873), .A3(n9433), .ZN(n9438) );
  INV_X1 U10582 ( .A(n9434), .ZN(n9436) );
  NAND4_X1 U10583 ( .A1(n9438), .A2(n9437), .A3(n9436), .A4(n9435), .ZN(n9642)
         );
  MUX2_X1 U10584 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9642), .S(n9911), .Z(
        P1_U3539) );
  INV_X1 U10585 ( .A(n9884), .ZN(n9673) );
  AOI22_X1 U10586 ( .A1(n9440), .A2(n9888), .B1(n9887), .B2(n9439), .ZN(n9441)
         );
  OAI211_X1 U10587 ( .C1(n9673), .C2(n9443), .A(n9442), .B(n9441), .ZN(n9643)
         );
  MUX2_X1 U10588 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9643), .S(n9911), .Z(
        P1_U3538) );
  AOI21_X1 U10589 ( .B1(n9887), .B2(n9445), .A(n9444), .ZN(n9446) );
  OAI211_X1 U10590 ( .C1(n9448), .C2(n9892), .A(n9447), .B(n9446), .ZN(n9644)
         );
  MUX2_X1 U10591 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9644), .S(n9911), .Z(
        P1_U3537) );
  MUX2_X1 U10592 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9449), .S(n9897), .Z(
        P1_U3522) );
  MUX2_X1 U10593 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9450), .S(n9897), .Z(n9628) );
  OAI22_X1 U10594 ( .A1(P1_D_REG_21__SCAN_IN), .A2(keyinput104), .B1(
        keyinput95), .B2(P2_REG3_REG_15__SCAN_IN), .ZN(n9451) );
  AOI221_X1 U10595 ( .B1(P1_D_REG_21__SCAN_IN), .B2(keyinput104), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput95), .A(n9451), .ZN(n9458) );
  OAI22_X1 U10596 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(keyinput98), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(keyinput86), .ZN(n9452) );
  AOI221_X1 U10597 ( .B1(P2_IR_REG_15__SCAN_IN), .B2(keyinput98), .C1(
        keyinput86), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n9452), .ZN(n9457) );
  OAI22_X1 U10598 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(keyinput68), .B1(keyinput76), .B2(P2_REG2_REG_23__SCAN_IN), .ZN(n9453) );
  AOI221_X1 U10599 ( .B1(P2_IR_REG_7__SCAN_IN), .B2(keyinput68), .C1(
        P2_REG2_REG_23__SCAN_IN), .C2(keyinput76), .A(n9453), .ZN(n9456) );
  OAI22_X1 U10600 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(keyinput121), .B1(
        keyinput120), .B2(P2_D_REG_4__SCAN_IN), .ZN(n9454) );
  AOI221_X1 U10601 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(keyinput121), .C1(
        P2_D_REG_4__SCAN_IN), .C2(keyinput120), .A(n9454), .ZN(n9455) );
  NAND4_X1 U10602 ( .A1(n9458), .A2(n9457), .A3(n9456), .A4(n9455), .ZN(n9486)
         );
  OAI22_X1 U10603 ( .A1(P1_STATE_REG_SCAN_IN), .A2(keyinput66), .B1(
        keyinput118), .B2(P2_REG0_REG_30__SCAN_IN), .ZN(n9459) );
  AOI221_X1 U10604 ( .B1(P1_STATE_REG_SCAN_IN), .B2(keyinput66), .C1(
        P2_REG0_REG_30__SCAN_IN), .C2(keyinput118), .A(n9459), .ZN(n9466) );
  OAI22_X1 U10605 ( .A1(P2_REG1_REG_5__SCAN_IN), .A2(keyinput103), .B1(
        keyinput84), .B2(P2_REG1_REG_3__SCAN_IN), .ZN(n9460) );
  AOI221_X1 U10606 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(keyinput103), .C1(
        P2_REG1_REG_3__SCAN_IN), .C2(keyinput84), .A(n9460), .ZN(n9465) );
  OAI22_X1 U10607 ( .A1(SI_9_), .A2(keyinput64), .B1(keyinput113), .B2(
        P1_ADDR_REG_11__SCAN_IN), .ZN(n9461) );
  AOI221_X1 U10608 ( .B1(SI_9_), .B2(keyinput64), .C1(P1_ADDR_REG_11__SCAN_IN), 
        .C2(keyinput113), .A(n9461), .ZN(n9464) );
  OAI22_X1 U10609 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(keyinput78), .B1(
        P2_ADDR_REG_0__SCAN_IN), .B2(keyinput99), .ZN(n9462) );
  AOI221_X1 U10610 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(keyinput78), .C1(
        keyinput99), .C2(P2_ADDR_REG_0__SCAN_IN), .A(n9462), .ZN(n9463) );
  NAND4_X1 U10611 ( .A1(n9466), .A2(n9465), .A3(n9464), .A4(n9463), .ZN(n9485)
         );
  OAI22_X1 U10612 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(keyinput90), .B1(
        P2_ADDR_REG_12__SCAN_IN), .B2(keyinput77), .ZN(n9467) );
  AOI221_X1 U10613 ( .B1(P1_REG3_REG_8__SCAN_IN), .B2(keyinput90), .C1(
        keyinput77), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n9467), .ZN(n9474) );
  OAI22_X1 U10614 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(keyinput65), .B1(
        keyinput119), .B2(P2_REG1_REG_7__SCAN_IN), .ZN(n9468) );
  AOI221_X1 U10615 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(keyinput65), .C1(
        P2_REG1_REG_7__SCAN_IN), .C2(keyinput119), .A(n9468), .ZN(n9473) );
  OAI22_X1 U10616 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(keyinput74), .B1(
        keyinput70), .B2(P1_REG2_REG_6__SCAN_IN), .ZN(n9469) );
  AOI221_X1 U10617 ( .B1(P2_DATAO_REG_18__SCAN_IN), .B2(keyinput74), .C1(
        P1_REG2_REG_6__SCAN_IN), .C2(keyinput70), .A(n9469), .ZN(n9472) );
  OAI22_X1 U10618 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput75), .B1(
        keyinput85), .B2(P1_REG1_REG_28__SCAN_IN), .ZN(n9470) );
  AOI221_X1 U10619 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput75), .C1(
        P1_REG1_REG_28__SCAN_IN), .C2(keyinput85), .A(n9470), .ZN(n9471) );
  NAND4_X1 U10620 ( .A1(n9474), .A2(n9473), .A3(n9472), .A4(n9471), .ZN(n9484)
         );
  OAI22_X1 U10621 ( .A1(P1_REG2_REG_29__SCAN_IN), .A2(keyinput108), .B1(
        keyinput83), .B2(P2_D_REG_2__SCAN_IN), .ZN(n9475) );
  AOI221_X1 U10622 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(keyinput108), .C1(
        P2_D_REG_2__SCAN_IN), .C2(keyinput83), .A(n9475), .ZN(n9482) );
  OAI22_X1 U10623 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(keyinput69), .B1(
        P2_REG1_REG_6__SCAN_IN), .B2(keyinput82), .ZN(n9476) );
  AOI221_X1 U10624 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(keyinput69), .C1(
        keyinput82), .C2(P2_REG1_REG_6__SCAN_IN), .A(n9476), .ZN(n9481) );
  OAI22_X1 U10625 ( .A1(P2_D_REG_13__SCAN_IN), .A2(keyinput80), .B1(
        P2_REG2_REG_21__SCAN_IN), .B2(keyinput106), .ZN(n9477) );
  AOI221_X1 U10626 ( .B1(P2_D_REG_13__SCAN_IN), .B2(keyinput80), .C1(
        keyinput106), .C2(P2_REG2_REG_21__SCAN_IN), .A(n9477), .ZN(n9480) );
  OAI22_X1 U10627 ( .A1(SI_12_), .A2(keyinput72), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(keyinput89), .ZN(n9478) );
  AOI221_X1 U10628 ( .B1(SI_12_), .B2(keyinput72), .C1(keyinput89), .C2(
        P2_REG3_REG_28__SCAN_IN), .A(n9478), .ZN(n9479) );
  NAND4_X1 U10629 ( .A1(n9482), .A2(n9481), .A3(n9480), .A4(n9479), .ZN(n9483)
         );
  NOR4_X1 U10630 ( .A1(n9486), .A2(n9485), .A3(n9484), .A4(n9483), .ZN(n9535)
         );
  AOI22_X1 U10631 ( .A1(n9488), .A2(keyinput109), .B1(keyinput111), .B2(n9583), 
        .ZN(n9487) );
  OAI221_X1 U10632 ( .B1(n9488), .B2(keyinput109), .C1(n9583), .C2(keyinput111), .A(n9487), .ZN(n9498) );
  INV_X1 U10633 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n9929) );
  INV_X1 U10634 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9833) );
  AOI22_X1 U10635 ( .A1(n9929), .A2(keyinput116), .B1(n9833), .B2(keyinput87), 
        .ZN(n9489) );
  OAI221_X1 U10636 ( .B1(n9929), .B2(keyinput116), .C1(n9833), .C2(keyinput87), 
        .A(n9489), .ZN(n9497) );
  INV_X1 U10637 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9928) );
  AOI22_X1 U10638 ( .A1(n9928), .A2(keyinput91), .B1(keyinput67), .B2(n9491), 
        .ZN(n9490) );
  OAI221_X1 U10639 ( .B1(n9928), .B2(keyinput91), .C1(n9491), .C2(keyinput67), 
        .A(n9490), .ZN(n9496) );
  INV_X1 U10640 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9494) );
  INV_X1 U10641 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9493) );
  AOI22_X1 U10642 ( .A1(n9494), .A2(keyinput81), .B1(n9493), .B2(keyinput125), 
        .ZN(n9492) );
  OAI221_X1 U10643 ( .B1(n9494), .B2(keyinput81), .C1(n9493), .C2(keyinput125), 
        .A(n9492), .ZN(n9495) );
  NOR4_X1 U10644 ( .A1(n9498), .A2(n9497), .A3(n9496), .A4(n9495), .ZN(n9534)
         );
  AOI22_X1 U10645 ( .A1(n6983), .A2(keyinput122), .B1(keyinput123), .B2(n7568), 
        .ZN(n9499) );
  OAI221_X1 U10646 ( .B1(n6983), .B2(keyinput122), .C1(n7568), .C2(keyinput123), .A(n9499), .ZN(n9506) );
  INV_X1 U10647 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n9927) );
  AOI22_X1 U10648 ( .A1(n9927), .A2(keyinput88), .B1(n9501), .B2(keyinput102), 
        .ZN(n9500) );
  OAI221_X1 U10649 ( .B1(n9927), .B2(keyinput88), .C1(n9501), .C2(keyinput102), 
        .A(n9500), .ZN(n9505) );
  INV_X1 U10650 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9604) );
  AOI22_X1 U10651 ( .A1(n9604), .A2(keyinput92), .B1(keyinput79), .B2(n9503), 
        .ZN(n9502) );
  OAI221_X1 U10652 ( .B1(n9604), .B2(keyinput92), .C1(n9503), .C2(keyinput79), 
        .A(n9502), .ZN(n9504) );
  NOR3_X1 U10653 ( .A1(n9506), .A2(n9505), .A3(n9504), .ZN(n9532) );
  XNOR2_X1 U10654 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput117), .ZN(n9510) );
  XNOR2_X1 U10655 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(keyinput112), .ZN(n9509)
         );
  XNOR2_X1 U10656 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput110), .ZN(n9508)
         );
  XNOR2_X1 U10657 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput126), .ZN(n9507) );
  NAND4_X1 U10658 ( .A1(n9510), .A2(n9509), .A3(n9508), .A4(n9507), .ZN(n9516)
         );
  XNOR2_X1 U10659 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput107), .ZN(n9514) );
  XNOR2_X1 U10660 ( .A(P2_IR_REG_2__SCAN_IN), .B(keyinput94), .ZN(n9513) );
  XNOR2_X1 U10661 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput101), .ZN(n9512) );
  XNOR2_X1 U10662 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput73), .ZN(n9511) );
  NAND4_X1 U10663 ( .A1(n9514), .A2(n9513), .A3(n9512), .A4(n9511), .ZN(n9515)
         );
  NOR2_X1 U10664 ( .A1(n9516), .A2(n9515), .ZN(n9531) );
  AOI22_X1 U10665 ( .A1(n5720), .A2(keyinput114), .B1(n9586), .B2(keyinput105), 
        .ZN(n9517) );
  OAI221_X1 U10666 ( .B1(n5720), .B2(keyinput114), .C1(n9586), .C2(keyinput105), .A(n9517), .ZN(n9523) );
  XNOR2_X1 U10667 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput124), .ZN(n9521) );
  XNOR2_X1 U10668 ( .A(SI_19_), .B(keyinput115), .ZN(n9520) );
  XNOR2_X1 U10669 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput97), .ZN(n9519) );
  XNOR2_X1 U10670 ( .A(P1_REG1_REG_15__SCAN_IN), .B(keyinput96), .ZN(n9518) );
  NAND4_X1 U10671 ( .A1(n9521), .A2(n9520), .A3(n9519), .A4(n9518), .ZN(n9522)
         );
  NOR2_X1 U10672 ( .A1(n9523), .A2(n9522), .ZN(n9530) );
  AOI22_X1 U10673 ( .A1(n9602), .A2(keyinput127), .B1(keyinput93), .B2(n6028), 
        .ZN(n9524) );
  OAI221_X1 U10674 ( .B1(n9602), .B2(keyinput127), .C1(n6028), .C2(keyinput93), 
        .A(n9524), .ZN(n9528) );
  AOI22_X1 U10675 ( .A1(n5750), .A2(keyinput100), .B1(n9526), .B2(keyinput71), 
        .ZN(n9525) );
  OAI221_X1 U10676 ( .B1(n5750), .B2(keyinput100), .C1(n9526), .C2(keyinput71), 
        .A(n9525), .ZN(n9527) );
  NOR2_X1 U10677 ( .A1(n9528), .A2(n9527), .ZN(n9529) );
  AND4_X1 U10678 ( .A1(n9532), .A2(n9531), .A3(n9530), .A4(n9529), .ZN(n9533)
         );
  NAND3_X1 U10679 ( .A1(n9535), .A2(n9534), .A3(n9533), .ZN(n9626) );
  AOI22_X1 U10680 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput53), .B1(SI_12_), 
        .B2(keyinput8), .ZN(n9536) );
  OAI221_X1 U10681 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput53), .C1(SI_12_), 
        .C2(keyinput8), .A(n9536), .ZN(n9543) );
  AOI22_X1 U10682 ( .A1(P2_D_REG_16__SCAN_IN), .A2(keyinput27), .B1(
        P2_D_REG_4__SCAN_IN), .B2(keyinput56), .ZN(n9537) );
  OAI221_X1 U10683 ( .B1(P2_D_REG_16__SCAN_IN), .B2(keyinput27), .C1(
        P2_D_REG_4__SCAN_IN), .C2(keyinput56), .A(n9537), .ZN(n9542) );
  AOI22_X1 U10684 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput15), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput25), .ZN(n9538) );
  OAI221_X1 U10685 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput15), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput25), .A(n9538), .ZN(n9541) );
  AOI22_X1 U10686 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(keyinput14), .B1(
        P2_IR_REG_7__SCAN_IN), .B2(keyinput4), .ZN(n9539) );
  OAI221_X1 U10687 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(keyinput14), .C1(
        P2_IR_REG_7__SCAN_IN), .C2(keyinput4), .A(n9539), .ZN(n9540) );
  NOR4_X1 U10688 ( .A1(n9543), .A2(n9542), .A3(n9541), .A4(n9540), .ZN(n9625)
         );
  AOI22_X1 U10689 ( .A1(P1_D_REG_16__SCAN_IN), .A2(keyinput23), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(keyinput48), .ZN(n9544) );
  OAI221_X1 U10690 ( .B1(P1_D_REG_16__SCAN_IN), .B2(keyinput23), .C1(
        P1_DATAO_REG_25__SCAN_IN), .C2(keyinput48), .A(n9544), .ZN(n9551) );
  AOI22_X1 U10691 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput7), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(keyinput38), .ZN(n9545) );
  OAI221_X1 U10692 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput7), .C1(
        P1_DATAO_REG_8__SCAN_IN), .C2(keyinput38), .A(n9545), .ZN(n9550) );
  AOI22_X1 U10693 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(keyinput6), .B1(
        P1_STATE_REG_SCAN_IN), .B2(keyinput2), .ZN(n9546) );
  OAI221_X1 U10694 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(keyinput6), .C1(
        P1_STATE_REG_SCAN_IN), .C2(keyinput2), .A(n9546), .ZN(n9549) );
  AOI22_X1 U10695 ( .A1(P1_REG0_REG_23__SCAN_IN), .A2(keyinput61), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(keyinput11), .ZN(n9547) );
  OAI221_X1 U10696 ( .B1(P1_REG0_REG_23__SCAN_IN), .B2(keyinput61), .C1(
        P2_DATAO_REG_8__SCAN_IN), .C2(keyinput11), .A(n9547), .ZN(n9548) );
  NOR4_X1 U10697 ( .A1(n9551), .A2(n9550), .A3(n9549), .A4(n9548), .ZN(n9624)
         );
  INV_X1 U10698 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9553) );
  AOI22_X1 U10699 ( .A1(n9553), .A2(keyinput21), .B1(keyinput36), .B2(n5750), 
        .ZN(n9552) );
  OAI221_X1 U10700 ( .B1(n9553), .B2(keyinput21), .C1(n5750), .C2(keyinput36), 
        .A(n9552), .ZN(n9563) );
  INV_X1 U10701 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n9556) );
  INV_X1 U10702 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9555) );
  AOI22_X1 U10703 ( .A1(n9556), .A2(keyinput34), .B1(n9555), .B2(keyinput44), 
        .ZN(n9554) );
  OAI221_X1 U10704 ( .B1(n9556), .B2(keyinput34), .C1(n9555), .C2(keyinput44), 
        .A(n9554), .ZN(n9562) );
  AOI22_X1 U10705 ( .A1(n6794), .A2(keyinput18), .B1(n7029), .B2(keyinput1), 
        .ZN(n9557) );
  OAI221_X1 U10706 ( .B1(n6794), .B2(keyinput18), .C1(n7029), .C2(keyinput1), 
        .A(n9557), .ZN(n9561) );
  AOI22_X1 U10707 ( .A1(n9559), .A2(keyinput30), .B1(keyinput52), .B2(n9929), 
        .ZN(n9558) );
  OAI221_X1 U10708 ( .B1(n9559), .B2(keyinput30), .C1(n9929), .C2(keyinput52), 
        .A(n9558), .ZN(n9560) );
  NOR4_X1 U10709 ( .A1(n9563), .A2(n9562), .A3(n9561), .A4(n9560), .ZN(n9622)
         );
  AOI22_X1 U10710 ( .A1(P2_D_REG_13__SCAN_IN), .A2(keyinput16), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(keyinput10), .ZN(n9564) );
  OAI221_X1 U10711 ( .B1(P2_D_REG_13__SCAN_IN), .B2(keyinput16), .C1(
        P2_DATAO_REG_18__SCAN_IN), .C2(keyinput10), .A(n9564), .ZN(n9571) );
  AOI22_X1 U10712 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(keyinput35), .B1(
        P2_REG1_REG_3__SCAN_IN), .B2(keyinput20), .ZN(n9565) );
  OAI221_X1 U10713 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(keyinput35), .C1(
        P2_REG1_REG_3__SCAN_IN), .C2(keyinput20), .A(n9565), .ZN(n9570) );
  AOI22_X1 U10714 ( .A1(P2_D_REG_22__SCAN_IN), .A2(keyinput24), .B1(
        P1_REG3_REG_8__SCAN_IN), .B2(keyinput26), .ZN(n9566) );
  OAI221_X1 U10715 ( .B1(P2_D_REG_22__SCAN_IN), .B2(keyinput24), .C1(
        P1_REG3_REG_8__SCAN_IN), .C2(keyinput26), .A(n9566), .ZN(n9569) );
  AOI22_X1 U10716 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(keyinput46), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(keyinput45), .ZN(n9567) );
  OAI221_X1 U10717 ( .B1(P1_DATAO_REG_2__SCAN_IN), .B2(keyinput46), .C1(
        P1_DATAO_REG_18__SCAN_IN), .C2(keyinput45), .A(n9567), .ZN(n9568) );
  NOR4_X1 U10718 ( .A1(n9571), .A2(n9570), .A3(n9569), .A4(n9568), .ZN(n9621)
         );
  AOI22_X1 U10719 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(keyinput49), .B1(
        P2_REG1_REG_5__SCAN_IN), .B2(keyinput39), .ZN(n9572) );
  OAI221_X1 U10720 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(keyinput49), .C1(
        P2_REG1_REG_5__SCAN_IN), .C2(keyinput39), .A(n9572), .ZN(n9579) );
  AOI22_X1 U10721 ( .A1(SI_9_), .A2(keyinput0), .B1(SI_19_), .B2(keyinput51), 
        .ZN(n9573) );
  OAI221_X1 U10722 ( .B1(SI_9_), .B2(keyinput0), .C1(SI_19_), .C2(keyinput51), 
        .A(n9573), .ZN(n9578) );
  AOI22_X1 U10723 ( .A1(P2_REG1_REG_22__SCAN_IN), .A2(keyinput17), .B1(
        P1_REG2_REG_0__SCAN_IN), .B2(keyinput5), .ZN(n9574) );
  OAI221_X1 U10724 ( .B1(P2_REG1_REG_22__SCAN_IN), .B2(keyinput17), .C1(
        P1_REG2_REG_0__SCAN_IN), .C2(keyinput5), .A(n9574), .ZN(n9577) );
  AOI22_X1 U10725 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(keyinput22), .B1(
        P1_IR_REG_25__SCAN_IN), .B2(keyinput33), .ZN(n9575) );
  OAI221_X1 U10726 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(keyinput22), .C1(
        P1_IR_REG_25__SCAN_IN), .C2(keyinput33), .A(n9575), .ZN(n9576) );
  NOR4_X1 U10727 ( .A1(n9579), .A2(n9578), .A3(n9577), .A4(n9576), .ZN(n9620)
         );
  INV_X1 U10728 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9581) );
  AOI22_X1 U10729 ( .A1(n9581), .A2(keyinput57), .B1(keyinput59), .B2(n7568), 
        .ZN(n9580) );
  OAI221_X1 U10730 ( .B1(n9581), .B2(keyinput57), .C1(n7568), .C2(keyinput59), 
        .A(n9580), .ZN(n9589) );
  INV_X1 U10731 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9584) );
  AOI22_X1 U10732 ( .A1(n9584), .A2(keyinput12), .B1(n9583), .B2(keyinput47), 
        .ZN(n9582) );
  OAI221_X1 U10733 ( .B1(n9584), .B2(keyinput12), .C1(n9583), .C2(keyinput47), 
        .A(n9582), .ZN(n9588) );
  AOI22_X1 U10734 ( .A1(n5967), .A2(keyinput42), .B1(n9586), .B2(keyinput41), 
        .ZN(n9585) );
  OAI221_X1 U10735 ( .B1(n5967), .B2(keyinput42), .C1(n9586), .C2(keyinput41), 
        .A(n9585), .ZN(n9587) );
  NOR3_X1 U10736 ( .A1(n9589), .A2(n9588), .A3(n9587), .ZN(n9618) );
  INV_X1 U10737 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9832) );
  AOI22_X1 U10738 ( .A1(n9832), .A2(keyinput40), .B1(keyinput54), .B2(n9591), 
        .ZN(n9590) );
  OAI221_X1 U10739 ( .B1(n9832), .B2(keyinput40), .C1(n9591), .C2(keyinput54), 
        .A(n9590), .ZN(n9597) );
  XNOR2_X1 U10740 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput43), .ZN(n9595) );
  XNOR2_X1 U10741 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput62), .ZN(n9594) );
  XNOR2_X1 U10742 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput37), .ZN(n9593) );
  XNOR2_X1 U10743 ( .A(P2_REG0_REG_22__SCAN_IN), .B(keyinput3), .ZN(n9592) );
  NAND4_X1 U10744 ( .A1(n9595), .A2(n9594), .A3(n9593), .A4(n9592), .ZN(n9596)
         );
  NOR2_X1 U10745 ( .A1(n9597), .A2(n9596), .ZN(n9617) );
  INV_X1 U10746 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n9599) );
  AOI22_X1 U10747 ( .A1(n9599), .A2(keyinput13), .B1(n5883), .B2(keyinput31), 
        .ZN(n9598) );
  OAI221_X1 U10748 ( .B1(n9599), .B2(keyinput13), .C1(n5883), .C2(keyinput31), 
        .A(n9598), .ZN(n9607) );
  AOI22_X1 U10749 ( .A1(n9602), .A2(keyinput63), .B1(keyinput32), .B2(n9601), 
        .ZN(n9600) );
  OAI221_X1 U10750 ( .B1(n9602), .B2(keyinput63), .C1(n9601), .C2(keyinput32), 
        .A(n9600), .ZN(n9606) );
  AOI22_X1 U10751 ( .A1(P2_REG0_REG_27__SCAN_IN), .A2(keyinput29), .B1(n9604), 
        .B2(keyinput28), .ZN(n9603) );
  OAI221_X1 U10752 ( .B1(P2_REG0_REG_27__SCAN_IN), .B2(keyinput29), .C1(n9604), 
        .C2(keyinput28), .A(n9603), .ZN(n9605) );
  NOR3_X1 U10753 ( .A1(n9607), .A2(n9606), .A3(n9605), .ZN(n9616) );
  INV_X1 U10754 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9930) );
  AOI22_X1 U10755 ( .A1(n5720), .A2(keyinput50), .B1(n9930), .B2(keyinput19), 
        .ZN(n9608) );
  OAI221_X1 U10756 ( .B1(n5720), .B2(keyinput50), .C1(n9930), .C2(keyinput19), 
        .A(n9608), .ZN(n9614) );
  XNOR2_X1 U10757 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput60), .ZN(n9612) );
  XNOR2_X1 U10758 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput9), .ZN(n9611) );
  XNOR2_X1 U10759 ( .A(keyinput58), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n9610) );
  XNOR2_X1 U10760 ( .A(keyinput55), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n9609) );
  NAND4_X1 U10761 ( .A1(n9612), .A2(n9611), .A3(n9610), .A4(n9609), .ZN(n9613)
         );
  NOR2_X1 U10762 ( .A1(n9614), .A2(n9613), .ZN(n9615) );
  AND4_X1 U10763 ( .A1(n9618), .A2(n9617), .A3(n9616), .A4(n9615), .ZN(n9619)
         );
  AND4_X1 U10764 ( .A1(n9622), .A2(n9621), .A3(n9620), .A4(n9619), .ZN(n9623)
         );
  NAND4_X1 U10765 ( .A1(n9626), .A2(n9625), .A3(n9624), .A4(n9623), .ZN(n9627)
         );
  XNOR2_X1 U10766 ( .A(n9628), .B(n9627), .ZN(P1_U3521) );
  MUX2_X1 U10767 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9629), .S(n9897), .Z(
        P1_U3520) );
  MUX2_X1 U10768 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9630), .S(n9897), .Z(
        P1_U3519) );
  MUX2_X1 U10769 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9631), .S(n9897), .Z(
        P1_U3518) );
  MUX2_X1 U10770 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9632), .S(n9897), .Z(
        P1_U3517) );
  MUX2_X1 U10771 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9633), .S(n9897), .Z(
        P1_U3516) );
  MUX2_X1 U10772 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9634), .S(n9897), .Z(
        P1_U3515) );
  MUX2_X1 U10773 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9635), .S(n9897), .Z(
        P1_U3514) );
  MUX2_X1 U10774 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9636), .S(n9897), .Z(
        P1_U3513) );
  MUX2_X1 U10775 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9637), .S(n9897), .Z(
        P1_U3512) );
  MUX2_X1 U10776 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9638), .S(n9897), .Z(
        P1_U3511) );
  MUX2_X1 U10777 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9639), .S(n9897), .Z(
        P1_U3510) );
  MUX2_X1 U10778 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9640), .S(n9897), .Z(
        P1_U3508) );
  MUX2_X1 U10779 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9641), .S(n9897), .Z(
        P1_U3505) );
  MUX2_X1 U10780 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9642), .S(n9897), .Z(
        P1_U3502) );
  MUX2_X1 U10781 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9643), .S(n9897), .Z(
        P1_U3499) );
  MUX2_X1 U10782 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9644), .S(n9897), .Z(
        P1_U3496) );
  NOR4_X1 U10783 ( .A1(n9645), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n5122), .ZN(n9646) );
  AOI21_X1 U10784 ( .B1(n9647), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9646), .ZN(
        n9648) );
  OAI21_X1 U10785 ( .B1(n9649), .B2(n9653), .A(n9648), .ZN(P1_U3322) );
  AOI22_X1 U10786 ( .A1(n9651), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9650), .ZN(n9652) );
  OAI21_X1 U10787 ( .B1(n9654), .B2(n9653), .A(n9652), .ZN(P1_U3323) );
  MUX2_X1 U10788 ( .A(n9656), .B(n9655), .S(P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10789 ( .A1(n9920), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9668) );
  OAI211_X1 U10790 ( .C1(n9659), .C2(n9658), .A(n9914), .B(n9657), .ZN(n9660)
         );
  OAI21_X1 U10791 ( .B1(n9915), .B2(n9661), .A(n9660), .ZN(n9662) );
  INV_X1 U10792 ( .A(n9662), .ZN(n9667) );
  OAI211_X1 U10793 ( .C1(n9665), .C2(n9664), .A(n9912), .B(n9663), .ZN(n9666)
         );
  NAND3_X1 U10794 ( .A1(n9668), .A2(n9667), .A3(n9666), .ZN(P2_U3247) );
  INV_X1 U10795 ( .A(n9674), .ZN(n9676) );
  AOI211_X1 U10796 ( .C1(n9887), .C2(n9671), .A(n9670), .B(n9669), .ZN(n9672)
         );
  OAI21_X1 U10797 ( .B1(n9674), .B2(n9673), .A(n9672), .ZN(n9675) );
  AOI21_X1 U10798 ( .B1(n9719), .B2(n9676), .A(n9675), .ZN(n9679) );
  INV_X1 U10799 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9677) );
  AOI22_X1 U10800 ( .A1(n9897), .A2(n9679), .B1(n9677), .B2(n9895), .ZN(
        P1_U3484) );
  AOI22_X1 U10801 ( .A1(n9911), .A2(n9679), .B1(n9678), .B2(n9909), .ZN(
        P1_U3533) );
  XNOR2_X1 U10802 ( .A(n9681), .B(n9680), .ZN(n9732) );
  AND2_X1 U10803 ( .A1(n4828), .A2(n9697), .ZN(n9683) );
  OR2_X1 U10804 ( .A1(n9683), .A2(n9682), .ZN(n9730) );
  INV_X1 U10805 ( .A(n9730), .ZN(n9684) );
  AOI22_X1 U10806 ( .A1(n9732), .A2(n9707), .B1(n9706), .B2(n9684), .ZN(n9700)
         );
  INV_X1 U10807 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9687) );
  OAI22_X1 U10808 ( .A1(n9725), .A2(n9687), .B1(n9686), .B2(n9685), .ZN(n9696)
         );
  XNOR2_X1 U10809 ( .A(n9689), .B(n9688), .ZN(n9693) );
  OAI22_X1 U10810 ( .A1(n9711), .A2(n9712), .B1(n9690), .B2(n9710), .ZN(n9691)
         );
  INV_X1 U10811 ( .A(n9691), .ZN(n9692) );
  OAI21_X1 U10812 ( .B1(n9693), .B2(n9716), .A(n9692), .ZN(n9694) );
  AOI21_X1 U10813 ( .B1(n9732), .B2(n9719), .A(n9694), .ZN(n9734) );
  NOR2_X1 U10814 ( .A1(n9734), .A2(n9309), .ZN(n9695) );
  AOI211_X1 U10815 ( .C1(n9698), .C2(n9697), .A(n9696), .B(n9695), .ZN(n9699)
         );
  NAND2_X1 U10816 ( .A1(n9700), .A2(n9699), .ZN(P1_U3278) );
  XNOR2_X1 U10817 ( .A(n9701), .B(n9708), .ZN(n9738) );
  OR2_X1 U10818 ( .A1(n9702), .A2(n9735), .ZN(n9703) );
  NAND2_X1 U10819 ( .A1(n9704), .A2(n9703), .ZN(n9736) );
  INV_X1 U10820 ( .A(n9736), .ZN(n9705) );
  AOI22_X1 U10821 ( .A1(n9738), .A2(n9707), .B1(n9706), .B2(n9705), .ZN(n9728)
         );
  XNOR2_X1 U10822 ( .A(n9709), .B(n9708), .ZN(n9717) );
  OAI22_X1 U10823 ( .A1(n9713), .A2(n9712), .B1(n9711), .B2(n9710), .ZN(n9714)
         );
  INV_X1 U10824 ( .A(n9714), .ZN(n9715) );
  OAI21_X1 U10825 ( .B1(n9717), .B2(n9716), .A(n9715), .ZN(n9718) );
  AOI21_X1 U10826 ( .B1(n9738), .B2(n9719), .A(n9718), .ZN(n9740) );
  INV_X1 U10827 ( .A(n9740), .ZN(n9726) );
  AOI22_X1 U10828 ( .A1(n9309), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9721), .B2(
        n9720), .ZN(n9722) );
  OAI21_X1 U10829 ( .B1(n9735), .B2(n9723), .A(n9722), .ZN(n9724) );
  AOI21_X1 U10830 ( .B1(n9726), .B2(n9725), .A(n9724), .ZN(n9727) );
  NAND2_X1 U10831 ( .A1(n9728), .A2(n9727), .ZN(P1_U3280) );
  OAI22_X1 U10832 ( .A1(n9730), .A2(n9854), .B1(n9729), .B2(n9852), .ZN(n9731)
         );
  AOI21_X1 U10833 ( .B1(n9732), .B2(n9884), .A(n9731), .ZN(n9733) );
  AND2_X1 U10834 ( .A1(n9734), .A2(n9733), .ZN(n9743) );
  AOI22_X1 U10835 ( .A1(n9911), .A2(n9743), .B1(n7158), .B2(n9909), .ZN(
        P1_U3536) );
  OAI22_X1 U10836 ( .A1(n9736), .A2(n9854), .B1(n9735), .B2(n9852), .ZN(n9737)
         );
  AOI21_X1 U10837 ( .B1(n9738), .B2(n9884), .A(n9737), .ZN(n9739) );
  AND2_X1 U10838 ( .A1(n9740), .A2(n9739), .ZN(n9745) );
  AOI22_X1 U10839 ( .A1(n9911), .A2(n9745), .B1(n9741), .B2(n9909), .ZN(
        P1_U3534) );
  INV_X1 U10840 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9742) );
  AOI22_X1 U10841 ( .A1(n9897), .A2(n9743), .B1(n9742), .B2(n9895), .ZN(
        P1_U3493) );
  INV_X1 U10842 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9744) );
  AOI22_X1 U10843 ( .A1(n9897), .A2(n9745), .B1(n9744), .B2(n9895), .ZN(
        P1_U3487) );
  XNOR2_X1 U10844 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10845 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10846 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9764) );
  MUX2_X1 U10847 ( .A(n9747), .B(n9746), .S(n6565), .Z(n9749) );
  OAI211_X1 U10848 ( .C1(n9749), .C2(n5639), .A(P1_U4006), .B(n9748), .ZN(
        n9780) );
  NAND2_X1 U10849 ( .A1(n9827), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n9758) );
  NAND2_X1 U10850 ( .A1(n9825), .A2(n9750), .ZN(n9757) );
  MUX2_X1 U10851 ( .A(n6575), .B(P1_REG2_REG_2__SCAN_IN), .S(n9750), .Z(n9753)
         );
  INV_X1 U10852 ( .A(n9751), .ZN(n9752) );
  NAND2_X1 U10853 ( .A1(n9753), .A2(n9752), .ZN(n9754) );
  NAND3_X1 U10854 ( .A1(n9798), .A2(n9755), .A3(n9754), .ZN(n9756) );
  AND4_X1 U10855 ( .A1(n9780), .A2(n9758), .A3(n9757), .A4(n9756), .ZN(n9763)
         );
  OAI211_X1 U10856 ( .C1(n9761), .C2(n9760), .A(n9823), .B(n9759), .ZN(n9762)
         );
  OAI211_X1 U10857 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9764), .A(n9763), .B(
        n9762), .ZN(P1_U3243) );
  INV_X1 U10858 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9772) );
  OAI21_X1 U10859 ( .B1(n9767), .B2(n9766), .A(n9765), .ZN(n9768) );
  NAND2_X1 U10860 ( .A1(n9798), .A2(n9768), .ZN(n9771) );
  NAND2_X1 U10861 ( .A1(n9825), .A2(n9769), .ZN(n9770) );
  OAI211_X1 U10862 ( .C1(n9773), .C2(n9772), .A(n9771), .B(n9770), .ZN(n9774)
         );
  INV_X1 U10863 ( .A(n9774), .ZN(n9782) );
  OAI21_X1 U10864 ( .B1(n9777), .B2(n9776), .A(n9775), .ZN(n9778) );
  NAND2_X1 U10865 ( .A1(n9823), .A2(n9778), .ZN(n9779) );
  NAND4_X1 U10866 ( .A1(n9782), .A2(n9781), .A3(n9780), .A4(n9779), .ZN(
        P1_U3245) );
  AOI22_X1 U10867 ( .A1(n9827), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n9783), .B2(
        n9825), .ZN(n9795) );
  NOR2_X1 U10868 ( .A1(n9785), .A2(n9784), .ZN(n9786) );
  OAI21_X1 U10869 ( .B1(n9787), .B2(n9786), .A(n9798), .ZN(n9793) );
  NAND2_X1 U10870 ( .A1(n9789), .A2(n9788), .ZN(n9790) );
  NAND3_X1 U10871 ( .A1(n9823), .A2(n9791), .A3(n9790), .ZN(n9792) );
  NAND4_X1 U10872 ( .A1(n9795), .A2(n9794), .A3(n9793), .A4(n9792), .ZN(
        P1_U3246) );
  AND4_X1 U10873 ( .A1(n9805), .A2(P1_REG1_REG_8__SCAN_IN), .A3(n9807), .A4(
        n9823), .ZN(n9796) );
  AOI211_X1 U10874 ( .C1(n9827), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9797), .B(
        n9796), .ZN(n9812) );
  INV_X1 U10875 ( .A(n9807), .ZN(n9802) );
  NAND2_X1 U10876 ( .A1(n9802), .A2(n4481), .ZN(n9800) );
  OAI211_X1 U10877 ( .C1(n9801), .C2(n9800), .A(n9799), .B(n9798), .ZN(n9811)
         );
  NAND2_X1 U10878 ( .A1(n9802), .A2(n9907), .ZN(n9804) );
  OAI211_X1 U10879 ( .C1(n9805), .C2(n9804), .A(n9803), .B(n9823), .ZN(n9810)
         );
  OAI211_X1 U10880 ( .C1(n9808), .C2(n5639), .A(n9807), .B(n9806), .ZN(n9809)
         );
  NAND4_X1 U10881 ( .A1(n9812), .A2(n9811), .A3(n9810), .A4(n9809), .ZN(
        P1_U3249) );
  OAI21_X1 U10882 ( .B1(n9815), .B2(n9814), .A(n9813), .ZN(n9824) );
  INV_X1 U10883 ( .A(n9816), .ZN(n9822) );
  AOI211_X1 U10884 ( .C1(n9820), .C2(n9819), .A(n9818), .B(n9817), .ZN(n9821)
         );
  AOI211_X1 U10885 ( .C1(n9824), .C2(n9823), .A(n9822), .B(n9821), .ZN(n9829)
         );
  AOI22_X1 U10886 ( .A1(n9827), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(n9826), .B2(
        n9825), .ZN(n9828) );
  NAND2_X1 U10887 ( .A1(n9829), .A2(n9828), .ZN(P1_U3251) );
  INV_X1 U10888 ( .A(n9830), .ZN(n9831) );
  AND2_X1 U10889 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9835), .ZN(P1_U3292) );
  AND2_X1 U10890 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9835), .ZN(P1_U3293) );
  AND2_X1 U10891 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9835), .ZN(P1_U3294) );
  AND2_X1 U10892 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9835), .ZN(P1_U3295) );
  AND2_X1 U10893 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9835), .ZN(P1_U3296) );
  AND2_X1 U10894 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9835), .ZN(P1_U3297) );
  AND2_X1 U10895 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9835), .ZN(P1_U3298) );
  AND2_X1 U10896 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9835), .ZN(P1_U3299) );
  AND2_X1 U10897 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9835), .ZN(P1_U3300) );
  AND2_X1 U10898 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9835), .ZN(P1_U3301) );
  INV_X1 U10899 ( .A(n9835), .ZN(n9834) );
  NOR2_X1 U10900 ( .A1(n9834), .A2(n9832), .ZN(P1_U3302) );
  AND2_X1 U10901 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9835), .ZN(P1_U3303) );
  AND2_X1 U10902 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9835), .ZN(P1_U3304) );
  AND2_X1 U10903 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9835), .ZN(P1_U3305) );
  AND2_X1 U10904 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9835), .ZN(P1_U3306) );
  NOR2_X1 U10905 ( .A1(n9834), .A2(n9833), .ZN(P1_U3307) );
  AND2_X1 U10906 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9835), .ZN(P1_U3308) );
  AND2_X1 U10907 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9835), .ZN(P1_U3309) );
  AND2_X1 U10908 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9835), .ZN(P1_U3310) );
  AND2_X1 U10909 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9835), .ZN(P1_U3311) );
  AND2_X1 U10910 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9835), .ZN(P1_U3312) );
  AND2_X1 U10911 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9835), .ZN(P1_U3313) );
  AND2_X1 U10912 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9835), .ZN(P1_U3314) );
  AND2_X1 U10913 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9835), .ZN(P1_U3315) );
  AND2_X1 U10914 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9835), .ZN(P1_U3316) );
  AND2_X1 U10915 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9835), .ZN(P1_U3317) );
  AND2_X1 U10916 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9835), .ZN(P1_U3318) );
  AND2_X1 U10917 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9835), .ZN(P1_U3319) );
  AND2_X1 U10918 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9835), .ZN(P1_U3320) );
  AND2_X1 U10919 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9835), .ZN(P1_U3321) );
  AOI21_X1 U10920 ( .B1(P1_D_REG_1__SCAN_IN), .B2(n9837), .A(n9836), .ZN(n9838) );
  INV_X1 U10921 ( .A(n9838), .ZN(P1_U3441) );
  OAI21_X1 U10922 ( .B1(n9840), .B2(n9854), .A(n9839), .ZN(n9842) );
  AOI211_X1 U10923 ( .C1(n9873), .C2(n9843), .A(n9842), .B(n9841), .ZN(n9898)
         );
  INV_X1 U10924 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9844) );
  AOI22_X1 U10925 ( .A1(n9897), .A2(n9898), .B1(n9844), .B2(n9895), .ZN(
        P1_U3463) );
  NAND2_X1 U10926 ( .A1(n9845), .A2(n9888), .ZN(n9846) );
  OAI21_X1 U10927 ( .B1(n9847), .B2(n9852), .A(n9846), .ZN(n9849) );
  AOI211_X1 U10928 ( .C1(n9884), .C2(n9850), .A(n9849), .B(n9848), .ZN(n9900)
         );
  INV_X1 U10929 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9851) );
  AOI22_X1 U10930 ( .A1(n9897), .A2(n9900), .B1(n9851), .B2(n9895), .ZN(
        P1_U3466) );
  OAI22_X1 U10931 ( .A1(n9855), .A2(n9854), .B1(n9853), .B2(n9852), .ZN(n9858)
         );
  INV_X1 U10932 ( .A(n9856), .ZN(n9857) );
  AOI211_X1 U10933 ( .C1(n9859), .C2(n9873), .A(n9858), .B(n9857), .ZN(n9902)
         );
  INV_X1 U10934 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9860) );
  AOI22_X1 U10935 ( .A1(n9897), .A2(n9902), .B1(n9860), .B2(n9895), .ZN(
        P1_U3469) );
  AOI21_X1 U10936 ( .B1(n9862), .B2(n9888), .A(n9861), .ZN(n9863) );
  OAI211_X1 U10937 ( .C1(n9865), .C2(n9881), .A(n9864), .B(n9863), .ZN(n9866)
         );
  AOI21_X1 U10938 ( .B1(n9884), .B2(n9867), .A(n9866), .ZN(n9904) );
  INV_X1 U10939 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9868) );
  AOI22_X1 U10940 ( .A1(n9897), .A2(n9904), .B1(n9868), .B2(n9895), .ZN(
        P1_U3472) );
  NAND3_X1 U10941 ( .A1(n9871), .A2(n9870), .A3(n9869), .ZN(n9872) );
  AOI21_X1 U10942 ( .B1(n9874), .B2(n9873), .A(n9872), .ZN(n9906) );
  INV_X1 U10943 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9875) );
  AOI22_X1 U10944 ( .A1(n9897), .A2(n9906), .B1(n9875), .B2(n9895), .ZN(
        P1_U3475) );
  INV_X1 U10945 ( .A(n9880), .ZN(n9883) );
  AOI211_X1 U10946 ( .C1(n9888), .C2(n9878), .A(n9877), .B(n9876), .ZN(n9879)
         );
  OAI21_X1 U10947 ( .B1(n9881), .B2(n9880), .A(n9879), .ZN(n9882) );
  AOI21_X1 U10948 ( .B1(n9884), .B2(n9883), .A(n9882), .ZN(n9908) );
  INV_X1 U10949 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9885) );
  AOI22_X1 U10950 ( .A1(n9897), .A2(n9908), .B1(n9885), .B2(n9895), .ZN(
        P1_U3478) );
  AOI22_X1 U10951 ( .A1(n9889), .A2(n9888), .B1(n9887), .B2(n9886), .ZN(n9890)
         );
  OAI211_X1 U10952 ( .C1(n9893), .C2(n9892), .A(n9891), .B(n9890), .ZN(n9894)
         );
  INV_X1 U10953 ( .A(n9894), .ZN(n9910) );
  INV_X1 U10954 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9896) );
  AOI22_X1 U10955 ( .A1(n9897), .A2(n9910), .B1(n9896), .B2(n9895), .ZN(
        P1_U3481) );
  AOI22_X1 U10956 ( .A1(n9911), .A2(n9898), .B1(n6595), .B2(n9909), .ZN(
        P1_U3526) );
  AOI22_X1 U10957 ( .A1(n9911), .A2(n9900), .B1(n9899), .B2(n9909), .ZN(
        P1_U3527) );
  AOI22_X1 U10958 ( .A1(n9911), .A2(n9902), .B1(n9901), .B2(n9909), .ZN(
        P1_U3528) );
  AOI22_X1 U10959 ( .A1(n9911), .A2(n9904), .B1(n9903), .B2(n9909), .ZN(
        P1_U3529) );
  AOI22_X1 U10960 ( .A1(n9911), .A2(n9906), .B1(n9905), .B2(n9909), .ZN(
        P1_U3530) );
  AOI22_X1 U10961 ( .A1(n9911), .A2(n9908), .B1(n9907), .B2(n9909), .ZN(
        P1_U3531) );
  AOI22_X1 U10962 ( .A1(n9911), .A2(n9910), .B1(n6605), .B2(n9909), .ZN(
        P1_U3532) );
  AOI22_X1 U10963 ( .A1(n9912), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9914), .ZN(n9924) );
  INV_X1 U10964 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9913) );
  NAND2_X1 U10965 ( .A1(n9914), .A2(n9913), .ZN(n9916) );
  OAI211_X1 U10966 ( .C1(n9917), .C2(P2_REG2_REG_0__SCAN_IN), .A(n9916), .B(
        n9915), .ZN(n9918) );
  INV_X1 U10967 ( .A(n9918), .ZN(n9922) );
  AOI22_X1 U10968 ( .A1(n9920), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9921) );
  OAI221_X1 U10969 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9924), .C1(n9923), .C2(
        n9922), .A(n9921), .ZN(P2_U3245) );
  NOR2_X1 U10970 ( .A1(n9926), .A2(n9925), .ZN(n9931) );
  AND2_X1 U10971 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9934), .ZN(P2_U3297) );
  AND2_X1 U10972 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9934), .ZN(P2_U3298) );
  AND2_X1 U10973 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9934), .ZN(P2_U3299) );
  AND2_X1 U10974 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9934), .ZN(P2_U3300) );
  AND2_X1 U10975 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9934), .ZN(P2_U3301) );
  AND2_X1 U10976 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9934), .ZN(P2_U3302) );
  AND2_X1 U10977 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9934), .ZN(P2_U3303) );
  AND2_X1 U10978 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9934), .ZN(P2_U3304) );
  AND2_X1 U10979 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9934), .ZN(P2_U3305) );
  NOR2_X1 U10980 ( .A1(n9931), .A2(n9927), .ZN(P2_U3306) );
  AND2_X1 U10981 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9934), .ZN(P2_U3307) );
  AND2_X1 U10982 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9934), .ZN(P2_U3308) );
  AND2_X1 U10983 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9934), .ZN(P2_U3309) );
  AND2_X1 U10984 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9934), .ZN(P2_U3310) );
  AND2_X1 U10985 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9934), .ZN(P2_U3311) );
  NOR2_X1 U10986 ( .A1(n9931), .A2(n9928), .ZN(P2_U3312) );
  AND2_X1 U10987 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9934), .ZN(P2_U3313) );
  AND2_X1 U10988 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9934), .ZN(P2_U3314) );
  AND2_X1 U10989 ( .A1(n9934), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3315) );
  AND2_X1 U10990 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9934), .ZN(P2_U3316) );
  NOR2_X1 U10991 ( .A1(n9931), .A2(n9929), .ZN(P2_U3317) );
  AND2_X1 U10992 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9934), .ZN(P2_U3318) );
  AND2_X1 U10993 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9934), .ZN(P2_U3319) );
  AND2_X1 U10994 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9934), .ZN(P2_U3320) );
  AND2_X1 U10995 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9934), .ZN(P2_U3321) );
  AND2_X1 U10996 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9934), .ZN(P2_U3322) );
  AND2_X1 U10997 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9934), .ZN(P2_U3323) );
  AND2_X1 U10998 ( .A1(n9934), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3324) );
  AND2_X1 U10999 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9934), .ZN(P2_U3325) );
  NOR2_X1 U11000 ( .A1(n9931), .A2(n9930), .ZN(P2_U3326) );
  AOI22_X1 U11001 ( .A1(n9937), .A2(n9933), .B1(n9932), .B2(n9934), .ZN(
        P2_U3437) );
  AOI22_X1 U11002 ( .A1(n9937), .A2(n9936), .B1(n9935), .B2(n9934), .ZN(
        P2_U3438) );
  AOI22_X1 U11003 ( .A1(n9940), .A2(n9985), .B1(n9939), .B2(n9938), .ZN(n9941)
         );
  AND2_X1 U11004 ( .A1(n9942), .A2(n9941), .ZN(n9989) );
  INV_X1 U11005 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9943) );
  AOI22_X1 U11006 ( .A1(n9988), .A2(n9989), .B1(n9943), .B2(n9987), .ZN(
        P2_U3451) );
  OAI21_X1 U11007 ( .B1(n9945), .B2(n9980), .A(n9944), .ZN(n9948) );
  INV_X1 U11008 ( .A(n9946), .ZN(n9947) );
  AOI211_X1 U11009 ( .C1(n9985), .C2(n9949), .A(n9948), .B(n9947), .ZN(n9991)
         );
  INV_X1 U11010 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9950) );
  AOI22_X1 U11011 ( .A1(n9988), .A2(n9991), .B1(n9950), .B2(n9987), .ZN(
        P2_U3454) );
  INV_X1 U11012 ( .A(n9951), .ZN(n9953) );
  OAI22_X1 U11013 ( .A1(n9953), .A2(n9981), .B1(n9952), .B2(n9980), .ZN(n9956)
         );
  INV_X1 U11014 ( .A(n9954), .ZN(n9955) );
  AOI211_X1 U11015 ( .C1(n9985), .C2(n9957), .A(n9956), .B(n9955), .ZN(n9993)
         );
  AOI22_X1 U11016 ( .A1(n9988), .A2(n9993), .B1(n5720), .B2(n9987), .ZN(
        P2_U3463) );
  OAI211_X1 U11017 ( .C1(n9960), .C2(n9980), .A(n9959), .B(n9958), .ZN(n9961)
         );
  AOI21_X1 U11018 ( .B1(n9985), .B2(n9962), .A(n9961), .ZN(n9995) );
  AOI22_X1 U11019 ( .A1(n9988), .A2(n9995), .B1(n5735), .B2(n9987), .ZN(
        P2_U3466) );
  OAI211_X1 U11020 ( .C1(n9965), .C2(n9980), .A(n9964), .B(n9963), .ZN(n9966)
         );
  AOI21_X1 U11021 ( .B1(n9985), .B2(n9967), .A(n9966), .ZN(n9996) );
  AOI22_X1 U11022 ( .A1(n9988), .A2(n9996), .B1(n5755), .B2(n9987), .ZN(
        P2_U3469) );
  INV_X1 U11023 ( .A(n9968), .ZN(n9973) );
  OAI22_X1 U11024 ( .A1(n9970), .A2(n9981), .B1(n9969), .B2(n9980), .ZN(n9972)
         );
  AOI211_X1 U11025 ( .C1(n9979), .C2(n9973), .A(n9972), .B(n9971), .ZN(n9997)
         );
  AOI22_X1 U11026 ( .A1(n9988), .A2(n9997), .B1(n5782), .B2(n9987), .ZN(
        P2_U3475) );
  OAI22_X1 U11027 ( .A1(n9975), .A2(n9981), .B1(n9974), .B2(n9980), .ZN(n9977)
         );
  AOI211_X1 U11028 ( .C1(n9979), .C2(n9978), .A(n9977), .B(n9976), .ZN(n9998)
         );
  AOI22_X1 U11029 ( .A1(n9988), .A2(n9998), .B1(n5810), .B2(n9987), .ZN(
        P2_U3481) );
  OAI22_X1 U11030 ( .A1(n9982), .A2(n9981), .B1(n4495), .B2(n9980), .ZN(n9984)
         );
  AOI211_X1 U11031 ( .C1(n9986), .C2(n9985), .A(n9984), .B(n9983), .ZN(n10000)
         );
  AOI22_X1 U11032 ( .A1(n9988), .A2(n10000), .B1(n5841), .B2(n9987), .ZN(
        P2_U3487) );
  AOI22_X1 U11033 ( .A1(n10001), .A2(n9989), .B1(n9913), .B2(n9999), .ZN(
        P2_U3520) );
  AOI22_X1 U11034 ( .A1(n10001), .A2(n9991), .B1(n9990), .B2(n9999), .ZN(
        P2_U3521) );
  INV_X1 U11035 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9992) );
  AOI22_X1 U11036 ( .A1(n10001), .A2(n9993), .B1(n9992), .B2(n9999), .ZN(
        P2_U3524) );
  INV_X1 U11037 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9994) );
  AOI22_X1 U11038 ( .A1(n10001), .A2(n9995), .B1(n9994), .B2(n9999), .ZN(
        P2_U3525) );
  AOI22_X1 U11039 ( .A1(n10001), .A2(n9996), .B1(n6794), .B2(n9999), .ZN(
        P2_U3526) );
  AOI22_X1 U11040 ( .A1(n10001), .A2(n9997), .B1(n6841), .B2(n9999), .ZN(
        P2_U3528) );
  AOI22_X1 U11041 ( .A1(n10001), .A2(n9998), .B1(n7174), .B2(n9999), .ZN(
        P2_U3530) );
  AOI22_X1 U11042 ( .A1(n10001), .A2(n10000), .B1(n7563), .B2(n9999), .ZN(
        P2_U3532) );
  INV_X1 U11043 ( .A(n10002), .ZN(n10003) );
  NAND2_X1 U11044 ( .A1(n10004), .A2(n10003), .ZN(n10005) );
  XOR2_X1 U11045 ( .A(n10006), .B(n10005), .Z(ADD_1071_U5) );
  XOR2_X1 U11046 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11047 ( .B1(n10009), .B2(n10008), .A(n10007), .ZN(ADD_1071_U56) );
  OAI21_X1 U11048 ( .B1(n10012), .B2(n10011), .A(n10010), .ZN(ADD_1071_U57) );
  OAI21_X1 U11049 ( .B1(n10015), .B2(n10014), .A(n10013), .ZN(ADD_1071_U58) );
  OAI21_X1 U11050 ( .B1(n10018), .B2(n10017), .A(n10016), .ZN(ADD_1071_U59) );
  OAI21_X1 U11051 ( .B1(n10021), .B2(n10020), .A(n10019), .ZN(ADD_1071_U60) );
  OAI21_X1 U11052 ( .B1(n10024), .B2(n10023), .A(n10022), .ZN(ADD_1071_U61) );
  AOI21_X1 U11053 ( .B1(n10027), .B2(n10026), .A(n10025), .ZN(ADD_1071_U62) );
  AOI21_X1 U11054 ( .B1(n10030), .B2(n10029), .A(n10028), .ZN(ADD_1071_U63) );
  XOR2_X1 U11055 ( .A(n10031), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11056 ( .A1(n10033), .A2(n10032), .ZN(n10034) );
  XOR2_X1 U11057 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10034), .Z(ADD_1071_U51) );
  OAI21_X1 U11058 ( .B1(n10037), .B2(n10036), .A(n10035), .ZN(n10038) );
  XNOR2_X1 U11059 ( .A(n10038), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11060 ( .B1(n10041), .B2(n10040), .A(n10039), .ZN(ADD_1071_U47) );
  XOR2_X1 U11061 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10042), .Z(ADD_1071_U48) );
  XOR2_X1 U11062 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10043), .Z(ADD_1071_U49) );
  XOR2_X1 U11063 ( .A(n10045), .B(n10044), .Z(ADD_1071_U54) );
  XOR2_X1 U11064 ( .A(n10047), .B(n10046), .Z(ADD_1071_U53) );
  XNOR2_X1 U11065 ( .A(n10049), .B(n10048), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4826 ( .A(n5880), .Z(n6096) );
  CLKBUF_X1 U4981 ( .A(n5673), .Z(n5691) );
  NAND2_X1 U5321 ( .A1(n6769), .A2(n6617), .ZN(n5773) );
  CLKBUF_X1 U7085 ( .A(n5209), .Z(n6343) );
endmodule

