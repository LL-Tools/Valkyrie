

module b17_C_gen_AntiSAT_k_128_4 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, 
        keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, 
        keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, 
        keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, 
        keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, 
        keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, 
        keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, 
        keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, 
        keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, 
        keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, 
        keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, 
        keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, 
        keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, 
        keyinput_g61, keyinput_g62, keyinput_g63, U355, U356, U357, U358, U359, 
        U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, 
        U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, 
        U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, 
        U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, 
        U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, 
        U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, 
        U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, 
        U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9669, n9671, n9672, n9673, n9674, n9675, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
         n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
         n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
         n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982,
         n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
         n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
         n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
         n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
         n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
         n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
         n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
         n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
         n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
         n21119, n21120, n21121, n21122, n21123;

  NAND3_X1 U11100 ( .A1(n15514), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15498) );
  AOI211_X1 U11101 ( .C1(n19792), .C2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19789), .ZN(n19790) );
  INV_X1 U11102 ( .A(n20307), .ZN(n20292) );
  AOI211_X1 U11103 ( .C1(n10739), .C2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n12899), .B(n12898), .ZN(n12900) );
  AND2_X1 U11104 ( .A1(n13056), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17812) );
  NOR2_X1 U11105 ( .A1(n18964), .A2(n18972), .ZN(n18359) );
  CLKBUF_X1 U11106 ( .A(n12706), .Z(n15344) );
  CLKBUF_X2 U11107 ( .A(n13243), .Z(n19299) );
  CLKBUF_X2 U11108 ( .A(n9673), .Z(n16135) );
  INV_X1 U11109 ( .A(n17968), .ZN(n18057) );
  CLKBUF_X3 U11110 ( .A(n11791), .Z(n9684) );
  NAND2_X1 U11111 ( .A1(n12354), .A2(n12353), .ZN(n12357) );
  NAND2_X1 U11112 ( .A1(n12350), .A2(n12349), .ZN(n12352) );
  OR2_X1 U11113 ( .A1(n11989), .A2(n9722), .ZN(n19857) );
  AOI211_X2 U11114 ( .C1(n17490), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n13097), .B(n13096), .ZN(n18493) );
  XNOR2_X1 U11115 ( .A(n13489), .B(n12347), .ZN(n13570) );
  NAND2_X1 U11116 ( .A1(n10138), .A2(n11987), .ZN(n12039) );
  NAND2_X1 U11117 ( .A1(n13490), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13489) );
  OAI21_X1 U11118 ( .B1(n14237), .B2(n12400), .A(n12338), .ZN(n13490) );
  NAND2_X1 U11119 ( .A1(n11086), .A2(n11085), .ZN(n11169) );
  INV_X2 U11120 ( .A(n12951), .ZN(n9685) );
  CLKBUF_X1 U11121 ( .A(n10504), .Z(n12677) );
  INV_X2 U11122 ( .A(n9756), .ZN(n15895) );
  CLKBUF_X1 U11123 ( .A(n11145), .Z(n11099) );
  CLKBUF_X2 U11124 ( .A(n12956), .Z(n17465) );
  INV_X1 U11125 ( .A(n12956), .ZN(n17485) );
  INV_X2 U11126 ( .A(n15864), .ZN(n17490) );
  CLKBUF_X1 U11127 ( .A(n10643), .Z(n9719) );
  NAND2_X1 U11128 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18974) );
  NAND3_X1 U11129 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15945) );
  CLKBUF_X2 U11130 ( .A(n11072), .Z(n11060) );
  NAND2_X1 U11131 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19130), .ZN(
        n12921) );
  CLKBUF_X2 U11132 ( .A(n10933), .Z(n11699) );
  INV_X2 U11133 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19146) );
  INV_X2 U11134 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19130) );
  INV_X4 U11135 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19139) );
  INV_X2 U11136 ( .A(n13992), .ZN(n13596) );
  CLKBUF_X2 U11137 ( .A(n10655), .Z(n13415) );
  INV_X2 U11139 ( .A(n10885), .ZN(n12446) );
  CLKBUF_X1 U11140 ( .A(n10656), .Z(n12549) );
  INV_X2 U11141 ( .A(n12504), .ZN(n9853) );
  AND2_X1 U11142 ( .A1(n11035), .A2(n9710), .ZN(n13378) );
  NAND2_X1 U11144 ( .A1(n10657), .A2(n10655), .ZN(n10631) );
  BUF_X1 U11146 ( .A(n10943), .Z(n9679) );
  INV_X1 U11147 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9656) );
  AND2_X2 U11148 ( .A1(n10907), .A2(n14061), .ZN(n11144) );
  AND2_X2 U11149 ( .A1(n14061), .A2(n13508), .ZN(n11656) );
  AND2_X1 U11150 ( .A1(n14065), .A2(n10908), .ZN(n11093) );
  AND2_X2 U11151 ( .A1(n14065), .A2(n10907), .ZN(n11143) );
  AND2_X2 U11152 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13508) );
  AND2_X2 U11153 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15788) );
  NAND2_X1 U11154 ( .A1(n10630), .A2(n9656), .ZN(n9657) );
  NAND2_X1 U11155 ( .A1(n10629), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9658) );
  NAND2_X1 U11156 ( .A1(n12309), .A2(n12093), .ZN(n12306) );
  INV_X1 U11157 ( .A(n16609), .ZN(n9659) );
  NAND2_X1 U11158 ( .A1(n10635), .A2(n12468), .ZN(n10646) );
  NAND2_X2 U11159 ( .A1(n9858), .A2(n9859), .ZN(n12502) );
  OAI22_X1 U11161 ( .A1(n12010), .A2(n12071), .B1(n12009), .B2(n12008), .ZN(
        n12011) );
  NAND2_X1 U11162 ( .A1(n18967), .A2(n18976), .ZN(n9660) );
  INV_X1 U11163 ( .A(n18966), .ZN(n9661) );
  AND2_X1 U11164 ( .A1(n9660), .A2(n9661), .ZN(n18988) );
  OR2_X1 U11165 ( .A1(n16687), .A2(n18151), .ZN(n9662) );
  AOI21_X1 U11166 ( .B1(n13168), .B2(n13159), .A(n13251), .ZN(n18976) );
  OR2_X1 U11167 ( .A1(n16815), .A2(n18498), .ZN(n18151) );
  NAND2_X1 U11168 ( .A1(n14846), .A2(n14870), .ZN(n9663) );
  NAND2_X1 U11169 ( .A1(n14846), .A2(n14870), .ZN(n9664) );
  CLKBUF_X1 U11170 ( .A(n13777), .Z(n9665) );
  CLKBUF_X1 U11171 ( .A(n13606), .Z(n9666) );
  INV_X1 U11174 ( .A(n14198), .ZN(n9669) );
  NAND2_X1 U11175 ( .A1(n14846), .A2(n14870), .ZN(n12424) );
  XNOR2_X1 U11176 ( .A(n12357), .B(n12355), .ZN(n13777) );
  XNOR2_X1 U11177 ( .A(n12352), .B(n12351), .ZN(n13606) );
  XNOR2_X1 U11178 ( .A(n11169), .B(n11170), .ZN(n14237) );
  INV_X1 U11180 ( .A(n21123), .ZN(n9671) );
  INV_X1 U11181 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10704) );
  CLKBUF_X3 U11182 ( .A(n10624), .Z(n9708) );
  AND2_X1 U11183 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12269) );
  NAND2_X1 U11186 ( .A1(n12528), .A2(n9737), .ZN(n9952) );
  CLKBUF_X3 U11187 ( .A(n10621), .Z(n12716) );
  OR2_X1 U11188 ( .A1(n10727), .A2(n10726), .ZN(n10728) );
  INV_X1 U11189 ( .A(n12977), .ZN(n17467) );
  AND2_X1 U11190 ( .A1(n12175), .A2(n10874), .ZN(n12200) );
  INV_X1 U11192 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10223) );
  INV_X1 U11193 ( .A(n12959), .ZN(n9704) );
  INV_X4 U11194 ( .A(n17373), .ZN(n17430) );
  NAND2_X1 U11195 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18977) );
  INV_X1 U11196 ( .A(n17470), .ZN(n17488) );
  OR2_X1 U11197 ( .A1(n10182), .A2(n12197), .ZN(n19232) );
  AND2_X1 U11198 ( .A1(n16615), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12463) );
  NOR2_X1 U11199 ( .A1(n11976), .A2(n13472), .ZN(n11964) );
  OR2_X1 U11200 ( .A1(n17180), .A2(n12927), .ZN(n17429) );
  CLKBUF_X2 U11201 ( .A(n10999), .Z(n13384) );
  INV_X2 U11202 ( .A(n10648), .ZN(n12030) );
  AND2_X1 U11203 ( .A1(n15469), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15443) );
  NAND2_X1 U11204 ( .A1(n18147), .A2(n18105), .ZN(n18078) );
  NAND2_X1 U11205 ( .A1(n10072), .A2(n9772), .ZN(n13047) );
  NOR2_X2 U11206 ( .A1(n19171), .A2(n18280), .ZN(n18953) );
  INV_X1 U11207 ( .A(n20268), .ZN(n16093) );
  NAND2_X1 U11208 ( .A1(n9909), .A2(n9907), .ZN(n16815) );
  NAND2_X1 U11209 ( .A1(n18041), .A2(n18256), .ZN(n17954) );
  OAI21_X1 U11210 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19168), .A(n16815), 
        .ZN(n18147) );
  XOR2_X1 U11211 ( .A(n11164), .B(n11163), .Z(n9672) );
  INV_X2 U11212 ( .A(n14059), .ZN(n10938) );
  AND2_X1 U11213 ( .A1(n12403), .A2(n12402), .ZN(n9673) );
  AND2_X2 U11214 ( .A1(n12716), .A2(n10283), .ZN(n9717) );
  INV_X4 U11215 ( .A(n15804), .ZN(n10622) );
  OAI21_X2 U11216 ( .B1(n12280), .B2(n14025), .A(n12293), .ZN(n9696) );
  OAI21_X2 U11217 ( .B1(n9943), .B2(n9944), .A(n9790), .ZN(n15445) );
  AND2_X2 U11218 ( .A1(n12146), .A2(n10031), .ZN(n10030) );
  AND2_X1 U11220 ( .A1(n14061), .A2(n13508), .ZN(n9674) );
  AND2_X2 U11221 ( .A1(n14061), .A2(n13508), .ZN(n9675) );
  AND2_X2 U11222 ( .A1(n10653), .A2(n10652), .ZN(n12528) );
  INV_X2 U11224 ( .A(n10657), .ZN(n12465) );
  AOI22_X2 U11225 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19648), .B1(
        n19594), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11972) );
  BUF_X2 U11226 ( .A(n10943), .Z(n9680) );
  AND2_X1 U11227 ( .A1(n10906), .A2(n14061), .ZN(n10943) );
  INV_X4 U11228 ( .A(n12733), .ZN(n10621) );
  NAND4_X1 U11229 ( .A1(n19146), .A2(n19130), .A3(n19139), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9681) );
  NAND4_X1 U11230 ( .A1(n19146), .A2(n19130), .A3(n19139), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9682) );
  NOR3_X4 U11231 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n17180), .ZN(n12970) );
  NAND2_X2 U11232 ( .A1(n19146), .A2(n12924), .ZN(n17180) );
  BUF_X2 U11233 ( .A(n12473), .Z(n9683) );
  NAND2_X2 U11234 ( .A1(n10044), .A2(n11046), .ZN(n11115) );
  INV_X1 U11235 ( .A(n18004), .ZN(n17990) );
  NOR2_X2 U11236 ( .A1(n19134), .A2(n18078), .ZN(n18004) );
  CLKBUF_X1 U11237 ( .A(n15267), .Z(n15268) );
  OR2_X1 U11238 ( .A1(n13059), .A2(n18057), .ZN(n13058) );
  CLKBUF_X1 U11239 ( .A(n15323), .Z(n15335) );
  AND2_X1 U11240 ( .A1(n17812), .A2(n9748), .ZN(n10069) );
  OR2_X1 U11241 ( .A1(n13054), .A2(n10171), .ZN(n13055) );
  AND2_X1 U11242 ( .A1(n12056), .A2(n12055), .ZN(n12141) );
  AND2_X1 U11243 ( .A1(n15101), .A2(n14229), .ZN(n16270) );
  NOR2_X1 U11244 ( .A1(n18989), .A2(n16038), .ZN(n17683) );
  CLKBUF_X1 U11245 ( .A(n14091), .Z(n20698) );
  NAND2_X1 U11247 ( .A1(n10019), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18009) );
  NAND2_X1 U11248 ( .A1(n11091), .A2(n12401), .ZN(n11122) );
  AND2_X1 U11249 ( .A1(n13441), .A2(n13440), .ZN(n13443) );
  NAND2_X1 U11250 ( .A1(n9693), .A2(n11117), .ZN(n13795) );
  NAND2_X1 U11251 ( .A1(n18359), .A2(n18988), .ZN(n18280) );
  AND2_X1 U11252 ( .A1(n10011), .A2(n9788), .ZN(n13045) );
  CLKBUF_X2 U11253 ( .A(n10374), .Z(n14501) );
  INV_X1 U11254 ( .A(n18493), .ZN(n17689) );
  NAND2_X1 U11255 ( .A1(n10273), .A2(n10272), .ZN(n10647) );
  INV_X2 U11256 ( .A(n13802), .ZN(n13989) );
  NAND2_X1 U11257 ( .A1(n12983), .A2(n12982), .ZN(n17682) );
  INV_X1 U11258 ( .A(n16615), .ZN(n20199) );
  AND4_X1 U11259 ( .A1(n11025), .A2(n11024), .A3(n11023), .A4(n11022), .ZN(
        n11026) );
  AND3_X1 U11260 ( .A1(n10919), .A2(n10920), .A3(n10921), .ZN(n9971) );
  INV_X4 U11261 ( .A(n12943), .ZN(n17489) );
  CLKBUF_X2 U11262 ( .A(n11059), .Z(n11521) );
  BUF_X2 U11263 ( .A(n11093), .Z(n11697) );
  CLKBUF_X2 U11264 ( .A(n11406), .Z(n11522) );
  CLKBUF_X2 U11265 ( .A(n10948), .Z(n9711) );
  CLKBUF_X2 U11266 ( .A(n11698), .Z(n11675) );
  INV_X1 U11267 ( .A(n12959), .ZN(n9688) );
  CLKBUF_X2 U11268 ( .A(n11485), .Z(n11527) );
  AND2_X2 U11269 ( .A1(n12717), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10513) );
  BUF_X4 U11270 ( .A(n11098), .Z(n9686) );
  AND2_X1 U11271 ( .A1(n10900), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10906) );
  INV_X4 U11272 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12924) );
  INV_X1 U11273 ( .A(n15668), .ZN(n15514) );
  NAND2_X1 U11274 ( .A1(n15691), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16435) );
  NAND2_X1 U11275 ( .A1(n15691), .A2(n9956), .ZN(n15668) );
  AND2_X1 U11276 ( .A1(n15709), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16446) );
  AND2_X1 U11277 ( .A1(n14822), .A2(n14821), .ZN(n14831) );
  AND2_X2 U11278 ( .A1(n12423), .A2(n14847), .ZN(n14830) );
  OAI21_X1 U11279 ( .B1(n10166), .B2(n14653), .A(n9725), .ZN(n14874) );
  OR2_X1 U11280 ( .A1(n14823), .A2(n14820), .ZN(n14822) );
  NOR2_X1 U11281 ( .A1(n15268), .A2(n9775), .ZN(n15322) );
  NAND2_X1 U11282 ( .A1(n15742), .A2(n10145), .ZN(n15708) );
  AND2_X1 U11283 ( .A1(n15742), .A2(n10143), .ZN(n15469) );
  AND2_X2 U11284 ( .A1(n14676), .A2(n14722), .ZN(n14664) );
  CLKBUF_X1 U11285 ( .A(n14342), .Z(n9695) );
  XNOR2_X1 U11286 ( .A(n14506), .B(n14505), .ZN(n16309) );
  XNOR2_X1 U11287 ( .A(n12754), .B(n9852), .ZN(n12753) );
  OR2_X1 U11288 ( .A1(n15299), .A2(n15298), .ZN(n16314) );
  OR2_X1 U11289 ( .A1(n15307), .A2(n15296), .ZN(n16336) );
  OAI211_X1 U11290 ( .C1(n16678), .C2(n13057), .A(n13058), .B(n10003), .ZN(
        n13063) );
  INV_X1 U11291 ( .A(n9935), .ZN(n10034) );
  NAND2_X1 U11292 ( .A1(n10047), .A2(n10048), .ZN(n16169) );
  NOR2_X1 U11293 ( .A1(n15970), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13059) );
  NOR2_X1 U11294 ( .A1(n15284), .A2(n9813), .ZN(n10077) );
  AND2_X1 U11295 ( .A1(n12298), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12305) );
  AOI21_X1 U11296 ( .B1(n9731), .B2(n9942), .A(n9781), .ZN(n9937) );
  AND2_X1 U11297 ( .A1(n12205), .A2(n9947), .ZN(n9946) );
  OAI21_X1 U11298 ( .B1(n12379), .B2(n10050), .A(n16174), .ZN(n10049) );
  AOI21_X1 U11299 ( .B1(n12410), .B2(n12409), .A(n9760), .ZN(n10058) );
  NOR2_X2 U11300 ( .A1(n13974), .A2(n14145), .ZN(n14294) );
  AND2_X1 U11301 ( .A1(n12141), .A2(n12034), .ZN(n10146) );
  OR2_X1 U11302 ( .A1(n14922), .A2(n12413), .ZN(n14906) );
  OR2_X1 U11303 ( .A1(n12230), .A2(n10075), .ZN(n15151) );
  NAND2_X1 U11304 ( .A1(n9897), .A2(n12408), .ZN(n12409) );
  NAND2_X1 U11305 ( .A1(n12376), .A2(n12375), .ZN(n12378) );
  INV_X1 U11306 ( .A(n9673), .ZN(n16158) );
  OR2_X1 U11307 ( .A1(n12373), .A2(n12400), .ZN(n12376) );
  NOR2_X1 U11308 ( .A1(n12227), .A2(n12226), .ZN(n12230) );
  NOR2_X1 U11309 ( .A1(n13565), .A2(n13688), .ZN(n13687) );
  NOR2_X1 U11310 ( .A1(n14605), .A2(n14587), .ZN(n14586) );
  AND2_X1 U11311 ( .A1(n11281), .A2(n11253), .ZN(n12372) );
  XNOR2_X1 U11312 ( .A(n12403), .B(n11283), .ZN(n12390) );
  OR2_X1 U11313 ( .A1(n11989), .A2(n19541), .ZN(n12060) );
  NOR2_X1 U11314 ( .A1(n18054), .A2(n18370), .ZN(n18053) );
  OR2_X1 U11315 ( .A1(n12192), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12221) );
  CLKBUF_X1 U11316 ( .A(n11932), .Z(n14800) );
  NAND2_X1 U11317 ( .A1(n9892), .A2(n9891), .ZN(n12403) );
  AND2_X1 U11318 ( .A1(n18055), .A2(n10022), .ZN(n17868) );
  NAND2_X1 U11319 ( .A1(n12346), .A2(n12345), .ZN(n12347) );
  AND2_X1 U11320 ( .A1(n11184), .A2(n11183), .ZN(n11204) );
  OR2_X1 U11321 ( .A1(n12570), .A2(n12569), .ZN(n13465) );
  INV_X1 U11322 ( .A(n14963), .ZN(n15053) );
  NAND2_X2 U11323 ( .A1(n14743), .A2(n13702), .ZN(n14793) );
  AOI21_X1 U11324 ( .B1(n10022), .B2(n17968), .A(n18285), .ZN(n10021) );
  INV_X2 U11325 ( .A(n14743), .ZN(n14783) );
  AOI21_X1 U11326 ( .B1(n13413), .B2(n13411), .A(n12561), .ZN(n13478) );
  NAND2_X1 U11327 ( .A1(n13623), .A2(n13622), .ZN(n15101) );
  NAND2_X1 U11328 ( .A1(n11203), .A2(n11202), .ZN(n13841) );
  CLKBUF_X1 U11329 ( .A(n9714), .Z(n9721) );
  XNOR2_X1 U11330 ( .A(n11122), .B(n11120), .ZN(n11162) );
  NAND2_X1 U11331 ( .A1(n13048), .A2(n17968), .ZN(n18033) );
  NAND2_X2 U11332 ( .A1(n20324), .A2(n13384), .ZN(n14742) );
  OAI22_X1 U11333 ( .A1(n13495), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n12331), 
        .B2(n11191), .ZN(n11154) );
  XNOR2_X1 U11334 ( .A(n14079), .B(n13905), .ZN(n14132) );
  OR2_X1 U11335 ( .A1(n18953), .A2(n9793), .ZN(n9909) );
  OR2_X1 U11336 ( .A1(n11137), .A2(n11136), .ZN(n11138) );
  XNOR2_X1 U11337 ( .A(n11963), .B(n11958), .ZN(n12556) );
  NAND2_X1 U11338 ( .A1(n11137), .A2(n11136), .ZN(n14079) );
  NOR2_X1 U11339 ( .A1(n18369), .A2(n18471), .ZN(n18470) );
  AND2_X1 U11340 ( .A1(n12097), .A2(n10096), .ZN(n12155) );
  XNOR2_X1 U11341 ( .A(n9888), .B(n11126), .ZN(n20450) );
  XNOR2_X1 U11342 ( .A(n10750), .B(n10748), .ZN(n11943) );
  OAI211_X1 U11343 ( .C1(n14204), .C2(n12441), .A(n11135), .B(n11134), .ZN(
        n11136) );
  NAND2_X1 U11344 ( .A1(n18976), .A2(n13250), .ZN(n18972) );
  NAND2_X1 U11345 ( .A1(n10677), .A2(n10181), .ZN(n10726) );
  NAND2_X1 U11346 ( .A1(n10745), .A2(n10744), .ZN(n10750) );
  NAND2_X1 U11347 ( .A1(n10724), .A2(n10723), .ZN(n11953) );
  NAND2_X1 U11348 ( .A1(n10872), .A2(n10871), .ZN(n12130) );
  OR2_X1 U11349 ( .A1(n11132), .A2(n14074), .ZN(n11189) );
  NAND2_X1 U11350 ( .A1(n15934), .A2(n15933), .ZN(n13251) );
  AND4_X1 U11351 ( .A1(n10722), .A2(n10721), .A3(n10720), .A4(n10719), .ZN(
        n10723) );
  NOR2_X2 U11352 ( .A1(n18498), .A2(n17782), .ZN(n17783) );
  OR2_X2 U11353 ( .A1(n17727), .A2(n19014), .ZN(n17792) );
  AND2_X1 U11354 ( .A1(n13506), .A2(n11915), .ZN(n9700) );
  AND2_X1 U11355 ( .A1(n13506), .A2(n11915), .ZN(n13604) );
  NAND2_X1 U11356 ( .A1(n13450), .A2(n13451), .ZN(n13449) );
  NAND2_X1 U11357 ( .A1(n10699), .A2(n9734), .ZN(n9953) );
  AND3_X1 U11358 ( .A1(n10857), .A2(n10110), .A3(n12105), .ZN(n12125) );
  OAI21_X1 U11359 ( .B1(n10714), .B2(n10713), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10722) );
  NAND2_X1 U11360 ( .A1(n15935), .A2(n15933), .ZN(n16814) );
  OAI21_X1 U11361 ( .B1(n10742), .B2(n10673), .A(n10672), .ZN(n10674) );
  OAI21_X1 U11362 ( .B1(n11048), .B2(n11030), .A(n13989), .ZN(n11041) );
  AND2_X2 U11363 ( .A1(n13503), .A2(n11042), .ZN(n11906) );
  NOR2_X1 U11364 ( .A1(n12102), .A2(n10111), .ZN(n10110) );
  AND2_X2 U11365 ( .A1(n12508), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10845) );
  NAND2_X1 U11366 ( .A1(n10654), .A2(n10703), .ZN(n10742) );
  AND2_X1 U11367 ( .A1(n12501), .A2(n10686), .ZN(n10712) );
  AND3_X1 U11368 ( .A1(n10396), .A2(n10395), .A3(n10394), .ZN(n13729) );
  AND3_X1 U11369 ( .A1(n10865), .A2(n10864), .A3(n10863), .ZN(n12102) );
  AOI21_X1 U11370 ( .B1(n10005), .B2(n10004), .A(n13034), .ZN(n18111) );
  MUX2_X1 U11371 ( .A(n10357), .B(n10356), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n13451) );
  AND2_X1 U11372 ( .A1(n10002), .A2(n10342), .ZN(n10358) );
  NOR2_X1 U11373 ( .A1(n17667), .A2(n13015), .ZN(n13039) );
  AND2_X1 U11374 ( .A1(n11038), .A2(n11784), .ZN(n11723) );
  AND2_X1 U11375 ( .A1(n11034), .A2(n11052), .ZN(n10119) );
  CLKBUF_X1 U11377 ( .A(n11784), .Z(n14523) );
  AND4_X1 U11378 ( .A1(n12489), .A2(n12488), .A3(n10644), .A4(n13415), .ZN(
        n10645) );
  AND2_X1 U11379 ( .A1(n12446), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10703) );
  AND2_X2 U11380 ( .A1(n10276), .A2(n10855), .ZN(n10534) );
  AND2_X1 U11381 ( .A1(n11031), .A2(n13384), .ZN(n11052) );
  INV_X4 U11382 ( .A(n11785), .ZN(n11808) );
  NAND2_X1 U11383 ( .A1(n12866), .A2(n10276), .ZN(n10566) );
  AND2_X1 U11384 ( .A1(n12469), .A2(n13415), .ZN(n9858) );
  NAND2_X1 U11385 ( .A1(n11191), .A2(n11190), .ZN(n11740) );
  NAND2_X1 U11386 ( .A1(n10659), .A2(n10658), .ZN(n12497) );
  OR2_X1 U11388 ( .A1(n9699), .A2(n11803), .ZN(n13611) );
  AND2_X1 U11389 ( .A1(n10191), .A2(n13812), .ZN(n12342) );
  OR2_X1 U11390 ( .A1(n10390), .A2(n10389), .ZN(n12031) );
  OR2_X1 U11391 ( .A1(n12969), .A2(n12968), .ZN(n13016) );
  AND2_X1 U11392 ( .A1(n12950), .A2(n12949), .ZN(n17667) );
  AND2_X1 U11393 ( .A1(n10647), .A2(n19920), .ZN(n10276) );
  OR2_X1 U11394 ( .A1(n10327), .A2(n10326), .ZN(n16586) );
  NAND2_X1 U11395 ( .A1(n9844), .A2(n9839), .ZN(n10642) );
  INV_X1 U11396 ( .A(n10647), .ZN(n9687) );
  INV_X2 U11397 ( .A(U212), .ZN(n16764) );
  INV_X2 U11398 ( .A(n16707), .ZN(n16767) );
  CLKBUF_X2 U11399 ( .A(n10641), .Z(n19565) );
  AND4_X1 U11400 ( .A1(n12981), .A2(n12980), .A3(n12979), .A4(n12978), .ZN(
        n12982) );
  NAND4_X2 U11401 ( .A1(n10996), .A2(n10995), .A3(n10994), .A4(n10993), .ZN(
        n13802) );
  OR2_X1 U11402 ( .A1(n10976), .A2(n10975), .ZN(n10999) );
  NOR2_X1 U11403 ( .A1(n10914), .A2(n10913), .ZN(n10191) );
  AND4_X1 U11404 ( .A1(n11020), .A2(n11019), .A3(n11018), .A4(n11017), .ZN(
        n11027) );
  AND4_X1 U11405 ( .A1(n11016), .A2(n11015), .A3(n11014), .A4(n11013), .ZN(
        n11028) );
  AND4_X1 U11406 ( .A1(n11012), .A2(n11011), .A3(n11010), .A4(n11009), .ZN(
        n11029) );
  AND4_X1 U11407 ( .A1(n10992), .A2(n10991), .A3(n10990), .A4(n10989), .ZN(
        n10993) );
  AND4_X1 U11408 ( .A1(n10988), .A2(n10987), .A3(n10986), .A4(n10985), .ZN(
        n10994) );
  AND4_X1 U11409 ( .A1(n10984), .A2(n10983), .A3(n10982), .A4(n10981), .ZN(
        n10995) );
  AND4_X1 U11410 ( .A1(n10980), .A2(n10979), .A3(n10978), .A4(n10977), .ZN(
        n10996) );
  AND4_X1 U11411 ( .A1(n10947), .A2(n10946), .A3(n10945), .A4(n10944), .ZN(
        n10964) );
  AND4_X1 U11412 ( .A1(n10956), .A2(n10955), .A3(n10954), .A4(n10953), .ZN(
        n10962) );
  NOR2_X1 U11413 ( .A1(n16486), .A2(n10204), .ZN(n10207) );
  NAND2_X2 U11414 ( .A1(n19116), .A2(n19047), .ZN(n19101) );
  AND2_X2 U11415 ( .A1(n9712), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10348) );
  AND2_X1 U11416 ( .A1(n10608), .A2(n10607), .ZN(n10612) );
  AND4_X1 U11417 ( .A1(n10952), .A2(n10951), .A3(n10950), .A4(n10949), .ZN(
        n10963) );
  INV_X1 U11418 ( .A(n9755), .ZN(n17448) );
  CLKBUF_X3 U11419 ( .A(n12849), .Z(n9712) );
  INV_X2 U11420 ( .A(n12984), .ZN(n17288) );
  NOR2_X1 U11421 ( .A1(n19134), .A2(n18148), .ZN(n19166) );
  AND2_X2 U11422 ( .A1(n12830), .A2(n10282), .ZN(n12678) );
  INV_X1 U11423 ( .A(n10200), .ZN(n9959) );
  INV_X2 U11424 ( .A(n19181), .ZN(n19116) );
  AND2_X2 U11425 ( .A1(n10622), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10397) );
  AND2_X2 U11426 ( .A1(n12717), .A2(n10283), .ZN(n10514) );
  INV_X2 U11427 ( .A(n16804), .ZN(n16806) );
  BUF_X2 U11428 ( .A(n10624), .Z(n9709) );
  INV_X2 U11429 ( .A(n20916), .ZN(n20875) );
  NOR2_X1 U11430 ( .A1(n19134), .A2(n19030), .ZN(n17173) );
  AND2_X2 U11431 ( .A1(n10906), .A2(n14062), .ZN(n11098) );
  BUF_X2 U11432 ( .A(n10624), .Z(n9707) );
  AND2_X4 U11433 ( .A1(n10907), .A2(n14062), .ZN(n10970) );
  AND2_X2 U11434 ( .A1(n14064), .A2(n13508), .ZN(n11072) );
  INV_X4 U11435 ( .A(n17429), .ZN(n9689) );
  NAND3_X1 U11436 ( .A1(n9993), .A2(n9992), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10277) );
  OR3_X1 U11437 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18974), .ZN(n17373) );
  NAND2_X2 U11438 ( .A1(n12924), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12926) );
  AND2_X2 U11439 ( .A1(n14061), .A2(n10908), .ZN(n11485) );
  NOR2_X1 U11441 ( .A1(n16507), .A2(n9961), .ZN(n9960) );
  INV_X1 U11442 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10282) );
  CLKBUF_X1 U11445 ( .A(n10030), .Z(n9691) );
  AOI21_X2 U11446 ( .B1(n13049), .B2(n17969), .A(n18057), .ZN(n17941) );
  NOR2_X1 U11447 ( .A1(n10656), .A2(n10632), .ZN(n12473) );
  INV_X2 U11448 ( .A(n10277), .ZN(n10609) );
  INV_X1 U11449 ( .A(n10277), .ZN(n12849) );
  AND2_X2 U11450 ( .A1(n9853), .A2(n19565), .ZN(n12495) );
  INV_X1 U11451 ( .A(n15975), .ZN(n9692) );
  XOR2_X1 U11452 ( .A(n9888), .B(n11126), .Z(n9693) );
  NAND2_X1 U11453 ( .A1(n11000), .A2(n10190), .ZN(n15974) );
  NAND2_X1 U11454 ( .A1(n9889), .A2(n11110), .ZN(n9888) );
  OAI21_X2 U11455 ( .B1(n11113), .B2(n11112), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11126) );
  NOR2_X2 U11456 ( .A1(n13435), .A2(n13433), .ZN(n13434) );
  INV_X1 U11457 ( .A(n15808), .ZN(n9694) );
  OR2_X1 U11458 ( .A1(n10090), .A2(n10091), .ZN(n9697) );
  NAND2_X1 U11459 ( .A1(n9697), .A2(n12294), .ZN(n12280) );
  INV_X2 U11460 ( .A(n15599), .ZN(n10085) );
  NAND2_X2 U11461 ( .A1(n12164), .A2(n12163), .ZN(n15715) );
  AND4_X1 U11462 ( .A1(n11986), .A2(n11985), .A3(n11984), .A4(n11983), .ZN(
        n11995) );
  NAND2_X1 U11463 ( .A1(n15535), .A2(n15534), .ZN(n15533) );
  INV_X1 U11464 ( .A(n12142), .ZN(n12140) );
  XNOR2_X1 U11465 ( .A(n12142), .B(n12141), .ZN(n12298) );
  XNOR2_X1 U11466 ( .A(n17682), .B(n13031), .ZN(n18138) );
  AND2_X2 U11467 ( .A1(n9850), .A2(n13948), .ZN(n12575) );
  NAND2_X2 U11468 ( .A1(n12800), .A2(n12799), .ZN(n15247) );
  NAND2_X1 U11469 ( .A1(n11043), .A2(n13604), .ZN(n9698) );
  NAND2_X1 U11470 ( .A1(n11035), .A2(n9710), .ZN(n9699) );
  NAND2_X1 U11471 ( .A1(n11043), .A2(n9700), .ZN(n10043) );
  NAND3_X1 U11472 ( .A1(n9691), .A2(n15536), .A3(n12145), .ZN(n9701) );
  CLKBUF_X1 U11473 ( .A(n14021), .Z(n9702) );
  NAND3_X1 U11474 ( .A1(n10030), .A2(n15536), .A3(n12145), .ZN(n10029) );
  INV_X1 U11475 ( .A(n12339), .ZN(n11163) );
  AOI21_X1 U11476 ( .B1(n12339), .B2(n11162), .A(n11123), .ZN(n11183) );
  AND2_X1 U11477 ( .A1(n11115), .A2(n11114), .ZN(n11116) );
  AND2_X1 U11478 ( .A1(n14064), .A2(n10906), .ZN(n11059) );
  AND4_X1 U11479 ( .A1(n10960), .A2(n10959), .A3(n10958), .A4(n10957), .ZN(
        n10961) );
  INV_X1 U11481 ( .A(n14059), .ZN(n9703) );
  NAND2_X2 U11482 ( .A1(n10246), .A2(n10247), .ZN(n10655) );
  OR2_X1 U11483 ( .A1(n12865), .A2(n10657), .ZN(n12469) );
  OR2_X1 U11484 ( .A1(n12927), .A2(n12926), .ZN(n12959) );
  AOI21_X1 U11485 ( .B1(n15503), .B2(n15500), .A(n15501), .ZN(n15491) );
  OR2_X2 U11486 ( .A1(n14091), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9773) );
  NOR2_X2 U11487 ( .A1(n16389), .A2(n16391), .ZN(n16390) );
  NOR2_X2 U11488 ( .A1(n16532), .A2(n9814), .ZN(n14366) );
  NOR2_X2 U11489 ( .A1(n16383), .A2(n16382), .ZN(n16381) );
  NOR2_X2 U11490 ( .A1(n16390), .A2(n12707), .ZN(n16383) );
  AND3_X2 U11491 ( .A1(n10029), .A2(n10034), .A3(n10027), .ZN(n12164) );
  INV_X2 U11492 ( .A(n10647), .ZN(n10648) );
  BUF_X8 U11493 ( .A(n10970), .Z(n9706) );
  AND2_X1 U11494 ( .A1(n10680), .A2(n10632), .ZN(n12865) );
  AND2_X2 U11495 ( .A1(n10339), .A2(n10338), .ZN(n10680) );
  NAND2_X2 U11496 ( .A1(n10614), .A2(n10613), .ZN(n10657) );
  NOR2_X2 U11497 ( .A1(n16381), .A2(n12731), .ZN(n12754) );
  XNOR2_X2 U11498 ( .A(n12706), .B(n12704), .ZN(n16389) );
  OR2_X2 U11499 ( .A1(n12092), .A2(n12302), .ZN(n12309) );
  OAI211_X2 U11500 ( .C1(n12889), .C2(n12888), .A(n12887), .B(n15375), .ZN(
        n12896) );
  INV_X1 U11501 ( .A(n10191), .ZN(n11036) );
  NAND2_X1 U11502 ( .A1(n10191), .A2(n11037), .ZN(n14060) );
  NAND2_X2 U11503 ( .A1(n11906), .A2(n13596), .ZN(n13506) );
  NAND2_X2 U11504 ( .A1(n13238), .A2(n13641), .ZN(n16532) );
  NOR2_X4 U11505 ( .A1(n13446), .A2(n13237), .ZN(n13238) );
  XNOR2_X2 U11506 ( .A(n11962), .B(n11961), .ZN(n9714) );
  XNOR2_X2 U11507 ( .A(n11155), .B(n11184), .ZN(n12329) );
  OAI211_X1 U11508 ( .C1(n10057), .C2(n14391), .A(n10055), .B(n9738), .ZN(
        n9893) );
  NAND2_X2 U11509 ( .A1(n14830), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14841) );
  BUF_X4 U11510 ( .A(n11002), .Z(n9710) );
  NAND4_X2 U11511 ( .A1(n10962), .A2(n10963), .A3(n10964), .A4(n10961), .ZN(
        n11002) );
  NAND2_X2 U11512 ( .A1(n13971), .A2(n12579), .ZN(n14142) );
  AND2_X1 U11513 ( .A1(n14064), .A2(n10908), .ZN(n10948) );
  NAND2_X2 U11514 ( .A1(n10998), .A2(n11002), .ZN(n11032) );
  INV_X1 U11515 ( .A(n9722), .ZN(n9713) );
  OR2_X1 U11516 ( .A1(n11132), .A2(n11133), .ZN(n11135) );
  BUF_X4 U11517 ( .A(n11098), .Z(n11633) );
  INV_X4 U11518 ( .A(n9719), .ZN(n10855) );
  NAND2_X2 U11519 ( .A1(n14897), .A2(n14896), .ZN(n14879) );
  XNOR2_X2 U11520 ( .A(n10726), .B(n10725), .ZN(n11957) );
  AOI211_X2 U11521 ( .C1(n19537), .C2(n19254), .A(n15676), .B(n15675), .ZN(
        n15678) );
  OAI21_X2 U11522 ( .B1(n12306), .B2(n12162), .A(n14120), .ZN(n14345) );
  NOR2_X4 U11523 ( .A1(n13923), .A2(n12578), .ZN(n13971) );
  NAND2_X2 U11524 ( .A1(n12577), .A2(n12576), .ZN(n13923) );
  NOR2_X2 U11525 ( .A1(n13727), .A2(n13729), .ZN(n13945) );
  NOR2_X4 U11526 ( .A1(n14612), .A2(n14614), .ZN(n14602) );
  INV_X1 U11527 ( .A(n9672), .ZN(n9715) );
  INV_X1 U11528 ( .A(n9672), .ZN(n9716) );
  AND2_X1 U11529 ( .A1(n12716), .A2(n10283), .ZN(n9718) );
  AND2_X1 U11530 ( .A1(n13802), .A2(n13992), .ZN(n11791) );
  AND3_X2 U11531 ( .A1(n10221), .A2(n10222), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10624) );
  BUF_X4 U11532 ( .A(n10643), .Z(n9720) );
  INV_X1 U11533 ( .A(n10632), .ZN(n10643) );
  AND2_X2 U11534 ( .A1(n14299), .A2(n10153), .ZN(n12706) );
  NOR2_X4 U11535 ( .A1(n14142), .A2(n14292), .ZN(n14299) );
  BUF_X4 U11536 ( .A(n9714), .Z(n9722) );
  NOR2_X1 U11537 ( .A1(n18498), .A2(n17782), .ZN(n9723) );
  AOI211_X2 U11538 ( .C1(n15895), .C2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n13087), .B(n13086), .ZN(n18498) );
  AND4_X1 U11539 ( .A1(n10308), .A2(n10307), .A3(n10306), .A4(n10305), .ZN(
        n10309) );
  NAND2_X1 U11540 ( .A1(n11204), .A2(n10121), .ZN(n11252) );
  AND2_X1 U11541 ( .A1(n13841), .A2(n11238), .ZN(n10121) );
  NOR2_X2 U11542 ( .A1(n11001), .A2(n20806), .ZN(n11396) );
  AOI21_X1 U11543 ( .B1(n10621), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(n9994), .ZN(n10230) );
  NOR2_X1 U11544 ( .A1(n10277), .A2(n9995), .ZN(n9994) );
  INV_X1 U11545 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11991) );
  NAND2_X1 U11546 ( .A1(n9842), .A2(n9778), .ZN(n9837) );
  NAND2_X1 U11547 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n9842) );
  NAND2_X1 U11548 ( .A1(n10609), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n9843) );
  AND2_X1 U11549 ( .A1(n11274), .A2(n11273), .ZN(n11280) );
  OAI211_X1 U11550 ( .C1(n13180), .C2(n13166), .A(n9913), .B(n9912), .ZN(n9911) );
  NAND2_X1 U11551 ( .A1(n9914), .A2(n18509), .ZN(n9913) );
  NAND2_X1 U11552 ( .A1(n13163), .A2(n13178), .ZN(n9912) );
  NOR2_X1 U11553 ( .A1(n14710), .A2(n10125), .ZN(n10124) );
  INV_X1 U11554 ( .A(n14666), .ZN(n10125) );
  INV_X1 U11555 ( .A(n11713), .ZN(n11688) );
  INV_X1 U11556 ( .A(n14732), .ZN(n10134) );
  NOR2_X1 U11557 ( .A1(n9673), .A2(n9809), .ZN(n9897) );
  NAND2_X1 U11558 ( .A1(n11785), .A2(n9684), .ZN(n11898) );
  INV_X1 U11559 ( .A(n14060), .ZN(n11780) );
  NAND2_X1 U11560 ( .A1(n20450), .A2(n11116), .ZN(n11128) );
  OR2_X1 U11561 ( .A1(n10583), .A2(n10581), .ZN(n10571) );
  INV_X1 U11562 ( .A(n10856), .ZN(n10111) );
  NAND2_X1 U11563 ( .A1(n12267), .A2(n10855), .ZN(n10857) );
  NAND2_X1 U11564 ( .A1(n10240), .A2(n10282), .ZN(n10247) );
  INV_X1 U11565 ( .A(n12497), .ZN(n12491) );
  INV_X1 U11566 ( .A(n15332), .ZN(n9997) );
  AND4_X1 U11567 ( .A1(n10300), .A2(n10299), .A3(n10298), .A4(n10297), .ZN(
        n10311) );
  AND4_X1 U11568 ( .A1(n10296), .A2(n10295), .A3(n10294), .A4(n10293), .ZN(
        n10312) );
  NAND2_X1 U11569 ( .A1(n12091), .A2(n12090), .ZN(n12302) );
  NAND2_X1 U11570 ( .A1(n12568), .A2(n12567), .ZN(n12570) );
  AND2_X1 U11571 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12569) );
  NOR2_X1 U11572 ( .A1(n19130), .A2(n12922), .ZN(n12956) );
  AND2_X1 U11573 ( .A1(n10070), .A2(n18200), .ZN(n10015) );
  NOR2_X1 U11574 ( .A1(n17660), .A2(n13041), .ZN(n13043) );
  OAI21_X1 U11575 ( .B1(n13075), .B2(n13074), .A(n13184), .ZN(n13253) );
  NAND2_X1 U11576 ( .A1(n9862), .A2(n15940), .ZN(n16036) );
  NAND2_X1 U11577 ( .A1(n9864), .A2(n9863), .ZN(n9862) );
  NAND2_X1 U11578 ( .A1(n17729), .A2(n19171), .ZN(n9863) );
  NAND2_X1 U11579 ( .A1(n16082), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13990) );
  INV_X1 U11580 ( .A(n14107), .ZN(n11261) );
  NOR2_X1 U11581 ( .A1(n12427), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9896) );
  INV_X1 U11582 ( .A(n12428), .ZN(n9895) );
  INV_X1 U11583 ( .A(n10061), .ZN(n10060) );
  AND2_X1 U11584 ( .A1(n9659), .A2(n16608), .ZN(n13344) );
  NOR2_X1 U11585 ( .A1(n12511), .A2(n12510), .ZN(n16607) );
  NOR2_X2 U11586 ( .A1(n15430), .A2(n15275), .ZN(n15277) );
  AOI21_X1 U11587 ( .B1(n10085), .B2(n9768), .A(n15391), .ZN(n9934) );
  AND2_X1 U11588 ( .A1(n12487), .A2(n13350), .ZN(n12538) );
  INV_X1 U11589 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19920) );
  OAI22_X1 U11590 ( .A1(n15942), .A2(n15943), .B1(n15908), .B2(n15907), .ZN(
        n16034) );
  INV_X2 U11591 ( .A(n12977), .ZN(n17431) );
  NAND2_X1 U11592 ( .A1(n17897), .A2(n10015), .ZN(n10018) );
  AND2_X1 U11593 ( .A1(n13344), .A2(n13350), .ZN(n20198) );
  NAND2_X1 U11594 ( .A1(n12467), .A2(n12278), .ZN(n13269) );
  OR2_X1 U11595 ( .A1(n19757), .A2(n12007), .ZN(n9856) );
  INV_X1 U11596 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11967) );
  NAND2_X1 U11597 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n9840) );
  NAND2_X1 U11598 ( .A1(n9847), .A2(n9777), .ZN(n9835) );
  NAND2_X1 U11599 ( .A1(n11731), .A2(n11730), .ZN(n11736) );
  NAND2_X1 U11600 ( .A1(n11227), .A2(n11226), .ZN(n11238) );
  NOR2_X1 U11601 ( .A1(n10901), .A2(n20222), .ZN(n9890) );
  INV_X1 U11602 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9993) );
  AND2_X1 U11603 ( .A1(n15464), .A2(n10178), .ZN(n12199) );
  NAND2_X1 U11604 ( .A1(n11998), .A2(n11997), .ZN(n10087) );
  NAND2_X1 U11605 ( .A1(n10834), .A2(n10704), .ZN(n9861) );
  NAND2_X1 U11606 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10594) );
  NAND2_X1 U11607 ( .A1(n9712), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n10595) );
  INV_X1 U11608 ( .A(n9875), .ZN(n9874) );
  NAND2_X1 U11609 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n9873) );
  NAND2_X1 U11610 ( .A1(n13039), .A2(n13188), .ZN(n13041) );
  NAND2_X1 U11611 ( .A1(n13035), .A2(n13190), .ZN(n13015) );
  NAND2_X1 U11612 ( .A1(n14573), .A2(n10132), .ZN(n10131) );
  INV_X1 U11613 ( .A(n14591), .ZN(n10132) );
  NAND2_X1 U11614 ( .A1(n14452), .A2(n11357), .ZN(n14436) );
  AND2_X1 U11615 ( .A1(n14277), .A2(n14324), .ZN(n10120) );
  INV_X1 U11616 ( .A(n11396), .ZN(n11420) );
  NOR2_X1 U11617 ( .A1(n14713), .A2(n9986), .ZN(n9985) );
  INV_X1 U11618 ( .A(n14656), .ZN(n9986) );
  INV_X1 U11619 ( .A(n12409), .ZN(n10056) );
  OR2_X1 U11620 ( .A1(n11071), .A2(n11070), .ZN(n12404) );
  NOR2_X1 U11621 ( .A1(n11089), .A2(n20222), .ZN(n11090) );
  NAND2_X1 U11622 ( .A1(n11035), .A2(n12404), .ZN(n11089) );
  NAND2_X1 U11623 ( .A1(n11035), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11191) );
  NAND2_X1 U11624 ( .A1(n10043), .A2(n10042), .ZN(n10044) );
  NAND2_X1 U11625 ( .A1(n11128), .A2(n11127), .ZN(n11137) );
  OR2_X1 U11626 ( .A1(n11126), .A2(n11125), .ZN(n11127) );
  INV_X1 U11627 ( .A(n14089), .ZN(n14311) );
  NOR2_X1 U11628 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16631) );
  AND2_X1 U11629 ( .A1(n10870), .A2(n10869), .ZN(n12124) );
  INV_X1 U11630 ( .A(n10674), .ZN(n10676) );
  AND2_X1 U11631 ( .A1(n19578), .A2(n12550), .ZN(n12797) );
  AND2_X1 U11632 ( .A1(n9801), .A2(n10154), .ZN(n10153) );
  INV_X1 U11633 ( .A(n15345), .ZN(n10154) );
  AND2_X1 U11634 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13948) );
  AND2_X1 U11635 ( .A1(n9802), .A2(n10113), .ZN(n10112) );
  INV_X1 U11636 ( .A(n14431), .ZN(n10113) );
  INV_X1 U11637 ( .A(n12308), .ZN(n10142) );
  INV_X1 U11638 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9961) );
  NAND2_X1 U11639 ( .A1(n15260), .A2(n10108), .ZN(n10107) );
  INV_X1 U11640 ( .A(n15251), .ZN(n10108) );
  NOR2_X1 U11641 ( .A1(n15597), .A2(n15393), .ZN(n10084) );
  INV_X1 U11642 ( .A(n15175), .ZN(n10079) );
  NOR2_X1 U11643 ( .A1(n12318), .A2(n10144), .ZN(n10143) );
  INV_X1 U11644 ( .A(n10145), .ZN(n10144) );
  NAND2_X1 U11645 ( .A1(n10000), .A2(n15693), .ZN(n9999) );
  INV_X1 U11646 ( .A(n16533), .ZN(n10000) );
  AND2_X1 U11647 ( .A1(n15717), .A2(n15714), .ZN(n15454) );
  NOR2_X1 U11648 ( .A1(n10433), .A2(n10432), .ZN(n12089) );
  OR2_X1 U11649 ( .A1(n11960), .A2(n11941), .ZN(n11942) );
  AND2_X1 U11650 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12551) );
  AND2_X1 U11651 ( .A1(n12494), .A2(n10651), .ZN(n10652) );
  AND2_X1 U11652 ( .A1(n9683), .A2(n10647), .ZN(n10649) );
  NAND3_X1 U11653 ( .A1(n10634), .A2(n12472), .A3(n10633), .ZN(n10683) );
  NAND2_X1 U11654 ( .A1(n9954), .A2(n9955), .ZN(n11989) );
  AND2_X1 U11655 ( .A1(n19559), .A2(n13423), .ZN(n9955) );
  NAND2_X1 U11656 ( .A1(n19139), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12927) );
  NAND2_X1 U11657 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10067) );
  INV_X1 U11658 ( .A(n12989), .ZN(n10068) );
  INV_X1 U11659 ( .A(n12990), .ZN(n10065) );
  NOR2_X1 U11660 ( .A1(n12921), .A2(n17180), .ZN(n13023) );
  NOR2_X1 U11661 ( .A1(n18143), .A2(n9928), .ZN(n9927) );
  AND2_X1 U11662 ( .A1(n10015), .A2(n10017), .ZN(n10014) );
  NAND2_X1 U11663 ( .A1(n18057), .A2(n18180), .ZN(n10017) );
  XNOR2_X1 U11664 ( .A(n13015), .B(n10063), .ZN(n13037) );
  INV_X1 U11665 ( .A(n17667), .ZN(n10063) );
  XNOR2_X1 U11666 ( .A(n13016), .B(n17682), .ZN(n13033) );
  INV_X1 U11667 ( .A(n9911), .ZN(n9910) );
  AND2_X1 U11668 ( .A1(n14564), .A2(n14574), .ZN(n9990) );
  INV_X1 U11669 ( .A(n13597), .ZN(n13521) );
  AND2_X1 U11670 ( .A1(n13504), .A2(n11725), .ZN(n13622) );
  OAI21_X1 U11671 ( .B1(n13374), .B2(n11918), .A(n11917), .ZN(n13529) );
  OR2_X1 U11672 ( .A1(n11690), .A2(n14815), .ZN(n11691) );
  OR2_X1 U11673 ( .A1(n11691), .A2(n14811), .ZN(n12439) );
  AND2_X1 U11674 ( .A1(n14602), .A2(n10126), .ZN(n14562) );
  NOR2_X1 U11675 ( .A1(n10128), .A2(n10127), .ZN(n10126) );
  INV_X1 U11676 ( .A(n10185), .ZN(n10127) );
  NAND2_X1 U11677 ( .A1(n10130), .A2(n10129), .ZN(n10128) );
  NAND2_X1 U11678 ( .A1(n11648), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11690) );
  NAND2_X1 U11679 ( .A1(n11606), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11646) );
  NAND2_X1 U11680 ( .A1(n9894), .A2(n9831), .ZN(n12420) );
  INV_X1 U11681 ( .A(n14897), .ZN(n9894) );
  AND2_X1 U11682 ( .A1(n11501), .A2(n11500), .ZN(n14666) );
  AND2_X1 U11683 ( .A1(n11481), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11482) );
  INV_X1 U11684 ( .A(n14686), .ZN(n10136) );
  INV_X1 U11685 ( .A(n14437), .ZN(n10135) );
  NAND2_X1 U11686 ( .A1(n11279), .A2(n11278), .ZN(n14152) );
  AND2_X1 U11687 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n11231), .ZN(
        n11254) );
  INV_X1 U11688 ( .A(n13790), .ZN(n11236) );
  AOI21_X1 U11689 ( .B1(n12372), .B2(n11396), .A(n11260), .ZN(n14107) );
  NAND2_X1 U11690 ( .A1(n13694), .A2(n11182), .ZN(n13645) );
  OR2_X1 U11691 ( .A1(n20897), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12441) );
  NAND2_X1 U11692 ( .A1(n12359), .A2(n12358), .ZN(n13929) );
  AND2_X1 U11693 ( .A1(n13623), .A2(n13614), .ZN(n14961) );
  INV_X1 U11694 ( .A(n11032), .ZN(n11000) );
  NAND2_X1 U11695 ( .A1(n9901), .A2(n9900), .ZN(n9899) );
  INV_X1 U11696 ( .A(n13508), .ZN(n9901) );
  INV_X1 U11697 ( .A(n10908), .ZN(n9900) );
  INV_X1 U11698 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14074) );
  AND2_X1 U11699 ( .A1(n13794), .A2(n15112), .ZN(n20413) );
  AND2_X1 U11700 ( .A1(n14097), .A2(n13903), .ZN(n20549) );
  INV_X1 U11701 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20661) );
  INV_X1 U11702 ( .A(n20698), .ZN(n20616) );
  AND2_X1 U11703 ( .A1(n14097), .A2(n13841), .ZN(n20747) );
  INV_X1 U11704 ( .A(n20545), .ZN(n20748) );
  NOR2_X1 U11705 ( .A1(n13521), .A2(n16023), .ZN(n15999) );
  NAND2_X1 U11706 ( .A1(n10854), .A2(n10853), .ZN(n12267) );
  NAND2_X1 U11707 ( .A1(n10885), .A2(n10852), .ZN(n10853) );
  NAND2_X1 U11708 ( .A1(n12289), .A2(n12537), .ZN(n10854) );
  AND2_X1 U11709 ( .A1(n12230), .A2(n10879), .ZN(n12233) );
  AND2_X1 U11710 ( .A1(n9764), .A2(n10097), .ZN(n10096) );
  NAND2_X1 U11711 ( .A1(n12097), .A2(n10873), .ZN(n12099) );
  NAND2_X1 U11712 ( .A1(n12803), .A2(n10159), .ZN(n10158) );
  INV_X1 U11713 ( .A(n15257), .ZN(n10159) );
  INV_X1 U11714 ( .A(n15247), .ZN(n9854) );
  AND3_X1 U11715 ( .A1(n10537), .A2(n10536), .A3(n10535), .ZN(n14042) );
  AND2_X1 U11716 ( .A1(n13946), .A2(n14047), .ZN(n9996) );
  NOR2_X1 U11717 ( .A1(n10218), .A2(n15379), .ZN(n10219) );
  NOR2_X1 U11718 ( .A1(n15285), .A2(n15286), .ZN(n10807) );
  OR2_X1 U11719 ( .A1(n14492), .A2(n14493), .ZN(n14495) );
  NOR2_X1 U11720 ( .A1(n14495), .A2(n13543), .ZN(n13567) );
  AOI21_X1 U11721 ( .B1(n11940), .B2(n9735), .A(n9785), .ZN(n10081) );
  NAND2_X1 U11722 ( .A1(n10085), .A2(n9733), .ZN(n15419) );
  INV_X1 U11723 ( .A(n15612), .ZN(n9998) );
  OR2_X1 U11724 ( .A1(n12253), .A2(n12252), .ZN(n15595) );
  OR2_X1 U11725 ( .A1(n15142), .A2(n15428), .ZN(n15430) );
  INV_X1 U11726 ( .A(n15435), .ZN(n9942) );
  AOI21_X1 U11727 ( .B1(n15435), .B2(n9941), .A(n9765), .ZN(n9940) );
  INV_X1 U11728 ( .A(n15446), .ZN(n9941) );
  INV_X1 U11729 ( .A(n9946), .ZN(n9944) );
  NAND2_X1 U11730 ( .A1(n10100), .A2(n14009), .ZN(n10099) );
  INV_X1 U11731 ( .A(n10102), .ZN(n10100) );
  AND3_X1 U11732 ( .A1(n10292), .A2(n10291), .A3(n10290), .ZN(n13435) );
  NOR2_X1 U11733 ( .A1(n10033), .A2(n10032), .ZN(n10031) );
  INV_X1 U11734 ( .A(n15540), .ZN(n10033) );
  OAI21_X1 U11735 ( .B1(n14345), .B2(n12150), .A(n9936), .ZN(n9935) );
  AND2_X1 U11736 ( .A1(n15539), .A2(n15756), .ZN(n9936) );
  NAND2_X1 U11737 ( .A1(n12304), .A2(n12303), .ZN(n14343) );
  NAND2_X1 U11738 ( .A1(n16498), .A2(n9736), .ZN(n12300) );
  INV_X1 U11739 ( .A(n12508), .ZN(n15789) );
  AOI21_X1 U11740 ( .B1(n12556), .B2(n12562), .A(n12555), .ZN(n13413) );
  OR2_X1 U11741 ( .A1(n13467), .A2(n13466), .ZN(n13477) );
  OR2_X1 U11742 ( .A1(n20154), .A2(n20177), .ZN(n19695) );
  INV_X1 U11743 ( .A(n19596), .ZN(n19820) );
  NAND2_X1 U11744 ( .A1(n15796), .A2(n20166), .ZN(n19696) );
  INV_X1 U11745 ( .A(n12060), .ZN(n14164) );
  INV_X1 U11746 ( .A(n12549), .ZN(n19578) );
  NAND2_X1 U11747 ( .A1(n13747), .A2(n20201), .ZN(n19915) );
  OR2_X1 U11748 ( .A1(n16634), .A2(n13746), .ZN(n13747) );
  INV_X1 U11749 ( .A(n19915), .ZN(n19995) );
  AND2_X1 U11750 ( .A1(n20184), .A2(n10587), .ZN(n16608) );
  NOR2_X1 U11751 ( .A1(n12466), .A2(n12464), .ZN(n13745) );
  NOR2_X1 U11752 ( .A1(n20184), .A2(n13393), .ZN(n12464) );
  OR2_X1 U11753 ( .A1(n18974), .A2(n12921), .ZN(n9756) );
  AOI21_X1 U11754 ( .B1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B2(n17465), .A(
        n13022), .ZN(n13028) );
  AOI21_X1 U11755 ( .B1(n16036), .B2(n16035), .A(n19020), .ZN(n17537) );
  NAND2_X1 U11756 ( .A1(n18525), .A2(n17538), .ZN(n18989) );
  INV_X1 U11757 ( .A(n17537), .ZN(n16038) );
  INV_X1 U11758 ( .A(n18498), .ZN(n19171) );
  NAND2_X1 U11759 ( .A1(n10071), .A2(n9762), .ZN(n10070) );
  NAND2_X1 U11760 ( .A1(n17868), .A2(n13052), .ZN(n10071) );
  NAND2_X1 U11761 ( .A1(n17885), .A2(n18196), .ZN(n17858) );
  OAI21_X1 U11762 ( .B1(n18056), .B2(n10023), .A(n10021), .ZN(n10024) );
  NAND2_X1 U11763 ( .A1(n18055), .A2(n13047), .ZN(n17979) );
  INV_X1 U11764 ( .A(n13047), .ZN(n13048) );
  NAND2_X1 U11765 ( .A1(n10072), .A2(n10020), .ZN(n10019) );
  INV_X1 U11766 ( .A(n13046), .ZN(n10020) );
  NAND2_X1 U11767 ( .A1(n18056), .A2(n18057), .ZN(n18055) );
  NAND2_X1 U11768 ( .A1(n18088), .A2(n10009), .ZN(n10008) );
  NAND2_X1 U11769 ( .A1(n10010), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10009) );
  INV_X1 U11770 ( .A(n18089), .ZN(n10010) );
  NAND2_X1 U11771 ( .A1(n18089), .A2(n13040), .ZN(n10007) );
  NOR2_X1 U11772 ( .A1(n15956), .A2(n15937), .ZN(n16689) );
  OR2_X1 U11773 ( .A1(n18137), .A2(n13032), .ZN(n10004) );
  INV_X1 U11774 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18443) );
  NOR2_X1 U11775 ( .A1(n18138), .A2(n18145), .ZN(n18137) );
  NAND2_X1 U11776 ( .A1(n13171), .A2(n13172), .ZN(n13250) );
  AOI21_X1 U11777 ( .B1(n13077), .B2(n13076), .A(n13253), .ZN(n18957) );
  INV_X1 U11778 ( .A(n13174), .ZN(n18525) );
  NOR2_X1 U11779 ( .A1(n13802), .A2(n13992), .ZN(n13371) );
  NAND2_X1 U11780 ( .A1(n16008), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20219) );
  NAND2_X1 U11781 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20906) );
  OR2_X1 U11782 ( .A1(n20904), .A2(n13983), .ZN(n16082) );
  INV_X1 U11783 ( .A(n16059), .ZN(n14782) );
  INV_X1 U11784 ( .A(n16181), .ZN(n16180) );
  AND2_X1 U11785 ( .A1(n12436), .A2(n20696), .ZN(n14887) );
  XNOR2_X1 U11786 ( .A(n10040), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14971) );
  NAND2_X1 U11787 ( .A1(n12430), .A2(n10041), .ZN(n10040) );
  NAND2_X1 U11788 ( .A1(n9895), .A2(n9744), .ZN(n10041) );
  NOR2_X2 U11789 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20696) );
  AND2_X1 U11790 ( .A1(n13985), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16008) );
  AND3_X1 U11791 ( .A1(n16608), .A2(n10654), .A3(n12278), .ZN(n13275) );
  NAND2_X1 U11792 ( .A1(n16318), .A2(n16319), .ZN(n16317) );
  INV_X1 U11793 ( .A(n19387), .ZN(n19366) );
  NOR2_X1 U11794 ( .A1(n15241), .A2(n12897), .ZN(n12901) );
  NAND2_X1 U11795 ( .A1(n12575), .A2(n10160), .ZN(n19405) );
  NOR2_X1 U11796 ( .A1(n10163), .A2(n10161), .ZN(n10160) );
  INV_X1 U11797 ( .A(n13636), .ZN(n10161) );
  NAND2_X1 U11798 ( .A1(n12864), .A2(n12863), .ZN(n19428) );
  NAND2_X1 U11799 ( .A1(n12862), .A2(n13350), .ZN(n12864) );
  AND2_X1 U11800 ( .A1(n19428), .A2(n19584), .ZN(n19417) );
  XNOR2_X1 U11801 ( .A(n9958), .B(n10192), .ZN(n12904) );
  NAND2_X1 U11802 ( .A1(n10219), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9958) );
  NAND2_X1 U11803 ( .A1(n10095), .A2(n10093), .ZN(n10092) );
  INV_X1 U11804 ( .A(n10094), .ZN(n10093) );
  OR2_X1 U11805 ( .A1(n12325), .A2(n19501), .ZN(n10095) );
  OAI21_X1 U11806 ( .B1(n16506), .B2(n10638), .A(n12324), .ZN(n10094) );
  AND2_X1 U11807 ( .A1(n12319), .A2(n12030), .ZN(n19507) );
  NOR2_X1 U11808 ( .A1(n14509), .A2(n9758), .ZN(n14510) );
  XNOR2_X1 U11809 ( .A(n12263), .B(n10172), .ZN(n12539) );
  INV_X1 U11810 ( .A(n20166), .ZN(n20169) );
  NOR2_X1 U11811 ( .A1(n11955), .A2(n12553), .ZN(n9857) );
  INV_X1 U11812 ( .A(n17136), .ZN(n17194) );
  INV_X1 U11813 ( .A(n17568), .ZN(n17564) );
  NOR2_X1 U11814 ( .A1(n17578), .A2(n9870), .ZN(n9869) );
  NOR3_X1 U11815 ( .A1(n17612), .A2(n17579), .A3(n17536), .ZN(n17574) );
  NAND2_X1 U11816 ( .A1(n17616), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17612) );
  NOR2_X2 U11817 ( .A1(n18525), .A2(n17680), .ZN(n17610) );
  NOR2_X1 U11818 ( .A1(n17623), .A2(n17793), .ZN(n17616) );
  AND2_X1 U11819 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17658), .ZN(n17646) );
  INV_X1 U11820 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18400) );
  INV_X1 U11821 ( .A(n17173), .ZN(n19028) );
  NAND2_X1 U11822 ( .A1(n10622), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n9841) );
  INV_X1 U11823 ( .A(n11964), .ZN(n12074) );
  NAND2_X1 U11824 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n9855) );
  INV_X1 U11825 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10260) );
  OR2_X1 U11826 ( .A1(n12733), .A2(n10259), .ZN(n10263) );
  OAI21_X1 U11827 ( .B1(n17470), .B2(n18933), .A(n9876), .ZN(n9875) );
  NAND2_X1 U11828 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n9876) );
  INV_X1 U11829 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n9903) );
  INV_X1 U11830 ( .A(n11741), .ZN(n11737) );
  NOR2_X1 U11831 ( .A1(n11251), .A2(n10123), .ZN(n10122) );
  INV_X1 U11832 ( .A(n11238), .ZN(n10123) );
  OR2_X1 U11833 ( .A1(n11272), .A2(n11271), .ZN(n12392) );
  INV_X1 U11834 ( .A(n11280), .ZN(n9891) );
  INV_X1 U11835 ( .A(n11281), .ZN(n9892) );
  OR2_X1 U11836 ( .A1(n11225), .A2(n11224), .ZN(n12365) );
  AND2_X1 U11837 ( .A1(n13802), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11087) );
  INV_X1 U11838 ( .A(n11090), .ZN(n12401) );
  NOR2_X1 U11839 ( .A1(n11151), .A2(n11150), .ZN(n12331) );
  NOR2_X1 U11840 ( .A1(n10900), .A2(n20222), .ZN(n10042) );
  NAND2_X1 U11841 ( .A1(n10119), .A2(n11035), .ZN(n13499) );
  INV_X1 U11842 ( .A(n11001), .ZN(n10998) );
  NAND2_X1 U11843 ( .A1(n13989), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11190) );
  AOI21_X1 U11844 ( .B1(n11736), .B2(n11735), .A(n11732), .ZN(n11766) );
  NAND2_X1 U11845 ( .A1(n11050), .A2(n11035), .ZN(n11006) );
  NAND2_X1 U11846 ( .A1(n13378), .A2(n11036), .ZN(n11005) );
  INV_X1 U11847 ( .A(n11762), .ZN(n11768) );
  NOR2_X1 U11848 ( .A1(n10118), .A2(n12178), .ZN(n10117) );
  INV_X1 U11849 ( .A(n10877), .ZN(n10118) );
  INV_X1 U11850 ( .A(n12235), .ZN(n10076) );
  AOI22_X1 U11851 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10232) );
  AOI22_X1 U11852 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10328) );
  INV_X1 U11853 ( .A(n15417), .ZN(n10083) );
  NOR2_X1 U11854 ( .A1(n16551), .A2(n15749), .ZN(n10145) );
  NAND2_X1 U11855 ( .A1(n12035), .A2(n12034), .ZN(n12142) );
  OR3_X1 U11856 ( .A1(n10365), .A2(n10080), .A3(n10368), .ZN(n10851) );
  INV_X1 U11857 ( .A(n10366), .ZN(n10368) );
  NOR2_X1 U11858 ( .A1(n12865), .A2(n9687), .ZN(n10709) );
  NAND2_X1 U11859 ( .A1(n10253), .A2(n10252), .ZN(n10257) );
  OR2_X1 U11860 ( .A1(n12733), .A2(n11967), .ZN(n10255) );
  AND2_X1 U11861 ( .A1(n19513), .A2(n11963), .ZN(n11990) );
  OAI21_X1 U11862 ( .B1(n9838), .B2(n9837), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9839) );
  OAI21_X1 U11863 ( .B1(n9836), .B2(n9835), .A(n10282), .ZN(n9844) );
  NOR2_X1 U11864 ( .A1(n17667), .A2(n13201), .ZN(n13189) );
  NAND2_X1 U11865 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18487), .ZN(
        n13182) );
  AOI21_X1 U11866 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n19005), .A(
        n13073), .ZN(n13184) );
  AND2_X1 U11867 ( .A1(n9906), .A2(n9905), .ZN(n13079) );
  NAND2_X1 U11868 ( .A1(n9730), .A2(n9902), .ZN(n9905) );
  NAND2_X1 U11869 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n9906) );
  NOR2_X1 U11870 ( .A1(n12924), .A2(n9903), .ZN(n9902) );
  INV_X1 U11871 ( .A(n14563), .ZN(n10129) );
  INV_X1 U11872 ( .A(n10131), .ZN(n10130) );
  NAND2_X1 U11873 ( .A1(n9743), .A2(n11466), .ZN(n10133) );
  NOR2_X1 U11874 ( .A1(n12429), .A2(n10062), .ZN(n10061) );
  NAND2_X1 U11875 ( .A1(n11879), .A2(n9985), .ZN(n9984) );
  NAND2_X1 U11876 ( .A1(n10046), .A2(n10045), .ZN(n14846) );
  AOI21_X1 U11877 ( .B1(n15065), .B2(n14943), .A(n14942), .ZN(n10045) );
  AND2_X1 U11878 ( .A1(n14905), .A2(n12416), .ZN(n16127) );
  INV_X1 U11879 ( .A(n14693), .ZN(n9989) );
  NOR2_X1 U11880 ( .A1(n9810), .A2(n9728), .ZN(n9982) );
  NOR2_X1 U11881 ( .A1(n13792), .A2(n9830), .ZN(n9973) );
  OR2_X1 U11882 ( .A1(n11201), .A2(n11200), .ZN(n12361) );
  INV_X1 U11883 ( .A(n14961), .ZN(n13629) );
  NAND2_X1 U11884 ( .A1(n11087), .A2(n11033), .ZN(n11762) );
  INV_X1 U11885 ( .A(n12340), .ZN(n11118) );
  NOR2_X1 U11886 ( .A1(n11762), .A2(n12400), .ZN(n11764) );
  INV_X1 U11887 ( .A(n13589), .ZN(n13522) );
  NOR2_X1 U11888 ( .A1(n10116), .A2(n12177), .ZN(n10115) );
  INV_X1 U11889 ( .A(n10117), .ZN(n10116) );
  INV_X1 U11890 ( .A(n12098), .ZN(n10098) );
  INV_X1 U11891 ( .A(n13340), .ZN(n13267) );
  OR2_X1 U11892 ( .A1(n12754), .A2(n12755), .ZN(n12756) );
  AOI21_X1 U11893 ( .B1(n10699), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10700), 
        .ZN(n10701) );
  AND2_X1 U11894 ( .A1(n16631), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10700) );
  NOR2_X1 U11895 ( .A1(n9799), .A2(n10156), .ZN(n10155) );
  NOR2_X1 U11896 ( .A1(n16425), .A2(n9967), .ZN(n9966) );
  NOR2_X1 U11897 ( .A1(n19230), .A2(n9970), .ZN(n9969) );
  INV_X1 U11898 ( .A(n15522), .ZN(n10114) );
  NAND2_X1 U11899 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n10212), .ZN(
        n10211) );
  NOR2_X1 U11900 ( .A1(n16457), .A2(n9964), .ZN(n9963) );
  INV_X1 U11901 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n9964) );
  NOR2_X1 U11902 ( .A1(n15436), .A2(n15619), .ZN(n10148) );
  NAND2_X1 U11903 ( .A1(n15454), .A2(n16464), .ZN(n9947) );
  NAND2_X1 U11904 ( .A1(n9946), .A2(n9948), .ZN(n9945) );
  INV_X1 U11905 ( .A(n15454), .ZN(n9948) );
  NAND2_X1 U11906 ( .A1(n15454), .A2(n16450), .ZN(n10035) );
  NAND2_X1 U11907 ( .A1(n10103), .A2(n10780), .ZN(n10102) );
  INV_X1 U11908 ( .A(n13242), .ZN(n10103) );
  NOR2_X1 U11909 ( .A1(n15708), .A2(n16535), .ZN(n15709) );
  NOR2_X1 U11910 ( .A1(n15744), .A2(n10028), .ZN(n10027) );
  INV_X1 U11911 ( .A(n15727), .ZN(n10028) );
  NAND2_X1 U11912 ( .A1(n16496), .A2(n16495), .ZN(n12146) );
  INV_X1 U11913 ( .A(n10087), .ZN(n10090) );
  INV_X1 U11914 ( .A(n10851), .ZN(n12289) );
  OR2_X1 U11915 ( .A1(n12282), .A2(n9720), .ZN(n10860) );
  AOI21_X1 U11916 ( .B1(n10707), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10706), 
        .ZN(n10708) );
  NOR2_X1 U11917 ( .A1(n10632), .A2(n10655), .ZN(n10659) );
  AOI22_X1 U11918 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10616) );
  AND2_X1 U11919 ( .A1(n19513), .A2(n11957), .ZN(n11978) );
  NAND3_X1 U11920 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20157), .A3(n19995), 
        .ZN(n13752) );
  NAND2_X1 U11921 ( .A1(n10598), .A2(n10597), .ZN(n10641) );
  NAND4_X1 U11922 ( .A1(n10174), .A2(n10596), .A3(n10595), .A4(n10594), .ZN(
        n10597) );
  AOI22_X1 U11923 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10596) );
  AOI22_X1 U11924 ( .A1(n9712), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n10621), .ZN(n10606) );
  AOI22_X1 U11925 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10607) );
  NOR3_X1 U11926 ( .A1(n13121), .A2(n9877), .A3(n9872), .ZN(n13122) );
  NOR2_X1 U11927 ( .A1(n12951), .A2(n9878), .ZN(n9877) );
  NAND3_X1 U11928 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n19146), .ZN(n12922) );
  INV_X1 U11929 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17471) );
  NAND2_X1 U11930 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12960) );
  OR2_X1 U11931 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15945), .ZN(
        n17486) );
  NAND2_X1 U11932 ( .A1(n16814), .A2(n13162), .ZN(n15934) );
  INV_X1 U11933 ( .A(n17947), .ZN(n9916) );
  AND2_X1 U11934 ( .A1(n17984), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9919) );
  INV_X1 U11935 ( .A(n16842), .ZN(n9918) );
  INV_X1 U11936 ( .A(n18047), .ZN(n9917) );
  AND2_X1 U11937 ( .A1(n18363), .A2(n18021), .ZN(n10074) );
  AND2_X1 U11938 ( .A1(n13016), .A2(n17682), .ZN(n13035) );
  OAI211_X1 U11939 ( .C1(n13141), .C2(n18528), .A(n13158), .B(n13157), .ZN(
        n13174) );
  INV_X1 U11940 ( .A(n13023), .ZN(n12919) );
  AOI221_X1 U11941 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19134), .C1(n19183), 
        .C2(P3_STATE2_REG_1__SCAN_IN), .A(n19147), .ZN(n18490) );
  INV_X1 U11942 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16075) );
  INV_X1 U11943 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16099) );
  AOI21_X1 U11944 ( .B1(n13563), .B2(n9684), .A(n11794), .ZN(n13616) );
  AND2_X1 U11945 ( .A1(n14817), .A2(n13980), .ZN(n11670) );
  AND2_X1 U11946 ( .A1(n11647), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11648) );
  AND2_X1 U11947 ( .A1(n11605), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11606) );
  OR2_X1 U11948 ( .A1(n14851), .A2(n11177), .ZN(n11609) );
  AND2_X1 U11949 ( .A1(n14862), .A2(n13980), .ZN(n11585) );
  NOR2_X1 U11950 ( .A1(n11564), .A2(n14873), .ZN(n11565) );
  AND2_X1 U11951 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n11517), .ZN(
        n11518) );
  AND2_X1 U11952 ( .A1(n11484), .A2(n11483), .ZN(n14722) );
  NOR2_X1 U11953 ( .A1(n11452), .A2(n16075), .ZN(n11481) );
  CLKBUF_X1 U11954 ( .A(n14676), .Z(n14677) );
  NOR2_X1 U11955 ( .A1(n11405), .A2(n11358), .ZN(n11423) );
  NAND2_X1 U11956 ( .A1(n11374), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11405) );
  CLKBUF_X1 U11957 ( .A(n14437), .Z(n14438) );
  AND2_X1 U11958 ( .A1(n11337), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11338) );
  NAND2_X1 U11959 ( .A1(n14153), .A2(n9825), .ZN(n14375) );
  NAND2_X1 U11960 ( .A1(n11308), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11333) );
  AND2_X1 U11961 ( .A1(n11285), .A2(n11284), .ZN(n11308) );
  AND2_X1 U11962 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11284) );
  AND2_X1 U11963 ( .A1(n11254), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11285) );
  NOR2_X1 U11964 ( .A1(n11208), .A2(n11207), .ZN(n11231) );
  CLKBUF_X1 U11965 ( .A(n13642), .Z(n13643) );
  INV_X1 U11966 ( .A(n13696), .ZN(n11180) );
  AND2_X1 U11967 ( .A1(n14586), .A2(n14574), .ZN(n14576) );
  OR2_X1 U11968 ( .A1(n9754), .A2(n14603), .ZN(n14605) );
  AND2_X1 U11969 ( .A1(n11891), .A2(n11890), .ZN(n14587) );
  NOR2_X1 U11970 ( .A1(n9752), .A2(n9983), .ZN(n14654) );
  INV_X1 U11971 ( .A(n9985), .ZN(n9983) );
  AND2_X1 U11972 ( .A1(n11870), .A2(n11869), .ZN(n14713) );
  NOR2_X1 U11973 ( .A1(n9752), .A2(n14713), .ZN(n14714) );
  NOR2_X1 U11974 ( .A1(n14736), .A2(n14679), .ZN(n14725) );
  AND2_X1 U11975 ( .A1(n11858), .A2(n11857), .ZN(n14733) );
  NAND2_X1 U11976 ( .A1(n14465), .A2(n9987), .ZN(n14736) );
  AND2_X1 U11977 ( .A1(n9803), .A2(n9988), .ZN(n9987) );
  INV_X1 U11978 ( .A(n14733), .ZN(n9988) );
  NAND2_X1 U11979 ( .A1(n14465), .A2(n9803), .ZN(n14734) );
  NAND2_X1 U11980 ( .A1(n14465), .A2(n14464), .ZN(n14692) );
  NOR2_X1 U11981 ( .A1(n14459), .A2(n14441), .ZN(n14465) );
  AND2_X1 U11982 ( .A1(n11848), .A2(n11847), .ZN(n14457) );
  NAND2_X1 U11983 ( .A1(n9981), .A2(n9979), .ZN(n14459) );
  AND2_X1 U11984 ( .A1(n9982), .A2(n9980), .ZN(n9979) );
  INV_X1 U11985 ( .A(n14457), .ZN(n9980) );
  NAND2_X1 U11986 ( .A1(n9981), .A2(n9982), .ZN(n15091) );
  NOR2_X1 U11987 ( .A1(n14338), .A2(n9728), .ZN(n16105) );
  NAND2_X1 U11988 ( .A1(n14391), .A2(n12409), .ZN(n10054) );
  NAND2_X1 U11989 ( .A1(n10053), .A2(n10058), .ZN(n10052) );
  INV_X1 U11990 ( .A(n14391), .ZN(n10053) );
  AND2_X1 U11991 ( .A1(n11833), .A2(n11832), .ZN(n14339) );
  NOR2_X1 U11992 ( .A1(n14338), .A2(n14339), .ZN(n14380) );
  INV_X1 U11993 ( .A(n9897), .ZN(n14389) );
  INV_X1 U11994 ( .A(n10049), .ZN(n10048) );
  OR2_X1 U11995 ( .A1(n13647), .A2(n9976), .ZN(n14279) );
  NAND2_X1 U11996 ( .A1(n9974), .A2(n9972), .ZN(n9976) );
  INV_X1 U11997 ( .A(n13648), .ZN(n9974) );
  AND2_X1 U11998 ( .A1(n14108), .A2(n9973), .ZN(n9972) );
  NOR2_X1 U11999 ( .A1(n13647), .A2(n9975), .ZN(n16282) );
  NAND2_X1 U12000 ( .A1(n9978), .A2(n14108), .ZN(n9975) );
  NOR2_X1 U12001 ( .A1(n13647), .A2(n9977), .ZN(n14109) );
  INV_X1 U12002 ( .A(n9978), .ZN(n9977) );
  OR2_X1 U12003 ( .A1(n13647), .A2(n13648), .ZN(n13791) );
  AND2_X1 U12004 ( .A1(n13602), .A2(n13601), .ZN(n13623) );
  INV_X1 U12005 ( .A(n11084), .ZN(n11085) );
  NAND2_X1 U12006 ( .A1(n11172), .A2(n20222), .ZN(n11086) );
  INV_X1 U12007 ( .A(n11340), .ZN(n13843) );
  AND2_X1 U12008 ( .A1(n20706), .A2(n14311), .ZN(n20619) );
  INV_X1 U12009 ( .A(n13827), .ZN(n13874) );
  INV_X1 U12010 ( .A(n20703), .ZN(n20516) );
  AND2_X1 U12011 ( .A1(n9716), .A2(n14198), .ZN(n20670) );
  AND2_X1 U12012 ( .A1(n9716), .A2(n9669), .ZN(n20610) );
  OR2_X1 U12013 ( .A1(n14077), .A2(n14076), .ZN(n15996) );
  AND2_X1 U12014 ( .A1(n10866), .A2(n10861), .ZN(n12458) );
  OR2_X1 U12015 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n12238), .ZN(n12242) );
  NAND2_X1 U12016 ( .A1(n12890), .A2(n12241), .ZN(n12250) );
  NAND2_X1 U12017 ( .A1(n12235), .A2(n12242), .ZN(n12890) );
  NAND2_X1 U12018 ( .A1(n12194), .A2(n12219), .ZN(n12227) );
  NAND2_X1 U12019 ( .A1(n12097), .A2(n9764), .ZN(n12152) );
  INV_X1 U12020 ( .A(n12128), .ZN(n10872) );
  NAND2_X1 U12021 ( .A1(n10857), .A2(n10856), .ZN(n12106) );
  XNOR2_X1 U12022 ( .A(n12778), .B(n9824), .ZN(n9849) );
  NAND2_X1 U12023 ( .A1(n13691), .A2(n10164), .ZN(n10163) );
  AND2_X1 U12024 ( .A1(n9746), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10164) );
  NOR2_X1 U12025 ( .A1(n9767), .A2(n10150), .ZN(n10149) );
  INV_X1 U12026 ( .A(n12571), .ZN(n10150) );
  AND2_X1 U12027 ( .A1(n9720), .A2(n13415), .ZN(n12866) );
  INV_X1 U12028 ( .A(n12463), .ZN(n13393) );
  INV_X1 U12029 ( .A(n15293), .ZN(n13751) );
  NAND2_X1 U12030 ( .A1(n10194), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10218) );
  AND2_X1 U12031 ( .A1(n10196), .A2(n9965), .ZN(n10194) );
  AND2_X1 U12032 ( .A1(n9747), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9965) );
  NAND2_X1 U12033 ( .A1(n10196), .A2(n9747), .ZN(n10217) );
  NAND2_X1 U12034 ( .A1(n10196), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10216) );
  NOR2_X1 U12035 ( .A1(n15437), .A2(n10197), .ZN(n10196) );
  AND2_X1 U12036 ( .A1(n10214), .A2(n9968), .ZN(n10198) );
  AND2_X1 U12037 ( .A1(n9742), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9968) );
  NAND2_X1 U12038 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n10198), .ZN(
        n10197) );
  NAND2_X1 U12039 ( .A1(n10214), .A2(n9742), .ZN(n10215) );
  NOR2_X1 U12040 ( .A1(n10211), .A2(n15516), .ZN(n10214) );
  NAND2_X1 U12041 ( .A1(n10214), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10213) );
  AND2_X1 U12042 ( .A1(n14294), .A2(n10112), .ZN(n15505) );
  NAND2_X1 U12043 ( .A1(n14294), .A2(n9802), .ZN(n15524) );
  AND2_X1 U12044 ( .A1(n10209), .A2(n9962), .ZN(n10212) );
  AND2_X1 U12045 ( .A1(n9741), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9962) );
  NAND2_X1 U12046 ( .A1(n10209), .A2(n9741), .ZN(n10210) );
  NAND2_X1 U12047 ( .A1(n10209), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10208) );
  NOR2_X1 U12048 ( .A1(n16473), .A2(n10206), .ZN(n10209) );
  NOR2_X1 U12049 ( .A1(n15733), .A2(n10102), .ZN(n14010) );
  NAND2_X1 U12050 ( .A1(n10101), .A2(n10780), .ZN(n15735) );
  INV_X1 U12051 ( .A(n15733), .ZN(n10101) );
  NAND2_X1 U12052 ( .A1(n9959), .A2(n9811), .ZN(n10204) );
  AOI21_X2 U12053 ( .B1(n14342), .B2(n10140), .A(n10139), .ZN(n15535) );
  AND2_X1 U12054 ( .A1(n15764), .A2(n15763), .ZN(n10139) );
  AND2_X1 U12055 ( .A1(n12313), .A2(n12314), .ZN(n15534) );
  NAND2_X1 U12056 ( .A1(n9959), .A2(n9960), .ZN(n10202) );
  AND2_X1 U12057 ( .A1(n9959), .A2(n9739), .ZN(n10205) );
  NOR2_X1 U12058 ( .A1(n10200), .A2(n16507), .ZN(n10203) );
  INV_X1 U12059 ( .A(n19368), .ZN(n10755) );
  NAND2_X1 U12060 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10199) );
  NOR2_X1 U12061 ( .A1(n10199), .A2(n14035), .ZN(n10201) );
  INV_X1 U12062 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14035) );
  NAND2_X1 U12063 ( .A1(n15277), .A2(n10104), .ZN(n15241) );
  AND2_X1 U12064 ( .A1(n10106), .A2(n15266), .ZN(n10104) );
  NOR2_X1 U12065 ( .A1(n10107), .A2(n10109), .ZN(n10106) );
  INV_X1 U12066 ( .A(n15239), .ZN(n10109) );
  INV_X1 U12067 ( .A(n10107), .ZN(n10105) );
  NAND2_X1 U12068 ( .A1(n15259), .A2(n15260), .ZN(n15262) );
  INV_X1 U12069 ( .A(n15419), .ZN(n15392) );
  AND2_X1 U12070 ( .A1(n9751), .A2(n9834), .ZN(n10147) );
  NAND2_X1 U12071 ( .A1(n9938), .A2(n9937), .ZN(n15599) );
  INV_X1 U12072 ( .A(n15143), .ZN(n10078) );
  NAND2_X1 U12073 ( .A1(n15443), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15444) );
  AND2_X1 U12074 ( .A1(n10550), .A2(n10549), .ZN(n15176) );
  INV_X1 U12075 ( .A(n10037), .ZN(n10036) );
  OAI21_X1 U12076 ( .B1(n9724), .B2(n15463), .A(n15464), .ZN(n10037) );
  AND2_X1 U12077 ( .A1(n10546), .A2(n10545), .ZN(n14425) );
  NAND2_X1 U12078 ( .A1(n15510), .A2(n15463), .ZN(n15503) );
  INV_X1 U12079 ( .A(n14302), .ZN(n10001) );
  NOR2_X1 U12080 ( .A1(n15671), .A2(n16432), .ZN(n9956) );
  OR2_X1 U12081 ( .A1(n16532), .A2(n9999), .ZN(n15692) );
  NOR2_X1 U12082 ( .A1(n16532), .A2(n16533), .ZN(n16531) );
  INV_X1 U12083 ( .A(n15744), .ZN(n10026) );
  CLKBUF_X1 U12084 ( .A(n13433), .Z(n16559) );
  AND2_X1 U12085 ( .A1(n10439), .A2(n10438), .ZN(n13438) );
  NAND2_X1 U12086 ( .A1(n14051), .A2(n10435), .ZN(n13441) );
  NAND2_X1 U12087 ( .A1(n9950), .A2(n9949), .ZN(n16498) );
  AND2_X1 U12088 ( .A1(n11946), .A2(n11942), .ZN(n11950) );
  INV_X1 U12089 ( .A(n12035), .ZN(n12294) );
  NAND2_X1 U12090 ( .A1(n13579), .A2(n13578), .ZN(n13577) );
  NAND2_X1 U12091 ( .A1(n12542), .A2(n19920), .ZN(n12566) );
  INV_X1 U12092 ( .A(n13243), .ZN(n19372) );
  CLKBUF_X1 U12093 ( .A(n10699), .Z(n15803) );
  NOR2_X1 U12094 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15790) );
  NOR2_X1 U12095 ( .A1(n15796), .A2(n20169), .ZN(n19596) );
  AND2_X1 U12096 ( .A1(n9721), .A2(n13416), .ZN(n10138) );
  INV_X1 U12097 ( .A(n12039), .ZN(n13962) );
  INV_X1 U12098 ( .A(n19695), .ZN(n19753) );
  NOR2_X2 U12099 ( .A1(n13751), .A2(n13752), .ZN(n19587) );
  NAND2_X1 U12100 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19995), .ZN(n19583) );
  INV_X1 U12101 ( .A(n19760), .ZN(n20151) );
  NAND2_X1 U12102 ( .A1(n13349), .A2(n13348), .ZN(n16620) );
  INV_X1 U12103 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20065) );
  NOR2_X1 U12104 ( .A1(n18978), .A2(n13251), .ZN(n18954) );
  NOR2_X1 U12105 ( .A1(n16863), .A2(n16862), .ZN(n16861) );
  NOR2_X1 U12106 ( .A1(n16876), .A2(n16875), .ZN(n16874) );
  NOR2_X1 U12107 ( .A1(n17876), .A2(n16935), .ZN(n16934) );
  NOR2_X1 U12108 ( .A1(n17888), .A2(n16944), .ZN(n16943) );
  NOR2_X1 U12109 ( .A1(n17182), .A2(n16843), .ZN(n16957) );
  NOR2_X1 U12110 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17116), .ZN(n17088) );
  AND2_X1 U12111 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17311), .ZN(n17285) );
  NAND2_X1 U12112 ( .A1(n9881), .A2(n9879), .ZN(n17538) );
  NOR2_X1 U12113 ( .A1(n13126), .A2(n9880), .ZN(n9879) );
  INV_X1 U12114 ( .A(n13125), .ZN(n9881) );
  AND2_X1 U12115 ( .A1(n15828), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n9880) );
  INV_X1 U12116 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17464) );
  OAI211_X1 U12117 ( .C1(n17470), .C2(n18523), .A(n13002), .B(n13001), .ZN(
        n13188) );
  NAND2_X1 U12118 ( .A1(n17431), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12939) );
  NOR2_X1 U12119 ( .A1(n10066), .A2(n10065), .ZN(n10064) );
  NAND2_X1 U12120 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12973) );
  OR2_X1 U12121 ( .A1(n9756), .A2(n17344), .ZN(n10168) );
  INV_X1 U12122 ( .A(n17726), .ZN(n17690) );
  INV_X1 U12123 ( .A(n17727), .ZN(n17728) );
  NAND2_X1 U12124 ( .A1(n16660), .A2(n9925), .ZN(n9930) );
  NOR2_X1 U12125 ( .A1(n9926), .A2(n9931), .ZN(n9925) );
  INV_X1 U12126 ( .A(n9927), .ZN(n9926) );
  NOR2_X1 U12127 ( .A1(n13220), .A2(n17797), .ZN(n16660) );
  AND2_X1 U12128 ( .A1(n17900), .A2(n9818), .ZN(n17825) );
  INV_X1 U12129 ( .A(n17837), .ZN(n9920) );
  NOR2_X1 U12130 ( .A1(n17878), .A2(n9922), .ZN(n9921) );
  INV_X1 U12131 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9922) );
  NAND2_X1 U12132 ( .A1(n17900), .A2(n9732), .ZN(n17836) );
  NAND2_X1 U12133 ( .A1(n17900), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17877) );
  NOR2_X1 U12134 ( .A1(n17912), .A2(n17913), .ZN(n17900) );
  NOR2_X1 U12135 ( .A1(n18047), .A2(n16842), .ZN(n17985) );
  AND2_X1 U12136 ( .A1(n18086), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18011) );
  AND2_X1 U12137 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18106) );
  NOR2_X1 U12138 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19183), .ZN(n17987) );
  AOI21_X1 U12139 ( .B1(n13059), .B2(n17968), .A(n10069), .ZN(n16015) );
  NOR2_X1 U12140 ( .A1(n16015), .A2(n16655), .ZN(n16014) );
  NAND2_X1 U12141 ( .A1(n17812), .A2(n18057), .ZN(n16688) );
  INV_X1 U12142 ( .A(n18165), .ZN(n17802) );
  NAND2_X1 U12143 ( .A1(n10013), .A2(n10012), .ZN(n10016) );
  NAND2_X1 U12144 ( .A1(n18057), .A2(n10017), .ZN(n10012) );
  NAND2_X1 U12145 ( .A1(n17897), .A2(n10014), .ZN(n10013) );
  AND2_X1 U12146 ( .A1(n9829), .A2(n17997), .ZN(n10073) );
  AND2_X1 U12147 ( .A1(n18022), .A2(n10074), .ZN(n17996) );
  AND2_X1 U12148 ( .A1(n18311), .A2(n18417), .ZN(n18321) );
  NOR2_X1 U12149 ( .A1(n18076), .A2(n18399), .ZN(n18075) );
  INV_X1 U12150 ( .A(n18127), .ZN(n10005) );
  INV_X1 U12151 ( .A(n18976), .ZN(n18979) );
  NOR2_X2 U12152 ( .A1(n19185), .A2(n15943), .ZN(n18964) );
  NOR2_X1 U12153 ( .A1(n12924), .A2(n18977), .ZN(n18970) );
  INV_X1 U12154 ( .A(n13250), .ZN(n9865) );
  AOI211_X1 U12155 ( .C1(n17488), .C2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n13148), .B(n13147), .ZN(n18514) );
  NOR2_X1 U12156 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18490), .ZN(n18857) );
  INV_X1 U12157 ( .A(n17538), .ZN(n18520) );
  INV_X1 U12158 ( .A(n18717), .ZN(n18891) );
  AOI21_X1 U12159 ( .B1(n18953), .B2(n18957), .A(n9793), .ZN(n18962) );
  OAI211_X1 U12160 ( .C1(n19170), .C2(n19171), .A(n19165), .B(n16812), .ZN(
        n19013) );
  AND2_X1 U12161 ( .A1(n16082), .A2(n14002), .ZN(n20307) );
  AND2_X1 U12162 ( .A1(n16082), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20306) );
  INV_X1 U12163 ( .A(n20259), .ZN(n20309) );
  INV_X1 U12164 ( .A(n16082), .ZN(n20301) );
  AND2_X1 U12165 ( .A1(n14000), .A2(n13994), .ZN(n20303) );
  NAND2_X1 U12166 ( .A1(n14000), .A2(n13998), .ZN(n20259) );
  AND2_X1 U12167 ( .A1(n14000), .A2(n13999), .ZN(n20304) );
  XNOR2_X1 U12168 ( .A(n9991), .B(n14524), .ZN(n14934) );
  INV_X1 U12169 ( .A(n14737), .ZN(n20320) );
  NAND2_X2 U12170 ( .A1(n11782), .A2(n11781), .ZN(n20324) );
  NAND2_X1 U12171 ( .A1(n20324), .A2(n14537), .ZN(n14737) );
  INV_X1 U12172 ( .A(n14767), .ZN(n14799) );
  NOR2_X1 U12173 ( .A1(n14783), .A2(n13702), .ZN(n14477) );
  NAND2_X1 U12174 ( .A1(n11921), .A2(n11920), .ZN(n14743) );
  NAND2_X1 U12175 ( .A1(n13529), .A2(n13601), .ZN(n11921) );
  INV_X1 U12176 ( .A(n14477), .ZN(n14490) );
  AND2_X1 U12177 ( .A1(n13540), .A2(n13539), .ZN(n20328) );
  INV_X1 U12178 ( .A(n13650), .ZN(n20369) );
  NOR2_X2 U12179 ( .A1(n20368), .A2(n13596), .ZN(n13681) );
  AND2_X1 U12180 ( .A1(n12439), .A2(n11692), .ZN(n14809) );
  INV_X1 U12181 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14873) );
  OAI21_X1 U12182 ( .B1(n14879), .B2(n14943), .A(n15065), .ZN(n14871) );
  AND2_X1 U12183 ( .A1(n14712), .A2(n14711), .ZN(n16059) );
  NAND2_X1 U12184 ( .A1(n10135), .A2(n9821), .ZN(n14731) );
  INV_X1 U12185 ( .A(n14887), .ZN(n16120) );
  OR2_X1 U12186 ( .A1(n16183), .A2(n12437), .ZN(n16187) );
  AND2_X1 U12187 ( .A1(n16187), .A2(n13491), .ZN(n16181) );
  INV_X1 U12188 ( .A(n16187), .ZN(n16173) );
  NAND2_X1 U12189 ( .A1(n9895), .A2(n9896), .ZN(n12914) );
  NAND2_X1 U12190 ( .A1(n12428), .A2(n14984), .ZN(n14806) );
  NOR2_X1 U12191 ( .A1(n12428), .A2(n12427), .ZN(n14807) );
  OR2_X1 U12192 ( .A1(n12441), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16238) );
  INV_X1 U12193 ( .A(n16286), .ZN(n16239) );
  NAND2_X1 U12194 ( .A1(n10051), .A2(n12379), .ZN(n16177) );
  NAND2_X1 U12195 ( .A1(n14224), .A2(n14225), .ZN(n10051) );
  INV_X1 U12196 ( .A(n16222), .ZN(n16289) );
  INV_X1 U12197 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n14105) );
  INV_X1 U12198 ( .A(n20696), .ZN(n20743) );
  CLKBUF_X1 U12199 ( .A(n13495), .Z(n13496) );
  NAND2_X1 U12200 ( .A1(n9763), .A2(n11206), .ZN(n15112) );
  NOR2_X1 U12201 ( .A1(n15112), .A2(n14097), .ZN(n20671) );
  NOR2_X1 U12202 ( .A1(n9692), .A2(n9899), .ZN(n15118) );
  NOR2_X1 U12203 ( .A1(n20888), .A2(n9899), .ZN(n15121) );
  NAND2_X1 U12204 ( .A1(n20700), .A2(n13985), .ZN(n20897) );
  OAI211_X1 U12205 ( .C1(n20696), .C2(n13891), .A(n13889), .B(n20748), .ZN(
        n20410) );
  OAI22_X1 U12206 ( .A1(n20520), .A2(n20519), .B1(n20706), .B2(n20518), .ZN(
        n20538) );
  INV_X1 U12207 ( .A(n20599), .ZN(n20576) );
  INV_X1 U12208 ( .A(n20548), .ZN(n20568) );
  OAI22_X1 U12209 ( .A1(n20624), .A2(n20623), .B1(n20622), .B2(n20621), .ZN(
        n20657) );
  NAND2_X1 U12210 ( .A1(n20671), .A2(n20670), .ZN(n20737) );
  INV_X1 U12211 ( .A(n20704), .ZN(n20734) );
  INV_X1 U12212 ( .A(n20611), .ZN(n20745) );
  INV_X1 U12213 ( .A(n20627), .ZN(n20756) );
  INV_X1 U12214 ( .A(n20631), .ZN(n20762) );
  INV_X1 U12215 ( .A(n20636), .ZN(n20768) );
  INV_X1 U12216 ( .A(n20640), .ZN(n20774) );
  INV_X1 U12217 ( .A(n20644), .ZN(n20780) );
  NAND2_X1 U12218 ( .A1(n20747), .A2(n20670), .ZN(n20791) );
  INV_X1 U12219 ( .A(n20649), .ZN(n20786) );
  AND2_X1 U12220 ( .A1(n20747), .A2(n20610), .ZN(n20788) );
  INV_X1 U12221 ( .A(n20791), .ZN(n20798) );
  OAI21_X1 U12222 ( .B1(n20750), .B2(n20749), .A(n20748), .ZN(n20799) );
  AND2_X1 U12223 ( .A1(n16004), .A2(n16003), .ZN(n16299) );
  INV_X1 U12224 ( .A(n16008), .ZN(n20804) );
  INV_X1 U12225 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20222) );
  INV_X1 U12226 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20700) );
  AND2_X1 U12227 ( .A1(n10575), .A2(n10574), .ZN(n20184) );
  AND2_X1 U12228 ( .A1(n16616), .A2(n20205), .ZN(n20189) );
  NAND2_X1 U12229 ( .A1(n16353), .A2(n16354), .ZN(n16352) );
  AND2_X1 U12230 ( .A1(n12236), .A2(n12235), .ZN(n16359) );
  NAND2_X1 U12231 ( .A1(n16362), .A2(n16363), .ZN(n16361) );
  OR2_X1 U12232 ( .A1(n13389), .A2(n16629), .ZN(n19381) );
  AOI22_X1 U12233 ( .A1(n12904), .A2(n20201), .B1(n10193), .B2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n13243) );
  INV_X1 U12234 ( .A(n19391), .ZN(n19360) );
  AND2_X1 U12235 ( .A1(n13275), .A2(n10891), .ZN(n19361) );
  INV_X1 U12236 ( .A(n19361), .ZN(n19382) );
  INV_X1 U12237 ( .A(n19389), .ZN(n19354) );
  OR2_X1 U12238 ( .A1(n20198), .A2(n10637), .ZN(n19387) );
  NOR2_X1 U12239 ( .A1(n10532), .A2(n10531), .ZN(n14292) );
  OR2_X1 U12240 ( .A1(n10500), .A2(n10499), .ZN(n14141) );
  OR2_X1 U12241 ( .A1(n10488), .A2(n10487), .ZN(n14016) );
  OR2_X1 U12242 ( .A1(n10475), .A2(n10474), .ZN(n14013) );
  OR2_X1 U12243 ( .A1(n10289), .A2(n10288), .ZN(n13636) );
  INV_X1 U12244 ( .A(n10164), .ZN(n10162) );
  INV_X1 U12245 ( .A(n19403), .ZN(n19411) );
  CLKBUF_X1 U12246 ( .A(n19415), .Z(n19406) );
  NAND2_X1 U12247 ( .A1(n19415), .A2(n13415), .ZN(n19403) );
  NOR2_X1 U12248 ( .A1(n10158), .A2(n9854), .ZN(n15256) );
  INV_X1 U12249 ( .A(n19417), .ZN(n15338) );
  NAND2_X1 U12250 ( .A1(n9851), .A2(n15272), .ZN(n15273) );
  NAND2_X1 U12251 ( .A1(n13945), .A2(n13946), .ZN(n14049) );
  AND2_X1 U12252 ( .A1(n15338), .A2(n15373), .ZN(n19437) );
  NOR2_X1 U12253 ( .A1(n13418), .A2(n13422), .ZN(n19394) );
  INV_X1 U12254 ( .A(n19428), .ZN(n19432) );
  OAI21_X1 U12255 ( .B1(n13391), .B2(n13390), .A(n13389), .ZN(n13392) );
  INV_X2 U12256 ( .A(n19445), .ZN(n19474) );
  INV_X1 U12257 ( .A(n13291), .ZN(n19486) );
  INV_X1 U12258 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15516) );
  NAND2_X1 U12259 ( .A1(n9695), .A2(n12308), .ZN(n15766) );
  AND2_X1 U12260 ( .A1(n16506), .A2(n19502), .ZN(n16494) );
  INV_X1 U12261 ( .A(n19507), .ZN(n19495) );
  INV_X1 U12262 ( .A(n19512), .ZN(n16436) );
  NAND2_X1 U12263 ( .A1(n13269), .A2(n12320), .ZN(n16506) );
  INV_X1 U12264 ( .A(n16506), .ZN(n19503) );
  AND2_X1 U12265 ( .A1(n16506), .A2(n20165), .ZN(n19512) );
  NAND2_X1 U12266 ( .A1(n16379), .A2(n19560), .ZN(n14513) );
  NAND2_X1 U12267 ( .A1(n15390), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15571) );
  NAND2_X1 U12268 ( .A1(n15144), .A2(n9823), .ZN(n15333) );
  NAND2_X1 U12269 ( .A1(n9939), .A2(n9940), .ZN(n15427) );
  OR2_X1 U12270 ( .A1(n12225), .A2(n9942), .ZN(n9939) );
  NOR2_X1 U12271 ( .A1(n15750), .A2(n15633), .ZN(n16046) );
  INV_X1 U12272 ( .A(n15701), .ZN(n16451) );
  AND2_X1 U12273 ( .A1(n13975), .A2(n13974), .ZN(n19306) );
  NAND2_X1 U12274 ( .A1(n10034), .A2(n9701), .ZN(n15746) );
  NAND2_X1 U12275 ( .A1(n12538), .A2(n12531), .ZN(n19554) );
  NAND2_X1 U12276 ( .A1(n12538), .A2(n12509), .ZN(n19533) );
  NAND2_X1 U12277 ( .A1(n19533), .A2(n12515), .ZN(n19549) );
  INV_X1 U12278 ( .A(n19554), .ZN(n19537) );
  INV_X1 U12279 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20182) );
  INV_X1 U12280 ( .A(n19394), .ZN(n20177) );
  INV_X1 U12281 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20163) );
  XNOR2_X1 U12282 ( .A(n13471), .B(n12552), .ZN(n20154) );
  OAI21_X1 U12283 ( .B1(n13477), .B2(n13469), .A(n13468), .ZN(n13471) );
  INV_X1 U12284 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16626) );
  INV_X1 U12285 ( .A(n13411), .ZN(n13412) );
  XNOR2_X1 U12286 ( .A(n13478), .B(n13477), .ZN(n15796) );
  INV_X1 U12287 ( .A(n20154), .ZN(n15819) );
  NOR2_X1 U12288 ( .A1(n19695), .A2(n19643), .ZN(n19691) );
  OAI21_X1 U12289 ( .B1(n19731), .B2(n19747), .A(n19995), .ZN(n19750) );
  NAND2_X1 U12290 ( .A1(n19753), .A2(n20151), .ZN(n19799) );
  OAI21_X1 U12291 ( .B1(n19790), .B2(n19812), .A(n19995), .ZN(n19815) );
  INV_X1 U12292 ( .A(n19799), .ZN(n19813) );
  INV_X1 U12293 ( .A(n19844), .ZN(n19845) );
  OAI21_X1 U12294 ( .B1(n19858), .B2(n19875), .A(n19995), .ZN(n19878) );
  NOR2_X1 U12295 ( .A1(n19786), .A2(n19643), .ZN(n19904) );
  NOR2_X1 U12296 ( .A1(n19818), .A2(n19643), .ZN(n19914) );
  OR2_X1 U12297 ( .A1(n19786), .A2(n19760), .ZN(n14162) );
  OAI21_X1 U12298 ( .B1(n14167), .B2(n14166), .A(n14165), .ZN(n19986) );
  INV_X1 U12299 ( .A(n14180), .ZN(n20002) );
  INV_X1 U12300 ( .A(n19926), .ZN(n20012) );
  INV_X1 U12301 ( .A(n19929), .ZN(n20019) );
  INV_X1 U12302 ( .A(n19935), .ZN(n20032) );
  INV_X1 U12303 ( .A(n19938), .ZN(n20039) );
  INV_X1 U12304 ( .A(n19612), .ZN(n20036) );
  INV_X1 U12305 ( .A(n14162), .ZN(n20055) );
  INV_X1 U12306 ( .A(n14332), .ZN(n20053) );
  INV_X1 U12307 ( .A(n19948), .ZN(n20054) );
  OR2_X1 U12308 ( .A1(n20064), .A2(n20065), .ZN(n16639) );
  NOR2_X1 U12309 ( .A1(n13745), .A2(n19920), .ZN(n16634) );
  NAND2_X1 U12310 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20074), .ZN(n20213) );
  NOR2_X1 U12311 ( .A1(n18954), .A2(n17727), .ZN(n19186) );
  NAND2_X1 U12312 ( .A1(n19169), .A2(n18955), .ZN(n17727) );
  AND2_X1 U12313 ( .A1(n9908), .A2(n19169), .ZN(n9907) );
  OR2_X1 U12314 ( .A1(n9793), .A2(n18957), .ZN(n9908) );
  NOR2_X1 U12315 ( .A1(n17830), .A2(n16895), .ZN(n16894) );
  NOR2_X1 U12316 ( .A1(n17849), .A2(n16918), .ZN(n16917) );
  NOR2_X1 U12317 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16967), .ZN(n16958) );
  AND2_X1 U12318 ( .A1(n17341), .A2(n16993), .ZN(n16987) );
  NOR2_X1 U12319 ( .A1(n19013), .A2(n13256), .ZN(n17155) );
  NAND4_X1 U12320 ( .A1(n18375), .A2(n13259), .A3(n19028), .A4(n19018), .ZN(
        n17196) );
  NOR2_X1 U12321 ( .A1(n16928), .A2(n17263), .ZN(n17269) );
  NOR4_X1 U12322 ( .A1(n17341), .A2(n15910), .A3(n17520), .A4(n17340), .ZN(
        n17328) );
  NAND4_X1 U12323 ( .A1(n19169), .A2(n19171), .A3(n17689), .A4(n16034), .ZN(
        n17520) );
  AOI21_X1 U12324 ( .B1(n17545), .B2(n17680), .A(n9887), .ZN(n9886) );
  NOR2_X1 U12325 ( .A1(n17673), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n9887) );
  INV_X1 U12326 ( .A(P3_EAX_REG_31__SCAN_IN), .ZN(n9885) );
  INV_X1 U12327 ( .A(n17545), .ZN(n17540) );
  NOR2_X1 U12328 ( .A1(n17753), .A2(n17554), .ZN(n17548) );
  NOR2_X1 U12329 ( .A1(n17749), .A2(n17563), .ZN(n17557) );
  NAND2_X1 U12330 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17564), .ZN(n17563) );
  NAND2_X1 U12331 ( .A1(n17574), .A2(n9749), .ZN(n17568) );
  NAND2_X1 U12332 ( .A1(n9868), .A2(n9866), .ZN(n17623) );
  NOR2_X1 U12333 ( .A1(n17535), .A2(n9867), .ZN(n9866) );
  INV_X1 U12334 ( .A(n17652), .ZN(n9868) );
  NOR2_X1 U12335 ( .A1(n17779), .A2(n17645), .ZN(n17640) );
  NOR2_X1 U12336 ( .A1(n17621), .A2(n17673), .ZN(n17658) );
  AOI211_X2 U12337 ( .C1(n15895), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n12936), .B(n12935), .ZN(n17660) );
  INV_X1 U12338 ( .A(n13016), .ZN(n17675) );
  INV_X1 U12339 ( .A(n17683), .ZN(n17676) );
  INV_X1 U12340 ( .A(n17684), .ZN(n17679) );
  NOR2_X1 U12341 ( .A1(n13020), .A2(n13019), .ZN(n13029) );
  NOR2_X1 U12342 ( .A1(n16037), .A2(n16038), .ZN(n17684) );
  NOR2_X1 U12343 ( .A1(n19166), .A2(n17690), .ZN(n17703) );
  CLKBUF_X1 U12344 ( .A(n17703), .Z(n17723) );
  CLKBUF_X1 U12346 ( .A(n17790), .Z(n17782) );
  OAI211_X1 U12347 ( .C1(n18498), .C2(n19165), .A(n17729), .B(n17728), .ZN(
        n17790) );
  OAI21_X1 U12348 ( .B1(n17812), .B2(n17968), .A(n16699), .ZN(n17808) );
  NAND2_X1 U12349 ( .A1(n18041), .A2(n9832), .ZN(n17820) );
  INV_X1 U12350 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17991) );
  INV_X1 U12351 ( .A(n18058), .ZN(n18044) );
  NOR2_X2 U12352 ( .A1(n17656), .A2(n18151), .ZN(n18058) );
  INV_X1 U12353 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18065) );
  AND2_X1 U12354 ( .A1(n18106), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18086) );
  INV_X1 U12355 ( .A(n18147), .ZN(n18118) );
  INV_X1 U12356 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18117) );
  NAND2_X1 U12357 ( .A1(n18857), .A2(n15932), .ZN(n18717) );
  INV_X1 U12358 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18133) );
  NOR2_X2 U12359 ( .A1(n19171), .A2(n16815), .ZN(n18136) );
  INV_X1 U12360 ( .A(n18136), .ZN(n18152) );
  NOR2_X1 U12361 ( .A1(n16680), .A2(n18395), .ZN(n16681) );
  NAND2_X1 U12362 ( .A1(n10018), .A2(n17968), .ZN(n17841) );
  NAND2_X1 U12363 ( .A1(n17897), .A2(n10070), .ZN(n17848) );
  INV_X1 U12364 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19183) );
  NAND2_X1 U12365 ( .A1(n18022), .A2(n9829), .ZN(n17955) );
  NAND2_X1 U12366 ( .A1(n18022), .A2(n18363), .ZN(n18017) );
  NAND2_X1 U12367 ( .A1(n18009), .A2(n13047), .ZN(n18396) );
  NOR3_X2 U12368 ( .A1(n17656), .A2(n18959), .A3(n18460), .ZN(n18391) );
  INV_X1 U12369 ( .A(n10072), .ZN(n18067) );
  NAND2_X1 U12370 ( .A1(n10008), .A2(n10007), .ZN(n18074) );
  NAND2_X1 U12371 ( .A1(n18088), .A2(n18089), .ZN(n18087) );
  INV_X1 U12372 ( .A(n10004), .ZN(n18128) );
  INV_X1 U12373 ( .A(n18468), .ZN(n18476) );
  INV_X1 U12374 ( .A(n18458), .ZN(n18474) );
  INV_X1 U12375 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18487) );
  INV_X1 U12376 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18996) );
  INV_X1 U12377 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19001) );
  INV_X1 U12378 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19004) );
  AOI211_X1 U12379 ( .C1(n19169), .C2(n18987), .A(n18492), .B(n15944), .ZN(
        n19152) );
  INV_X1 U12380 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18963) );
  INV_X1 U12381 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18501) );
  INV_X1 U12382 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18528) );
  INV_X1 U12383 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18740) );
  INV_X1 U12384 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n18806) );
  NAND2_X1 U12385 ( .A1(n19045), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19181) );
  AND2_X2 U12386 ( .A1(n11931), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n13800)
         );
  CLKBUF_X1 U12387 ( .A(n16797), .Z(n16801) );
  OAI21_X1 U12388 ( .B1(n14971), .B2(n20226), .A(n9783), .ZN(P1_U2968) );
  INV_X1 U12389 ( .A(n10640), .ZN(n10898) );
  NOR2_X1 U12390 ( .A1(n12885), .A2(n12884), .ZN(n12886) );
  INV_X1 U12391 ( .A(n12905), .ZN(n12908) );
  OR2_X1 U12392 ( .A1(n12323), .A2(n10092), .ZN(n12326) );
  OR2_X1 U12393 ( .A1(n16867), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9915) );
  AOI211_X1 U12394 ( .C1(n16857), .C2(n17173), .A(n16856), .B(n16855), .ZN(
        n16860) );
  OAI21_X1 U12395 ( .B1(n17539), .B2(P3_EAX_REG_31__SCAN_IN), .A(n9882), .ZN(
        P3_U2704) );
  NOR2_X1 U12396 ( .A1(n9884), .A2(n9883), .ZN(n9882) );
  AND2_X1 U12397 ( .A1(n17610), .A2(BUF2_REG_31__SCAN_IN), .ZN(n9883) );
  NOR2_X1 U12398 ( .A1(n9886), .A2(n9885), .ZN(n9884) );
  NAND2_X1 U12399 ( .A1(n17574), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n17573) );
  OR3_X1 U12400 ( .A1(n19025), .A2(n19024), .A3(n19023), .ZN(n19026) );
  AOI21_X1 U12401 ( .B1(n10058), .B2(n10056), .A(n9766), .ZN(n10055) );
  OR2_X1 U12402 ( .A1(n10039), .A2(n10038), .ZN(n9724) );
  NAND2_X2 U12403 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12925), .ZN(
        n12943) );
  NAND3_X2 U12404 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15804) );
  INV_X1 U12405 ( .A(n18009), .ZN(n13224) );
  NAND2_X1 U12406 ( .A1(n14664), .A2(n9805), .ZN(n9725) );
  NAND2_X1 U12407 ( .A1(n14602), .A2(n10185), .ZN(n14590) );
  OR2_X1 U12408 ( .A1(n14590), .A2(n10131), .ZN(n9726) );
  AND2_X1 U12409 ( .A1(n15443), .A2(n10148), .ZN(n9727) );
  NOR2_X1 U12410 ( .A1(n15284), .A2(n9798), .ZN(n15141) );
  NAND2_X1 U12411 ( .A1(n14664), .A2(n14666), .ZN(n14665) );
  OR2_X1 U12412 ( .A1(n14339), .A2(n11835), .ZN(n9728) );
  AND2_X1 U12413 ( .A1(n12778), .A2(n9824), .ZN(n9729) );
  NAND2_X1 U12414 ( .A1(n10052), .A2(n10055), .ZN(n14903) );
  NOR2_X1 U12415 ( .A1(n15284), .A2(n15483), .ZN(n15174) );
  AND2_X1 U12416 ( .A1(n9904), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9730) );
  AND2_X1 U12417 ( .A1(n9940), .A2(n9771), .ZN(n9731) );
  AND2_X1 U12418 ( .A1(n9921), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9732) );
  AND2_X1 U12419 ( .A1(n10083), .A2(n12237), .ZN(n9733) );
  INV_X1 U12420 ( .A(n14375), .ZN(n14451) );
  AND2_X1 U12421 ( .A1(n10885), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9734) );
  AND2_X1 U12422 ( .A1(n10738), .A2(n11959), .ZN(n9735) );
  AND2_X1 U12423 ( .A1(n9951), .A2(n16499), .ZN(n9736) );
  INV_X1 U12424 ( .A(n11941), .ZN(n11959) );
  NAND2_X1 U12425 ( .A1(n10731), .A2(n10730), .ZN(n11941) );
  AND2_X1 U12426 ( .A1(n12495), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9737) );
  NOR2_X1 U12427 ( .A1(n12415), .A2(n16132), .ZN(n9738) );
  NAND2_X1 U12428 ( .A1(n9698), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11132) );
  AND2_X1 U12429 ( .A1(n9960), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9739) );
  INV_X1 U12430 ( .A(n13384), .ZN(n14537) );
  AND2_X1 U12431 ( .A1(n11952), .A2(n11956), .ZN(n19513) );
  OR2_X1 U12432 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n11177) );
  NAND2_X1 U12433 ( .A1(n12538), .A2(n20189), .ZN(n19556) );
  NAND2_X1 U12434 ( .A1(n14299), .A2(n9801), .ZN(n15280) );
  NOR2_X1 U12435 ( .A1(n16532), .A2(n9804), .ZN(n9740) );
  AND2_X1 U12436 ( .A1(n9963), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9741) );
  AND2_X1 U12437 ( .A1(n9969), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9742) );
  AND2_X1 U12438 ( .A1(n10134), .A2(n9821), .ZN(n9743) );
  AND2_X1 U12439 ( .A1(n17537), .A2(n17578), .ZN(n17641) );
  INV_X2 U12440 ( .A(n17641), .ZN(n17680) );
  INV_X1 U12441 ( .A(n15500), .ZN(n10038) );
  AND2_X1 U12442 ( .A1(n9896), .A2(n14945), .ZN(n9744) );
  AND2_X1 U12443 ( .A1(n10115), .A2(n16401), .ZN(n9745) );
  AND2_X1 U12444 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9746) );
  AND2_X1 U12445 ( .A1(n9966), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9747) );
  AND2_X1 U12446 ( .A1(n18057), .A2(n15966), .ZN(n9748) );
  AND2_X1 U12447 ( .A1(n9869), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n9749) );
  NAND3_X1 U12448 ( .A1(n10222), .A2(n10221), .A3(n9992), .ZN(n12733) );
  AND2_X1 U12449 ( .A1(n16644), .A2(n18256), .ZN(n9750) );
  AND2_X1 U12450 ( .A1(n10148), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9751) );
  OR2_X1 U12451 ( .A1(n14727), .A2(n14667), .ZN(n9752) );
  INV_X2 U12452 ( .A(n17486), .ZN(n17393) );
  INV_X2 U12453 ( .A(n12919), .ZN(n15828) );
  AND2_X1 U12454 ( .A1(n18041), .A2(n9750), .ZN(n9753) );
  AND2_X2 U12455 ( .A1(n9712), .A2(n10282), .ZN(n10360) );
  NAND2_X1 U12456 ( .A1(n15742), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15724) );
  OR3_X1 U12457 ( .A1(n9752), .A2(n9984), .A3(n14615), .ZN(n9754) );
  AND2_X1 U12458 ( .A1(n14664), .A2(n10124), .ZN(n14653) );
  OR2_X1 U12459 ( .A1(n18974), .A2(n12927), .ZN(n9755) );
  NOR2_X1 U12460 ( .A1(n14437), .A2(n14463), .ZN(n14462) );
  NAND2_X1 U12461 ( .A1(n12145), .A2(n12146), .ZN(n14344) );
  AND4_X1 U12462 ( .A1(n13027), .A2(n13026), .A3(n13025), .A4(n13024), .ZN(
        n9757) );
  NAND2_X2 U12463 ( .A1(n13043), .A2(n16687), .ZN(n17968) );
  AND3_X1 U12464 ( .A1(n14508), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n10193), .ZN(n9758) );
  NAND2_X1 U12465 ( .A1(n10054), .A2(n10058), .ZN(n14927) );
  AND4_X1 U12466 ( .A1(n10937), .A2(n10936), .A3(n10935), .A4(n10934), .ZN(
        n9759) );
  AND2_X1 U12467 ( .A1(n16135), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9760) );
  AND4_X1 U12468 ( .A1(n10918), .A2(n10917), .A3(n10916), .A4(n10915), .ZN(
        n9761) );
  OR3_X1 U12469 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17870), .ZN(n9762) );
  NAND2_X1 U12470 ( .A1(n11204), .A2(n13841), .ZN(n9763) );
  AND2_X1 U12471 ( .A1(n10873), .A2(n10098), .ZN(n9764) );
  NAND2_X1 U12472 ( .A1(n12225), .A2(n15446), .ZN(n15434) );
  AND3_X1 U12473 ( .A1(n12229), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n12162), .ZN(n9765) );
  NAND2_X1 U12474 ( .A1(n15443), .A2(n9751), .ZN(n15413) );
  INV_X1 U12475 ( .A(n12552), .ZN(n13470) );
  XNOR2_X1 U12476 ( .A(n15241), .B(n12897), .ZN(n12322) );
  NAND2_X1 U12477 ( .A1(n13174), .A2(n17538), .ZN(n15947) );
  INV_X1 U12478 ( .A(n15947), .ZN(n13166) );
  AND2_X1 U12479 ( .A1(n15065), .A2(n16259), .ZN(n9766) );
  NAND2_X2 U12481 ( .A1(n9687), .A2(n16615), .ZN(n10885) );
  NAND2_X1 U12482 ( .A1(n15247), .A2(n12803), .ZN(n15255) );
  AND2_X1 U12483 ( .A1(n12574), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n9767) );
  AND2_X1 U12484 ( .A1(n9733), .A2(n15559), .ZN(n9768) );
  AND3_X1 U12485 ( .A1(n12961), .A2(n12960), .A3(n10170), .ZN(n9769) );
  AND2_X1 U12486 ( .A1(n13416), .A2(n19541), .ZN(n9770) );
  NAND2_X1 U12487 ( .A1(n10135), .A2(n9743), .ZN(n10137) );
  OR2_X1 U12488 ( .A1(n15425), .A2(n15610), .ZN(n9771) );
  NOR2_X1 U12489 ( .A1(n13046), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9772) );
  AND2_X1 U12490 ( .A1(n15157), .A2(n15158), .ZN(n15144) );
  NOR2_X1 U12491 ( .A1(n15062), .A2(n12419), .ZN(n9774) );
  AND2_X1 U12492 ( .A1(n9849), .A2(n15269), .ZN(n9775) );
  INV_X1 U12493 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9992) );
  AND2_X1 U12494 ( .A1(n9919), .A2(n9916), .ZN(n9776) );
  INV_X1 U12495 ( .A(n16175), .ZN(n10050) );
  AND2_X1 U12496 ( .A1(n9848), .A2(n9845), .ZN(n9777) );
  AOI211_X1 U12497 ( .C1(n15895), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n13117), .B(n13116), .ZN(n18509) );
  AND2_X1 U12498 ( .A1(n9843), .A2(n9841), .ZN(n9778) );
  AND4_X1 U12499 ( .A1(n12988), .A2(n12987), .A3(n12986), .A4(n12985), .ZN(
        n9779) );
  AND2_X1 U12500 ( .A1(n14225), .A2(n16175), .ZN(n9780) );
  AND2_X1 U12501 ( .A1(n15425), .A2(n15610), .ZN(n9781) );
  AND2_X1 U12502 ( .A1(n15387), .A2(n15386), .ZN(n9782) );
  AND2_X1 U12503 ( .A1(n12445), .A2(n12444), .ZN(n9783) );
  INV_X1 U12504 ( .A(n12306), .ZN(n9951) );
  INV_X1 U12505 ( .A(n10023), .ZN(n10022) );
  NAND2_X1 U12506 ( .A1(n13047), .A2(n18256), .ZN(n10023) );
  AND2_X1 U12507 ( .A1(n15305), .A2(n10564), .ZN(n15296) );
  INV_X1 U12508 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10221) );
  AND4_X1 U12509 ( .A1(n10251), .A2(n10250), .A3(n10249), .A4(n10248), .ZN(
        n9784) );
  AND2_X1 U12510 ( .A1(n12570), .A2(n12569), .ZN(n13466) );
  NAND2_X1 U12511 ( .A1(n10737), .A2(n10736), .ZN(n11960) );
  NAND2_X1 U12512 ( .A1(n15144), .A2(n15145), .ZN(n15146) );
  NOR2_X1 U12513 ( .A1(n14590), .A2(n14591), .ZN(n14572) );
  NOR2_X1 U12514 ( .A1(n10750), .A2(n10749), .ZN(n9785) );
  INV_X1 U12515 ( .A(n10058), .ZN(n10057) );
  INV_X1 U12516 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10222) );
  AND2_X1 U12517 ( .A1(n15259), .A2(n10105), .ZN(n9786) );
  XNOR2_X1 U12518 ( .A(n13418), .B(n12559), .ZN(n13411) );
  NOR3_X1 U12519 ( .A1(n17820), .A2(n16647), .A3(n16646), .ZN(n9787) );
  INV_X1 U12520 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10283) );
  INV_X1 U12521 ( .A(n17682), .ZN(n13195) );
  NAND2_X1 U12522 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13042), .ZN(
        n9788) );
  AND3_X1 U12523 ( .A1(n10034), .A2(n9701), .A3(n10026), .ZN(n9789) );
  AND2_X1 U12524 ( .A1(n9945), .A2(n12218), .ZN(n9790) );
  AND2_X1 U12525 ( .A1(n10703), .A2(n12495), .ZN(n9791) );
  NOR2_X1 U12526 ( .A1(n12921), .A2(n12926), .ZN(n12962) );
  INV_X1 U12527 ( .A(n12962), .ZN(n12977) );
  INV_X1 U12528 ( .A(n10742), .ZN(n10757) );
  BUF_X1 U12529 ( .A(n10742), .Z(n10848) );
  INV_X1 U12530 ( .A(n11173), .ZN(n11403) );
  INV_X1 U12531 ( .A(n11403), .ZN(n11497) );
  AND4_X2 U12532 ( .A1(n10312), .A2(n10311), .A3(n10310), .A4(n10309), .ZN(
        n12101) );
  NAND2_X1 U12533 ( .A1(n12558), .A2(n12557), .ZN(n13418) );
  NAND2_X1 U12534 ( .A1(n13812), .A2(n13992), .ZN(n11803) );
  NAND2_X1 U12535 ( .A1(n17897), .A2(n17884), .ZN(n17885) );
  NAND2_X1 U12536 ( .A1(n13972), .A2(n13973), .ZN(n13974) );
  AND2_X1 U12537 ( .A1(n14299), .A2(n10155), .ZN(n9792) );
  NAND2_X1 U12538 ( .A1(n14294), .A2(n14295), .ZN(n14293) );
  AND2_X1 U12539 ( .A1(n16689), .A2(n18958), .ZN(n9793) );
  OR2_X1 U12540 ( .A1(n15483), .A2(n10079), .ZN(n9794) );
  AND2_X1 U12541 ( .A1(n10209), .A2(n9963), .ZN(n9795) );
  AND2_X1 U12542 ( .A1(n10214), .A2(n9969), .ZN(n9796) );
  INV_X1 U12543 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n20201) );
  INV_X1 U12544 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20156) );
  AND3_X1 U12545 ( .A1(n9917), .A2(n9776), .A3(n9918), .ZN(n9797) );
  OR2_X1 U12546 ( .A1(n9794), .A2(n15154), .ZN(n9798) );
  OR2_X1 U12547 ( .A1(n10187), .A2(n12631), .ZN(n9799) );
  AND2_X1 U12548 ( .A1(n14153), .A2(n10120), .ZN(n9800) );
  AND3_X1 U12549 ( .A1(n11293), .A2(n14152), .A3(n14151), .ZN(n14153) );
  NOR2_X1 U12550 ( .A1(n15733), .A2(n10099), .ZN(n13972) );
  AND2_X1 U12551 ( .A1(n10155), .A2(n15281), .ZN(n9801) );
  AND2_X1 U12552 ( .A1(n14295), .A2(n10114), .ZN(n9802) );
  AND2_X1 U12553 ( .A1(n14464), .A2(n9989), .ZN(n9803) );
  OR2_X1 U12554 ( .A1(n9999), .A2(n14042), .ZN(n9804) );
  AND2_X1 U12555 ( .A1(n10166), .A2(n10124), .ZN(n9805) );
  AND2_X1 U12556 ( .A1(n17574), .A2(n9869), .ZN(n9806) );
  INV_X1 U12557 ( .A(n15489), .ZN(n10039) );
  INV_X1 U12558 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11133) );
  OR2_X1 U12559 ( .A1(n15284), .A2(n9794), .ZN(n9807) );
  OR2_X1 U12560 ( .A1(n9752), .A2(n9984), .ZN(n9808) );
  NOR2_X1 U12561 ( .A1(n12407), .A2(n12406), .ZN(n9809) );
  NAND2_X1 U12562 ( .A1(n15092), .A2(n16106), .ZN(n9810) );
  AND2_X1 U12563 ( .A1(n9739), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9811) );
  INV_X1 U12564 ( .A(n9864), .ZN(n18978) );
  NAND2_X1 U12565 ( .A1(n18976), .A2(n9865), .ZN(n9864) );
  INV_X1 U12566 ( .A(n12553), .ZN(n12562) );
  NAND2_X1 U12567 ( .A1(n20201), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12553) );
  AND2_X1 U12568 ( .A1(n14153), .A2(n14277), .ZN(n9812) );
  OR2_X1 U12569 ( .A1(n9798), .A2(n10078), .ZN(n9813) );
  OR2_X1 U12570 ( .A1(n9804), .A2(n10001), .ZN(n9814) );
  AND2_X1 U12571 ( .A1(n10061), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9815) );
  AND2_X1 U12572 ( .A1(n10112), .A2(n15504), .ZN(n9816) );
  AND2_X1 U12573 ( .A1(n9805), .A2(n14643), .ZN(n9817) );
  AND2_X1 U12574 ( .A1(n9732), .A2(n9920), .ZN(n9818) );
  AND2_X1 U12575 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_EBX_REG_3__SCAN_IN), 
        .ZN(n9819) );
  INV_X1 U12576 ( .A(n9924), .ZN(n17182) );
  NOR2_X1 U12577 ( .A1(n13648), .A2(n13792), .ZN(n9978) );
  AND3_X1 U12578 ( .A1(n9898), .A2(n13384), .A3(n13802), .ZN(n13338) );
  NAND2_X1 U12579 ( .A1(n12538), .A2(n12521), .ZN(n19540) );
  INV_X1 U12580 ( .A(n19540), .ZN(n19560) );
  NOR2_X1 U12581 ( .A1(n13545), .A2(n10163), .ZN(n13635) );
  NAND2_X1 U12582 ( .A1(n12575), .A2(n9746), .ZN(n13546) );
  INV_X1 U12583 ( .A(n12064), .ZN(n14186) );
  NAND2_X1 U12584 ( .A1(n12528), .A2(n12495), .ZN(n10705) );
  AND2_X1 U12585 ( .A1(n17900), .A2(n9921), .ZN(n9820) );
  AND2_X1 U12586 ( .A1(n9709), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10504) );
  INV_X1 U12587 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n9995) );
  NOR2_X1 U12588 ( .A1(n10136), .A2(n14463), .ZN(n9821) );
  INV_X1 U12589 ( .A(n12575), .ZN(n13545) );
  AND2_X1 U12590 ( .A1(n10196), .A2(n9966), .ZN(n9822) );
  AND2_X1 U12591 ( .A1(n9998), .A2(n15145), .ZN(n9823) );
  INV_X1 U12592 ( .A(n15757), .ZN(n10032) );
  INV_X1 U12593 ( .A(n19169), .ZN(n19020) );
  NOR2_X1 U12594 ( .A1(n18302), .A2(n18290), .ZN(n18256) );
  OR2_X1 U12595 ( .A1(n14279), .A2(n11828), .ZN(n14338) );
  INV_X1 U12596 ( .A(n14338), .ZN(n9981) );
  AND2_X1 U12597 ( .A1(n12775), .A2(n12796), .ZN(n9824) );
  NOR2_X1 U12598 ( .A1(n13545), .A2(n10162), .ZN(n13689) );
  AND2_X1 U12599 ( .A1(n10120), .A2(n14376), .ZN(n9825) );
  OR2_X1 U12600 ( .A1(n10407), .A2(n10406), .ZN(n12034) );
  AND2_X1 U12601 ( .A1(n9823), .A2(n9997), .ZN(n9826) );
  INV_X1 U12602 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15171) );
  INV_X1 U12603 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n9923) );
  AND2_X1 U12604 ( .A1(n16660), .A2(n9927), .ZN(n9827) );
  AND2_X1 U12605 ( .A1(n16660), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9828) );
  AND2_X1 U12606 ( .A1(n10074), .A2(n17981), .ZN(n9829) );
  NAND2_X1 U12607 ( .A1(n11817), .A2(n11816), .ZN(n9830) );
  INV_X1 U12608 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9928) );
  INV_X2 U12609 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15781) );
  AND4_X1 U12610 ( .A1(n16218), .A2(n15045), .A3(n15044), .A4(n14954), .ZN(
        n9831) );
  INV_X1 U12611 ( .A(n18977), .ZN(n9904) );
  AND2_X1 U12612 ( .A1(n9750), .A2(n16645), .ZN(n9832) );
  INV_X1 U12613 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n9929) );
  INV_X1 U12614 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n9870) );
  INV_X1 U12615 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n9871) );
  INV_X1 U12616 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n9931) );
  INV_X1 U12617 ( .A(n14984), .ZN(n10062) );
  INV_X1 U12618 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n9878) );
  INV_X1 U12619 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n9967) );
  AND2_X1 U12620 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n19135), .ZN(
        n9833) );
  INV_X1 U12621 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9970) );
  AND2_X1 U12622 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n9834) );
  INV_X1 U12623 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10097) );
  NOR2_X1 U12624 ( .A1(n16687), .A2(n18151), .ZN(n18008) );
  AOI211_X1 U12625 ( .C1(n17490), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n13010), .B(n13009), .ZN(n13011) );
  OR3_X1 U12626 ( .A1(n12261), .A2(n12101), .A3(n12527), .ZN(n12887) );
  OR2_X1 U12627 ( .A1(n16372), .A2(n12101), .ZN(n15425) );
  NOR2_X1 U12628 ( .A1(n15151), .A2(n12101), .ZN(n12228) );
  NOR2_X1 U12629 ( .A1(n19232), .A2(n12101), .ZN(n12215) );
  OR2_X1 U12630 ( .A1(n19322), .A2(n12101), .ZN(n12172) );
  NOR3_X2 U12631 ( .A1(n19023), .A2(n18996), .A3(n18621), .ZN(n18595) );
  AOI211_X2 U12632 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(n18888), .A(n18799), 
        .B(n18798), .ZN(n18826) );
  AOI22_X2 U12633 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n13871), .B1(DATAI_24_), 
        .B2(n13870), .ZN(n20754) );
  NOR2_X1 U12634 ( .A1(n13800), .A2(n16120), .ZN(n13870) );
  NOR2_X1 U12635 ( .A1(n16120), .A2(n13799), .ZN(n13871) );
  NOR3_X2 U12636 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19023), .A3(
        n18713), .ZN(n18685) );
  NOR2_X1 U12637 ( .A1(n13170), .A2(n15948), .ZN(n18967) );
  NAND2_X1 U12638 ( .A1(n13171), .A2(n15948), .ZN(n15935) );
  NOR2_X1 U12639 ( .A1(n13162), .A2(n15948), .ZN(n13180) );
  INV_X1 U12640 ( .A(n15948), .ZN(n18503) );
  NAND3_X1 U12641 ( .A1(n10602), .A2(n9846), .A3(n10601), .ZN(n9836) );
  NAND3_X1 U12642 ( .A1(n10600), .A2(n9840), .A3(n10599), .ZN(n9838) );
  NAND2_X1 U12643 ( .A1(n10622), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n9845) );
  NAND2_X1 U12644 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n9846) );
  NAND2_X1 U12645 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n9847) );
  NAND2_X1 U12646 ( .A1(n12849), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n9848) );
  NOR2_X1 U12647 ( .A1(n9849), .A2(n15269), .ZN(n15267) );
  NAND3_X1 U12648 ( .A1(n12573), .A2(n12572), .A3(n10149), .ZN(n9850) );
  INV_X1 U12649 ( .A(n12753), .ZN(n9851) );
  INV_X1 U12650 ( .A(n12755), .ZN(n9852) );
  OAI21_X1 U12651 ( .B1(n12502), .B2(n9853), .A(n10690), .ZN(n10697) );
  NAND2_X1 U12652 ( .A1(n12508), .A2(n9819), .ZN(n10741) );
  INV_X1 U12653 ( .A(n10845), .ZN(n10834) );
  NAND2_X1 U12654 ( .A1(n10845), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10675) );
  NAND2_X1 U12655 ( .A1(n10845), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10720) );
  NAND2_X1 U12656 ( .A1(n10845), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10733) );
  AND2_X1 U12657 ( .A1(n9855), .A2(n9856), .ZN(n12013) );
  NAND2_X1 U12658 ( .A1(n9857), .A2(n11952), .ZN(n12558) );
  AND2_X1 U12659 ( .A1(n12471), .A2(n9859), .ZN(n12478) );
  NAND3_X1 U12660 ( .A1(n10688), .A2(n10687), .A3(n10657), .ZN(n9859) );
  OAI22_X2 U12661 ( .A1(n19492), .A2(n19490), .B1(n19520), .B2(n19363), .ZN(
        n16496) );
  NAND2_X1 U12662 ( .A1(n14022), .A2(n12123), .ZN(n19492) );
  NAND2_X2 U12663 ( .A1(n15715), .A2(n15454), .ZN(n15701) );
  OR2_X2 U12664 ( .A1(n15512), .A2(n15513), .ZN(n15510) );
  NAND2_X1 U12665 ( .A1(n9860), .A2(n10708), .ZN(n11954) );
  OAI21_X1 U12666 ( .B1(n10747), .B2(n9791), .A(n9861), .ZN(n9860) );
  NAND3_X1 U12667 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_8__SCAN_IN), 
        .A3(P3_EAX_REG_13__SCAN_IN), .ZN(n9867) );
  NAND3_X1 U12668 ( .A1(n13120), .A2(n9874), .A3(n9873), .ZN(n9872) );
  NAND2_X1 U12669 ( .A1(n9698), .A2(n9890), .ZN(n9889) );
  NAND4_X1 U12670 ( .A1(n13841), .A2(n11184), .A3(n11183), .A4(n10122), .ZN(
        n11281) );
  XNOR2_X2 U12671 ( .A(n11154), .B(n11153), .ZN(n11184) );
  NAND2_X2 U12672 ( .A1(n9893), .A2(n9774), .ZN(n14897) );
  NAND2_X1 U12673 ( .A1(n9898), .A2(n13384), .ZN(n13589) );
  AND3_X2 U12674 ( .A1(n12342), .A2(n11743), .A3(n10965), .ZN(n9898) );
  INV_X1 U12675 ( .A(n9898), .ZN(n13379) );
  AND2_X2 U12676 ( .A1(n10908), .A2(n14062), .ZN(n11145) );
  OAI21_X1 U12677 ( .B1(n15996), .B2(n10908), .A(n14087), .ZN(n14101) );
  NAND2_X2 U12678 ( .A1(n9730), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n17470) );
  INV_X1 U12679 ( .A(n18151), .ZN(n18140) );
  NAND2_X1 U12680 ( .A1(n13167), .A2(n9910), .ZN(n15936) );
  INV_X1 U12681 ( .A(n13168), .ZN(n9914) );
  NAND3_X1 U12682 ( .A1(n16860), .A2(n16859), .A3(n9915), .ZN(P3_U2641) );
  NAND4_X1 U12683 ( .A1(n9917), .A2(n9776), .A3(n9918), .A4(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17912) );
  NAND3_X1 U12684 ( .A1(n9917), .A2(n9918), .A3(n9919), .ZN(n17945) );
  XOR2_X1 U12685 ( .A(n9930), .B(n9929), .Z(n9924) );
  NAND2_X2 U12686 ( .A1(n9932), .A2(n20199), .ZN(n12468) );
  INV_X1 U12687 ( .A(n10683), .ZN(n9932) );
  OR2_X1 U12688 ( .A1(n12256), .A2(n15396), .ZN(n9933) );
  NAND2_X1 U12689 ( .A1(n9933), .A2(n9934), .ZN(n15377) );
  NAND2_X2 U12690 ( .A1(n11987), .A2(n9770), .ZN(n12064) );
  AND2_X2 U12691 ( .A1(n13472), .A2(n13423), .ZN(n11987) );
  NAND2_X1 U12692 ( .A1(n12225), .A2(n9731), .ZN(n9938) );
  INV_X1 U12693 ( .A(n12164), .ZN(n9943) );
  NAND2_X1 U12694 ( .A1(n12297), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9949) );
  NAND2_X1 U12695 ( .A1(n12296), .A2(n9696), .ZN(n9950) );
  NAND2_X1 U12696 ( .A1(n16498), .A2(n16499), .ZN(n16497) );
  NAND2_X1 U12697 ( .A1(n10739), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10677) );
  NAND2_X2 U12698 ( .A1(n9953), .A2(n9952), .ZN(n10739) );
  OR2_X2 U12699 ( .A1(n10646), .A2(n10645), .ZN(n10699) );
  NAND3_X1 U12700 ( .A1(n13416), .A2(n9954), .A3(n13423), .ZN(n11968) );
  INV_X1 U12701 ( .A(n13472), .ZN(n9954) );
  XNOR2_X1 U12702 ( .A(n12035), .B(n12034), .ZN(n19493) );
  AND2_X2 U12703 ( .A1(n10090), .A2(n10091), .ZN(n12035) );
  NAND2_X1 U12704 ( .A1(n15668), .A2(n9957), .ZN(n15670) );
  NAND2_X1 U12705 ( .A1(n19556), .A2(n12515), .ZN(n9957) );
  INV_X1 U12706 ( .A(n11803), .ZN(n11785) );
  NAND3_X2 U12707 ( .A1(n9761), .A2(n9971), .A3(n10922), .ZN(n13812) );
  NAND2_X1 U12708 ( .A1(n14586), .A2(n9990), .ZN(n14520) );
  MUX2_X1 U12709 ( .A(n14521), .B(n11808), .S(n14520), .Z(n9991) );
  NAND2_X1 U12710 ( .A1(n13945), .A2(n9996), .ZN(n14051) );
  AND2_X2 U12711 ( .A1(n15144), .A2(n9826), .ZN(n15323) );
  INV_X2 U12712 ( .A(n10566), .ZN(n10544) );
  NAND3_X1 U12713 ( .A1(n12866), .A2(n10276), .A3(P2_REIP_REG_1__SCAN_IN), 
        .ZN(n10002) );
  NOR2_X1 U12714 ( .A1(n13060), .A2(n9833), .ZN(n10003) );
  XNOR2_X1 U12715 ( .A(n13033), .B(n18443), .ZN(n18127) );
  INV_X1 U12716 ( .A(n18073), .ZN(n10006) );
  NAND3_X1 U12717 ( .A1(n10008), .A2(n10006), .A3(n10007), .ZN(n10011) );
  INV_X1 U12718 ( .A(n10011), .ZN(n18072) );
  INV_X1 U12719 ( .A(n10018), .ZN(n17847) );
  OAI21_X1 U12720 ( .B1(n17842), .B2(n18180), .A(n10016), .ZN(n17824) );
  NAND2_X1 U12721 ( .A1(n10024), .A2(n13050), .ZN(n13051) );
  AND2_X2 U12722 ( .A1(n10025), .A2(n9683), .ZN(n10692) );
  NAND2_X1 U12723 ( .A1(n10025), .A2(n12472), .ZN(n12264) );
  NOR2_X2 U12724 ( .A1(n10631), .A2(n10615), .ZN(n10025) );
  AND2_X2 U12725 ( .A1(n10621), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12620) );
  AND2_X2 U12726 ( .A1(n15701), .A2(n10035), .ZN(n15455) );
  OAI21_X1 U12727 ( .B1(n15510), .B2(n9724), .A(n10036), .ZN(n15482) );
  XNOR2_X2 U12728 ( .A(n11115), .B(n11058), .ZN(n11172) );
  NAND2_X1 U12729 ( .A1(n14879), .A2(n15065), .ZN(n10046) );
  NAND2_X1 U12730 ( .A1(n14224), .A2(n9780), .ZN(n10047) );
  OAI21_X1 U12731 ( .B1(n14391), .B2(n12410), .A(n12409), .ZN(n14409) );
  NAND2_X1 U12732 ( .A1(n14830), .A2(n9815), .ZN(n10059) );
  NAND2_X2 U12733 ( .A1(n12426), .A2(n14841), .ZN(n12428) );
  OAI21_X1 U12734 ( .B1(n12426), .B2(n10060), .A(n10059), .ZN(n12913) );
  NAND3_X1 U12735 ( .A1(n9779), .A2(n12991), .A3(n10064), .ZN(n13190) );
  NAND3_X1 U12736 ( .A1(n10068), .A2(n12992), .A3(n10067), .ZN(n10066) );
  NOR3_X2 U12737 ( .A1(n17847), .A2(n18197), .A3(n17858), .ZN(n17842) );
  NAND2_X2 U12738 ( .A1(n17936), .A2(n17968), .ZN(n17897) );
  OR2_X2 U12739 ( .A1(n18068), .A2(n18400), .ZN(n10072) );
  AND2_X2 U12740 ( .A1(n18022), .A2(n10073), .ZN(n17969) );
  NAND4_X1 U12741 ( .A1(n19146), .A2(n19130), .A3(n19139), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15864) );
  AND2_X1 U12742 ( .A1(n12227), .A2(n12226), .ZN(n10075) );
  AND2_X2 U12743 ( .A1(n12165), .A2(n12189), .ZN(n12175) );
  AND2_X2 U12744 ( .A1(n12161), .A2(n12167), .ZN(n12165) );
  OR2_X2 U12745 ( .A1(n12166), .A2(n10076), .ZN(n12161) );
  INV_X1 U12746 ( .A(n10077), .ZN(n15142) );
  NAND3_X1 U12747 ( .A1(n10369), .A2(n10370), .A3(n10367), .ZN(n10080) );
  NAND2_X1 U12748 ( .A1(n11962), .A2(n11951), .ZN(n10082) );
  NAND2_X1 U12749 ( .A1(n10082), .A2(n10081), .ZN(n19369) );
  AND3_X2 U12750 ( .A1(n10085), .A2(n10084), .A3(n10083), .ZN(n15388) );
  OR2_X1 U12751 ( .A1(n15599), .A2(n15597), .ZN(n15416) );
  NAND2_X1 U12752 ( .A1(n12033), .A2(n12032), .ZN(n10091) );
  INV_X1 U12753 ( .A(n10091), .ZN(n10089) );
  NAND3_X1 U12754 ( .A1(n10088), .A2(n10086), .A3(n15209), .ZN(n12122) );
  NAND3_X1 U12755 ( .A1(n10087), .A2(n10091), .A3(n12101), .ZN(n10086) );
  NAND3_X1 U12756 ( .A1(n10089), .A2(n10090), .A3(n12101), .ZN(n10088) );
  AND2_X1 U12757 ( .A1(n15277), .A2(n15266), .ZN(n15259) );
  NAND3_X1 U12758 ( .A1(n10857), .A2(n12105), .A3(n10856), .ZN(n12107) );
  NAND2_X1 U12759 ( .A1(n14294), .A2(n9816), .ZN(n15285) );
  AND2_X1 U12760 ( .A1(n12200), .A2(n10115), .ZN(n12197) );
  NAND2_X1 U12761 ( .A1(n12200), .A2(n9745), .ZN(n12192) );
  NAND2_X1 U12762 ( .A1(n12200), .A2(n10117), .ZN(n12180) );
  NAND2_X1 U12763 ( .A1(n12200), .A2(n10877), .ZN(n12185) );
  AND2_X2 U12764 ( .A1(n14664), .A2(n9817), .ZN(n14627) );
  NOR2_X2 U12765 ( .A1(n14437), .A2(n10133), .ZN(n14676) );
  INV_X1 U12766 ( .A(n10137), .ZN(n14675) );
  AOI21_X1 U12767 ( .B1(n10141), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n10142), .ZN(n10140) );
  INV_X1 U12768 ( .A(n15764), .ZN(n10141) );
  NAND2_X2 U12769 ( .A1(n15533), .A2(n12314), .ZN(n15742) );
  NAND2_X1 U12770 ( .A1(n12035), .A2(n10146), .ZN(n12092) );
  AND2_X2 U12771 ( .A1(n15443), .A2(n10147), .ZN(n15409) );
  NAND3_X1 U12772 ( .A1(n12573), .A2(n12572), .A3(n12571), .ZN(n10152) );
  OR2_X1 U12773 ( .A1(n10152), .A2(n10151), .ZN(n13951) );
  NAND2_X1 U12774 ( .A1(n13950), .A2(n13949), .ZN(n10151) );
  NAND2_X1 U12775 ( .A1(n14299), .A2(n14301), .ZN(n14300) );
  INV_X1 U12776 ( .A(n14301), .ZN(n10156) );
  NAND2_X1 U12777 ( .A1(n10157), .A2(n15249), .ZN(n15243) );
  NAND2_X1 U12778 ( .A1(n10158), .A2(n15247), .ZN(n10157) );
  AOI21_X1 U12779 ( .B1(n12536), .B2(n19507), .A(n12326), .ZN(n12327) );
  NAND2_X1 U12780 ( .A1(n15460), .A2(n15459), .ZN(n15527) );
  INV_X1 U12781 ( .A(n12912), .ZN(n14561) );
  NAND2_X1 U12782 ( .A1(n12912), .A2(n11783), .ZN(n11905) );
  XNOR2_X1 U12784 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11735) );
  AND2_X2 U12785 ( .A1(n11133), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14064) );
  NAND2_X1 U12786 ( .A1(n15419), .A2(n15393), .ZN(n15387) );
  AND2_X2 U12787 ( .A1(n11987), .A2(n19559), .ZN(n11988) );
  NAND2_X1 U12788 ( .A1(n14627), .A2(n14629), .ZN(n14612) );
  AND2_X1 U12789 ( .A1(n9714), .A2(n11978), .ZN(n11980) );
  OAI22_X1 U12790 ( .A1(n10585), .A2(n10569), .B1(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n20163), .ZN(n10583) );
  AND2_X1 U12791 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20163), .ZN(
        n10569) );
  INV_X1 U12792 ( .A(n13789), .ZN(n11262) );
  NOR2_X1 U12793 ( .A1(n11954), .A2(n11953), .ZN(n11955) );
  NAND2_X1 U12794 ( .A1(n11954), .A2(n11953), .ZN(n11952) );
  AND2_X1 U12795 ( .A1(n11906), .A2(n13992), .ZN(n15977) );
  NAND2_X1 U12796 ( .A1(n12339), .A2(n13992), .ZN(n12346) );
  NAND2_X1 U12797 ( .A1(n9710), .A2(n13992), .ZN(n12400) );
  INV_X1 U12798 ( .A(n9710), .ZN(n11743) );
  NOR2_X1 U12799 ( .A1(n9692), .A2(n20222), .ZN(n11713) );
  NOR2_X1 U12800 ( .A1(n15703), .A2(n16429), .ZN(n10165) );
  INV_X1 U12801 ( .A(n13794), .ZN(n14097) );
  INV_X1 U12802 ( .A(n12329), .ZN(n13794) );
  AND2_X1 U12803 ( .A1(n11538), .A2(n11537), .ZN(n10166) );
  INV_X1 U12804 ( .A(n14653), .ZN(n14712) );
  INV_X1 U12805 ( .A(n11177), .ZN(n13980) );
  OR2_X1 U12806 ( .A1(n12306), .A2(n12305), .ZN(n10167) );
  INV_X1 U12807 ( .A(n12865), .ZN(n10678) );
  OR2_X1 U12808 ( .A1(n9756), .A2(n17418), .ZN(n10169) );
  OR2_X1 U12809 ( .A1(n12959), .A2(n17447), .ZN(n10170) );
  AND2_X1 U12810 ( .A1(n18057), .A2(n15963), .ZN(n10171) );
  OR2_X1 U12811 ( .A1(n12888), .A2(n12262), .ZN(n10172) );
  NAND2_X1 U12812 ( .A1(n15274), .A2(n12756), .ZN(n12778) );
  INV_X1 U12813 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11332) );
  OR2_X1 U12814 ( .A1(n13269), .A2(n12030), .ZN(n19510) );
  AND3_X1 U12815 ( .A1(n10604), .A2(n10283), .A3(n10603), .ZN(n10173) );
  AND3_X1 U12816 ( .A1(n10593), .A2(n10592), .A3(n10283), .ZN(n10174) );
  NOR2_X1 U12817 ( .A1(n9716), .A2(n14198), .ZN(n10175) );
  OR2_X1 U12818 ( .A1(n12004), .A2(n12003), .ZN(n10176) );
  AND2_X1 U12819 ( .A1(n11006), .A2(n13384), .ZN(n10177) );
  AND3_X1 U12820 ( .A1(n12191), .A2(n15463), .A3(n15700), .ZN(n10178) );
  NOR2_X1 U12821 ( .A1(n20662), .A2(n20661), .ZN(n10179) );
  OR2_X1 U12822 ( .A1(n20324), .A2(n14558), .ZN(n10180) );
  INV_X1 U12823 ( .A(n14742), .ZN(n11783) );
  AND2_X1 U12824 ( .A1(n10676), .A2(n10675), .ZN(n10181) );
  INV_X1 U12825 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13040) );
  INV_X1 U12826 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n13985) );
  AND2_X1 U12827 ( .A1(n12180), .A2(n12177), .ZN(n10182) );
  INV_X1 U12828 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12246) );
  AND2_X1 U12829 ( .A1(n10242), .A2(n10241), .ZN(n10183) );
  AND2_X1 U12830 ( .A1(n17533), .A2(n17578), .ZN(n17530) );
  INV_X2 U12831 ( .A(n17530), .ZN(n17525) );
  INV_X1 U12832 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10192) );
  AND3_X1 U12833 ( .A1(n10589), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10588), .ZN(n10184) );
  AND2_X1 U12834 ( .A1(n11628), .A2(n11627), .ZN(n10185) );
  INV_X1 U12835 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13031) );
  INV_X1 U12836 ( .A(n10274), .ZN(n10373) );
  AND2_X1 U12837 ( .A1(n15725), .A2(n15726), .ZN(n10186) );
  INV_X1 U12838 ( .A(n12730), .ZN(n12704) );
  INV_X1 U12839 ( .A(n12101), .ZN(n12162) );
  INV_X1 U12840 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20806) );
  NAND2_X1 U12841 ( .A1(n17987), .A2(n18147), .ZN(n17899) );
  OR2_X1 U12842 ( .A1(n15362), .A2(n14421), .ZN(n10187) );
  INV_X1 U12843 ( .A(n20071), .ZN(n19342) );
  AND3_X1 U12844 ( .A1(n13228), .A2(n13227), .A3(n13226), .ZN(n10188) );
  AND4_X1 U12845 ( .A1(n10942), .A2(n10941), .A3(n10940), .A4(n10939), .ZN(
        n10189) );
  AND2_X2 U12846 ( .A1(n14065), .A2(n13508), .ZN(n11406) );
  AND2_X1 U12847 ( .A1(n11033), .A2(n10999), .ZN(n10190) );
  INV_X1 U12848 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11726) );
  OR3_X1 U12849 ( .A1(n11759), .A2(n11758), .A3(n11907), .ZN(n11760) );
  NOR2_X1 U12850 ( .A1(n11122), .A2(n11121), .ZN(n11123) );
  INV_X1 U12851 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10259) );
  NAND2_X1 U12852 ( .A1(n9720), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10856) );
  NAND2_X1 U12853 ( .A1(n10655), .A2(n12465), .ZN(n10679) );
  AOI22_X1 U12854 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10592) );
  AND2_X1 U12855 ( .A1(n11766), .A2(n11765), .ZN(n11910) );
  OR2_X1 U12856 ( .A1(n11248), .A2(n11247), .ZN(n12382) );
  NAND2_X1 U12857 ( .A1(n11003), .A2(n10191), .ZN(n11004) );
  AND3_X1 U12858 ( .A1(n11108), .A2(n11107), .A3(n11106), .ZN(n11120) );
  INV_X1 U12859 ( .A(n10679), .ZN(n10651) );
  NAND2_X1 U12860 ( .A1(n10622), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10254) );
  INV_X1 U12861 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n11733) );
  INV_X1 U12862 ( .A(n11045), .ZN(n11046) );
  INV_X1 U12863 ( .A(n14678), .ZN(n11466) );
  AND2_X1 U12864 ( .A1(n11250), .A2(n11249), .ZN(n11251) );
  OR2_X1 U12865 ( .A1(n11105), .A2(n11104), .ZN(n12340) );
  NAND2_X1 U12866 ( .A1(n15974), .A2(n13812), .ZN(n11008) );
  AND2_X1 U12867 ( .A1(n10571), .A2(n10570), .ZN(n10580) );
  CLKBUF_X3 U12868 ( .A(n10623), .Z(n12830) );
  NOR2_X1 U12869 ( .A1(n12030), .A2(n20201), .ZN(n12550) );
  INV_X1 U12870 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12245) );
  INV_X1 U12871 ( .A(n16464), .ZN(n12163) );
  AND4_X1 U12872 ( .A1(n10304), .A2(n10303), .A3(n10302), .A4(n10301), .ZN(
        n10310) );
  AOI21_X1 U12873 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n19001), .A(
        n13065), .ZN(n13066) );
  NOR2_X1 U12874 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n11733), .ZN(
        n11765) );
  OR2_X1 U12875 ( .A1(n11723), .A2(n11722), .ZN(n13608) );
  INV_X1 U12876 ( .A(n11604), .ZN(n11605) );
  AND2_X1 U12877 ( .A1(n14439), .A2(n14435), .ZN(n11404) );
  NOR2_X1 U12878 ( .A1(n13384), .A2(n20806), .ZN(n11173) );
  INV_X1 U12879 ( .A(n14106), .ZN(n11293) );
  INV_X1 U12880 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11207) );
  OR2_X1 U12881 ( .A1(n11083), .A2(n11082), .ZN(n12341) );
  INV_X1 U12882 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11729) );
  INV_X1 U12883 ( .A(n11162), .ZN(n11164) );
  INV_X1 U12884 ( .A(n10580), .ZN(n10573) );
  INV_X1 U12885 ( .A(n12127), .ZN(n10871) );
  AND2_X1 U12886 ( .A1(n14143), .A2(n14141), .ZN(n12579) );
  INV_X1 U12887 ( .A(n19404), .ZN(n12576) );
  NAND2_X1 U12888 ( .A1(n12246), .A2(n12245), .ZN(n12247) );
  OR2_X1 U12889 ( .A1(n12101), .A2(n19289), .ZN(n12206) );
  INV_X1 U12890 ( .A(n19565), .ZN(n12492) );
  NAND3_X1 U12891 ( .A1(n9713), .A2(n11990), .A3(n13472), .ZN(n12079) );
  AOI21_X1 U12892 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18996), .A(
        n13064), .ZN(n13069) );
  INV_X1 U12893 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17452) );
  NAND2_X1 U12894 ( .A1(n18057), .A2(n18285), .ZN(n13050) );
  INV_X1 U12895 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13137) );
  INV_X1 U12896 ( .A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17316) );
  AND2_X1 U12897 ( .A1(n18503), .A2(n13165), .ZN(n13161) );
  AOI21_X1 U12898 ( .B1(n11766), .B2(n11734), .A(n11765), .ZN(n11912) );
  OR2_X1 U12899 ( .A1(n16285), .A2(n13982), .ZN(n13983) );
  OR2_X1 U12900 ( .A1(n14059), .A2(n11021), .ZN(n11022) );
  NOR2_X1 U12901 ( .A1(n12439), .A2(n12910), .ZN(n12440) );
  OR2_X1 U12902 ( .A1(n14834), .A2(n11177), .ZN(n11652) );
  AND2_X1 U12903 ( .A1(n11569), .A2(n11568), .ZN(n14643) );
  NAND2_X1 U12904 ( .A1(n11356), .A2(n11355), .ZN(n11357) );
  NAND2_X1 U12905 ( .A1(n13522), .A2(n11791), .ZN(n11915) );
  NAND2_X1 U12906 ( .A1(n11189), .A2(n11188), .ZN(n13905) );
  OAI211_X1 U12907 ( .C1(n11762), .C2(n20376), .A(n11089), .B(n11088), .ZN(
        n11170) );
  NAND2_X1 U12908 ( .A1(n14132), .A2(n20222), .ZN(n11203) );
  NAND2_X1 U12909 ( .A1(n10885), .A2(n10650), .ZN(n12494) );
  AND2_X1 U12910 ( .A1(n10558), .A2(n10557), .ZN(n15332) );
  INV_X1 U12911 ( .A(n16427), .ZN(n15459) );
  AND2_X1 U12912 ( .A1(n10556), .A2(n10555), .ZN(n15612) );
  NOR2_X1 U12913 ( .A1(n15366), .A2(n15176), .ZN(n15157) );
  INV_X1 U12914 ( .A(n15732), .ZN(n10780) );
  NAND3_X1 U12916 ( .A1(n15817), .A2(n11978), .A3(n19541), .ZN(n13744) );
  AOI22_X1 U12917 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n18996), .B2(n19146), .ZN(
        n13185) );
  AND2_X1 U12918 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12954) );
  INV_X1 U12919 ( .A(n13021), .ZN(n13022) );
  INV_X1 U12920 ( .A(n18256), .ZN(n15959) );
  NOR2_X1 U12921 ( .A1(n13206), .A2(n18091), .ZN(n13208) );
  NOR2_X1 U12922 ( .A1(n18533), .A2(n17689), .ZN(n13168) );
  NOR2_X1 U12923 ( .A1(n18533), .A2(n18509), .ZN(n13175) );
  INV_X1 U12924 ( .A(n11516), .ZN(n11517) );
  INV_X1 U12925 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14690) );
  INV_X1 U12926 ( .A(n20306), .ZN(n20254) );
  NOR2_X1 U12927 ( .A1(n13990), .A2(n13989), .ZN(n14000) );
  INV_X1 U12928 ( .A(n12433), .ZN(n12434) );
  NAND2_X1 U12929 ( .A1(n11565), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11604) );
  OR2_X1 U12930 ( .A1(n11437), .A2(n14690), .ZN(n11452) );
  NOR2_X1 U12931 ( .A1(n11399), .A2(n16099), .ZN(n11374) );
  NOR2_X1 U12932 ( .A1(n11333), .A2(n11332), .ZN(n11337) );
  OAI211_X1 U12933 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n13985), .A(n20888), 
        .B(n20804), .ZN(n13801) );
  OR2_X1 U12934 ( .A1(n13530), .A2(n13529), .ZN(n15979) );
  INV_X1 U12936 ( .A(n20732), .ZN(n13883) );
  AND2_X1 U12937 ( .A1(n14246), .A2(n14245), .ZN(n15127) );
  INV_X1 U12938 ( .A(n14237), .ZN(n14198) );
  INV_X1 U12939 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n10997) );
  INV_X1 U12940 ( .A(n10893), .ZN(n10894) );
  OR2_X1 U12941 ( .A1(n12099), .A2(n9720), .ZN(n12235) );
  OR2_X1 U12942 ( .A1(n19366), .A2(n19920), .ZN(n19391) );
  INV_X1 U12943 ( .A(n15272), .ZN(n12752) );
  AND3_X1 U12944 ( .A1(n10478), .A2(n10477), .A3(n10476), .ZN(n13237) );
  OAI21_X1 U12945 ( .B1(n12875), .B2(n12874), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n15293) );
  OR2_X1 U12946 ( .A1(n15394), .A2(n15393), .ZN(n15395) );
  AND3_X1 U12947 ( .A1(n10503), .A2(n10502), .A3(n10501), .ZN(n16533) );
  NAND2_X1 U12948 ( .A1(n12312), .A2(n12311), .ZN(n12314) );
  INV_X1 U12949 ( .A(n19517), .ZN(n19350) );
  INV_X1 U12950 ( .A(n12264), .ZN(n16616) );
  INV_X1 U12951 ( .A(n15796), .ZN(n20158) );
  NAND2_X1 U12952 ( .A1(n15819), .A2(n20177), .ZN(n19727) );
  NAND2_X1 U12953 ( .A1(n15796), .A2(n20169), .ZN(n19760) );
  NAND2_X1 U12954 ( .A1(n20158), .A2(n20169), .ZN(n19643) );
  INV_X1 U12955 ( .A(n20157), .ZN(n20150) );
  NOR2_X1 U12956 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17046), .ZN(n17027) );
  NAND2_X1 U12957 ( .A1(n19186), .A2(n17689), .ZN(n13256) );
  INV_X1 U12958 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17447) );
  INV_X1 U12959 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17372) );
  INV_X1 U12960 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17418) );
  INV_X1 U12961 ( .A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17402) );
  OR2_X1 U12962 ( .A1(n12955), .A2(n12954), .ZN(n12969) );
  OR2_X1 U12963 ( .A1(n16685), .A2(n18152), .ZN(n13228) );
  NOR2_X1 U12964 ( .A1(n18000), .A2(n17991), .ZN(n17984) );
  INV_X1 U12965 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18049) );
  NOR2_X1 U12966 ( .A1(n17840), .A2(n15963), .ZN(n18155) );
  NOR2_X1 U12967 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n13014), .ZN(
        n17886) );
  NOR2_X1 U12968 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18057), .ZN(
        n17927) );
  OR2_X1 U12969 ( .A1(n17997), .A2(n17956), .ZN(n18290) );
  INV_X1 U12970 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18370) );
  INV_X1 U12971 ( .A(n18964), .ZN(n18983) );
  INV_X1 U12972 ( .A(n18668), .ZN(n18669) );
  INV_X1 U12973 ( .A(n17987), .ZN(n18148) );
  NAND2_X1 U12974 ( .A1(n11777), .A2(n11776), .ZN(n13597) );
  INV_X1 U12975 ( .A(n20219), .ZN(n13601) );
  NAND2_X1 U12976 ( .A1(n11518), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11564) );
  AND2_X1 U12977 ( .A1(n16082), .A2(n13986), .ZN(n20268) );
  NOR2_X1 U12978 ( .A1(n20301), .A2(n20223), .ZN(n20288) );
  INV_X1 U12979 ( .A(n20324), .ZN(n14740) );
  INV_X1 U12980 ( .A(n11936), .ZN(n11937) );
  OR2_X1 U12981 ( .A1(n11919), .A2(n13987), .ZN(n11920) );
  INV_X1 U12982 ( .A(n13800), .ZN(n13799) );
  NAND2_X1 U12983 ( .A1(n11482), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11516) );
  NAND2_X1 U12984 ( .A1(n11338), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11399) );
  AND3_X1 U12985 ( .A1(n13523), .A2(n12431), .A3(n13597), .ZN(n16183) );
  OR2_X1 U12986 ( .A1(n15027), .A2(n16209), .ZN(n14968) );
  AND2_X1 U12987 ( .A1(n14968), .A2(n14967), .ZN(n15007) );
  OR3_X1 U12988 ( .A1(n15031), .A2(n14966), .A3(n14965), .ZN(n15027) );
  INV_X1 U12989 ( .A(n16270), .ZN(n16209) );
  AND2_X1 U12990 ( .A1(n13623), .A2(n15977), .ZN(n14963) );
  INV_X2 U12991 ( .A(n16238), .ZN(n16285) );
  AND2_X1 U12992 ( .A1(n13623), .A2(n13621), .ZN(n16286) );
  NAND2_X1 U12993 ( .A1(n20222), .A2(n13801), .ZN(n14089) );
  NAND2_X1 U12994 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n13597), .ZN(n20888) );
  AND2_X1 U12995 ( .A1(n20413), .A2(n10175), .ZN(n20409) );
  OAI22_X1 U12996 ( .A1(n20420), .A2(n20419), .B1(n20621), .B2(n20518), .ZN(
        n20444) );
  OAI21_X1 U12997 ( .B1(n14203), .B2(n20491), .A(n20516), .ZN(n20492) );
  INV_X1 U12998 ( .A(n14199), .ZN(n20508) );
  INV_X1 U12999 ( .A(n20571), .ZN(n20561) );
  OAI211_X1 U13000 ( .C1(n20594), .C2(n20700), .A(n20579), .B(n20619), .ZN(
        n20596) );
  AND2_X1 U13001 ( .A1(n20671), .A2(n10175), .ZN(n20606) );
  INV_X1 U13003 ( .A(n20737), .ZN(n20695) );
  OAI22_X1 U13004 ( .A1(n20708), .A2(n20707), .B1(n20706), .B2(n20705), .ZN(
        n20733) );
  AND2_X1 U13005 ( .A1(n20747), .A2(n10175), .ZN(n20732) );
  OAI21_X1 U13006 ( .B1(n20700), .B2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n14311), .ZN(n20545) );
  AND2_X1 U13007 ( .A1(n20747), .A2(n21122), .ZN(n15130) );
  OAI211_X1 U13008 ( .C1(n15128), .C2(n14241), .A(n20516), .B(n20617), .ZN(
        n15126) );
  NOR2_X1 U13009 ( .A1(n13827), .A2(n14537), .ZN(n20794) );
  INV_X1 U13010 ( .A(n20872), .ZN(n20852) );
  AND2_X1 U13011 ( .A1(n20875), .A2(n10997), .ZN(n20849) );
  INV_X1 U13012 ( .A(n16639), .ZN(n13350) );
  OAI21_X1 U13013 ( .B1(n12261), .B2(n19362), .A(n10894), .ZN(n10895) );
  INV_X1 U13014 ( .A(n19362), .ZN(n19385) );
  INV_X1 U13015 ( .A(n19517), .ZN(n19324) );
  INV_X1 U13016 ( .A(n19381), .ZN(n19305) );
  AND2_X1 U13017 ( .A1(n20198), .A2(n10850), .ZN(n19389) );
  OR2_X1 U13018 ( .A1(n10449), .A2(n10448), .ZN(n13691) );
  INV_X1 U13019 ( .A(n15369), .ZN(n16412) );
  NOR2_X1 U13020 ( .A1(n14398), .A2(n14399), .ZN(n14423) );
  AND2_X1 U13021 ( .A1(n19428), .A2(n13426), .ZN(n19434) );
  INV_X1 U13022 ( .A(n13277), .ZN(n19482) );
  INV_X1 U13023 ( .A(n19510), .ZN(n12279) );
  INV_X1 U13024 ( .A(n15683), .ZN(n19400) );
  AND2_X1 U13025 ( .A1(n15735), .A2(n15734), .ZN(n19407) );
  AND2_X1 U13026 ( .A1(n14492), .A2(n19370), .ZN(n19523) );
  NAND2_X1 U13027 ( .A1(n15571), .A2(n15395), .ZN(n15398) );
  OR2_X1 U13028 ( .A1(n15722), .A2(n15631), .ZN(n16524) );
  AND2_X1 U13029 ( .A1(n14147), .A2(n14146), .ZN(n19294) );
  INV_X1 U13030 ( .A(n19556), .ZN(n16577) );
  AND2_X1 U13031 ( .A1(n12538), .A2(n20187), .ZN(n19551) );
  NOR2_X2 U13032 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20157) );
  OAI21_X1 U13033 ( .B1(n14194), .B2(n14193), .A(n14192), .ZN(n19589) );
  NOR2_X2 U13034 ( .A1(n19820), .A2(n19727), .ZN(n19619) );
  INV_X1 U13035 ( .A(n19623), .ZN(n19639) );
  NOR2_X1 U13036 ( .A1(n19727), .A2(n19643), .ZN(n19668) );
  NOR2_X1 U13037 ( .A1(n19727), .A2(n19696), .ZN(n19713) );
  NOR2_X1 U13038 ( .A1(n19760), .A2(n19727), .ZN(n19782) );
  OAI21_X1 U13039 ( .B1(n19796), .B2(n19795), .A(n19794), .ZN(n19814) );
  NAND2_X1 U13040 ( .A1(n20154), .A2(n20177), .ZN(n19786) );
  OAI21_X1 U13041 ( .B1(n19942), .B2(n19920), .A(n19919), .ZN(n19944) );
  NOR2_X2 U13042 ( .A1(n13753), .A2(n13752), .ZN(n19588) );
  INV_X1 U13043 ( .A(n15825), .ZN(n19985) );
  INV_X1 U13044 ( .A(n19831), .ZN(n20005) );
  INV_X1 U13045 ( .A(n19932), .ZN(n20026) );
  INV_X1 U13046 ( .A(n19941), .ZN(n20045) );
  AND2_X1 U13047 ( .A1(n20173), .A2(n12275), .ZN(n16628) );
  NAND2_X1 U13048 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20174) );
  AND3_X1 U13049 ( .A1(n20074), .A2(n20132), .A3(n20083), .ZN(n20208) );
  NOR2_X1 U13050 ( .A1(n17689), .A2(n18498), .ZN(n13162) );
  NOR2_X1 U13051 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16927), .ZN(n16916) );
  NOR2_X1 U13052 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16947), .ZN(n16933) );
  NOR2_X1 U13053 ( .A1(n16994), .A2(P3_EBX_REG_17__SCAN_IN), .ZN(n16993) );
  NOR2_X1 U13054 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17070), .ZN(n17053) );
  NOR2_X1 U13055 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17076), .ZN(n17075) );
  NOR2_X1 U13056 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17142), .ZN(n17120) );
  INV_X1 U13057 ( .A(n17159), .ZN(n17183) );
  INV_X1 U13058 ( .A(n17155), .ZN(n17187) );
  NOR2_X1 U13059 ( .A1(n16948), .A2(n17298), .ZN(n17270) );
  INV_X1 U13060 ( .A(n18533), .ZN(n17578) );
  INV_X1 U13061 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17513) );
  NOR2_X1 U13062 ( .A1(n17735), .A2(n17605), .ZN(n17600) );
  AOI21_X1 U13063 ( .B1(n15934), .B2(n19014), .A(n19038), .ZN(n17688) );
  NOR2_X1 U13064 ( .A1(n15962), .A2(n17872), .ZN(n17834) );
  INV_X1 U13065 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18269) );
  INV_X1 U13066 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17997) );
  INV_X1 U13067 ( .A(n18375), .ZN(n18369) );
  INV_X1 U13068 ( .A(n18471), .ZN(n18460) );
  NOR2_X1 U13069 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19125), .ZN(
        n19147) );
  CLKBUF_X1 U13070 ( .A(n18581), .Z(n18594) );
  INV_X1 U13071 ( .A(n18638), .ZN(n18640) );
  INV_X1 U13072 ( .A(n18906), .ZN(n18803) );
  INV_X1 U13073 ( .A(n18842), .ZN(n18849) );
  CLKBUF_X1 U13074 ( .A(n18884), .Z(n18877) );
  AND2_X1 U13075 ( .A1(n18891), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18922) );
  INV_X1 U13076 ( .A(n18880), .ZN(n18935) );
  NOR2_X1 U13077 ( .A1(n19025), .A2(n19183), .ZN(n19169) );
  INV_X1 U13078 ( .A(n13751), .ZN(n13753) );
  NAND2_X1 U13079 ( .A1(n13357), .A2(n13459), .ZN(n20904) );
  INV_X1 U13080 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21095) );
  INV_X1 U13081 ( .A(n20303), .ZN(n20274) );
  INV_X1 U13082 ( .A(n20304), .ZN(n20289) );
  OR2_X1 U13083 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16304), .ZN(n20327) );
  INV_X1 U13084 ( .A(n20328), .ZN(n20356) );
  OR2_X1 U13085 ( .A1(n20368), .A2(n13992), .ZN(n13650) );
  INV_X1 U13086 ( .A(n16183), .ZN(n20226) );
  NAND2_X1 U13087 ( .A1(n13623), .A2(n13605), .ZN(n16222) );
  AOI211_X2 U13088 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n14317), .A(n14315), 
        .B(n14314), .ZN(n20397) );
  NAND2_X1 U13089 ( .A1(n20413), .A2(n21122), .ZN(n20442) );
  NAND2_X1 U13090 ( .A1(n20413), .A2(n20610), .ZN(n20479) );
  NAND2_X1 U13091 ( .A1(n20413), .A2(n20670), .ZN(n20495) );
  NAND2_X1 U13092 ( .A1(n20549), .A2(n21122), .ZN(n20531) );
  NAND2_X1 U13093 ( .A1(n20549), .A2(n20610), .ZN(n20571) );
  NAND2_X1 U13094 ( .A1(n20549), .A2(n20670), .ZN(n20599) );
  NAND2_X1 U13095 ( .A1(n20671), .A2(n21122), .ZN(n20655) );
  NAND2_X1 U13096 ( .A1(n20671), .A2(n20610), .ZN(n20684) );
  INV_X1 U13097 ( .A(n20775), .ZN(n20724) );
  AOI21_X1 U13098 ( .B1(n15114), .B2(n20694), .A(n20545), .ZN(n13887) );
  INV_X1 U13099 ( .A(n20497), .ZN(n20766) );
  INV_X1 U13100 ( .A(n20788), .ZN(n20802) );
  NOR2_X1 U13101 ( .A1(n20875), .A2(n20817), .ZN(n20884) );
  INV_X1 U13102 ( .A(n20852), .ZN(n20868) );
  INV_X1 U13103 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20074) );
  INV_X1 U13104 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19595) );
  AOI21_X1 U13105 ( .B1(n10896), .B2(n19389), .A(n10895), .ZN(n10897) );
  NAND2_X1 U13106 ( .A1(n20198), .A2(n10886), .ZN(n19362) );
  XNOR2_X1 U13107 ( .A(n13413), .B(n13412), .ZN(n20166) );
  NAND2_X1 U13108 ( .A1(n19428), .A2(n12865), .ZN(n15373) );
  NAND2_X1 U13109 ( .A1(n19477), .A2(n20195), .ZN(n19445) );
  OR2_X1 U13110 ( .A1(n19477), .A2(n13393), .ZN(n19439) );
  NAND2_X1 U13111 ( .A1(n13392), .A2(n20208), .ZN(n19477) );
  NAND2_X1 U13112 ( .A1(n13275), .A2(n12030), .ZN(n13389) );
  INV_X1 U13113 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16425) );
  INV_X1 U13114 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19279) );
  INV_X1 U13115 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16457) );
  INV_X1 U13116 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16486) );
  INV_X1 U13117 ( .A(n16494), .ZN(n19501) );
  INV_X1 U13118 ( .A(n19551), .ZN(n16589) );
  INV_X1 U13119 ( .A(n19549), .ZN(n16593) );
  AOI211_X2 U13120 ( .C1(n14188), .C2(n14193), .A(n14187), .B(n19915), .ZN(
        n19593) );
  NAND2_X1 U13121 ( .A1(n19596), .A2(n19753), .ZN(n19623) );
  INV_X1 U13122 ( .A(n19668), .ZN(n19664) );
  INV_X1 U13123 ( .A(n19691), .ZN(n19686) );
  INV_X1 U13124 ( .A(n19713), .ZN(n19724) );
  INV_X1 U13125 ( .A(n19782), .ZN(n19780) );
  OR2_X1 U13126 ( .A1(n19820), .A2(n19786), .ZN(n19844) );
  INV_X1 U13127 ( .A(n19904), .ZN(n19881) );
  INV_X1 U13128 ( .A(n19914), .ZN(n19947) );
  AOI211_X2 U13129 ( .C1(n13836), .C2(n13835), .A(n19915), .B(n13834), .ZN(
        n19970) );
  AOI211_X2 U13130 ( .C1(n14159), .C2(n14166), .A(n14158), .B(n19915), .ZN(
        n19990) );
  NOR2_X1 U13131 ( .A1(n19997), .A2(n19996), .ZN(n20059) );
  NOR2_X1 U13132 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16633) );
  INV_X1 U13133 ( .A(n20146), .ZN(n20073) );
  CLKBUF_X1 U13134 ( .A(n20136), .Z(n20131) );
  INV_X2 U13135 ( .A(n20213), .ZN(n20216) );
  INV_X1 U13136 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16812) );
  INV_X1 U13137 ( .A(n13258), .ZN(n17136) );
  NAND2_X1 U13138 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17196), .ZN(n17159) );
  INV_X1 U13139 ( .A(n17193), .ZN(n17192) );
  NOR2_X1 U13140 ( .A1(n16908), .A2(n17253), .ZN(n17258) );
  INV_X1 U13141 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17389) );
  INV_X1 U13142 ( .A(n17520), .ZN(n17533) );
  INV_X1 U13143 ( .A(n16687), .ZN(n17656) );
  NAND2_X1 U13144 ( .A1(n17690), .A2(n17689), .ZN(n17707) );
  NAND2_X1 U13145 ( .A1(n17728), .A2(n17688), .ZN(n17726) );
  INV_X1 U13146 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18021) );
  INV_X1 U13147 ( .A(n18139), .ZN(n18130) );
  INV_X1 U13148 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18143) );
  OR3_X1 U13149 ( .A1(n16699), .A2(n18380), .A3(n17807), .ZN(n16700) );
  INV_X1 U13150 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18285) );
  INV_X1 U13151 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18302) );
  INV_X1 U13152 ( .A(n18391), .ZN(n18380) );
  AND2_X1 U13153 ( .A1(n17197), .A2(n16810), .ZN(n19168) );
  INV_X1 U13154 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18523) );
  INV_X1 U13155 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18537) );
  INV_X1 U13156 ( .A(n18616), .ZN(n18615) );
  INV_X1 U13157 ( .A(n18707), .ZN(n18694) );
  INV_X1 U13158 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18722) );
  INV_X1 U13159 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18733) );
  INV_X1 U13160 ( .A(n18766), .ZN(n18761) );
  INV_X1 U13161 ( .A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18802) );
  INV_X1 U13162 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18825) );
  INV_X1 U13163 ( .A(n18909), .ZN(n18836) );
  INV_X1 U13164 ( .A(n18945), .ZN(n18888) );
  INV_X1 U13165 ( .A(n18869), .ZN(n18925) );
  INV_X1 U13166 ( .A(n18876), .ZN(n18941) );
  INV_X1 U13167 ( .A(n19122), .ZN(n19119) );
  INV_X1 U13168 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19045) );
  NOR2_X1 U13169 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13234), .ZN(n16797)
         );
  INV_X1 U13170 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20093) );
  OR4_X1 U13171 ( .A1(n13249), .A2(n13248), .A3(n13247), .A4(n13246), .ZN(
        P2_U2844) );
  INV_X1 U13172 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10193) );
  INV_X1 U13173 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15437) );
  INV_X1 U13174 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n19230) );
  INV_X1 U13175 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16473) );
  INV_X1 U13176 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16492) );
  INV_X1 U13177 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16507) );
  NAND2_X1 U13178 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n10201), .ZN(
        n10200) );
  NAND2_X1 U13179 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n10207), .ZN(
        n10206) );
  INV_X1 U13180 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10195) );
  INV_X1 U13181 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15379) );
  OAI21_X1 U13182 ( .B1(n10194), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n10218), .ZN(n16333) );
  AOI21_X1 U13183 ( .B1(n10217), .B2(n10195), .A(n10194), .ZN(n15408) );
  INV_X1 U13184 ( .A(n15408), .ZN(n16343) );
  OAI21_X1 U13185 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n10196), .A(
        n10216), .ZN(n16371) );
  AOI21_X1 U13186 ( .B1(n15437), .B2(n10197), .A(n10196), .ZN(n15440) );
  INV_X1 U13187 ( .A(n15440), .ZN(n15137) );
  OAI21_X1 U13188 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n10198), .A(
        n10197), .ZN(n15449) );
  AOI21_X1 U13189 ( .B1(n15171), .B2(n10215), .A(n10198), .ZN(n15471) );
  AOI21_X1 U13190 ( .B1(n10213), .B2(n19230), .A(n9796), .ZN(n19229) );
  AOI21_X1 U13191 ( .B1(n15516), .B2(n10211), .A(n10214), .ZN(n15517) );
  AOI21_X1 U13192 ( .B1(n19279), .B2(n10210), .A(n10212), .ZN(n19277) );
  AOI21_X1 U13193 ( .B1(n16457), .B2(n10208), .A(n9795), .ZN(n19301) );
  AOI21_X1 U13194 ( .B1(n16473), .B2(n10206), .A(n10209), .ZN(n16463) );
  AOI21_X1 U13195 ( .B1(n16486), .B2(n10204), .A(n10207), .ZN(n16479) );
  AOI21_X1 U13196 ( .B1(n16492), .B2(n10202), .A(n10205), .ZN(n19347) );
  AOI21_X1 U13197 ( .B1(n16507), .B2(n10200), .A(n10203), .ZN(n16493) );
  AOI21_X1 U13198 ( .B1(n14035), .B2(n10199), .A(n10201), .ZN(n15206) );
  INV_X1 U13199 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16585) );
  INV_X1 U13200 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19515) );
  AOI22_X1 U13201 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16585), .B1(n19515), 
        .B2(n20201), .ZN(n15774) );
  INV_X1 U13202 ( .A(n15774), .ZN(n19398) );
  INV_X1 U13203 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15229) );
  OAI22_X1 U13204 ( .A1(n20201), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n15229), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15227) );
  AND2_X1 U13205 ( .A1(n19398), .A2(n15227), .ZN(n15219) );
  OAI21_X1 U13206 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n10199), .ZN(n15221) );
  NAND2_X1 U13207 ( .A1(n15219), .A2(n15221), .ZN(n15204) );
  NOR2_X1 U13208 ( .A1(n15206), .A2(n15204), .ZN(n19371) );
  OAI21_X1 U13209 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n10201), .A(
        n10200), .ZN(n19500) );
  NAND2_X1 U13210 ( .A1(n19371), .A2(n19500), .ZN(n15193) );
  NOR2_X1 U13211 ( .A1(n16493), .A2(n15193), .ZN(n14114) );
  OAI21_X1 U13212 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n10203), .A(
        n10202), .ZN(n14346) );
  NAND2_X1 U13213 ( .A1(n14114), .A2(n14346), .ZN(n19346) );
  NOR2_X1 U13214 ( .A1(n19347), .A2(n19346), .ZN(n19338) );
  OAI21_X1 U13215 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n10205), .A(
        n10204), .ZN(n19339) );
  NAND2_X1 U13216 ( .A1(n19338), .A2(n19339), .ZN(n15182) );
  NOR2_X1 U13217 ( .A1(n16479), .A2(n15182), .ZN(n19327) );
  OAI21_X1 U13218 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n10207), .A(
        n10206), .ZN(n19328) );
  NAND2_X1 U13219 ( .A1(n19327), .A2(n19328), .ZN(n13235) );
  NOR2_X1 U13220 ( .A1(n16463), .A2(n13235), .ZN(n19313) );
  OAI21_X1 U13221 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n10209), .A(
        n10208), .ZN(n19314) );
  NAND2_X1 U13222 ( .A1(n19313), .A2(n19314), .ZN(n19298) );
  NOR2_X1 U13223 ( .A1(n19301), .A2(n19298), .ZN(n19291) );
  OAI21_X1 U13224 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n9795), .A(
        n10210), .ZN(n19292) );
  NAND2_X1 U13225 ( .A1(n19291), .A2(n19292), .ZN(n19275) );
  NOR2_X1 U13226 ( .A1(n19277), .A2(n19275), .ZN(n19268) );
  OAI21_X1 U13227 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n10212), .A(
        n10211), .ZN(n19269) );
  NAND2_X1 U13228 ( .A1(n19268), .A2(n19269), .ZN(n19256) );
  NOR2_X1 U13229 ( .A1(n15517), .A2(n19256), .ZN(n19245) );
  OAI21_X1 U13230 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n10214), .A(
        n10213), .ZN(n19246) );
  NAND2_X1 U13231 ( .A1(n19245), .A2(n19246), .ZN(n19227) );
  NOR2_X1 U13232 ( .A1(n19229), .A2(n19227), .ZN(n19223) );
  OAI21_X1 U13233 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n9796), .A(
        n10215), .ZN(n19226) );
  NAND2_X1 U13234 ( .A1(n19223), .A2(n19226), .ZN(n15168) );
  OAI21_X1 U13235 ( .B1(n15471), .B2(n15168), .A(n19299), .ZN(n15153) );
  NAND2_X1 U13236 ( .A1(n15449), .A2(n15153), .ZN(n15152) );
  NAND2_X1 U13237 ( .A1(n19299), .A2(n15152), .ZN(n15136) );
  NAND2_X1 U13238 ( .A1(n15137), .A2(n15136), .ZN(n15135) );
  NAND2_X1 U13239 ( .A1(n19299), .A2(n15135), .ZN(n16370) );
  NAND2_X1 U13240 ( .A1(n16371), .A2(n16370), .ZN(n16369) );
  NAND2_X1 U13241 ( .A1(n19299), .A2(n16369), .ZN(n16362) );
  AOI21_X1 U13242 ( .B1(n16425), .B2(n10216), .A(n9822), .ZN(n16418) );
  INV_X1 U13243 ( .A(n16418), .ZN(n16363) );
  NAND2_X1 U13244 ( .A1(n19299), .A2(n16361), .ZN(n16353) );
  OAI21_X1 U13245 ( .B1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n9822), .A(
        n10217), .ZN(n16354) );
  NAND2_X1 U13246 ( .A1(n19299), .A2(n16352), .ZN(n16342) );
  NAND2_X1 U13247 ( .A1(n16343), .A2(n16342), .ZN(n16341) );
  NAND2_X1 U13248 ( .A1(n13243), .A2(n16341), .ZN(n16332) );
  NAND2_X1 U13249 ( .A1(n16333), .A2(n16332), .ZN(n16331) );
  NAND2_X1 U13250 ( .A1(n19299), .A2(n16331), .ZN(n16318) );
  AOI21_X1 U13251 ( .B1(n15379), .B2(n10218), .A(n10219), .ZN(n15382) );
  INV_X1 U13252 ( .A(n15382), .ZN(n16319) );
  NAND2_X1 U13253 ( .A1(n19299), .A2(n16317), .ZN(n10220) );
  XNOR2_X1 U13254 ( .A(n10219), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12325) );
  NOR3_X1 U13255 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n16033) );
  NAND2_X1 U13256 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n16033), .ZN(n20071) );
  NAND2_X1 U13257 ( .A1(n12325), .A2(n10220), .ZN(n16312) );
  OAI211_X1 U13258 ( .C1(n10220), .C2(n12325), .A(n19342), .B(n16312), .ZN(
        n10899) );
  AND3_X4 U13259 ( .A1(n15781), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U13260 ( .A1(n9709), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10227) );
  AOI22_X1 U13261 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10609), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10226) );
  AND2_X4 U13262 ( .A1(n12269), .A2(n10221), .ZN(n12717) );
  AOI22_X1 U13263 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10225) );
  AND2_X4 U13264 ( .A1(n15788), .A2(n10222), .ZN(n12805) );
  AND3_X4 U13265 ( .A1(n10223), .A2(n10704), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10623) );
  AOI22_X1 U13266 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10224) );
  NAND4_X1 U13267 ( .A1(n10227), .A2(n10226), .A3(n10225), .A4(n10224), .ZN(
        n10228) );
  NAND2_X1 U13268 ( .A1(n10228), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10235) );
  AOI22_X1 U13269 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10231) );
  AOI22_X1 U13270 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10229) );
  NAND4_X1 U13271 ( .A1(n10232), .A2(n10231), .A3(n10230), .A4(n10229), .ZN(
        n10233) );
  NAND2_X1 U13272 ( .A1(n10233), .A2(n10282), .ZN(n10234) );
  NAND2_X2 U13273 ( .A1(n10235), .A2(n10234), .ZN(n10632) );
  AOI22_X1 U13274 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n9709), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10239) );
  AOI22_X1 U13275 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10609), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10238) );
  AOI22_X1 U13276 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12805), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10237) );
  AOI22_X1 U13277 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10236) );
  NAND4_X1 U13278 ( .A1(n10239), .A2(n10238), .A3(n10237), .A4(n10236), .ZN(
        n10240) );
  AOI22_X1 U13279 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10242) );
  AOI22_X1 U13280 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10241) );
  AOI22_X1 U13281 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10609), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10244) );
  AOI22_X1 U13282 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10243) );
  NAND3_X1 U13283 ( .A1(n10183), .A2(n10244), .A3(n10243), .ZN(n10245) );
  NAND2_X1 U13284 ( .A1(n10245), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10246) );
  NAND2_X1 U13285 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10251) );
  NAND2_X1 U13286 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10250) );
  NAND2_X1 U13287 ( .A1(n10623), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10249) );
  NAND2_X1 U13288 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10248) );
  NAND2_X1 U13289 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10253) );
  OR2_X1 U13290 ( .A1(n10277), .A2(n11991), .ZN(n10252) );
  NAND2_X1 U13291 ( .A1(n10255), .A2(n10254), .ZN(n10256) );
  NOR2_X1 U13292 ( .A1(n10257), .A2(n10256), .ZN(n10258) );
  NAND3_X1 U13293 ( .A1(n9784), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10258), .ZN(n10273) );
  NAND2_X1 U13294 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10264) );
  OR2_X1 U13295 ( .A1(n10277), .A2(n10260), .ZN(n10262) );
  NAND2_X1 U13296 ( .A1(n10622), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10261) );
  NAND4_X1 U13297 ( .A1(n10264), .A2(n10263), .A3(n10262), .A4(n10261), .ZN(
        n10270) );
  NAND2_X1 U13298 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10268) );
  NAND2_X1 U13299 ( .A1(n9709), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10267) );
  NAND2_X1 U13300 ( .A1(n10623), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10266) );
  NAND2_X1 U13301 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10265) );
  NAND4_X1 U13302 ( .A1(n10268), .A2(n10267), .A3(n10266), .A4(n10265), .ZN(
        n10269) );
  NOR2_X1 U13303 ( .A1(n10270), .A2(n10269), .ZN(n10271) );
  NAND2_X1 U13304 ( .A1(n10271), .A2(n10283), .ZN(n10272) );
  INV_X1 U13305 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20133) );
  NOR2_X1 U13306 ( .A1(n13415), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10274) );
  NOR2_X1 U13307 ( .A1(n10647), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10374) );
  AOI22_X1 U13308 ( .A1(n14502), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10275) );
  OAI21_X1 U13309 ( .B1(n10566), .B2(n20133), .A(n10275), .ZN(n14500) );
  NAND2_X1 U13310 ( .A1(n10544), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10292) );
  INV_X2 U13311 ( .A(n10373), .ZN(n14502) );
  AOI22_X1 U13312 ( .A1(n14502), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n14501), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10291) );
  AOI22_X1 U13313 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10360), .B1(
        n12620), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10281) );
  AOI22_X1 U13314 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n9717), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10280) );
  AOI22_X1 U13315 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10397), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10279) );
  AND2_X2 U13316 ( .A1(n10622), .A2(n10282), .ZN(n15815) );
  AOI22_X1 U13317 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10513), .B1(
        n15815), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10278) );
  NAND4_X1 U13318 ( .A1(n10281), .A2(n10280), .A3(n10279), .A4(n10278), .ZN(
        n10289) );
  AND2_X2 U13319 ( .A1(n12805), .A2(n10282), .ZN(n12675) );
  AND2_X2 U13320 ( .A1(n12805), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10507) );
  AOI22_X1 U13321 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12675), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10287) );
  AND2_X2 U13322 ( .A1(n9708), .A2(n10282), .ZN(n12676) );
  AOI22_X1 U13323 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12676), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10286) );
  AND2_X2 U13324 ( .A1(n12830), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10505) );
  AND2_X1 U13325 ( .A1(n10620), .A2(n10283), .ZN(n10508) );
  AOI22_X1 U13326 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n10505), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10285) );
  AND2_X2 U13327 ( .A1(n10620), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10506) );
  AOI22_X1 U13328 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12678), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10284) );
  NAND4_X1 U13329 ( .A1(n10287), .A2(n10286), .A3(n10285), .A4(n10284), .ZN(
        n10288) );
  NAND2_X1 U13330 ( .A1(n10534), .A2(n13636), .ZN(n10290) );
  NAND2_X1 U13331 ( .A1(n12620), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10296) );
  NAND2_X1 U13332 ( .A1(n10360), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10295) );
  NAND2_X1 U13333 ( .A1(n9718), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10294) );
  NAND2_X1 U13334 ( .A1(n10348), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10293) );
  NAND2_X1 U13335 ( .A1(n12677), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10300) );
  NAND2_X1 U13336 ( .A1(n12676), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10299) );
  NAND2_X1 U13337 ( .A1(n10505), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10298) );
  NAND2_X1 U13338 ( .A1(n10508), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10297) );
  NAND2_X1 U13339 ( .A1(n10507), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10304) );
  NAND2_X1 U13340 ( .A1(n12675), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10303) );
  NAND2_X1 U13341 ( .A1(n12678), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10302) );
  NAND2_X1 U13342 ( .A1(n10506), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10301) );
  NAND2_X1 U13343 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10308) );
  NAND2_X1 U13344 ( .A1(n10514), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10307) );
  NAND2_X1 U13345 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10306) );
  NAND2_X1 U13346 ( .A1(n15815), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10305) );
  INV_X1 U13347 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n10313) );
  OR2_X1 U13348 ( .A1(n10566), .A2(n10313), .ZN(n10317) );
  INV_X1 U13349 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19478) );
  NAND2_X1 U13350 ( .A1(n10648), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10314) );
  OAI211_X1 U13351 ( .C1(n19478), .C2(n13415), .A(n10314), .B(n19920), .ZN(
        n10315) );
  INV_X1 U13352 ( .A(n10315), .ZN(n10316) );
  NAND2_X1 U13353 ( .A1(n10317), .A2(n10316), .ZN(n13429) );
  AOI22_X1 U13354 ( .A1(n12620), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10321) );
  AOI22_X1 U13355 ( .A1(n9717), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U13356 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U13357 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15815), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10318) );
  NAND4_X1 U13358 ( .A1(n10321), .A2(n10320), .A3(n10319), .A4(n10318), .ZN(
        n10327) );
  AOI22_X1 U13359 ( .A1(n12675), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10325) );
  AOI22_X1 U13360 ( .A1(n12676), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U13361 ( .A1(n10505), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10323) );
  AOI22_X1 U13362 ( .A1(n12678), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10322) );
  NAND4_X1 U13363 ( .A1(n10325), .A2(n10324), .A3(n10323), .A4(n10322), .ZN(
        n10326) );
  NAND2_X1 U13364 ( .A1(n10534), .A2(n16586), .ZN(n10341) );
  AOI22_X1 U13365 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10609), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10331) );
  AOI22_X1 U13366 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U13367 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10329) );
  NAND4_X1 U13368 ( .A1(n10331), .A2(n10330), .A3(n10329), .A4(n10328), .ZN(
        n10332) );
  NAND2_X1 U13369 ( .A1(n10332), .A2(n10282), .ZN(n10339) );
  AOI22_X1 U13370 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13371 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10609), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U13372 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U13373 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10333) );
  NAND4_X1 U13374 ( .A1(n10336), .A2(n10335), .A3(n10334), .A4(n10333), .ZN(
        n10337) );
  NAND2_X1 U13375 ( .A1(n10337), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10338) );
  NAND2_X1 U13376 ( .A1(n12865), .A2(n10374), .ZN(n10371) );
  NAND2_X1 U13377 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10340) );
  NAND4_X1 U13378 ( .A1(n10341), .A2(n10373), .A3(n10371), .A4(n10340), .ZN(
        n13428) );
  NAND2_X1 U13379 ( .A1(n13429), .A2(n13428), .ZN(n13427) );
  AOI22_X1 U13380 ( .A1(n10274), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n10374), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10342) );
  INV_X1 U13381 ( .A(n10358), .ZN(n10343) );
  XNOR2_X1 U13382 ( .A(n13427), .B(n10343), .ZN(n13450) );
  AOI22_X1 U13383 ( .A1(n12620), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10397), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10347) );
  AOI22_X1 U13384 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10514), .B1(
        n10505), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U13385 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10507), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10345) );
  AOI22_X1 U13386 ( .A1(n10360), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10344) );
  NAND4_X1 U13387 ( .A1(n10347), .A2(n10346), .A3(n10345), .A4(n10344), .ZN(
        n10354) );
  AOI22_X1 U13388 ( .A1(n9718), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12676), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10352) );
  AOI22_X1 U13389 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10513), .B1(
        n12675), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10351) );
  AOI22_X1 U13390 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12678), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U13391 ( .A1(n10348), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15815), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10349) );
  NAND4_X1 U13392 ( .A1(n10352), .A2(n10351), .A3(n10350), .A4(n10349), .ZN(
        n10353) );
  NOR2_X1 U13393 ( .A1(n10354), .A2(n10353), .ZN(n12282) );
  NAND2_X1 U13394 ( .A1(n10678), .A2(n13415), .ZN(n13425) );
  OAI21_X1 U13395 ( .B1(n10860), .B2(n10648), .A(n13425), .ZN(n10355) );
  INV_X1 U13396 ( .A(n10355), .ZN(n10357) );
  INV_X1 U13397 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10356) );
  NAND2_X1 U13398 ( .A1(n10358), .A2(n13427), .ZN(n10359) );
  NAND2_X1 U13399 ( .A1(n13449), .A2(n10359), .ZN(n10378) );
  AOI22_X1 U13400 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12678), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10370) );
  AOI22_X1 U13401 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10360), .B1(
        n12620), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10364) );
  AOI22_X1 U13402 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n9717), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10363) );
  AOI22_X1 U13403 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10397), .B1(
        n10513), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U13404 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10514), .B1(
        n15815), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10361) );
  NAND4_X1 U13405 ( .A1(n10364), .A2(n10363), .A3(n10362), .A4(n10361), .ZN(
        n10365) );
  AOI22_X1 U13406 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12676), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10369) );
  AOI22_X1 U13407 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12675), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U13408 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n10505), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10367) );
  NAND2_X1 U13409 ( .A1(n10534), .A2(n10851), .ZN(n10372) );
  OAI211_X1 U13410 ( .C1(n19920), .C2(n20163), .A(n10372), .B(n10371), .ZN(
        n10377) );
  XNOR2_X1 U13411 ( .A(n10378), .B(n10377), .ZN(n13579) );
  NAND2_X1 U13412 ( .A1(n10544), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U13413 ( .A1(n14502), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n14501), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10375) );
  AND2_X1 U13414 ( .A1(n10376), .A2(n10375), .ZN(n13578) );
  INV_X1 U13415 ( .A(n10377), .ZN(n10379) );
  NAND2_X1 U13416 ( .A1(n10379), .A2(n10378), .ZN(n10380) );
  NAND2_X1 U13417 ( .A1(n13577), .A2(n10380), .ZN(n13727) );
  AOI22_X1 U13418 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n9717), .B1(
        n12620), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10384) );
  AOI22_X1 U13419 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10360), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10383) );
  AOI22_X1 U13420 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10397), .B1(
        n10513), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10382) );
  AOI22_X1 U13421 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10514), .B1(
        n15815), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10381) );
  NAND4_X1 U13422 ( .A1(n10384), .A2(n10383), .A3(n10382), .A4(n10381), .ZN(
        n10390) );
  AOI22_X1 U13423 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12675), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10388) );
  AOI22_X1 U13424 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12676), .B1(
        n10505), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10387) );
  AOI22_X1 U13425 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10504), .B1(
        n12678), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U13426 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10508), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10385) );
  NAND4_X1 U13427 ( .A1(n10388), .A2(n10387), .A3(n10386), .A4(n10385), .ZN(
        n10389) );
  NAND2_X1 U13428 ( .A1(n10534), .A2(n12031), .ZN(n10393) );
  NOR2_X1 U13429 ( .A1(n20156), .A2(n19920), .ZN(n10391) );
  AOI21_X1 U13430 ( .B1(n14501), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10391), .ZN(n10392) );
  AND2_X1 U13431 ( .A1(n10393), .A2(n10392), .ZN(n10396) );
  NAND2_X1 U13432 ( .A1(n10544), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10395) );
  NAND2_X1 U13433 ( .A1(n14502), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10394) );
  AOI22_X1 U13434 ( .A1(n10544), .A2(P2_REIP_REG_4__SCAN_IN), .B1(n14502), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n10409) );
  AOI22_X1 U13435 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10360), .B1(
        n12620), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10401) );
  AOI22_X1 U13436 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n9717), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10400) );
  AOI22_X1 U13437 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10397), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10399) );
  INV_X1 U13438 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n20035) );
  AOI22_X1 U13439 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n15815), .B1(
        n10513), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10398) );
  NAND4_X1 U13440 ( .A1(n10401), .A2(n10400), .A3(n10399), .A4(n10398), .ZN(
        n10407) );
  AOI22_X1 U13441 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12675), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10405) );
  AOI22_X1 U13442 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12676), .B1(
        n10504), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10404) );
  AOI22_X1 U13443 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10505), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10403) );
  AOI22_X1 U13444 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12678), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10402) );
  NAND4_X1 U13445 ( .A1(n10405), .A2(n10404), .A3(n10403), .A4(n10402), .ZN(
        n10406) );
  AOI22_X1 U13446 ( .A1(n10534), .A2(n12034), .B1(n14501), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10408) );
  NAND2_X1 U13447 ( .A1(n10409), .A2(n10408), .ZN(n13946) );
  NAND2_X1 U13448 ( .A1(n10544), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n10423) );
  AOI22_X1 U13449 ( .A1(n14502), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n14501), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10422) );
  AOI22_X1 U13450 ( .A1(n12620), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U13451 ( .A1(n9718), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10412) );
  AOI22_X1 U13452 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10411) );
  AOI22_X1 U13453 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15815), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10410) );
  NAND4_X1 U13454 ( .A1(n10413), .A2(n10412), .A3(n10411), .A4(n10410), .ZN(
        n10419) );
  AOI22_X1 U13455 ( .A1(n12675), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10417) );
  AOI22_X1 U13456 ( .A1(n12676), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10416) );
  AOI22_X1 U13457 ( .A1(n12677), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10505), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10415) );
  AOI22_X1 U13458 ( .A1(n12678), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10414) );
  NAND4_X1 U13459 ( .A1(n10417), .A2(n10416), .A3(n10415), .A4(n10414), .ZN(
        n10418) );
  NOR2_X1 U13460 ( .A1(n10419), .A2(n10418), .ZN(n12054) );
  INV_X1 U13461 ( .A(n12054), .ZN(n10420) );
  NAND2_X1 U13462 ( .A1(n10534), .A2(n10420), .ZN(n10421) );
  NAND3_X1 U13463 ( .A1(n10423), .A2(n10422), .A3(n10421), .ZN(n14047) );
  AOI22_X1 U13464 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10360), .B1(
        n12620), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10427) );
  AOI22_X1 U13465 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n9717), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10426) );
  AOI22_X1 U13466 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10514), .B1(
        n10397), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10425) );
  AOI22_X1 U13467 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n15815), .B1(
        n10513), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10424) );
  NAND4_X1 U13468 ( .A1(n10427), .A2(n10426), .A3(n10425), .A4(n10424), .ZN(
        n10433) );
  AOI22_X1 U13469 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12675), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10431) );
  AOI22_X1 U13470 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12676), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10430) );
  AOI22_X1 U13471 ( .A1(n10505), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10429) );
  AOI22_X1 U13472 ( .A1(n12678), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10428) );
  NAND4_X1 U13473 ( .A1(n10431), .A2(n10430), .A3(n10429), .A4(n10428), .ZN(
        n10432) );
  INV_X1 U13474 ( .A(n12089), .ZN(n10434) );
  NAND2_X1 U13475 ( .A1(n10534), .A2(n10434), .ZN(n10435) );
  NAND2_X1 U13476 ( .A1(n10544), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n10437) );
  AOI22_X1 U13477 ( .A1(n14502), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n14501), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10436) );
  NAND2_X1 U13478 ( .A1(n10437), .A2(n10436), .ZN(n13440) );
  AOI21_X1 U13479 ( .B1(n10534), .B2(n12162), .A(n13443), .ZN(n13439) );
  NAND2_X1 U13480 ( .A1(n10544), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n10439) );
  AOI22_X1 U13481 ( .A1(n14502), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n14501), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10438) );
  NOR2_X2 U13482 ( .A1(n13439), .A2(n13438), .ZN(n16557) );
  NAND2_X1 U13483 ( .A1(n10544), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U13484 ( .A1(n14502), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n14501), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10451) );
  AOI22_X1 U13485 ( .A1(n12620), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9718), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U13486 ( .A1(n10360), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10442) );
  AOI22_X1 U13487 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10441) );
  AOI22_X1 U13488 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15815), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10440) );
  NAND4_X1 U13489 ( .A1(n10443), .A2(n10442), .A3(n10441), .A4(n10440), .ZN(
        n10449) );
  AOI22_X1 U13490 ( .A1(n12675), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10447) );
  AOI22_X1 U13491 ( .A1(n12677), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10505), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10446) );
  AOI22_X1 U13492 ( .A1(n12676), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10445) );
  AOI22_X1 U13493 ( .A1(n12678), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10444) );
  NAND4_X1 U13494 ( .A1(n10447), .A2(n10446), .A3(n10445), .A4(n10444), .ZN(
        n10448) );
  NAND2_X1 U13495 ( .A1(n10534), .A2(n13691), .ZN(n10450) );
  NAND3_X1 U13496 ( .A1(n10452), .A2(n10451), .A3(n10450), .ZN(n16558) );
  NAND2_X1 U13497 ( .A1(n16557), .A2(n16558), .ZN(n13433) );
  NAND2_X1 U13498 ( .A1(n10544), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n10465) );
  AOI22_X1 U13499 ( .A1(n14502), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10464) );
  AOI22_X1 U13500 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n9717), .B1(
        n12620), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10456) );
  AOI22_X1 U13501 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10360), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10455) );
  AOI22_X1 U13502 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10513), .B1(
        n10397), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10454) );
  AOI22_X1 U13503 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n10514), .B1(
        n15815), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10453) );
  NAND4_X1 U13504 ( .A1(n10456), .A2(n10455), .A3(n10454), .A4(n10453), .ZN(
        n10462) );
  AOI22_X1 U13505 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12675), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10460) );
  AOI22_X1 U13506 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12676), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10459) );
  AOI22_X1 U13507 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n12677), .B1(
        n10505), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U13508 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12678), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10457) );
  NAND4_X1 U13509 ( .A1(n10460), .A2(n10459), .A3(n10458), .A4(n10457), .ZN(
        n10461) );
  NOR2_X1 U13510 ( .A1(n10462), .A2(n10461), .ZN(n19404) );
  NAND2_X1 U13511 ( .A1(n10534), .A2(n12576), .ZN(n10463) );
  NAND3_X1 U13512 ( .A1(n10465), .A2(n10464), .A3(n10463), .ZN(n13445) );
  NAND2_X1 U13513 ( .A1(n13434), .A2(n13445), .ZN(n13446) );
  NAND2_X1 U13514 ( .A1(n10544), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n10478) );
  AOI22_X1 U13515 ( .A1(n14502), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10477) );
  AOI22_X1 U13516 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10360), .B1(
        n12620), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10469) );
  AOI22_X1 U13517 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n9718), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10468) );
  AOI22_X1 U13518 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10397), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10467) );
  INV_X1 U13519 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19573) );
  AOI22_X1 U13520 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n15815), .B1(
        n10513), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10466) );
  NAND4_X1 U13521 ( .A1(n10469), .A2(n10468), .A3(n10467), .A4(n10466), .ZN(
        n10475) );
  AOI22_X1 U13522 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12675), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10473) );
  AOI22_X1 U13523 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12676), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U13524 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n10505), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10471) );
  AOI22_X1 U13525 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12678), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10470) );
  NAND4_X1 U13526 ( .A1(n10473), .A2(n10472), .A3(n10471), .A4(n10470), .ZN(
        n10474) );
  NAND2_X1 U13527 ( .A1(n10534), .A2(n14013), .ZN(n10476) );
  AOI22_X1 U13528 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n9717), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10482) );
  AOI22_X1 U13529 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10360), .B1(
        n12620), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10481) );
  AOI22_X1 U13530 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10513), .B1(
        n10397), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10480) );
  AOI22_X1 U13531 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10514), .B1(
        n15815), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10479) );
  NAND4_X1 U13532 ( .A1(n10482), .A2(n10481), .A3(n10480), .A4(n10479), .ZN(
        n10488) );
  AOI22_X1 U13533 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12675), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U13534 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12676), .B1(
        n10505), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13535 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12678), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U13536 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12677), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10483) );
  NAND4_X1 U13537 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n10483), .ZN(
        n10487) );
  AOI22_X1 U13538 ( .A1(n10544), .A2(P2_REIP_REG_12__SCAN_IN), .B1(n10534), 
        .B2(n14016), .ZN(n10490) );
  AOI22_X1 U13539 ( .A1(n14502), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10489) );
  NAND2_X1 U13540 ( .A1(n10490), .A2(n10489), .ZN(n13641) );
  NAND2_X1 U13541 ( .A1(n10544), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n10503) );
  AOI22_X1 U13542 ( .A1(n14502), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10502) );
  AOI22_X1 U13543 ( .A1(n12620), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10494) );
  AOI22_X1 U13544 ( .A1(n9718), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10493) );
  AOI22_X1 U13545 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13546 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15815), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10491) );
  NAND4_X1 U13547 ( .A1(n10494), .A2(n10493), .A3(n10492), .A4(n10491), .ZN(
        n10500) );
  AOI22_X1 U13548 ( .A1(n12675), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10498) );
  AOI22_X1 U13549 ( .A1(n12676), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10497) );
  AOI22_X1 U13550 ( .A1(n10505), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10496) );
  AOI22_X1 U13551 ( .A1(n12678), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10495) );
  NAND4_X1 U13552 ( .A1(n10498), .A2(n10497), .A3(n10496), .A4(n10495), .ZN(
        n10499) );
  NAND2_X1 U13553 ( .A1(n10534), .A2(n14141), .ZN(n10501) );
  INV_X1 U13554 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12067) );
  INV_X1 U13555 ( .A(n10504), .ZN(n12637) );
  INV_X1 U13556 ( .A(n10505), .ZN(n12635) );
  INV_X1 U13557 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12061) );
  OAI22_X1 U13558 ( .A1(n12067), .A2(n12637), .B1(n12635), .B2(n12061), .ZN(
        n10512) );
  INV_X1 U13559 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12066) );
  INV_X1 U13560 ( .A(n12676), .ZN(n12639) );
  INV_X1 U13561 ( .A(n10506), .ZN(n12643) );
  INV_X1 U13562 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12070) );
  OAI22_X1 U13563 ( .A1(n12066), .A2(n12639), .B1(n12643), .B2(n12070), .ZN(
        n10511) );
  INV_X1 U13564 ( .A(n12675), .ZN(n12642) );
  INV_X1 U13565 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12072) );
  INV_X1 U13566 ( .A(n10507), .ZN(n12640) );
  INV_X1 U13567 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12073) );
  OAI22_X1 U13568 ( .A1(n12642), .A2(n12072), .B1(n12640), .B2(n12073), .ZN(
        n10510) );
  INV_X1 U13569 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12059) );
  INV_X1 U13570 ( .A(n12678), .ZN(n12645) );
  INV_X1 U13571 ( .A(n10508), .ZN(n12633) );
  INV_X1 U13572 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12075) );
  OAI22_X1 U13573 ( .A1(n12059), .A2(n12645), .B1(n12633), .B2(n12075), .ZN(
        n10509) );
  NOR4_X1 U13574 ( .A1(n10512), .A2(n10511), .A3(n10510), .A4(n10509), .ZN(
        n10520) );
  AOI22_X1 U13575 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n9717), .B1(
        n12620), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10519) );
  AOI22_X1 U13576 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10360), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10518) );
  INV_X1 U13577 ( .A(n10513), .ZN(n12654) );
  INV_X1 U13578 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19582) );
  NOR2_X1 U13579 ( .A1(n12654), .A2(n19582), .ZN(n10516) );
  INV_X1 U13580 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12065) );
  INV_X1 U13581 ( .A(n10514), .ZN(n12651) );
  INV_X1 U13582 ( .A(n15815), .ZN(n12653) );
  INV_X1 U13583 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12080) );
  OAI22_X1 U13584 ( .A1(n12065), .A2(n12651), .B1(n12653), .B2(n12080), .ZN(
        n10515) );
  AOI211_X1 U13585 ( .C1(n10397), .C2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n10516), .B(n10515), .ZN(n10517) );
  NAND4_X1 U13586 ( .A1(n10520), .A2(n10519), .A3(n10518), .A4(n10517), .ZN(
        n14143) );
  AOI22_X1 U13587 ( .A1(n14143), .A2(n10534), .B1(P2_REIP_REG_14__SCAN_IN), 
        .B2(n10544), .ZN(n10522) );
  AOI22_X1 U13588 ( .A1(n14502), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10521) );
  NAND2_X1 U13589 ( .A1(n10522), .A2(n10521), .ZN(n15693) );
  NAND2_X1 U13590 ( .A1(n10544), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13591 ( .A1(n14502), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13592 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10360), .B1(
        n12620), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U13593 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n9717), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10525) );
  AOI22_X1 U13594 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10397), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10524) );
  INV_X1 U13595 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19592) );
  AOI22_X1 U13596 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n15815), .B1(
        n10513), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10523) );
  NAND4_X1 U13597 ( .A1(n10526), .A2(n10525), .A3(n10524), .A4(n10523), .ZN(
        n10532) );
  AOI22_X1 U13598 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12675), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10530) );
  AOI22_X1 U13599 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12676), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10529) );
  AOI22_X1 U13600 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n10505), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10528) );
  AOI22_X1 U13601 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12678), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10527) );
  NAND4_X1 U13602 ( .A1(n10530), .A2(n10529), .A3(n10528), .A4(n10527), .ZN(
        n10531) );
  INV_X1 U13603 ( .A(n14292), .ZN(n10533) );
  NAND2_X1 U13604 ( .A1(n10534), .A2(n10533), .ZN(n10535) );
  NAND2_X1 U13605 ( .A1(n10544), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10539) );
  AOI22_X1 U13606 ( .A1(n14502), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10538) );
  NAND2_X1 U13607 ( .A1(n10539), .A2(n10538), .ZN(n14302) );
  NAND2_X1 U13608 ( .A1(n10544), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U13609 ( .A1(n14502), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10540) );
  NAND2_X1 U13610 ( .A1(n10541), .A2(n10540), .ZN(n14365) );
  AND2_X2 U13611 ( .A1(n14366), .A2(n14365), .ZN(n14401) );
  NAND2_X1 U13612 ( .A1(n10544), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n10543) );
  AOI22_X1 U13613 ( .A1(n14502), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10542) );
  NAND2_X1 U13614 ( .A1(n10543), .A2(n10542), .ZN(n14400) );
  NAND2_X1 U13615 ( .A1(n14401), .A2(n14400), .ZN(n14424) );
  NAND2_X1 U13616 ( .A1(n10544), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n10546) );
  AOI22_X1 U13617 ( .A1(n14502), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10545) );
  NOR2_X2 U13618 ( .A1(n14424), .A2(n14425), .ZN(n15364) );
  NAND2_X1 U13619 ( .A1(n10544), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n10548) );
  AOI22_X1 U13620 ( .A1(n14502), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10547) );
  NAND2_X1 U13621 ( .A1(n10548), .A2(n10547), .ZN(n15365) );
  NAND2_X1 U13622 ( .A1(n15364), .A2(n15365), .ZN(n15366) );
  NAND2_X1 U13623 ( .A1(n10544), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n10550) );
  AOI22_X1 U13624 ( .A1(n14502), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10549) );
  NAND2_X1 U13625 ( .A1(n10544), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n10552) );
  AOI22_X1 U13626 ( .A1(n14502), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10551) );
  NAND2_X1 U13627 ( .A1(n10552), .A2(n10551), .ZN(n15158) );
  NAND2_X1 U13628 ( .A1(n10544), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n10554) );
  AOI22_X1 U13629 ( .A1(n14502), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10553) );
  NAND2_X1 U13630 ( .A1(n10554), .A2(n10553), .ZN(n15145) );
  NAND2_X1 U13631 ( .A1(n10544), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U13632 ( .A1(n14502), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10555) );
  NAND2_X1 U13633 ( .A1(n10544), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n10558) );
  AOI22_X1 U13634 ( .A1(n14502), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10557) );
  INV_X1 U13635 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20124) );
  AOI22_X1 U13636 ( .A1(n14502), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10559) );
  OAI21_X1 U13637 ( .B1(n10566), .B2(n20124), .A(n10559), .ZN(n15324) );
  NAND2_X1 U13638 ( .A1(n15323), .A2(n15324), .ZN(n15326) );
  NAND2_X1 U13639 ( .A1(n10544), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n10561) );
  AOI22_X1 U13640 ( .A1(n14502), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10560) );
  AND2_X1 U13641 ( .A1(n10561), .A2(n10560), .ZN(n15315) );
  NOR2_X2 U13642 ( .A1(n15326), .A2(n15315), .ZN(n15305) );
  NAND2_X1 U13643 ( .A1(n10544), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n10563) );
  AOI22_X1 U13644 ( .A1(n14502), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10562) );
  AND2_X1 U13645 ( .A1(n10563), .A2(n10562), .ZN(n15306) );
  INV_X1 U13646 ( .A(n15306), .ZN(n10564) );
  INV_X1 U13647 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U13648 ( .A1(n14502), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10565) );
  OAI21_X1 U13649 ( .B1(n10566), .B2(n10841), .A(n10565), .ZN(n15297) );
  AND2_X2 U13650 ( .A1(n15296), .A2(n15297), .ZN(n15299) );
  XOR2_X1 U13651 ( .A(n14500), .B(n15299), .Z(n12880) );
  INV_X1 U13652 ( .A(n12880), .ZN(n10639) );
  MUX2_X1 U13653 ( .A(n10356), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12266) );
  NAND2_X1 U13654 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20182), .ZN(
        n12112) );
  INV_X1 U13655 ( .A(n12112), .ZN(n10567) );
  NAND2_X1 U13656 ( .A1(n12266), .A2(n10567), .ZN(n10577) );
  NAND2_X1 U13657 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n10356), .ZN(
        n10568) );
  NAND2_X1 U13658 ( .A1(n10577), .A2(n10568), .ZN(n10585) );
  MUX2_X1 U13659 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n20156), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10581) );
  NAND2_X1 U13660 ( .A1(n20156), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10570) );
  NAND2_X1 U13661 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12270), .ZN(
        n10572) );
  NAND2_X1 U13662 ( .A1(n10573), .A2(n10572), .ZN(n10575) );
  NAND2_X1 U13663 ( .A1(n16626), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10574) );
  INV_X1 U13664 ( .A(n12266), .ZN(n10576) );
  NAND2_X1 U13665 ( .A1(n10576), .A2(n12112), .ZN(n10578) );
  AND2_X1 U13666 ( .A1(n10578), .A2(n10577), .ZN(n12449) );
  NOR2_X1 U13667 ( .A1(n16626), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10579) );
  NAND2_X1 U13668 ( .A1(n10580), .A2(n10579), .ZN(n10866) );
  INV_X1 U13669 ( .A(n10581), .ZN(n10582) );
  XNOR2_X1 U13670 ( .A(n10583), .B(n10582), .ZN(n10861) );
  XOR2_X1 U13671 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .Z(n10584) );
  XNOR2_X1 U13672 ( .A(n10585), .B(n10584), .ZN(n12451) );
  NAND2_X1 U13673 ( .A1(n12458), .A2(n12451), .ZN(n12273) );
  INV_X1 U13674 ( .A(n12273), .ZN(n10586) );
  NAND2_X1 U13675 ( .A1(n12449), .A2(n10586), .ZN(n10587) );
  AOI22_X1 U13676 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10591) );
  AOI22_X1 U13677 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U13678 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10588) );
  AOI22_X1 U13679 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10590) );
  NAND3_X1 U13680 ( .A1(n10591), .A2(n10184), .A3(n10590), .ZN(n10598) );
  AOI22_X1 U13681 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U13682 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10600) );
  AOI22_X1 U13683 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10599) );
  AOI22_X1 U13684 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10602) );
  AOI22_X1 U13685 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10601) );
  NAND2_X1 U13686 ( .A1(n10641), .A2(n10642), .ZN(n10615) );
  AOI22_X1 U13687 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10605) );
  AOI22_X1 U13688 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10604) );
  AOI22_X1 U13689 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10603) );
  NAND3_X1 U13690 ( .A1(n10606), .A2(n10605), .A3(n10173), .ZN(n10614) );
  AOI22_X1 U13691 ( .A1(n9709), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10608) );
  AOI22_X1 U13692 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10609), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10611) );
  AOI22_X1 U13693 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10610) );
  NAND4_X1 U13694 ( .A1(n10612), .A2(n10611), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A4(n10610), .ZN(n10613) );
  AOI22_X1 U13696 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9707), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13697 ( .A1(n10623), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10618) );
  AOI22_X1 U13698 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10609), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10617) );
  NAND4_X1 U13699 ( .A1(n10619), .A2(n10618), .A3(n10617), .A4(n10616), .ZN(
        n10630) );
  AOI22_X1 U13700 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10628) );
  AOI22_X1 U13701 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10609), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10627) );
  AOI22_X1 U13702 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10626) );
  AOI22_X1 U13703 ( .A1(n9709), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10625) );
  NAND4_X1 U13704 ( .A1(n10628), .A2(n10627), .A3(n10626), .A4(n10625), .ZN(
        n10629) );
  NAND2_X1 U13705 ( .A1(n15777), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20064) );
  AND2_X1 U13706 ( .A1(n16615), .A2(n13350), .ZN(n12278) );
  NAND2_X2 U13707 ( .A1(n20216), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n20132) );
  NOR2_X1 U13708 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19196) );
  INV_X1 U13709 ( .A(n19196), .ZN(n20083) );
  NAND2_X1 U13710 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20202) );
  NAND2_X1 U13711 ( .A1(n20208), .A2(n20202), .ZN(n13340) );
  NAND2_X1 U13712 ( .A1(n19595), .A2(n13267), .ZN(n16629) );
  INV_X1 U13713 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10638) );
  NAND2_X1 U13714 ( .A1(n10692), .A2(n16615), .ZN(n10635) );
  INV_X1 U13715 ( .A(n10631), .ZN(n10634) );
  INV_X2 U13716 ( .A(n10680), .ZN(n10656) );
  AND2_X2 U13717 ( .A1(n10656), .A2(n10632), .ZN(n12472) );
  NOR2_X1 U13718 ( .A1(n10641), .A2(n10642), .ZN(n10633) );
  NAND2_X1 U13719 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20065), .ZN(n20067) );
  NOR2_X1 U13720 ( .A1(n20064), .A2(n20067), .ZN(n16627) );
  NAND2_X1 U13721 ( .A1(n20157), .A2(n15777), .ZN(n19193) );
  INV_X1 U13722 ( .A(n19193), .ZN(n13271) );
  AND2_X2 U13723 ( .A1(n13271), .A2(n20201), .ZN(n19517) );
  NOR2_X1 U13724 ( .A1(n16627), .A2(n19517), .ZN(n10636) );
  NAND2_X1 U13725 ( .A1(n20071), .A2(n10636), .ZN(n10637) );
  OAI22_X1 U13726 ( .A1(n10639), .A2(n19381), .B1(n10638), .B2(n19391), .ZN(
        n10640) );
  AND2_X1 U13727 ( .A1(n19565), .A2(n10647), .ZN(n12489) );
  NOR2_X1 U13728 ( .A1(n12504), .A2(n16615), .ZN(n12488) );
  AND2_X1 U13729 ( .A1(n12549), .A2(n9720), .ZN(n10644) );
  MUX2_X1 U13730 ( .A(n12865), .B(n10649), .S(n9853), .Z(n10653) );
  NAND2_X1 U13731 ( .A1(n20199), .A2(n10647), .ZN(n10650) );
  BUF_X1 U13732 ( .A(n10739), .Z(n10779) );
  NAND2_X1 U13733 ( .A1(n10779), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10665) );
  INV_X1 U13734 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n10662) );
  AND2_X1 U13735 ( .A1(n10657), .A2(n10656), .ZN(n10658) );
  AND3_X2 U13736 ( .A1(n12491), .A2(n12446), .A3(n12495), .ZN(n12508) );
  NAND2_X1 U13737 ( .A1(n10838), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10661) );
  NAND2_X1 U13738 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10660) );
  OAI211_X1 U13739 ( .C1(n10848), .C2(n10662), .A(n10661), .B(n10660), .ZN(
        n10663) );
  INV_X1 U13740 ( .A(n10663), .ZN(n10664) );
  NAND2_X1 U13741 ( .A1(n10665), .A2(n10664), .ZN(n15143) );
  NAND2_X1 U13742 ( .A1(n10779), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10671) );
  INV_X1 U13743 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n10668) );
  NAND2_X1 U13744 ( .A1(n10838), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10667) );
  NAND2_X1 U13745 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10666) );
  OAI211_X1 U13746 ( .C1(n10848), .C2(n10668), .A(n10667), .B(n10666), .ZN(
        n10669) );
  INV_X1 U13747 ( .A(n10669), .ZN(n10670) );
  NAND2_X1 U13748 ( .A1(n10671), .A2(n10670), .ZN(n14295) );
  INV_X1 U13749 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10673) );
  NAND2_X1 U13750 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10672) );
  NAND2_X1 U13751 ( .A1(n10678), .A2(n12504), .ZN(n10682) );
  OAI21_X1 U13752 ( .B1(n10680), .B2(n12465), .A(n10679), .ZN(n10681) );
  INV_X1 U13753 ( .A(n12472), .ZN(n10687) );
  NAND4_X1 U13754 ( .A1(n10682), .A2(n10681), .A3(n19565), .A4(n10687), .ZN(
        n10684) );
  NAND3_X1 U13755 ( .A1(n10684), .A2(n10683), .A3(n20199), .ZN(n12501) );
  NAND2_X1 U13756 ( .A1(n10709), .A2(n12497), .ZN(n10685) );
  NAND2_X1 U13757 ( .A1(n10685), .A2(n20199), .ZN(n10686) );
  INV_X1 U13758 ( .A(n9683), .ZN(n10688) );
  OAI21_X1 U13759 ( .B1(n12504), .B2(n12497), .A(n12446), .ZN(n10689) );
  INV_X1 U13760 ( .A(n10689), .ZN(n10690) );
  NOR2_X1 U13761 ( .A1(n12492), .A2(n10647), .ZN(n10691) );
  NAND2_X1 U13762 ( .A1(n12264), .A2(n10691), .ZN(n10694) );
  INV_X1 U13763 ( .A(n10692), .ZN(n10693) );
  NAND2_X1 U13764 ( .A1(n10694), .A2(n10693), .ZN(n10718) );
  INV_X1 U13765 ( .A(n10718), .ZN(n10695) );
  NAND2_X1 U13766 ( .A1(n10695), .A2(n16615), .ZN(n10696) );
  NAND3_X1 U13767 ( .A1(n10696), .A2(n10697), .A3(n10712), .ZN(n10698) );
  AND2_X2 U13768 ( .A1(n10698), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10747) );
  NAND2_X1 U13769 ( .A1(n10747), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10702) );
  AND2_X2 U13770 ( .A1(n10702), .A2(n10701), .ZN(n10725) );
  INV_X1 U13771 ( .A(n10705), .ZN(n10707) );
  INV_X1 U13772 ( .A(n16631), .ZN(n10716) );
  NOR2_X1 U13773 ( .A1(n10716), .A2(n20182), .ZN(n10706) );
  NAND2_X1 U13774 ( .A1(n10739), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10724) );
  INV_X1 U13775 ( .A(n12502), .ZN(n10711) );
  INV_X1 U13776 ( .A(n10709), .ZN(n12496) );
  AOI21_X1 U13777 ( .B1(n12496), .B2(n12497), .A(n12504), .ZN(n10710) );
  AOI21_X1 U13778 ( .B1(n10711), .B2(n12504), .A(n10710), .ZN(n10714) );
  INV_X1 U13779 ( .A(n10712), .ZN(n10713) );
  NAND2_X1 U13780 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10715) );
  NAND2_X1 U13781 ( .A1(n10716), .A2(n10715), .ZN(n10717) );
  AOI21_X1 U13782 ( .B1(n10757), .B2(P2_REIP_REG_0__SCAN_IN), .A(n10717), .ZN(
        n10721) );
  NAND2_X1 U13783 ( .A1(n10695), .A2(n12463), .ZN(n10719) );
  NAND2_X1 U13784 ( .A1(n11957), .A2(n11952), .ZN(n10729) );
  INV_X1 U13785 ( .A(n10725), .ZN(n10727) );
  NAND2_X2 U13786 ( .A1(n10729), .A2(n10728), .ZN(n11962) );
  NAND2_X1 U13787 ( .A1(n10747), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10731) );
  AOI21_X1 U13788 ( .B1(n20201), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10730) );
  INV_X1 U13789 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n10734) );
  NAND2_X1 U13790 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10732) );
  OAI211_X1 U13791 ( .C1(n10742), .C2(n10734), .A(n10733), .B(n10732), .ZN(
        n10735) );
  INV_X1 U13792 ( .A(n10735), .ZN(n10737) );
  NAND2_X1 U13793 ( .A1(n10739), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10736) );
  INV_X1 U13794 ( .A(n11960), .ZN(n10738) );
  NAND2_X1 U13795 ( .A1(n10739), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10745) );
  INV_X1 U13796 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n14034) );
  NAND2_X1 U13797 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10740) );
  OAI211_X1 U13798 ( .C1(n10742), .C2(n14034), .A(n10741), .B(n10740), .ZN(
        n10743) );
  INV_X1 U13799 ( .A(n10743), .ZN(n10744) );
  AND2_X1 U13800 ( .A1(n16631), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10746) );
  AOI21_X2 U13801 ( .B1(n10747), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10746), .ZN(n10748) );
  INV_X1 U13802 ( .A(n10748), .ZN(n10749) );
  INV_X1 U13803 ( .A(n19369), .ZN(n10756) );
  INV_X1 U13804 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n10753) );
  NAND2_X1 U13805 ( .A1(n10838), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n10752) );
  NAND2_X1 U13806 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10751) );
  OAI211_X1 U13807 ( .C1(n10848), .C2(n10753), .A(n10752), .B(n10751), .ZN(
        n10754) );
  AOI21_X1 U13808 ( .B1(n10779), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n10754), .ZN(n19368) );
  NAND2_X1 U13809 ( .A1(n10756), .A2(n10755), .ZN(n14492) );
  INV_X1 U13810 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n10760) );
  NAND2_X1 U13811 ( .A1(n10838), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n10759) );
  NAND2_X1 U13812 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10758) );
  OAI211_X1 U13813 ( .C1(n10848), .C2(n10760), .A(n10759), .B(n10758), .ZN(
        n10761) );
  AOI21_X1 U13814 ( .B1(n10779), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n10761), .ZN(n14493) );
  NAND2_X1 U13815 ( .A1(n10838), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n10763) );
  NAND2_X1 U13816 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10762) );
  OAI211_X1 U13817 ( .C1(n10848), .C2(n20096), .A(n10763), .B(n10762), .ZN(
        n10764) );
  AOI21_X1 U13818 ( .B1(n10779), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n10764), .ZN(n13543) );
  INV_X1 U13819 ( .A(n10779), .ZN(n10813) );
  INV_X1 U13820 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15763) );
  INV_X1 U13821 ( .A(n10848), .ZN(n10830) );
  AOI22_X1 U13822 ( .A1(n10830), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10766) );
  NAND2_X1 U13823 ( .A1(n10838), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n10765) );
  OAI211_X1 U13824 ( .C1(n10813), .C2(n15763), .A(n10766), .B(n10765), .ZN(
        n13566) );
  NAND2_X1 U13825 ( .A1(n13567), .A2(n13566), .ZN(n13565) );
  INV_X1 U13826 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n10767) );
  INV_X1 U13827 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n19334) );
  OAI22_X1 U13828 ( .A1(n10848), .A2(n10767), .B1(n15777), .B2(n19334), .ZN(
        n10769) );
  INV_X1 U13829 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12310) );
  NOR2_X1 U13830 ( .A1(n10813), .A2(n12310), .ZN(n10768) );
  AOI211_X1 U13831 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n10838), .A(n10769), .B(
        n10768), .ZN(n13688) );
  NAND2_X1 U13832 ( .A1(n10779), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10774) );
  INV_X1 U13833 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n15185) );
  NAND2_X1 U13834 ( .A1(n10838), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10771) );
  NAND2_X1 U13835 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10770) );
  OAI211_X1 U13836 ( .C1(n10848), .C2(n15185), .A(n10771), .B(n10770), .ZN(
        n10772) );
  INV_X1 U13837 ( .A(n10772), .ZN(n10773) );
  NAND2_X1 U13838 ( .A1(n10774), .A2(n10773), .ZN(n13637) );
  NAND2_X1 U13839 ( .A1(n13687), .A2(n13637), .ZN(n15733) );
  INV_X1 U13840 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n10777) );
  NAND2_X1 U13841 ( .A1(n10838), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10776) );
  NAND2_X1 U13842 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10775) );
  OAI211_X1 U13843 ( .C1(n10848), .C2(n10777), .A(n10776), .B(n10775), .ZN(
        n10778) );
  AOI21_X1 U13844 ( .B1(n10779), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n10778), .ZN(n15732) );
  INV_X1 U13845 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n10783) );
  NAND2_X1 U13846 ( .A1(n10845), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10782) );
  NAND2_X1 U13847 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10781) );
  OAI211_X1 U13848 ( .C1(n10848), .C2(n10783), .A(n10782), .B(n10781), .ZN(
        n10784) );
  AOI21_X1 U13849 ( .B1(n10779), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n10784), .ZN(n13242) );
  INV_X1 U13850 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n10787) );
  NAND2_X1 U13851 ( .A1(n10779), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10786) );
  AOI22_X1 U13852 ( .A1(n10830), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n10785) );
  OAI211_X1 U13853 ( .C1(n10787), .C2(n10834), .A(n10786), .B(n10785), .ZN(
        n14009) );
  INV_X1 U13854 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10790) );
  NAND2_X1 U13855 ( .A1(n10779), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10789) );
  AOI22_X1 U13856 ( .A1(n10830), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n10788) );
  OAI211_X1 U13857 ( .C1(n10790), .C2(n10834), .A(n10789), .B(n10788), .ZN(
        n13973) );
  INV_X1 U13858 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n10793) );
  NAND2_X1 U13859 ( .A1(n10838), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10792) );
  NAND2_X1 U13860 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10791) );
  OAI211_X1 U13861 ( .C1(n10848), .C2(n10793), .A(n10792), .B(n10791), .ZN(
        n10794) );
  AOI21_X1 U13862 ( .B1(n10779), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n10794), .ZN(n14145) );
  INV_X1 U13863 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n15684) );
  NAND2_X1 U13864 ( .A1(n10838), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10796) );
  NAND2_X1 U13865 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10795) );
  OAI211_X1 U13866 ( .C1(n10848), .C2(n15684), .A(n10796), .B(n10795), .ZN(
        n10797) );
  AOI21_X1 U13867 ( .B1(n10779), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10797), .ZN(n15522) );
  INV_X1 U13868 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n15672) );
  NAND2_X1 U13869 ( .A1(n10845), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10799) );
  NAND2_X1 U13870 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10798) );
  OAI211_X1 U13871 ( .C1(n10848), .C2(n15672), .A(n10799), .B(n10798), .ZN(
        n10800) );
  AOI21_X1 U13872 ( .B1(n10779), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10800), .ZN(n14431) );
  INV_X1 U13873 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U13874 ( .A1(n10830), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n10802) );
  NAND2_X1 U13875 ( .A1(n10838), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10801) );
  OAI211_X1 U13876 ( .C1(n10813), .C2(n10803), .A(n10802), .B(n10801), .ZN(
        n15504) );
  INV_X1 U13877 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n15493) );
  NAND2_X1 U13878 ( .A1(n10838), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10805) );
  NAND2_X1 U13879 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10804) );
  OAI211_X1 U13880 ( .C1(n10848), .C2(n15493), .A(n10805), .B(n10804), .ZN(
        n10806) );
  AOI21_X1 U13881 ( .B1(n10779), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n10806), .ZN(n15286) );
  INV_X1 U13882 ( .A(n10807), .ZN(n15284) );
  INV_X1 U13883 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20115) );
  NAND2_X1 U13884 ( .A1(n10838), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10809) );
  NAND2_X1 U13885 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10808) );
  OAI211_X1 U13886 ( .C1(n10848), .C2(n20115), .A(n10809), .B(n10808), .ZN(
        n10810) );
  AOI21_X1 U13887 ( .B1(n10779), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n10810), .ZN(n15483) );
  INV_X1 U13888 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15470) );
  AOI22_X1 U13889 ( .A1(n10830), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n10812) );
  NAND2_X1 U13890 ( .A1(n10838), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10811) );
  OAI211_X1 U13891 ( .C1(n10813), .C2(n15470), .A(n10812), .B(n10811), .ZN(
        n15175) );
  INV_X1 U13892 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n10816) );
  NAND2_X1 U13893 ( .A1(n10838), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10815) );
  NAND2_X1 U13894 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10814) );
  OAI211_X1 U13895 ( .C1(n10848), .C2(n10816), .A(n10815), .B(n10814), .ZN(
        n10817) );
  AOI21_X1 U13896 ( .B1(n10779), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n10817), .ZN(n15154) );
  INV_X1 U13897 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n10820) );
  NAND2_X1 U13898 ( .A1(n10838), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10819) );
  NAND2_X1 U13899 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10818) );
  OAI211_X1 U13900 ( .C1(n10848), .C2(n10820), .A(n10819), .B(n10818), .ZN(
        n10821) );
  AOI21_X1 U13901 ( .B1(n10779), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n10821), .ZN(n15428) );
  INV_X1 U13902 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20122) );
  NAND2_X1 U13903 ( .A1(n10838), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10823) );
  NAND2_X1 U13904 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10822) );
  OAI211_X1 U13905 ( .C1(n10848), .C2(n20122), .A(n10823), .B(n10822), .ZN(
        n10824) );
  AOI21_X1 U13906 ( .B1(n10779), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n10824), .ZN(n15275) );
  NAND2_X1 U13907 ( .A1(n10779), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10829) );
  NAND2_X1 U13908 ( .A1(n10838), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10826) );
  NAND2_X1 U13909 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10825) );
  OAI211_X1 U13910 ( .C1(n10848), .C2(n20124), .A(n10826), .B(n10825), .ZN(
        n10827) );
  INV_X1 U13911 ( .A(n10827), .ZN(n10828) );
  NAND2_X1 U13912 ( .A1(n10829), .A2(n10828), .ZN(n15266) );
  INV_X1 U13913 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n10833) );
  NAND2_X1 U13914 ( .A1(n10779), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10832) );
  AOI22_X1 U13915 ( .A1(n10830), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n10831) );
  OAI211_X1 U13916 ( .C1(n10834), .C2(n10833), .A(n10832), .B(n10831), .ZN(
        n15260) );
  INV_X1 U13917 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20128) );
  NAND2_X1 U13918 ( .A1(n10838), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10836) );
  NAND2_X1 U13919 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10835) );
  OAI211_X1 U13920 ( .C1(n10848), .C2(n20128), .A(n10836), .B(n10835), .ZN(
        n10837) );
  AOI21_X1 U13921 ( .B1(n10779), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n10837), .ZN(n15251) );
  NAND2_X1 U13922 ( .A1(n10779), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10844) );
  NAND2_X1 U13923 ( .A1(n10838), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10840) );
  NAND2_X1 U13924 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10839) );
  OAI211_X1 U13925 ( .C1(n10848), .C2(n10841), .A(n10840), .B(n10839), .ZN(
        n10842) );
  INV_X1 U13926 ( .A(n10842), .ZN(n10843) );
  NAND2_X1 U13927 ( .A1(n10844), .A2(n10843), .ZN(n15239) );
  NAND2_X1 U13928 ( .A1(n10845), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10847) );
  NAND2_X1 U13929 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10846) );
  OAI211_X1 U13930 ( .C1(n10848), .C2(n20133), .A(n10847), .B(n10846), .ZN(
        n10849) );
  AOI21_X1 U13931 ( .B1(n10779), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n10849), .ZN(n12897) );
  INV_X1 U13932 ( .A(n12322), .ZN(n10896) );
  NAND2_X1 U13933 ( .A1(n20202), .A2(n19595), .ZN(n10887) );
  NOR2_X1 U13934 ( .A1(n10885), .A2(n10887), .ZN(n10850) );
  INV_X1 U13935 ( .A(n12451), .ZN(n10852) );
  INV_X1 U13936 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n15230) );
  INV_X1 U13937 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n10858) );
  NAND3_X1 U13938 ( .A1(n9720), .A2(n15230), .A3(n10858), .ZN(n10859) );
  NAND2_X1 U13939 ( .A1(n10860), .A2(n10859), .ZN(n12105) );
  NOR2_X1 U13940 ( .A1(n10885), .A2(n9720), .ZN(n12115) );
  NAND2_X1 U13941 ( .A1(n12115), .A2(n12031), .ZN(n10865) );
  AND2_X1 U13942 ( .A1(n10885), .A2(n10855), .ZN(n12114) );
  NAND2_X1 U13943 ( .A1(n12114), .A2(n10861), .ZN(n10864) );
  INV_X1 U13944 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10862) );
  NAND2_X1 U13945 ( .A1(n9720), .A2(n10862), .ZN(n10863) );
  INV_X1 U13946 ( .A(n10866), .ZN(n10868) );
  INV_X1 U13947 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n19414) );
  NOR2_X1 U13948 ( .A1(n10855), .A2(n19414), .ZN(n10867) );
  AOI21_X1 U13949 ( .B1(n12114), .B2(n10868), .A(n10867), .ZN(n10870) );
  INV_X1 U13950 ( .A(n12034), .ZN(n12295) );
  NAND2_X1 U13951 ( .A1(n12115), .A2(n12295), .ZN(n10869) );
  NAND2_X1 U13952 ( .A1(n12125), .A2(n12124), .ZN(n12128) );
  MUX2_X1 U13953 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n12054), .S(n10855), .Z(
        n12127) );
  MUX2_X1 U13954 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n12089), .S(n10855), .Z(
        n12094) );
  NOR2_X2 U13955 ( .A1(n12130), .A2(n12094), .ZN(n12097) );
  MUX2_X1 U13956 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n12101), .S(n10855), .Z(
        n12096) );
  INV_X1 U13957 ( .A(n12096), .ZN(n10873) );
  INV_X1 U13958 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n19335) );
  NOR2_X1 U13959 ( .A1(n10855), .A2(n19335), .ZN(n12098) );
  INV_X1 U13960 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n19410) );
  NAND2_X1 U13961 ( .A1(n12155), .A2(n19410), .ZN(n12158) );
  NOR2_X2 U13962 ( .A1(n12158), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n12166) );
  NAND2_X1 U13963 ( .A1(n9720), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12167) );
  NAND2_X1 U13964 ( .A1(n9720), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12189) );
  OAI21_X1 U13965 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n9720), .ZN(n10874) );
  INV_X1 U13966 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n12181) );
  INV_X1 U13967 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10875) );
  NAND2_X1 U13968 ( .A1(n12181), .A2(n10875), .ZN(n10876) );
  NAND2_X1 U13969 ( .A1(n9720), .A2(n10876), .ZN(n10877) );
  INV_X1 U13970 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n19241) );
  NOR2_X1 U13971 ( .A1(n10855), .A2(n19241), .ZN(n12178) );
  INV_X1 U13972 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n19231) );
  NOR2_X1 U13973 ( .A1(n10855), .A2(n19231), .ZN(n12177) );
  INV_X1 U13974 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n16401) );
  NAND2_X1 U13975 ( .A1(n12221), .A2(n12235), .ZN(n12194) );
  NAND2_X1 U13976 ( .A1(n9720), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12219) );
  INV_X1 U13977 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10878) );
  NOR2_X1 U13978 ( .A1(n10855), .A2(n10878), .ZN(n12226) );
  INV_X1 U13979 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10879) );
  INV_X1 U13980 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n10880) );
  NAND2_X1 U13981 ( .A1(n12233), .A2(n10880), .ZN(n12238) );
  NAND2_X1 U13982 ( .A1(n9720), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12241) );
  INV_X1 U13983 ( .A(n12250), .ZN(n10881) );
  NAND2_X1 U13984 ( .A1(n9720), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12248) );
  NAND2_X1 U13985 ( .A1(n10881), .A2(n12248), .ZN(n12257) );
  INV_X1 U13986 ( .A(n12257), .ZN(n10882) );
  NAND2_X1 U13987 ( .A1(n9720), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12258) );
  NAND2_X1 U13988 ( .A1(n10882), .A2(n12258), .ZN(n12891) );
  NAND2_X1 U13989 ( .A1(n9720), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10883) );
  XNOR2_X1 U13990 ( .A(n12891), .B(n10883), .ZN(n12260) );
  INV_X1 U13991 ( .A(n12260), .ZN(n12261) );
  NAND2_X1 U13992 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n10887), .ZN(n10884) );
  NOR2_X1 U13993 ( .A1(n10885), .A2(n10884), .ZN(n10886) );
  INV_X1 U13994 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n10892) );
  INV_X1 U13995 ( .A(n10887), .ZN(n10888) );
  NOR2_X1 U13996 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n10888), .ZN(n10889) );
  OAI22_X1 U13997 ( .A1(n12030), .A2(n10889), .B1(P2_STATEBS16_REG_SCAN_IN), 
        .B2(n13340), .ZN(n10890) );
  INV_X1 U13998 ( .A(n10890), .ZN(n10891) );
  OAI22_X1 U13999 ( .A1(n10892), .A2(n19382), .B1(n20133), .B2(n19387), .ZN(
        n10893) );
  NAND3_X1 U14000 ( .A1(n10899), .A2(n10898), .A3(n10897), .ZN(P2_U2825) );
  INV_X1 U14001 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10900) );
  NOR2_X4 U14002 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14061) );
  AOI22_X1 U14003 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11072), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10905) );
  NOR2_X2 U14004 ( .A1(n11133), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14065) );
  INV_X1 U14005 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10901) );
  AND2_X2 U14006 ( .A1(n10901), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10907) );
  AOI22_X1 U14007 ( .A1(n11098), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11143), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10904) );
  AOI22_X1 U14008 ( .A1(n10948), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10903) );
  AOI22_X1 U14009 ( .A1(n11145), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10902) );
  NAND4_X1 U14010 ( .A1(n10905), .A2(n10904), .A3(n10903), .A4(n10902), .ZN(
        n10914) );
  AOI22_X1 U14011 ( .A1(n10933), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10912) );
  AND2_X2 U14012 ( .A1(n10906), .A2(n14065), .ZN(n11698) );
  AOI22_X1 U14013 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11698), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U14014 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11144), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U14015 ( .A1(n11485), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11656), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10909) );
  NAND4_X1 U14016 ( .A1(n10912), .A2(n10911), .A3(n10910), .A4(n10909), .ZN(
        n10913) );
  AOI22_X1 U14017 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11698), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10918) );
  AOI22_X1 U14018 ( .A1(n9680), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11072), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10917) );
  AOI22_X1 U14019 ( .A1(n10933), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U14020 ( .A1(n11485), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U14021 ( .A1(n10948), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11143), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U14022 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10921) );
  AOI22_X1 U14023 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10920) );
  INV_X2 U14024 ( .A(n14059), .ZN(n11700) );
  AOI22_X1 U14025 ( .A1(n11145), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10919) );
  AOI22_X1 U14026 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10926) );
  AOI22_X1 U14027 ( .A1(n11098), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11143), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10925) );
  AOI22_X1 U14028 ( .A1(n10948), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11144), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U14029 ( .A1(n10933), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11485), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10923) );
  NAND4_X1 U14030 ( .A1(n10926), .A2(n10925), .A3(n10924), .A4(n10923), .ZN(
        n10932) );
  AOI22_X1 U14031 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9674), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10930) );
  AOI22_X1 U14032 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U14033 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11072), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U14034 ( .A1(n10943), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9703), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10927) );
  NAND4_X1 U14035 ( .A1(n10930), .A2(n10928), .A3(n10929), .A4(n10927), .ZN(
        n10931) );
  OR2_X2 U14036 ( .A1(n10932), .A2(n10931), .ZN(n11001) );
  AOI22_X1 U14037 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11698), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U14038 ( .A1(n9680), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11072), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10936) );
  AOI22_X1 U14039 ( .A1(n10933), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11093), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10935) );
  AOI22_X1 U14040 ( .A1(n11485), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U14041 ( .A1(n10948), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11143), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U14042 ( .A1(n11098), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U14043 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10970), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U14044 ( .A1(n11145), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9703), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10939) );
  NAND2_X2 U14045 ( .A1(n9759), .A2(n10189), .ZN(n11033) );
  INV_X2 U14046 ( .A(n11033), .ZN(n11035) );
  INV_X1 U14047 ( .A(n11006), .ZN(n10965) );
  NAND2_X1 U14048 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10947) );
  NAND2_X1 U14049 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10946) );
  NAND2_X1 U14050 ( .A1(n10943), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10945) );
  NAND2_X1 U14051 ( .A1(n11072), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10944) );
  NAND2_X1 U14052 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10952) );
  NAND2_X1 U14053 ( .A1(n10948), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10951) );
  NAND2_X1 U14054 ( .A1(n11098), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10950) );
  NAND2_X1 U14055 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10949) );
  NAND2_X1 U14056 ( .A1(n10933), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10956) );
  NAND2_X1 U14057 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10955) );
  NAND2_X1 U14058 ( .A1(n11656), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10954) );
  NAND2_X1 U14059 ( .A1(n11485), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10953) );
  NAND2_X1 U14060 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10960) );
  NAND2_X1 U14061 ( .A1(n10970), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10959) );
  NAND2_X1 U14062 ( .A1(n11145), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10958) );
  NAND2_X1 U14063 ( .A1(n10938), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10957) );
  AOI22_X1 U14064 ( .A1(n10948), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11143), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10969) );
  AOI22_X1 U14065 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11406), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10968) );
  AOI22_X1 U14066 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11485), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10967) );
  AOI22_X1 U14067 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10966) );
  NAND4_X1 U14068 ( .A1(n10969), .A2(n10968), .A3(n10967), .A4(n10966), .ZN(
        n10976) );
  AOI22_X1 U14069 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11072), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10974) );
  AOI22_X1 U14070 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10973) );
  AOI22_X1 U14071 ( .A1(n10933), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11656), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10972) );
  AOI22_X1 U14072 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10971) );
  NAND4_X1 U14073 ( .A1(n10974), .A2(n10973), .A3(n10972), .A4(n10971), .ZN(
        n10975) );
  NAND2_X1 U14074 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10980) );
  NAND2_X1 U14075 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10979) );
  NAND2_X1 U14076 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10978) );
  NAND2_X1 U14077 ( .A1(n11072), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10977) );
  NAND2_X1 U14078 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10984) );
  NAND2_X1 U14079 ( .A1(n10948), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10983) );
  NAND2_X1 U14080 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10982) );
  NAND2_X1 U14081 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10981) );
  NAND2_X1 U14082 ( .A1(n10933), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10988) );
  NAND2_X1 U14083 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10987) );
  NAND2_X1 U14084 ( .A1(n11656), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10986) );
  NAND2_X1 U14085 ( .A1(n11485), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10985) );
  NAND2_X1 U14086 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10992) );
  NAND2_X1 U14087 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10991) );
  NAND2_X1 U14088 ( .A1(n11145), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10990) );
  NAND2_X1 U14089 ( .A1(n11700), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10989) );
  XNOR2_X1 U14090 ( .A(n10997), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n13375) );
  NAND2_X1 U14091 ( .A1(n13338), .A2(n13375), .ZN(n11111) );
  NAND2_X1 U14092 ( .A1(n11001), .A2(n9710), .ZN(n11003) );
  NAND2_X1 U14093 ( .A1(n11005), .A2(n11004), .ZN(n11007) );
  AND3_X2 U14094 ( .A1(n11008), .A2(n11007), .A3(n10177), .ZN(n13503) );
  INV_X1 U14095 ( .A(n13503), .ZN(n11048) );
  INV_X1 U14096 ( .A(n13812), .ZN(n11037) );
  NAND2_X1 U14097 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11012) );
  NAND2_X1 U14098 ( .A1(n11059), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11011) );
  NAND2_X1 U14099 ( .A1(n9680), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11010) );
  NAND2_X1 U14100 ( .A1(n11072), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11009) );
  NAND2_X1 U14101 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11016) );
  NAND2_X1 U14102 ( .A1(n10948), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11015) );
  NAND2_X1 U14103 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11014) );
  NAND2_X1 U14104 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11013) );
  NAND2_X1 U14105 ( .A1(n10933), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11020) );
  NAND2_X1 U14106 ( .A1(n11093), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11019) );
  NAND2_X1 U14107 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11018) );
  NAND2_X1 U14108 ( .A1(n11485), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11017) );
  NAND2_X1 U14109 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11025) );
  NAND2_X1 U14110 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11024) );
  NAND2_X1 U14111 ( .A1(n11145), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11023) );
  INV_X1 U14112 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11021) );
  NAND4_X4 U14113 ( .A1(n11029), .A2(n11028), .A3(n11027), .A4(n11026), .ZN(
        n13992) );
  NAND2_X1 U14114 ( .A1(n14060), .A2(n13596), .ZN(n11030) );
  NAND2_X1 U14115 ( .A1(n11743), .A2(n11001), .ZN(n11031) );
  OR2_X1 U14116 ( .A1(n11032), .A2(n11033), .ZN(n11034) );
  NAND2_X1 U14117 ( .A1(n13499), .A2(n15974), .ZN(n11040) );
  NAND2_X2 U14118 ( .A1(n13596), .A2(n13802), .ZN(n20910) );
  NAND2_X1 U14119 ( .A1(n11036), .A2(n13802), .ZN(n11720) );
  OAI211_X1 U14120 ( .C1(n11035), .C2(n20910), .A(n13611), .B(n11720), .ZN(
        n11053) );
  INV_X1 U14121 ( .A(n12342), .ZN(n11038) );
  NAND2_X1 U14122 ( .A1(n11037), .A2(n13802), .ZN(n11807) );
  NAND2_X1 U14123 ( .A1(n11807), .A2(n11803), .ZN(n11784) );
  NOR2_X1 U14124 ( .A1(n11053), .A2(n11723), .ZN(n11039) );
  AND4_X2 U14125 ( .A1(n11111), .A2(n11039), .A3(n11040), .A4(n11041), .ZN(
        n11043) );
  NOR2_X1 U14126 ( .A1(n9699), .A2(n13802), .ZN(n11042) );
  INV_X1 U14127 ( .A(n12441), .ZN(n11044) );
  MUX2_X1 U14128 ( .A(n20804), .B(n11044), .S(n14105), .Z(n11045) );
  INV_X1 U14129 ( .A(n13371), .ZN(n13987) );
  NAND3_X1 U14130 ( .A1(n13987), .A2(n11032), .A3(n13812), .ZN(n11047) );
  NAND2_X1 U14131 ( .A1(n11048), .A2(n11047), .ZN(n11057) );
  NAND2_X1 U14132 ( .A1(n13989), .A2(n13992), .ZN(n13984) );
  NOR2_X1 U14133 ( .A1(n20897), .A2(n20222), .ZN(n11049) );
  AND2_X1 U14134 ( .A1(n13984), .A2(n11049), .ZN(n11051) );
  NAND2_X1 U14135 ( .A1(n11780), .A2(n11050), .ZN(n13609) );
  OAI211_X1 U14136 ( .C1(n11052), .C2(n20910), .A(n11051), .B(n13609), .ZN(
        n11054) );
  NOR2_X1 U14137 ( .A1(n11054), .A2(n11053), .ZN(n11056) );
  NAND3_X1 U14138 ( .A1(n13499), .A2(n13992), .A3(n15974), .ZN(n11055) );
  NAND3_X1 U14139 ( .A1(n11057), .A2(n11056), .A3(n11055), .ZN(n11114) );
  INV_X1 U14140 ( .A(n11114), .ZN(n11058) );
  AOI22_X1 U14141 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11675), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11064) );
  AOI22_X1 U14142 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11063) );
  AOI22_X1 U14143 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11062) );
  AOI22_X1 U14144 ( .A1(n11485), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11656), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11061) );
  NAND4_X1 U14145 ( .A1(n11064), .A2(n11063), .A3(n11062), .A4(n11061), .ZN(
        n11071) );
  BUF_X1 U14146 ( .A(n11143), .Z(n11065) );
  AOI22_X1 U14147 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11069) );
  AOI22_X1 U14148 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11068) );
  AOI22_X1 U14149 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11067) );
  INV_X1 U14150 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n20396) );
  AOI22_X1 U14151 ( .A1(n11145), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11066) );
  NAND4_X1 U14152 ( .A1(n11069), .A2(n11068), .A3(n11067), .A4(n11066), .ZN(
        n11070) );
  NOR2_X1 U14153 ( .A1(n11191), .A2(n12404), .ZN(n11092) );
  BUF_X1 U14154 ( .A(n9679), .Z(n11543) );
  AOI22_X1 U14155 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n11543), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11076) );
  AOI22_X1 U14156 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n11065), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11075) );
  AOI22_X1 U14157 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n9711), .B1(n9706), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11074) );
  AOI22_X1 U14158 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11656), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11073) );
  NAND4_X1 U14159 ( .A1(n11076), .A2(n11075), .A3(n11074), .A4(n11073), .ZN(
        n11083) );
  AOI22_X1 U14160 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11698), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11081) );
  BUF_X1 U14161 ( .A(n11144), .Z(n11077) );
  AOI22_X1 U14162 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n9686), .B1(
        n11077), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11080) );
  AOI22_X1 U14163 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11485), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11079) );
  AOI22_X1 U14164 ( .A1(n11145), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11078) );
  NAND4_X1 U14165 ( .A1(n11081), .A2(n11080), .A3(n11079), .A4(n11078), .ZN(
        n11082) );
  MUX2_X1 U14166 ( .A(n11090), .B(n11092), .S(n12341), .Z(n11084) );
  INV_X1 U14167 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20376) );
  INV_X1 U14168 ( .A(n11087), .ZN(n11746) );
  OAI21_X1 U14169 ( .B1(n20222), .B2(n12341), .A(n11746), .ZN(n11088) );
  NAND2_X1 U14170 ( .A1(n11169), .A2(n11170), .ZN(n11091) );
  INV_X1 U14171 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20379) );
  OR2_X1 U14172 ( .A1(n11762), .A2(n20379), .ZN(n11108) );
  INV_X1 U14173 ( .A(n11092), .ZN(n11107) );
  AOI22_X1 U14174 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11097) );
  AOI22_X1 U14175 ( .A1(n11675), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11096) );
  AOI22_X1 U14176 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11077), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11095) );
  AOI22_X1 U14177 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11485), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11094) );
  NAND4_X1 U14178 ( .A1(n11097), .A2(n11096), .A3(n11095), .A4(n11094), .ZN(
        n11105) );
  AOI22_X1 U14179 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11103) );
  AOI22_X1 U14180 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11102) );
  AOI22_X1 U14181 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11101) );
  AOI22_X1 U14182 ( .A1(n11099), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11100) );
  NAND4_X1 U14183 ( .A1(n11103), .A2(n11102), .A3(n11101), .A4(n11100), .ZN(
        n11104) );
  OR2_X1 U14184 ( .A1(n11190), .A2(n11118), .ZN(n11106) );
  NAND2_X1 U14185 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11130) );
  OAI21_X1 U14186 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n11130), .ZN(n20574) );
  NAND2_X1 U14187 ( .A1(n20804), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11124) );
  OAI21_X1 U14188 ( .B1(n12441), .B2(n20574), .A(n11124), .ZN(n11109) );
  INV_X1 U14189 ( .A(n11109), .ZN(n11110) );
  INV_X1 U14190 ( .A(n9700), .ZN(n11113) );
  AND2_X1 U14191 ( .A1(n11001), .A2(n13384), .ZN(n11934) );
  NAND4_X1 U14192 ( .A1(n11780), .A2(n13371), .A3(n11743), .A4(n11934), .ZN(
        n13620) );
  NAND2_X1 U14193 ( .A1(n11111), .A2(n13620), .ZN(n11112) );
  INV_X1 U14194 ( .A(n11116), .ZN(n11117) );
  NAND2_X1 U14195 ( .A1(n11128), .A2(n13795), .ZN(n14091) );
  OR2_X1 U14196 ( .A1(n11191), .A2(n11118), .ZN(n11119) );
  AND2_X2 U14197 ( .A1(n9773), .A2(n11119), .ZN(n12339) );
  INV_X1 U14198 ( .A(n11120), .ZN(n11121) );
  INV_X1 U14199 ( .A(n11183), .ZN(n11155) );
  AND2_X1 U14200 ( .A1(n11124), .A2(n10901), .ZN(n11125) );
  INV_X1 U14201 ( .A(n11130), .ZN(n11129) );
  NAND2_X1 U14202 ( .A1(n11129), .A2(n11729), .ZN(n20662) );
  NAND2_X1 U14203 ( .A1(n11130), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11131) );
  AND2_X1 U14204 ( .A1(n20662), .A2(n11131), .ZN(n14204) );
  NAND2_X1 U14205 ( .A1(n20804), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11134) );
  NAND2_X1 U14206 ( .A1(n11138), .A2(n14079), .ZN(n13495) );
  AOI22_X1 U14207 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11698), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11142) );
  AOI22_X1 U14208 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11141) );
  AOI22_X1 U14209 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11140) );
  AOI22_X1 U14210 ( .A1(n11485), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11139) );
  NAND4_X1 U14211 ( .A1(n11142), .A2(n11141), .A3(n11140), .A4(n11139), .ZN(
        n11151) );
  AOI22_X1 U14212 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11149) );
  AOI22_X1 U14213 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11148) );
  AOI22_X1 U14214 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11147) );
  AOI22_X1 U14215 ( .A1(n11099), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11146) );
  NAND4_X1 U14216 ( .A1(n11149), .A2(n11148), .A3(n11147), .A4(n11146), .ZN(
        n11150) );
  INV_X1 U14217 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20382) );
  OAI22_X1 U14218 ( .A1(n11762), .A2(n20382), .B1(n11190), .B2(n12331), .ZN(
        n11152) );
  INV_X1 U14219 ( .A(n11152), .ZN(n11153) );
  NAND2_X1 U14220 ( .A1(n12329), .A2(n11396), .ZN(n11160) );
  NAND2_X1 U14221 ( .A1(n11934), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11213) );
  XNOR2_X1 U14222 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20305) );
  NAND2_X1 U14223 ( .A1(n20806), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11340) );
  AOI21_X1 U14224 ( .B1(n13980), .B2(n20305), .A(n13843), .ZN(n11157) );
  NAND2_X1 U14225 ( .A1(n11497), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11156) );
  OAI211_X1 U14226 ( .C1(n11213), .C2(n11133), .A(n11157), .B(n11156), .ZN(
        n11158) );
  INV_X1 U14227 ( .A(n11158), .ZN(n11159) );
  NAND2_X1 U14228 ( .A1(n11160), .A2(n11159), .ZN(n11161) );
  NAND2_X1 U14229 ( .A1(n13843), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11182) );
  NAND2_X1 U14230 ( .A1(n11161), .A2(n11182), .ZN(n13697) );
  INV_X1 U14231 ( .A(n13697), .ZN(n11181) );
  NAND2_X1 U14232 ( .A1(n9715), .A2(n11396), .ZN(n11168) );
  AOI22_X1 U14233 ( .A1(n11497), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20806), .ZN(n11166) );
  INV_X1 U14234 ( .A(n11213), .ZN(n11228) );
  NAND2_X1 U14235 ( .A1(n11228), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11165) );
  AND2_X1 U14236 ( .A1(n11166), .A2(n11165), .ZN(n11167) );
  NAND2_X1 U14237 ( .A1(n11168), .A2(n11167), .ZN(n13562) );
  NAND2_X1 U14238 ( .A1(n14237), .A2(n11050), .ZN(n11171) );
  NAND2_X1 U14239 ( .A1(n11171), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13487) );
  NAND2_X1 U14240 ( .A1(n11173), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11175) );
  NAND2_X1 U14241 ( .A1(n20806), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11174) );
  OAI211_X1 U14242 ( .C1(n11213), .C2(n10900), .A(n11175), .B(n11174), .ZN(
        n11176) );
  AOI21_X1 U14243 ( .B1(n11172), .B2(n11396), .A(n11176), .ZN(n13488) );
  OR2_X1 U14244 ( .A1(n13487), .A2(n13488), .ZN(n13485) );
  INV_X1 U14245 ( .A(n13488), .ZN(n11178) );
  OR2_X1 U14246 ( .A1(n11178), .A2(n11177), .ZN(n11179) );
  NAND2_X1 U14247 ( .A1(n13485), .A2(n11179), .ZN(n13561) );
  NAND2_X1 U14248 ( .A1(n13562), .A2(n13561), .ZN(n13696) );
  NAND2_X1 U14249 ( .A1(n11181), .A2(n11180), .ZN(n13694) );
  NAND3_X1 U14250 ( .A1(n20661), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20547) );
  INV_X1 U14251 ( .A(n20547), .ZN(n11185) );
  NAND2_X1 U14252 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11185), .ZN(
        n20542) );
  NAND2_X1 U14253 ( .A1(n20661), .A2(n20542), .ZN(n11186) );
  NAND3_X1 U14254 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20741) );
  INV_X1 U14255 ( .A(n20741), .ZN(n20749) );
  NAND2_X1 U14256 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20749), .ZN(
        n20742) );
  NAND2_X1 U14257 ( .A1(n11186), .A2(n20742), .ZN(n20573) );
  OAI22_X1 U14258 ( .A1(n12441), .A2(n20573), .B1(n16008), .B2(n20661), .ZN(
        n11187) );
  INV_X1 U14259 ( .A(n11187), .ZN(n11188) );
  AOI22_X1 U14260 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11675), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11195) );
  AOI22_X1 U14261 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11194) );
  AOI22_X1 U14262 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11656), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11193) );
  AOI22_X1 U14263 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11099), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11192) );
  NAND4_X1 U14264 ( .A1(n11195), .A2(n11194), .A3(n11193), .A4(n11192), .ZN(
        n11201) );
  AOI22_X1 U14265 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11199) );
  AOI22_X1 U14266 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11077), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11198) );
  AOI22_X1 U14267 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11197) );
  AOI22_X1 U14268 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11196) );
  NAND4_X1 U14269 ( .A1(n11199), .A2(n11198), .A3(n11197), .A4(n11196), .ZN(
        n11200) );
  AOI22_X1 U14270 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11768), .B1(
        n11740), .B2(n12361), .ZN(n11202) );
  INV_X1 U14271 ( .A(n11204), .ZN(n11205) );
  INV_X1 U14272 ( .A(n13841), .ZN(n13903) );
  NAND2_X1 U14273 ( .A1(n11205), .A2(n13903), .ZN(n11206) );
  NAND2_X1 U14274 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11208) );
  INV_X1 U14275 ( .A(n11208), .ZN(n11210) );
  INV_X1 U14276 ( .A(n11231), .ZN(n11209) );
  OAI21_X1 U14277 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11210), .A(
        n11209), .ZN(n14131) );
  AOI22_X1 U14278 ( .A1(n13980), .A2(n14131), .B1(n13843), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11212) );
  NAND2_X1 U14279 ( .A1(n11497), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11211) );
  OAI211_X1 U14280 ( .C1(n11213), .C2(n14074), .A(n11212), .B(n11211), .ZN(
        n11214) );
  INV_X1 U14281 ( .A(n11214), .ZN(n11215) );
  OAI21_X1 U14282 ( .B1(n15112), .B2(n11420), .A(n11215), .ZN(n13644) );
  NAND2_X1 U14283 ( .A1(n13645), .A2(n13644), .ZN(n13642) );
  INV_X1 U14284 ( .A(n13642), .ZN(n11237) );
  AOI22_X1 U14285 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11675), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11219) );
  AOI22_X1 U14286 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11218) );
  AOI22_X1 U14287 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11217) );
  AOI22_X1 U14288 ( .A1(n11527), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11656), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11216) );
  NAND4_X1 U14289 ( .A1(n11219), .A2(n11218), .A3(n11217), .A4(n11216), .ZN(
        n11225) );
  AOI22_X1 U14290 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11223) );
  AOI22_X1 U14291 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11222) );
  AOI22_X1 U14292 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11221) );
  INV_X1 U14293 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n20388) );
  AOI22_X1 U14294 ( .A1(n11099), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11220) );
  NAND4_X1 U14295 ( .A1(n11223), .A2(n11222), .A3(n11221), .A4(n11220), .ZN(
        n11224) );
  NAND2_X1 U14296 ( .A1(n11740), .A2(n12365), .ZN(n11227) );
  OR2_X1 U14297 ( .A1(n11762), .A2(n20388), .ZN(n11226) );
  XNOR2_X1 U14298 ( .A(n9763), .B(n11238), .ZN(n12360) );
  NAND2_X1 U14299 ( .A1(n11228), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11234) );
  INV_X1 U14300 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11229) );
  AOI21_X1 U14301 ( .B1(n11229), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11230) );
  AOI21_X1 U14302 ( .B1(n11497), .B2(P1_EAX_REG_4__SCAN_IN), .A(n11230), .ZN(
        n11233) );
  NOR2_X1 U14303 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n11231), .ZN(
        n11232) );
  NOR2_X1 U14304 ( .A1(n11254), .A2(n11232), .ZN(n13930) );
  AOI22_X1 U14305 ( .A1(n11234), .A2(n11233), .B1(n13980), .B2(n13930), .ZN(
        n11235) );
  AOI21_X1 U14306 ( .B1(n12360), .B2(n11396), .A(n11235), .ZN(n13790) );
  NAND2_X1 U14307 ( .A1(n11237), .A2(n11236), .ZN(n13789) );
  AOI22_X1 U14308 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11675), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11242) );
  AOI22_X1 U14309 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11241) );
  AOI22_X1 U14310 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9686), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11240) );
  AOI22_X1 U14311 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11239) );
  NAND4_X1 U14312 ( .A1(n11242), .A2(n11241), .A3(n11240), .A4(n11239), .ZN(
        n11248) );
  AOI22_X1 U14313 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11246) );
  AOI22_X1 U14314 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11245) );
  AOI22_X1 U14315 ( .A1(n11527), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11244) );
  AOI22_X1 U14316 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11099), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11243) );
  NAND4_X1 U14317 ( .A1(n11246), .A2(n11245), .A3(n11244), .A4(n11243), .ZN(
        n11247) );
  NAND2_X1 U14318 ( .A1(n11740), .A2(n12382), .ZN(n11250) );
  INV_X1 U14319 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14323) );
  OR2_X1 U14320 ( .A1(n11762), .A2(n14323), .ZN(n11249) );
  NAND2_X1 U14321 ( .A1(n11252), .A2(n11251), .ZN(n11253) );
  INV_X1 U14322 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11259) );
  INV_X1 U14323 ( .A(n11285), .ZN(n11257) );
  INV_X1 U14324 ( .A(n11254), .ZN(n11255) );
  INV_X1 U14325 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16188) );
  NAND2_X1 U14326 ( .A1(n11255), .A2(n16188), .ZN(n11256) );
  NAND2_X1 U14327 ( .A1(n11257), .A2(n11256), .ZN(n20282) );
  AOI22_X1 U14328 ( .A1(n20282), .A2(n13980), .B1(n13843), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11258) );
  OAI21_X1 U14329 ( .B1(n11403), .B2(n11259), .A(n11258), .ZN(n11260) );
  NAND2_X1 U14330 ( .A1(n11262), .A2(n11261), .ZN(n14106) );
  NAND2_X1 U14331 ( .A1(n11768), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11274) );
  AOI22_X1 U14332 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11675), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11266) );
  AOI22_X1 U14333 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11265) );
  AOI22_X1 U14334 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11264) );
  AOI22_X1 U14335 ( .A1(n11527), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11656), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11263) );
  NAND4_X1 U14336 ( .A1(n11266), .A2(n11265), .A3(n11264), .A4(n11263), .ZN(
        n11272) );
  AOI22_X1 U14337 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11270) );
  AOI22_X1 U14338 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11269) );
  AOI22_X1 U14339 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11268) );
  INV_X1 U14340 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20391) );
  AOI22_X1 U14341 ( .A1(n11099), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11267) );
  NAND4_X1 U14342 ( .A1(n11270), .A2(n11269), .A3(n11268), .A4(n11267), .ZN(
        n11271) );
  NAND2_X1 U14343 ( .A1(n11740), .A2(n12392), .ZN(n11273) );
  NAND2_X1 U14344 ( .A1(n11281), .A2(n11280), .ZN(n12380) );
  NAND2_X1 U14345 ( .A1(n12380), .A2(n11396), .ZN(n11279) );
  XNOR2_X1 U14346 ( .A(n11285), .B(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n20272) );
  NAND2_X1 U14347 ( .A1(n20272), .A2(n13980), .ZN(n11276) );
  NAND2_X1 U14348 ( .A1(n13843), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11275) );
  NAND2_X1 U14349 ( .A1(n11276), .A2(n11275), .ZN(n11277) );
  AOI21_X1 U14350 ( .B1(n11497), .B2(P1_EAX_REG_6__SCAN_IN), .A(n11277), .ZN(
        n11278) );
  NAND2_X1 U14351 ( .A1(n11740), .A2(n12404), .ZN(n11282) );
  OAI21_X1 U14352 ( .B1(n20396), .B2(n11762), .A(n11282), .ZN(n11283) );
  NAND2_X1 U14353 ( .A1(n12390), .A2(n11396), .ZN(n11292) );
  INV_X1 U14354 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20253) );
  INV_X1 U14355 ( .A(n11308), .ZN(n11288) );
  NAND2_X1 U14356 ( .A1(n11285), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11286) );
  NAND2_X1 U14357 ( .A1(n11286), .A2(n20253), .ZN(n11287) );
  NAND2_X1 U14358 ( .A1(n11288), .A2(n11287), .ZN(n20264) );
  NAND2_X1 U14359 ( .A1(n20264), .A2(n13980), .ZN(n11289) );
  OAI21_X1 U14360 ( .B1(n20253), .B2(n11340), .A(n11289), .ZN(n11290) );
  AOI21_X1 U14361 ( .B1(n11497), .B2(P1_EAX_REG_7__SCAN_IN), .A(n11290), .ZN(
        n11291) );
  NAND2_X1 U14362 ( .A1(n11292), .A2(n11291), .ZN(n14151) );
  AOI22_X1 U14363 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11297) );
  AOI22_X1 U14364 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n9711), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11296) );
  AOI22_X1 U14365 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n9686), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11295) );
  AOI22_X1 U14366 ( .A1(n11060), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11099), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11294) );
  NAND4_X1 U14367 ( .A1(n11297), .A2(n11296), .A3(n11295), .A4(n11294), .ZN(
        n11303) );
  AOI22_X1 U14368 ( .A1(n11675), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U14369 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n11077), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11300) );
  AOI22_X1 U14370 ( .A1(n11527), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11656), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11299) );
  AOI22_X1 U14371 ( .A1(n9680), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11298) );
  NAND4_X1 U14372 ( .A1(n11301), .A2(n11300), .A3(n11299), .A4(n11298), .ZN(
        n11302) );
  OAI21_X1 U14373 ( .B1(n11303), .B2(n11302), .A(n11396), .ZN(n11307) );
  NAND2_X1 U14374 ( .A1(n11497), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11306) );
  NAND2_X1 U14375 ( .A1(n13843), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11305) );
  XNOR2_X1 U14376 ( .A(n11308), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14392) );
  NAND2_X1 U14377 ( .A1(n14392), .A2(n13980), .ZN(n11304) );
  NAND4_X1 U14378 ( .A1(n11307), .A2(n11306), .A3(n11305), .A4(n11304), .ZN(
        n14277) );
  XNOR2_X1 U14379 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n11333), .ZN(
        n20246) );
  AOI22_X1 U14380 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11675), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11312) );
  AOI22_X1 U14381 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11311) );
  AOI22_X1 U14382 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11656), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11310) );
  AOI22_X1 U14383 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11099), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11309) );
  NAND4_X1 U14384 ( .A1(n11312), .A2(n11311), .A3(n11310), .A4(n11309), .ZN(
        n11318) );
  AOI22_X1 U14385 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11316) );
  AOI22_X1 U14386 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11077), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11315) );
  AOI22_X1 U14387 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11314) );
  AOI22_X1 U14388 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11313) );
  NAND4_X1 U14389 ( .A1(n11316), .A2(n11315), .A3(n11314), .A4(n11313), .ZN(
        n11317) );
  OR2_X1 U14390 ( .A1(n11318), .A2(n11317), .ZN(n11319) );
  AOI22_X1 U14391 ( .A1(n11396), .A2(n11319), .B1(n13843), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11321) );
  NAND2_X1 U14392 ( .A1(n11497), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11320) );
  OAI211_X1 U14393 ( .C1(n20246), .C2(n11177), .A(n11321), .B(n11320), .ZN(
        n14324) );
  AOI22_X1 U14394 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11675), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14395 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U14396 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11323) );
  AOI22_X1 U14397 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11322) );
  NAND4_X1 U14398 ( .A1(n11325), .A2(n11324), .A3(n11323), .A4(n11322), .ZN(
        n11331) );
  AOI22_X1 U14399 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11329) );
  AOI22_X1 U14400 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11328) );
  AOI22_X1 U14401 ( .A1(n11527), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11327) );
  AOI22_X1 U14402 ( .A1(n11099), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11326) );
  NAND4_X1 U14403 ( .A1(n11329), .A2(n11328), .A3(n11327), .A4(n11326), .ZN(
        n11330) );
  NOR2_X1 U14404 ( .A1(n11331), .A2(n11330), .ZN(n11336) );
  XNOR2_X1 U14405 ( .A(n11337), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14929) );
  NAND2_X1 U14406 ( .A1(n14929), .A2(n13980), .ZN(n11335) );
  AOI22_X1 U14407 ( .A1(n11497), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n13843), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11334) );
  OAI211_X1 U14408 ( .C1(n11336), .C2(n11420), .A(n11335), .B(n11334), .ZN(
        n14376) );
  INV_X1 U14409 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11341) );
  OAI21_X1 U14410 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11338), .A(
        n11399), .ZN(n16166) );
  NAND2_X1 U14411 ( .A1(n16166), .A2(n13980), .ZN(n11339) );
  OAI21_X1 U14412 ( .B1(n11341), .B2(n11340), .A(n11339), .ZN(n11342) );
  AOI21_X1 U14413 ( .B1(n11497), .B2(P1_EAX_REG_11__SCAN_IN), .A(n11342), .ZN(
        n11343) );
  INV_X1 U14414 ( .A(n11343), .ZN(n14453) );
  NAND2_X1 U14415 ( .A1(n14451), .A2(n14453), .ZN(n14452) );
  INV_X1 U14416 ( .A(n14375), .ZN(n11356) );
  AOI22_X1 U14417 ( .A1(n11060), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11347) );
  AOI22_X1 U14418 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11346) );
  AOI22_X1 U14419 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11144), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11345) );
  AOI22_X1 U14420 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11656), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11344) );
  NAND4_X1 U14421 ( .A1(n11347), .A2(n11346), .A3(n11345), .A4(n11344), .ZN(
        n11353) );
  AOI22_X1 U14422 ( .A1(n11675), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11543), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11351) );
  AOI22_X1 U14423 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U14424 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11349) );
  AOI22_X1 U14425 ( .A1(n11145), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11348) );
  NAND4_X1 U14426 ( .A1(n11351), .A2(n11350), .A3(n11349), .A4(n11348), .ZN(
        n11352) );
  OR2_X1 U14427 ( .A1(n11353), .A2(n11352), .ZN(n11354) );
  NAND2_X1 U14428 ( .A1(n11396), .A2(n11354), .ZN(n14476) );
  INV_X1 U14429 ( .A(n14476), .ZN(n11355) );
  INV_X1 U14430 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11358) );
  XNOR2_X1 U14431 ( .A(n11405), .B(n11358), .ZN(n14910) );
  AOI22_X1 U14432 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11543), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U14433 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11361) );
  AOI22_X1 U14434 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11360) );
  AOI22_X1 U14435 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11359) );
  NAND4_X1 U14436 ( .A1(n11362), .A2(n11361), .A3(n11360), .A4(n11359), .ZN(
        n11368) );
  AOI22_X1 U14437 ( .A1(n11675), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11366) );
  AOI22_X1 U14438 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11077), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11365) );
  AOI22_X1 U14439 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U14440 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11099), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11363) );
  NAND4_X1 U14441 ( .A1(n11366), .A2(n11365), .A3(n11364), .A4(n11363), .ZN(
        n11367) );
  NOR2_X1 U14442 ( .A1(n11368), .A2(n11367), .ZN(n11371) );
  NAND2_X1 U14443 ( .A1(n11497), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11370) );
  NAND2_X1 U14444 ( .A1(n13843), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11369) );
  OAI211_X1 U14445 ( .C1(n11420), .C2(n11371), .A(n11370), .B(n11369), .ZN(
        n11372) );
  AOI21_X1 U14446 ( .B1(n14910), .B2(n13980), .A(n11372), .ZN(n11373) );
  INV_X1 U14447 ( .A(n11373), .ZN(n14439) );
  XOR2_X1 U14448 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11374), .Z(
        n16096) );
  AOI22_X1 U14449 ( .A1(n11675), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U14450 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11377) );
  AOI22_X1 U14451 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11376) );
  AOI22_X1 U14452 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11099), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11375) );
  NAND4_X1 U14453 ( .A1(n11378), .A2(n11377), .A3(n11376), .A4(n11375), .ZN(
        n11384) );
  AOI22_X1 U14454 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11382) );
  AOI22_X1 U14455 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11381) );
  AOI22_X1 U14456 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11380) );
  AOI22_X1 U14457 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11379) );
  NAND4_X1 U14458 ( .A1(n11382), .A2(n11381), .A3(n11380), .A4(n11379), .ZN(
        n11383) );
  OR2_X1 U14459 ( .A1(n11384), .A2(n11383), .ZN(n11385) );
  AOI22_X1 U14460 ( .A1(n11396), .A2(n11385), .B1(n13843), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11387) );
  NAND2_X1 U14461 ( .A1(n11497), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11386) );
  OAI211_X1 U14462 ( .C1(n16096), .C2(n11177), .A(n11387), .B(n11386), .ZN(
        n14455) );
  INV_X1 U14463 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14488) );
  AOI22_X1 U14464 ( .A1(n11675), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14465 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11077), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11390) );
  AOI22_X1 U14466 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11389) );
  AOI22_X1 U14467 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11388) );
  NAND4_X1 U14468 ( .A1(n11391), .A2(n11390), .A3(n11389), .A4(n11388), .ZN(
        n11398) );
  AOI22_X1 U14469 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14470 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11394) );
  AOI22_X1 U14471 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14472 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11099), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11392) );
  NAND4_X1 U14473 ( .A1(n11395), .A2(n11394), .A3(n11393), .A4(n11392), .ZN(
        n11397) );
  OAI21_X1 U14474 ( .B1(n11398), .B2(n11397), .A(n11396), .ZN(n11402) );
  XNOR2_X1 U14475 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11399), .ZN(
        n16154) );
  INV_X1 U14476 ( .A(n16154), .ZN(n11400) );
  AOI22_X1 U14477 ( .A1(n13843), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n13980), .B2(n11400), .ZN(n11401) );
  OAI211_X1 U14478 ( .C1(n11403), .C2(n14488), .A(n11402), .B(n11401), .ZN(
        n14484) );
  AND2_X1 U14479 ( .A1(n14455), .A2(n14484), .ZN(n14435) );
  NAND2_X1 U14480 ( .A1(n14436), .A2(n11404), .ZN(n14437) );
  XOR2_X1 U14481 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n11423), .Z(
        n16148) );
  INV_X1 U14482 ( .A(n16148), .ZN(n11422) );
  AOI22_X1 U14483 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11675), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14484 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11409) );
  AOI22_X1 U14485 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11408) );
  AOI22_X1 U14486 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11407) );
  NAND4_X1 U14487 ( .A1(n11410), .A2(n11409), .A3(n11408), .A4(n11407), .ZN(
        n11416) );
  AOI22_X1 U14488 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14489 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11413) );
  AOI22_X1 U14490 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11412) );
  AOI22_X1 U14491 ( .A1(n11099), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11411) );
  NAND4_X1 U14492 ( .A1(n11414), .A2(n11413), .A3(n11412), .A4(n11411), .ZN(
        n11415) );
  NOR2_X1 U14493 ( .A1(n11416), .A2(n11415), .ZN(n11419) );
  NAND2_X1 U14494 ( .A1(n11497), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11418) );
  NAND2_X1 U14495 ( .A1(n13843), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11417) );
  OAI211_X1 U14496 ( .C1(n11420), .C2(n11419), .A(n11418), .B(n11417), .ZN(
        n11421) );
  AOI21_X1 U14497 ( .B1(n11422), .B2(n13980), .A(n11421), .ZN(n14463) );
  NAND2_X1 U14498 ( .A1(n11423), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11437) );
  XNOR2_X1 U14499 ( .A(n11437), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16143) );
  AOI21_X1 U14500 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14690), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11424) );
  AOI21_X1 U14501 ( .B1(n11497), .B2(P1_EAX_REG_16__SCAN_IN), .A(n11424), .ZN(
        n11436) );
  AOI22_X1 U14502 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U14503 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14504 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n11522), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11426) );
  AOI22_X1 U14505 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n9706), .B1(
        n11077), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11425) );
  NAND4_X1 U14506 ( .A1(n11428), .A2(n11427), .A3(n11426), .A4(n11425), .ZN(
        n11434) );
  AOI22_X1 U14507 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11675), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11432) );
  AOI22_X1 U14508 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n9711), .B1(
        n11633), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U14509 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n11527), .B1(
        n11656), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11430) );
  AOI22_X1 U14510 ( .A1(n11099), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11429) );
  NAND4_X1 U14511 ( .A1(n11432), .A2(n11431), .A3(n11430), .A4(n11429), .ZN(
        n11433) );
  OAI21_X1 U14512 ( .B1(n11434), .B2(n11433), .A(n11713), .ZN(n11435) );
  AOI22_X1 U14513 ( .A1(n16143), .A2(n13980), .B1(n11436), .B2(n11435), .ZN(
        n14686) );
  XNOR2_X1 U14514 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11452), .ZN(
        n16139) );
  INV_X1 U14515 ( .A(n16139), .ZN(n11451) );
  AOI22_X1 U14516 ( .A1(n11675), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11543), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U14517 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11440) );
  AOI22_X1 U14518 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11077), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11439) );
  AOI22_X1 U14519 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11438) );
  NAND4_X1 U14520 ( .A1(n11441), .A2(n11440), .A3(n11439), .A4(n11438), .ZN(
        n11447) );
  AOI22_X1 U14521 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11445) );
  AOI22_X1 U14522 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11444) );
  AOI22_X1 U14523 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11656), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11443) );
  AOI22_X1 U14524 ( .A1(n11099), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11442) );
  NAND4_X1 U14525 ( .A1(n11445), .A2(n11444), .A3(n11443), .A4(n11442), .ZN(
        n11446) );
  NOR2_X1 U14526 ( .A1(n11447), .A2(n11446), .ZN(n11449) );
  AOI22_X1 U14527 ( .A1(n11497), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n13843), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11448) );
  OAI21_X1 U14528 ( .B1(n11688), .B2(n11449), .A(n11448), .ZN(n11450) );
  AOI21_X1 U14529 ( .B1(n11451), .B2(n13980), .A(n11450), .ZN(n14732) );
  XNOR2_X1 U14530 ( .A(n11481), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14899) );
  AOI22_X1 U14531 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11456) );
  AOI22_X1 U14532 ( .A1(n11675), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11455) );
  AOI22_X1 U14533 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11656), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U14534 ( .A1(n11060), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11453) );
  NAND4_X1 U14535 ( .A1(n11456), .A2(n11455), .A3(n11454), .A4(n11453), .ZN(
        n11462) );
  AOI22_X1 U14536 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14537 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11459) );
  AOI22_X1 U14538 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11458) );
  AOI22_X1 U14539 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11457) );
  NAND4_X1 U14540 ( .A1(n11460), .A2(n11459), .A3(n11458), .A4(n11457), .ZN(
        n11461) );
  OAI21_X1 U14541 ( .B1(n11462), .B2(n11461), .A(n11713), .ZN(n11464) );
  AOI22_X1 U14542 ( .A1(n11497), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n20806), .ZN(n11463) );
  AOI21_X1 U14543 ( .B1(n11464), .B2(n11463), .A(n13980), .ZN(n11465) );
  AOI21_X1 U14544 ( .B1(n14899), .B2(n13980), .A(n11465), .ZN(n14678) );
  AOI22_X1 U14545 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11470) );
  AOI22_X1 U14546 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11633), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11469) );
  AOI22_X1 U14547 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11468) );
  AOI22_X1 U14548 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11467) );
  NAND4_X1 U14549 ( .A1(n11470), .A2(n11469), .A3(n11468), .A4(n11467), .ZN(
        n11476) );
  AOI22_X1 U14550 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11675), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U14551 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11473) );
  AOI22_X1 U14552 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11472) );
  AOI22_X1 U14553 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11099), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11471) );
  NAND4_X1 U14554 ( .A1(n11474), .A2(n11473), .A3(n11472), .A4(n11471), .ZN(
        n11475) );
  NOR2_X1 U14555 ( .A1(n11476), .A2(n11475), .ZN(n11480) );
  NAND2_X1 U14556 ( .A1(n20806), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11477) );
  NAND2_X1 U14557 ( .A1(n11177), .A2(n11477), .ZN(n11478) );
  AOI21_X1 U14558 ( .B1(n11497), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11478), .ZN(
        n11479) );
  OAI21_X1 U14559 ( .B1(n11688), .B2(n11480), .A(n11479), .ZN(n11484) );
  OAI21_X1 U14560 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n11482), .A(
        n11516), .ZN(n16125) );
  OR2_X1 U14561 ( .A1(n11177), .A2(n16125), .ZN(n11483) );
  AOI22_X1 U14562 ( .A1(n11675), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11543), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11489) );
  AOI22_X1 U14563 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9686), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11488) );
  AOI22_X1 U14564 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11487) );
  AOI22_X1 U14565 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11486) );
  NAND4_X1 U14566 ( .A1(n11489), .A2(n11488), .A3(n11487), .A4(n11486), .ZN(
        n11495) );
  AOI22_X1 U14567 ( .A1(n11060), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11493) );
  AOI22_X1 U14568 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11492) );
  AOI22_X1 U14569 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11656), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U14570 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11099), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11490) );
  NAND4_X1 U14571 ( .A1(n11493), .A2(n11492), .A3(n11491), .A4(n11490), .ZN(
        n11494) );
  NOR2_X1 U14572 ( .A1(n11495), .A2(n11494), .ZN(n11499) );
  INV_X1 U14573 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14889) );
  AOI21_X1 U14574 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14889), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11496) );
  AOI21_X1 U14575 ( .B1(n11497), .B2(P1_EAX_REG_20__SCAN_IN), .A(n11496), .ZN(
        n11498) );
  OAI21_X1 U14576 ( .B1(n11688), .B2(n11499), .A(n11498), .ZN(n11501) );
  XNOR2_X1 U14577 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n11516), .ZN(
        n14891) );
  NAND2_X1 U14578 ( .A1(n13980), .A2(n14891), .ZN(n11500) );
  AOI22_X1 U14579 ( .A1(n11675), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11543), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U14580 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U14581 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U14582 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11099), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11502) );
  NAND4_X1 U14583 ( .A1(n11505), .A2(n11504), .A3(n11503), .A4(n11502), .ZN(
        n11511) );
  AOI22_X1 U14584 ( .A1(n11072), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11509) );
  AOI22_X1 U14585 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U14586 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U14587 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11506) );
  NAND4_X1 U14588 ( .A1(n11509), .A2(n11508), .A3(n11507), .A4(n11506), .ZN(
        n11510) );
  NOR2_X1 U14589 ( .A1(n11511), .A2(n11510), .ZN(n11515) );
  NAND2_X1 U14590 ( .A1(n20806), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11512) );
  NAND2_X1 U14591 ( .A1(n11177), .A2(n11512), .ZN(n11513) );
  AOI21_X1 U14592 ( .B1(n11497), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11513), .ZN(
        n11514) );
  OAI21_X1 U14593 ( .B1(n11688), .B2(n11515), .A(n11514), .ZN(n11520) );
  OAI21_X1 U14594 ( .B1(n11518), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n11564), .ZN(n16061) );
  OR2_X1 U14595 ( .A1(n16061), .A2(n11177), .ZN(n11519) );
  NAND2_X1 U14596 ( .A1(n11520), .A2(n11519), .ZN(n14710) );
  AOI22_X1 U14597 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11072), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14598 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11525) );
  AOI22_X1 U14599 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11144), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U14600 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11523) );
  NAND4_X1 U14601 ( .A1(n11526), .A2(n11525), .A3(n11524), .A4(n11523), .ZN(
        n11533) );
  AOI22_X1 U14602 ( .A1(n11675), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11543), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U14603 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11530) );
  AOI22_X1 U14604 ( .A1(n11527), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11656), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11529) );
  AOI22_X1 U14605 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11528) );
  NAND4_X1 U14606 ( .A1(n11531), .A2(n11530), .A3(n11529), .A4(n11528), .ZN(
        n11532) );
  NOR2_X1 U14607 ( .A1(n11533), .A2(n11532), .ZN(n11536) );
  AOI21_X1 U14608 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14873), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11534) );
  AOI21_X1 U14609 ( .B1(n11497), .B2(P1_EAX_REG_22__SCAN_IN), .A(n11534), .ZN(
        n11535) );
  OAI21_X1 U14610 ( .B1(n11688), .B2(n11536), .A(n11535), .ZN(n11538) );
  XNOR2_X1 U14611 ( .A(n11564), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14877) );
  NAND2_X1 U14612 ( .A1(n14877), .A2(n13980), .ZN(n11537) );
  AOI22_X1 U14613 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11675), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11542) );
  AOI22_X1 U14614 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n9686), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11541) );
  AOI22_X1 U14615 ( .A1(n11527), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11540) );
  AOI22_X1 U14616 ( .A1(n9706), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11539) );
  NAND4_X1 U14617 ( .A1(n11542), .A2(n11541), .A3(n11540), .A4(n11539), .ZN(
        n11549) );
  AOI22_X1 U14618 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11547) );
  AOI22_X1 U14619 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n11543), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11546) );
  AOI22_X1 U14620 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n9711), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U14621 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11099), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11544) );
  NAND4_X1 U14622 ( .A1(n11547), .A2(n11546), .A3(n11545), .A4(n11544), .ZN(
        n11548) );
  NOR2_X1 U14623 ( .A1(n11549), .A2(n11548), .ZN(n11570) );
  AOI22_X1 U14624 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U14625 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11552) );
  AOI22_X1 U14626 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11656), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U14627 ( .A1(n11543), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11099), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11550) );
  NAND4_X1 U14628 ( .A1(n11553), .A2(n11552), .A3(n11551), .A4(n11550), .ZN(
        n11559) );
  AOI22_X1 U14629 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U14630 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11144), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U14631 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U14632 ( .A1(n11060), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11554) );
  NAND4_X1 U14633 ( .A1(n11557), .A2(n11556), .A3(n11555), .A4(n11554), .ZN(
        n11558) );
  NOR2_X1 U14634 ( .A1(n11559), .A2(n11558), .ZN(n11571) );
  XNOR2_X1 U14635 ( .A(n11570), .B(n11571), .ZN(n11563) );
  NAND2_X1 U14636 ( .A1(n20806), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11560) );
  NAND2_X1 U14637 ( .A1(n11177), .A2(n11560), .ZN(n11561) );
  AOI21_X1 U14638 ( .B1(n11497), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11561), .ZN(
        n11562) );
  OAI21_X1 U14639 ( .B1(n11688), .B2(n11563), .A(n11562), .ZN(n11569) );
  INV_X1 U14640 ( .A(n11565), .ZN(n11566) );
  INV_X1 U14641 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14646) );
  NAND2_X1 U14642 ( .A1(n11566), .A2(n14646), .ZN(n11567) );
  NAND2_X1 U14643 ( .A1(n11604), .A2(n11567), .ZN(n14866) );
  OR2_X1 U14644 ( .A1(n14866), .A2(n11177), .ZN(n11568) );
  NOR2_X1 U14645 ( .A1(n11571), .A2(n11570), .ZN(n11599) );
  AOI22_X1 U14646 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11675), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U14647 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11574) );
  AOI22_X1 U14648 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U14649 ( .A1(n11527), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11572) );
  NAND4_X1 U14650 ( .A1(n11575), .A2(n11574), .A3(n11573), .A4(n11572), .ZN(
        n11581) );
  AOI22_X1 U14651 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14652 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14653 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U14654 ( .A1(n11099), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11576) );
  NAND4_X1 U14655 ( .A1(n11579), .A2(n11578), .A3(n11577), .A4(n11576), .ZN(
        n11580) );
  OR2_X1 U14656 ( .A1(n11581), .A2(n11580), .ZN(n11598) );
  INV_X1 U14657 ( .A(n11598), .ZN(n11582) );
  XNOR2_X1 U14658 ( .A(n11599), .B(n11582), .ZN(n11583) );
  NAND2_X1 U14659 ( .A1(n11583), .A2(n11713), .ZN(n11587) );
  INV_X1 U14660 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14858) );
  OAI21_X1 U14661 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14858), .A(n11177), 
        .ZN(n11584) );
  AOI21_X1 U14662 ( .B1(n11173), .B2(P1_EAX_REG_24__SCAN_IN), .A(n11584), .ZN(
        n11586) );
  XNOR2_X1 U14663 ( .A(n11604), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14862) );
  AOI21_X1 U14664 ( .B1(n11587), .B2(n11586), .A(n11585), .ZN(n14629) );
  AOI22_X1 U14665 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11591) );
  AOI22_X1 U14666 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11144), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11590) );
  AOI22_X1 U14667 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U14668 ( .A1(n11675), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11588) );
  NAND4_X1 U14669 ( .A1(n11591), .A2(n11590), .A3(n11589), .A4(n11588), .ZN(
        n11597) );
  AOI22_X1 U14670 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U14671 ( .A1(n11633), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U14672 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11593) );
  AOI22_X1 U14673 ( .A1(n9680), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11592) );
  NAND4_X1 U14674 ( .A1(n11595), .A2(n11594), .A3(n11593), .A4(n11592), .ZN(
        n11596) );
  NOR2_X1 U14675 ( .A1(n11597), .A2(n11596), .ZN(n11612) );
  NAND2_X1 U14676 ( .A1(n11599), .A2(n11598), .ZN(n11611) );
  XNOR2_X1 U14677 ( .A(n11612), .B(n11611), .ZN(n11603) );
  NAND2_X1 U14678 ( .A1(n20806), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11600) );
  NAND2_X1 U14679 ( .A1(n11177), .A2(n11600), .ZN(n11601) );
  AOI21_X1 U14680 ( .B1(n11173), .B2(P1_EAX_REG_25__SCAN_IN), .A(n11601), .ZN(
        n11602) );
  OAI21_X1 U14681 ( .B1(n11603), .B2(n11688), .A(n11602), .ZN(n11610) );
  INV_X1 U14682 ( .A(n11606), .ZN(n11607) );
  INV_X1 U14683 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14617) );
  NAND2_X1 U14684 ( .A1(n11607), .A2(n14617), .ZN(n11608) );
  NAND2_X1 U14685 ( .A1(n11646), .A2(n11608), .ZN(n14851) );
  NAND2_X1 U14686 ( .A1(n11610), .A2(n11609), .ZN(n14614) );
  NOR2_X1 U14687 ( .A1(n11612), .A2(n11611), .ZN(n11641) );
  AOI22_X1 U14688 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11698), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11616) );
  AOI22_X1 U14689 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11072), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U14690 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11614) );
  AOI22_X1 U14691 ( .A1(n11527), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11613) );
  NAND4_X1 U14692 ( .A1(n11616), .A2(n11615), .A3(n11614), .A4(n11613), .ZN(
        n11622) );
  AOI22_X1 U14693 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11143), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11620) );
  AOI22_X1 U14694 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U14695 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14696 ( .A1(n11099), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10938), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11617) );
  NAND4_X1 U14697 ( .A1(n11620), .A2(n11619), .A3(n11618), .A4(n11617), .ZN(
        n11621) );
  OR2_X1 U14698 ( .A1(n11622), .A2(n11621), .ZN(n11640) );
  XNOR2_X1 U14699 ( .A(n11641), .B(n11640), .ZN(n11626) );
  NAND2_X1 U14700 ( .A1(n20806), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11623) );
  NAND2_X1 U14701 ( .A1(n11177), .A2(n11623), .ZN(n11624) );
  AOI21_X1 U14702 ( .B1(n11173), .B2(P1_EAX_REG_26__SCAN_IN), .A(n11624), .ZN(
        n11625) );
  OAI21_X1 U14703 ( .B1(n11626), .B2(n11688), .A(n11625), .ZN(n11628) );
  XNOR2_X1 U14704 ( .A(n11646), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14840) );
  NAND2_X1 U14705 ( .A1(n14840), .A2(n13980), .ZN(n11627) );
  AOI22_X1 U14706 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11632) );
  AOI22_X1 U14707 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11144), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11631) );
  AOI22_X1 U14708 ( .A1(n11527), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9674), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U14709 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11629) );
  NAND4_X1 U14710 ( .A1(n11632), .A2(n11631), .A3(n11630), .A4(n11629), .ZN(
        n11639) );
  AOI22_X1 U14711 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11699), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11637) );
  AOI22_X1 U14712 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U14713 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U14714 ( .A1(n11060), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11145), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11634) );
  NAND4_X1 U14715 ( .A1(n11637), .A2(n11636), .A3(n11635), .A4(n11634), .ZN(
        n11638) );
  NOR2_X1 U14716 ( .A1(n11639), .A2(n11638), .ZN(n11655) );
  NAND2_X1 U14717 ( .A1(n11641), .A2(n11640), .ZN(n11654) );
  XNOR2_X1 U14718 ( .A(n11655), .B(n11654), .ZN(n11645) );
  NAND2_X1 U14719 ( .A1(n20806), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11642) );
  NAND2_X1 U14720 ( .A1(n11177), .A2(n11642), .ZN(n11643) );
  AOI21_X1 U14721 ( .B1(n11497), .B2(P1_EAX_REG_27__SCAN_IN), .A(n11643), .ZN(
        n11644) );
  OAI21_X1 U14722 ( .B1(n11645), .B2(n11688), .A(n11644), .ZN(n11653) );
  INV_X1 U14723 ( .A(n11646), .ZN(n11647) );
  INV_X1 U14724 ( .A(n11648), .ZN(n11650) );
  INV_X1 U14725 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11649) );
  NAND2_X1 U14726 ( .A1(n11650), .A2(n11649), .ZN(n11651) );
  NAND2_X1 U14727 ( .A1(n11690), .A2(n11651), .ZN(n14834) );
  NAND2_X1 U14728 ( .A1(n11653), .A2(n11652), .ZN(n14591) );
  NOR2_X1 U14729 ( .A1(n11655), .A2(n11654), .ZN(n11674) );
  AOI22_X1 U14730 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11698), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14731 ( .A1(n9680), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11060), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14732 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U14733 ( .A1(n11527), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11656), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11657) );
  NAND4_X1 U14734 ( .A1(n11660), .A2(n11659), .A3(n11658), .A4(n11657), .ZN(
        n11666) );
  AOI22_X1 U14735 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U14736 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U14737 ( .A1(n11144), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11662) );
  AOI22_X1 U14738 ( .A1(n11099), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11661) );
  NAND4_X1 U14739 ( .A1(n11664), .A2(n11663), .A3(n11662), .A4(n11661), .ZN(
        n11665) );
  OR2_X1 U14740 ( .A1(n11666), .A2(n11665), .ZN(n11673) );
  INV_X1 U14741 ( .A(n11673), .ZN(n11667) );
  XNOR2_X1 U14742 ( .A(n11674), .B(n11667), .ZN(n11668) );
  NAND2_X1 U14743 ( .A1(n11668), .A2(n11713), .ZN(n11672) );
  INV_X1 U14744 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14815) );
  AOI21_X1 U14745 ( .B1(n14815), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11669) );
  AOI21_X1 U14746 ( .B1(n11173), .B2(P1_EAX_REG_28__SCAN_IN), .A(n11669), .ZN(
        n11671) );
  XNOR2_X1 U14747 ( .A(n11690), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14817) );
  AOI21_X1 U14748 ( .B1(n11672), .B2(n11671), .A(n11670), .ZN(n14573) );
  NAND2_X1 U14749 ( .A1(n11674), .A2(n11673), .ZN(n11695) );
  AOI22_X1 U14750 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11675), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14751 ( .A1(n11098), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11144), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14752 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U14753 ( .A1(n11145), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11676) );
  NAND4_X1 U14754 ( .A1(n11679), .A2(n11678), .A3(n11677), .A4(n11676), .ZN(
        n11685) );
  AOI22_X1 U14755 ( .A1(n9680), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11072), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14756 ( .A1(n11143), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U14757 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U14758 ( .A1(n11697), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11656), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11680) );
  NAND4_X1 U14759 ( .A1(n11683), .A2(n11682), .A3(n11681), .A4(n11680), .ZN(
        n11684) );
  NOR2_X1 U14760 ( .A1(n11685), .A2(n11684), .ZN(n11696) );
  XNOR2_X1 U14761 ( .A(n11695), .B(n11696), .ZN(n11689) );
  INV_X1 U14762 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14811) );
  AOI21_X1 U14763 ( .B1(n14811), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11686) );
  AOI21_X1 U14764 ( .B1(n11173), .B2(P1_EAX_REG_29__SCAN_IN), .A(n11686), .ZN(
        n11687) );
  OAI21_X1 U14765 ( .B1(n11689), .B2(n11688), .A(n11687), .ZN(n11694) );
  NAND2_X1 U14766 ( .A1(n11691), .A2(n14811), .ZN(n11692) );
  NAND2_X1 U14767 ( .A1(n14809), .A2(n13980), .ZN(n11693) );
  NAND2_X1 U14768 ( .A1(n11694), .A2(n11693), .ZN(n14563) );
  NOR2_X1 U14769 ( .A1(n11696), .A2(n11695), .ZN(n11712) );
  AOI22_X1 U14770 ( .A1(n11698), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11697), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11704) );
  AOI22_X1 U14771 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9706), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11703) );
  AOI22_X1 U14772 ( .A1(n11699), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11527), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11702) );
  AOI22_X1 U14773 ( .A1(n11060), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11700), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11701) );
  NAND4_X1 U14774 ( .A1(n11704), .A2(n11703), .A3(n11702), .A4(n11701), .ZN(
        n11710) );
  AOI22_X1 U14775 ( .A1(n9711), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11143), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U14776 ( .A1(n11098), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11522), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11707) );
  AOI22_X1 U14777 ( .A1(n11521), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9675), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11706) );
  AOI22_X1 U14778 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11099), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11705) );
  NAND4_X1 U14779 ( .A1(n11708), .A2(n11707), .A3(n11706), .A4(n11705), .ZN(
        n11709) );
  NOR2_X1 U14780 ( .A1(n11710), .A2(n11709), .ZN(n11711) );
  XNOR2_X1 U14781 ( .A(n11712), .B(n11711), .ZN(n11714) );
  NAND2_X1 U14782 ( .A1(n11714), .A2(n11713), .ZN(n11718) );
  INV_X1 U14783 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12910) );
  AOI21_X1 U14784 ( .B1(n12910), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11715) );
  AOI21_X1 U14785 ( .B1(n11173), .B2(P1_EAX_REG_30__SCAN_IN), .A(n11715), .ZN(
        n11717) );
  XNOR2_X1 U14786 ( .A(n12439), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14555) );
  AND2_X1 U14787 ( .A1(n14555), .A2(n13980), .ZN(n11716) );
  AOI21_X1 U14788 ( .B1(n11718), .B2(n11717), .A(n11716), .ZN(n12432) );
  INV_X1 U14789 ( .A(n12432), .ZN(n11719) );
  XNOR2_X1 U14790 ( .A(n14562), .B(n11719), .ZN(n12912) );
  INV_X1 U14791 ( .A(n13984), .ZN(n13520) );
  NAND2_X1 U14792 ( .A1(n13520), .A2(n9699), .ZN(n11721) );
  NAND2_X1 U14793 ( .A1(n11721), .A2(n11720), .ZN(n11722) );
  INV_X1 U14794 ( .A(n13611), .ZN(n11724) );
  NOR2_X1 U14795 ( .A1(n13608), .A2(n11724), .ZN(n13504) );
  NAND2_X1 U14796 ( .A1(n10119), .A2(n14060), .ZN(n13500) );
  OR2_X1 U14797 ( .A1(n11032), .A2(n13596), .ZN(n13497) );
  NOR2_X1 U14798 ( .A1(n13500), .A2(n13497), .ZN(n11725) );
  MUX2_X1 U14799 ( .A(n11726), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11738) );
  NAND2_X1 U14800 ( .A1(n14105), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11741) );
  NAND2_X1 U14801 ( .A1(n11738), .A2(n11737), .ZN(n11728) );
  NAND2_X1 U14802 ( .A1(n11726), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11727) );
  NAND2_X1 U14803 ( .A1(n11728), .A2(n11727), .ZN(n11753) );
  MUX2_X1 U14804 ( .A(n11729), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11752) );
  NAND2_X1 U14805 ( .A1(n11753), .A2(n11752), .ZN(n11731) );
  NAND2_X1 U14806 ( .A1(n11729), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11730) );
  NOR2_X1 U14807 ( .A1(n14074), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11732) );
  NAND2_X1 U14808 ( .A1(n11733), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11734) );
  NAND2_X1 U14809 ( .A1(n11764), .A2(n11912), .ZN(n11777) );
  NAND2_X1 U14810 ( .A1(n11912), .A2(n11740), .ZN(n11775) );
  XNOR2_X1 U14811 ( .A(n11736), .B(n11735), .ZN(n11909) );
  XNOR2_X1 U14812 ( .A(n11738), .B(n11737), .ZN(n11908) );
  AOI22_X1 U14813 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n11743), .B1(n11740), 
        .B2(n13992), .ZN(n11751) );
  INV_X1 U14814 ( .A(n11751), .ZN(n11739) );
  NOR2_X1 U14815 ( .A1(n11908), .A2(n11739), .ZN(n11749) );
  INV_X1 U14816 ( .A(n11740), .ZN(n11759) );
  OAI21_X1 U14817 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14105), .A(
        n11741), .ZN(n11742) );
  NOR2_X1 U14818 ( .A1(n11759), .A2(n11742), .ZN(n11748) );
  INV_X1 U14819 ( .A(n11742), .ZN(n11745) );
  NAND2_X1 U14820 ( .A1(n11743), .A2(n13802), .ZN(n11744) );
  NAND2_X1 U14821 ( .A1(n11744), .A2(n13596), .ZN(n11758) );
  OAI211_X1 U14822 ( .C1(n9699), .C2(n11746), .A(n11745), .B(n11758), .ZN(
        n11747) );
  OAI21_X1 U14823 ( .B1(n11764), .B2(n11748), .A(n11747), .ZN(n11750) );
  NAND2_X1 U14824 ( .A1(n11749), .A2(n11750), .ZN(n11757) );
  NAND2_X1 U14825 ( .A1(n11751), .A2(n13992), .ZN(n11770) );
  OAI211_X1 U14826 ( .C1(n11751), .C2(n11750), .A(n11908), .B(n11770), .ZN(
        n11756) );
  XNOR2_X1 U14827 ( .A(n11753), .B(n11752), .ZN(n11907) );
  NAND2_X1 U14828 ( .A1(n11768), .A2(n11907), .ZN(n11754) );
  OAI211_X1 U14829 ( .C1(n11759), .C2(n11907), .A(n11754), .B(n11758), .ZN(
        n11755) );
  NAND3_X1 U14830 ( .A1(n11757), .A2(n11756), .A3(n11755), .ZN(n11761) );
  AOI22_X1 U14831 ( .A1(n11762), .A2(n11909), .B1(n11761), .B2(n11760), .ZN(
        n11763) );
  AOI21_X1 U14832 ( .B1(n11764), .B2(n11909), .A(n11763), .ZN(n11772) );
  INV_X1 U14833 ( .A(n11910), .ZN(n11767) );
  NOR2_X1 U14834 ( .A1(n11768), .A2(n11767), .ZN(n11771) );
  NAND2_X1 U14835 ( .A1(n11768), .A2(n11910), .ZN(n11769) );
  OAI22_X1 U14836 ( .A1(n11772), .A2(n11771), .B1(n11770), .B2(n11769), .ZN(
        n11773) );
  AOI21_X1 U14837 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20222), .A(
        n11773), .ZN(n11774) );
  NAND2_X1 U14838 ( .A1(n11775), .A2(n11774), .ZN(n11776) );
  NAND3_X1 U14839 ( .A1(n13622), .A2(n13601), .A3(n13521), .ZN(n11782) );
  NOR2_X1 U14840 ( .A1(n11033), .A2(n20219), .ZN(n11779) );
  NOR2_X1 U14841 ( .A1(n13384), .A2(n9710), .ZN(n11778) );
  NAND4_X1 U14842 ( .A1(n11780), .A2(n11779), .A3(n11778), .A4(n11001), .ZN(
        n11919) );
  INV_X1 U14843 ( .A(n9684), .ZN(n14522) );
  OR2_X1 U14844 ( .A1(n11919), .A2(n14522), .ZN(n11781) );
  AOI22_X1 U14845 ( .A1(n14523), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n14522), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14521) );
  MUX2_X1 U14846 ( .A(n11892), .B(n11808), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n11787) );
  NAND2_X1 U14847 ( .A1(n14522), .A2(n11785), .ZN(n11786) );
  OAI211_X1 U14848 ( .C1(n14523), .C2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n11787), .B(n11786), .ZN(n11793) );
  INV_X1 U14849 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n11788) );
  OR2_X1 U14850 ( .A1(n11797), .A2(n11788), .ZN(n11790) );
  NAND2_X1 U14851 ( .A1(n11785), .A2(n11788), .ZN(n11789) );
  NAND2_X1 U14852 ( .A1(n11790), .A2(n11789), .ZN(n11792) );
  XNOR2_X1 U14853 ( .A(n11793), .B(n11792), .ZN(n13563) );
  INV_X1 U14854 ( .A(n11792), .ZN(n13715) );
  AND2_X1 U14855 ( .A1(n11793), .A2(n13715), .ZN(n11794) );
  MUX2_X1 U14856 ( .A(n11892), .B(n11808), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n11795) );
  OAI21_X1 U14857 ( .B1(n14523), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n11795), .ZN(n13618) );
  INV_X1 U14858 ( .A(n13618), .ZN(n11796) );
  NAND2_X1 U14859 ( .A1(n13616), .A2(n11796), .ZN(n13647) );
  OR2_X1 U14860 ( .A1(n11898), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n11802) );
  INV_X1 U14861 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12355) );
  NAND2_X1 U14862 ( .A1(n11797), .A2(n12355), .ZN(n11800) );
  INV_X1 U14863 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n11798) );
  NAND2_X1 U14864 ( .A1(n9684), .A2(n11798), .ZN(n11799) );
  NAND3_X1 U14865 ( .A1(n11800), .A2(n11808), .A3(n11799), .ZN(n11801) );
  AND2_X1 U14866 ( .A1(n11802), .A2(n11801), .ZN(n13648) );
  INV_X1 U14867 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n20290) );
  NAND2_X1 U14868 ( .A1(n9684), .A2(n20290), .ZN(n11805) );
  NAND2_X1 U14869 ( .A1(n11808), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11804) );
  NAND3_X1 U14870 ( .A1(n11797), .A2(n11805), .A3(n11804), .ZN(n11806) );
  OAI21_X1 U14871 ( .B1(n11892), .B2(P1_EBX_REG_4__SCAN_IN), .A(n11806), .ZN(
        n13792) );
  OR2_X1 U14872 ( .A1(n11898), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n11813) );
  NAND2_X1 U14873 ( .A1(n11808), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11809) );
  NAND2_X1 U14874 ( .A1(n11797), .A2(n11809), .ZN(n11811) );
  INV_X1 U14875 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n14111) );
  NAND2_X1 U14876 ( .A1(n9684), .A2(n14111), .ZN(n11810) );
  NAND2_X1 U14877 ( .A1(n11811), .A2(n11810), .ZN(n11812) );
  NAND2_X1 U14878 ( .A1(n11813), .A2(n11812), .ZN(n14108) );
  INV_X1 U14879 ( .A(n11892), .ZN(n11836) );
  INV_X1 U14880 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20323) );
  NAND2_X1 U14881 ( .A1(n11836), .A2(n20323), .ZN(n11817) );
  NAND2_X1 U14882 ( .A1(n9684), .A2(n20323), .ZN(n11815) );
  NAND2_X1 U14883 ( .A1(n11808), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11814) );
  NAND3_X1 U14884 ( .A1(n11797), .A2(n11815), .A3(n11814), .ZN(n11816) );
  INV_X1 U14885 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n11818) );
  NAND2_X1 U14886 ( .A1(n11836), .A2(n11818), .ZN(n11822) );
  NAND2_X1 U14887 ( .A1(n9684), .A2(n11818), .ZN(n11820) );
  NAND2_X1 U14888 ( .A1(n11808), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11819) );
  NAND3_X1 U14889 ( .A1(n11797), .A2(n11820), .A3(n11819), .ZN(n11821) );
  AND2_X1 U14890 ( .A1(n11822), .A2(n11821), .ZN(n14280) );
  OR2_X1 U14891 ( .A1(n11898), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n11827) );
  NAND2_X1 U14892 ( .A1(n11808), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11823) );
  NAND2_X1 U14893 ( .A1(n11797), .A2(n11823), .ZN(n11825) );
  INV_X1 U14894 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n14155) );
  NAND2_X1 U14895 ( .A1(n9684), .A2(n14155), .ZN(n11824) );
  NAND2_X1 U14896 ( .A1(n11825), .A2(n11824), .ZN(n11826) );
  NAND2_X1 U14897 ( .A1(n11827), .A2(n11826), .ZN(n14281) );
  NAND2_X1 U14898 ( .A1(n14280), .A2(n14281), .ZN(n11828) );
  OR2_X1 U14899 ( .A1(n11898), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n11833) );
  NAND2_X1 U14900 ( .A1(n11808), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11829) );
  NAND2_X1 U14901 ( .A1(n11797), .A2(n11829), .ZN(n11831) );
  INV_X1 U14902 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n14341) );
  NAND2_X1 U14903 ( .A1(n9684), .A2(n14341), .ZN(n11830) );
  NAND2_X1 U14904 ( .A1(n11831), .A2(n11830), .ZN(n11832) );
  MUX2_X1 U14905 ( .A(n11892), .B(n11808), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n11834) );
  OAI21_X1 U14906 ( .B1(n14523), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n11834), .ZN(n11835) );
  INV_X1 U14907 ( .A(n11835), .ZN(n14379) );
  INV_X1 U14908 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n16116) );
  NAND2_X1 U14909 ( .A1(n11836), .A2(n16116), .ZN(n11840) );
  NAND2_X1 U14910 ( .A1(n9684), .A2(n16116), .ZN(n11838) );
  NAND2_X1 U14911 ( .A1(n11808), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11837) );
  NAND3_X1 U14912 ( .A1(n11797), .A2(n11838), .A3(n11837), .ZN(n11839) );
  AND2_X1 U14913 ( .A1(n11840), .A2(n11839), .ZN(n15092) );
  OR2_X1 U14914 ( .A1(n11898), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n11844) );
  INV_X1 U14915 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16161) );
  NAND2_X1 U14916 ( .A1(n11797), .A2(n16161), .ZN(n11842) );
  INV_X1 U14917 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n16118) );
  NAND2_X1 U14918 ( .A1(n9684), .A2(n16118), .ZN(n11841) );
  NAND3_X1 U14919 ( .A1(n11842), .A2(n11808), .A3(n11841), .ZN(n11843) );
  NAND2_X1 U14920 ( .A1(n11844), .A2(n11843), .ZN(n16106) );
  OR2_X1 U14921 ( .A1(n11898), .A2(P1_EBX_REG_13__SCAN_IN), .ZN(n11848) );
  INV_X1 U14922 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16245) );
  NAND2_X1 U14923 ( .A1(n11797), .A2(n16245), .ZN(n11846) );
  INV_X1 U14924 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n16086) );
  NAND2_X1 U14925 ( .A1(n9684), .A2(n16086), .ZN(n11845) );
  NAND3_X1 U14926 ( .A1(n11846), .A2(n11808), .A3(n11845), .ZN(n11847) );
  MUX2_X1 U14927 ( .A(n11892), .B(n11808), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n11849) );
  OAI21_X1 U14928 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n14523), .A(
        n11849), .ZN(n14441) );
  OR2_X1 U14929 ( .A1(n11898), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n11853) );
  INV_X1 U14930 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15084) );
  NAND2_X1 U14931 ( .A1(n11797), .A2(n15084), .ZN(n11851) );
  INV_X1 U14932 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14469) );
  NAND2_X1 U14933 ( .A1(n9684), .A2(n14469), .ZN(n11850) );
  NAND3_X1 U14934 ( .A1(n11851), .A2(n11808), .A3(n11850), .ZN(n11852) );
  NAND2_X1 U14935 ( .A1(n11853), .A2(n11852), .ZN(n14464) );
  MUX2_X1 U14936 ( .A(n11892), .B(n11808), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n11854) );
  OAI21_X1 U14937 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n14523), .A(
        n11854), .ZN(n14693) );
  OR2_X1 U14938 ( .A1(n11898), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n11858) );
  INV_X1 U14939 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16137) );
  NAND2_X1 U14940 ( .A1(n11797), .A2(n16137), .ZN(n11856) );
  INV_X1 U14941 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n16074) );
  NAND2_X1 U14942 ( .A1(n9684), .A2(n16074), .ZN(n11855) );
  NAND3_X1 U14943 ( .A1(n11856), .A2(n11808), .A3(n11855), .ZN(n11857) );
  MUX2_X1 U14944 ( .A(n11892), .B(n11808), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n11859) );
  OAI21_X1 U14945 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n14523), .A(
        n11859), .ZN(n14679) );
  OR2_X1 U14946 ( .A1(n11898), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n11863) );
  INV_X1 U14947 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14954) );
  NAND2_X1 U14948 ( .A1(n11797), .A2(n14954), .ZN(n11861) );
  INV_X1 U14949 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n16071) );
  NAND2_X1 U14950 ( .A1(n9684), .A2(n16071), .ZN(n11860) );
  NAND3_X1 U14951 ( .A1(n11861), .A2(n11808), .A3(n11860), .ZN(n11862) );
  NAND2_X1 U14952 ( .A1(n11863), .A2(n11862), .ZN(n14724) );
  NAND2_X1 U14953 ( .A1(n14725), .A2(n14724), .ZN(n14727) );
  INV_X1 U14954 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14719) );
  NAND2_X1 U14955 ( .A1(n9684), .A2(n14719), .ZN(n11865) );
  NAND2_X1 U14956 ( .A1(n11808), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11864) );
  NAND3_X1 U14957 ( .A1(n11797), .A2(n11865), .A3(n11864), .ZN(n11866) );
  OAI21_X1 U14958 ( .B1(n11892), .B2(P1_EBX_REG_20__SCAN_IN), .A(n11866), .ZN(
        n14667) );
  OR2_X1 U14959 ( .A1(n11898), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n11870) );
  INV_X1 U14960 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15045) );
  NAND2_X1 U14961 ( .A1(n11797), .A2(n15045), .ZN(n11868) );
  INV_X1 U14962 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14716) );
  NAND2_X1 U14963 ( .A1(n9684), .A2(n14716), .ZN(n11867) );
  NAND3_X1 U14964 ( .A1(n11868), .A2(n11808), .A3(n11867), .ZN(n11869) );
  MUX2_X1 U14965 ( .A(n11892), .B(n11808), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n11872) );
  OR2_X1 U14966 ( .A1(n14523), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11871) );
  AND2_X1 U14967 ( .A1(n11872), .A2(n11871), .ZN(n14656) );
  OR2_X1 U14968 ( .A1(n11898), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n11876) );
  INV_X1 U14969 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16197) );
  NAND2_X1 U14970 ( .A1(n11797), .A2(n16197), .ZN(n11874) );
  INV_X1 U14971 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14708) );
  NAND2_X1 U14972 ( .A1(n9684), .A2(n14708), .ZN(n11873) );
  NAND3_X1 U14973 ( .A1(n11874), .A2(n11808), .A3(n11873), .ZN(n11875) );
  AND2_X1 U14974 ( .A1(n11876), .A2(n11875), .ZN(n14633) );
  MUX2_X1 U14975 ( .A(n11892), .B(n11808), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n11878) );
  OR2_X1 U14976 ( .A1(n14523), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11877) );
  NAND2_X1 U14977 ( .A1(n11878), .A2(n11877), .ZN(n14634) );
  NOR2_X1 U14978 ( .A1(n14633), .A2(n14634), .ZN(n11879) );
  OR2_X1 U14979 ( .A1(n11898), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n11884) );
  NAND2_X1 U14980 ( .A1(n11808), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11880) );
  NAND2_X1 U14981 ( .A1(n11797), .A2(n11880), .ZN(n11882) );
  INV_X1 U14982 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14706) );
  NAND2_X1 U14983 ( .A1(n9684), .A2(n14706), .ZN(n11881) );
  NAND2_X1 U14984 ( .A1(n11882), .A2(n11881), .ZN(n11883) );
  AND2_X1 U14985 ( .A1(n11884), .A2(n11883), .ZN(n14615) );
  INV_X1 U14986 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14704) );
  NAND2_X1 U14987 ( .A1(n9684), .A2(n14704), .ZN(n11886) );
  NAND2_X1 U14988 ( .A1(n11808), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11885) );
  NAND3_X1 U14989 ( .A1(n11797), .A2(n11886), .A3(n11885), .ZN(n11887) );
  OAI21_X1 U14990 ( .B1(n11892), .B2(P1_EBX_REG_26__SCAN_IN), .A(n11887), .ZN(
        n14603) );
  OR2_X1 U14991 ( .A1(n11898), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n11891) );
  INV_X1 U14992 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15002) );
  NAND2_X1 U14993 ( .A1(n11797), .A2(n15002), .ZN(n11889) );
  INV_X1 U14994 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14703) );
  NAND2_X1 U14995 ( .A1(n9684), .A2(n14703), .ZN(n11888) );
  NAND3_X1 U14996 ( .A1(n11889), .A2(n11808), .A3(n11888), .ZN(n11890) );
  MUX2_X1 U14997 ( .A(n11892), .B(n11808), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n11894) );
  OR2_X1 U14998 ( .A1(n14523), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11893) );
  AND2_X1 U14999 ( .A1(n11894), .A2(n11893), .ZN(n14574) );
  OR2_X1 U15000 ( .A1(n14523), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11897) );
  INV_X1 U15001 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n11895) );
  NAND2_X1 U15002 ( .A1(n9684), .A2(n11895), .ZN(n11896) );
  NAND2_X1 U15003 ( .A1(n11897), .A2(n11896), .ZN(n11900) );
  OAI22_X1 U15004 ( .A1(n11900), .A2(n11785), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n11898), .ZN(n14564) );
  NAND2_X1 U15005 ( .A1(n14520), .A2(n11785), .ZN(n11901) );
  INV_X1 U15006 ( .A(n14576), .ZN(n11899) );
  AOI22_X1 U15007 ( .A1(n11901), .A2(n11900), .B1(n11899), .B2(n11808), .ZN(
        n11902) );
  XOR2_X1 U15008 ( .A(n14521), .B(n11902), .Z(n14551) );
  INV_X1 U15009 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14558) );
  OAI21_X1 U15010 ( .B1(n14551), .B2(n14737), .A(n10180), .ZN(n11903) );
  INV_X1 U15011 ( .A(n11903), .ZN(n11904) );
  NAND2_X1 U15012 ( .A1(n11905), .A2(n11904), .ZN(P1_U2842) );
  NOR4_X1 U15013 ( .A1(n11910), .A2(n11909), .A3(n11908), .A4(n11907), .ZN(
        n11911) );
  OR2_X1 U15014 ( .A1(n11912), .A2(n11911), .ZN(n13593) );
  INV_X1 U15015 ( .A(n13593), .ZN(n11913) );
  NAND2_X1 U15016 ( .A1(n11906), .A2(n11913), .ZN(n13374) );
  NAND2_X1 U15017 ( .A1(n13596), .A2(n20906), .ZN(n11918) );
  INV_X1 U15018 ( .A(n20906), .ZN(n16022) );
  NAND2_X1 U15019 ( .A1(n9692), .A2(n13989), .ZN(n11914) );
  AND3_X1 U15020 ( .A1(n10119), .A2(n12342), .A3(n11914), .ZN(n13523) );
  NAND2_X1 U15021 ( .A1(n13523), .A2(n13371), .ZN(n13509) );
  OAI21_X1 U15022 ( .B1(n11915), .B2(n16022), .A(n13509), .ZN(n11916) );
  NAND2_X1 U15023 ( .A1(n11916), .A2(n13597), .ZN(n11917) );
  NAND2_X1 U15024 ( .A1(n11032), .A2(n13384), .ZN(n13702) );
  NOR3_X4 U15025 ( .A1(n14783), .A2(n14537), .A3(n9710), .ZN(n14802) );
  NOR4_X1 U15026 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n11925) );
  NOR4_X1 U15027 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n11924) );
  NOR4_X1 U15028 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n11923) );
  NOR4_X1 U15029 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n11922) );
  AND4_X1 U15030 ( .A1(n11925), .A2(n11924), .A3(n11923), .A4(n11922), .ZN(
        n11930) );
  NOR4_X1 U15031 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n11928) );
  NOR4_X1 U15032 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n11927) );
  NOR4_X1 U15033 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n11926) );
  INV_X1 U15034 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20825) );
  AND4_X1 U15035 ( .A1(n11928), .A2(n11927), .A3(n11926), .A4(n20825), .ZN(
        n11929) );
  NAND2_X1 U15036 ( .A1(n11930), .A2(n11929), .ZN(n11931) );
  MUX2_X1 U15037 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n13800), .Z(
        n14449) );
  INV_X1 U15038 ( .A(n11934), .ZN(n13588) );
  NOR3_X1 U15039 ( .A1(n14783), .A2(n13800), .A3(n13588), .ZN(n11932) );
  AOI22_X1 U15040 ( .A1(n14802), .A2(n14449), .B1(n14800), .B2(DATAI_30_), 
        .ZN(n11933) );
  INV_X1 U15041 ( .A(n11933), .ZN(n11938) );
  AND2_X1 U15042 ( .A1(n11934), .A2(n13800), .ZN(n11935) );
  NAND2_X1 U15043 ( .A1(n14743), .A2(n11935), .ZN(n14767) );
  AOI22_X1 U15044 ( .A1(n14799), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14783), .ZN(n11936) );
  NOR2_X1 U15045 ( .A1(n11938), .A2(n11937), .ZN(n11939) );
  OAI21_X1 U15046 ( .B1(n14561), .B2(n14793), .A(n11939), .ZN(P1_U2874) );
  NAND2_X1 U15047 ( .A1(n11960), .A2(n11941), .ZN(n11945) );
  AND2_X1 U15048 ( .A1(n11940), .A2(n11945), .ZN(n11951) );
  INV_X1 U15049 ( .A(n11943), .ZN(n11946) );
  NAND2_X1 U15050 ( .A1(n11943), .A2(n11942), .ZN(n11944) );
  OR2_X2 U15051 ( .A1(n11962), .A2(n11944), .ZN(n11949) );
  AND2_X1 U15052 ( .A1(n11946), .A2(n11945), .ZN(n11947) );
  NAND2_X1 U15053 ( .A1(n11962), .A2(n11947), .ZN(n11948) );
  OAI211_X2 U15054 ( .C1(n11951), .C2(n11950), .A(n11949), .B(n11948), .ZN(
        n12548) );
  BUF_X4 U15055 ( .A(n12548), .Z(n13472) );
  INV_X1 U15056 ( .A(n11955), .ZN(n11956) );
  INV_X1 U15057 ( .A(n11957), .ZN(n11963) );
  INV_X1 U15058 ( .A(n11952), .ZN(n11958) );
  INV_X1 U15059 ( .A(n19559), .ZN(n13416) );
  XNOR2_X1 U15060 ( .A(n11960), .B(n11959), .ZN(n11961) );
  OR2_X2 U15061 ( .A1(n11968), .A2(n9722), .ZN(n19792) );
  INV_X1 U15062 ( .A(n19513), .ZN(n13423) );
  NAND2_X1 U15063 ( .A1(n13962), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11966) );
  NAND2_X1 U15064 ( .A1(n9714), .A2(n11990), .ZN(n11976) );
  NAND2_X1 U15065 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11965) );
  OAI211_X1 U15066 ( .C1(n19792), .C2(n11967), .A(n11966), .B(n11965), .ZN(
        n11975) );
  INV_X1 U15067 ( .A(n11968), .ZN(n11969) );
  INV_X2 U15068 ( .A(n9722), .ZN(n19541) );
  NAND2_X2 U15069 ( .A1(n11969), .A2(n9721), .ZN(n19910) );
  INV_X1 U15070 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11973) );
  NAND3_X2 U15071 ( .A1(n13472), .A2(n11978), .A3(n9713), .ZN(n12021) );
  INV_X1 U15072 ( .A(n12021), .ZN(n19648) );
  INV_X1 U15073 ( .A(n12079), .ZN(n19594) );
  INV_X1 U15074 ( .A(n13472), .ZN(n15817) );
  INV_X1 U15075 ( .A(n13744), .ZN(n11970) );
  NAND2_X1 U15076 ( .A1(n11970), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11971) );
  OAI211_X1 U15077 ( .C1(n19910), .C2(n11973), .A(n11972), .B(n11971), .ZN(
        n11974) );
  NOR2_X1 U15078 ( .A1(n11975), .A2(n11974), .ZN(n11996) );
  INV_X1 U15079 ( .A(n19857), .ZN(n19851) );
  NAND2_X1 U15080 ( .A1(n19851), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11986) );
  INV_X1 U15081 ( .A(n11976), .ZN(n11977) );
  NAND2_X1 U15082 ( .A1(n11977), .A2(n13472), .ZN(n12071) );
  INV_X1 U15083 ( .A(n12071), .ZN(n19701) );
  NAND2_X1 U15084 ( .A1(n11980), .A2(n13472), .ZN(n19757) );
  INV_X1 U15085 ( .A(n19757), .ZN(n11979) );
  AOI22_X1 U15086 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19701), .B1(
        n11979), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11985) );
  INV_X1 U15087 ( .A(n11980), .ZN(n11981) );
  OR2_X2 U15088 ( .A1(n13472), .A2(n11981), .ZN(n12009) );
  INV_X1 U15089 ( .A(n12009), .ZN(n11982) );
  NAND2_X1 U15090 ( .A1(n11982), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11984) );
  NAND2_X1 U15091 ( .A1(n14186), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11983) );
  NAND2_X2 U15092 ( .A1(n11988), .A2(n19541), .ZN(n14176) );
  INV_X1 U15093 ( .A(n14176), .ZN(n14171) );
  NAND2_X2 U15094 ( .A1(n11988), .A2(n9722), .ZN(n19730) );
  INV_X1 U15095 ( .A(n19730), .ZN(n19725) );
  AOI22_X1 U15096 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n14171), .B1(
        n19725), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11994) );
  NAND3_X1 U15097 ( .A1(n15817), .A2(n11990), .A3(n19541), .ZN(n19822) );
  OAI21_X1 U15098 ( .B1(n19822), .B2(n11991), .A(n10648), .ZN(n11992) );
  AOI21_X1 U15099 ( .B1(n14164), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n11992), .ZN(n11993) );
  NAND4_X1 U15100 ( .A1(n11996), .A2(n11995), .A3(n11994), .A4(n11993), .ZN(
        n11998) );
  NAND2_X1 U15101 ( .A1(n16586), .A2(n12030), .ZN(n12281) );
  OR2_X1 U15102 ( .A1(n12282), .A2(n12281), .ZN(n12287) );
  NAND2_X1 U15103 ( .A1(n12287), .A2(n12289), .ZN(n11997) );
  INV_X1 U15104 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12000) );
  INV_X1 U15105 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11999) );
  OAI22_X1 U15106 ( .A1(n12000), .A2(n19857), .B1(n19730), .B2(n11999), .ZN(
        n12004) );
  INV_X1 U15107 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12002) );
  INV_X1 U15108 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12001) );
  OAI22_X1 U15109 ( .A1(n12002), .A2(n12060), .B1(n14176), .B2(n12001), .ZN(
        n12003) );
  INV_X1 U15110 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12005) );
  OAI22_X1 U15111 ( .A1(n12005), .A2(n19792), .B1(n12064), .B2(n19573), .ZN(
        n12015) );
  INV_X1 U15112 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12007) );
  INV_X1 U15113 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12006) );
  INV_X1 U15114 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12010) );
  INV_X1 U15115 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12008) );
  INV_X1 U15116 ( .A(n12011), .ZN(n12012) );
  NAND2_X1 U15117 ( .A1(n12013), .A2(n12012), .ZN(n12014) );
  NOR2_X1 U15118 ( .A1(n12015), .A2(n12014), .ZN(n12028) );
  INV_X1 U15119 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12017) );
  INV_X1 U15120 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12016) );
  OAI22_X1 U15121 ( .A1(n12017), .A2(n19910), .B1(n12039), .B2(n12016), .ZN(
        n12018) );
  INV_X1 U15122 ( .A(n12018), .ZN(n12027) );
  INV_X1 U15123 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12020) );
  INV_X1 U15124 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12019) );
  OAI22_X1 U15125 ( .A1(n19822), .A2(n12020), .B1(n12079), .B2(n12019), .ZN(
        n12025) );
  INV_X1 U15126 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12023) );
  INV_X1 U15127 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12022) );
  OAI22_X1 U15128 ( .A1(n13744), .A2(n12023), .B1(n12021), .B2(n12022), .ZN(
        n12024) );
  NOR2_X1 U15129 ( .A1(n12025), .A2(n12024), .ZN(n12026) );
  NAND3_X1 U15130 ( .A1(n12028), .A2(n12027), .A3(n12026), .ZN(n12029) );
  OAI21_X1 U15131 ( .B1(n10176), .B2(n12029), .A(n10648), .ZN(n12033) );
  NAND2_X1 U15132 ( .A1(n12031), .A2(n12030), .ZN(n12032) );
  INV_X1 U15133 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12652) );
  INV_X1 U15134 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12641) );
  OAI22_X1 U15135 ( .A1(n12652), .A2(n19857), .B1(n19730), .B2(n12641), .ZN(
        n12038) );
  INV_X1 U15136 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14170) );
  INV_X1 U15137 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12036) );
  OAI22_X1 U15138 ( .A1(n14170), .A2(n12060), .B1(n14176), .B2(n12036), .ZN(
        n12037) );
  NOR2_X1 U15139 ( .A1(n12038), .A2(n12037), .ZN(n12053) );
  INV_X1 U15140 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12041) );
  INV_X1 U15141 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12040) );
  OAI22_X1 U15142 ( .A1(n12041), .A2(n19910), .B1(n12039), .B2(n12040), .ZN(
        n12043) );
  INV_X1 U15143 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12632) );
  INV_X1 U15144 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14197) );
  OAI22_X1 U15145 ( .A1(n12632), .A2(n19792), .B1(n12064), .B2(n14197), .ZN(
        n12042) );
  NOR2_X1 U15146 ( .A1(n12043), .A2(n12042), .ZN(n12052) );
  INV_X1 U15147 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12644) );
  INV_X1 U15148 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12636) );
  OAI22_X1 U15149 ( .A1(n12644), .A2(n19757), .B1(n12074), .B2(n12636), .ZN(
        n12045) );
  INV_X1 U15150 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12638) );
  INV_X1 U15151 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12634) );
  OAI22_X1 U15152 ( .A1(n12638), .A2(n12071), .B1(n12009), .B2(n12634), .ZN(
        n12044) );
  NOR2_X1 U15153 ( .A1(n12045), .A2(n12044), .ZN(n12051) );
  INV_X1 U15154 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12650) );
  OAI22_X1 U15155 ( .A1(n19822), .A2(n12650), .B1(n12079), .B2(n9995), .ZN(
        n12049) );
  INV_X1 U15156 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12047) );
  INV_X1 U15157 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12046) );
  OAI22_X1 U15158 ( .A1(n13744), .A2(n12047), .B1(n12021), .B2(n12046), .ZN(
        n12048) );
  NOR2_X1 U15159 ( .A1(n12049), .A2(n12048), .ZN(n12050) );
  NAND4_X1 U15160 ( .A1(n12053), .A2(n12052), .A3(n12051), .A4(n12050), .ZN(
        n12056) );
  NAND2_X1 U15161 ( .A1(n12054), .A2(n12030), .ZN(n12055) );
  INV_X1 U15162 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12058) );
  INV_X1 U15163 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12057) );
  OAI22_X1 U15164 ( .A1(n12058), .A2(n19857), .B1(n14176), .B2(n12057), .ZN(
        n12063) );
  OAI22_X1 U15165 ( .A1(n12061), .A2(n12060), .B1(n19730), .B2(n12059), .ZN(
        n12062) );
  NOR2_X1 U15166 ( .A1(n12063), .A2(n12062), .ZN(n12088) );
  OAI22_X1 U15167 ( .A1(n12065), .A2(n19792), .B1(n12064), .B2(n19582), .ZN(
        n12069) );
  OAI22_X1 U15168 ( .A1(n12067), .A2(n19910), .B1(n12039), .B2(n12066), .ZN(
        n12068) );
  NOR2_X1 U15169 ( .A1(n12069), .A2(n12068), .ZN(n12087) );
  OAI22_X1 U15170 ( .A1(n12072), .A2(n12071), .B1(n12009), .B2(n12070), .ZN(
        n12077) );
  OAI22_X1 U15171 ( .A1(n12075), .A2(n19757), .B1(n12074), .B2(n12073), .ZN(
        n12076) );
  NOR2_X1 U15172 ( .A1(n12077), .A2(n12076), .ZN(n12086) );
  INV_X1 U15173 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12078) );
  OAI22_X1 U15174 ( .A1(n19822), .A2(n12080), .B1(n12079), .B2(n12078), .ZN(
        n12084) );
  INV_X1 U15175 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12082) );
  INV_X1 U15176 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12081) );
  OAI22_X1 U15177 ( .A1(n13744), .A2(n12082), .B1(n12021), .B2(n12081), .ZN(
        n12083) );
  NOR2_X1 U15178 ( .A1(n12084), .A2(n12083), .ZN(n12085) );
  NAND4_X1 U15179 ( .A1(n12088), .A2(n12087), .A3(n12086), .A4(n12085), .ZN(
        n12091) );
  NAND2_X1 U15180 ( .A1(n12089), .A2(n12030), .ZN(n12090) );
  NAND2_X1 U15181 ( .A1(n12092), .A2(n12302), .ZN(n12093) );
  AND2_X1 U15182 ( .A1(n12130), .A2(n12094), .ZN(n12095) );
  OR2_X1 U15183 ( .A1(n12095), .A2(n12097), .ZN(n14120) );
  NAND2_X1 U15184 ( .A1(n14345), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15536) );
  XNOR2_X1 U15185 ( .A(n12097), .B(n12096), .ZN(n19349) );
  NAND2_X1 U15186 ( .A1(n19349), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15757) );
  NAND2_X1 U15187 ( .A1(n12099), .A2(n12098), .ZN(n12100) );
  NAND2_X1 U15188 ( .A1(n12152), .A2(n12100), .ZN(n19336) );
  NOR2_X1 U15189 ( .A1(n19336), .A2(n12101), .ZN(n12148) );
  NAND2_X1 U15190 ( .A1(n12148), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15540) );
  INV_X1 U15191 ( .A(n12125), .ZN(n12104) );
  NAND2_X1 U15192 ( .A1(n12107), .A2(n12102), .ZN(n12103) );
  NAND2_X1 U15193 ( .A1(n12104), .A2(n12103), .ZN(n15209) );
  NAND2_X1 U15194 ( .A1(n12122), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14021) );
  INV_X1 U15195 ( .A(n12105), .ZN(n12111) );
  NAND2_X1 U15196 ( .A1(n12111), .A2(n12106), .ZN(n12108) );
  NAND2_X1 U15197 ( .A1(n12108), .A2(n12107), .ZN(n15216) );
  XNOR2_X1 U15198 ( .A(n15216), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13362) );
  AND2_X1 U15199 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n12109) );
  NAND2_X1 U15200 ( .A1(n9720), .A2(n12109), .ZN(n12110) );
  NAND2_X1 U15201 ( .A1(n12111), .A2(n12110), .ZN(n15234) );
  INV_X1 U15202 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15780) );
  OAI21_X1 U15203 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20182), .A(
        n12112), .ZN(n12448) );
  INV_X1 U15204 ( .A(n12448), .ZN(n12265) );
  NOR2_X1 U15205 ( .A1(n10855), .A2(n10858), .ZN(n12113) );
  AOI21_X1 U15206 ( .B1(n12114), .B2(n12265), .A(n12113), .ZN(n12117) );
  NAND2_X1 U15207 ( .A1(n12115), .A2(n16586), .ZN(n12116) );
  NAND2_X1 U15208 ( .A1(n12117), .A2(n12116), .ZN(n19384) );
  NAND2_X1 U15209 ( .A1(n19384), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16584) );
  OAI21_X1 U15210 ( .B1(n15234), .B2(n15780), .A(n16584), .ZN(n12119) );
  NAND2_X1 U15211 ( .A1(n15234), .A2(n15780), .ZN(n12118) );
  AND2_X1 U15212 ( .A1(n12119), .A2(n12118), .ZN(n13361) );
  NAND2_X1 U15213 ( .A1(n13362), .A2(n13361), .ZN(n13360) );
  INV_X1 U15214 ( .A(n15216), .ZN(n12120) );
  NAND2_X1 U15215 ( .A1(n12120), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12121) );
  AND2_X1 U15216 ( .A1(n13360), .A2(n12121), .ZN(n14023) );
  NAND2_X1 U15217 ( .A1(n14021), .A2(n14023), .ZN(n12123) );
  OR2_X2 U15218 ( .A1(n12122), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14022) );
  OR2_X1 U15219 ( .A1(n12125), .A2(n12124), .ZN(n12126) );
  NAND2_X1 U15220 ( .A1(n12126), .A2(n12128), .ZN(n19363) );
  INV_X1 U15221 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19520) );
  XNOR2_X1 U15222 ( .A(n19363), .B(n19520), .ZN(n19490) );
  NAND2_X1 U15223 ( .A1(n12128), .A2(n12127), .ZN(n12129) );
  NAND2_X1 U15224 ( .A1(n12130), .A2(n12129), .ZN(n15200) );
  AND2_X1 U15225 ( .A1(n15200), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12133) );
  INV_X1 U15226 ( .A(n12133), .ZN(n12131) );
  INV_X1 U15227 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16582) );
  NAND2_X1 U15228 ( .A1(n12101), .A2(n16582), .ZN(n12135) );
  MUX2_X1 U15229 ( .A(n12131), .B(n12135), .S(n12141), .Z(n12139) );
  OAI21_X1 U15230 ( .B1(n12101), .B2(n16582), .A(n15200), .ZN(n12132) );
  OAI21_X1 U15231 ( .B1(n15200), .B2(n16582), .A(n12132), .ZN(n12138) );
  NAND2_X1 U15232 ( .A1(n12141), .A2(n12133), .ZN(n12134) );
  OAI21_X1 U15233 ( .B1(n12141), .B2(n12135), .A(n12134), .ZN(n12136) );
  NAND2_X1 U15234 ( .A1(n12140), .A2(n12136), .ZN(n12137) );
  OAI211_X1 U15235 ( .C1(n12140), .C2(n12139), .A(n12138), .B(n12137), .ZN(
        n16495) );
  NAND2_X1 U15236 ( .A1(n12298), .A2(n12101), .ZN(n12143) );
  NAND2_X1 U15237 ( .A1(n12143), .A2(n15200), .ZN(n12144) );
  NAND2_X1 U15238 ( .A1(n12144), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12145) );
  INV_X1 U15239 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12512) );
  NAND3_X1 U15240 ( .A1(n15540), .A2(n12512), .A3(n15757), .ZN(n12150) );
  INV_X1 U15241 ( .A(n19349), .ZN(n12147) );
  NAND2_X1 U15242 ( .A1(n12147), .A2(n15763), .ZN(n15756) );
  INV_X1 U15243 ( .A(n12148), .ZN(n12149) );
  NAND2_X1 U15244 ( .A1(n12149), .A2(n12310), .ZN(n15539) );
  NAND2_X1 U15245 ( .A1(n12152), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12151) );
  MUX2_X1 U15246 ( .A(n12152), .B(n12151), .S(n9720), .Z(n12153) );
  INV_X1 U15247 ( .A(n12153), .ZN(n12154) );
  NOR2_X1 U15248 ( .A1(n12154), .A2(n12155), .ZN(n15181) );
  AOI21_X1 U15249 ( .B1(n15181), .B2(n12162), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15744) );
  NAND2_X1 U15250 ( .A1(n9720), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12156) );
  MUX2_X1 U15251 ( .A(n12156), .B(P2_EBX_REG_10__SCAN_IN), .S(n12155), .Z(
        n12157) );
  NAND2_X1 U15252 ( .A1(n12157), .A2(n12235), .ZN(n19322) );
  INV_X1 U15253 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15731) );
  NAND2_X1 U15254 ( .A1(n12172), .A2(n15731), .ZN(n15727) );
  NAND2_X1 U15255 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n12158), .ZN(n12159) );
  NOR2_X1 U15256 ( .A1(n10855), .A2(n12159), .ZN(n12160) );
  NOR2_X1 U15257 ( .A1(n12161), .A2(n12160), .ZN(n12169) );
  AOI21_X1 U15258 ( .B1(n12169), .B2(n12162), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16464) );
  NOR2_X1 U15259 ( .A1(n12167), .A2(n12166), .ZN(n12168) );
  NOR2_X1 U15260 ( .A1(n12165), .A2(n12168), .ZN(n19310) );
  AND2_X1 U15261 ( .A1(n19310), .A2(n12162), .ZN(n12188) );
  NAND2_X1 U15262 ( .A1(n12188), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15717) );
  INV_X1 U15263 ( .A(n12169), .ZN(n13241) );
  INV_X1 U15264 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16546) );
  OR2_X1 U15265 ( .A1(n12101), .A2(n16546), .ZN(n12170) );
  OR2_X1 U15266 ( .A1(n13241), .A2(n12170), .ZN(n16465) );
  INV_X1 U15267 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15749) );
  NOR2_X1 U15268 ( .A1(n12101), .A2(n15749), .ZN(n12171) );
  NAND2_X1 U15269 ( .A1(n15181), .A2(n12171), .ZN(n15725) );
  OR2_X1 U15270 ( .A1(n15731), .A2(n12172), .ZN(n15726) );
  AND2_X1 U15271 ( .A1(n16465), .A2(n10186), .ZN(n15714) );
  INV_X1 U15272 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15696) );
  INV_X1 U15273 ( .A(n12175), .ZN(n12173) );
  NAND2_X1 U15274 ( .A1(n12173), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12174) );
  MUX2_X1 U15275 ( .A(n12174), .B(n12173), .S(n10855), .Z(n12176) );
  INV_X1 U15276 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n14150) );
  NAND2_X1 U15277 ( .A1(n12175), .A2(n14150), .ZN(n12201) );
  NAND2_X1 U15278 ( .A1(n12176), .A2(n12201), .ZN(n19289) );
  NAND2_X1 U15279 ( .A1(n15696), .A2(n12206), .ZN(n15702) );
  NOR2_X1 U15280 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n12215), .ZN(
        n15490) );
  NAND2_X1 U15281 ( .A1(n12185), .A2(n12178), .ZN(n12179) );
  NAND2_X1 U15282 ( .A1(n12180), .A2(n12179), .ZN(n19242) );
  NOR2_X1 U15283 ( .A1(n19242), .A2(n12101), .ZN(n12209) );
  NOR2_X1 U15284 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n12209), .ZN(
        n15501) );
  NOR2_X2 U15285 ( .A1(n15490), .A2(n15501), .ZN(n15464) );
  NAND2_X1 U15286 ( .A1(n9720), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12182) );
  NAND2_X1 U15287 ( .A1(n12200), .A2(n12181), .ZN(n12184) );
  OAI211_X1 U15288 ( .C1(n12200), .C2(n12182), .A(n12235), .B(n12184), .ZN(
        n19265) );
  OR2_X1 U15289 ( .A1(n19265), .A2(n12101), .ZN(n12210) );
  INV_X1 U15290 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15671) );
  XNOR2_X1 U15291 ( .A(n12210), .B(n15671), .ZN(n15529) );
  INV_X1 U15292 ( .A(n15529), .ZN(n12191) );
  NOR2_X1 U15293 ( .A1(n10855), .A2(n10875), .ZN(n12183) );
  NAND2_X1 U15294 ( .A1(n12184), .A2(n12183), .ZN(n12186) );
  NAND2_X1 U15295 ( .A1(n12186), .A2(n12185), .ZN(n19252) );
  OR2_X1 U15296 ( .A1(n19252), .A2(n12101), .ZN(n12187) );
  INV_X1 U15297 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15679) );
  NAND2_X1 U15298 ( .A1(n12187), .A2(n15679), .ZN(n15463) );
  NOR2_X1 U15299 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n12188), .ZN(
        n16450) );
  INV_X1 U15300 ( .A(n16450), .ZN(n15716) );
  INV_X1 U15301 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16536) );
  INV_X1 U15302 ( .A(n12189), .ZN(n12190) );
  XNOR2_X1 U15303 ( .A(n12165), .B(n12190), .ZN(n19302) );
  NAND2_X1 U15304 ( .A1(n19302), .A2(n12162), .ZN(n12213) );
  NAND2_X1 U15305 ( .A1(n16536), .A2(n12213), .ZN(n16448) );
  AND2_X1 U15306 ( .A1(n15716), .A2(n16448), .ZN(n15700) );
  AND3_X1 U15307 ( .A1(n12192), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n9720), .ZN(
        n12193) );
  NOR2_X1 U15308 ( .A1(n12194), .A2(n12193), .ZN(n15167) );
  NAND2_X1 U15309 ( .A1(n15167), .A2(n12162), .ZN(n12195) );
  NAND2_X1 U15310 ( .A1(n12195), .A2(n15470), .ZN(n15465) );
  NOR2_X1 U15311 ( .A1(n10855), .A2(n16401), .ZN(n12196) );
  XNOR2_X1 U15312 ( .A(n12197), .B(n12196), .ZN(n19221) );
  NAND2_X1 U15313 ( .A1(n19221), .A2(n12162), .ZN(n12214) );
  INV_X1 U15314 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15636) );
  AND2_X1 U15315 ( .A1(n12214), .A2(n15636), .ZN(n15479) );
  INV_X1 U15316 ( .A(n15479), .ZN(n12198) );
  NAND4_X1 U15317 ( .A1(n15702), .A2(n12199), .A3(n15465), .A4(n12198), .ZN(
        n12204) );
  INV_X1 U15318 ( .A(n12200), .ZN(n12203) );
  NAND3_X1 U15319 ( .A1(n12201), .A2(P2_EBX_REG_15__SCAN_IN), .A3(n9720), .ZN(
        n12202) );
  NAND2_X1 U15320 ( .A1(n12203), .A2(n12202), .ZN(n19280) );
  NOR2_X1 U15321 ( .A1(n12101), .A2(n19280), .ZN(n12207) );
  NOR2_X1 U15322 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n12207), .ZN(
        n16427) );
  NOR2_X1 U15323 ( .A1(n12204), .A2(n16427), .ZN(n12205) );
  NOR2_X1 U15324 ( .A1(n15696), .A2(n12206), .ZN(n15703) );
  AND2_X1 U15325 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n12207), .ZN(
        n16426) );
  OR2_X1 U15326 ( .A1(n15703), .A2(n16426), .ZN(n15456) );
  NOR2_X1 U15327 ( .A1(n12101), .A2(n15470), .ZN(n12208) );
  NAND2_X1 U15328 ( .A1(n15167), .A2(n12208), .ZN(n15466) );
  NAND2_X1 U15329 ( .A1(n12209), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15500) );
  INV_X1 U15330 ( .A(n12210), .ZN(n12211) );
  NAND2_X1 U15331 ( .A1(n12211), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15461) );
  OR2_X1 U15332 ( .A1(n12101), .A2(n15679), .ZN(n12212) );
  OR2_X1 U15333 ( .A1(n19252), .A2(n12212), .ZN(n15462) );
  OR2_X1 U15334 ( .A1(n12213), .A2(n16536), .ZN(n16449) );
  AND4_X1 U15335 ( .A1(n15500), .A2(n15461), .A3(n15462), .A4(n16449), .ZN(
        n12216) );
  OR2_X1 U15336 ( .A1(n12214), .A2(n15636), .ZN(n15478) );
  NAND2_X1 U15337 ( .A1(n12215), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15489) );
  NAND4_X1 U15338 ( .A1(n15466), .A2(n12216), .A3(n15478), .A4(n15489), .ZN(
        n12217) );
  NOR2_X1 U15339 ( .A1(n15456), .A2(n12217), .ZN(n12218) );
  INV_X1 U15340 ( .A(n12219), .ZN(n12220) );
  NAND2_X1 U15341 ( .A1(n12221), .A2(n12220), .ZN(n12222) );
  NAND2_X1 U15342 ( .A1(n12227), .A2(n12222), .ZN(n15166) );
  OR2_X1 U15343 ( .A1(n15166), .A2(n12101), .ZN(n12223) );
  INV_X1 U15344 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15619) );
  NAND2_X1 U15345 ( .A1(n12223), .A2(n15619), .ZN(n15447) );
  NAND2_X1 U15346 ( .A1(n15445), .A2(n15447), .ZN(n12225) );
  OR2_X1 U15347 ( .A1(n12101), .A2(n15619), .ZN(n12224) );
  OR2_X1 U15348 ( .A1(n15166), .A2(n12224), .ZN(n15446) );
  INV_X1 U15349 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15436) );
  XNOR2_X1 U15350 ( .A(n12228), .B(n15436), .ZN(n15435) );
  INV_X1 U15351 ( .A(n15151), .ZN(n12229) );
  NAND2_X1 U15352 ( .A1(n9720), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12231) );
  MUX2_X1 U15353 ( .A(n12231), .B(P2_EBX_REG_24__SCAN_IN), .S(n12230), .Z(
        n12232) );
  NAND2_X1 U15354 ( .A1(n12232), .A2(n12235), .ZN(n16372) );
  INV_X1 U15355 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15610) );
  NAND2_X1 U15356 ( .A1(n9720), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12234) );
  MUX2_X1 U15357 ( .A(n12234), .B(P2_EBX_REG_25__SCAN_IN), .S(n12233), .Z(
        n12236) );
  AOI21_X1 U15358 ( .B1(n16359), .B2(n12162), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15597) );
  INV_X1 U15359 ( .A(n15597), .ZN(n12237) );
  NAND2_X1 U15360 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n12238), .ZN(n12239) );
  NOR2_X1 U15361 ( .A1(n10855), .A2(n12239), .ZN(n12240) );
  NOR2_X1 U15362 ( .A1(n12890), .A2(n12240), .ZN(n16348) );
  NAND2_X1 U15363 ( .A1(n16348), .A2(n12162), .ZN(n12254) );
  INV_X1 U15364 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15588) );
  XNOR2_X1 U15365 ( .A(n12254), .B(n15588), .ZN(n15417) );
  INV_X1 U15366 ( .A(n12241), .ZN(n12243) );
  NAND2_X1 U15367 ( .A1(n12243), .A2(n12242), .ZN(n12244) );
  AND2_X1 U15368 ( .A1(n12250), .A2(n12244), .ZN(n16337) );
  NAND2_X1 U15369 ( .A1(n16337), .A2(n12162), .ZN(n15393) );
  NOR2_X1 U15370 ( .A1(n15388), .A2(n12247), .ZN(n12256) );
  INV_X1 U15371 ( .A(n12248), .ZN(n12249) );
  NAND2_X1 U15372 ( .A1(n12250), .A2(n12249), .ZN(n12251) );
  AND2_X1 U15373 ( .A1(n12257), .A2(n12251), .ZN(n16330) );
  NAND2_X1 U15374 ( .A1(n16330), .A2(n12162), .ZN(n15396) );
  AND2_X1 U15375 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15559) );
  INV_X1 U15376 ( .A(n16359), .ZN(n12253) );
  INV_X1 U15377 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15604) );
  OR2_X1 U15378 ( .A1(n12101), .A2(n15604), .ZN(n12252) );
  OR2_X1 U15379 ( .A1(n12254), .A2(n15588), .ZN(n12255) );
  NAND2_X1 U15380 ( .A1(n15595), .A2(n12255), .ZN(n15391) );
  XOR2_X1 U15381 ( .A(n12258), .B(n12257), .Z(n12259) );
  INV_X1 U15382 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15550) );
  OAI21_X1 U15383 ( .B1(n12259), .B2(n12101), .A(n15550), .ZN(n15376) );
  NAND2_X1 U15384 ( .A1(n15377), .A2(n15376), .ZN(n12889) );
  INV_X1 U15385 ( .A(n12259), .ZN(n16313) );
  NAND3_X1 U15386 ( .A1(n16313), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12162), .ZN(n15375) );
  NAND2_X1 U15387 ( .A1(n12889), .A2(n15375), .ZN(n12263) );
  AOI21_X1 U15388 ( .B1(n12260), .B2(n12162), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12888) );
  INV_X1 U15389 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12527) );
  INV_X1 U15390 ( .A(n12887), .ZN(n12262) );
  AND2_X1 U15391 ( .A1(n12030), .A2(n16615), .ZN(n20205) );
  NAND2_X1 U15392 ( .A1(n12266), .A2(n12265), .ZN(n12455) );
  NAND2_X1 U15393 ( .A1(n12267), .A2(n12455), .ZN(n12268) );
  NAND2_X1 U15394 ( .A1(n12268), .A2(n12458), .ZN(n20185) );
  NAND3_X1 U15395 ( .A1(n20189), .A2(n20184), .A3(n20185), .ZN(n12277) );
  NAND2_X1 U15396 ( .A1(n9694), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12271) );
  INV_X1 U15397 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12270) );
  NAND2_X1 U15398 ( .A1(n12271), .A2(n12270), .ZN(n13353) );
  NOR2_X1 U15399 ( .A1(n15777), .A2(P2_FLUSH_REG_SCAN_IN), .ZN(n12272) );
  OAI21_X1 U15400 ( .B1(n10506), .B2(n13353), .A(n12272), .ZN(n20173) );
  OAI21_X1 U15401 ( .B1(n12448), .B2(n12273), .A(n16608), .ZN(n12274) );
  NAND2_X1 U15402 ( .A1(n15777), .A2(n12274), .ZN(n12275) );
  NAND3_X1 U15403 ( .A1(n16616), .A2(n16628), .A3(n10648), .ZN(n12276) );
  NAND2_X1 U15404 ( .A1(n12277), .A2(n12276), .ZN(n12467) );
  NAND2_X1 U15405 ( .A1(n12539), .A2(n12279), .ZN(n12328) );
  INV_X1 U15406 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12286) );
  NAND2_X1 U15407 ( .A1(n12281), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16588) );
  INV_X1 U15408 ( .A(n16588), .ZN(n12283) );
  XNOR2_X1 U15409 ( .A(n12282), .B(n16586), .ZN(n12284) );
  NAND2_X1 U15410 ( .A1(n12283), .A2(n12284), .ZN(n12285) );
  XNOR2_X1 U15411 ( .A(n16588), .B(n12284), .ZN(n13329) );
  NAND2_X1 U15412 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13329), .ZN(
        n13330) );
  NAND2_X1 U15413 ( .A1(n12285), .A2(n13330), .ZN(n12290) );
  XNOR2_X1 U15414 ( .A(n12286), .B(n12290), .ZN(n13366) );
  INV_X1 U15415 ( .A(n12287), .ZN(n12288) );
  XOR2_X1 U15416 ( .A(n12289), .B(n12288), .Z(n13365) );
  NAND2_X1 U15417 ( .A1(n13366), .A2(n13365), .ZN(n13364) );
  NAND2_X1 U15418 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12290), .ZN(
        n12291) );
  NAND2_X1 U15419 ( .A1(n13364), .A2(n12291), .ZN(n12292) );
  XNOR2_X1 U15420 ( .A(n12292), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14025) );
  NAND2_X1 U15421 ( .A1(n12292), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12293) );
  NAND2_X1 U15422 ( .A1(n19493), .A2(n19520), .ZN(n12296) );
  INV_X1 U15423 ( .A(n19493), .ZN(n12297) );
  INV_X1 U15424 ( .A(n12298), .ZN(n12299) );
  NAND2_X1 U15425 ( .A1(n12299), .A2(n16582), .ZN(n16499) );
  NAND2_X1 U15426 ( .A1(n10167), .A2(n16497), .ZN(n12301) );
  NAND2_X1 U15427 ( .A1(n12301), .A2(n12300), .ZN(n12304) );
  NAND2_X1 U15428 ( .A1(n12305), .A2(n12302), .ZN(n12303) );
  NAND2_X1 U15429 ( .A1(n14343), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14342) );
  INV_X1 U15430 ( .A(n12305), .ZN(n16501) );
  NAND2_X1 U15431 ( .A1(n16497), .A2(n16501), .ZN(n12307) );
  NAND2_X1 U15432 ( .A1(n12307), .A2(n9951), .ZN(n12308) );
  XNOR2_X1 U15433 ( .A(n12309), .B(n12101), .ZN(n15764) );
  OAI21_X1 U15434 ( .B1(n12309), .B2(n12101), .A(n12310), .ZN(n12313) );
  INV_X1 U15435 ( .A(n12309), .ZN(n12312) );
  NOR2_X1 U15436 ( .A1(n12101), .A2(n12310), .ZN(n12311) );
  AND2_X1 U15437 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15628) );
  INV_X1 U15438 ( .A(n15628), .ZN(n16551) );
  NAND3_X1 U15439 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15659) );
  INV_X1 U15440 ( .A(n15659), .ZN(n12315) );
  NAND2_X1 U15441 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n12315), .ZN(
        n15635) );
  NAND2_X1 U15442 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12316) );
  NOR2_X1 U15443 ( .A1(n15635), .A2(n12316), .ZN(n12317) );
  AND3_X1 U15444 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15634) );
  AND2_X1 U15445 ( .A1(n12317), .A2(n15634), .ZN(n16047) );
  INV_X1 U15446 ( .A(n16047), .ZN(n12318) );
  NAND2_X1 U15447 ( .A1(n15409), .A2(n15559), .ZN(n15399) );
  NOR2_X2 U15448 ( .A1(n15399), .A2(n15550), .ZN(n15383) );
  XNOR2_X1 U15449 ( .A(n15383), .B(n12527), .ZN(n12536) );
  INV_X1 U15450 ( .A(n13269), .ZN(n12319) );
  NOR2_X1 U15451 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15799) );
  OR2_X1 U15452 ( .A1(n20157), .A2(n15799), .ZN(n20164) );
  NAND2_X1 U15453 ( .A1(n20164), .A2(n20201), .ZN(n12320) );
  NAND2_X1 U15454 ( .A1(n19595), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12321) );
  NAND2_X1 U15455 ( .A1(n12553), .A2(n12321), .ZN(n19502) );
  NOR2_X1 U15456 ( .A1(n19324), .A2(n20133), .ZN(n12526) );
  INV_X1 U15457 ( .A(n12526), .ZN(n12324) );
  AND2_X1 U15458 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20165) );
  NOR2_X1 U15459 ( .A1(n12322), .A2(n16436), .ZN(n12323) );
  NAND2_X1 U15460 ( .A1(n12328), .A2(n12327), .ZN(P2_U2984) );
  INV_X1 U15461 ( .A(n12400), .ZN(n12389) );
  NAND2_X1 U15462 ( .A1(n12329), .A2(n12389), .ZN(n12335) );
  NAND2_X1 U15463 ( .A1(n12341), .A2(n12340), .ZN(n12330) );
  NAND2_X1 U15464 ( .A1(n12330), .A2(n12331), .ZN(n12362) );
  OAI21_X1 U15465 ( .B1(n12331), .B2(n12330), .A(n12362), .ZN(n12333) );
  INV_X1 U15466 ( .A(n20910), .ZN(n12405) );
  NAND2_X1 U15467 ( .A1(n13989), .A2(n13812), .ZN(n12336) );
  INV_X1 U15468 ( .A(n12336), .ZN(n12332) );
  AOI21_X1 U15469 ( .B1(n12333), .B2(n12405), .A(n12332), .ZN(n12334) );
  NAND2_X1 U15470 ( .A1(n12335), .A2(n12334), .ZN(n13607) );
  OAI21_X1 U15471 ( .B1(n20910), .B2(n12341), .A(n12336), .ZN(n12337) );
  INV_X1 U15472 ( .A(n12337), .ZN(n12338) );
  XNOR2_X1 U15473 ( .A(n12341), .B(n12340), .ZN(n12343) );
  OAI211_X1 U15474 ( .C1(n12343), .C2(n20910), .A(n12342), .B(n9710), .ZN(
        n12344) );
  INV_X1 U15475 ( .A(n12344), .ZN(n12345) );
  NAND2_X1 U15476 ( .A1(n13570), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12350) );
  INV_X1 U15477 ( .A(n12347), .ZN(n12348) );
  OR2_X1 U15478 ( .A1(n13489), .A2(n12348), .ZN(n12349) );
  INV_X1 U15479 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12351) );
  NAND2_X1 U15480 ( .A1(n13607), .A2(n13606), .ZN(n12354) );
  NAND2_X1 U15481 ( .A1(n12352), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12353) );
  XNOR2_X1 U15482 ( .A(n12362), .B(n12361), .ZN(n12356) );
  OAI22_X1 U15483 ( .A1(n15112), .A2(n12400), .B1(n20910), .B2(n12356), .ZN(
        n13778) );
  NAND2_X1 U15484 ( .A1(n13777), .A2(n13778), .ZN(n12359) );
  NAND2_X1 U15485 ( .A1(n12357), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12358) );
  NAND2_X1 U15486 ( .A1(n12360), .A2(n12389), .ZN(n12368) );
  NAND2_X1 U15487 ( .A1(n12362), .A2(n12361), .ZN(n12364) );
  INV_X1 U15488 ( .A(n12364), .ZN(n12366) );
  INV_X1 U15489 ( .A(n12365), .ZN(n12363) );
  OR2_X1 U15490 ( .A1(n12364), .A2(n12363), .ZN(n12381) );
  OAI211_X1 U15491 ( .C1(n12366), .C2(n12365), .A(n12405), .B(n12381), .ZN(
        n12367) );
  NAND2_X1 U15492 ( .A1(n12368), .A2(n12367), .ZN(n12369) );
  INV_X1 U15493 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13938) );
  XNOR2_X1 U15494 ( .A(n12369), .B(n13938), .ZN(n13928) );
  NAND2_X1 U15495 ( .A1(n13929), .A2(n13928), .ZN(n12371) );
  NAND2_X1 U15496 ( .A1(n12369), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12370) );
  NAND2_X2 U15497 ( .A1(n12371), .A2(n12370), .ZN(n14224) );
  INV_X1 U15498 ( .A(n12372), .ZN(n12373) );
  XNOR2_X1 U15499 ( .A(n12381), .B(n12382), .ZN(n12374) );
  NAND2_X1 U15500 ( .A1(n12374), .A2(n12405), .ZN(n12375) );
  INV_X1 U15501 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12377) );
  XNOR2_X1 U15502 ( .A(n12378), .B(n12377), .ZN(n14225) );
  NAND2_X1 U15503 ( .A1(n12378), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12379) );
  NAND3_X1 U15504 ( .A1(n12403), .A2(n12380), .A3(n12389), .ZN(n12386) );
  INV_X1 U15505 ( .A(n12381), .ZN(n12383) );
  NAND2_X1 U15506 ( .A1(n12383), .A2(n12382), .ZN(n12391) );
  XNOR2_X1 U15507 ( .A(n12391), .B(n12392), .ZN(n12384) );
  NAND2_X1 U15508 ( .A1(n12384), .A2(n12405), .ZN(n12385) );
  AND2_X1 U15509 ( .A1(n12386), .A2(n12385), .ZN(n12387) );
  INV_X1 U15510 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16293) );
  NAND2_X1 U15511 ( .A1(n12387), .A2(n16293), .ZN(n16175) );
  INV_X1 U15512 ( .A(n12387), .ZN(n12388) );
  NAND2_X1 U15513 ( .A1(n12388), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16174) );
  NAND2_X1 U15514 ( .A1(n12390), .A2(n12389), .ZN(n12396) );
  INV_X1 U15515 ( .A(n12391), .ZN(n12393) );
  NAND2_X1 U15516 ( .A1(n12393), .A2(n12392), .ZN(n12407) );
  XNOR2_X1 U15517 ( .A(n12407), .B(n12404), .ZN(n12394) );
  NAND2_X1 U15518 ( .A1(n12394), .A2(n12405), .ZN(n12395) );
  NAND2_X1 U15519 ( .A1(n12396), .A2(n12395), .ZN(n16167) );
  OR2_X1 U15520 ( .A1(n16167), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12397) );
  NAND2_X1 U15521 ( .A1(n16169), .A2(n12397), .ZN(n12399) );
  NAND2_X1 U15522 ( .A1(n16167), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12398) );
  NAND2_X2 U15523 ( .A1(n12399), .A2(n12398), .ZN(n14391) );
  NOR2_X1 U15524 ( .A1(n12401), .A2(n12400), .ZN(n12402) );
  NAND2_X1 U15525 ( .A1(n12405), .A2(n12404), .ZN(n12406) );
  AND2_X1 U15526 ( .A1(n14389), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12410) );
  INV_X1 U15527 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12408) );
  INV_X2 U15528 ( .A(n9673), .ZN(n15065) );
  INV_X1 U15529 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16259) );
  NAND2_X1 U15530 ( .A1(n9673), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14905) );
  NAND2_X1 U15531 ( .A1(n15065), .A2(n16245), .ZN(n12411) );
  NAND2_X1 U15532 ( .A1(n14905), .A2(n12411), .ZN(n14922) );
  INV_X1 U15533 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14937) );
  NAND2_X1 U15534 ( .A1(n16158), .A2(n14937), .ZN(n14920) );
  NAND2_X1 U15535 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12412) );
  NAND2_X1 U15536 ( .A1(n15065), .A2(n12412), .ZN(n14917) );
  NAND2_X1 U15537 ( .A1(n14920), .A2(n14917), .ZN(n12413) );
  INV_X1 U15538 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16233) );
  AND2_X1 U15539 ( .A1(n16158), .A2(n16233), .ZN(n12414) );
  NOR2_X1 U15540 ( .A1(n14906), .A2(n12414), .ZN(n16130) );
  OAI21_X1 U15541 ( .B1(n16135), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16130), .ZN(n12415) );
  XNOR2_X1 U15542 ( .A(n15065), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15067) );
  NAND2_X1 U15543 ( .A1(n16158), .A2(n15084), .ZN(n15077) );
  NAND2_X1 U15544 ( .A1(n15067), .A2(n15077), .ZN(n16132) );
  NAND2_X1 U15545 ( .A1(n16135), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12416) );
  NAND2_X1 U15546 ( .A1(n16161), .A2(n16260), .ZN(n14904) );
  OAI21_X1 U15547 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n14904), .A(
        n16135), .ZN(n12417) );
  NAND2_X1 U15548 ( .A1(n16127), .A2(n12417), .ZN(n15062) );
  NOR2_X1 U15549 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15072) );
  AND2_X1 U15550 ( .A1(n15072), .A2(n16137), .ZN(n12418) );
  NOR2_X1 U15551 ( .A1(n15065), .A2(n12418), .ZN(n12419) );
  XNOR2_X1 U15552 ( .A(n15065), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14896) );
  NAND3_X1 U15553 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14943) );
  INV_X1 U15554 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16218) );
  INV_X1 U15555 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15044) );
  NAND2_X1 U15556 ( .A1(n12420), .A2(n16135), .ZN(n14870) );
  AND2_X1 U15557 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15018) );
  AND2_X1 U15558 ( .A1(n15018), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15012) );
  NAND2_X1 U15559 ( .A1(n12424), .A2(n15012), .ZN(n14818) );
  NOR2_X1 U15560 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12421) );
  AND2_X1 U15561 ( .A1(n12421), .A2(n16197), .ZN(n14819) );
  NAND2_X1 U15562 ( .A1(n16135), .A2(n14819), .ZN(n12422) );
  NAND2_X1 U15563 ( .A1(n14818), .A2(n12422), .ZN(n12423) );
  NAND2_X1 U15564 ( .A1(n9663), .A2(n16135), .ZN(n14847) );
  INV_X1 U15565 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15011) );
  INV_X1 U15566 ( .A(n14819), .ZN(n12425) );
  OAI21_X1 U15567 ( .B1(n9664), .B2(n12425), .A(n16135), .ZN(n12426) );
  NOR2_X1 U15568 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14993) );
  NAND2_X1 U15569 ( .A1(n16135), .A2(n14993), .ZN(n12427) );
  INV_X1 U15570 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14983) );
  AND2_X1 U15571 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14984) );
  NAND2_X1 U15572 ( .A1(n15065), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12429) );
  NAND2_X1 U15573 ( .A1(n12913), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12430) );
  NOR2_X1 U15574 ( .A1(n9699), .A2(n20219), .ZN(n12431) );
  NAND2_X1 U15575 ( .A1(n14562), .A2(n12432), .ZN(n12435) );
  AOI22_X1 U15576 ( .A1(n11173), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13843), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12433) );
  XNOR2_X2 U15577 ( .A(n12435), .B(n12434), .ZN(n14539) );
  NAND3_X1 U15578 ( .A1(n20222), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16298) );
  INV_X1 U15579 ( .A(n16298), .ZN(n12436) );
  NAND2_X1 U15580 ( .A1(n14539), .A2(n14887), .ZN(n12445) );
  NAND2_X1 U15581 ( .A1(n20743), .A2(n12441), .ZN(n20905) );
  AND2_X1 U15582 ( .A1(n20905), .A2(n20222), .ZN(n12437) );
  NAND2_X1 U15583 ( .A1(n20222), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16002) );
  NAND2_X1 U15584 ( .A1(n21095), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12438) );
  NAND2_X1 U15585 ( .A1(n16002), .A2(n12438), .ZN(n13491) );
  XNOR2_X1 U15586 ( .A(n12440), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14001) );
  INV_X1 U15587 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21032) );
  NOR2_X1 U15588 ( .A1(n16238), .A2(n21032), .ZN(n14947) );
  AOI21_X1 U15589 ( .B1(n16173), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14947), .ZN(n12442) );
  OAI21_X1 U15590 ( .B1(n16180), .B2(n14001), .A(n12442), .ZN(n12443) );
  INV_X1 U15591 ( .A(n12443), .ZN(n12444) );
  NOR2_X1 U15592 ( .A1(n12463), .A2(n12030), .ZN(n12447) );
  MUX2_X1 U15593 ( .A(n12447), .B(n12537), .S(n12451), .Z(n12457) );
  NAND2_X1 U15594 ( .A1(n12030), .A2(n12448), .ZN(n12450) );
  NAND2_X1 U15595 ( .A1(n12450), .A2(n12449), .ZN(n12453) );
  NAND2_X1 U15596 ( .A1(n12030), .A2(n12451), .ZN(n12452) );
  NAND2_X1 U15597 ( .A1(n12453), .A2(n12452), .ZN(n12454) );
  AOI22_X1 U15598 ( .A1(n12537), .A2(n12455), .B1(n12454), .B2(n20199), .ZN(
        n12456) );
  NOR2_X1 U15599 ( .A1(n12457), .A2(n12456), .ZN(n12459) );
  MUX2_X1 U15600 ( .A(n12537), .B(n12459), .S(n12458), .Z(n12461) );
  INV_X1 U15601 ( .A(n20184), .ZN(n12460) );
  NOR2_X1 U15602 ( .A1(n12461), .A2(n12460), .ZN(n12462) );
  MUX2_X1 U15603 ( .A(n12462), .B(n12270), .S(n20201), .Z(n12466) );
  INV_X1 U15604 ( .A(n13745), .ZN(n16612) );
  NAND2_X1 U15605 ( .A1(n16612), .A2(n10648), .ZN(n13391) );
  OAI211_X1 U15606 ( .C1(n12466), .C2(n16615), .A(n13391), .B(n12465), .ZN(
        n12486) );
  INV_X1 U15607 ( .A(n13391), .ZN(n13342) );
  NAND3_X1 U15608 ( .A1(n13342), .A2(n12492), .A3(n13267), .ZN(n12485) );
  INV_X1 U15609 ( .A(n12467), .ZN(n12483) );
  NAND2_X1 U15610 ( .A1(n12469), .A2(n19565), .ZN(n12470) );
  NAND2_X1 U15611 ( .A1(n12468), .A2(n12470), .ZN(n12479) );
  INV_X1 U15612 ( .A(n12495), .ZN(n12471) );
  OAI21_X1 U15613 ( .B1(n12472), .B2(n9683), .A(n13415), .ZN(n12474) );
  NAND2_X1 U15614 ( .A1(n12474), .A2(n20205), .ZN(n12503) );
  NAND2_X1 U15615 ( .A1(n12465), .A2(n12030), .ZN(n12510) );
  NAND2_X1 U15616 ( .A1(n12510), .A2(n20199), .ZN(n12475) );
  NAND2_X1 U15617 ( .A1(n12475), .A2(n13415), .ZN(n12476) );
  NAND2_X1 U15618 ( .A1(n12476), .A2(n19565), .ZN(n12477) );
  NAND4_X1 U15619 ( .A1(n12479), .A2(n12478), .A3(n12503), .A4(n12477), .ZN(
        n12511) );
  AND3_X1 U15620 ( .A1(n16608), .A2(n10654), .A3(n13267), .ZN(n12480) );
  NOR2_X1 U15621 ( .A1(n12511), .A2(n12480), .ZN(n13346) );
  INV_X1 U15622 ( .A(n20202), .ZN(n20196) );
  NOR2_X1 U15623 ( .A1(n12489), .A2(n20196), .ZN(n12481) );
  OAI211_X1 U15624 ( .C1(n10654), .C2(n12030), .A(n16608), .B(n12481), .ZN(
        n12482) );
  AND3_X1 U15625 ( .A1(n12483), .A2(n13346), .A3(n12482), .ZN(n12484) );
  NAND3_X1 U15626 ( .A1(n12486), .A2(n12485), .A3(n12484), .ZN(n12487) );
  AND2_X1 U15627 ( .A1(n12489), .A2(n12488), .ZN(n12490) );
  NAND2_X1 U15628 ( .A1(n12491), .A2(n12490), .ZN(n12861) );
  NAND2_X1 U15629 ( .A1(n12492), .A2(n16615), .ZN(n12493) );
  AND2_X1 U15630 ( .A1(n12861), .A2(n12493), .ZN(n12500) );
  INV_X1 U15631 ( .A(n12494), .ZN(n13274) );
  OAI21_X1 U15632 ( .B1(n12495), .B2(n12465), .A(n13274), .ZN(n12499) );
  NAND3_X1 U15633 ( .A1(n12497), .A2(n12496), .A3(n12495), .ZN(n12498) );
  AND4_X1 U15634 ( .A1(n12501), .A2(n12500), .A3(n12499), .A4(n12498), .ZN(
        n12507) );
  NAND2_X1 U15635 ( .A1(n12502), .A2(n10648), .ZN(n15771) );
  NAND2_X1 U15636 ( .A1(n15771), .A2(n12503), .ZN(n12505) );
  NAND2_X1 U15637 ( .A1(n12505), .A2(n12504), .ZN(n12506) );
  AND2_X1 U15638 ( .A1(n12507), .A2(n12506), .ZN(n15795) );
  NAND2_X1 U15639 ( .A1(n15795), .A2(n15789), .ZN(n12509) );
  NAND2_X1 U15640 ( .A1(n12538), .A2(n16607), .ZN(n12515) );
  NAND2_X1 U15641 ( .A1(n15559), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12525) );
  NAND2_X1 U15642 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16514) );
  NAND4_X1 U15643 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n15628), .A4(n16047), .ZN(
        n12523) );
  INV_X1 U15644 ( .A(n12523), .ZN(n12518) );
  NOR2_X1 U15645 ( .A1(n19520), .A2(n16582), .ZN(n16571) );
  INV_X1 U15646 ( .A(n16571), .ZN(n14351) );
  NOR2_X1 U15647 ( .A1(n12512), .A2(n14351), .ZN(n12517) );
  NOR2_X1 U15648 ( .A1(n15780), .A2(n16585), .ZN(n19564) );
  NOR2_X1 U15649 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19564), .ZN(
        n19531) );
  NAND2_X1 U15650 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19564), .ZN(
        n12514) );
  OAI22_X1 U15651 ( .A1(n19531), .A2(n12515), .B1(n19533), .B2(n12514), .ZN(
        n14027) );
  NAND2_X1 U15652 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14027), .ZN(
        n19521) );
  INV_X1 U15653 ( .A(n19521), .ZN(n12513) );
  NAND2_X1 U15654 ( .A1(n12517), .A2(n12513), .ZN(n12522) );
  AOI21_X1 U15655 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n12522), .ZN(n16561) );
  INV_X1 U15656 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14028) );
  INV_X1 U15657 ( .A(n12514), .ZN(n19532) );
  INV_X1 U15658 ( .A(n12515), .ZN(n19535) );
  NOR2_X1 U15659 ( .A1(n12538), .A2(n19517), .ZN(n19552) );
  AOI21_X1 U15660 ( .B1(n19535), .B2(n19531), .A(n19552), .ZN(n12516) );
  OAI21_X1 U15661 ( .B1(n19532), .B2(n19533), .A(n12516), .ZN(n14029) );
  AOI21_X1 U15662 ( .B1(n14028), .B2(n19549), .A(n14029), .ZN(n19519) );
  OAI21_X1 U15663 ( .B1(n16593), .B2(n12517), .A(n19519), .ZN(n16565) );
  NOR2_X1 U15664 ( .A1(n16561), .A2(n16565), .ZN(n15748) );
  OAI21_X1 U15665 ( .B1(n16593), .B2(n12518), .A(n15748), .ZN(n16509) );
  AOI21_X1 U15666 ( .B1(n16514), .B2(n19549), .A(n16509), .ZN(n15609) );
  INV_X1 U15667 ( .A(n15609), .ZN(n12519) );
  AOI21_X1 U15668 ( .B1(n15610), .B2(n19549), .A(n12519), .ZN(n15605) );
  OAI21_X1 U15669 ( .B1(n9834), .B2(n16593), .A(n15605), .ZN(n15577) );
  AOI21_X1 U15670 ( .B1(n19549), .B2(n12525), .A(n15577), .ZN(n14498) );
  NOR2_X1 U15671 ( .A1(n14498), .A2(n12527), .ZN(n12535) );
  NAND2_X1 U15672 ( .A1(n15803), .A2(n12030), .ZN(n12520) );
  NAND2_X1 U15673 ( .A1(n12520), .A2(n10705), .ZN(n12521) );
  AND2_X1 U15674 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15584) );
  INV_X1 U15675 ( .A(n12522), .ZN(n15761) );
  NAND3_X1 U15676 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(n15761), .ZN(n15750) );
  NOR2_X1 U15677 ( .A1(n12523), .A2(n15750), .ZN(n16515) );
  NAND3_X1 U15678 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n16515), .ZN(n15611) );
  INV_X1 U15679 ( .A(n15611), .ZN(n15587) );
  AND2_X1 U15680 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15587), .ZN(
        n12524) );
  NAND2_X1 U15681 ( .A1(n15584), .A2(n12524), .ZN(n15549) );
  NOR2_X1 U15682 ( .A1(n15549), .A2(n12525), .ZN(n14508) );
  AOI21_X1 U15683 ( .B1(n14508), .B2(n12527), .A(n12526), .ZN(n12533) );
  AND2_X1 U15684 ( .A1(n12528), .A2(n10718), .ZN(n16613) );
  INV_X1 U15685 ( .A(n16613), .ZN(n12530) );
  NAND2_X1 U15686 ( .A1(n9659), .A2(n10648), .ZN(n12529) );
  NAND2_X1 U15687 ( .A1(n12530), .A2(n12529), .ZN(n12531) );
  NAND2_X1 U15688 ( .A1(n19537), .A2(n12880), .ZN(n12532) );
  OAI211_X1 U15689 ( .C1(n12322), .C2(n19540), .A(n12533), .B(n12532), .ZN(
        n12534) );
  AOI211_X1 U15690 ( .C1(n12536), .C2(n16577), .A(n12535), .B(n12534), .ZN(
        n12541) );
  AND2_X1 U15691 ( .A1(n16616), .A2(n12537), .ZN(n20187) );
  NAND2_X1 U15692 ( .A1(n12539), .A2(n19551), .ZN(n12540) );
  NAND2_X1 U15693 ( .A1(n12541), .A2(n12540), .ZN(P2_U3016) );
  NAND2_X1 U15694 ( .A1(n12549), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12542) );
  NAND2_X1 U15695 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19991) );
  INV_X1 U15696 ( .A(n19991), .ZN(n12543) );
  NAND2_X1 U15697 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12543), .ZN(
        n12563) );
  INV_X1 U15698 ( .A(n12563), .ZN(n12544) );
  NAND2_X1 U15699 ( .A1(n12544), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19993) );
  NAND2_X1 U15700 ( .A1(n20156), .A2(n12563), .ZN(n12545) );
  AND3_X1 U15701 ( .A1(n19993), .A2(n20157), .A3(n12545), .ZN(n12546) );
  AOI21_X1 U15702 ( .B1(n12566), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12546), .ZN(n12547) );
  OAI21_X2 U15703 ( .B1(n12548), .B2(n12553), .A(n12547), .ZN(n12574) );
  OAI21_X1 U15704 ( .B1(n12574), .B2(n12551), .A(n13950), .ZN(n12552) );
  NAND2_X1 U15705 ( .A1(n12566), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12554) );
  NAND2_X1 U15706 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10356), .ZN(
        n19819) );
  NAND2_X1 U15707 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20182), .ZN(
        n19850) );
  NAND2_X1 U15708 ( .A1(n19819), .A2(n19850), .ZN(n14173) );
  NAND2_X1 U15709 ( .A1(n20157), .A2(n14173), .ZN(n19853) );
  NAND2_X1 U15710 ( .A1(n12554), .A2(n19853), .ZN(n12555) );
  AOI22_X1 U15711 ( .A1(n12566), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20157), .B2(n20182), .ZN(n12557) );
  NAND2_X1 U15712 ( .A1(n12797), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12559) );
  INV_X1 U15713 ( .A(n12559), .ZN(n12560) );
  NOR2_X1 U15714 ( .A1(n13418), .A2(n12560), .ZN(n12561) );
  NAND2_X1 U15715 ( .A1(n9714), .A2(n12562), .ZN(n12568) );
  NAND2_X1 U15716 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19755) );
  NAND2_X1 U15717 ( .A1(n19755), .A2(n20163), .ZN(n12564) );
  NAND2_X1 U15718 ( .A1(n12564), .A2(n12563), .ZN(n13957) );
  NOR2_X1 U15719 ( .A1(n20150), .A2(n13957), .ZN(n12565) );
  AOI21_X1 U15720 ( .B1(n12566), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12565), .ZN(n12567) );
  NAND3_X1 U15721 ( .A1(n13470), .A2(n13478), .A3(n13465), .ZN(n12573) );
  NAND2_X1 U15722 ( .A1(n13470), .A2(n13466), .ZN(n12572) );
  NAND2_X1 U15723 ( .A1(n12549), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12571) );
  INV_X1 U15724 ( .A(n19405), .ZN(n12577) );
  NAND2_X1 U15725 ( .A1(n14013), .A2(n14016), .ZN(n12578) );
  AOI22_X1 U15726 ( .A1(n12620), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12583) );
  AOI22_X1 U15727 ( .A1(n9718), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12582) );
  AOI22_X1 U15728 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12581) );
  AOI22_X1 U15729 ( .A1(n10513), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15815), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12580) );
  NAND4_X1 U15730 ( .A1(n12583), .A2(n12582), .A3(n12581), .A4(n12580), .ZN(
        n12589) );
  AOI22_X1 U15731 ( .A1(n12675), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12587) );
  AOI22_X1 U15732 ( .A1(n12676), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12586) );
  AOI22_X1 U15733 ( .A1(n10505), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U15734 ( .A1(n12678), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12584) );
  NAND4_X1 U15735 ( .A1(n12587), .A2(n12586), .A3(n12585), .A4(n12584), .ZN(
        n12588) );
  OR2_X1 U15736 ( .A1(n12589), .A2(n12588), .ZN(n14301) );
  AOI22_X1 U15737 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10360), .B1(
        n12620), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12593) );
  AOI22_X1 U15738 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n9718), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12592) );
  AOI22_X1 U15739 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10397), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U15740 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10513), .B1(
        n15815), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12590) );
  NAND4_X1 U15741 ( .A1(n12593), .A2(n12592), .A3(n12591), .A4(n12590), .ZN(
        n12599) );
  AOI22_X1 U15742 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12675), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12597) );
  AOI22_X1 U15743 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12676), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12596) );
  AOI22_X1 U15744 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n10505), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U15745 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n12678), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12594) );
  NAND4_X1 U15746 ( .A1(n12597), .A2(n12596), .A3(n12595), .A4(n12594), .ZN(
        n12598) );
  NOR2_X1 U15747 ( .A1(n12599), .A2(n12598), .ZN(n15362) );
  AOI22_X1 U15748 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10360), .B1(
        n12620), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12603) );
  AOI22_X1 U15749 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n9718), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12602) );
  AOI22_X1 U15750 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10397), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12601) );
  AOI22_X1 U15751 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10513), .B1(
        n15815), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12600) );
  NAND4_X1 U15752 ( .A1(n12603), .A2(n12602), .A3(n12601), .A4(n12600), .ZN(
        n12609) );
  AOI22_X1 U15753 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12676), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12607) );
  AOI22_X1 U15754 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12675), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12606) );
  AOI22_X1 U15755 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n10505), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12605) );
  AOI22_X1 U15756 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12678), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12604) );
  NAND4_X1 U15757 ( .A1(n12607), .A2(n12606), .A3(n12605), .A4(n12604), .ZN(
        n12608) );
  NOR2_X1 U15758 ( .A1(n12609), .A2(n12608), .ZN(n14421) );
  AOI22_X1 U15759 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10360), .B1(
        n12620), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12613) );
  AOI22_X1 U15760 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n9717), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12612) );
  AOI22_X1 U15761 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10397), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12611) );
  AOI22_X1 U15762 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10513), .B1(
        n15815), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12610) );
  NAND4_X1 U15763 ( .A1(n12613), .A2(n12612), .A3(n12611), .A4(n12610), .ZN(
        n12619) );
  AOI22_X1 U15764 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12675), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12617) );
  AOI22_X1 U15765 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12676), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12616) );
  AOI22_X1 U15766 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10505), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12615) );
  AOI22_X1 U15767 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12678), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12614) );
  NAND4_X1 U15768 ( .A1(n12617), .A2(n12616), .A3(n12615), .A4(n12614), .ZN(
        n12618) );
  OR2_X1 U15769 ( .A1(n12619), .A2(n12618), .ZN(n14363) );
  AOI22_X1 U15770 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10360), .B1(
        n12620), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12624) );
  AOI22_X1 U15771 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n9718), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12623) );
  AOI22_X1 U15772 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10397), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12622) );
  AOI22_X1 U15773 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10513), .B1(
        n15815), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12621) );
  NAND4_X1 U15774 ( .A1(n12624), .A2(n12623), .A3(n12622), .A4(n12621), .ZN(
        n12630) );
  AOI22_X1 U15775 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12675), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12628) );
  AOI22_X1 U15776 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12676), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12627) );
  AOI22_X1 U15777 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n10505), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12626) );
  AOI22_X1 U15778 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n12678), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12625) );
  NAND4_X1 U15779 ( .A1(n12628), .A2(n12627), .A3(n12626), .A4(n12625), .ZN(
        n12629) );
  OR2_X1 U15780 ( .A1(n12630), .A2(n12629), .ZN(n14397) );
  NAND2_X1 U15781 ( .A1(n14363), .A2(n14397), .ZN(n12631) );
  OAI22_X1 U15782 ( .A1(n12635), .A2(n12634), .B1(n12633), .B2(n12632), .ZN(
        n12649) );
  OAI22_X1 U15783 ( .A1(n12639), .A2(n12638), .B1(n12637), .B2(n12636), .ZN(
        n12648) );
  OAI22_X1 U15784 ( .A1(n12642), .A2(n12641), .B1(n12640), .B2(n14170), .ZN(
        n12647) );
  OAI22_X1 U15785 ( .A1(n12645), .A2(n12644), .B1(n12643), .B2(n14197), .ZN(
        n12646) );
  NOR4_X1 U15786 ( .A1(n12649), .A2(n12648), .A3(n12647), .A4(n12646), .ZN(
        n12660) );
  AOI22_X1 U15787 ( .A1(n12620), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10360), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12659) );
  AOI22_X1 U15788 ( .A1(n9717), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12658) );
  NOR2_X1 U15789 ( .A1(n12651), .A2(n12650), .ZN(n12656) );
  OAI22_X1 U15790 ( .A1(n12654), .A2(n9995), .B1(n12653), .B2(n12652), .ZN(
        n12655) );
  AOI211_X1 U15791 ( .C1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .C2(n10397), .A(
        n12656), .B(n12655), .ZN(n12657) );
  NAND4_X1 U15792 ( .A1(n12660), .A2(n12659), .A3(n12658), .A4(n12657), .ZN(
        n15281) );
  AOI22_X1 U15793 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10360), .B1(
        n12620), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12664) );
  AOI22_X1 U15794 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n9718), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U15795 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10397), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12662) );
  AOI22_X1 U15796 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10513), .B1(
        n15815), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12661) );
  NAND4_X1 U15797 ( .A1(n12664), .A2(n12663), .A3(n12662), .A4(n12661), .ZN(
        n12670) );
  AOI22_X1 U15798 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12675), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12668) );
  AOI22_X1 U15799 ( .A1(n12676), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12667) );
  AOI22_X1 U15800 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10505), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12666) );
  AOI22_X1 U15801 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12678), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12665) );
  NAND4_X1 U15802 ( .A1(n12668), .A2(n12667), .A3(n12666), .A4(n12665), .ZN(
        n12669) );
  NOR2_X1 U15803 ( .A1(n12670), .A2(n12669), .ZN(n15345) );
  AOI22_X1 U15804 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n9717), .B1(
        n12620), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12674) );
  AOI22_X1 U15805 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10360), .B1(
        n10348), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12673) );
  AOI22_X1 U15806 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10397), .B1(
        n10513), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12672) );
  AOI22_X1 U15807 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n15815), .B1(
        n10514), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12671) );
  NAND4_X1 U15808 ( .A1(n12674), .A2(n12673), .A3(n12672), .A4(n12671), .ZN(
        n12684) );
  AOI22_X1 U15809 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12675), .B1(
        n10507), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12682) );
  AOI22_X1 U15810 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12676), .B1(
        n10505), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12681) );
  AOI22_X1 U15811 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n12677), .B1(
        n10506), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12680) );
  AOI22_X1 U15812 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12678), .B1(
        n10508), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12679) );
  NAND4_X1 U15813 ( .A1(n12682), .A2(n12681), .A3(n12680), .A4(n12679), .ZN(
        n12683) );
  NOR2_X1 U15814 ( .A1(n12684), .A2(n12683), .ZN(n12702) );
  INV_X1 U15815 ( .A(n12702), .ZN(n12701) );
  AOI22_X1 U15816 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12691) );
  AOI22_X1 U15817 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12690) );
  NAND2_X1 U15818 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12688) );
  NAND2_X1 U15819 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12687) );
  NAND2_X1 U15820 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12686) );
  NAND2_X1 U15821 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12685) );
  AND4_X1 U15822 ( .A1(n12688), .A2(n12687), .A3(n12686), .A4(n12685), .ZN(
        n12689) );
  XNOR2_X1 U15823 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12846) );
  NAND4_X1 U15824 ( .A1(n12691), .A2(n12690), .A3(n12689), .A4(n12846), .ZN(
        n12700) );
  AOI22_X1 U15825 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12698) );
  INV_X1 U15826 ( .A(n12846), .ZN(n12852) );
  AOI22_X1 U15827 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12697) );
  NAND2_X1 U15828 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12695) );
  NAND2_X1 U15829 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12694) );
  NAND2_X1 U15830 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12693) );
  NAND2_X1 U15831 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12692) );
  AND4_X1 U15832 ( .A1(n12695), .A2(n12694), .A3(n12693), .A4(n12692), .ZN(
        n12696) );
  NAND4_X1 U15833 ( .A1(n12698), .A2(n12852), .A3(n12697), .A4(n12696), .ZN(
        n12699) );
  NAND2_X1 U15834 ( .A1(n12700), .A2(n12699), .ZN(n12729) );
  INV_X1 U15835 ( .A(n12729), .ZN(n12705) );
  NAND2_X1 U15836 ( .A1(n12701), .A2(n12705), .ZN(n12708) );
  OAI21_X1 U15837 ( .B1(n12030), .B2(n12729), .A(n12702), .ZN(n12703) );
  OAI21_X1 U15838 ( .B1(n12708), .B2(n12030), .A(n12703), .ZN(n12730) );
  NAND2_X1 U15839 ( .A1(n12030), .A2(n12705), .ZN(n16391) );
  AND2_X1 U15840 ( .A1(n15344), .A2(n12704), .ZN(n12707) );
  INV_X1 U15841 ( .A(n12708), .ZN(n12727) );
  AOI22_X1 U15842 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12715) );
  AOI22_X1 U15843 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12714) );
  NAND2_X1 U15844 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12712) );
  NAND2_X1 U15845 ( .A1(n9709), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12711) );
  NAND2_X1 U15846 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12710) );
  NAND2_X1 U15847 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12709) );
  AND4_X1 U15848 ( .A1(n12712), .A2(n12711), .A3(n12710), .A4(n12709), .ZN(
        n12713) );
  NAND4_X1 U15849 ( .A1(n12715), .A2(n12714), .A3(n12713), .A4(n12846), .ZN(
        n12726) );
  AOI22_X1 U15850 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12724) );
  AOI22_X1 U15851 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12723) );
  NAND2_X1 U15852 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12721) );
  NAND2_X1 U15853 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12720) );
  NAND2_X1 U15854 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12719) );
  NAND2_X1 U15855 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12718) );
  AND4_X1 U15856 ( .A1(n12721), .A2(n12720), .A3(n12719), .A4(n12718), .ZN(
        n12722) );
  NAND4_X1 U15857 ( .A1(n12724), .A2(n12852), .A3(n12723), .A4(n12722), .ZN(
        n12725) );
  AND2_X1 U15858 ( .A1(n12726), .A2(n12725), .ZN(n12728) );
  NAND2_X1 U15859 ( .A1(n12727), .A2(n12728), .ZN(n12732) );
  OAI211_X1 U15860 ( .C1(n12727), .C2(n12728), .A(n12797), .B(n12732), .ZN(
        n16382) );
  NAND2_X1 U15861 ( .A1(n12030), .A2(n12728), .ZN(n16384) );
  NOR3_X1 U15862 ( .A1(n12730), .A2(n12729), .A3(n16384), .ZN(n12731) );
  INV_X1 U15863 ( .A(n12732), .ZN(n12750) );
  AOI22_X1 U15864 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12740) );
  AOI22_X1 U15865 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12739) );
  NAND2_X1 U15866 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12737) );
  NAND2_X1 U15867 ( .A1(n9709), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12736) );
  NAND2_X1 U15868 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12735) );
  NAND2_X1 U15869 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n12734) );
  AND4_X1 U15870 ( .A1(n12737), .A2(n12736), .A3(n12735), .A4(n12734), .ZN(
        n12738) );
  NAND4_X1 U15871 ( .A1(n12740), .A2(n12739), .A3(n12738), .A4(n12846), .ZN(
        n12749) );
  AOI22_X1 U15872 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12747) );
  AOI22_X1 U15873 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12746) );
  NAND2_X1 U15874 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12744) );
  NAND2_X1 U15875 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12743) );
  NAND2_X1 U15876 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12742) );
  NAND2_X1 U15877 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12741) );
  AND4_X1 U15878 ( .A1(n12744), .A2(n12743), .A3(n12742), .A4(n12741), .ZN(
        n12745) );
  NAND4_X1 U15879 ( .A1(n12747), .A2(n12852), .A3(n12746), .A4(n12745), .ZN(
        n12748) );
  AND2_X1 U15880 ( .A1(n12749), .A2(n12748), .ZN(n12751) );
  NAND2_X1 U15881 ( .A1(n12750), .A2(n12751), .ZN(n12774) );
  OAI211_X1 U15882 ( .C1(n12750), .C2(n12751), .A(n12797), .B(n12774), .ZN(
        n12755) );
  NAND2_X1 U15883 ( .A1(n12030), .A2(n12751), .ZN(n15272) );
  NAND2_X1 U15884 ( .A1(n12753), .A2(n12752), .ZN(n15274) );
  AOI22_X1 U15885 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12763) );
  AOI22_X1 U15886 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12762) );
  NAND2_X1 U15887 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12760) );
  NAND2_X1 U15888 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12759) );
  NAND2_X1 U15889 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12758) );
  NAND2_X1 U15890 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12757) );
  AND4_X1 U15891 ( .A1(n12760), .A2(n12759), .A3(n12758), .A4(n12757), .ZN(
        n12761) );
  NAND4_X1 U15892 ( .A1(n12763), .A2(n12762), .A3(n12761), .A4(n12846), .ZN(
        n12772) );
  AOI22_X1 U15893 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12770) );
  AOI22_X1 U15894 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12769) );
  NAND2_X1 U15895 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12767) );
  NAND2_X1 U15896 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12766) );
  NAND2_X1 U15897 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12765) );
  NAND2_X1 U15898 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12764) );
  AND4_X1 U15899 ( .A1(n12767), .A2(n12766), .A3(n12765), .A4(n12764), .ZN(
        n12768) );
  NAND4_X1 U15900 ( .A1(n12770), .A2(n12852), .A3(n12769), .A4(n12768), .ZN(
        n12771) );
  NAND2_X1 U15901 ( .A1(n12772), .A2(n12771), .ZN(n12776) );
  INV_X1 U15902 ( .A(n12797), .ZN(n12773) );
  AOI21_X1 U15903 ( .B1(n12774), .B2(n12776), .A(n12773), .ZN(n12775) );
  OR2_X1 U15904 ( .A1(n12774), .A2(n12776), .ZN(n12796) );
  INV_X1 U15905 ( .A(n12776), .ZN(n12777) );
  NAND2_X1 U15906 ( .A1(n12030), .A2(n12777), .ZN(n15269) );
  NOR2_X2 U15907 ( .A1(n15267), .A2(n9729), .ZN(n12802) );
  INV_X1 U15908 ( .A(n12802), .ZN(n12800) );
  AOI22_X1 U15909 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12785) );
  AOI22_X1 U15910 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12784) );
  NAND2_X1 U15911 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12782) );
  NAND2_X1 U15912 ( .A1(n9709), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12781) );
  NAND2_X1 U15913 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12780) );
  NAND2_X1 U15914 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12779) );
  AND4_X1 U15915 ( .A1(n12782), .A2(n12781), .A3(n12780), .A4(n12779), .ZN(
        n12783) );
  NAND4_X1 U15916 ( .A1(n12785), .A2(n12784), .A3(n12783), .A4(n12846), .ZN(
        n12794) );
  AOI22_X1 U15917 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12792) );
  AOI22_X1 U15918 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12791) );
  NAND2_X1 U15919 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12789) );
  NAND2_X1 U15920 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12788) );
  NAND2_X1 U15921 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12787) );
  NAND2_X1 U15922 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12786) );
  AND4_X1 U15923 ( .A1(n12789), .A2(n12788), .A3(n12787), .A4(n12786), .ZN(
        n12790) );
  NAND4_X1 U15924 ( .A1(n12792), .A2(n12852), .A3(n12791), .A4(n12790), .ZN(
        n12793) );
  NAND2_X1 U15925 ( .A1(n12794), .A2(n12793), .ZN(n12795) );
  INV_X1 U15926 ( .A(n12795), .ZN(n12804) );
  INV_X1 U15927 ( .A(n12796), .ZN(n12798) );
  OR2_X1 U15928 ( .A1(n12796), .A2(n12795), .ZN(n15248) );
  OAI211_X1 U15929 ( .C1(n12804), .C2(n12798), .A(n15248), .B(n12797), .ZN(
        n12801) );
  INV_X1 U15930 ( .A(n12801), .ZN(n12799) );
  NAND2_X1 U15931 ( .A1(n12802), .A2(n12801), .ZN(n12803) );
  NAND2_X1 U15932 ( .A1(n12030), .A2(n12804), .ZN(n15257) );
  AOI22_X1 U15933 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12812) );
  AOI22_X1 U15934 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12811) );
  NAND2_X1 U15935 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12809) );
  NAND2_X1 U15936 ( .A1(n9709), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12808) );
  NAND2_X1 U15937 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12807) );
  NAND2_X1 U15938 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12806) );
  AND4_X1 U15939 ( .A1(n12809), .A2(n12808), .A3(n12807), .A4(n12806), .ZN(
        n12810) );
  NAND4_X1 U15940 ( .A1(n12812), .A2(n12811), .A3(n12810), .A4(n12846), .ZN(
        n12821) );
  AOI22_X1 U15941 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12819) );
  AOI22_X1 U15942 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12818) );
  NAND2_X1 U15943 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12816) );
  NAND2_X1 U15944 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12815) );
  NAND2_X1 U15945 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12814) );
  NAND2_X1 U15946 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12813) );
  AND4_X1 U15947 ( .A1(n12816), .A2(n12815), .A3(n12814), .A4(n12813), .ZN(
        n12817) );
  NAND4_X1 U15948 ( .A1(n12819), .A2(n12852), .A3(n12818), .A4(n12817), .ZN(
        n12820) );
  AND2_X1 U15949 ( .A1(n12821), .A2(n12820), .ZN(n15249) );
  NAND2_X1 U15950 ( .A1(n10648), .A2(n15249), .ZN(n12822) );
  NOR2_X1 U15951 ( .A1(n15248), .A2(n12822), .ZN(n12841) );
  AOI22_X1 U15952 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12829) );
  AOI22_X1 U15953 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12828) );
  NAND2_X1 U15954 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12826) );
  NAND2_X1 U15955 ( .A1(n9708), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12825) );
  NAND2_X1 U15956 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12824) );
  NAND2_X1 U15957 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12823) );
  AND4_X1 U15958 ( .A1(n12826), .A2(n12825), .A3(n12824), .A4(n12823), .ZN(
        n12827) );
  NAND4_X1 U15959 ( .A1(n12829), .A2(n12828), .A3(n12827), .A4(n12846), .ZN(
        n12839) );
  AOI22_X1 U15960 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12837) );
  AOI22_X1 U15961 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12836) );
  NAND2_X1 U15962 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12834) );
  NAND2_X1 U15963 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12833) );
  NAND2_X1 U15964 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12832) );
  NAND2_X1 U15965 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12831) );
  AND4_X1 U15966 ( .A1(n12834), .A2(n12833), .A3(n12832), .A4(n12831), .ZN(
        n12835) );
  NAND4_X1 U15967 ( .A1(n12837), .A2(n12852), .A3(n12836), .A4(n12835), .ZN(
        n12838) );
  AND2_X1 U15968 ( .A1(n12839), .A2(n12838), .ZN(n12840) );
  NAND2_X1 U15969 ( .A1(n12841), .A2(n12840), .ZN(n12842) );
  OAI21_X1 U15970 ( .B1(n12841), .B2(n12840), .A(n12842), .ZN(n15244) );
  NOR2_X1 U15971 ( .A1(n15243), .A2(n15244), .ZN(n15242) );
  INV_X1 U15972 ( .A(n12842), .ZN(n12843) );
  NOR2_X1 U15973 ( .A1(n15242), .A2(n12843), .ZN(n12860) );
  AOI22_X1 U15974 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12845) );
  AOI22_X1 U15975 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12844) );
  NAND2_X1 U15976 ( .A1(n12845), .A2(n12844), .ZN(n12858) );
  AOI22_X1 U15977 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12830), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12848) );
  AOI22_X1 U15978 ( .A1(n9707), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12847) );
  NAND3_X1 U15979 ( .A1(n12848), .A2(n12847), .A3(n12846), .ZN(n12857) );
  AOI22_X1 U15980 ( .A1(n12716), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9712), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12851) );
  AOI22_X1 U15981 ( .A1(n12717), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12850) );
  NAND2_X1 U15982 ( .A1(n12851), .A2(n12850), .ZN(n12856) );
  AOI22_X1 U15983 ( .A1(n12805), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9709), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12854) );
  AOI22_X1 U15984 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12853) );
  NAND3_X1 U15985 ( .A1(n12854), .A2(n12853), .A3(n12852), .ZN(n12855) );
  OAI22_X1 U15986 ( .A1(n12858), .A2(n12857), .B1(n12856), .B2(n12855), .ZN(
        n12859) );
  XNOR2_X1 U15987 ( .A(n12860), .B(n12859), .ZN(n14536) );
  NAND2_X1 U15988 ( .A1(n16612), .A2(n16607), .ZN(n13347) );
  NAND2_X1 U15989 ( .A1(n13347), .A2(n12861), .ZN(n12862) );
  AND2_X1 U15990 ( .A1(n12494), .A2(n20202), .ZN(n13343) );
  NAND2_X1 U15991 ( .A1(n20198), .A2(n13343), .ZN(n12863) );
  INV_X1 U15992 ( .A(n13415), .ZN(n19584) );
  NAND2_X1 U15993 ( .A1(n19428), .A2(n12866), .ZN(n15369) );
  NOR4_X1 U15994 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12870) );
  NOR4_X1 U15995 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12869) );
  NOR4_X1 U15996 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12868) );
  NOR4_X1 U15997 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12867) );
  NAND4_X1 U15998 ( .A1(n12870), .A2(n12869), .A3(n12868), .A4(n12867), .ZN(
        n12875) );
  NOR4_X1 U15999 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12873) );
  NOR4_X1 U16000 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12872) );
  NOR4_X1 U16001 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12871) );
  NAND4_X1 U16002 ( .A1(n12873), .A2(n12872), .A3(n12871), .A4(n20093), .ZN(
        n12874) );
  INV_X1 U16003 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16737) );
  OR2_X1 U16004 ( .A1(n15293), .A2(n16737), .ZN(n12877) );
  NAND2_X1 U16005 ( .A1(n15293), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12876) );
  AND2_X1 U16006 ( .A1(n12877), .A2(n12876), .ZN(n19422) );
  INV_X1 U16007 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12878) );
  OAI22_X1 U16008 ( .A1(n15369), .A2(n19422), .B1(n19428), .B2(n12878), .ZN(
        n12879) );
  AOI21_X1 U16009 ( .B1(n19417), .B2(n12880), .A(n12879), .ZN(n12881) );
  INV_X1 U16010 ( .A(n12881), .ZN(n12885) );
  NAND3_X1 U16011 ( .A1(n19428), .A2(n12549), .A3(n13415), .ZN(n12882) );
  NOR2_X2 U16012 ( .A1(n12882), .A2(n13751), .ZN(n19418) );
  NOR2_X2 U16013 ( .A1(n12882), .A2(n13753), .ZN(n19419) );
  AOI22_X1 U16014 ( .A1(n19418), .A2(BUF2_REG_30__SCAN_IN), .B1(n19419), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n12883) );
  INV_X1 U16015 ( .A(n12883), .ZN(n12884) );
  OAI21_X1 U16016 ( .B1(n14536), .B2(n15373), .A(n12886), .ZN(P2_U2889) );
  INV_X1 U16017 ( .A(n12890), .ZN(n12893) );
  NOR2_X1 U16018 ( .A1(n12891), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12892) );
  MUX2_X1 U16019 ( .A(n12893), .B(n12892), .S(n9720), .Z(n16305) );
  NAND2_X1 U16020 ( .A1(n16305), .A2(n12162), .ZN(n12894) );
  XNOR2_X1 U16021 ( .A(n12894), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12895) );
  XNOR2_X1 U16022 ( .A(n12896), .B(n12895), .ZN(n14519) );
  AND2_X1 U16023 ( .A1(n10838), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12899) );
  INV_X1 U16024 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20135) );
  OAI22_X1 U16025 ( .A1(n10848), .A2(n20135), .B1(n15777), .B2(n10192), .ZN(
        n12898) );
  XNOR2_X1 U16026 ( .A(n12901), .B(n12900), .ZN(n16379) );
  NAND2_X1 U16027 ( .A1(n19517), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14507) );
  OAI21_X1 U16028 ( .B1(n16506), .B2(n10192), .A(n14507), .ZN(n12902) );
  AOI21_X1 U16029 ( .B1(n16379), .B2(n19512), .A(n12902), .ZN(n12903) );
  OAI21_X1 U16030 ( .B1(n12904), .B2(n19501), .A(n12903), .ZN(n12905) );
  NAND2_X1 U16031 ( .A1(n15383), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12906) );
  XNOR2_X2 U16032 ( .A(n12906), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14516) );
  NAND2_X1 U16033 ( .A1(n14516), .A2(n19507), .ZN(n12907) );
  OAI211_X1 U16034 ( .C1(n14519), .C2(n19510), .A(n12908), .B(n12907), .ZN(
        P2_U2983) );
  NAND2_X1 U16035 ( .A1(n16181), .A2(n14555), .ZN(n12909) );
  NAND2_X1 U16036 ( .A1(n16285), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14972) );
  OAI211_X1 U16037 ( .C1(n12910), .C2(n16187), .A(n12909), .B(n14972), .ZN(
        n12911) );
  AOI21_X1 U16038 ( .B1(n12912), .B2(n14887), .A(n12911), .ZN(n12918) );
  INV_X1 U16039 ( .A(n12913), .ZN(n12915) );
  NAND2_X1 U16040 ( .A1(n12915), .A2(n12914), .ZN(n12916) );
  XNOR2_X1 U16041 ( .A(n12916), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14980) );
  NAND2_X1 U16043 ( .A1(n12917), .A2(n12918), .ZN(P1_U2969) );
  INV_X1 U16044 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19135) );
  NOR2_X1 U16045 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n19135), .ZN(
        n16678) );
  NAND2_X1 U16046 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16647) );
  INV_X1 U16047 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16671) );
  NOR2_X1 U16048 ( .A1(n16647), .A2(n16671), .ZN(n15966) );
  INV_X1 U16049 ( .A(n15966), .ZN(n16016) );
  AOI22_X1 U16050 ( .A1(n15828), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12920) );
  OAI21_X1 U16051 ( .B1(n17429), .B2(n18740), .A(n12920), .ZN(n12936) );
  OR2_X2 U16052 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12922), .ZN(
        n12984) );
  NOR3_X2 U16053 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n12926), .ZN(n12952) );
  BUF_X4 U16054 ( .A(n12952), .Z(n17482) );
  AOI22_X1 U16055 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12934) );
  AOI22_X1 U16056 ( .A1(n17490), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12923) );
  OAI21_X1 U16057 ( .B1(n17470), .B2(n18528), .A(n12923), .ZN(n12932) );
  NOR3_X1 U16058 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n12924), .ZN(n12925) );
  INV_X1 U16059 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12930) );
  NOR3_X1 U16060 ( .A1(n19130), .A2(n19139), .A3(n17180), .ZN(n13017) );
  INV_X1 U16061 ( .A(n13017), .ZN(n12951) );
  INV_X1 U16062 ( .A(n12970), .ZN(n13141) );
  INV_X2 U16063 ( .A(n13141), .ZN(n17449) );
  AOI22_X1 U16064 ( .A1(n9685), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12929) );
  INV_X2 U16065 ( .A(n9755), .ZN(n15894) );
  AOI22_X1 U16066 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12928) );
  OAI211_X1 U16067 ( .C1(n12943), .C2(n12930), .A(n12929), .B(n12928), .ZN(
        n12931) );
  AOI211_X1 U16068 ( .C1(n17393), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n12932), .B(n12931), .ZN(n12933) );
  OAI211_X1 U16069 ( .C1(n12977), .C2(n17402), .A(n12934), .B(n12933), .ZN(
        n12935) );
  INV_X1 U16070 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12938) );
  AOI22_X1 U16071 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9704), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12937) );
  OAI21_X1 U16072 ( .B1(n17373), .B2(n12938), .A(n12937), .ZN(n12942) );
  AOI22_X1 U16073 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12940) );
  NAND3_X1 U16074 ( .A1(n12940), .A2(n10169), .A3(n12939), .ZN(n12941) );
  NOR2_X1 U16075 ( .A1(n12942), .A2(n12941), .ZN(n12950) );
  INV_X1 U16076 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18517) );
  AOI22_X1 U16077 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12944) );
  OAI21_X1 U16078 ( .B1(n17470), .B2(n18517), .A(n12944), .ZN(n12948) );
  INV_X1 U16079 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17300) );
  AOI22_X1 U16080 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13023), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12946) );
  AOI22_X1 U16081 ( .A1(n9685), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12945) );
  OAI211_X1 U16082 ( .C1(n15864), .C2(n17300), .A(n12946), .B(n12945), .ZN(
        n12947) );
  AOI211_X1 U16083 ( .C1(n17393), .C2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n12948), .B(n12947), .ZN(n12949) );
  INV_X1 U16084 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17337) );
  AOI22_X1 U16085 ( .A1(n17430), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12952), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12953) );
  OAI21_X1 U16086 ( .B1(n12951), .B2(n17337), .A(n12953), .ZN(n12955) );
  INV_X1 U16087 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15841) );
  AOI22_X1 U16088 ( .A1(n17490), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12957) );
  OAI21_X1 U16089 ( .B1(n17485), .B2(n15841), .A(n12957), .ZN(n12958) );
  INV_X1 U16090 ( .A(n12958), .ZN(n12967) );
  AOI22_X1 U16091 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12961) );
  INV_X1 U16092 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18506) );
  AOI22_X1 U16093 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12970), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12964) );
  AOI22_X1 U16094 ( .A1(n12962), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13023), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12963) );
  OAI211_X1 U16095 ( .C1(n17470), .C2(n18506), .A(n12964), .B(n12963), .ZN(
        n12965) );
  INV_X1 U16096 ( .A(n12965), .ZN(n12966) );
  NAND3_X1 U16097 ( .A1(n12967), .A2(n9769), .A3(n12966), .ZN(n12968) );
  AOI22_X1 U16098 ( .A1(n12970), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17430), .ZN(n12972) );
  AOI22_X1 U16099 ( .A1(n13017), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n13023), .ZN(n12971) );
  OAI211_X1 U16100 ( .C1(n18501), .C2(n17470), .A(n12972), .B(n12971), .ZN(
        n12976) );
  AOI22_X1 U16101 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n17465), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n12952), .ZN(n12974) );
  INV_X1 U16102 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17344) );
  NAND3_X1 U16103 ( .A1(n12974), .A2(n12973), .A3(n10168), .ZN(n12975) );
  NOR2_X1 U16104 ( .A1(n12976), .A2(n12975), .ZN(n12983) );
  AOI22_X1 U16105 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n17448), .ZN(n12981) );
  AOI22_X1 U16106 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17467), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12980) );
  AOI22_X1 U16107 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17489), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12979) );
  NAND2_X1 U16108 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17288), .ZN(
        n12978) );
  AOI22_X1 U16109 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12992) );
  AOI22_X1 U16110 ( .A1(n17431), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12970), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12991) );
  AOI22_X1 U16111 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12990) );
  INV_X1 U16112 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18512) );
  INV_X1 U16113 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17428) );
  OAI22_X1 U16114 ( .A1(n17470), .A2(n18512), .B1(n12943), .B2(n17428), .ZN(
        n12989) );
  AOI22_X1 U16115 ( .A1(n9685), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9704), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12988) );
  AOI22_X1 U16116 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12987) );
  AOI22_X1 U16117 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13023), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12986) );
  NAND2_X1 U16118 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12985) );
  AOI22_X1 U16119 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13002) );
  INV_X1 U16120 ( .A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13124) );
  AOI22_X1 U16121 ( .A1(n12970), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12994) );
  AOI22_X1 U16122 ( .A1(n17430), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12993) );
  OAI211_X1 U16123 ( .C1(n12943), .C2(n13124), .A(n12994), .B(n12993), .ZN(
        n13000) );
  AOI22_X1 U16124 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17431), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12998) );
  AOI22_X1 U16125 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12997) );
  AOI22_X1 U16126 ( .A1(n9685), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9704), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12996) );
  NAND2_X1 U16127 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12995) );
  NAND4_X1 U16128 ( .A1(n12998), .A2(n12997), .A3(n12996), .A4(n12995), .ZN(
        n12999) );
  AOI211_X1 U16129 ( .C1(n17490), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n13000), .B(n12999), .ZN(n13001) );
  INV_X1 U16130 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13013) );
  AOI22_X1 U16131 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13012) );
  AOI22_X1 U16132 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13004) );
  AOI22_X1 U16133 ( .A1(n17431), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13003) );
  OAI211_X1 U16134 ( .C1(n17470), .C2(n18537), .A(n13004), .B(n13003), .ZN(
        n13010) );
  AOI22_X1 U16135 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13008) );
  AOI22_X1 U16136 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9685), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13007) );
  AOI22_X1 U16137 ( .A1(n15828), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13006) );
  NAND2_X1 U16138 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n13005) );
  NAND4_X1 U16139 ( .A1(n13008), .A2(n13007), .A3(n13006), .A4(n13005), .ZN(
        n13009) );
  OAI211_X1 U16140 ( .C1(n12943), .C2(n13013), .A(n13012), .B(n13011), .ZN(
        n16687) );
  INV_X1 U16141 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18180) );
  INV_X1 U16142 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18248) );
  NAND2_X1 U16143 ( .A1(n17927), .A2(n18248), .ZN(n13014) );
  INV_X1 U16144 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18220) );
  NAND2_X1 U16145 ( .A1(n17886), .A2(n18220), .ZN(n17870) );
  NAND2_X1 U16146 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18350) );
  NOR2_X1 U16147 ( .A1(n18350), .A2(n18021), .ZN(n18335) );
  NAND3_X1 U16148 ( .A1(n18335), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17956) );
  AND2_X1 U16149 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13037), .ZN(
        n13038) );
  AOI22_X1 U16150 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13030) );
  INV_X1 U16151 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18496) );
  INV_X1 U16152 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17357) );
  OAI22_X1 U16153 ( .A1(n17470), .A2(n18496), .B1(n12943), .B2(n17357), .ZN(
        n13020) );
  AOI22_X1 U16154 ( .A1(n13017), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13018) );
  INV_X1 U16155 ( .A(n13018), .ZN(n13019) );
  AOI22_X1 U16156 ( .A1(n17431), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13021) );
  AOI22_X1 U16157 ( .A1(n12970), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13027) );
  AOI22_X1 U16158 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9688), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13026) );
  AOI22_X1 U16159 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13023), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13025) );
  NAND2_X1 U16160 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13024) );
  NAND4_X2 U16161 ( .A1(n13030), .A2(n13029), .A3(n13028), .A4(n9757), .ZN(
        n18146) );
  NAND2_X1 U16162 ( .A1(n18146), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18145) );
  NOR2_X1 U16163 ( .A1(n17682), .A2(n13031), .ZN(n13032) );
  NOR2_X1 U16164 ( .A1(n18443), .A2(n13033), .ZN(n13034) );
  INV_X1 U16165 ( .A(n13190), .ZN(n17670) );
  XOR2_X1 U16166 ( .A(n17670), .B(n13035), .Z(n18112) );
  NOR2_X1 U16167 ( .A1(n18111), .A2(n18112), .ZN(n13036) );
  NAND2_X1 U16168 ( .A1(n18111), .A2(n18112), .ZN(n18110) );
  OAI21_X1 U16169 ( .B1(n13036), .B2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n18110), .ZN(n18103) );
  XNOR2_X1 U16170 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n13037), .ZN(
        n18104) );
  NOR2_X1 U16171 ( .A1(n18103), .A2(n18104), .ZN(n18102) );
  NOR2_X2 U16172 ( .A1(n13038), .A2(n18102), .ZN(n18088) );
  INV_X1 U16173 ( .A(n13188), .ZN(n17663) );
  XOR2_X1 U16174 ( .A(n17663), .B(n13039), .Z(n18089) );
  XOR2_X1 U16175 ( .A(n17660), .B(n13041), .Z(n13042) );
  XNOR2_X1 U16176 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n13042), .ZN(
        n18073) );
  OAI21_X1 U16177 ( .B1(n13043), .B2(n16687), .A(n17968), .ZN(n13044) );
  NOR2_X1 U16178 ( .A1(n13045), .A2(n13044), .ZN(n13046) );
  XNOR2_X1 U16179 ( .A(n13045), .B(n13044), .ZN(n18068) );
  INV_X1 U16180 ( .A(n18396), .ZN(n18056) );
  NOR2_X1 U16181 ( .A1(n18285), .A2(n18269), .ZN(n18261) );
  INV_X1 U16182 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17921) );
  NAND2_X1 U16183 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18221) );
  NOR3_X1 U16184 ( .A1(n17921), .A2(n18220), .A3(n18221), .ZN(n13053) );
  NAND2_X1 U16185 ( .A1(n18261), .A2(n13053), .ZN(n18158) );
  INV_X1 U16186 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18157) );
  NOR2_X1 U16187 ( .A1(n18158), .A2(n18157), .ZN(n16644) );
  NAND2_X1 U16188 ( .A1(n16644), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17855) );
  INV_X1 U16189 ( .A(n17855), .ZN(n13052) );
  NOR2_X1 U16190 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n13049) );
  NOR2_X2 U16191 ( .A1(n18033), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18022) );
  INV_X1 U16192 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18363) );
  INV_X1 U16193 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17981) );
  NOR2_X1 U16194 ( .A1(n17941), .A2(n13051), .ZN(n17937) );
  NAND2_X1 U16195 ( .A1(n17937), .A2(n18269), .ZN(n17936) );
  AND2_X1 U16196 ( .A1(n13053), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18196) );
  NAND2_X1 U16197 ( .A1(n18261), .A2(n17868), .ZN(n17884) );
  INV_X1 U16198 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18197) );
  NOR2_X1 U16199 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17824), .ZN(
        n17823) );
  NOR2_X1 U16200 ( .A1(n17842), .A2(n17968), .ZN(n13054) );
  NAND2_X1 U16201 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15963) );
  NOR2_X1 U16202 ( .A1(n17823), .A2(n13055), .ZN(n13056) );
  INV_X1 U16203 ( .A(n10069), .ZN(n13057) );
  NOR2_X2 U16204 ( .A1(n13056), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16686) );
  INV_X1 U16205 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17803) );
  NAND2_X1 U16206 ( .A1(n16686), .A2(n17803), .ZN(n15970) );
  AOI22_X1 U16207 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18057), .B1(
        n17968), .B2(n19135), .ZN(n13060) );
  INV_X1 U16208 ( .A(n13058), .ZN(n13061) );
  INV_X1 U16209 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16655) );
  OAI21_X1 U16210 ( .B1(n13061), .B2(n16014), .A(n13060), .ZN(n13062) );
  NAND2_X1 U16211 ( .A1(n13063), .A2(n13062), .ZN(n16682) );
  OAI21_X1 U16212 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18487), .A(
        n13182), .ZN(n13181) );
  NOR2_X1 U16213 ( .A1(n13181), .A2(n13185), .ZN(n13077) );
  NOR2_X1 U16214 ( .A1(n13185), .A2(n13182), .ZN(n13064) );
  OAI22_X1 U16215 ( .A1(n19139), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n19001), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13068) );
  NOR2_X1 U16216 ( .A1(n13069), .A2(n13068), .ZN(n13065) );
  AOI22_X1 U16217 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18963), .B1(
        n13066), .B2(n19130), .ZN(n13070) );
  NOR2_X1 U16218 ( .A1(n13066), .A2(n19130), .ZN(n13071) );
  NAND2_X1 U16219 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18963), .ZN(
        n13067) );
  OAI22_X1 U16220 ( .A1(n13070), .A2(n19004), .B1(n13071), .B2(n13067), .ZN(
        n13074) );
  INV_X1 U16221 ( .A(n13074), .ZN(n13076) );
  XNOR2_X1 U16222 ( .A(n13069), .B(n13068), .ZN(n13075) );
  INV_X1 U16223 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19005) );
  OAI21_X1 U16224 ( .B1(n19004), .B2(n13071), .A(n13070), .ZN(n13072) );
  INV_X1 U16225 ( .A(n13072), .ZN(n13073) );
  AOI22_X1 U16226 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17431), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13078) );
  OAI21_X1 U16227 ( .B1(n12951), .B2(n18806), .A(n13078), .ZN(n13087) );
  AOI22_X1 U16228 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9704), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13085) );
  OAI22_X1 U16229 ( .A1(n9682), .A2(n17471), .B1(n17485), .B2(n17464), .ZN(
        n13083) );
  AOI22_X1 U16230 ( .A1(n15828), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13081) );
  AOI22_X1 U16231 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13080) );
  NAND3_X1 U16232 ( .A1(n13081), .A2(n13080), .A3(n13079), .ZN(n13082) );
  AOI211_X1 U16233 ( .C1(n17393), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n13083), .B(n13082), .ZN(n13084) );
  OAI211_X1 U16234 ( .C1(n13141), .C2(n18501), .A(n13085), .B(n13084), .ZN(
        n13086) );
  AOI22_X1 U16235 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13089) );
  AOI22_X1 U16236 ( .A1(n17467), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13088) );
  OAI211_X1 U16237 ( .C1(n12943), .C2(n18722), .A(n13089), .B(n13088), .ZN(
        n13097) );
  AOI22_X1 U16238 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13095) );
  AOI22_X1 U16239 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13090) );
  OAI21_X1 U16240 ( .B1(n12951), .B2(n18802), .A(n13090), .ZN(n13093) );
  INV_X1 U16241 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18900) );
  AOI22_X1 U16242 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13091) );
  OAI21_X1 U16243 ( .B1(n17470), .B2(n18900), .A(n13091), .ZN(n13092) );
  AOI211_X1 U16244 ( .C1(n15895), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n13093), .B(n13092), .ZN(n13094) );
  OAI211_X1 U16245 ( .C1(n12959), .C2(n17357), .A(n13095), .B(n13094), .ZN(
        n13096) );
  NOR2_X1 U16246 ( .A1(n19171), .A2(n18493), .ZN(n13160) );
  OR2_X1 U16247 ( .A1(n13162), .A2(n13160), .ZN(n19185) );
  AOI22_X1 U16248 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13098) );
  OAI21_X1 U16249 ( .B1(n12951), .B2(n18825), .A(n13098), .ZN(n13107) );
  AOI22_X1 U16250 ( .A1(n15828), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13105) );
  INV_X1 U16251 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17223) );
  INV_X1 U16252 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17374) );
  OAI22_X1 U16253 ( .A1(n17485), .A2(n17223), .B1(n17470), .B2(n17374), .ZN(
        n13103) );
  AOI22_X1 U16254 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13101) );
  AOI22_X1 U16255 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13100) );
  AOI22_X1 U16256 ( .A1(n17490), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13099) );
  NAND3_X1 U16257 ( .A1(n13101), .A2(n13100), .A3(n13099), .ZN(n13102) );
  AOI211_X1 U16258 ( .C1(n17393), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n13103), .B(n13102), .ZN(n13104) );
  OAI211_X1 U16259 ( .C1(n12984), .C2(n17372), .A(n13105), .B(n13104), .ZN(
        n13106) );
  AOI211_X4 U16260 ( .C1(n17431), .C2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n13107), .B(n13106), .ZN(n18533) );
  AOI22_X1 U16261 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9704), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13108) );
  OAI21_X1 U16262 ( .B1(n12919), .B2(n17316), .A(n13108), .ZN(n13117) );
  INV_X1 U16263 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18812) );
  AOI22_X1 U16264 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13115) );
  INV_X1 U16265 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18919) );
  AOI22_X1 U16266 ( .A1(n17490), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13109) );
  OAI21_X1 U16267 ( .B1(n17470), .B2(n18919), .A(n13109), .ZN(n13113) );
  INV_X1 U16268 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17315) );
  AOI22_X1 U16269 ( .A1(n17467), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13111) );
  AOI22_X1 U16270 ( .A1(n12970), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13110) );
  OAI211_X1 U16271 ( .C1(n12943), .C2(n17315), .A(n13111), .B(n13110), .ZN(
        n13112) );
  AOI211_X1 U16272 ( .C1(n17393), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n13113), .B(n13112), .ZN(n13114) );
  OAI211_X1 U16273 ( .C1(n12951), .C2(n18812), .A(n13115), .B(n13114), .ZN(
        n13116) );
  AOI22_X1 U16274 ( .A1(n17430), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13118) );
  OAI21_X1 U16275 ( .B1(n13141), .B2(n18523), .A(n13118), .ZN(n13126) );
  AOI22_X1 U16276 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13123) );
  INV_X1 U16277 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18736) );
  AOI22_X1 U16278 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13119) );
  OAI21_X1 U16279 ( .B1(n12943), .B2(n18736), .A(n13119), .ZN(n13121) );
  INV_X1 U16280 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18933) );
  AOI22_X1 U16281 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17431), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13120) );
  OAI211_X1 U16282 ( .C1(n12959), .C2(n13124), .A(n13123), .B(n13122), .ZN(
        n13125) );
  AOI22_X1 U16283 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13136) );
  AOI22_X1 U16284 ( .A1(n9685), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13128) );
  AOI22_X1 U16285 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17467), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13127) );
  OAI211_X1 U16286 ( .C1(n15864), .C2(n17452), .A(n13128), .B(n13127), .ZN(
        n13134) );
  AOI22_X1 U16287 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13132) );
  AOI22_X1 U16288 ( .A1(n17430), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13131) );
  AOI22_X1 U16289 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17488), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13130) );
  NAND2_X1 U16290 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n13129) );
  NAND4_X1 U16291 ( .A1(n13132), .A2(n13131), .A3(n13130), .A4(n13129), .ZN(
        n13133) );
  AOI211_X1 U16292 ( .C1(n17393), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n13134), .B(n13133), .ZN(n13135) );
  OAI211_X1 U16293 ( .C1(n9756), .C2(n13137), .A(n13136), .B(n13135), .ZN(
        n15948) );
  NOR2_X1 U16294 ( .A1(n18520), .A2(n15948), .ZN(n15952) );
  AOI22_X1 U16295 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13139) );
  AOI22_X1 U16296 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17467), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13138) );
  OAI211_X1 U16297 ( .C1(n12943), .C2(n18733), .A(n13139), .B(n13138), .ZN(
        n13148) );
  INV_X1 U16298 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15833) );
  AOI22_X1 U16299 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13146) );
  AOI22_X1 U16300 ( .A1(n17430), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13140) );
  OAI21_X1 U16301 ( .B1(n13141), .B2(n18517), .A(n13140), .ZN(n13144) );
  INV_X1 U16302 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17413) );
  AOI22_X1 U16303 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13142) );
  OAI21_X1 U16304 ( .B1(n9681), .B2(n17413), .A(n13142), .ZN(n13143) );
  AOI211_X1 U16305 ( .C1(n9685), .C2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A(
        n13144), .B(n13143), .ZN(n13145) );
  OAI211_X1 U16306 ( .C1(n17485), .C2(n15833), .A(n13146), .B(n13145), .ZN(
        n13147) );
  AOI22_X1 U16307 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13158) );
  AOI22_X1 U16308 ( .A1(n17431), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13150) );
  AOI22_X1 U16309 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9704), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13149) );
  OAI211_X1 U16310 ( .C1(n12943), .C2(n18740), .A(n13150), .B(n13149), .ZN(
        n13156) );
  AOI22_X1 U16311 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9685), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13154) );
  AOI22_X1 U16312 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13153) );
  AOI22_X1 U16313 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17488), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13152) );
  NAND2_X1 U16314 ( .A1(n17490), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n13151) );
  NAND4_X1 U16315 ( .A1(n13154), .A2(n13153), .A3(n13152), .A4(n13151), .ZN(
        n13155) );
  AOI211_X1 U16316 ( .C1(n17393), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n13156), .B(n13155), .ZN(n13157) );
  NOR2_X1 U16317 ( .A1(n18514), .A2(n13174), .ZN(n18968) );
  NAND3_X1 U16318 ( .A1(n13175), .A2(n15952), .A3(n18968), .ZN(n15943) );
  INV_X1 U16319 ( .A(n18509), .ZN(n13170) );
  NOR2_X1 U16320 ( .A1(n18525), .A2(n17538), .ZN(n13177) );
  NAND2_X1 U16321 ( .A1(n18967), .A2(n13177), .ZN(n15908) );
  NOR2_X1 U16322 ( .A1(n19171), .A2(n15908), .ZN(n13159) );
  INV_X1 U16323 ( .A(n18514), .ZN(n13178) );
  NOR2_X1 U16324 ( .A1(n13174), .A2(n13178), .ZN(n13165) );
  NAND4_X1 U16325 ( .A1(n13175), .A2(n18520), .A3(n13161), .A4(n17689), .ZN(
        n15933) );
  AND4_X1 U16326 ( .A1(n18509), .A2(n18514), .A3(n13168), .A4(n13166), .ZN(
        n13171) );
  NAND2_X1 U16327 ( .A1(n17578), .A2(n18989), .ZN(n16037) );
  NAND2_X1 U16328 ( .A1(n13160), .A2(n16037), .ZN(n15938) );
  OAI21_X1 U16329 ( .B1(n15952), .B2(n13161), .A(n15938), .ZN(n13169) );
  NAND2_X1 U16330 ( .A1(n17578), .A2(n15947), .ZN(n13163) );
  OAI21_X1 U16331 ( .B1(n15948), .B2(n17689), .A(n18989), .ZN(n13164) );
  OAI21_X1 U16332 ( .B1(n13166), .B2(n13165), .A(n13164), .ZN(n13167) );
  AOI21_X1 U16333 ( .B1(n13170), .B2(n13169), .A(n15936), .ZN(n13172) );
  OR3_X1 U16334 ( .A1(n18498), .A2(n13251), .A3(n13175), .ZN(n13173) );
  NAND2_X1 U16335 ( .A1(n13173), .A2(n13172), .ZN(n18966) );
  NOR2_X1 U16336 ( .A1(n18498), .A2(n15948), .ZN(n15950) );
  NAND2_X1 U16337 ( .A1(n15950), .A2(n13174), .ZN(n15956) );
  INV_X1 U16338 ( .A(n13175), .ZN(n13176) );
  AOI211_X1 U16339 ( .C1(n13178), .C2(n18989), .A(n13177), .B(n13176), .ZN(
        n13179) );
  NAND2_X1 U16340 ( .A1(n13180), .A2(n13179), .ZN(n15937) );
  INV_X1 U16341 ( .A(n13181), .ZN(n13187) );
  INV_X1 U16342 ( .A(n13182), .ZN(n13186) );
  NAND2_X1 U16343 ( .A1(n13186), .A2(n13185), .ZN(n13183) );
  OAI211_X1 U16344 ( .C1(n13186), .C2(n13185), .A(n13184), .B(n13183), .ZN(
        n13252) );
  OAI21_X1 U16345 ( .B1(n13187), .B2(n13252), .A(n13253), .ZN(n18958) );
  INV_X1 U16346 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19134) );
  NAND2_X1 U16347 ( .A1(n19134), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n19025) );
  NAND2_X1 U16348 ( .A1(n16682), .A2(n18058), .ZN(n13229) );
  NAND2_X1 U16349 ( .A1(n18146), .A2(n17682), .ZN(n13192) );
  NAND2_X1 U16350 ( .A1(n17675), .A2(n13192), .ZN(n13191) );
  NAND2_X1 U16351 ( .A1(n13191), .A2(n13190), .ZN(n13201) );
  NAND2_X1 U16352 ( .A1(n13189), .A2(n13188), .ZN(n13207) );
  NOR2_X1 U16353 ( .A1(n17660), .A2(n13207), .ZN(n13211) );
  NAND2_X1 U16354 ( .A1(n13211), .A2(n16687), .ZN(n13212) );
  XOR2_X1 U16355 ( .A(n13189), .B(n13188), .Z(n13205) );
  AND2_X1 U16356 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13205), .ZN(
        n13206) );
  XNOR2_X1 U16357 ( .A(n13191), .B(n13190), .ZN(n13199) );
  INV_X1 U16358 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18427) );
  NOR2_X1 U16359 ( .A1(n13199), .A2(n18427), .ZN(n13200) );
  XOR2_X1 U16360 ( .A(n17675), .B(n13192), .Z(n13193) );
  NOR2_X1 U16361 ( .A1(n13193), .A2(n18443), .ZN(n13198) );
  XNOR2_X1 U16362 ( .A(n18443), .B(n13193), .ZN(n18126) );
  INV_X1 U16363 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19149) );
  NOR2_X1 U16364 ( .A1(n13195), .A2(n19149), .ZN(n13197) );
  INV_X1 U16365 ( .A(n18146), .ZN(n13196) );
  NAND3_X1 U16366 ( .A1(n13196), .A2(n13195), .A3(n19149), .ZN(n13194) );
  OAI221_X1 U16367 ( .B1(n13197), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n13196), .C2(n13195), .A(n13194), .ZN(n18125) );
  NOR2_X1 U16368 ( .A1(n18126), .A2(n18125), .ZN(n18124) );
  NOR2_X1 U16369 ( .A1(n13198), .A2(n18124), .ZN(n18116) );
  XNOR2_X1 U16370 ( .A(n13199), .B(n18427), .ZN(n18115) );
  NOR2_X1 U16371 ( .A1(n18116), .A2(n18115), .ZN(n18114) );
  NOR2_X1 U16372 ( .A1(n13200), .A2(n18114), .ZN(n13202) );
  XNOR2_X1 U16373 ( .A(n13201), .B(n17667), .ZN(n13203) );
  NOR2_X1 U16374 ( .A1(n13202), .A2(n13203), .ZN(n13204) );
  INV_X1 U16375 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18432) );
  XNOR2_X1 U16376 ( .A(n13203), .B(n13202), .ZN(n18099) );
  NOR2_X1 U16377 ( .A1(n18432), .A2(n18099), .ZN(n18098) );
  NOR2_X1 U16378 ( .A1(n13204), .A2(n18098), .ZN(n18093) );
  XNOR2_X1 U16379 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n13205), .ZN(
        n18092) );
  NOR2_X1 U16380 ( .A1(n18093), .A2(n18092), .ZN(n18091) );
  XNOR2_X1 U16381 ( .A(n13207), .B(n17660), .ZN(n13209) );
  NOR2_X1 U16382 ( .A1(n13208), .A2(n13209), .ZN(n13210) );
  XNOR2_X1 U16383 ( .A(n13209), .B(n13208), .ZN(n18076) );
  INV_X1 U16384 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18399) );
  NOR2_X1 U16385 ( .A1(n13210), .A2(n18075), .ZN(n13213) );
  XOR2_X1 U16386 ( .A(n13211), .B(n17656), .Z(n13214) );
  NAND2_X1 U16387 ( .A1(n13213), .A2(n13214), .ZN(n18061) );
  NAND2_X1 U16388 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18061), .ZN(
        n13216) );
  NOR2_X1 U16389 ( .A1(n13212), .A2(n13216), .ZN(n13218) );
  INV_X1 U16390 ( .A(n13212), .ZN(n13217) );
  OR2_X1 U16391 ( .A1(n13214), .A2(n13213), .ZN(n18062) );
  OAI21_X1 U16392 ( .B1(n13217), .B2(n13216), .A(n18062), .ZN(n13215) );
  AOI21_X1 U16393 ( .B1(n13217), .B2(n13216), .A(n13215), .ZN(n18054) );
  NOR2_X2 U16394 ( .A1(n13218), .A2(n18053), .ZN(n18345) );
  NOR2_X2 U16395 ( .A1(n18345), .A2(n15959), .ZN(n18287) );
  INV_X1 U16396 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18200) );
  NOR2_X1 U16397 ( .A1(n17855), .A2(n18200), .ZN(n18179) );
  NAND2_X1 U16398 ( .A1(n18287), .A2(n18179), .ZN(n17840) );
  NAND3_X1 U16399 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15966), .A3(
        n18155), .ZN(n13219) );
  XOR2_X1 U16400 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13219), .Z(
        n16685) );
  NOR2_X1 U16401 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19184) );
  INV_X1 U16402 ( .A(n19184), .ZN(n17197) );
  INV_X1 U16403 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19125) );
  NAND2_X1 U16404 ( .A1(n19183), .A2(n19125), .ZN(n16810) );
  NAND2_X1 U16405 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18105) );
  NAND2_X1 U16406 ( .A1(n18011), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18047) );
  NOR2_X1 U16407 ( .A1(n18065), .A2(n18049), .ZN(n18045) );
  NAND4_X1 U16408 ( .A1(n18045), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16842) );
  INV_X1 U16409 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18000) );
  NAND2_X1 U16410 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17947) );
  NAND2_X1 U16411 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17913) );
  NAND2_X1 U16412 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17878) );
  NAND2_X1 U16413 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17837) );
  NAND2_X1 U16414 ( .A1(n17825), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13220) );
  NAND2_X1 U16415 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17797) );
  INV_X1 U16416 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19106) );
  INV_X1 U16417 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19174) );
  NAND3_X2 U16418 ( .A1(n19184), .A2(n19174), .A3(n19183), .ZN(n18375) );
  NOR2_X1 U16419 ( .A1(n19106), .A2(n18375), .ZN(n16677) );
  NOR3_X1 U16420 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n16812), .ZN(n15932) );
  OAI21_X1 U16421 ( .B1(n18143), .B2(n17899), .A(n18717), .ZN(n17983) );
  NAND2_X1 U16422 ( .A1(n9828), .A2(n17983), .ZN(n16650) );
  XOR2_X1 U16423 ( .A(n9929), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(n13222) );
  NOR2_X1 U16424 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17899), .ZN(
        n16663) );
  INV_X1 U16425 ( .A(n13220), .ZN(n17796) );
  NAND2_X1 U16426 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17796), .ZN(
        n16832) );
  OR2_X1 U16427 ( .A1(n16832), .A2(n17797), .ZN(n16830) );
  NOR2_X1 U16428 ( .A1(n18717), .A2(n9828), .ZN(n16659) );
  AOI211_X1 U16429 ( .C1(n16830), .C2(n17987), .A(n18118), .B(n16659), .ZN(
        n13221) );
  INV_X1 U16430 ( .A(n13221), .ZN(n16661) );
  NOR2_X1 U16431 ( .A1(n16663), .A2(n16661), .ZN(n16649) );
  OAI22_X1 U16432 ( .A1(n16650), .A2(n13222), .B1(n16649), .B2(n9929), .ZN(
        n13223) );
  AOI211_X1 U16433 ( .C1(n18004), .C2(n9924), .A(n16677), .B(n13223), .ZN(
        n13227) );
  INV_X1 U16434 ( .A(n15963), .ZN(n18162) );
  INV_X1 U16435 ( .A(n18179), .ZN(n15962) );
  NAND2_X1 U16436 ( .A1(n18256), .A2(n13224), .ZN(n17872) );
  NAND2_X1 U16437 ( .A1(n18162), .A2(n17834), .ZN(n18165) );
  NAND3_X1 U16438 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15966), .A3(
        n19135), .ZN(n16674) );
  NAND2_X1 U16439 ( .A1(n15966), .A2(n17802), .ZN(n16657) );
  OAI21_X1 U16440 ( .B1(n16655), .B2(n16657), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13225) );
  OAI21_X1 U16441 ( .B1(n18165), .B2(n16674), .A(n13225), .ZN(n16679) );
  NAND2_X1 U16442 ( .A1(n16679), .A2(n18008), .ZN(n13226) );
  NAND2_X1 U16443 ( .A1(n13229), .A2(n10188), .ZN(P3_U2799) );
  NOR2_X1 U16444 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13231) );
  NOR4_X1 U16445 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13230) );
  NAND4_X1 U16446 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13231), .A4(n13230), .ZN(n13234) );
  INV_X1 U16447 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n20967) );
  INV_X1 U16448 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20994) );
  NOR4_X1 U16449 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), .A3(
        n20967), .A4(n20994), .ZN(n13233) );
  NOR4_X1 U16450 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n13232)
         );
  NAND3_X1 U16451 ( .A1(n13800), .A2(n13233), .A3(n13232), .ZN(U214) );
  NOR2_X1 U16452 ( .A1(n13753), .A2(n13234), .ZN(n16705) );
  NAND2_X1 U16453 ( .A1(n16705), .A2(U214), .ZN(U212) );
  NAND2_X1 U16454 ( .A1(n19342), .A2(n13243), .ZN(n19397) );
  AOI211_X1 U16455 ( .C1(n16463), .C2(n13235), .A(n19313), .B(n19397), .ZN(
        n13249) );
  INV_X1 U16456 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13924) );
  AOI22_X1 U16457 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19360), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n19366), .ZN(n13236) );
  OAI211_X1 U16458 ( .C1(n13924), .C2(n19382), .A(n13236), .B(n19324), .ZN(
        n13248) );
  NAND2_X1 U16459 ( .A1(n13237), .A2(n13446), .ZN(n13240) );
  INV_X1 U16460 ( .A(n13238), .ZN(n13239) );
  NAND2_X1 U16461 ( .A1(n13240), .A2(n13239), .ZN(n19431) );
  OAI22_X1 U16462 ( .A1(n13241), .A2(n19362), .B1(n19381), .B2(n19431), .ZN(
        n13247) );
  AOI21_X1 U16463 ( .B1(n13242), .B2(n15735), .A(n14010), .ZN(n16549) );
  INV_X1 U16464 ( .A(n16549), .ZN(n13245) );
  NAND2_X1 U16465 ( .A1(n19372), .A2(n19342), .ZN(n19390) );
  INV_X1 U16466 ( .A(n16463), .ZN(n13244) );
  OAI22_X1 U16467 ( .A1(n13245), .A2(n19354), .B1(n19390), .B2(n13244), .ZN(
        n13246) );
  INV_X1 U16468 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17532) );
  INV_X1 U16469 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17526) );
  NAND2_X1 U16470 ( .A1(n17532), .A2(n17526), .ZN(n13255) );
  NOR3_X1 U16471 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17175) );
  NAND2_X1 U16472 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n19165) );
  NAND2_X1 U16473 ( .A1(n13253), .A2(n13252), .ZN(n18955) );
  NAND2_X1 U16474 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n19171), .ZN(n13254) );
  AOI211_X4 U16475 ( .C1(n16812), .C2(n19165), .A(n13256), .B(n13254), .ZN(
        n17193) );
  AOI211_X1 U16476 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n13255), .A(n17175), .B(
        n17192), .ZN(n13265) );
  INV_X1 U16477 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19153) );
  INV_X1 U16478 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19049) );
  NOR2_X1 U16479 ( .A1(n19153), .A2(n19049), .ZN(n17167) );
  NAND2_X2 U16480 ( .A1(n19116), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19109) );
  OAI211_X1 U16481 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n19045), .B(n19109), .ZN(n19038) );
  INV_X1 U16482 ( .A(n19038), .ZN(n19170) );
  AOI211_X1 U16483 ( .C1(n19153), .C2(n19049), .A(n17167), .B(n17187), .ZN(
        n13264) );
  INV_X1 U16484 ( .A(n19186), .ZN(n13259) );
  NAND3_X1 U16485 ( .A1(n19174), .A2(n19183), .A3(n16812), .ZN(n19030) );
  NOR2_X2 U16486 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19125), .ZN(n19023) );
  INV_X1 U16487 ( .A(n19023), .ZN(n18893) );
  OR2_X1 U16488 ( .A1(n19025), .A2(n18893), .ZN(n19018) );
  INV_X1 U16489 ( .A(n19013), .ZN(n13257) );
  AOI211_X1 U16490 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n19171), .A(n13257), .B(
        n13256), .ZN(n13258) );
  INV_X1 U16491 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17519) );
  OAI22_X1 U16492 ( .A1(n18133), .A2(n17159), .B1(n17136), .B2(n17519), .ZN(
        n13263) );
  NOR2_X1 U16493 ( .A1(n9924), .A2(n19028), .ZN(n17125) );
  INV_X1 U16494 ( .A(n17125), .ZN(n16979) );
  AOI22_X1 U16495 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18133), .B1(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18143), .ZN(n18129) );
  INV_X1 U16496 ( .A(n17196), .ZN(n17181) );
  AOI21_X1 U16497 ( .B1(n18974), .B2(n19139), .A(n18970), .ZN(n19136) );
  NOR2_X1 U16498 ( .A1(n17689), .A2(n13259), .ZN(n19188) );
  AOI22_X1 U16499 ( .A1(n17181), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n19136), 
        .B2(n19188), .ZN(n13261) );
  INV_X1 U16500 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17110) );
  NAND2_X1 U16501 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17110), .ZN(
        n17150) );
  INV_X1 U16502 ( .A(n17150), .ZN(n16989) );
  AOI21_X1 U16503 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n16989), .A(
        n17182), .ZN(n17170) );
  OAI211_X1 U16504 ( .C1(n16989), .C2(n18129), .A(n17173), .B(n17170), .ZN(
        n13260) );
  OAI211_X1 U16505 ( .C1(n16979), .C2(n18129), .A(n13261), .B(n13260), .ZN(
        n13262) );
  OR4_X1 U16506 ( .A1(n13265), .A2(n13264), .A3(n13263), .A4(n13262), .ZN(
        P3_U2669) );
  NOR2_X1 U16507 ( .A1(n12468), .A2(n16639), .ZN(n13388) );
  AND2_X1 U16508 ( .A1(n13388), .A2(n16608), .ZN(n19393) );
  INV_X1 U16509 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n20215) );
  INV_X1 U16510 ( .A(n13275), .ZN(n13266) );
  OAI211_X1 U16511 ( .C1(n19393), .C2(n20215), .A(n13266), .B(n19193), .ZN(
        P2_U2814) );
  INV_X1 U16512 ( .A(n13344), .ZN(n13268) );
  NOR3_X1 U16513 ( .A1(n13268), .A2(n13343), .A3(n13267), .ZN(n16617) );
  NOR2_X1 U16514 ( .A1(n16617), .A2(n16639), .ZN(n20192) );
  INV_X1 U16515 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13270) );
  OAI21_X1 U16516 ( .B1(n20192), .B2(n13270), .A(n13269), .ZN(P2_U2819) );
  INV_X1 U16517 ( .A(n20198), .ZN(n13273) );
  OAI21_X1 U16518 ( .B1(n13271), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n13273), 
        .ZN(n13272) );
  OAI21_X1 U16519 ( .B1(n13274), .B2(n13273), .A(n13272), .ZN(P2_U3612) );
  INV_X1 U16520 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n14046) );
  INV_X1 U16521 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13276) );
  OAI21_X1 U16522 ( .B1(n12030), .B2(n20202), .A(n13275), .ZN(n13287) );
  INV_X1 U16523 ( .A(n13287), .ZN(n13291) );
  NAND3_X1 U16524 ( .A1(n13275), .A2(n20202), .A3(n10648), .ZN(n13277) );
  AOI22_X1 U16525 ( .A1(n13751), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13753), .ZN(n14043) );
  OAI222_X1 U16526 ( .A1(n14046), .A2(n13389), .B1(n13276), .B2(n13291), .C1(
        n13277), .C2(n14043), .ZN(P2_U2982) );
  INV_X2 U16527 ( .A(n13389), .ZN(n19487) );
  AOI22_X1 U16528 ( .A1(n19487), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n13287), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13279) );
  AOI22_X1 U16529 ( .A1(n13751), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n13753), .ZN(n15309) );
  INV_X1 U16530 ( .A(n15309), .ZN(n13278) );
  NAND2_X1 U16531 ( .A1(n19482), .A2(n13278), .ZN(n13283) );
  NAND2_X1 U16532 ( .A1(n13279), .A2(n13283), .ZN(P2_U2979) );
  AOI22_X1 U16533 ( .A1(n19487), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n13287), 
        .B2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13282) );
  INV_X1 U16534 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16745) );
  OR2_X1 U16535 ( .A1(n15293), .A2(n16745), .ZN(n13281) );
  NAND2_X1 U16536 ( .A1(n15293), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13280) );
  NAND2_X1 U16537 ( .A1(n13281), .A2(n13280), .ZN(n15327) );
  NAND2_X1 U16538 ( .A1(n19482), .A2(n15327), .ZN(n13298) );
  NAND2_X1 U16539 ( .A1(n13282), .A2(n13298), .ZN(P2_U2962) );
  AOI22_X1 U16540 ( .A1(n19487), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n13287), 
        .B2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13284) );
  NAND2_X1 U16541 ( .A1(n13284), .A2(n13283), .ZN(P2_U2964) );
  AOI22_X1 U16542 ( .A1(n19487), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13287), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n13285) );
  AOI22_X1 U16543 ( .A1(n13751), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13753), .ZN(n19574) );
  INV_X1 U16544 ( .A(n19574), .ZN(n13952) );
  NAND2_X1 U16545 ( .A1(n19482), .A2(n13952), .ZN(n13320) );
  NAND2_X1 U16546 ( .A1(n13285), .A2(n13320), .ZN(P2_U2971) );
  AOI22_X1 U16547 ( .A1(n19487), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13287), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13286) );
  OAI22_X1 U16548 ( .A1(n13753), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13751), .ZN(n19586) );
  INV_X1 U16549 ( .A(n19586), .ZN(n16411) );
  NAND2_X1 U16550 ( .A1(n19482), .A2(n16411), .ZN(n13300) );
  NAND2_X1 U16551 ( .A1(n13286), .A2(n13300), .ZN(P2_U2959) );
  AOI22_X1 U16552 ( .A1(n19487), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n13287), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13290) );
  INV_X1 U16553 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16747) );
  OR2_X1 U16554 ( .A1(n15293), .A2(n16747), .ZN(n13289) );
  NAND2_X1 U16555 ( .A1(n15293), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13288) );
  NAND2_X1 U16556 ( .A1(n13289), .A2(n13288), .ZN(n15340) );
  NAND2_X1 U16557 ( .A1(n19482), .A2(n15340), .ZN(n13306) );
  NAND2_X1 U16558 ( .A1(n13290), .A2(n13306), .ZN(P2_U2961) );
  INV_X1 U16559 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19460) );
  INV_X1 U16560 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16749) );
  INV_X1 U16561 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17655) );
  AOI22_X1 U16562 ( .A1(n13751), .A2(n16749), .B1(n17655), .B2(n13753), .ZN(
        n19433) );
  NAND2_X1 U16563 ( .A1(n19482), .A2(n19433), .ZN(n13318) );
  NAND2_X1 U16564 ( .A1(n19486), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13292) );
  OAI211_X1 U16565 ( .C1(n19460), .C2(n13389), .A(n13318), .B(n13292), .ZN(
        P2_U2975) );
  INV_X1 U16566 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19454) );
  INV_X1 U16567 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16743) );
  OR2_X1 U16568 ( .A1(n15293), .A2(n16743), .ZN(n13294) );
  NAND2_X1 U16569 ( .A1(n15293), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13293) );
  NAND2_X1 U16570 ( .A1(n13294), .A2(n13293), .ZN(n19429) );
  NAND2_X1 U16571 ( .A1(n19482), .A2(n19429), .ZN(n13297) );
  NAND2_X1 U16572 ( .A1(n19486), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13295) );
  OAI211_X1 U16573 ( .C1(n19454), .C2(n13389), .A(n13297), .B(n13295), .ZN(
        P2_U2978) );
  INV_X1 U16574 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n13404) );
  NAND2_X1 U16575 ( .A1(n19486), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13296) );
  OAI211_X1 U16576 ( .C1(n13404), .C2(n13389), .A(n13297), .B(n13296), .ZN(
        P2_U2963) );
  AOI22_X1 U16577 ( .A1(n19487), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n19486), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13299) );
  NAND2_X1 U16578 ( .A1(n13299), .A2(n13298), .ZN(P2_U2977) );
  AOI22_X1 U16579 ( .A1(n19487), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n19486), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n13301) );
  NAND2_X1 U16580 ( .A1(n13301), .A2(n13300), .ZN(P2_U2974) );
  AOI22_X1 U16581 ( .A1(n19487), .A2(P2_EAX_REG_0__SCAN_IN), .B1(n19486), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n13303) );
  AOI22_X1 U16582 ( .A1(n13751), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13753), .ZN(n14305) );
  INV_X1 U16583 ( .A(n14305), .ZN(n13302) );
  NAND2_X1 U16584 ( .A1(n19482), .A2(n13302), .ZN(n13308) );
  NAND2_X1 U16585 ( .A1(n13303), .A2(n13308), .ZN(P2_U2967) );
  AOI22_X1 U16586 ( .A1(n19487), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n19486), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n13305) );
  AOI22_X1 U16587 ( .A1(n13751), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13753), .ZN(n19579) );
  INV_X1 U16588 ( .A(n19579), .ZN(n13304) );
  NAND2_X1 U16589 ( .A1(n19482), .A2(n13304), .ZN(n13314) );
  NAND2_X1 U16590 ( .A1(n13305), .A2(n13314), .ZN(P2_U2973) );
  AOI22_X1 U16591 ( .A1(n19487), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n19486), .B2(
        P2_LWORD_REG_9__SCAN_IN), .ZN(n13307) );
  NAND2_X1 U16592 ( .A1(n13307), .A2(n13306), .ZN(P2_U2976) );
  AOI22_X1 U16593 ( .A1(n19487), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13309) );
  NAND2_X1 U16594 ( .A1(n13309), .A2(n13308), .ZN(P2_U2952) );
  AOI22_X1 U16595 ( .A1(n19487), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n19486), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13310) );
  AOI22_X1 U16596 ( .A1(n13751), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13753), .ZN(n19566) );
  INV_X1 U16597 ( .A(n19566), .ZN(n13583) );
  NAND2_X1 U16598 ( .A1(n19482), .A2(n13583), .ZN(n13326) );
  NAND2_X1 U16599 ( .A1(n13310), .A2(n13326), .ZN(P2_U2969) );
  AOI22_X1 U16600 ( .A1(n19487), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13311) );
  AOI22_X1 U16601 ( .A1(n13751), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13753), .ZN(n15353) );
  INV_X1 U16602 ( .A(n15353), .ZN(n14053) );
  NAND2_X1 U16603 ( .A1(n19482), .A2(n14053), .ZN(n13312) );
  NAND2_X1 U16604 ( .A1(n13311), .A2(n13312), .ZN(P2_U2957) );
  AOI22_X1 U16605 ( .A1(n19487), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n19486), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n13313) );
  NAND2_X1 U16606 ( .A1(n13313), .A2(n13312), .ZN(P2_U2972) );
  AOI22_X1 U16607 ( .A1(n19487), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13315) );
  NAND2_X1 U16608 ( .A1(n13315), .A2(n13314), .ZN(P2_U2958) );
  AOI22_X1 U16609 ( .A1(n19487), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n19486), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13316) );
  AOI22_X1 U16610 ( .A1(n13751), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13753), .ZN(n19570) );
  INV_X1 U16611 ( .A(n19570), .ZN(n13732) );
  NAND2_X1 U16612 ( .A1(n19482), .A2(n13732), .ZN(n13322) );
  NAND2_X1 U16613 ( .A1(n13316), .A2(n13322), .ZN(P2_U2970) );
  AOI22_X1 U16614 ( .A1(n19487), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13317) );
  AOI22_X1 U16615 ( .A1(n13751), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13753), .ZN(n14369) );
  INV_X1 U16616 ( .A(n14369), .ZN(n13454) );
  NAND2_X1 U16617 ( .A1(n19482), .A2(n13454), .ZN(n13324) );
  NAND2_X1 U16618 ( .A1(n13317), .A2(n13324), .ZN(P2_U2953) );
  AOI22_X1 U16619 ( .A1(n19487), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13319) );
  NAND2_X1 U16620 ( .A1(n13319), .A2(n13318), .ZN(P2_U2960) );
  AOI22_X1 U16621 ( .A1(n19487), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13321) );
  NAND2_X1 U16622 ( .A1(n13321), .A2(n13320), .ZN(P2_U2956) );
  AOI22_X1 U16623 ( .A1(n19487), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13323) );
  NAND2_X1 U16624 ( .A1(n13323), .A2(n13322), .ZN(P2_U2955) );
  AOI22_X1 U16625 ( .A1(n19487), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n19486), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13325) );
  NAND2_X1 U16626 ( .A1(n13325), .A2(n13324), .ZN(P2_U2968) );
  AOI22_X1 U16627 ( .A1(n19487), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13327) );
  NAND2_X1 U16628 ( .A1(n13327), .A2(n13326), .ZN(P2_U2954) );
  XNOR2_X1 U16629 ( .A(n16584), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13328) );
  XNOR2_X1 U16630 ( .A(n15234), .B(n13328), .ZN(n19550) );
  OR2_X1 U16631 ( .A1(n13329), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13331) );
  NAND2_X1 U16632 ( .A1(n13331), .A2(n13330), .ZN(n19555) );
  INV_X1 U16633 ( .A(n19555), .ZN(n13332) );
  AND2_X1 U16634 ( .A1(n19517), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n19558) );
  AOI21_X1 U16635 ( .B1(n19507), .B2(n13332), .A(n19558), .ZN(n13334) );
  NAND2_X1 U16636 ( .A1(n16494), .A2(n15229), .ZN(n13333) );
  OAI211_X1 U16637 ( .C1(n15229), .C2(n16506), .A(n13334), .B(n13333), .ZN(
        n13335) );
  AOI21_X1 U16638 ( .B1(n12279), .B2(n19550), .A(n13335), .ZN(n13336) );
  OAI21_X1 U16639 ( .B1(n13416), .B2(n16436), .A(n13336), .ZN(P2_U3013) );
  INV_X1 U16640 ( .A(n13374), .ZN(n13337) );
  NAND2_X1 U16641 ( .A1(n13337), .A2(n13601), .ZN(n13357) );
  INV_X1 U16642 ( .A(n13357), .ZN(n13339) );
  INV_X1 U16643 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21011) );
  NAND3_X1 U16644 ( .A1(n13338), .A2(n13601), .A3(n13597), .ZN(n13459) );
  NAND2_X1 U16645 ( .A1(n20696), .A2(n13985), .ZN(n20223) );
  OAI211_X1 U16646 ( .C1(n13339), .C2(n21011), .A(n13459), .B(n20223), .ZN(
        P1_U2801) );
  NOR2_X1 U16647 ( .A1(n12468), .A2(n13340), .ZN(n13341) );
  NAND2_X1 U16648 ( .A1(n13342), .A2(n13341), .ZN(n13349) );
  NAND2_X1 U16649 ( .A1(n13745), .A2(n16613), .ZN(n13414) );
  NAND2_X1 U16650 ( .A1(n13344), .A2(n13343), .ZN(n13345) );
  AND4_X1 U16651 ( .A1(n13347), .A2(n13346), .A3(n13414), .A4(n13345), .ZN(
        n13348) );
  NAND2_X1 U16652 ( .A1(n16620), .A2(n13350), .ZN(n13352) );
  NOR2_X1 U16653 ( .A1(n20201), .A2(n20174), .ZN(n16641) );
  AOI22_X1 U16654 ( .A1(n20201), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n16641), 
        .B2(P2_FLUSH_REG_SCAN_IN), .ZN(n13351) );
  NAND2_X1 U16655 ( .A1(n13352), .A2(n13351), .ZN(n15820) );
  INV_X1 U16656 ( .A(n13353), .ZN(n13354) );
  NOR3_X1 U16657 ( .A1(n12468), .A2(n13354), .A3(n10648), .ZN(n16614) );
  NAND3_X1 U16658 ( .A1(n15820), .A2(n15799), .A3(n16614), .ZN(n13355) );
  OAI21_X1 U16659 ( .B1(n15820), .B2(n12270), .A(n13355), .ZN(P2_U3595) );
  INV_X1 U16660 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n13356) );
  AND2_X1 U16661 ( .A1(n20223), .A2(n13356), .ZN(n13359) );
  OAI21_X1 U16662 ( .B1(n11785), .B2(n13371), .A(n20904), .ZN(n13358) );
  OAI21_X1 U16663 ( .B1(n13359), .B2(n20904), .A(n13358), .ZN(P1_U3487) );
  OAI21_X1 U16664 ( .B1(n13362), .B2(n13361), .A(n13360), .ZN(n13363) );
  INV_X1 U16665 ( .A(n13363), .ZN(n19545) );
  OAI21_X1 U16666 ( .B1(n13366), .B2(n13365), .A(n13364), .ZN(n19548) );
  NOR2_X1 U16667 ( .A1(n19324), .A2(n10734), .ZN(n19536) );
  NOR2_X1 U16668 ( .A1(n19501), .A2(n15221), .ZN(n13367) );
  AOI211_X1 U16669 ( .C1(n19503), .C2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n19536), .B(n13367), .ZN(n13368) );
  OAI21_X1 U16670 ( .B1(n19548), .B2(n19495), .A(n13368), .ZN(n13369) );
  AOI21_X1 U16671 ( .B1(n12279), .B2(n19545), .A(n13369), .ZN(n13370) );
  OAI21_X1 U16672 ( .B1(n19541), .B2(n16436), .A(n13370), .ZN(P2_U3012) );
  INV_X1 U16673 ( .A(n13338), .ZN(n13373) );
  NOR2_X1 U16674 ( .A1(n13597), .A2(n13371), .ZN(n13372) );
  AOI21_X1 U16675 ( .B1(n13374), .B2(n13373), .A(n13372), .ZN(n20218) );
  INV_X1 U16676 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20814) );
  NAND2_X1 U16677 ( .A1(n13375), .A2(n20814), .ZN(n16023) );
  INV_X1 U16678 ( .A(n16023), .ZN(n13587) );
  NOR2_X1 U16679 ( .A1(n9684), .A2(n13587), .ZN(n13376) );
  NAND2_X1 U16680 ( .A1(n13987), .A2(n13376), .ZN(n13377) );
  NAND2_X1 U16681 ( .A1(n13377), .A2(n20906), .ZN(n20908) );
  NAND2_X1 U16682 ( .A1(n20218), .A2(n20908), .ZN(n15993) );
  AND2_X1 U16683 ( .A1(n15993), .A2(n13601), .ZN(n20227) );
  INV_X1 U16684 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n21056) );
  NAND2_X1 U16685 ( .A1(n13523), .A2(n13378), .ZN(n15991) );
  AND2_X1 U16686 ( .A1(n13509), .A2(n15991), .ZN(n13603) );
  OAI21_X1 U16687 ( .B1(n13989), .B2(n13379), .A(n13603), .ZN(n13380) );
  NAND2_X1 U16688 ( .A1(n13380), .A2(n13521), .ZN(n13383) );
  NAND2_X1 U16689 ( .A1(n11906), .A2(n13593), .ZN(n13382) );
  NAND2_X1 U16690 ( .A1(n13622), .A2(n13597), .ZN(n13381) );
  NAND3_X1 U16691 ( .A1(n13383), .A2(n13382), .A3(n13381), .ZN(n13385) );
  NAND2_X1 U16692 ( .A1(n13385), .A2(n13384), .ZN(n15990) );
  INV_X1 U16693 ( .A(n15990), .ZN(n13386) );
  NAND2_X1 U16694 ( .A1(n20227), .A2(n13386), .ZN(n13387) );
  OAI21_X1 U16695 ( .B1(n20227), .B2(n21056), .A(n13387), .ZN(P1_U3484) );
  INV_X1 U16696 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n14403) );
  INV_X1 U16697 ( .A(n13388), .ZN(n13390) );
  OR2_X1 U16698 ( .A1(n20174), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20195) );
  INV_X2 U16699 ( .A(n20195), .ZN(n19475) );
  AOI22_X1 U16700 ( .A1(n19475), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13394) );
  OAI21_X1 U16701 ( .B1(n14403), .B2(n19439), .A(n13394), .ZN(P2_U2933) );
  INV_X1 U16702 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14368) );
  AOI22_X1 U16703 ( .A1(n19475), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13395) );
  OAI21_X1 U16704 ( .B1(n14368), .B2(n19439), .A(n13395), .ZN(P2_U2934) );
  INV_X1 U16705 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14426) );
  AOI22_X1 U16706 ( .A1(n19475), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13396) );
  OAI21_X1 U16707 ( .B1(n14426), .B2(n19439), .A(n13396), .ZN(P2_U2932) );
  INV_X1 U16708 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n15336) );
  AOI22_X1 U16709 ( .A1(n19475), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13397) );
  OAI21_X1 U16710 ( .B1(n15336), .B2(n19439), .A(n13397), .ZN(P2_U2926) );
  INV_X1 U16711 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13399) );
  AOI22_X1 U16712 ( .A1(n19475), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13398) );
  OAI21_X1 U16713 ( .B1(n13399), .B2(n19439), .A(n13398), .ZN(P2_U2927) );
  INV_X1 U16714 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n14304) );
  AOI22_X1 U16715 ( .A1(n19475), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13400) );
  OAI21_X1 U16716 ( .B1(n14304), .B2(n19439), .A(n13400), .ZN(P2_U2935) );
  INV_X1 U16717 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n15346) );
  AOI22_X1 U16718 ( .A1(n19475), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13401) );
  OAI21_X1 U16719 ( .B1(n15346), .B2(n19439), .A(n13401), .ZN(P2_U2929) );
  INV_X1 U16720 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n15308) );
  AOI22_X1 U16721 ( .A1(n19475), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13402) );
  OAI21_X1 U16722 ( .B1(n15308), .B2(n19439), .A(n13402), .ZN(P2_U2923) );
  AOI22_X1 U16723 ( .A1(n19475), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13403) );
  OAI21_X1 U16724 ( .B1(n13404), .B2(n19439), .A(n13403), .ZN(P2_U2924) );
  INV_X1 U16725 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13406) );
  AOI22_X1 U16726 ( .A1(n19475), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13405) );
  OAI21_X1 U16727 ( .B1(n13406), .B2(n19439), .A(n13405), .ZN(P2_U2925) );
  INV_X1 U16728 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n13408) );
  AOI22_X1 U16729 ( .A1(n19475), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13407) );
  OAI21_X1 U16730 ( .B1(n13408), .B2(n19439), .A(n13407), .ZN(P2_U2928) );
  INV_X1 U16731 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15352) );
  AOI22_X1 U16732 ( .A1(n19475), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13409) );
  OAI21_X1 U16733 ( .B1(n15352), .B2(n19439), .A(n13409), .ZN(P2_U2930) );
  INV_X1 U16734 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n15368) );
  AOI22_X1 U16735 ( .A1(n19475), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13410) );
  OAI21_X1 U16736 ( .B1(n15368), .B2(n19439), .A(n13410), .ZN(P2_U2931) );
  AOI21_X2 U16737 ( .B1(n13414), .B2(n15789), .A(n16639), .ZN(n19415) );
  MUX2_X1 U16738 ( .A(n15230), .B(n13416), .S(n19406), .Z(n13417) );
  OAI21_X1 U16739 ( .B1(n20166), .B2(n19403), .A(n13417), .ZN(P2_U2886) );
  INV_X1 U16740 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13420) );
  AND2_X1 U16741 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19920), .ZN(n13419) );
  OAI211_X1 U16742 ( .C1(n12030), .C2(n13420), .A(n19578), .B(n13419), .ZN(
        n13421) );
  INV_X1 U16743 ( .A(n13421), .ZN(n13422) );
  MUX2_X1 U16744 ( .A(n10858), .B(n13423), .S(n19406), .Z(n13424) );
  OAI21_X1 U16745 ( .B1(n20177), .B2(n19403), .A(n13424), .ZN(P2_U2887) );
  INV_X1 U16746 ( .A(n13425), .ZN(n13426) );
  INV_X1 U16747 ( .A(n19434), .ZN(n14044) );
  OAI21_X1 U16748 ( .B1(n13429), .B2(n13428), .A(n13427), .ZN(n19380) );
  INV_X1 U16749 ( .A(n19380), .ZN(n16583) );
  NOR2_X1 U16750 ( .A1(n20177), .A2(n19380), .ZN(n13453) );
  INV_X1 U16751 ( .A(n13453), .ZN(n13430) );
  INV_X1 U16752 ( .A(n15373), .ZN(n16413) );
  OAI211_X1 U16753 ( .C1(n19394), .C2(n16583), .A(n13430), .B(n16413), .ZN(
        n13432) );
  AOI22_X1 U16754 ( .A1(n19417), .A2(n16583), .B1(n19432), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n13431) );
  OAI211_X1 U16755 ( .C1(n14305), .C2(n14044), .A(n13432), .B(n13431), .ZN(
        P2_U2919) );
  AOI21_X1 U16756 ( .B1(n13435), .B2(n16559), .A(n13434), .ZN(n13436) );
  INV_X1 U16757 ( .A(n13436), .ZN(n15752) );
  AOI22_X1 U16758 ( .A1(n19434), .A2(n15340), .B1(n19432), .B2(
        P2_EAX_REG_9__SCAN_IN), .ZN(n13437) );
  OAI21_X1 U16759 ( .B1(n19437), .B2(n15752), .A(n13437), .ZN(P2_U2910) );
  XOR2_X1 U16760 ( .A(n13439), .B(n13438), .Z(n15762) );
  INV_X1 U16761 ( .A(n15762), .ZN(n19355) );
  INV_X1 U16762 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19462) );
  OAI222_X1 U16763 ( .A1(n19355), .A2(n19437), .B1(n14044), .B2(n19586), .C1(
        n19428), .C2(n19462), .ZN(P2_U2912) );
  INV_X1 U16764 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n13444) );
  NOR2_X1 U16765 ( .A1(n13441), .A2(n13440), .ZN(n13442) );
  OR2_X1 U16766 ( .A1(n13443), .A2(n13442), .ZN(n14357) );
  OAI222_X1 U16767 ( .A1(n13444), .A2(n19428), .B1(n14044), .B2(n19579), .C1(
        n14357), .C2(n19437), .ZN(P2_U2913) );
  INV_X1 U16768 ( .A(n15327), .ZN(n13448) );
  OR2_X1 U16769 ( .A1(n13445), .A2(n13434), .ZN(n13447) );
  NAND2_X1 U16770 ( .A1(n13447), .A2(n13446), .ZN(n19333) );
  INV_X1 U16771 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19456) );
  OAI222_X1 U16772 ( .A1(n14044), .A2(n13448), .B1(n19333), .B2(n19437), .C1(
        n19428), .C2(n19456), .ZN(P2_U2909) );
  OAI21_X1 U16773 ( .B1(n13451), .B2(n13450), .A(n13449), .ZN(n20171) );
  INV_X1 U16774 ( .A(n20171), .ZN(n19553) );
  NAND2_X1 U16775 ( .A1(n20166), .A2(n19553), .ZN(n13574) );
  OAI21_X1 U16776 ( .B1(n20166), .B2(n19553), .A(n13574), .ZN(n13452) );
  NOR2_X1 U16777 ( .A1(n13452), .A2(n13453), .ZN(n13576) );
  AOI21_X1 U16778 ( .B1(n13453), .B2(n13452), .A(n13576), .ZN(n13457) );
  AOI22_X1 U16779 ( .A1(n19417), .A2(n20171), .B1(n19432), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n13456) );
  NAND2_X1 U16780 ( .A1(n19434), .A2(n13454), .ZN(n13455) );
  OAI211_X1 U16781 ( .C1(n13457), .C2(n15373), .A(n13456), .B(n13455), .ZN(
        P2_U2918) );
  AND2_X1 U16782 ( .A1(n20910), .A2(n16022), .ZN(n13458) );
  OR2_X2 U16783 ( .A1(n13459), .A2(n13458), .ZN(n20368) );
  INV_X1 U16784 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13765) );
  NAND2_X1 U16785 ( .A1(n20368), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13460) );
  MUX2_X1 U16786 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n13800), .Z(
        n14757) );
  NAND2_X1 U16787 ( .A1(n13681), .A2(n14757), .ZN(n20360) );
  OAI211_X1 U16788 ( .C1(n13650), .C2(n13765), .A(n13460), .B(n20360), .ZN(
        P1_U2947) );
  INV_X1 U16789 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13558) );
  NAND2_X1 U16790 ( .A1(n20368), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n13461) );
  MUX2_X1 U16791 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n13800), .Z(
        n14750) );
  NAND2_X1 U16792 ( .A1(n13681), .A2(n14750), .ZN(n20364) );
  OAI211_X1 U16793 ( .C1(n13650), .C2(n13558), .A(n13461), .B(n20364), .ZN(
        P1_U2949) );
  INV_X1 U16794 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13552) );
  NAND2_X1 U16795 ( .A1(n20368), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13462) );
  MUX2_X1 U16796 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n13800), .Z(
        n14753) );
  NAND2_X1 U16797 ( .A1(n13681), .A2(n14753), .ZN(n20362) );
  OAI211_X1 U16798 ( .C1(n13650), .C2(n13552), .A(n13462), .B(n20362), .ZN(
        P1_U2948) );
  INV_X1 U16799 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13556) );
  NAND2_X1 U16800 ( .A1(n20368), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13463) );
  MUX2_X1 U16801 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n13800), .Z(
        n14760) );
  NAND2_X1 U16802 ( .A1(n13681), .A2(n14760), .ZN(n20358) );
  OAI211_X1 U16803 ( .C1(n13650), .C2(n13556), .A(n13463), .B(n20358), .ZN(
        P1_U2946) );
  INV_X1 U16804 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13542) );
  NAND2_X1 U16805 ( .A1(n20368), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13464) );
  NAND2_X1 U16806 ( .A1(n13681), .A2(n14449), .ZN(n20370) );
  OAI211_X1 U16807 ( .C1(n13650), .C2(n13542), .A(n13464), .B(n20370), .ZN(
        P1_U2951) );
  INV_X1 U16808 ( .A(n13465), .ZN(n13467) );
  INV_X1 U16809 ( .A(n13478), .ZN(n13469) );
  INV_X1 U16810 ( .A(n13466), .ZN(n13468) );
  MUX2_X1 U16811 ( .A(n13472), .B(n10862), .S(n16392), .Z(n13473) );
  OAI21_X1 U16812 ( .B1(n15819), .B2(n19403), .A(n13473), .ZN(P2_U2884) );
  INV_X1 U16813 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14480) );
  INV_X1 U16814 ( .A(n13681), .ZN(n13476) );
  INV_X1 U16815 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13474) );
  NOR2_X1 U16816 ( .A1(n13799), .A2(n13474), .ZN(n13475) );
  AOI21_X1 U16817 ( .B1(DATAI_15_), .B2(n13799), .A(n13475), .ZN(n14481) );
  INV_X1 U16818 ( .A(n20368), .ZN(n13651) );
  INV_X1 U16819 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20326) );
  OAI222_X1 U16820 ( .A1(n13650), .A2(n14480), .B1(n13476), .B2(n14481), .C1(
        n13651), .C2(n20326), .ZN(P1_U2967) );
  MUX2_X1 U16821 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n9722), .S(n19406), .Z(n13479) );
  AOI21_X1 U16822 ( .B1(n15796), .B2(n19411), .A(n13479), .ZN(n13480) );
  INV_X1 U16823 ( .A(n13480), .ZN(P2_U2885) );
  INV_X1 U16824 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13554) );
  NAND2_X1 U16825 ( .A1(n20368), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13482) );
  NOR2_X1 U16826 ( .A1(n13800), .A2(DATAI_8_), .ZN(n13481) );
  AOI21_X1 U16827 ( .B1(n13800), .B2(n16749), .A(n13481), .ZN(n14764) );
  NAND2_X1 U16828 ( .A1(n13681), .A2(n14764), .ZN(n13483) );
  OAI211_X1 U16829 ( .C1(n13650), .C2(n13554), .A(n13482), .B(n13483), .ZN(
        P1_U2945) );
  INV_X1 U16830 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20342) );
  NAND2_X1 U16831 ( .A1(n20368), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13484) );
  OAI211_X1 U16832 ( .C1(n13650), .C2(n20342), .A(n13484), .B(n13483), .ZN(
        P1_U2960) );
  INV_X1 U16833 ( .A(n13485), .ZN(n13486) );
  AOI21_X1 U16834 ( .B1(n13488), .B2(n13487), .A(n13486), .ZN(n13988) );
  OAI21_X1 U16835 ( .B1(n13490), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13489), .ZN(n13723) );
  NAND2_X1 U16836 ( .A1(n16285), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13716) );
  OAI21_X1 U16837 ( .B1(n16173), .B2(n13491), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13492) );
  OAI211_X1 U16838 ( .C1(n13723), .C2(n20226), .A(n13716), .B(n13492), .ZN(
        n13493) );
  AOI21_X1 U16839 ( .B1(n13988), .B2(n14887), .A(n13493), .ZN(n13494) );
  INV_X1 U16840 ( .A(n13494), .ZN(P1_U2999) );
  AND2_X1 U16841 ( .A1(n13497), .A2(n13802), .ZN(n13498) );
  AND2_X1 U16842 ( .A1(n13499), .A2(n13498), .ZN(n13524) );
  INV_X1 U16843 ( .A(n13524), .ZN(n13502) );
  NAND2_X1 U16844 ( .A1(n13500), .A2(n13992), .ZN(n13501) );
  OAI211_X1 U16845 ( .C1(n13503), .C2(n13987), .A(n13502), .B(n13501), .ZN(
        n13613) );
  NAND2_X1 U16846 ( .A1(n13504), .A2(n9710), .ZN(n13505) );
  NOR2_X1 U16847 ( .A1(n13613), .A2(n13505), .ZN(n13507) );
  NAND2_X1 U16848 ( .A1(n13507), .A2(n13506), .ZN(n15976) );
  INV_X1 U16849 ( .A(n15976), .ZN(n13515) );
  XNOR2_X1 U16850 ( .A(n13508), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13517) );
  NOR2_X1 U16851 ( .A1(n14060), .A2(n13517), .ZN(n13511) );
  INV_X1 U16852 ( .A(n13509), .ZN(n13510) );
  OR2_X1 U16853 ( .A1(n13622), .A2(n13510), .ZN(n14070) );
  AOI22_X1 U16854 ( .A1(n13515), .A2(n13511), .B1(n14070), .B2(n13517), .ZN(
        n13514) );
  NAND2_X1 U16855 ( .A1(n15977), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13512) );
  NAND2_X1 U16856 ( .A1(n15977), .A2(n10901), .ZN(n15117) );
  MUX2_X1 U16857 ( .A(n13512), .B(n15117), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13513) );
  OAI211_X1 U16858 ( .C1(n13496), .C2(n13515), .A(n13514), .B(n13513), .ZN(
        n14057) );
  INV_X1 U16859 ( .A(n20897), .ZN(n13519) );
  INV_X1 U16860 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13705) );
  NOR2_X1 U16861 ( .A1(n13985), .A2(n13705), .ZN(n15122) );
  INV_X1 U16862 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13624) );
  INV_X1 U16863 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13516) );
  AOI22_X1 U16864 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13624), .B2(n13516), .ZN(
        n15120) );
  INV_X1 U16865 ( .A(n20888), .ZN(n16010) );
  INV_X1 U16866 ( .A(n13517), .ZN(n13518) );
  AOI222_X1 U16867 ( .A1(n14057), .A2(n13519), .B1(n15122), .B2(n15120), .C1(
        n16010), .C2(n13518), .ZN(n13536) );
  AOI22_X1 U16868 ( .A1(n13622), .A2(n13521), .B1(n10191), .B2(n13520), .ZN(
        n13528) );
  OAI211_X1 U16869 ( .C1(n15977), .C2(n13522), .A(n15999), .B(n20906), .ZN(
        n13527) );
  INV_X1 U16870 ( .A(n11906), .ZN(n13526) );
  INV_X1 U16871 ( .A(n13523), .ZN(n13525) );
  AOI21_X1 U16872 ( .B1(n13526), .B2(n13525), .A(n13524), .ZN(n13600) );
  NAND3_X1 U16873 ( .A1(n13528), .A2(n13527), .A3(n13600), .ZN(n13530) );
  NAND2_X1 U16874 ( .A1(n15979), .A2(n13601), .ZN(n13534) );
  INV_X1 U16875 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20957) );
  NAND2_X1 U16876 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16304) );
  NOR3_X1 U16877 ( .A1(n20222), .A2(n20957), .A3(n16304), .ZN(n13532) );
  NOR2_X1 U16878 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20700), .ZN(n13531) );
  NOR2_X1 U16879 ( .A1(n13532), .A2(n13531), .ZN(n13533) );
  NAND2_X1 U16880 ( .A1(n13534), .A2(n13533), .ZN(n20892) );
  INV_X1 U16881 ( .A(n20892), .ZN(n20894) );
  NAND2_X1 U16882 ( .A1(n20894), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13535) );
  OAI21_X1 U16883 ( .B1(n13536), .B2(n20894), .A(n13535), .ZN(P1_U3472) );
  INV_X1 U16884 ( .A(n15977), .ZN(n13537) );
  NAND2_X1 U16885 ( .A1(n13338), .A2(n13596), .ZN(n16001) );
  NAND2_X1 U16886 ( .A1(n13537), .A2(n16001), .ZN(n13540) );
  INV_X1 U16887 ( .A(n15999), .ZN(n13538) );
  NOR2_X1 U16888 ( .A1(n20219), .A2(n13538), .ZN(n13539) );
  NAND2_X1 U16889 ( .A1(n20328), .A2(n13802), .ZN(n13775) );
  NOR2_X4 U16890 ( .A1(n20328), .A2(n20907), .ZN(n20340) );
  INV_X2 U16891 ( .A(n20327), .ZN(n20907) );
  AOI22_X1 U16892 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20340), .B1(n20907), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13541) );
  OAI21_X1 U16893 ( .B1(n13542), .B2(n13775), .A(n13541), .ZN(P1_U2906) );
  AND2_X1 U16894 ( .A1(n14495), .A2(n13543), .ZN(n13544) );
  OR2_X1 U16895 ( .A1(n13544), .A2(n13567), .ZN(n14353) );
  NOR2_X1 U16896 ( .A1(n13545), .A2(n14197), .ZN(n13547) );
  OAI211_X1 U16897 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13547), .A(
        n13546), .B(n19411), .ZN(n13549) );
  NAND2_X1 U16898 ( .A1(n16392), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13548) );
  OAI211_X1 U16899 ( .C1(n14353), .C2(n16392), .A(n13549), .B(n13548), .ZN(
        P2_U2881) );
  INV_X1 U16900 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14744) );
  AOI22_X1 U16901 ( .A1(n20907), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13550) );
  OAI21_X1 U16902 ( .B1(n14744), .B2(n13775), .A(n13550), .ZN(P1_U2907) );
  AOI22_X1 U16903 ( .A1(n20907), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13551) );
  OAI21_X1 U16904 ( .B1(n13552), .B2(n13775), .A(n13551), .ZN(P1_U2909) );
  AOI22_X1 U16905 ( .A1(n20907), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13553) );
  OAI21_X1 U16906 ( .B1(n13554), .B2(n13775), .A(n13553), .ZN(P1_U2912) );
  AOI22_X1 U16907 ( .A1(n20907), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13555) );
  OAI21_X1 U16908 ( .B1(n13556), .B2(n13775), .A(n13555), .ZN(P1_U2911) );
  AOI22_X1 U16909 ( .A1(n20907), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13557) );
  OAI21_X1 U16910 ( .B1(n13558), .B2(n13775), .A(n13557), .ZN(P1_U2908) );
  INV_X1 U16911 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13560) );
  AOI22_X1 U16912 ( .A1(n20907), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13559) );
  OAI21_X1 U16913 ( .B1(n13560), .B2(n13775), .A(n13559), .ZN(P1_U2913) );
  OAI21_X1 U16914 ( .B1(n13562), .B2(n13561), .A(n13696), .ZN(n13703) );
  XNOR2_X1 U16915 ( .A(n13563), .B(n9684), .ZN(n14545) );
  AOI22_X1 U16916 ( .A1(n20320), .A2(n14545), .B1(n14740), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13564) );
  OAI21_X1 U16917 ( .B1(n13703), .B2(n14742), .A(n13564), .ZN(P1_U2871) );
  XOR2_X1 U16918 ( .A(n13546), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13569)
         );
  INV_X1 U16919 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n19352) );
  OAI21_X1 U16920 ( .B1(n13567), .B2(n13566), .A(n13565), .ZN(n19353) );
  MUX2_X1 U16921 ( .A(n19352), .B(n19353), .S(n19406), .Z(n13568) );
  OAI21_X1 U16922 ( .B1(n13569), .B2(n19403), .A(n13568), .ZN(P2_U2880) );
  XNOR2_X1 U16923 ( .A(n13570), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13712) );
  INV_X1 U16924 ( .A(n13703), .ZN(n14542) );
  INV_X1 U16925 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20898) );
  NOR2_X1 U16926 ( .A1(n16238), .A2(n20898), .ZN(n13709) );
  AOI21_X1 U16927 ( .B1(n16173), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13709), .ZN(n13571) );
  OAI21_X1 U16928 ( .B1(n16180), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13571), .ZN(n13572) );
  AOI21_X1 U16929 ( .B1(n14542), .B2(n14887), .A(n13572), .ZN(n13573) );
  OAI21_X1 U16930 ( .B1(n13712), .B2(n20226), .A(n13573), .ZN(P1_U2998) );
  INV_X1 U16931 ( .A(n13574), .ZN(n13575) );
  NOR2_X1 U16932 ( .A1(n13576), .A2(n13575), .ZN(n13582) );
  OAI21_X1 U16933 ( .B1(n13579), .B2(n13578), .A(n13577), .ZN(n20161) );
  INV_X1 U16934 ( .A(n20161), .ZN(n13580) );
  NAND2_X1 U16935 ( .A1(n20158), .A2(n13580), .ZN(n13724) );
  OAI21_X1 U16936 ( .B1(n20158), .B2(n13580), .A(n13724), .ZN(n13581) );
  NOR2_X1 U16937 ( .A1(n13581), .A2(n13582), .ZN(n13726) );
  AOI21_X1 U16938 ( .B1(n13582), .B2(n13581), .A(n13726), .ZN(n13586) );
  AOI22_X1 U16939 ( .A1(n19417), .A2(n20161), .B1(n19432), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n13585) );
  NAND2_X1 U16940 ( .A1(n19434), .A2(n13583), .ZN(n13584) );
  OAI211_X1 U16941 ( .C1(n13586), .C2(n15373), .A(n13585), .B(n13584), .ZN(
        P2_U2917) );
  OAI21_X1 U16942 ( .B1(n13992), .B2(n13587), .A(n20906), .ZN(n13991) );
  OAI211_X1 U16943 ( .C1(n13589), .C2(n13991), .A(n13802), .B(n13588), .ZN(
        n13590) );
  NAND2_X1 U16944 ( .A1(n13590), .A2(n13597), .ZN(n13595) );
  NAND2_X1 U16945 ( .A1(n13992), .A2(n16023), .ZN(n13591) );
  NAND2_X1 U16946 ( .A1(n13591), .A2(n20906), .ZN(n13592) );
  OR2_X1 U16947 ( .A1(n13593), .A2(n13592), .ZN(n13594) );
  MUX2_X1 U16948 ( .A(n13595), .B(n13594), .S(n11036), .Z(n13599) );
  OR3_X1 U16949 ( .A1(n9692), .A2(n13597), .A3(n13596), .ZN(n13598) );
  NAND3_X1 U16950 ( .A1(n13600), .A2(n13599), .A3(n13598), .ZN(n13602) );
  OAI211_X1 U16951 ( .C1(n11035), .C2(n13620), .A(n9700), .B(n13603), .ZN(
        n13605) );
  XNOR2_X1 U16952 ( .A(n9666), .B(n13607), .ZN(n13701) );
  INV_X1 U16953 ( .A(n13608), .ZN(n13610) );
  OAI211_X1 U16954 ( .C1(n13611), .C2(n13802), .A(n13610), .B(n13609), .ZN(
        n13612) );
  OR2_X1 U16955 ( .A1(n13613), .A2(n13612), .ZN(n13614) );
  OAI22_X1 U16956 ( .A1(n16285), .A2(n13623), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13629), .ZN(n14952) );
  INV_X1 U16957 ( .A(n14952), .ZN(n15070) );
  NAND2_X1 U16958 ( .A1(n15053), .A2(n13629), .ZN(n15096) );
  NAND2_X1 U16959 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13615) );
  NAND2_X1 U16960 ( .A1(n15096), .A2(n13615), .ZN(n14228) );
  NAND2_X1 U16961 ( .A1(n15070), .A2(n14228), .ZN(n13633) );
  INV_X1 U16962 ( .A(n13616), .ZN(n13619) );
  INV_X1 U16963 ( .A(n13647), .ZN(n13617) );
  AOI21_X1 U16964 ( .B1(n13619), .B2(n13618), .A(n13617), .ZN(n20302) );
  OAI21_X1 U16965 ( .B1(n13620), .B2(n11033), .A(n16001), .ZN(n13621) );
  INV_X1 U16966 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20824) );
  NOR2_X1 U16967 ( .A1(n16238), .A2(n20824), .ZN(n13628) );
  NOR2_X1 U16968 ( .A1(n13705), .A2(n13624), .ZN(n13625) );
  AOI21_X1 U16969 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14227) );
  AOI21_X1 U16970 ( .B1(n13625), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n14227), .ZN(n13626) );
  NOR2_X1 U16971 ( .A1(n15101), .A2(n13626), .ZN(n13627) );
  AOI211_X1 U16972 ( .C1(n20302), .C2(n16286), .A(n13628), .B(n13627), .ZN(
        n13631) );
  OAI21_X1 U16973 ( .B1(n13629), .B2(n13705), .A(n15053), .ZN(n15103) );
  NAND3_X1 U16974 ( .A1(n15103), .A2(n12351), .A3(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13630) );
  NAND2_X1 U16975 ( .A1(n13631), .A2(n13630), .ZN(n13632) );
  AOI21_X1 U16976 ( .B1(n13633), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n13632), .ZN(n13634) );
  OAI21_X1 U16977 ( .B1(n16222), .B2(n13701), .A(n13634), .ZN(P1_U3029) );
  XNOR2_X1 U16978 ( .A(n13635), .B(n13636), .ZN(n13640) );
  OR2_X1 U16979 ( .A1(n13637), .A2(n13687), .ZN(n13638) );
  NAND2_X1 U16980 ( .A1(n15733), .A2(n13638), .ZN(n15751) );
  MUX2_X1 U16981 ( .A(n10097), .B(n15751), .S(n19406), .Z(n13639) );
  OAI21_X1 U16982 ( .B1(n13640), .B2(n19403), .A(n13639), .ZN(P2_U2878) );
  OAI21_X1 U16983 ( .B1(n13641), .B2(n13238), .A(n16532), .ZN(n19320) );
  INV_X1 U16984 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19452) );
  OAI222_X1 U16985 ( .A1(n14044), .A2(n15309), .B1(n19320), .B2(n19437), .C1(
        n19428), .C2(n19452), .ZN(P2_U2907) );
  OAI21_X1 U16986 ( .B1(n13645), .B2(n13644), .A(n13643), .ZN(n14137) );
  INV_X1 U16987 ( .A(n13791), .ZN(n13646) );
  AOI21_X1 U16988 ( .B1(n13648), .B2(n13647), .A(n13646), .ZN(n14135) );
  AOI22_X1 U16989 ( .A1(n14135), .A2(n20320), .B1(n14740), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n13649) );
  OAI21_X1 U16990 ( .B1(n14137), .B2(n14742), .A(n13649), .ZN(P1_U2869) );
  AOI22_X1 U16991 ( .A1(n20369), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20368), .ZN(n13653) );
  INV_X1 U16992 ( .A(DATAI_7_), .ZN(n21048) );
  INV_X1 U16993 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16751) );
  MUX2_X1 U16994 ( .A(n21048), .B(n16751), .S(n13800), .Z(n14770) );
  INV_X1 U16995 ( .A(n14770), .ZN(n13652) );
  NAND2_X1 U16996 ( .A1(n13681), .A2(n13652), .ZN(n13678) );
  NAND2_X1 U16997 ( .A1(n13653), .A2(n13678), .ZN(P1_U2959) );
  AOI22_X1 U16998 ( .A1(n20369), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20368), .ZN(n13656) );
  NAND2_X1 U16999 ( .A1(n13799), .A2(DATAI_5_), .ZN(n13655) );
  NAND2_X1 U17000 ( .A1(n13800), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13654) );
  AND2_X1 U17001 ( .A1(n13655), .A2(n13654), .ZN(n14112) );
  INV_X1 U17002 ( .A(n14112), .ZN(n14779) );
  NAND2_X1 U17003 ( .A1(n13681), .A2(n14779), .ZN(n13670) );
  NAND2_X1 U17004 ( .A1(n13656), .A2(n13670), .ZN(P1_U2957) );
  AOI22_X1 U17005 ( .A1(n20369), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20368), .ZN(n13658) );
  INV_X1 U17006 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16761) );
  NAND2_X1 U17007 ( .A1(n13800), .A2(n16761), .ZN(n13657) );
  OAI21_X1 U17008 ( .B1(n13800), .B2(DATAI_2_), .A(n13657), .ZN(n13818) );
  INV_X1 U17009 ( .A(n13818), .ZN(n14790) );
  NAND2_X1 U17010 ( .A1(n13681), .A2(n14790), .ZN(n13662) );
  NAND2_X1 U17011 ( .A1(n13658), .A2(n13662), .ZN(P1_U2954) );
  AOI22_X1 U17012 ( .A1(n20369), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20368), .ZN(n13659) );
  MUX2_X1 U17013 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n13800), .Z(
        n14746) );
  NAND2_X1 U17014 ( .A1(n13681), .A2(n14746), .ZN(n20366) );
  NAND2_X1 U17015 ( .A1(n13659), .A2(n20366), .ZN(P1_U2950) );
  AOI22_X1 U17016 ( .A1(n20369), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20368), .ZN(n13661) );
  INV_X1 U17017 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16768) );
  NAND2_X1 U17018 ( .A1(n13800), .A2(n16768), .ZN(n13660) );
  OAI21_X1 U17019 ( .B1(n13800), .B2(DATAI_0_), .A(n13660), .ZN(n13803) );
  INV_X1 U17020 ( .A(n13803), .ZN(n14801) );
  NAND2_X1 U17021 ( .A1(n13681), .A2(n14801), .ZN(n13676) );
  NAND2_X1 U17022 ( .A1(n13661), .A2(n13676), .ZN(P1_U2937) );
  AOI22_X1 U17023 ( .A1(n20369), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20368), .ZN(n13663) );
  NAND2_X1 U17024 ( .A1(n13663), .A2(n13662), .ZN(P1_U2939) );
  AOI22_X1 U17025 ( .A1(n20369), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20368), .ZN(n13665) );
  INV_X1 U17026 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16759) );
  NAND2_X1 U17027 ( .A1(n13800), .A2(n16759), .ZN(n13664) );
  OAI21_X1 U17028 ( .B1(n13800), .B2(DATAI_3_), .A(n13664), .ZN(n13813) );
  INV_X1 U17029 ( .A(n13813), .ZN(n14787) );
  NAND2_X1 U17030 ( .A1(n13681), .A2(n14787), .ZN(n13683) );
  NAND2_X1 U17031 ( .A1(n13665), .A2(n13683), .ZN(P1_U2955) );
  AOI22_X1 U17032 ( .A1(n20369), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20368), .ZN(n13667) );
  INV_X1 U17033 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16753) );
  NAND2_X1 U17034 ( .A1(n13800), .A2(n16753), .ZN(n13666) );
  OAI21_X1 U17035 ( .B1(n13800), .B2(DATAI_6_), .A(n13666), .ZN(n14140) );
  INV_X1 U17036 ( .A(n14140), .ZN(n14776) );
  NAND2_X1 U17037 ( .A1(n13681), .A2(n14776), .ZN(n13674) );
  NAND2_X1 U17038 ( .A1(n13667), .A2(n13674), .ZN(P1_U2958) );
  AOI22_X1 U17039 ( .A1(n20369), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20368), .ZN(n13669) );
  INV_X1 U17040 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16757) );
  NAND2_X1 U17041 ( .A1(n13800), .A2(n16757), .ZN(n13668) );
  OAI21_X1 U17042 ( .B1(n13800), .B2(DATAI_4_), .A(n13668), .ZN(n13853) );
  INV_X1 U17043 ( .A(n13853), .ZN(n14784) );
  NAND2_X1 U17044 ( .A1(n13681), .A2(n14784), .ZN(n13672) );
  NAND2_X1 U17045 ( .A1(n13669), .A2(n13672), .ZN(P1_U2941) );
  AOI22_X1 U17046 ( .A1(n20369), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20368), .ZN(n13671) );
  NAND2_X1 U17047 ( .A1(n13671), .A2(n13670), .ZN(P1_U2942) );
  AOI22_X1 U17048 ( .A1(n20369), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20368), .ZN(n13673) );
  NAND2_X1 U17049 ( .A1(n13673), .A2(n13672), .ZN(P1_U2956) );
  AOI22_X1 U17050 ( .A1(n20369), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20368), .ZN(n13675) );
  NAND2_X1 U17051 ( .A1(n13675), .A2(n13674), .ZN(P1_U2943) );
  AOI22_X1 U17052 ( .A1(n20369), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20368), .ZN(n13677) );
  NAND2_X1 U17053 ( .A1(n13677), .A2(n13676), .ZN(P1_U2952) );
  AOI22_X1 U17054 ( .A1(n20369), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20368), .ZN(n13679) );
  NAND2_X1 U17055 ( .A1(n13679), .A2(n13678), .ZN(P1_U2944) );
  AOI22_X1 U17056 ( .A1(n20369), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20368), .ZN(n13682) );
  INV_X1 U17057 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16763) );
  NAND2_X1 U17058 ( .A1(n13800), .A2(n16763), .ZN(n13680) );
  OAI21_X1 U17059 ( .B1(n13800), .B2(DATAI_1_), .A(n13680), .ZN(n13875) );
  INV_X1 U17060 ( .A(n13875), .ZN(n14795) );
  NAND2_X1 U17061 ( .A1(n13681), .A2(n14795), .ZN(n13685) );
  NAND2_X1 U17062 ( .A1(n13682), .A2(n13685), .ZN(P1_U2953) );
  AOI22_X1 U17063 ( .A1(n20369), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20368), .ZN(n13684) );
  NAND2_X1 U17064 ( .A1(n13684), .A2(n13683), .ZN(P1_U2940) );
  AOI22_X1 U17065 ( .A1(n20369), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20368), .ZN(n13686) );
  NAND2_X1 U17066 ( .A1(n13686), .A2(n13685), .ZN(P1_U2938) );
  AOI21_X1 U17067 ( .B1(n13688), .B2(n13565), .A(n13687), .ZN(n19341) );
  INV_X1 U17068 ( .A(n19341), .ZN(n15543) );
  INV_X1 U17069 ( .A(n13635), .ZN(n13690) );
  OAI211_X1 U17070 ( .C1(n13689), .C2(n13691), .A(n13690), .B(n19411), .ZN(
        n13693) );
  NAND2_X1 U17071 ( .A1(n16392), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13692) );
  OAI211_X1 U17072 ( .C1(n15543), .C2(n16392), .A(n13693), .B(n13692), .ZN(
        P2_U2879) );
  INV_X1 U17073 ( .A(n13694), .ZN(n13695) );
  AOI21_X1 U17074 ( .B1(n13697), .B2(n13696), .A(n13695), .ZN(n20315) );
  AOI22_X1 U17075 ( .A1(n16173), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n16285), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13698) );
  OAI21_X1 U17076 ( .B1(n16180), .B2(n20305), .A(n13698), .ZN(n13699) );
  AOI21_X1 U17077 ( .B1(n20315), .B2(n14887), .A(n13699), .ZN(n13700) );
  OAI21_X1 U17078 ( .B1(n20226), .B2(n13701), .A(n13700), .ZN(P1_U2997) );
  INV_X1 U17079 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20354) );
  OAI222_X1 U17080 ( .A1(n14490), .A2(n13875), .B1(n14743), .B2(n20354), .C1(
        n14793), .C2(n13703), .ZN(P1_U2903) );
  INV_X1 U17081 ( .A(n15096), .ZN(n14229) );
  NOR2_X1 U17082 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14963), .ZN(
        n13704) );
  NOR2_X1 U17083 ( .A1(n16270), .A2(n13704), .ZN(n13707) );
  INV_X1 U17084 ( .A(n15101), .ZN(n13717) );
  AOI21_X1 U17085 ( .B1(n13717), .B2(n13705), .A(n14952), .ZN(n13719) );
  INV_X1 U17086 ( .A(n13719), .ZN(n13706) );
  MUX2_X1 U17087 ( .A(n13707), .B(n13706), .S(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n13708) );
  INV_X1 U17088 ( .A(n13708), .ZN(n13711) );
  AOI21_X1 U17089 ( .B1(n16286), .B2(n14545), .A(n13709), .ZN(n13710) );
  OAI211_X1 U17090 ( .C1(n13712), .C2(n16222), .A(n13711), .B(n13710), .ZN(
        P1_U3030) );
  INV_X1 U17091 ( .A(n20315), .ZN(n13736) );
  AOI22_X1 U17092 ( .A1(n20302), .A2(n20320), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n14740), .ZN(n13713) );
  OAI21_X1 U17093 ( .B1(n13736), .B2(n14742), .A(n13713), .ZN(P1_U2870) );
  OR2_X1 U17094 ( .A1(n14523), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13714) );
  AND2_X1 U17095 ( .A1(n13715), .A2(n13714), .ZN(n13995) );
  INV_X1 U17096 ( .A(n13716), .ZN(n13721) );
  NOR3_X1 U17097 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13717), .A3(
        n14961), .ZN(n13718) );
  AOI21_X1 U17098 ( .B1(n15053), .B2(n13719), .A(n13718), .ZN(n13720) );
  AOI211_X1 U17099 ( .C1(n16286), .C2(n13995), .A(n13721), .B(n13720), .ZN(
        n13722) );
  OAI21_X1 U17100 ( .B1(n13723), .B2(n16222), .A(n13722), .ZN(P1_U3031) );
  INV_X1 U17101 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20350) );
  OAI222_X1 U17102 ( .A1(n14490), .A2(n13813), .B1(n14743), .B2(n20350), .C1(
        n14793), .C2(n14137), .ZN(P1_U2901) );
  INV_X1 U17103 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20357) );
  INV_X1 U17104 ( .A(n13988), .ZN(n13737) );
  OAI222_X1 U17105 ( .A1(n14490), .A2(n13803), .B1(n14743), .B2(n20357), .C1(
        n14793), .C2(n13737), .ZN(P1_U2904) );
  INV_X1 U17106 ( .A(n13724), .ZN(n13725) );
  NOR2_X1 U17107 ( .A1(n13726), .A2(n13725), .ZN(n13731) );
  INV_X1 U17108 ( .A(n13727), .ZN(n13728) );
  XNOR2_X1 U17109 ( .A(n13729), .B(n13728), .ZN(n20153) );
  XNOR2_X1 U17110 ( .A(n20154), .B(n20153), .ZN(n13730) );
  NOR2_X1 U17111 ( .A1(n13731), .A2(n13730), .ZN(n13943) );
  AOI21_X1 U17112 ( .B1(n13731), .B2(n13730), .A(n13943), .ZN(n13735) );
  AOI22_X1 U17113 ( .A1(n19434), .A2(n13732), .B1(n19432), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n13734) );
  NAND2_X1 U17114 ( .A1(n19417), .A2(n20153), .ZN(n13733) );
  OAI211_X1 U17115 ( .C1(n13735), .C2(n15373), .A(n13734), .B(n13733), .ZN(
        P2_U2916) );
  INV_X1 U17116 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20352) );
  OAI222_X1 U17117 ( .A1(n14490), .A2(n13818), .B1(n14743), .B2(n20352), .C1(
        n14793), .C2(n13736), .ZN(P1_U2902) );
  INV_X1 U17118 ( .A(n13995), .ZN(n13738) );
  OAI222_X1 U17119 ( .A1(n13738), .A2(n14737), .B1(n20324), .B2(n11788), .C1(
        n13737), .C2(n14742), .ZN(P1_U2872) );
  AND2_X1 U17120 ( .A1(n20154), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19992) );
  INV_X1 U17121 ( .A(n19643), .ZN(n13739) );
  NAND2_X1 U17122 ( .A1(n19992), .A2(n13739), .ZN(n13740) );
  NOR2_X1 U17123 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20156), .ZN(
        n19787) );
  INV_X1 U17124 ( .A(n19787), .ZN(n19854) );
  OR2_X1 U17125 ( .A1(n10356), .A2(n19854), .ZN(n13754) );
  NAND2_X1 U17126 ( .A1(n13740), .A2(n13754), .ZN(n13750) );
  INV_X1 U17127 ( .A(n19755), .ZN(n13741) );
  NAND2_X1 U17128 ( .A1(n19787), .A2(n13741), .ZN(n13742) );
  INV_X1 U17129 ( .A(n13742), .ZN(n19902) );
  AND2_X1 U17130 ( .A1(n13742), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13743) );
  NAND2_X1 U17131 ( .A1(n13744), .A2(n13743), .ZN(n13756) );
  INV_X1 U17132 ( .A(n16633), .ZN(n20200) );
  AND2_X1 U17133 ( .A1(n20200), .A2(n20174), .ZN(n13746) );
  OAI211_X1 U17134 ( .C1(n19902), .C2(n19920), .A(n13756), .B(n19995), .ZN(
        n13748) );
  INV_X1 U17135 ( .A(n13748), .ZN(n13749) );
  NAND2_X1 U17136 ( .A1(n13750), .A2(n13749), .ZN(n19898) );
  INV_X1 U17137 ( .A(n19898), .ZN(n19908) );
  INV_X1 U17138 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13759) );
  AOI22_X1 U17139 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19587), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19588), .ZN(n19926) );
  NAND2_X1 U17140 ( .A1(n20154), .A2(n19394), .ZN(n19818) );
  AOI22_X1 U17141 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19588), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19587), .ZN(n19864) );
  INV_X1 U17142 ( .A(n19864), .ZN(n20011) );
  AOI22_X1 U17143 ( .A1(n19904), .A2(n20012), .B1(n19914), .B2(n20011), .ZN(
        n13758) );
  OAI21_X1 U17144 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n13754), .A(n20065), 
        .ZN(n13755) );
  AND2_X1 U17145 ( .A1(n13756), .A2(n13755), .ZN(n19903) );
  NOR2_X2 U17146 ( .A1(n14369), .A2(n19915), .ZN(n20010) );
  NOR2_X2 U17147 ( .A1(n12030), .A2(n19583), .ZN(n20009) );
  AOI22_X1 U17148 ( .A1(n19903), .A2(n20010), .B1(n19902), .B2(n20009), .ZN(
        n13757) );
  OAI211_X1 U17149 ( .C1(n19908), .C2(n13759), .A(n13758), .B(n13757), .ZN(
        P2_U3137) );
  INV_X1 U17150 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13761) );
  AOI22_X1 U17151 ( .A1(n20907), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13760) );
  OAI21_X1 U17152 ( .B1(n13761), .B2(n13775), .A(n13760), .ZN(P1_U2917) );
  INV_X1 U17153 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13763) );
  AOI22_X1 U17154 ( .A1(n20907), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13762) );
  OAI21_X1 U17155 ( .B1(n13763), .B2(n13775), .A(n13762), .ZN(P1_U2919) );
  AOI22_X1 U17156 ( .A1(n20907), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13764) );
  OAI21_X1 U17157 ( .B1(n13765), .B2(n13775), .A(n13764), .ZN(P1_U2910) );
  INV_X1 U17158 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13767) );
  AOI22_X1 U17159 ( .A1(n20907), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13766) );
  OAI21_X1 U17160 ( .B1(n13767), .B2(n13775), .A(n13766), .ZN(P1_U2916) );
  INV_X1 U17161 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13769) );
  AOI22_X1 U17162 ( .A1(n20907), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13768) );
  OAI21_X1 U17163 ( .B1(n13769), .B2(n13775), .A(n13768), .ZN(P1_U2918) );
  INV_X1 U17164 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13771) );
  AOI22_X1 U17165 ( .A1(n20907), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13770) );
  OAI21_X1 U17166 ( .B1(n13771), .B2(n13775), .A(n13770), .ZN(P1_U2915) );
  INV_X1 U17167 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13773) );
  AOI22_X1 U17168 ( .A1(n20907), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13772) );
  OAI21_X1 U17169 ( .B1(n13773), .B2(n13775), .A(n13772), .ZN(P1_U2920) );
  INV_X1 U17170 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13776) );
  AOI22_X1 U17171 ( .A1(n20907), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13774) );
  OAI21_X1 U17172 ( .B1(n13776), .B2(n13775), .A(n13774), .ZN(P1_U2914) );
  XNOR2_X1 U17173 ( .A(n9665), .B(n13778), .ZN(n13788) );
  INV_X1 U17174 ( .A(n14227), .ZN(n13779) );
  OAI211_X1 U17175 ( .C1(n15101), .C2(n13779), .A(n15070), .B(n14228), .ZN(
        n13935) );
  NAND3_X1 U17176 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n15103), .ZN(n16266) );
  NAND2_X1 U17177 ( .A1(n15101), .A2(n16266), .ZN(n16232) );
  NAND2_X1 U17178 ( .A1(n13779), .A2(n16232), .ZN(n14232) );
  NAND2_X1 U17179 ( .A1(n14135), .A2(n16286), .ZN(n13780) );
  NAND2_X1 U17180 ( .A1(n16285), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n13784) );
  OAI211_X1 U17181 ( .C1(n14232), .C2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n13780), .B(n13784), .ZN(n13781) );
  AOI21_X1 U17182 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13935), .A(
        n13781), .ZN(n13782) );
  OAI21_X1 U17183 ( .B1(n16222), .B2(n13788), .A(n13782), .ZN(P1_U3028) );
  INV_X1 U17184 ( .A(n14137), .ZN(n13786) );
  NAND2_X1 U17185 ( .A1(n16173), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13783) );
  OAI211_X1 U17186 ( .C1(n16180), .C2(n14131), .A(n13784), .B(n13783), .ZN(
        n13785) );
  AOI21_X1 U17187 ( .B1(n13786), .B2(n14887), .A(n13785), .ZN(n13787) );
  OAI21_X1 U17188 ( .B1(n13788), .B2(n20226), .A(n13787), .ZN(P1_U2996) );
  AOI21_X1 U17189 ( .B1(n13790), .B2(n13643), .A(n11262), .ZN(n13933) );
  INV_X1 U17190 ( .A(n13933), .ZN(n20295) );
  AOI21_X1 U17191 ( .B1(n13792), .B2(n13791), .A(n14109), .ZN(n20298) );
  AOI22_X1 U17192 ( .A1(n20298), .A2(n20320), .B1(n14740), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n13793) );
  OAI21_X1 U17193 ( .B1(n20295), .B2(n14742), .A(n13793), .ZN(P1_U2868) );
  NAND3_X1 U17194 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11729), .A3(
        n11726), .ZN(n20572) );
  INV_X1 U17195 ( .A(n20572), .ZN(n13805) );
  INV_X1 U17196 ( .A(n20671), .ZN(n13796) );
  AND2_X1 U17197 ( .A1(n14132), .A2(n13496), .ZN(n20663) );
  INV_X1 U17198 ( .A(n13795), .ZN(n13906) );
  NOR2_X1 U17199 ( .A1(n14105), .A2(n20572), .ZN(n20605) );
  AOI21_X1 U17200 ( .B1(n20663), .B2(n13906), .A(n20605), .ZN(n13804) );
  OAI211_X1 U17201 ( .C1(n13796), .C2(n21095), .A(n20696), .B(n13804), .ZN(
        n13797) );
  OAI211_X1 U17202 ( .C1(n20696), .C2(n13805), .A(n13797), .B(n20748), .ZN(
        n20607) );
  INV_X1 U17203 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16734) );
  INV_X1 U17204 ( .A(n13871), .ZN(n13873) );
  INV_X1 U17205 ( .A(DATAI_16_), .ZN(n21029) );
  INV_X1 U17206 ( .A(n13870), .ZN(n13872) );
  OAI22_X1 U17207 ( .A1(n16734), .A2(n13873), .B1(n21029), .B2(n13872), .ZN(
        n20751) );
  INV_X1 U17208 ( .A(n20751), .ZN(n20612) );
  INV_X1 U17209 ( .A(n20754), .ZN(n20373) );
  NAND2_X1 U17210 ( .A1(n20606), .A2(n20373), .ZN(n13809) );
  NAND3_X1 U17211 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20222), .A3(n13801), 
        .ZN(n13827) );
  NAND2_X1 U17212 ( .A1(n13874), .A2(n13802), .ZN(n20611) );
  NOR2_X2 U17213 ( .A1(n13803), .A2(n14089), .ZN(n20744) );
  OR2_X1 U17214 ( .A1(n13804), .A2(n20743), .ZN(n13807) );
  NAND2_X1 U17215 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n13805), .ZN(n13806) );
  NAND2_X1 U17216 ( .A1(n13807), .A2(n13806), .ZN(n20604) );
  AOI22_X1 U17217 ( .A1(n20745), .A2(n20605), .B1(n20744), .B2(n20604), .ZN(
        n13808) );
  OAI211_X1 U17218 ( .C1(n20655), .C2(n20612), .A(n13809), .B(n13808), .ZN(
        n13810) );
  AOI21_X1 U17219 ( .B1(n20607), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n13810), .ZN(n13811) );
  INV_X1 U17220 ( .A(n13811), .ZN(P1_U3105) );
  INV_X1 U17221 ( .A(DATAI_19_), .ZN(n21014) );
  INV_X1 U17222 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16729) );
  OAI22_X1 U17223 ( .A1(n21014), .A2(n13872), .B1(n16729), .B2(n13873), .ZN(
        n20717) );
  INV_X1 U17224 ( .A(n20717), .ZN(n20772) );
  AOI22_X1 U17225 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n13871), .B1(DATAI_27_), 
        .B2(n13870), .ZN(n20720) );
  INV_X1 U17226 ( .A(n20720), .ZN(n20769) );
  NAND2_X1 U17227 ( .A1(n20606), .A2(n20769), .ZN(n13815) );
  NAND2_X1 U17228 ( .A1(n13874), .A2(n13812), .ZN(n20636) );
  NOR2_X2 U17229 ( .A1(n13813), .A2(n14089), .ZN(n20767) );
  AOI22_X1 U17230 ( .A1(n20768), .A2(n20605), .B1(n20767), .B2(n20604), .ZN(
        n13814) );
  OAI211_X1 U17231 ( .C1(n20655), .C2(n20772), .A(n13815), .B(n13814), .ZN(
        n13816) );
  AOI21_X1 U17232 ( .B1(n20607), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A(
        n13816), .ZN(n13817) );
  INV_X1 U17233 ( .A(n13817), .ZN(P1_U3108) );
  AOI22_X1 U17234 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n13871), .B1(DATAI_18_), 
        .B2(n13870), .ZN(n20635) );
  INV_X1 U17235 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16716) );
  INV_X1 U17236 ( .A(DATAI_26_), .ZN(n21008) );
  OAI22_X1 U17237 ( .A1(n16716), .A2(n13873), .B1(n21008), .B2(n13872), .ZN(
        n20497) );
  NAND2_X1 U17238 ( .A1(n20606), .A2(n20497), .ZN(n13820) );
  NAND2_X1 U17239 ( .A1(n13874), .A2(n11036), .ZN(n20631) );
  NOR2_X2 U17240 ( .A1(n13818), .A2(n14089), .ZN(n20761) );
  AOI22_X1 U17241 ( .A1(n20762), .A2(n20605), .B1(n20761), .B2(n20604), .ZN(
        n13819) );
  OAI211_X1 U17242 ( .C1(n20635), .C2(n20655), .A(n13820), .B(n13819), .ZN(
        n13821) );
  AOI21_X1 U17243 ( .B1(n20607), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n13821), .ZN(n13822) );
  INV_X1 U17244 ( .A(n13822), .ZN(P1_U3107) );
  INV_X1 U17245 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20348) );
  OAI222_X1 U17246 ( .A1(n20295), .A2(n14793), .B1(n14743), .B2(n20348), .C1(
        n14490), .C2(n13853), .ZN(P1_U2900) );
  AOI22_X1 U17247 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n13871), .B1(DATAI_21_), 
        .B2(n13870), .ZN(n20648) );
  INV_X1 U17248 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16710) );
  INV_X1 U17249 ( .A(DATAI_29_), .ZN(n20926) );
  OAI22_X1 U17250 ( .A1(n16710), .A2(n13873), .B1(n20926), .B2(n13872), .ZN(
        n20560) );
  NAND2_X1 U17251 ( .A1(n20606), .A2(n20560), .ZN(n13824) );
  NAND2_X1 U17252 ( .A1(n13874), .A2(n9710), .ZN(n20644) );
  NOR2_X2 U17253 ( .A1(n14112), .A2(n14089), .ZN(n20779) );
  AOI22_X1 U17254 ( .A1(n20780), .A2(n20605), .B1(n20779), .B2(n20604), .ZN(
        n13823) );
  OAI211_X1 U17255 ( .C1(n20648), .C2(n20655), .A(n13824), .B(n13823), .ZN(
        n13825) );
  AOI21_X1 U17256 ( .B1(n20607), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n13825), .ZN(n13826) );
  INV_X1 U17257 ( .A(n13826), .ZN(P1_U3110) );
  AOI22_X1 U17258 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n13871), .B1(DATAI_23_), 
        .B2(n13870), .ZN(n20693) );
  INV_X1 U17259 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16706) );
  INV_X1 U17260 ( .A(DATAI_31_), .ZN(n21049) );
  OAI22_X1 U17261 ( .A1(n16706), .A2(n13873), .B1(n21049), .B2(n13872), .ZN(
        n20688) );
  NAND2_X1 U17262 ( .A1(n20606), .A2(n20688), .ZN(n13829) );
  NOR2_X2 U17263 ( .A1(n14089), .A2(n14770), .ZN(n20796) );
  AOI22_X1 U17264 ( .A1(n20796), .A2(n20604), .B1(n20794), .B2(n20605), .ZN(
        n13828) );
  OAI211_X1 U17265 ( .C1(n20693), .C2(n20655), .A(n13829), .B(n13828), .ZN(
        n13830) );
  AOI21_X1 U17266 ( .B1(n20607), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n13830), .ZN(n13831) );
  INV_X1 U17267 ( .A(n13831), .ZN(P1_U3112) );
  NAND3_X1 U17268 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n10356), .ZN(n19911) );
  NOR2_X1 U17269 ( .A1(n20182), .A2(n19911), .ZN(n19964) );
  INV_X1 U17270 ( .A(n19964), .ZN(n13836) );
  OAI21_X1 U17271 ( .B1(n11964), .B2(n20065), .A(n19920), .ZN(n13835) );
  INV_X1 U17272 ( .A(n19696), .ZN(n13833) );
  INV_X1 U17273 ( .A(n19911), .ZN(n13832) );
  AOI21_X1 U17274 ( .B1(n19992), .B2(n13833), .A(n13832), .ZN(n13834) );
  INV_X1 U17275 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13840) );
  OR2_X1 U17276 ( .A1(n19818), .A2(n19696), .ZN(n15825) );
  AOI22_X1 U17277 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19588), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19587), .ZN(n19831) );
  NOR2_X2 U17278 ( .A1(n19786), .A2(n19696), .ZN(n19966) );
  AOI22_X1 U17279 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19588), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19587), .ZN(n19923) );
  INV_X1 U17280 ( .A(n19923), .ZN(n20004) );
  AOI22_X1 U17281 ( .A1(n19985), .A2(n20005), .B1(n19966), .B2(n20004), .ZN(
        n13839) );
  OAI21_X1 U17282 ( .B1(n11964), .B2(n19964), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13837) );
  OAI21_X1 U17283 ( .B1(n19911), .B2(n20150), .A(n13837), .ZN(n19965) );
  NOR2_X2 U17284 ( .A1(n14305), .A2(n19915), .ZN(n20003) );
  INV_X1 U17285 ( .A(n19583), .ZN(n14160) );
  NAND2_X1 U17286 ( .A1(n16615), .A2(n14160), .ZN(n14180) );
  AOI22_X1 U17287 ( .A1(n19965), .A2(n20003), .B1(n20002), .B2(n19964), .ZN(
        n13838) );
  OAI211_X1 U17288 ( .C1(n19970), .C2(n13840), .A(n13839), .B(n13838), .ZN(
        P2_U3152) );
  INV_X1 U17289 ( .A(n9716), .ZN(n13842) );
  NAND4_X1 U17290 ( .A1(n20747), .A2(n13843), .A3(n13842), .A4(n20700), .ZN(
        n15114) );
  NAND3_X1 U17291 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n11726), .ZN(n20694) );
  INV_X1 U17292 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13848) );
  NOR2_X1 U17293 ( .A1(n14105), .A2(n20694), .ZN(n13881) );
  INV_X1 U17294 ( .A(n13881), .ZN(n13844) );
  INV_X1 U17295 ( .A(n13905), .ZN(n14078) );
  OR2_X1 U17296 ( .A1(n13496), .A2(n14078), .ZN(n14238) );
  NOR2_X1 U17297 ( .A1(n14238), .A2(n20743), .ZN(n14242) );
  INV_X1 U17298 ( .A(n14242), .ZN(n20740) );
  OAI222_X1 U17299 ( .A1(n13844), .A2(n20743), .B1(n20806), .B2(n20694), .C1(
        n13795), .C2(n20740), .ZN(n13880) );
  AOI22_X1 U17300 ( .A1(n20768), .A2(n13881), .B1(n13880), .B2(n20767), .ZN(
        n13845) );
  OAI21_X1 U17301 ( .B1(n13883), .B2(n20720), .A(n13845), .ZN(n13846) );
  AOI21_X1 U17302 ( .B1(n15130), .B2(n20717), .A(n13846), .ZN(n13847) );
  OAI21_X1 U17303 ( .B1(n13887), .B2(n13848), .A(n13847), .ZN(P1_U3140) );
  INV_X1 U17304 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13852) );
  INV_X1 U17305 ( .A(DATAI_22_), .ZN(n21043) );
  INV_X1 U17306 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16724) );
  OAI22_X1 U17307 ( .A1(n21043), .A2(n13872), .B1(n16724), .B2(n13873), .ZN(
        n20727) );
  AOI22_X1 U17308 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n13871), .B1(DATAI_30_), 
        .B2(n13870), .ZN(n20730) );
  NAND2_X1 U17309 ( .A1(n13874), .A2(n11001), .ZN(n20649) );
  NOR2_X2 U17310 ( .A1(n14140), .A2(n14089), .ZN(n20785) );
  AOI22_X1 U17311 ( .A1(n20786), .A2(n13881), .B1(n13880), .B2(n20785), .ZN(
        n13849) );
  OAI21_X1 U17312 ( .B1(n13883), .B2(n20730), .A(n13849), .ZN(n13850) );
  AOI21_X1 U17313 ( .B1(n15130), .B2(n20727), .A(n13850), .ZN(n13851) );
  OAI21_X1 U17314 ( .B1(n13887), .B2(n13852), .A(n13851), .ZN(P1_U3143) );
  INV_X1 U17315 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13857) );
  AOI22_X1 U17316 ( .A1(DATAI_20_), .A2(n13870), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n13871), .ZN(n20778) );
  INV_X1 U17317 ( .A(n20778), .ZN(n20721) );
  INV_X1 U17318 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16712) );
  INV_X1 U17319 ( .A(DATAI_28_), .ZN(n21097) );
  OAI22_X1 U17320 ( .A1(n16712), .A2(n13873), .B1(n21097), .B2(n13872), .ZN(
        n20775) );
  NAND2_X1 U17321 ( .A1(n13874), .A2(n11033), .ZN(n20640) );
  NOR2_X2 U17322 ( .A1(n13853), .A2(n14089), .ZN(n20773) );
  AOI22_X1 U17323 ( .A1(n20774), .A2(n13881), .B1(n13880), .B2(n20773), .ZN(
        n13854) );
  OAI21_X1 U17324 ( .B1(n13883), .B2(n20724), .A(n13854), .ZN(n13855) );
  AOI21_X1 U17325 ( .B1(n15130), .B2(n20721), .A(n13855), .ZN(n13856) );
  OAI21_X1 U17326 ( .B1(n13887), .B2(n13857), .A(n13856), .ZN(P1_U3141) );
  INV_X1 U17327 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13861) );
  INV_X1 U17328 ( .A(n20648), .ZN(n20781) );
  INV_X1 U17329 ( .A(n20560), .ZN(n20784) );
  AOI22_X1 U17330 ( .A1(n20780), .A2(n13881), .B1(n13880), .B2(n20779), .ZN(
        n13858) );
  OAI21_X1 U17331 ( .B1(n13883), .B2(n20784), .A(n13858), .ZN(n13859) );
  AOI21_X1 U17332 ( .B1(n15130), .B2(n20781), .A(n13859), .ZN(n13860) );
  OAI21_X1 U17333 ( .B1(n13887), .B2(n13861), .A(n13860), .ZN(P1_U3142) );
  INV_X1 U17334 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13865) );
  INV_X1 U17335 ( .A(n20693), .ZN(n20797) );
  INV_X1 U17336 ( .A(n20688), .ZN(n20803) );
  AOI22_X1 U17337 ( .A1(n13880), .A2(n20796), .B1(n20794), .B2(n13881), .ZN(
        n13862) );
  OAI21_X1 U17338 ( .B1(n13883), .B2(n20803), .A(n13862), .ZN(n13863) );
  AOI21_X1 U17339 ( .B1(n15130), .B2(n20797), .A(n13863), .ZN(n13864) );
  OAI21_X1 U17340 ( .B1(n13887), .B2(n13865), .A(n13864), .ZN(P1_U3144) );
  INV_X1 U17341 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13869) );
  INV_X1 U17342 ( .A(n20635), .ZN(n20763) );
  AOI22_X1 U17343 ( .A1(n20762), .A2(n13881), .B1(n13880), .B2(n20761), .ZN(
        n13866) );
  OAI21_X1 U17344 ( .B1(n13883), .B2(n20766), .A(n13866), .ZN(n13867) );
  AOI21_X1 U17345 ( .B1(n15130), .B2(n20763), .A(n13867), .ZN(n13868) );
  OAI21_X1 U17346 ( .B1(n13887), .B2(n13869), .A(n13868), .ZN(P1_U3139) );
  INV_X1 U17347 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13879) );
  AOI22_X1 U17348 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n13871), .B1(DATAI_17_), 
        .B2(n13870), .ZN(n20760) );
  INV_X1 U17349 ( .A(n20760), .ZN(n20711) );
  INV_X1 U17350 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16718) );
  INV_X1 U17351 ( .A(DATAI_25_), .ZN(n21091) );
  OAI22_X1 U17352 ( .A1(n16718), .A2(n13873), .B1(n21091), .B2(n13872), .ZN(
        n20757) );
  INV_X1 U17353 ( .A(n20757), .ZN(n20714) );
  NAND2_X1 U17354 ( .A1(n13874), .A2(n13992), .ZN(n20627) );
  NOR2_X2 U17355 ( .A1(n13875), .A2(n14089), .ZN(n20755) );
  AOI22_X1 U17356 ( .A1(n20756), .A2(n13881), .B1(n13880), .B2(n20755), .ZN(
        n13876) );
  OAI21_X1 U17357 ( .B1(n13883), .B2(n20714), .A(n13876), .ZN(n13877) );
  AOI21_X1 U17358 ( .B1(n15130), .B2(n20711), .A(n13877), .ZN(n13878) );
  OAI21_X1 U17359 ( .B1(n13887), .B2(n13879), .A(n13878), .ZN(P1_U3138) );
  INV_X1 U17360 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13886) );
  AOI22_X1 U17361 ( .A1(n20745), .A2(n13881), .B1(n13880), .B2(n20744), .ZN(
        n13882) );
  OAI21_X1 U17362 ( .B1(n13883), .B2(n20754), .A(n13882), .ZN(n13884) );
  AOI21_X1 U17363 ( .B1(n20751), .B2(n15130), .A(n13884), .ZN(n13885) );
  OAI21_X1 U17364 ( .B1(n13887), .B2(n13886), .A(n13885), .ZN(P1_U3137) );
  NAND3_X1 U17365 ( .A1(n20661), .A2(n11729), .A3(n11726), .ZN(n14310) );
  INV_X1 U17366 ( .A(n14310), .ZN(n13891) );
  INV_X1 U17367 ( .A(n20413), .ZN(n20449) );
  INV_X1 U17368 ( .A(n13496), .ZN(n13888) );
  OR2_X1 U17369 ( .A1(n14132), .A2(n13888), .ZN(n14313) );
  INV_X1 U17370 ( .A(n14313), .ZN(n20452) );
  NOR2_X1 U17371 ( .A1(n14105), .A2(n14310), .ZN(n20407) );
  AOI21_X1 U17372 ( .B1(n20452), .B2(n13906), .A(n20407), .ZN(n13890) );
  OAI211_X1 U17373 ( .C1(n20449), .C2(n21095), .A(n20696), .B(n13890), .ZN(
        n13889) );
  NAND2_X1 U17374 ( .A1(n20410), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13895) );
  INV_X1 U17375 ( .A(n13890), .ZN(n13892) );
  AOI22_X1 U17376 ( .A1(n13892), .A2(n20696), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13891), .ZN(n20398) );
  INV_X1 U17377 ( .A(n20744), .ZN(n14255) );
  INV_X1 U17378 ( .A(n20407), .ZN(n13899) );
  OAI22_X1 U17379 ( .A1(n20398), .A2(n14255), .B1(n20611), .B2(n13899), .ZN(
        n13893) );
  AOI21_X1 U17380 ( .B1(n20409), .B2(n20373), .A(n13893), .ZN(n13894) );
  OAI211_X1 U17381 ( .C1(n20442), .C2(n20612), .A(n13895), .B(n13894), .ZN(
        P1_U3041) );
  NAND2_X1 U17382 ( .A1(n20410), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n13898) );
  INV_X1 U17383 ( .A(n20773), .ZN(n14247) );
  OAI22_X1 U17384 ( .A1(n20398), .A2(n14247), .B1(n20640), .B2(n13899), .ZN(
        n13896) );
  AOI21_X1 U17385 ( .B1(n20775), .B2(n20409), .A(n13896), .ZN(n13897) );
  OAI211_X1 U17386 ( .C1(n20778), .C2(n20442), .A(n13898), .B(n13897), .ZN(
        P1_U3045) );
  NAND2_X1 U17387 ( .A1(n20410), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13902) );
  INV_X1 U17388 ( .A(n20755), .ZN(n14251) );
  OAI22_X1 U17389 ( .A1(n20398), .A2(n14251), .B1(n20627), .B2(n13899), .ZN(
        n13900) );
  AOI21_X1 U17390 ( .B1(n20757), .B2(n20409), .A(n13900), .ZN(n13901) );
  OAI211_X1 U17391 ( .C1(n20760), .C2(n20442), .A(n13902), .B(n13901), .ZN(
        P1_U3042) );
  NAND2_X1 U17392 ( .A1(n20549), .A2(n10175), .ZN(n14199) );
  INV_X1 U17393 ( .A(n20796), .ZN(n14210) );
  NOR2_X1 U17394 ( .A1(n13496), .A2(n13905), .ZN(n20543) );
  NAND3_X1 U17395 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20661), .A3(
        n11726), .ZN(n14202) );
  NOR2_X1 U17396 ( .A1(n14105), .A2(n14202), .ZN(n20506) );
  AOI21_X1 U17397 ( .B1(n20543), .B2(n13906), .A(n20506), .ZN(n13909) );
  INV_X1 U17398 ( .A(n13909), .ZN(n13907) );
  INV_X1 U17399 ( .A(n14202), .ZN(n13913) );
  AOI22_X1 U17400 ( .A1(n13907), .A2(n20696), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13913), .ZN(n20496) );
  INV_X1 U17401 ( .A(n20794), .ZN(n20654) );
  INV_X1 U17402 ( .A(n20506), .ZN(n13919) );
  OAI22_X1 U17403 ( .A1(n14210), .A2(n20496), .B1(n20654), .B2(n13919), .ZN(
        n13908) );
  AOI21_X1 U17404 ( .B1(n20688), .B2(n20508), .A(n13908), .ZN(n13915) );
  INV_X1 U17405 ( .A(n20549), .ZN(n13911) );
  NAND2_X1 U17406 ( .A1(n20696), .A2(n21095), .ZN(n20614) );
  INV_X1 U17407 ( .A(n20614), .ZN(n13910) );
  OAI21_X1 U17408 ( .B1(n13911), .B2(n13910), .A(n13909), .ZN(n13912) );
  OAI211_X1 U17409 ( .C1(n20696), .C2(n13913), .A(n13912), .B(n20748), .ZN(
        n20509) );
  NAND2_X1 U17410 ( .A1(n20509), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n13914) );
  OAI211_X1 U17411 ( .C1(n20693), .C2(n20531), .A(n13915), .B(n13914), .ZN(
        P1_U3080) );
  NAND2_X1 U17412 ( .A1(n20509), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n13918) );
  OAI22_X1 U17413 ( .A1(n20496), .A2(n14255), .B1(n20611), .B2(n13919), .ZN(
        n13916) );
  AOI21_X1 U17414 ( .B1(n20508), .B2(n20373), .A(n13916), .ZN(n13917) );
  OAI211_X1 U17415 ( .C1(n20531), .C2(n20612), .A(n13918), .B(n13917), .ZN(
        P1_U3073) );
  NAND2_X1 U17416 ( .A1(n20509), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13922) );
  OAI22_X1 U17417 ( .A1(n20496), .A2(n14251), .B1(n20627), .B2(n13919), .ZN(
        n13920) );
  AOI21_X1 U17418 ( .B1(n20757), .B2(n20508), .A(n13920), .ZN(n13921) );
  OAI211_X1 U17419 ( .C1(n20760), .C2(n20531), .A(n13922), .B(n13921), .ZN(
        P1_U3074) );
  XOR2_X1 U17420 ( .A(n13923), .B(n14013), .Z(n13927) );
  NOR2_X1 U17421 ( .A1(n19406), .A2(n13924), .ZN(n13925) );
  AOI21_X1 U17422 ( .B1(n16549), .B2(n19406), .A(n13925), .ZN(n13926) );
  OAI21_X1 U17423 ( .B1(n13927), .B2(n19403), .A(n13926), .ZN(P2_U2876) );
  XNOR2_X1 U17424 ( .A(n13929), .B(n13928), .ZN(n13942) );
  INV_X1 U17425 ( .A(n13930), .ZN(n20293) );
  NAND2_X1 U17426 ( .A1(n16285), .A2(P1_REIP_REG_4__SCAN_IN), .ZN(n13937) );
  NAND2_X1 U17427 ( .A1(n16173), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13931) );
  OAI211_X1 U17428 ( .C1(n16180), .C2(n20293), .A(n13937), .B(n13931), .ZN(
        n13932) );
  AOI21_X1 U17429 ( .B1(n13933), .B2(n14887), .A(n13932), .ZN(n13934) );
  OAI21_X1 U17430 ( .B1(n20226), .B2(n13942), .A(n13934), .ZN(P1_U2995) );
  NAND2_X1 U17431 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13935), .ZN(
        n13936) );
  NAND2_X1 U17432 ( .A1(n13937), .A2(n13936), .ZN(n13940) );
  NOR2_X1 U17433 ( .A1(n13938), .A2(n12355), .ZN(n14410) );
  AOI211_X1 U17434 ( .C1(n13938), .C2(n12355), .A(n14410), .B(n14232), .ZN(
        n13939) );
  AOI211_X1 U17435 ( .C1(n16286), .C2(n20298), .A(n13940), .B(n13939), .ZN(
        n13941) );
  OAI21_X1 U17436 ( .B1(n16222), .B2(n13942), .A(n13941), .ZN(P1_U3027) );
  INV_X1 U17437 ( .A(n20153), .ZN(n13944) );
  AOI21_X1 U17438 ( .B1(n15819), .B2(n13944), .A(n13943), .ZN(n13947) );
  XOR2_X1 U17439 ( .A(n13945), .B(n13946), .Z(n19524) );
  NOR2_X1 U17440 ( .A1(n13947), .A2(n19524), .ZN(n14052) );
  INV_X1 U17441 ( .A(n13948), .ZN(n13949) );
  NAND2_X1 U17442 ( .A1(n13545), .A2(n13951), .ZN(n19367) );
  XNOR2_X1 U17443 ( .A(n14052), .B(n19367), .ZN(n13955) );
  AOI22_X1 U17444 ( .A1(n19434), .A2(n13952), .B1(n19432), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n13954) );
  NAND2_X1 U17445 ( .A1(n19524), .A2(n19417), .ZN(n13953) );
  OAI211_X1 U17446 ( .C1(n13955), .C2(n15373), .A(n13954), .B(n13953), .ZN(
        P2_U2915) );
  NAND2_X1 U17447 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20156), .ZN(
        n19754) );
  NOR3_X2 U17448 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19754), .ZN(n19689) );
  NOR2_X1 U17449 ( .A1(n20157), .A2(n19689), .ZN(n13956) );
  OAI21_X1 U17450 ( .B1(n12039), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n13956), 
        .ZN(n13961) );
  NOR2_X1 U17451 ( .A1(n13957), .A2(n14173), .ZN(n19909) );
  NAND2_X1 U17452 ( .A1(n19909), .A2(n20156), .ZN(n13964) );
  OAI21_X1 U17453 ( .B1(n19691), .B2(n19713), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13958) );
  AND2_X1 U17454 ( .A1(n13964), .A2(n13958), .ZN(n13959) );
  NOR2_X1 U17455 ( .A1(n19915), .A2(n13959), .ZN(n13960) );
  NAND2_X1 U17456 ( .A1(n13961), .A2(n13960), .ZN(n19692) );
  INV_X1 U17457 ( .A(n19692), .ZN(n19679) );
  INV_X1 U17458 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13970) );
  OAI21_X1 U17459 ( .B1(n13962), .B2(n19689), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13963) );
  OAI21_X1 U17460 ( .B1(n13964), .B2(n20150), .A(n13963), .ZN(n19690) );
  INV_X1 U17461 ( .A(n20009), .ZN(n13967) );
  INV_X1 U17462 ( .A(n19689), .ZN(n13966) );
  AOI22_X1 U17463 ( .A1(n19691), .A2(n20012), .B1(n19713), .B2(n20011), .ZN(
        n13965) );
  OAI21_X1 U17464 ( .B1(n13967), .B2(n13966), .A(n13965), .ZN(n13968) );
  AOI21_X1 U17465 ( .B1(n19690), .B2(n20010), .A(n13968), .ZN(n13969) );
  OAI21_X1 U17466 ( .B1(n19679), .B2(n13970), .A(n13969), .ZN(P2_U3081) );
  XNOR2_X1 U17467 ( .A(n13971), .B(n14141), .ZN(n13978) );
  OR2_X1 U17468 ( .A1(n13972), .A2(n13973), .ZN(n13975) );
  NOR2_X1 U17469 ( .A1(n19406), .A2(n10790), .ZN(n13976) );
  AOI21_X1 U17470 ( .B1(n19306), .B2(n19406), .A(n13976), .ZN(n13977) );
  OAI21_X1 U17471 ( .B1(n13978), .B2(n19403), .A(n13977), .ZN(P2_U2874) );
  NOR2_X1 U17472 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20911) );
  NAND2_X1 U17473 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20911), .ZN(n16300) );
  AND2_X1 U17474 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20222), .ZN(n13979) );
  NAND2_X1 U17475 ( .A1(n13980), .A2(n13979), .ZN(n13981) );
  OAI21_X1 U17476 ( .B1(n16300), .B2(n20222), .A(n13981), .ZN(n13982) );
  OR2_X1 U17477 ( .A1(n13990), .A2(n13984), .ZN(n20312) );
  INV_X1 U17478 ( .A(n11172), .ZN(n14102) );
  NOR2_X1 U17479 ( .A1(n14001), .A2(n13985), .ZN(n13986) );
  OAI21_X1 U17480 ( .B1(n13987), .B2(n13990), .A(n16093), .ZN(n20314) );
  NAND2_X1 U17481 ( .A1(n13988), .A2(n20314), .ZN(n14008) );
  NOR2_X1 U17482 ( .A1(n13991), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13998) );
  NAND2_X1 U17483 ( .A1(n20259), .A2(n16082), .ZN(n16083) );
  NAND2_X1 U17484 ( .A1(n16083), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n14006) );
  NAND2_X1 U17485 ( .A1(n13992), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13996) );
  AND2_X1 U17486 ( .A1(n20906), .A2(n21095), .ZN(n13993) );
  NOR2_X1 U17487 ( .A1(n13996), .A2(n13993), .ZN(n13994) );
  NAND2_X1 U17488 ( .A1(n20303), .A2(n13995), .ZN(n14005) );
  INV_X1 U17489 ( .A(n13996), .ZN(n13997) );
  NOR2_X1 U17490 ( .A1(n13998), .A2(n13997), .ZN(n13999) );
  NAND2_X1 U17491 ( .A1(n20304), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n14004) );
  AND2_X1 U17492 ( .A1(n14001), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14002) );
  OAI21_X1 U17493 ( .B1(n20306), .B2(n20307), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14003) );
  AND4_X1 U17494 ( .A1(n14006), .A2(n14005), .A3(n14004), .A4(n14003), .ZN(
        n14007) );
  OAI211_X1 U17495 ( .C1(n20312), .C2(n14102), .A(n14008), .B(n14007), .ZN(
        P1_U2840) );
  INV_X1 U17496 ( .A(n14009), .ZN(n14012) );
  INV_X1 U17497 ( .A(n14010), .ZN(n14011) );
  AOI21_X1 U17498 ( .B1(n14012), .B2(n14011), .A(n13972), .ZN(n19316) );
  INV_X1 U17499 ( .A(n19316), .ZN(n14020) );
  INV_X1 U17500 ( .A(n14013), .ZN(n14014) );
  NOR2_X1 U17501 ( .A1(n13923), .A2(n14014), .ZN(n14017) );
  INV_X1 U17502 ( .A(n13971), .ZN(n14015) );
  OAI211_X1 U17503 ( .C1(n14017), .C2(n14016), .A(n14015), .B(n19411), .ZN(
        n14019) );
  NAND2_X1 U17504 ( .A1(n16392), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14018) );
  OAI211_X1 U17505 ( .C1(n14020), .C2(n16392), .A(n14019), .B(n14018), .ZN(
        P2_U2875) );
  NAND2_X1 U17506 ( .A1(n14022), .A2(n9702), .ZN(n14024) );
  XNOR2_X1 U17507 ( .A(n14024), .B(n14023), .ZN(n14041) );
  XOR2_X1 U17508 ( .A(n12280), .B(n14025), .Z(n14039) );
  NOR2_X1 U17509 ( .A1(n14034), .A2(n19324), .ZN(n14026) );
  AOI221_X1 U17510 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14029), .C1(
        n14028), .C2(n14027), .A(n14026), .ZN(n14031) );
  NAND2_X1 U17511 ( .A1(n19537), .A2(n20153), .ZN(n14030) );
  OAI211_X1 U17512 ( .C1(n19540), .C2(n13472), .A(n14031), .B(n14030), .ZN(
        n14032) );
  AOI21_X1 U17513 ( .B1(n16577), .B2(n14039), .A(n14032), .ZN(n14033) );
  OAI21_X1 U17514 ( .B1(n14041), .B2(n16589), .A(n14033), .ZN(P2_U3043) );
  OAI22_X1 U17515 ( .A1(n16506), .A2(n14035), .B1(n14034), .B2(n19324), .ZN(
        n14036) );
  AOI21_X1 U17516 ( .B1(n16494), .B2(n15206), .A(n14036), .ZN(n14037) );
  OAI21_X1 U17517 ( .B1(n13472), .B2(n16436), .A(n14037), .ZN(n14038) );
  AOI21_X1 U17518 ( .B1(n14039), .B2(n19507), .A(n14038), .ZN(n14040) );
  OAI21_X1 U17519 ( .B1(n14041), .B2(n19510), .A(n14040), .ZN(P2_U3011) );
  AOI21_X1 U17520 ( .B1(n14042), .B2(n15692), .A(n9740), .ZN(n19283) );
  INV_X1 U17521 ( .A(n19283), .ZN(n14045) );
  OAI222_X1 U17522 ( .A1(n14046), .A2(n19428), .B1(n14045), .B2(n19437), .C1(
        n14044), .C2(n14043), .ZN(P2_U2904) );
  INV_X1 U17523 ( .A(n14047), .ZN(n14048) );
  NAND2_X1 U17524 ( .A1(n14049), .A2(n14048), .ZN(n14050) );
  AND2_X1 U17525 ( .A1(n14051), .A2(n14050), .ZN(n16572) );
  INV_X1 U17526 ( .A(n16572), .ZN(n14056) );
  OR3_X1 U17527 ( .A1(n14052), .A2(n15373), .A3(n19367), .ZN(n14055) );
  AOI22_X1 U17528 ( .A1(n19434), .A2(n14053), .B1(n19432), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n14054) );
  OAI211_X1 U17529 ( .C1(n19437), .C2(n14056), .A(n14055), .B(n14054), .ZN(
        P2_U2914) );
  NOR2_X1 U17530 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13985), .ZN(n14084) );
  MUX2_X1 U17531 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14057), .S(
        n15979), .Z(n15985) );
  AOI22_X1 U17532 ( .A1(n14084), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15985), .B2(n13985), .ZN(n14077) );
  INV_X1 U17533 ( .A(n14061), .ZN(n14058) );
  OAI211_X1 U17534 ( .C1(n13508), .C2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n14059), .B(n14058), .ZN(n20885) );
  OR3_X1 U17535 ( .A1(n15976), .A2(n14060), .A3(n20885), .ZN(n14072) );
  MUX2_X1 U17536 ( .A(n14061), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n13508), .Z(n14063) );
  NOR2_X1 U17537 ( .A1(n14063), .A2(n14062), .ZN(n14069) );
  INV_X1 U17538 ( .A(n14064), .ZN(n14067) );
  NAND2_X1 U17539 ( .A1(n14065), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14066) );
  NAND2_X1 U17540 ( .A1(n14067), .A2(n14066), .ZN(n14068) );
  AOI22_X1 U17541 ( .A1(n14070), .A2(n14069), .B1(n15977), .B2(n14068), .ZN(
        n14071) );
  OAI211_X1 U17542 ( .C1(n14074), .C2(n15117), .A(n14072), .B(n14071), .ZN(
        n14073) );
  AOI21_X1 U17543 ( .B1(n14132), .B2(n15976), .A(n14073), .ZN(n20886) );
  MUX2_X1 U17544 ( .A(n14074), .B(n20886), .S(n15979), .Z(n15986) );
  INV_X1 U17545 ( .A(n15986), .ZN(n14075) );
  AOI22_X1 U17546 ( .A1(n14075), .A2(n13985), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n14084), .ZN(n14076) );
  OR2_X1 U17547 ( .A1(n14079), .A2(n14078), .ZN(n14080) );
  INV_X1 U17548 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16296) );
  XNOR2_X1 U17549 ( .A(n14080), .B(n16296), .ZN(n20284) );
  OAI21_X1 U17550 ( .B1(n20284), .B2(n13506), .A(n15979), .ZN(n14083) );
  INV_X1 U17551 ( .A(n15979), .ZN(n14081) );
  NAND2_X1 U17552 ( .A1(n14081), .A2(n16296), .ZN(n14082) );
  NAND3_X1 U17553 ( .A1(n14083), .A2(n13985), .A3(n14082), .ZN(n14086) );
  NAND2_X1 U17554 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n14084), .ZN(
        n14085) );
  NAND2_X1 U17555 ( .A1(n14086), .A2(n14085), .ZN(n15995) );
  INV_X1 U17556 ( .A(n15995), .ZN(n14087) );
  NOR2_X1 U17557 ( .A1(n20222), .A2(n16304), .ZN(n14088) );
  OAI21_X1 U17558 ( .B1(n14101), .B2(P1_FLUSH_REG_SCAN_IN), .A(n14088), .ZN(
        n14090) );
  NAND2_X1 U17559 ( .A1(n14090), .A2(n14089), .ZN(n20372) );
  AND2_X1 U17560 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20700), .ZN(n15110) );
  OR2_X1 U17561 ( .A1(n9716), .A2(n20743), .ZN(n14092) );
  NAND2_X1 U17562 ( .A1(n14092), .A2(n20614), .ZN(n20666) );
  OAI21_X1 U17563 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n9716), .A(n20666), 
        .ZN(n14093) );
  OAI21_X1 U17564 ( .B1(n15110), .B2(n20698), .A(n14093), .ZN(n14094) );
  NAND2_X1 U17565 ( .A1(n20372), .A2(n14094), .ZN(n14095) );
  OAI21_X1 U17566 ( .B1(n20372), .B2(n11726), .A(n14095), .ZN(P1_U3477) );
  NOR2_X1 U17567 ( .A1(n13496), .A2(n15110), .ZN(n14099) );
  AND2_X1 U17568 ( .A1(n20696), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14096) );
  AND2_X1 U17569 ( .A1(n9716), .A2(n14096), .ZN(n20746) );
  MUX2_X1 U17570 ( .A(n20746), .B(n20666), .S(n14097), .Z(n14098) );
  OAI21_X1 U17571 ( .B1(n14099), .B2(n14098), .A(n20372), .ZN(n14100) );
  OAI21_X1 U17572 ( .B1(n11729), .B2(n20372), .A(n14100), .ZN(P1_U3476) );
  NOR2_X1 U17573 ( .A1(n14101), .A2(n16304), .ZN(n16006) );
  OAI22_X1 U17574 ( .A1(n9669), .A2(n20743), .B1(n14102), .B2(n15110), .ZN(
        n14103) );
  OAI21_X1 U17575 ( .B1(n16006), .B2(n14103), .A(n20372), .ZN(n14104) );
  OAI21_X1 U17576 ( .B1(n20372), .B2(n14105), .A(n14104), .ZN(P1_U3478) );
  AOI21_X1 U17577 ( .B1(n14107), .B2(n13789), .A(n11293), .ZN(n20280) );
  INV_X1 U17578 ( .A(n20280), .ZN(n14113) );
  NOR2_X1 U17579 ( .A1(n14109), .A2(n14108), .ZN(n14110) );
  OR2_X1 U17580 ( .A1(n16282), .A2(n14110), .ZN(n20273) );
  OAI222_X1 U17581 ( .A1(n14113), .A2(n14742), .B1(n20324), .B2(n14111), .C1(
        n14737), .C2(n20273), .ZN(P1_U2867) );
  OAI222_X1 U17582 ( .A1(n14113), .A2(n14793), .B1(n14490), .B2(n14112), .C1(
        n14743), .C2(n11259), .ZN(P1_U2899) );
  NOR2_X1 U17583 ( .A1(n19372), .A2(n14114), .ZN(n14115) );
  XNOR2_X1 U17584 ( .A(n14115), .B(n14346), .ZN(n14116) );
  NAND2_X1 U17585 ( .A1(n14116), .A2(n19342), .ZN(n14124) );
  INV_X1 U17586 ( .A(n14357), .ZN(n14122) );
  INV_X1 U17587 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20096) );
  OAI21_X1 U17588 ( .B1(n20096), .B2(n19387), .A(n19324), .ZN(n14117) );
  AOI21_X1 U17589 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19360), .A(
        n14117), .ZN(n14119) );
  NAND2_X1 U17590 ( .A1(n19361), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n14118) );
  OAI211_X1 U17591 ( .C1(n14120), .C2(n19362), .A(n14119), .B(n14118), .ZN(
        n14121) );
  AOI21_X1 U17592 ( .B1(n14122), .B2(n19305), .A(n14121), .ZN(n14123) );
  OAI211_X1 U17593 ( .C1(n14353), .C2(n19354), .A(n14124), .B(n14123), .ZN(
        P2_U2849) );
  INV_X1 U17594 ( .A(n20314), .ZN(n20294) );
  NAND2_X1 U17595 ( .A1(n20304), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n14130) );
  NAND3_X1 U17596 ( .A1(n20309), .A2(P1_REIP_REG_1__SCAN_IN), .A3(
        P1_REIP_REG_2__SCAN_IN), .ZN(n14127) );
  OAI221_X1 U17597 ( .B1(n20259), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n20259), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n16082), .ZN(n14125) );
  NAND2_X1 U17598 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n14125), .ZN(n14126) );
  OAI21_X1 U17599 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(n14127), .A(n14126), .ZN(
        n14128) );
  AOI21_X1 U17600 ( .B1(n20306), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n14128), .ZN(n14129) );
  OAI211_X1 U17601 ( .C1(n20292), .C2(n14131), .A(n14130), .B(n14129), .ZN(
        n14134) );
  INV_X1 U17602 ( .A(n14132), .ZN(n15111) );
  NOR2_X1 U17603 ( .A1(n15111), .A2(n20312), .ZN(n14133) );
  AOI211_X1 U17604 ( .C1(n14135), .C2(n20303), .A(n14134), .B(n14133), .ZN(
        n14136) );
  OAI21_X1 U17605 ( .B1(n14137), .B2(n20294), .A(n14136), .ZN(P1_U2837) );
  XNOR2_X1 U17606 ( .A(n14106), .B(n14152), .ZN(n20321) );
  INV_X1 U17607 ( .A(n20321), .ZN(n14139) );
  INV_X1 U17608 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n14138) );
  OAI222_X1 U17609 ( .A1(n14490), .A2(n14140), .B1(n14793), .B2(n14139), .C1(
        n14138), .C2(n14743), .ZN(P1_U2898) );
  AND2_X1 U17610 ( .A1(n13971), .A2(n14141), .ZN(n14144) );
  OAI211_X1 U17611 ( .C1(n14144), .C2(n14143), .A(n19411), .B(n14142), .ZN(
        n14149) );
  NAND2_X1 U17612 ( .A1(n14145), .A2(n13974), .ZN(n14147) );
  INV_X1 U17613 ( .A(n14294), .ZN(n14146) );
  NAND2_X1 U17614 ( .A1(n19415), .A2(n19294), .ZN(n14148) );
  OAI211_X1 U17615 ( .C1(n19406), .C2(n14150), .A(n14149), .B(n14148), .ZN(
        P2_U2873) );
  AOI21_X1 U17616 ( .B1(n11293), .B2(n14152), .A(n14151), .ZN(n14154) );
  OR2_X1 U17617 ( .A1(n14154), .A2(n14153), .ZN(n16170) );
  XNOR2_X1 U17618 ( .A(n14279), .B(n14281), .ZN(n20251) );
  INV_X1 U17619 ( .A(n20251), .ZN(n14156) );
  OAI222_X1 U17620 ( .A1(n16170), .A2(n14742), .B1(n14737), .B2(n14156), .C1(
        n14155), .C2(n20324), .ZN(P1_U2865) );
  INV_X1 U17621 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n20344) );
  OAI222_X1 U17622 ( .A1(n16170), .A2(n14793), .B1(n14490), .B2(n14770), .C1(
        n14743), .C2(n20344), .ZN(P1_U2897) );
  NOR3_X1 U17623 ( .A1(n20055), .A2(n19985), .A3(n20150), .ZN(n14157) );
  NOR2_X1 U17624 ( .A1(n20150), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20147) );
  NOR2_X1 U17625 ( .A1(n14157), .A2(n20147), .ZN(n14167) );
  INV_X1 U17626 ( .A(n14167), .ZN(n14159) );
  NOR3_X2 U17627 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20156), .A3(
        n19991), .ZN(n19984) );
  NOR2_X1 U17628 ( .A1(n19984), .A2(n19964), .ZN(n14166) );
  AOI211_X1 U17629 ( .C1(n14164), .C2(n19920), .A(n20157), .B(n19984), .ZN(
        n14158) );
  AOI22_X1 U17630 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19587), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19588), .ZN(n19938) );
  AOI22_X1 U17631 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19588), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19587), .ZN(n19897) );
  INV_X1 U17632 ( .A(n19984), .ZN(n14161) );
  NAND2_X1 U17633 ( .A1(n10855), .A2(n14160), .ZN(n19612) );
  OAI22_X1 U17634 ( .A1(n19897), .A2(n14162), .B1(n14161), .B2(n19612), .ZN(
        n14163) );
  AOI21_X1 U17635 ( .B1(n19985), .B2(n20039), .A(n14163), .ZN(n14169) );
  OAI21_X1 U17636 ( .B1(n14164), .B2(n19984), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14165) );
  NOR2_X2 U17637 ( .A1(n15353), .A2(n19915), .ZN(n20037) );
  NAND2_X1 U17638 ( .A1(n19986), .A2(n20037), .ZN(n14168) );
  OAI211_X1 U17639 ( .C1(n19990), .C2(n14170), .A(n14169), .B(n14168), .ZN(
        P2_U3165) );
  NOR2_X1 U17640 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n14185) );
  INV_X1 U17641 ( .A(n14185), .ZN(n19644) );
  NOR2_X1 U17642 ( .A1(n19850), .A2(n19644), .ZN(n19637) );
  INV_X1 U17643 ( .A(n19637), .ZN(n14179) );
  OAI21_X1 U17644 ( .B1(n14171), .B2(n20065), .A(n19920), .ZN(n14175) );
  AOI21_X1 U17645 ( .B1(n19623), .B2(n19664), .A(n19595), .ZN(n14172) );
  AOI21_X1 U17646 ( .B1(n14173), .B2(n14185), .A(n14172), .ZN(n14174) );
  AOI211_X1 U17647 ( .C1(n14179), .C2(n14175), .A(n19915), .B(n14174), .ZN(
        n19624) );
  INV_X1 U17648 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14183) );
  AND2_X1 U17649 ( .A1(n14176), .A2(n14179), .ZN(n14177) );
  OAI22_X1 U17650 ( .A1(n14177), .A2(n20065), .B1(n19644), .B2(n19853), .ZN(
        n19638) );
  AOI22_X1 U17651 ( .A1(n19668), .A2(n20005), .B1(n19639), .B2(n20004), .ZN(
        n14178) );
  OAI21_X1 U17652 ( .B1(n14180), .B2(n14179), .A(n14178), .ZN(n14181) );
  AOI21_X1 U17653 ( .B1(n19638), .B2(n20003), .A(n14181), .ZN(n14182) );
  OAI21_X1 U17654 ( .B1(n19624), .B2(n14183), .A(n14182), .ZN(P2_U3064) );
  OR2_X1 U17655 ( .A1(n19818), .A2(n19760), .ZN(n14332) );
  NOR3_X1 U17656 ( .A1(n20053), .A2(n19619), .A3(n20150), .ZN(n14184) );
  NOR2_X1 U17657 ( .A1(n14184), .A2(n20147), .ZN(n14194) );
  INV_X1 U17658 ( .A(n14194), .ZN(n14188) );
  NAND2_X1 U17659 ( .A1(n14185), .A2(n10356), .ZN(n19599) );
  NOR2_X1 U17660 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19599), .ZN(
        n19585) );
  INV_X1 U17661 ( .A(n19585), .ZN(n14189) );
  AND2_X1 U17662 ( .A1(n19993), .A2(n14189), .ZN(n14193) );
  AOI211_X1 U17663 ( .C1(n14186), .C2(n19920), .A(n20157), .B(n19585), .ZN(
        n14187) );
  INV_X1 U17664 ( .A(n19619), .ZN(n14190) );
  OAI22_X1 U17665 ( .A1(n19897), .A2(n14190), .B1(n19612), .B2(n14189), .ZN(
        n14191) );
  AOI21_X1 U17666 ( .B1(n20039), .B2(n20053), .A(n14191), .ZN(n14196) );
  OAI21_X1 U17667 ( .B1(n14186), .B2(n19585), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14192) );
  NAND2_X1 U17668 ( .A1(n19589), .A2(n20037), .ZN(n14195) );
  OAI211_X1 U17669 ( .C1(n19593), .C2(n14197), .A(n14196), .B(n14195), .ZN(
        P2_U3053) );
  AOI21_X1 U17670 ( .B1(n20495), .B2(n14199), .A(n21095), .ZN(n14200) );
  AOI21_X1 U17671 ( .B1(n20543), .B2(n20698), .A(n14200), .ZN(n14201) );
  NOR2_X1 U17672 ( .A1(n14201), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14203) );
  NOR2_X1 U17673 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14202), .ZN(
        n20491) );
  NAND2_X1 U17674 ( .A1(n14204), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20621) );
  NAND2_X1 U17675 ( .A1(n20621), .A2(n14311), .ZN(n20703) );
  NAND2_X1 U17676 ( .A1(n20492), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n14209) );
  INV_X1 U17677 ( .A(n20491), .ZN(n14220) );
  NOR2_X1 U17678 ( .A1(n20616), .A2(n20743), .ZN(n14206) );
  OR2_X1 U17679 ( .A1(n14204), .A2(n20806), .ZN(n20706) );
  INV_X1 U17680 ( .A(n20706), .ZN(n14244) );
  NAND2_X1 U17681 ( .A1(n20574), .A2(n20573), .ZN(n14317) );
  INV_X1 U17682 ( .A(n14317), .ZN(n14205) );
  AOI22_X1 U17683 ( .A1(n20543), .A2(n14206), .B1(n14244), .B2(n14205), .ZN(
        n20485) );
  INV_X1 U17684 ( .A(n20779), .ZN(n14271) );
  OAI22_X1 U17685 ( .A1(n20644), .A2(n14220), .B1(n20485), .B2(n14271), .ZN(
        n14207) );
  AOI21_X1 U17686 ( .B1(n20508), .B2(n20781), .A(n14207), .ZN(n14208) );
  OAI211_X1 U17687 ( .C1(n20495), .C2(n20784), .A(n14209), .B(n14208), .ZN(
        P1_U3070) );
  NAND2_X1 U17688 ( .A1(n20492), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n14213) );
  OAI22_X1 U17689 ( .A1(n14210), .A2(n20485), .B1(n20654), .B2(n14220), .ZN(
        n14211) );
  AOI21_X1 U17690 ( .B1(n20508), .B2(n20797), .A(n14211), .ZN(n14212) );
  OAI211_X1 U17691 ( .C1(n20495), .C2(n20803), .A(n14213), .B(n14212), .ZN(
        P1_U3072) );
  NAND2_X1 U17692 ( .A1(n20492), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n14216) );
  OAI22_X1 U17693 ( .A1(n20627), .A2(n14220), .B1(n20485), .B2(n14251), .ZN(
        n14214) );
  AOI21_X1 U17694 ( .B1(n20508), .B2(n20711), .A(n14214), .ZN(n14215) );
  OAI211_X1 U17695 ( .C1(n20495), .C2(n20714), .A(n14216), .B(n14215), .ZN(
        P1_U3066) );
  NAND2_X1 U17696 ( .A1(n20492), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n14219) );
  INV_X1 U17697 ( .A(n20761), .ZN(n14263) );
  OAI22_X1 U17698 ( .A1(n20631), .A2(n14220), .B1(n20485), .B2(n14263), .ZN(
        n14217) );
  AOI21_X1 U17699 ( .B1(n20508), .B2(n20763), .A(n14217), .ZN(n14218) );
  OAI211_X1 U17700 ( .C1(n20495), .C2(n20766), .A(n14219), .B(n14218), .ZN(
        P1_U3067) );
  NAND2_X1 U17701 ( .A1(n20492), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n14223) );
  OAI22_X1 U17702 ( .A1(n20640), .A2(n14220), .B1(n20485), .B2(n14247), .ZN(
        n14221) );
  AOI21_X1 U17703 ( .B1(n20508), .B2(n20721), .A(n14221), .ZN(n14222) );
  OAI211_X1 U17704 ( .C1(n20495), .C2(n20724), .A(n14223), .B(n14222), .ZN(
        P1_U3069) );
  XOR2_X1 U17705 ( .A(n14225), .B(n14224), .Z(n16184) );
  INV_X1 U17706 ( .A(n16184), .ZN(n14236) );
  NAND2_X1 U17707 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14410), .ZN(
        n14226) );
  NOR2_X1 U17708 ( .A1(n14227), .A2(n14226), .ZN(n14940) );
  OAI21_X1 U17709 ( .B1(n15101), .B2(n14940), .A(n15070), .ZN(n14411) );
  INV_X1 U17710 ( .A(n14411), .ZN(n15100) );
  OAI211_X1 U17711 ( .C1(n14229), .C2(n14410), .A(n15100), .B(n14228), .ZN(
        n16267) );
  NAND2_X1 U17712 ( .A1(n16285), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n16185) );
  OAI21_X1 U17713 ( .B1(n20273), .B2(n16239), .A(n16185), .ZN(n14234) );
  INV_X1 U17714 ( .A(n14410), .ZN(n14230) );
  NOR2_X1 U17715 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14230), .ZN(
        n16268) );
  INV_X1 U17716 ( .A(n16268), .ZN(n14231) );
  NOR2_X1 U17717 ( .A1(n14232), .A2(n14231), .ZN(n14233) );
  AOI211_X1 U17718 ( .C1(n16267), .C2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n14234), .B(n14233), .ZN(n14235) );
  OAI21_X1 U17719 ( .B1(n14236), .B2(n16222), .A(n14235), .ZN(P1_U3026) );
  NOR2_X1 U17720 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20741), .ZN(
        n15128) );
  OAI21_X1 U17721 ( .B1(n20788), .B2(n15130), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14240) );
  INV_X1 U17722 ( .A(n14238), .ZN(n20699) );
  NAND2_X1 U17723 ( .A1(n20699), .A2(n20616), .ZN(n14239) );
  AOI21_X1 U17724 ( .B1(n14240), .B2(n14239), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n14241) );
  OR2_X1 U17725 ( .A1(n20574), .A2(n20661), .ZN(n20622) );
  NAND2_X1 U17726 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20622), .ZN(n20617) );
  NAND2_X1 U17727 ( .A1(n15126), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n14250) );
  INV_X1 U17728 ( .A(n15128), .ZN(n14272) );
  NAND2_X1 U17729 ( .A1(n14242), .A2(n20616), .ZN(n14246) );
  INV_X1 U17730 ( .A(n20622), .ZN(n14243) );
  NAND2_X1 U17731 ( .A1(n14244), .A2(n14243), .ZN(n14245) );
  OAI22_X1 U17732 ( .A1(n20640), .A2(n14272), .B1(n15127), .B2(n14247), .ZN(
        n14248) );
  AOI21_X1 U17733 ( .B1(n15130), .B2(n20775), .A(n14248), .ZN(n14249) );
  OAI211_X1 U17734 ( .C1(n20778), .C2(n20802), .A(n14250), .B(n14249), .ZN(
        P1_U3149) );
  NAND2_X1 U17735 ( .A1(n15126), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n14254) );
  OAI22_X1 U17736 ( .A1(n20627), .A2(n14272), .B1(n15127), .B2(n14251), .ZN(
        n14252) );
  AOI21_X1 U17737 ( .B1(n15130), .B2(n20757), .A(n14252), .ZN(n14253) );
  OAI211_X1 U17738 ( .C1(n20760), .C2(n20802), .A(n14254), .B(n14253), .ZN(
        P1_U3146) );
  NAND2_X1 U17739 ( .A1(n15126), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n14258) );
  OAI22_X1 U17740 ( .A1(n20611), .A2(n14272), .B1(n15127), .B2(n14255), .ZN(
        n14256) );
  AOI21_X1 U17741 ( .B1(n15130), .B2(n20373), .A(n14256), .ZN(n14257) );
  OAI211_X1 U17742 ( .C1(n20612), .C2(n20802), .A(n14258), .B(n14257), .ZN(
        P1_U3145) );
  INV_X1 U17743 ( .A(n20727), .ZN(n20792) );
  NAND2_X1 U17744 ( .A1(n15126), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n14262) );
  INV_X1 U17745 ( .A(n20730), .ZN(n20787) );
  INV_X1 U17746 ( .A(n20785), .ZN(n14259) );
  OAI22_X1 U17747 ( .A1(n20649), .A2(n14272), .B1(n15127), .B2(n14259), .ZN(
        n14260) );
  AOI21_X1 U17748 ( .B1(n15130), .B2(n20787), .A(n14260), .ZN(n14261) );
  OAI211_X1 U17749 ( .C1(n20802), .C2(n20792), .A(n14262), .B(n14261), .ZN(
        P1_U3151) );
  NAND2_X1 U17750 ( .A1(n15126), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n14266) );
  OAI22_X1 U17751 ( .A1(n20631), .A2(n14272), .B1(n15127), .B2(n14263), .ZN(
        n14264) );
  AOI21_X1 U17752 ( .B1(n15130), .B2(n20497), .A(n14264), .ZN(n14265) );
  OAI211_X1 U17753 ( .C1(n20635), .C2(n20802), .A(n14266), .B(n14265), .ZN(
        P1_U3147) );
  NAND2_X1 U17754 ( .A1(n15126), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n14270) );
  INV_X1 U17755 ( .A(n20767), .ZN(n14267) );
  OAI22_X1 U17756 ( .A1(n20636), .A2(n14272), .B1(n15127), .B2(n14267), .ZN(
        n14268) );
  AOI21_X1 U17757 ( .B1(n15130), .B2(n20769), .A(n14268), .ZN(n14269) );
  OAI211_X1 U17758 ( .C1(n20802), .C2(n20772), .A(n14270), .B(n14269), .ZN(
        P1_U3148) );
  NAND2_X1 U17759 ( .A1(n15126), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n14275) );
  OAI22_X1 U17760 ( .A1(n20644), .A2(n14272), .B1(n15127), .B2(n14271), .ZN(
        n14273) );
  AOI21_X1 U17761 ( .B1(n15130), .B2(n20560), .A(n14273), .ZN(n14274) );
  OAI211_X1 U17762 ( .C1(n20648), .C2(n20802), .A(n14275), .B(n14274), .ZN(
        P1_U3150) );
  INV_X1 U17763 ( .A(n9812), .ZN(n14276) );
  OAI21_X1 U17764 ( .B1(n14153), .B2(n14277), .A(n14276), .ZN(n14396) );
  INV_X1 U17765 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20827) );
  NAND3_X1 U17766 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n20286) );
  NOR2_X1 U17767 ( .A1(n20827), .A2(n20286), .ZN(n20258) );
  NAND4_X1 U17768 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20258), .A3(
        P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n14278) );
  INV_X1 U17769 ( .A(n14278), .ZN(n14288) );
  INV_X1 U17770 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20835) );
  NOR2_X1 U17771 ( .A1(n20835), .A2(n14278), .ZN(n20241) );
  NOR2_X1 U17772 ( .A1(n20241), .A2(n20259), .ZN(n14287) );
  INV_X1 U17773 ( .A(n14279), .ZN(n16283) );
  AOI21_X1 U17774 ( .B1(n16283), .B2(n14281), .A(n14280), .ZN(n14282) );
  NOR2_X1 U17775 ( .A1(n14282), .A2(n9981), .ZN(n16265) );
  INV_X1 U17776 ( .A(n16265), .ZN(n14283) );
  OAI22_X1 U17777 ( .A1(n14283), .A2(n20274), .B1(n14392), .B2(n20292), .ZN(
        n14286) );
  NOR2_X1 U17778 ( .A1(n20301), .A2(n14287), .ZN(n20250) );
  AOI22_X1 U17779 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n20306), .B1(
        P1_EBX_REG_8__SCAN_IN), .B2(n20304), .ZN(n14284) );
  INV_X1 U17780 ( .A(n20288), .ZN(n20276) );
  OAI211_X1 U17781 ( .C1(n20250), .C2(n20835), .A(n14284), .B(n20276), .ZN(
        n14285) );
  AOI211_X1 U17782 ( .C1(n14288), .C2(n14287), .A(n14286), .B(n14285), .ZN(
        n14289) );
  OAI21_X1 U17783 ( .B1(n14396), .B2(n16093), .A(n14289), .ZN(P1_U2832) );
  AOI22_X1 U17784 ( .A1(n16265), .A2(n20320), .B1(n14740), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n14290) );
  OAI21_X1 U17785 ( .B1(n14396), .B2(n14742), .A(n14290), .ZN(P1_U2864) );
  AOI22_X1 U17786 ( .A1(n14477), .A2(n14764), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14783), .ZN(n14291) );
  OAI21_X1 U17787 ( .B1(n14396), .B2(n14793), .A(n14291), .ZN(P1_U2896) );
  XNOR2_X1 U17788 ( .A(n14142), .B(n14292), .ZN(n14298) );
  INV_X1 U17789 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n19278) );
  OR2_X1 U17790 ( .A1(n14295), .A2(n14294), .ZN(n14296) );
  NAND2_X1 U17791 ( .A1(n14293), .A2(n14296), .ZN(n16526) );
  MUX2_X1 U17792 ( .A(n19278), .B(n16526), .S(n19406), .Z(n14297) );
  OAI21_X1 U17793 ( .B1(n14298), .B2(n19403), .A(n14297), .ZN(P2_U2872) );
  OAI21_X1 U17794 ( .B1(n14299), .B2(n14301), .A(n14300), .ZN(n19399) );
  NOR2_X1 U17795 ( .A1(n14302), .A2(n9740), .ZN(n14303) );
  OR2_X1 U17796 ( .A1(n14366), .A2(n14303), .ZN(n19274) );
  INV_X1 U17797 ( .A(n19274), .ZN(n14307) );
  OAI22_X1 U17798 ( .A1(n15369), .A2(n14305), .B1(n14304), .B2(n19428), .ZN(
        n14306) );
  AOI21_X1 U17799 ( .B1(n19417), .B2(n14307), .A(n14306), .ZN(n14309) );
  AOI22_X1 U17800 ( .A1(n19418), .A2(BUF2_REG_16__SCAN_IN), .B1(n19419), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n14308) );
  OAI211_X1 U17801 ( .C1(n19399), .C2(n15373), .A(n14309), .B(n14308), .ZN(
        P2_U2903) );
  NOR2_X1 U17802 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14310), .ZN(
        n20392) );
  OAI21_X1 U17803 ( .B1(n20700), .B2(n20392), .A(n20619), .ZN(n14315) );
  OAI21_X1 U17804 ( .B1(n20409), .B2(n20798), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14312) );
  NAND2_X1 U17805 ( .A1(n14312), .A2(n20696), .ZN(n14319) );
  NOR2_X1 U17806 ( .A1(n14313), .A2(n20616), .ZN(n14316) );
  NOR2_X1 U17807 ( .A1(n14319), .A2(n14316), .ZN(n14314) );
  INV_X1 U17808 ( .A(n14316), .ZN(n14318) );
  OAI22_X1 U17809 ( .A1(n14319), .A2(n14318), .B1(n14317), .B2(n20621), .ZN(
        n20393) );
  AOI22_X1 U17810 ( .A1(n20409), .A2(n20781), .B1(n20392), .B2(n20780), .ZN(
        n14320) );
  OAI21_X1 U17811 ( .B1(n20784), .B2(n20791), .A(n14320), .ZN(n14321) );
  AOI21_X1 U17812 ( .B1(n20393), .B2(n20779), .A(n14321), .ZN(n14322) );
  OAI21_X1 U17813 ( .B1(n20397), .B2(n14323), .A(n14322), .ZN(P1_U3038) );
  NOR2_X1 U17814 ( .A1(n9812), .A2(n14324), .ZN(n14325) );
  OR2_X1 U17815 ( .A1(n9800), .A2(n14325), .ZN(n14417) );
  AOI22_X1 U17816 ( .A1(n14477), .A2(n14760), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14783), .ZN(n14326) );
  OAI21_X1 U17817 ( .B1(n14417), .B2(n14793), .A(n14326), .ZN(P1_U2895) );
  INV_X1 U17818 ( .A(n19589), .ZN(n14337) );
  INV_X1 U17819 ( .A(n20010), .ZN(n14330) );
  INV_X1 U17820 ( .A(n19593), .ZN(n14334) );
  AOI22_X1 U17821 ( .A1(n20011), .A2(n19619), .B1(n20009), .B2(n19585), .ZN(
        n14327) );
  OAI21_X1 U17822 ( .B1(n14332), .B2(n19926), .A(n14327), .ZN(n14328) );
  AOI21_X1 U17823 ( .B1(n14334), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A(
        n14328), .ZN(n14329) );
  OAI21_X1 U17824 ( .B1(n14337), .B2(n14330), .A(n14329), .ZN(P2_U3049) );
  INV_X1 U17825 ( .A(n20003), .ZN(n14336) );
  AOI22_X1 U17826 ( .A1(n20005), .A2(n19619), .B1(n20002), .B2(n19585), .ZN(
        n14331) );
  OAI21_X1 U17827 ( .B1(n19923), .B2(n14332), .A(n14331), .ZN(n14333) );
  AOI21_X1 U17828 ( .B1(n14334), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        n14333), .ZN(n14335) );
  OAI21_X1 U17829 ( .B1(n14337), .B2(n14336), .A(n14335), .ZN(P2_U3048) );
  AOI21_X1 U17830 ( .B1(n14339), .B2(n14338), .A(n14380), .ZN(n14340) );
  INV_X1 U17831 ( .A(n14340), .ZN(n20244) );
  OAI222_X1 U17832 ( .A1(n14417), .A2(n14742), .B1(n20324), .B2(n14341), .C1(
        n20244), .C2(n14737), .ZN(P1_U2863) );
  OAI21_X1 U17833 ( .B1(n14343), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n9695), .ZN(n14362) );
  XNOR2_X1 U17834 ( .A(n14345), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15537) );
  XNOR2_X1 U17835 ( .A(n14344), .B(n15537), .ZN(n14360) );
  OAI22_X1 U17836 ( .A1(n20096), .A2(n19324), .B1(n19501), .B2(n14346), .ZN(
        n14347) );
  AOI21_X1 U17837 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19503), .A(
        n14347), .ZN(n14348) );
  OAI21_X1 U17838 ( .B1(n16436), .B2(n14353), .A(n14348), .ZN(n14349) );
  AOI21_X1 U17839 ( .B1(n14360), .B2(n12279), .A(n14349), .ZN(n14350) );
  OAI21_X1 U17840 ( .B1(n19495), .B2(n14362), .A(n14350), .ZN(P2_U3008) );
  NOR2_X1 U17841 ( .A1(n14351), .A2(n19521), .ZN(n14352) );
  MUX2_X1 U17842 ( .A(n14352), .B(n16565), .S(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(n14359) );
  NAND2_X1 U17843 ( .A1(n19517), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n14356) );
  INV_X1 U17844 ( .A(n14353), .ZN(n14354) );
  NAND2_X1 U17845 ( .A1(n14354), .A2(n19560), .ZN(n14355) );
  OAI211_X1 U17846 ( .C1(n14357), .C2(n19554), .A(n14356), .B(n14355), .ZN(
        n14358) );
  AOI211_X1 U17847 ( .C1(n14360), .C2(n19551), .A(n14359), .B(n14358), .ZN(
        n14361) );
  OAI21_X1 U17848 ( .B1(n19556), .B2(n14362), .A(n14361), .ZN(P2_U3040) );
  INV_X1 U17849 ( .A(n14300), .ZN(n14364) );
  NAND2_X1 U17850 ( .A1(n14364), .A2(n14363), .ZN(n14398) );
  OAI21_X1 U17851 ( .B1(n14364), .B2(n14363), .A(n14398), .ZN(n14434) );
  NOR2_X1 U17852 ( .A1(n14366), .A2(n14365), .ZN(n14367) );
  NOR2_X1 U17853 ( .A1(n14401), .A2(n14367), .ZN(n19254) );
  OAI22_X1 U17854 ( .A1(n15369), .A2(n14369), .B1(n14368), .B2(n19428), .ZN(
        n14373) );
  INV_X1 U17855 ( .A(n19418), .ZN(n15357) );
  INV_X1 U17856 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n14371) );
  INV_X1 U17857 ( .A(n19419), .ZN(n15355) );
  INV_X1 U17858 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n14370) );
  OAI22_X1 U17859 ( .A1(n15357), .A2(n14371), .B1(n15355), .B2(n14370), .ZN(
        n14372) );
  AOI211_X1 U17860 ( .C1(n19417), .C2(n19254), .A(n14373), .B(n14372), .ZN(
        n14374) );
  OAI21_X1 U17861 ( .B1(n14434), .B2(n15373), .A(n14374), .ZN(P2_U2902) );
  OAI21_X1 U17862 ( .B1(n9800), .B2(n14376), .A(n14375), .ZN(n14933) );
  AOI22_X1 U17863 ( .A1(n14477), .A2(n14757), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n14783), .ZN(n14377) );
  OAI21_X1 U17864 ( .B1(n14933), .B2(n14793), .A(n14377), .ZN(P1_U2894) );
  INV_X1 U17865 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20840) );
  NAND2_X1 U17866 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n20241), .ZN(n14378) );
  NOR2_X1 U17867 ( .A1(n20840), .A2(n14378), .ZN(n16098) );
  NOR2_X1 U17868 ( .A1(n16098), .A2(n20259), .ZN(n16110) );
  NAND2_X1 U17869 ( .A1(n20840), .A2(n14378), .ZN(n14385) );
  INV_X1 U17870 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14387) );
  OAI22_X1 U17871 ( .A1(n20289), .A2(n14387), .B1(n14929), .B2(n20292), .ZN(
        n14384) );
  NOR2_X1 U17872 ( .A1(n14380), .A2(n14379), .ZN(n14381) );
  OR2_X1 U17873 ( .A1(n16105), .A2(n14381), .ZN(n14388) );
  INV_X1 U17874 ( .A(n14388), .ZN(n16255) );
  AOI22_X1 U17875 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n20306), .B1(
        n20303), .B2(n16255), .ZN(n14382) );
  OAI211_X1 U17876 ( .C1(n20840), .C2(n16082), .A(n14382), .B(n20276), .ZN(
        n14383) );
  AOI211_X1 U17877 ( .C1(n16110), .C2(n14385), .A(n14384), .B(n14383), .ZN(
        n14386) );
  OAI21_X1 U17878 ( .B1(n14933), .B2(n16093), .A(n14386), .ZN(P1_U2830) );
  OAI222_X1 U17879 ( .A1(n14388), .A2(n14737), .B1(n14387), .B2(n20324), .C1(
        n14742), .C2(n14933), .ZN(P1_U2862) );
  XNOR2_X1 U17880 ( .A(n14389), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14390) );
  XNOR2_X1 U17881 ( .A(n14391), .B(n14390), .ZN(n16271) );
  NAND2_X1 U17882 ( .A1(n16271), .A2(n16183), .ZN(n14395) );
  AND2_X1 U17883 ( .A1(n16285), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n16264) );
  NOR2_X1 U17884 ( .A1(n16180), .A2(n14392), .ZN(n14393) );
  AOI211_X1 U17885 ( .C1(n16173), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16264), .B(n14393), .ZN(n14394) );
  OAI211_X1 U17886 ( .C1(n16120), .C2(n14396), .A(n14395), .B(n14394), .ZN(
        P1_U2991) );
  INV_X1 U17887 ( .A(n14397), .ZN(n14399) );
  AOI21_X1 U17888 ( .B1(n14399), .B2(n14398), .A(n14423), .ZN(n16403) );
  INV_X1 U17889 ( .A(n16403), .ZN(n14407) );
  OR2_X1 U17890 ( .A1(n14401), .A2(n14400), .ZN(n14402) );
  NAND2_X1 U17891 ( .A1(n14402), .A2(n14424), .ZN(n19251) );
  INV_X1 U17892 ( .A(n19251), .ZN(n15657) );
  OAI22_X1 U17893 ( .A1(n15369), .A2(n19566), .B1(n14403), .B2(n19428), .ZN(
        n14404) );
  AOI21_X1 U17894 ( .B1(n19417), .B2(n15657), .A(n14404), .ZN(n14406) );
  AOI22_X1 U17895 ( .A1(n19418), .A2(BUF2_REG_18__SCAN_IN), .B1(n19419), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n14405) );
  OAI211_X1 U17896 ( .C1(n14407), .C2(n15373), .A(n14406), .B(n14405), .ZN(
        P2_U2901) );
  XNOR2_X1 U17897 ( .A(n16158), .B(n16259), .ZN(n14408) );
  XNOR2_X1 U17898 ( .A(n14409), .B(n14408), .ZN(n14420) );
  NAND2_X1 U17899 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16272) );
  NOR2_X1 U17900 ( .A1(n16293), .A2(n16272), .ZN(n14935) );
  NAND4_X1 U17901 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A4(n14410), .ZN(n15097) );
  AOI21_X1 U17902 ( .B1(n15096), .B2(n15097), .A(n14411), .ZN(n14412) );
  NOR2_X1 U17903 ( .A1(n16209), .A2(n14952), .ZN(n14955) );
  AOI21_X1 U17904 ( .B1(n14935), .B2(n14412), .A(n14955), .ZN(n16256) );
  INV_X1 U17905 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20837) );
  OAI22_X1 U17906 ( .A1(n20244), .A2(n16239), .B1(n20837), .B2(n16238), .ZN(
        n14413) );
  AOI21_X1 U17907 ( .B1(n16256), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n14413), .ZN(n14415) );
  NAND2_X1 U17908 ( .A1(n14940), .A2(n16232), .ZN(n16287) );
  NOR3_X1 U17909 ( .A1(n16293), .A2(n16272), .A3(n16287), .ZN(n16258) );
  NAND2_X1 U17910 ( .A1(n16258), .A2(n16259), .ZN(n14414) );
  OAI211_X1 U17911 ( .C1(n14420), .C2(n16222), .A(n14415), .B(n14414), .ZN(
        P1_U3022) );
  OAI22_X1 U17912 ( .A1(n16187), .A2(n11332), .B1(n16238), .B2(n20837), .ZN(
        n14416) );
  AOI21_X1 U17913 ( .B1(n16181), .B2(n20246), .A(n14416), .ZN(n14419) );
  INV_X1 U17914 ( .A(n14417), .ZN(n20247) );
  NAND2_X1 U17915 ( .A1(n20247), .A2(n14887), .ZN(n14418) );
  OAI211_X1 U17916 ( .C1(n14420), .C2(n20226), .A(n14419), .B(n14418), .ZN(
        P1_U2990) );
  INV_X1 U17917 ( .A(n14421), .ZN(n14422) );
  NAND2_X1 U17918 ( .A1(n14423), .A2(n14422), .ZN(n15363) );
  OAI21_X1 U17919 ( .B1(n14423), .B2(n14422), .A(n15363), .ZN(n15290) );
  AOI21_X1 U17920 ( .B1(n14425), .B2(n14424), .A(n15364), .ZN(n19234) );
  OAI22_X1 U17921 ( .A1(n15369), .A2(n19570), .B1(n14426), .B2(n19428), .ZN(
        n14429) );
  INV_X1 U17922 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n14427) );
  OAI22_X1 U17923 ( .A1(n15357), .A2(n14427), .B1(n15355), .B2(n16729), .ZN(
        n14428) );
  AOI211_X1 U17924 ( .C1(n19417), .C2(n19234), .A(n14429), .B(n14428), .ZN(
        n14430) );
  OAI21_X1 U17925 ( .B1(n15290), .B2(n15373), .A(n14430), .ZN(P2_U2900) );
  INV_X2 U17926 ( .A(n19406), .ZN(n16392) );
  AOI21_X1 U17927 ( .B1(n14431), .B2(n15524), .A(n15505), .ZN(n19255) );
  INV_X1 U17928 ( .A(n19255), .ZN(n15673) );
  NOR2_X1 U17929 ( .A1(n15673), .A2(n16392), .ZN(n14432) );
  AOI21_X1 U17930 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n16392), .A(n14432), .ZN(
        n14433) );
  OAI21_X1 U17931 ( .B1(n14434), .B2(n19403), .A(n14433), .ZN(P2_U2870) );
  NAND2_X1 U17932 ( .A1(n14436), .A2(n14435), .ZN(n14454) );
  INV_X1 U17933 ( .A(n14454), .ZN(n14440) );
  OAI21_X1 U17934 ( .B1(n14440), .B2(n14439), .A(n14438), .ZN(n14914) );
  AOI21_X1 U17935 ( .B1(n14441), .B2(n14459), .A(n14465), .ZN(n16229) );
  AOI22_X1 U17936 ( .A1(n16229), .A2(n20320), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n14740), .ZN(n14442) );
  OAI21_X1 U17937 ( .B1(n14914), .B2(n14742), .A(n14442), .ZN(P1_U2858) );
  INV_X1 U17938 ( .A(n14910), .ZN(n14447) );
  AOI22_X1 U17939 ( .A1(P1_EBX_REG_14__SCAN_IN), .A2(n20304), .B1(n20303), 
        .B2(n16229), .ZN(n14443) );
  OAI211_X1 U17940 ( .C1(n20254), .C2(n11358), .A(n14443), .B(n20276), .ZN(
        n14446) );
  INV_X1 U17941 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20845) );
  INV_X1 U17942 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20838) );
  NAND2_X1 U17943 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(n16098), .ZN(n16084) );
  NOR2_X1 U17944 ( .A1(n20838), .A2(n16084), .ZN(n16085) );
  NAND2_X1 U17945 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n16085), .ZN(n14471) );
  NOR2_X1 U17946 ( .A1(n20845), .A2(n14471), .ZN(n14525) );
  INV_X1 U17947 ( .A(n14525), .ZN(n14444) );
  AOI21_X1 U17948 ( .B1(n20309), .B2(n14444), .A(n20301), .ZN(n14688) );
  AOI221_X1 U17949 ( .B1(n20259), .B2(n20845), .C1(n14471), .C2(n20845), .A(
        n14688), .ZN(n14445) );
  AOI211_X1 U17950 ( .C1(n20307), .C2(n14447), .A(n14446), .B(n14445), .ZN(
        n14448) );
  OAI21_X1 U17951 ( .B1(n14914), .B2(n16093), .A(n14448), .ZN(P1_U2826) );
  AOI22_X1 U17952 ( .A1(n14477), .A2(n14449), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14783), .ZN(n14450) );
  OAI21_X1 U17953 ( .B1(n14914), .B2(n14793), .A(n14450), .ZN(P1_U2890) );
  OAI21_X1 U17954 ( .B1(n11356), .B2(n14453), .A(n14452), .ZN(n14475) );
  OAI21_X1 U17955 ( .B1(n14475), .B2(n14476), .A(n14452), .ZN(n14483) );
  AND2_X1 U17956 ( .A1(n14483), .A2(n14484), .ZN(n14485) );
  OAI21_X1 U17957 ( .B1(n14485), .B2(n14455), .A(n14454), .ZN(n16094) );
  AOI22_X1 U17958 ( .A1(n14477), .A2(n14746), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14783), .ZN(n14456) );
  OAI21_X1 U17959 ( .B1(n16094), .B2(n14793), .A(n14456), .ZN(P1_U2891) );
  NAND2_X1 U17960 ( .A1(n15091), .A2(n14457), .ZN(n14458) );
  NAND2_X1 U17961 ( .A1(n14459), .A2(n14458), .ZN(n16240) );
  OAI22_X1 U17962 ( .A1(n16240), .A2(n14737), .B1(n16086), .B2(n20324), .ZN(
        n14460) );
  INV_X1 U17963 ( .A(n14460), .ZN(n14461) );
  OAI21_X1 U17964 ( .B1(n16094), .B2(n14742), .A(n14461), .ZN(P1_U2859) );
  AOI21_X1 U17965 ( .B1(n14463), .B2(n14438), .A(n14462), .ZN(n16149) );
  OR2_X1 U17966 ( .A1(n14465), .A2(n14464), .ZN(n14466) );
  NAND2_X1 U17967 ( .A1(n14692), .A2(n14466), .ZN(n15081) );
  OAI22_X1 U17968 ( .A1(n15081), .A2(n14737), .B1(n14469), .B2(n20324), .ZN(
        n14467) );
  AOI21_X1 U17969 ( .B1(n16149), .B2(n11783), .A(n14467), .ZN(n14468) );
  INV_X1 U17970 ( .A(n14468), .ZN(P1_U2857) );
  INV_X1 U17971 ( .A(n16149), .ZN(n14482) );
  INV_X1 U17972 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20848) );
  OAI22_X1 U17973 ( .A1(n14469), .A2(n20289), .B1(n20848), .B2(n14688), .ZN(
        n14470) );
  AOI211_X1 U17974 ( .C1(n20306), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n20288), .B(n14470), .ZN(n14472) );
  NOR3_X1 U17975 ( .A1(n20259), .A2(n20845), .A3(n14471), .ZN(n16072) );
  NAND2_X1 U17976 ( .A1(n16072), .A2(n20848), .ZN(n14687) );
  OAI211_X1 U17977 ( .C1(n15081), .C2(n20274), .A(n14472), .B(n14687), .ZN(
        n14473) );
  AOI21_X1 U17978 ( .B1(n16148), .B2(n20307), .A(n14473), .ZN(n14474) );
  OAI21_X1 U17979 ( .B1(n14482), .B2(n16093), .A(n14474), .ZN(P1_U2825) );
  XOR2_X1 U17980 ( .A(n14476), .B(n14475), .Z(n16163) );
  INV_X1 U17981 ( .A(n16163), .ZN(n14479) );
  AOI22_X1 U17982 ( .A1(n14477), .A2(n14753), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n14783), .ZN(n14478) );
  OAI21_X1 U17983 ( .B1(n14479), .B2(n14793), .A(n14478), .ZN(P1_U2893) );
  OAI222_X1 U17984 ( .A1(n14482), .A2(n14793), .B1(n14490), .B2(n14481), .C1(
        n14743), .C2(n14480), .ZN(P1_U2889) );
  INV_X1 U17985 ( .A(n14483), .ZN(n14487) );
  INV_X1 U17986 ( .A(n14484), .ZN(n14486) );
  AOI21_X1 U17987 ( .B1(n14487), .B2(n14486), .A(n14485), .ZN(n16153) );
  INV_X1 U17988 ( .A(n16153), .ZN(n14491) );
  INV_X1 U17989 ( .A(n14750), .ZN(n14489) );
  OAI222_X1 U17990 ( .A1(n14491), .A2(n14793), .B1(n14490), .B2(n14489), .C1(
        n14488), .C2(n14743), .ZN(P1_U2892) );
  XOR2_X1 U17991 ( .A(n13545), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n14497)
         );
  NAND2_X1 U17992 ( .A1(n14492), .A2(n14493), .ZN(n14494) );
  NAND2_X1 U17993 ( .A1(n14495), .A2(n14494), .ZN(n16503) );
  INV_X1 U17994 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n15196) );
  MUX2_X1 U17995 ( .A(n16503), .B(n15196), .S(n16392), .Z(n14496) );
  OAI21_X1 U17996 ( .B1(n14497), .B2(n19403), .A(n14496), .ZN(P2_U2882) );
  OAI21_X1 U17997 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16593), .A(
        n14498), .ZN(n14499) );
  INV_X1 U17998 ( .A(n14499), .ZN(n14514) );
  NAND2_X1 U17999 ( .A1(n15299), .A2(n14500), .ZN(n14506) );
  NAND2_X1 U18000 ( .A1(n10544), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14504) );
  AOI22_X1 U18001 ( .A1(n14502), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n14501), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14503) );
  AND2_X1 U18002 ( .A1(n14504), .A2(n14503), .ZN(n14505) );
  INV_X1 U18003 ( .A(n14507), .ZN(n14509) );
  OAI21_X1 U18004 ( .B1(n16309), .B2(n19554), .A(n14510), .ZN(n14511) );
  INV_X1 U18005 ( .A(n14511), .ZN(n14512) );
  OAI211_X1 U18006 ( .C1(n14514), .C2(n10193), .A(n14513), .B(n14512), .ZN(
        n14515) );
  INV_X1 U18007 ( .A(n14515), .ZN(n14518) );
  NAND2_X1 U18008 ( .A1(n14516), .A2(n16577), .ZN(n14517) );
  OAI211_X1 U18009 ( .C1(n14519), .C2(n16589), .A(n14518), .B(n14517), .ZN(
        P2_U3015) );
  AOI22_X1 U18010 ( .A1(n14523), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n14522), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14524) );
  NAND2_X1 U18011 ( .A1(n14539), .A2(n20268), .ZN(n14533) );
  INV_X1 U18012 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21058) );
  INV_X1 U18013 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21098) );
  INV_X1 U18014 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21119) );
  NAND4_X1 U18015 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n14525), .A3(
        P1_REIP_REG_16__SCAN_IN), .A4(P1_REIP_REG_15__SCAN_IN), .ZN(n14681) );
  NAND2_X1 U18016 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n16062) );
  NOR3_X1 U18017 ( .A1(n21119), .A2(n14681), .A3(n16062), .ZN(n16054) );
  NAND2_X1 U18018 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n16054), .ZN(n14657) );
  OR2_X1 U18019 ( .A1(n21098), .A2(n14657), .ZN(n14645) );
  NOR2_X1 U18020 ( .A1(n21058), .A2(n14645), .ZN(n14631) );
  AND2_X1 U18021 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n14631), .ZN(n14618) );
  NAND3_X1 U18022 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .A3(n14618), .ZN(n14594) );
  INV_X1 U18023 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20866) );
  NOR2_X1 U18024 ( .A1(n14594), .A2(n20866), .ZN(n14577) );
  AND2_X1 U18025 ( .A1(n14577), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14579) );
  NAND2_X1 U18026 ( .A1(n16082), .A2(n14579), .ZN(n14526) );
  INV_X1 U18027 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21040) );
  AOI21_X1 U18028 ( .B1(n16083), .B2(n14526), .A(n21040), .ZN(n14569) );
  INV_X1 U18029 ( .A(n16083), .ZN(n14527) );
  AOI21_X1 U18030 ( .B1(n14569), .B2(P1_REIP_REG_30__SCAN_IN), .A(n14527), 
        .ZN(n14553) );
  INV_X1 U18031 ( .A(n14579), .ZN(n14528) );
  OR3_X1 U18032 ( .A1(n20259), .A2(n21040), .A3(n14528), .ZN(n14552) );
  NOR3_X1 U18033 ( .A1(n14552), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n20959), 
        .ZN(n14531) );
  INV_X1 U18034 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14700) );
  INV_X1 U18035 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14529) );
  OAI22_X1 U18036 ( .A1(n20289), .A2(n14700), .B1(n14529), .B2(n20254), .ZN(
        n14530) );
  AOI211_X1 U18037 ( .C1(n14553), .C2(P1_REIP_REG_31__SCAN_IN), .A(n14531), 
        .B(n14530), .ZN(n14532) );
  OAI211_X1 U18038 ( .C1(n14934), .C2(n20274), .A(n14533), .B(n14532), .ZN(
        P1_U2809) );
  NOR2_X1 U18039 ( .A1(n12322), .A2(n16392), .ZN(n14534) );
  AOI21_X1 U18040 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n16392), .A(n14534), .ZN(
        n14535) );
  OAI21_X1 U18041 ( .B1(n14536), .B2(n19403), .A(n14535), .ZN(P2_U2857) );
  AND2_X1 U18042 ( .A1(n14743), .A2(n14537), .ZN(n14538) );
  NAND2_X1 U18043 ( .A1(n14539), .A2(n14538), .ZN(n14541) );
  AOI22_X1 U18044 ( .A1(n14800), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14783), .ZN(n14540) );
  OAI211_X1 U18045 ( .C1(n14767), .C2(n16706), .A(n14541), .B(n14540), .ZN(
        P1_U2873) );
  NAND2_X1 U18046 ( .A1(n14542), .A2(n20314), .ZN(n14550) );
  NAND2_X1 U18047 ( .A1(n20304), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n14544) );
  AOI22_X1 U18048 ( .A1(n20306), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20301), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n14543) );
  OAI211_X1 U18049 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20292), .A(
        n14544), .B(n14543), .ZN(n14548) );
  NAND2_X1 U18050 ( .A1(n20303), .A2(n14545), .ZN(n14546) );
  OAI21_X1 U18051 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20259), .A(n14546), .ZN(
        n14547) );
  NOR2_X1 U18052 ( .A1(n14548), .A2(n14547), .ZN(n14549) );
  OAI211_X1 U18053 ( .C1(n20312), .C2(n20698), .A(n14550), .B(n14549), .ZN(
        P1_U2839) );
  INV_X1 U18054 ( .A(n14551), .ZN(n14974) );
  INV_X1 U18055 ( .A(n14552), .ZN(n14554) );
  OAI21_X1 U18056 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14554), .A(n14553), 
        .ZN(n14557) );
  AOI22_X1 U18057 ( .A1(n14555), .A2(n20307), .B1(n20306), .B2(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14556) );
  OAI211_X1 U18058 ( .C1(n20289), .C2(n14558), .A(n14557), .B(n14556), .ZN(
        n14559) );
  AOI21_X1 U18059 ( .B1(n14974), .B2(n20303), .A(n14559), .ZN(n14560) );
  OAI21_X1 U18060 ( .B1(n14561), .B2(n16093), .A(n14560), .ZN(P1_U2810) );
  AOI21_X1 U18061 ( .B1(n14563), .B2(n9726), .A(n14562), .ZN(n14813) );
  INV_X1 U18062 ( .A(n14813), .ZN(n14749) );
  INV_X1 U18063 ( .A(n14564), .ZN(n14565) );
  XNOR2_X1 U18064 ( .A(n14576), .B(n14565), .ZN(n14982) );
  AOI21_X1 U18065 ( .B1(n20309), .B2(n14579), .A(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14568) );
  AOI22_X1 U18066 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n20306), .B1(
        n20307), .B2(n14809), .ZN(n14567) );
  NAND2_X1 U18067 ( .A1(n20304), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14566) );
  OAI211_X1 U18068 ( .C1(n14569), .C2(n14568), .A(n14567), .B(n14566), .ZN(
        n14570) );
  AOI21_X1 U18069 ( .B1(n14982), .B2(n20303), .A(n14570), .ZN(n14571) );
  OAI21_X1 U18070 ( .B1(n14749), .B2(n16093), .A(n14571), .ZN(P1_U2811) );
  OAI21_X1 U18071 ( .B1(n14572), .B2(n14573), .A(n9726), .ZN(n14829) );
  NOR2_X1 U18072 ( .A1(n14586), .A2(n14574), .ZN(n14575) );
  OR2_X1 U18073 ( .A1(n14576), .A2(n14575), .ZN(n14997) );
  INV_X1 U18074 ( .A(n14997), .ZN(n14584) );
  NOR2_X1 U18075 ( .A1(n14577), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14578) );
  NOR3_X1 U18076 ( .A1(n20259), .A2(n14579), .A3(n14578), .ZN(n14583) );
  INV_X1 U18077 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14702) );
  AOI22_X1 U18078 ( .A1(n20306), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n20301), .B2(P1_REIP_REG_28__SCAN_IN), .ZN(n14581) );
  NAND2_X1 U18079 ( .A1(n20307), .A2(n14817), .ZN(n14580) );
  OAI211_X1 U18080 ( .C1(n20289), .C2(n14702), .A(n14581), .B(n14580), .ZN(
        n14582) );
  AOI211_X1 U18081 ( .C1(n14584), .C2(n20303), .A(n14583), .B(n14582), .ZN(
        n14585) );
  OAI21_X1 U18082 ( .B1(n14829), .B2(n16093), .A(n14585), .ZN(P1_U2812) );
  INV_X1 U18083 ( .A(n14586), .ZN(n14589) );
  NAND2_X1 U18084 ( .A1(n14605), .A2(n14587), .ZN(n14588) );
  NAND2_X1 U18085 ( .A1(n14589), .A2(n14588), .ZN(n15005) );
  AOI21_X1 U18086 ( .B1(n14591), .B2(n14590), .A(n14572), .ZN(n14836) );
  NAND2_X1 U18087 ( .A1(n14836), .A2(n20268), .ZN(n14601) );
  INV_X1 U18088 ( .A(n14594), .ZN(n14592) );
  NAND2_X1 U18089 ( .A1(n16082), .A2(n14592), .ZN(n14593) );
  AND2_X1 U18090 ( .A1(n16083), .A2(n14593), .ZN(n14606) );
  NAND2_X1 U18091 ( .A1(n20304), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n14598) );
  OR3_X1 U18092 ( .A1(n20259), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14594), .ZN(
        n14597) );
  INV_X1 U18093 ( .A(n14834), .ZN(n14595) );
  AOI22_X1 U18094 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n20306), .B1(
        n20307), .B2(n14595), .ZN(n14596) );
  NAND3_X1 U18095 ( .A1(n14598), .A2(n14597), .A3(n14596), .ZN(n14599) );
  AOI21_X1 U18096 ( .B1(n14606), .B2(P1_REIP_REG_27__SCAN_IN), .A(n14599), 
        .ZN(n14600) );
  OAI211_X1 U18097 ( .C1(n20274), .C2(n15005), .A(n14601), .B(n14600), .ZN(
        P1_U2813) );
  OAI21_X1 U18098 ( .B1(n14602), .B2(n10185), .A(n14590), .ZN(n14845) );
  NAND2_X1 U18099 ( .A1(n9754), .A2(n14603), .ZN(n14604) );
  NAND2_X1 U18100 ( .A1(n14605), .A2(n14604), .ZN(n14705) );
  INV_X1 U18101 ( .A(n14705), .ZN(n15016) );
  AND3_X1 U18102 ( .A1(n20309), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n14618), 
        .ZN(n14607) );
  OAI21_X1 U18103 ( .B1(n14607), .B2(P1_REIP_REG_26__SCAN_IN), .A(n14606), 
        .ZN(n14609) );
  AOI22_X1 U18104 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n20306), .B1(
        n20307), .B2(n14840), .ZN(n14608) );
  OAI211_X1 U18105 ( .C1(n14704), .C2(n20289), .A(n14609), .B(n14608), .ZN(
        n14610) );
  AOI21_X1 U18106 ( .B1(n15016), .B2(n20303), .A(n14610), .ZN(n14611) );
  OAI21_X1 U18107 ( .B1(n14845), .B2(n16093), .A(n14611), .ZN(P1_U2814) );
  BUF_X1 U18108 ( .A(n14612), .Z(n14613) );
  AOI21_X1 U18109 ( .B1(n14614), .B2(n14613), .A(n14602), .ZN(n14853) );
  NAND2_X1 U18110 ( .A1(n9808), .A2(n14615), .ZN(n14616) );
  NAND2_X1 U18111 ( .A1(n9754), .A2(n14616), .ZN(n15024) );
  OAI22_X1 U18112 ( .A1(n14617), .A2(n20254), .B1(n20292), .B2(n14851), .ZN(
        n14621) );
  INV_X1 U18113 ( .A(n14618), .ZN(n14619) );
  NOR3_X1 U18114 ( .A1(n20259), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n14619), 
        .ZN(n14620) );
  AOI211_X1 U18115 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n20304), .A(n14621), .B(
        n14620), .ZN(n14624) );
  NOR2_X1 U18116 ( .A1(n20259), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14630) );
  OR2_X1 U18117 ( .A1(n20259), .A2(n14631), .ZN(n14622) );
  NAND2_X1 U18118 ( .A1(n14622), .A2(n16082), .ZN(n14650) );
  OAI21_X1 U18119 ( .B1(n14630), .B2(n14650), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14623) );
  OAI211_X1 U18120 ( .C1(n15024), .C2(n20274), .A(n14624), .B(n14623), .ZN(
        n14625) );
  AOI21_X1 U18121 ( .B1(n14853), .B2(n20268), .A(n14625), .ZN(n14626) );
  INV_X1 U18122 ( .A(n14626), .ZN(P1_U2815) );
  BUF_X1 U18123 ( .A(n14627), .Z(n14628) );
  OAI21_X1 U18124 ( .B1(n14628), .B2(n14629), .A(n14613), .ZN(n14859) );
  INV_X1 U18125 ( .A(n14859), .ZN(n14640) );
  AOI22_X1 U18126 ( .A1(P1_EBX_REG_24__SCAN_IN), .A2(n20304), .B1(n14631), 
        .B2(n14630), .ZN(n14632) );
  OAI21_X1 U18127 ( .B1(n14858), .B2(n20254), .A(n14632), .ZN(n14639) );
  INV_X1 U18128 ( .A(n14633), .ZN(n14642) );
  NAND2_X1 U18129 ( .A1(n14654), .A2(n14642), .ZN(n14635) );
  NAND2_X1 U18130 ( .A1(n14635), .A2(n14634), .ZN(n14636) );
  NAND2_X1 U18131 ( .A1(n14636), .A2(n9808), .ZN(n15035) );
  AOI22_X1 U18132 ( .A1(n14650), .A2(P1_REIP_REG_24__SCAN_IN), .B1(n14862), 
        .B2(n20307), .ZN(n14637) );
  OAI21_X1 U18133 ( .B1(n15035), .B2(n20274), .A(n14637), .ZN(n14638) );
  AOI211_X1 U18134 ( .C1(n14640), .C2(n20268), .A(n14639), .B(n14638), .ZN(
        n14641) );
  INV_X1 U18135 ( .A(n14641), .ZN(P1_U2816) );
  XNOR2_X1 U18136 ( .A(n14654), .B(n14642), .ZN(n16192) );
  INV_X1 U18137 ( .A(n14643), .ZN(n14644) );
  AOI21_X1 U18138 ( .B1(n14644), .B2(n9725), .A(n14628), .ZN(n14868) );
  NAND2_X1 U18139 ( .A1(n14868), .A2(n20268), .ZN(n14652) );
  OAI21_X1 U18140 ( .B1(n20259), .B2(n14645), .A(n21058), .ZN(n14649) );
  OAI22_X1 U18141 ( .A1(n14646), .A2(n20254), .B1(n20292), .B2(n14866), .ZN(
        n14648) );
  NOR2_X1 U18142 ( .A1(n20289), .A2(n14708), .ZN(n14647) );
  AOI211_X1 U18143 ( .C1(n14650), .C2(n14649), .A(n14648), .B(n14647), .ZN(
        n14651) );
  OAI211_X1 U18144 ( .C1(n16192), .C2(n20274), .A(n14652), .B(n14651), .ZN(
        P1_U2817) );
  INV_X1 U18145 ( .A(n14654), .ZN(n14655) );
  OAI21_X1 U18146 ( .B1(n14656), .B2(n14714), .A(n14655), .ZN(n16201) );
  NOR2_X1 U18147 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n20259), .ZN(n16053) );
  OAI21_X1 U18148 ( .B1(n16054), .B2(n20259), .A(n16082), .ZN(n16052) );
  OAI21_X1 U18149 ( .B1(n16053), .B2(n16052), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14659) );
  OR3_X1 U18150 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n20259), .A3(n14657), .ZN(
        n14658) );
  OAI211_X1 U18151 ( .C1(n16201), .C2(n20274), .A(n14659), .B(n14658), .ZN(
        n14662) );
  AOI22_X1 U18152 ( .A1(n14877), .A2(n20307), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n20304), .ZN(n14660) );
  OAI21_X1 U18153 ( .B1(n14873), .B2(n20254), .A(n14660), .ZN(n14661) );
  NOR2_X1 U18154 ( .A1(n14662), .A2(n14661), .ZN(n14663) );
  OAI21_X1 U18155 ( .B1(n14874), .B2(n16093), .A(n14663), .ZN(P1_U2818) );
  OAI21_X1 U18156 ( .B1(n14664), .B2(n14666), .A(n14665), .ZN(n14895) );
  OR2_X1 U18157 ( .A1(n20259), .A2(n14681), .ZN(n16064) );
  OAI21_X1 U18158 ( .B1(n16062), .B2(n16064), .A(n21119), .ZN(n14673) );
  NAND2_X1 U18159 ( .A1(n14727), .A2(n14667), .ZN(n14668) );
  AND2_X1 U18160 ( .A1(n9752), .A2(n14668), .ZN(n16028) );
  INV_X1 U18161 ( .A(n16028), .ZN(n14671) );
  OAI22_X1 U18162 ( .A1(n14889), .A2(n20254), .B1(n14719), .B2(n20289), .ZN(
        n14669) );
  AOI21_X1 U18163 ( .B1(n20307), .B2(n14891), .A(n14669), .ZN(n14670) );
  OAI21_X1 U18164 ( .B1(n14671), .B2(n20274), .A(n14670), .ZN(n14672) );
  AOI21_X1 U18165 ( .B1(n14673), .B2(n16052), .A(n14672), .ZN(n14674) );
  OAI21_X1 U18166 ( .B1(n14895), .B2(n16093), .A(n14674), .ZN(P1_U2820) );
  AOI21_X1 U18167 ( .B1(n14678), .B2(n10137), .A(n14677), .ZN(n14901) );
  INV_X1 U18168 ( .A(n14901), .ZN(n14794) );
  AOI21_X1 U18169 ( .B1(n14679), .B2(n14736), .A(n14725), .ZN(n16214) );
  INV_X1 U18170 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14680) );
  OAI22_X1 U18171 ( .A1(n20289), .A2(n14680), .B1(n14899), .B2(n20292), .ZN(
        n14684) );
  INV_X1 U18172 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20855) );
  AOI21_X1 U18173 ( .B1(n20309), .B2(n14681), .A(n20301), .ZN(n16080) );
  AOI21_X1 U18174 ( .B1(n20306), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20288), .ZN(n14682) );
  OAI221_X1 U18175 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n16064), .C1(n20855), 
        .C2(n16080), .A(n14682), .ZN(n14683) );
  AOI211_X1 U18176 ( .C1(n16214), .C2(n20303), .A(n14684), .B(n14683), .ZN(
        n14685) );
  OAI21_X1 U18177 ( .B1(n14794), .B2(n16093), .A(n14685), .ZN(P1_U2822) );
  XOR2_X1 U18178 ( .A(n14686), .B(n14462), .Z(n16144) );
  INV_X1 U18179 ( .A(n16144), .ZN(n14805) );
  INV_X1 U18180 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20851) );
  AOI21_X1 U18181 ( .B1(n14688), .B2(n14687), .A(n20851), .ZN(n14698) );
  NAND3_X1 U18182 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n16072), .A3(n20851), 
        .ZN(n14689) );
  OAI211_X1 U18183 ( .C1(n20254), .C2(n14690), .A(n20276), .B(n14689), .ZN(
        n14697) );
  INV_X1 U18184 ( .A(n14734), .ZN(n14691) );
  AOI21_X1 U18185 ( .B1(n14693), .B2(n14692), .A(n14691), .ZN(n15074) );
  INV_X1 U18186 ( .A(n15074), .ZN(n14695) );
  AOI22_X1 U18187 ( .A1(n20304), .A2(P1_EBX_REG_16__SCAN_IN), .B1(n20307), 
        .B2(n16143), .ZN(n14694) );
  OAI21_X1 U18188 ( .B1(n14695), .B2(n20274), .A(n14694), .ZN(n14696) );
  NOR3_X1 U18189 ( .A1(n14698), .A2(n14697), .A3(n14696), .ZN(n14699) );
  OAI21_X1 U18190 ( .B1(n14805), .B2(n16093), .A(n14699), .ZN(P1_U2824) );
  OAI22_X1 U18191 ( .A1(n14934), .A2(n14737), .B1(n14700), .B2(n20324), .ZN(
        P1_U2841) );
  AOI22_X1 U18192 ( .A1(n14982), .A2(n20320), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14740), .ZN(n14701) );
  OAI21_X1 U18193 ( .B1(n14749), .B2(n14742), .A(n14701), .ZN(P1_U2843) );
  OAI222_X1 U18194 ( .A1(n14702), .A2(n20324), .B1(n14737), .B2(n14997), .C1(
        n14829), .C2(n14742), .ZN(P1_U2844) );
  INV_X1 U18195 ( .A(n14836), .ZN(n14756) );
  OAI222_X1 U18196 ( .A1(n14703), .A2(n20324), .B1(n14737), .B2(n15005), .C1(
        n14756), .C2(n14742), .ZN(P1_U2845) );
  OAI222_X1 U18197 ( .A1(n14705), .A2(n14737), .B1(n14704), .B2(n20324), .C1(
        n14845), .C2(n14742), .ZN(P1_U2846) );
  INV_X1 U18198 ( .A(n14853), .ZN(n14763) );
  OAI222_X1 U18199 ( .A1(n14706), .A2(n20324), .B1(n14737), .B2(n15024), .C1(
        n14763), .C2(n14742), .ZN(P1_U2847) );
  INV_X1 U18200 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14707) );
  OAI222_X1 U18201 ( .A1(n14742), .A2(n14859), .B1(n20324), .B2(n14707), .C1(
        n15035), .C2(n14737), .ZN(P1_U2848) );
  INV_X1 U18202 ( .A(n14868), .ZN(n14775) );
  OAI222_X1 U18203 ( .A1(n14775), .A2(n14742), .B1(n14737), .B2(n16192), .C1(
        n20324), .C2(n14708), .ZN(P1_U2849) );
  INV_X1 U18204 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14709) );
  OAI222_X1 U18205 ( .A1(n14874), .A2(n14742), .B1(n20324), .B2(n14709), .C1(
        n16201), .C2(n14737), .ZN(P1_U2850) );
  NAND2_X1 U18206 ( .A1(n14665), .A2(n14710), .ZN(n14711) );
  AND2_X1 U18207 ( .A1(n9752), .A2(n14713), .ZN(n14715) );
  OR2_X1 U18208 ( .A1(n14715), .A2(n14714), .ZN(n16057) );
  OAI22_X1 U18209 ( .A1(n16057), .A2(n14737), .B1(n14716), .B2(n20324), .ZN(
        n14717) );
  INV_X1 U18210 ( .A(n14717), .ZN(n14718) );
  OAI21_X1 U18211 ( .B1(n14782), .B2(n14742), .A(n14718), .ZN(P1_U2851) );
  NOR2_X1 U18212 ( .A1(n20324), .A2(n14719), .ZN(n14720) );
  AOI21_X1 U18213 ( .B1(n16028), .B2(n20320), .A(n14720), .ZN(n14721) );
  OAI21_X1 U18214 ( .B1(n14895), .B2(n14742), .A(n14721), .ZN(P1_U2852) );
  NOR2_X1 U18215 ( .A1(n14677), .A2(n14722), .ZN(n14723) );
  OR2_X1 U18216 ( .A1(n14664), .A2(n14723), .ZN(n16121) );
  OR2_X1 U18217 ( .A1(n14725), .A2(n14724), .ZN(n14726) );
  AND2_X1 U18218 ( .A1(n14727), .A2(n14726), .ZN(n16066) );
  NOR2_X1 U18219 ( .A1(n20324), .A2(n16071), .ZN(n14728) );
  AOI21_X1 U18220 ( .B1(n16066), .B2(n20320), .A(n14728), .ZN(n14729) );
  OAI21_X1 U18221 ( .B1(n16121), .B2(n14742), .A(n14729), .ZN(P1_U2853) );
  AOI22_X1 U18222 ( .A1(n16214), .A2(n20320), .B1(n14740), .B2(
        P1_EBX_REG_18__SCAN_IN), .ZN(n14730) );
  OAI21_X1 U18223 ( .B1(n14794), .B2(n14742), .A(n14730), .ZN(P1_U2854) );
  AOI21_X1 U18224 ( .B1(n14732), .B2(n14731), .A(n14675), .ZN(n16140) );
  INV_X1 U18225 ( .A(n16140), .ZN(n14798) );
  NAND2_X1 U18226 ( .A1(n14734), .A2(n14733), .ZN(n14735) );
  NAND2_X1 U18227 ( .A1(n14736), .A2(n14735), .ZN(n16221) );
  OAI22_X1 U18228 ( .A1(n16221), .A2(n14737), .B1(n16074), .B2(n20324), .ZN(
        n14738) );
  INV_X1 U18229 ( .A(n14738), .ZN(n14739) );
  OAI21_X1 U18230 ( .B1(n14798), .B2(n14742), .A(n14739), .ZN(P1_U2855) );
  AOI22_X1 U18231 ( .A1(n15074), .A2(n20320), .B1(n14740), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n14741) );
  OAI21_X1 U18232 ( .B1(n14805), .B2(n14742), .A(n14741), .ZN(P1_U2856) );
  OAI22_X1 U18233 ( .A1(n14767), .A2(n16710), .B1(n14744), .B2(n14743), .ZN(
        n14745) );
  INV_X1 U18234 ( .A(n14745), .ZN(n14748) );
  AOI22_X1 U18235 ( .A1(n14802), .A2(n14746), .B1(n14800), .B2(DATAI_29_), 
        .ZN(n14747) );
  OAI211_X1 U18236 ( .C1(n14749), .C2(n14793), .A(n14748), .B(n14747), .ZN(
        P1_U2875) );
  AOI22_X1 U18237 ( .A1(n14799), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14783), .ZN(n14752) );
  AOI22_X1 U18238 ( .A1(n14802), .A2(n14750), .B1(n14800), .B2(DATAI_28_), 
        .ZN(n14751) );
  OAI211_X1 U18239 ( .C1(n14829), .C2(n14793), .A(n14752), .B(n14751), .ZN(
        P1_U2876) );
  AOI22_X1 U18240 ( .A1(n14799), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n14783), .ZN(n14755) );
  AOI22_X1 U18241 ( .A1(n14802), .A2(n14753), .B1(n14800), .B2(DATAI_27_), 
        .ZN(n14754) );
  OAI211_X1 U18242 ( .C1(n14756), .C2(n14793), .A(n14755), .B(n14754), .ZN(
        P1_U2877) );
  AOI22_X1 U18243 ( .A1(n14799), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n14783), .ZN(n14759) );
  AOI22_X1 U18244 ( .A1(n14802), .A2(n14757), .B1(n14800), .B2(DATAI_26_), 
        .ZN(n14758) );
  OAI211_X1 U18245 ( .C1(n14845), .C2(n14793), .A(n14759), .B(n14758), .ZN(
        P1_U2878) );
  AOI22_X1 U18246 ( .A1(n14799), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n14783), .ZN(n14762) );
  AOI22_X1 U18247 ( .A1(n14802), .A2(n14760), .B1(n14800), .B2(DATAI_25_), 
        .ZN(n14761) );
  OAI211_X1 U18248 ( .C1(n14763), .C2(n14793), .A(n14762), .B(n14761), .ZN(
        P1_U2879) );
  AOI22_X1 U18249 ( .A1(n14799), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n14783), .ZN(n14766) );
  AOI22_X1 U18250 ( .A1(n14802), .A2(n14764), .B1(n14800), .B2(DATAI_24_), 
        .ZN(n14765) );
  OAI211_X1 U18251 ( .C1(n14859), .C2(n14793), .A(n14766), .B(n14765), .ZN(
        P1_U2880) );
  INV_X1 U18252 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16722) );
  NOR2_X1 U18253 ( .A1(n14767), .A2(n16722), .ZN(n14773) );
  INV_X1 U18254 ( .A(n14802), .ZN(n14771) );
  INV_X1 U18255 ( .A(n14800), .ZN(n14769) );
  INV_X1 U18256 ( .A(DATAI_23_), .ZN(n14768) );
  OAI22_X1 U18257 ( .A1(n14771), .A2(n14770), .B1(n14769), .B2(n14768), .ZN(
        n14772) );
  AOI211_X1 U18258 ( .C1(n14783), .C2(P1_EAX_REG_23__SCAN_IN), .A(n14773), .B(
        n14772), .ZN(n14774) );
  OAI21_X1 U18259 ( .B1(n14775), .B2(n14793), .A(n14774), .ZN(P1_U2881) );
  AOI22_X1 U18260 ( .A1(n14799), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n14783), .ZN(n14778) );
  AOI22_X1 U18261 ( .A1(n14802), .A2(n14776), .B1(n14800), .B2(DATAI_22_), 
        .ZN(n14777) );
  OAI211_X1 U18262 ( .C1(n14874), .C2(n14793), .A(n14778), .B(n14777), .ZN(
        P1_U2882) );
  AOI22_X1 U18263 ( .A1(n14799), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n14783), .ZN(n14781) );
  AOI22_X1 U18264 ( .A1(n14802), .A2(n14779), .B1(n14800), .B2(DATAI_21_), 
        .ZN(n14780) );
  OAI211_X1 U18265 ( .C1(n14782), .C2(n14793), .A(n14781), .B(n14780), .ZN(
        P1_U2883) );
  AOI22_X1 U18266 ( .A1(n14799), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n14783), .ZN(n14786) );
  AOI22_X1 U18267 ( .A1(n14802), .A2(n14784), .B1(n14800), .B2(DATAI_20_), 
        .ZN(n14785) );
  OAI211_X1 U18268 ( .C1(n14895), .C2(n14793), .A(n14786), .B(n14785), .ZN(
        P1_U2884) );
  AOI22_X1 U18269 ( .A1(n14799), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14783), .ZN(n14789) );
  AOI22_X1 U18270 ( .A1(n14802), .A2(n14787), .B1(n14800), .B2(DATAI_19_), 
        .ZN(n14788) );
  OAI211_X1 U18271 ( .C1(n16121), .C2(n14793), .A(n14789), .B(n14788), .ZN(
        P1_U2885) );
  AOI22_X1 U18272 ( .A1(n14799), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n14783), .ZN(n14792) );
  AOI22_X1 U18273 ( .A1(n14802), .A2(n14790), .B1(n14800), .B2(DATAI_18_), 
        .ZN(n14791) );
  OAI211_X1 U18274 ( .C1(n14794), .C2(n14793), .A(n14792), .B(n14791), .ZN(
        P1_U2886) );
  AOI22_X1 U18275 ( .A1(n14799), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14783), .ZN(n14797) );
  AOI22_X1 U18276 ( .A1(n14802), .A2(n14795), .B1(n14800), .B2(DATAI_17_), 
        .ZN(n14796) );
  OAI211_X1 U18277 ( .C1(n14798), .C2(n14793), .A(n14797), .B(n14796), .ZN(
        P1_U2887) );
  AOI22_X1 U18278 ( .A1(n14799), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n14783), .ZN(n14804) );
  AOI22_X1 U18279 ( .A1(n14802), .A2(n14801), .B1(n14800), .B2(DATAI_16_), 
        .ZN(n14803) );
  OAI211_X1 U18280 ( .C1(n14805), .C2(n14793), .A(n14804), .B(n14803), .ZN(
        P1_U2888) );
  MUX2_X1 U18281 ( .A(n16158), .B(n14807), .S(n14806), .Z(n14808) );
  XNOR2_X1 U18282 ( .A(n14808), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14991) );
  NAND2_X1 U18283 ( .A1(n16181), .A2(n14809), .ZN(n14810) );
  NAND2_X1 U18284 ( .A1(n16285), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14985) );
  OAI211_X1 U18285 ( .C1(n14811), .C2(n16187), .A(n14810), .B(n14985), .ZN(
        n14812) );
  AOI21_X1 U18286 ( .B1(n14813), .B2(n14887), .A(n14812), .ZN(n14814) );
  OAI21_X1 U18287 ( .B1(n14991), .B2(n20226), .A(n14814), .ZN(P1_U2970) );
  NAND2_X1 U18288 ( .A1(n16285), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14996) );
  OAI21_X1 U18289 ( .B1(n16187), .B2(n14815), .A(n14996), .ZN(n14816) );
  AOI21_X1 U18290 ( .B1(n14817), .B2(n16181), .A(n14816), .ZN(n14828) );
  NAND2_X1 U18291 ( .A1(n14847), .A2(n14818), .ZN(n14823) );
  AND2_X1 U18292 ( .A1(n14819), .A2(n15011), .ZN(n14820) );
  NAND2_X1 U18293 ( .A1(n15065), .A2(n15011), .ZN(n14821) );
  INV_X1 U18294 ( .A(n14823), .ZN(n14824) );
  MUX2_X1 U18295 ( .A(n16158), .B(n14824), .S(n15002), .Z(n14825) );
  NAND2_X1 U18296 ( .A1(n14831), .A2(n14825), .ZN(n14826) );
  XNOR2_X1 U18297 ( .A(n14826), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14992) );
  NAND2_X1 U18298 ( .A1(n14992), .A2(n16183), .ZN(n14827) );
  OAI211_X1 U18299 ( .C1(n14829), .C2(n16120), .A(n14828), .B(n14827), .ZN(
        P1_U2971) );
  NAND2_X1 U18300 ( .A1(n14831), .A2(n14830), .ZN(n14832) );
  XNOR2_X1 U18301 ( .A(n14832), .B(n15002), .ZN(n15009) );
  NOR2_X1 U18302 ( .A1(n16238), .A2(n20866), .ZN(n15001) );
  AOI21_X1 U18303 ( .B1(n16173), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15001), .ZN(n14833) );
  OAI21_X1 U18304 ( .B1(n16180), .B2(n14834), .A(n14833), .ZN(n14835) );
  AOI21_X1 U18305 ( .B1(n14836), .B2(n14887), .A(n14835), .ZN(n14837) );
  OAI21_X1 U18306 ( .B1(n20226), .B2(n15009), .A(n14837), .ZN(P1_U2972) );
  INV_X1 U18307 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14838) );
  NAND2_X1 U18308 ( .A1(n16285), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15013) );
  OAI21_X1 U18309 ( .B1(n16187), .B2(n14838), .A(n15013), .ZN(n14839) );
  AOI21_X1 U18310 ( .B1(n14840), .B2(n16181), .A(n14839), .ZN(n14844) );
  INV_X1 U18311 ( .A(n14830), .ZN(n14842) );
  NAND2_X1 U18312 ( .A1(n14842), .A2(n15011), .ZN(n15010) );
  NAND3_X1 U18313 ( .A1(n14841), .A2(n15010), .A3(n16183), .ZN(n14843) );
  OAI211_X1 U18314 ( .C1(n14845), .C2(n16120), .A(n14844), .B(n14843), .ZN(
        P1_U2973) );
  AOI21_X1 U18315 ( .B1(n14846), .B2(n15065), .A(n16197), .ZN(n14855) );
  MUX2_X1 U18316 ( .A(n16135), .B(n14855), .S(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .Z(n14848) );
  OAI211_X1 U18317 ( .C1(n16158), .C2(n16197), .A(n14848), .B(n14847), .ZN(
        n14849) );
  XOR2_X1 U18318 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n14849), .Z(
        n15029) );
  NAND2_X1 U18319 ( .A1(n16285), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n15023) );
  NAND2_X1 U18320 ( .A1(n16173), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14850) );
  OAI211_X1 U18321 ( .C1(n16180), .C2(n14851), .A(n15023), .B(n14850), .ZN(
        n14852) );
  AOI21_X1 U18322 ( .B1(n14853), .B2(n14887), .A(n14852), .ZN(n14854) );
  OAI21_X1 U18323 ( .B1(n20226), .B2(n15029), .A(n14854), .ZN(P1_U2974) );
  NOR2_X1 U18324 ( .A1(n9664), .A2(n15065), .ZN(n14856) );
  MUX2_X1 U18325 ( .A(n14856), .B(n16158), .S(n14855), .Z(n14857) );
  XNOR2_X1 U18326 ( .A(n14857), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15040) );
  NAND2_X1 U18327 ( .A1(n16285), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15034) );
  OAI21_X1 U18328 ( .B1(n16187), .B2(n14858), .A(n15034), .ZN(n14861) );
  NOR2_X1 U18329 ( .A1(n14859), .A2(n16120), .ZN(n14860) );
  AOI211_X1 U18330 ( .C1(n16181), .C2(n14862), .A(n14861), .B(n14860), .ZN(
        n14863) );
  OAI21_X1 U18331 ( .B1(n15040), .B2(n20226), .A(n14863), .ZN(P1_U2975) );
  XNOR2_X1 U18332 ( .A(n16158), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14864) );
  XNOR2_X1 U18333 ( .A(n9663), .B(n14864), .ZN(n16191) );
  AOI22_X1 U18334 ( .A1(n16173), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n16285), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n14865) );
  OAI21_X1 U18335 ( .B1(n16180), .B2(n14866), .A(n14865), .ZN(n14867) );
  AOI21_X1 U18336 ( .B1(n14868), .B2(n14887), .A(n14867), .ZN(n14869) );
  OAI21_X1 U18337 ( .B1(n16191), .B2(n20226), .A(n14869), .ZN(P1_U2976) );
  NAND2_X1 U18338 ( .A1(n14871), .A2(n14870), .ZN(n14872) );
  XOR2_X1 U18339 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n14872), .Z(
        n16200) );
  OAI22_X1 U18340 ( .A1(n16187), .A2(n14873), .B1(n16238), .B2(n21098), .ZN(
        n14876) );
  NOR2_X1 U18341 ( .A1(n14874), .A2(n16120), .ZN(n14875) );
  AOI211_X1 U18342 ( .C1(n16181), .C2(n14877), .A(n14876), .B(n14875), .ZN(
        n14878) );
  OAI21_X1 U18343 ( .B1(n20226), .B2(n16200), .A(n14878), .ZN(P1_U2977) );
  OR3_X1 U18344 ( .A1(n14879), .A2(n16135), .A3(n14954), .ZN(n14883) );
  NAND2_X1 U18345 ( .A1(n16135), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14880) );
  NAND2_X1 U18346 ( .A1(n14879), .A2(n14880), .ZN(n15052) );
  NAND2_X1 U18347 ( .A1(n16135), .A2(n14954), .ZN(n14881) );
  OAI21_X1 U18348 ( .B1(n15052), .B2(n14881), .A(n14883), .ZN(n14892) );
  NAND3_X1 U18349 ( .A1(n14892), .A2(n16135), .A3(n15044), .ZN(n14882) );
  OAI21_X1 U18350 ( .B1(n14883), .B2(n15044), .A(n14882), .ZN(n14884) );
  XNOR2_X1 U18351 ( .A(n14884), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15050) );
  NAND2_X1 U18352 ( .A1(n16285), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15046) );
  NAND2_X1 U18353 ( .A1(n16173), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14885) );
  OAI211_X1 U18354 ( .C1(n16180), .C2(n16061), .A(n15046), .B(n14885), .ZN(
        n14886) );
  AOI21_X1 U18355 ( .B1(n16059), .B2(n14887), .A(n14886), .ZN(n14888) );
  OAI21_X1 U18356 ( .B1(n15050), .B2(n20226), .A(n14888), .ZN(P1_U2978) );
  NOR2_X1 U18357 ( .A1(n16238), .A2(n21119), .ZN(n16025) );
  NOR2_X1 U18358 ( .A1(n16187), .A2(n14889), .ZN(n14890) );
  AOI211_X1 U18359 ( .C1(n16181), .C2(n14891), .A(n16025), .B(n14890), .ZN(
        n14894) );
  XNOR2_X1 U18360 ( .A(n14892), .B(n15044), .ZN(n16029) );
  NAND2_X1 U18361 ( .A1(n16029), .A2(n16183), .ZN(n14893) );
  OAI211_X1 U18362 ( .C1(n14895), .C2(n16120), .A(n14894), .B(n14893), .ZN(
        P1_U2979) );
  OAI21_X1 U18363 ( .B1(n14897), .B2(n14896), .A(n14879), .ZN(n16213) );
  AOI22_X1 U18364 ( .A1(n16173), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n16285), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14898) );
  OAI21_X1 U18365 ( .B1(n14899), .B2(n16180), .A(n14898), .ZN(n14900) );
  AOI21_X1 U18366 ( .B1(n14901), .B2(n14887), .A(n14900), .ZN(n14902) );
  OAI21_X1 U18367 ( .B1(n20226), .B2(n16213), .A(n14902), .ZN(P1_U2981) );
  NAND2_X1 U18368 ( .A1(n16135), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14919) );
  NAND2_X1 U18369 ( .A1(n16135), .A2(n14904), .ZN(n14915) );
  NAND3_X1 U18370 ( .A1(n14903), .A2(n14919), .A3(n14915), .ZN(n16131) );
  INV_X1 U18371 ( .A(n16131), .ZN(n14907) );
  OAI21_X1 U18372 ( .B1(n14907), .B2(n14906), .A(n14905), .ZN(n14909) );
  XNOR2_X1 U18373 ( .A(n15065), .B(n16233), .ZN(n14908) );
  XNOR2_X1 U18374 ( .A(n14909), .B(n14908), .ZN(n16231) );
  NAND2_X1 U18375 ( .A1(n16231), .A2(n16183), .ZN(n14913) );
  AND2_X1 U18376 ( .A1(n16285), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n16228) );
  NOR2_X1 U18377 ( .A1(n16180), .A2(n14910), .ZN(n14911) );
  AOI211_X1 U18378 ( .C1(n16173), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16228), .B(n14911), .ZN(n14912) );
  OAI211_X1 U18379 ( .C1(n16120), .C2(n14914), .A(n14913), .B(n14912), .ZN(
        P1_U2985) );
  INV_X1 U18380 ( .A(n14903), .ZN(n14918) );
  INV_X1 U18381 ( .A(n14915), .ZN(n14916) );
  AOI21_X1 U18382 ( .B1(n14918), .B2(n14917), .A(n14916), .ZN(n15089) );
  AND2_X1 U18383 ( .A1(n14919), .A2(n14920), .ZN(n15088) );
  NAND2_X1 U18384 ( .A1(n15089), .A2(n15088), .ZN(n15087) );
  NAND2_X1 U18385 ( .A1(n15087), .A2(n14920), .ZN(n14921) );
  XOR2_X1 U18386 ( .A(n14922), .B(n14921), .Z(n16242) );
  NAND2_X1 U18387 ( .A1(n16242), .A2(n16183), .ZN(n14926) );
  INV_X1 U18388 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14923) );
  OAI22_X1 U18389 ( .A1(n16187), .A2(n14923), .B1(n16238), .B2(n20844), .ZN(
        n14924) );
  AOI21_X1 U18390 ( .B1(n16096), .B2(n16181), .A(n14924), .ZN(n14925) );
  OAI211_X1 U18391 ( .C1(n16120), .C2(n16094), .A(n14926), .B(n14925), .ZN(
        P1_U2986) );
  MUX2_X1 U18392 ( .A(n14927), .B(n14903), .S(n16158), .Z(n14928) );
  XNOR2_X1 U18393 ( .A(n14928), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16257) );
  NAND2_X1 U18394 ( .A1(n16257), .A2(n16183), .ZN(n14932) );
  AND2_X1 U18395 ( .A1(n16285), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n16254) );
  NOR2_X1 U18396 ( .A1(n16180), .A2(n14929), .ZN(n14930) );
  AOI211_X1 U18397 ( .C1(n16173), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16254), .B(n14930), .ZN(n14931) );
  OAI211_X1 U18398 ( .C1(n16120), .C2(n14933), .A(n14932), .B(n14931), .ZN(
        P1_U2989) );
  INV_X1 U18399 ( .A(n14934), .ZN(n14948) );
  NAND3_X1 U18400 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n14935), .ZN(n15098) );
  INV_X1 U18401 ( .A(n15098), .ZN(n14936) );
  NAND2_X1 U18402 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14936), .ZN(
        n15095) );
  NOR2_X1 U18403 ( .A1(n14937), .A2(n15095), .ZN(n14939) );
  INV_X1 U18404 ( .A(n15097), .ZN(n14938) );
  NAND2_X1 U18405 ( .A1(n14939), .A2(n14938), .ZN(n15069) );
  INV_X1 U18406 ( .A(n15069), .ZN(n14949) );
  NAND2_X1 U18407 ( .A1(n14940), .A2(n14939), .ZN(n14950) );
  NAND3_X1 U18408 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14961), .A3(
        n14949), .ZN(n14941) );
  OAI21_X1 U18409 ( .B1(n14950), .B2(n15101), .A(n14941), .ZN(n15041) );
  AOI21_X1 U18410 ( .B1(n14963), .B2(n14949), .A(n15041), .ZN(n16246) );
  NOR2_X1 U18411 ( .A1(n16246), .A2(n16245), .ZN(n16190) );
  INV_X1 U18412 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16126) );
  NOR2_X1 U18413 ( .A1(n15084), .A2(n16126), .ZN(n16220) );
  NAND3_X1 U18414 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n16220), .ZN(n16211) );
  NOR2_X1 U18415 ( .A1(n16218), .A2(n16211), .ZN(n14951) );
  INV_X1 U18416 ( .A(n14951), .ZN(n14944) );
  INV_X1 U18417 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14942) );
  NOR3_X1 U18418 ( .A1(n14944), .A2(n14943), .A3(n14942), .ZN(n15030) );
  NAND2_X1 U18419 ( .A1(n16190), .A2(n15030), .ZN(n15033) );
  INV_X1 U18420 ( .A(n15012), .ZN(n14962) );
  NOR3_X1 U18421 ( .A1(n15033), .A2(n15011), .A3(n14962), .ZN(n15003) );
  NAND3_X1 U18422 ( .A1(n15003), .A2(n14984), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14975) );
  INV_X1 U18423 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14945) );
  NOR3_X1 U18424 ( .A1(n14975), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14945), .ZN(n14946) );
  AOI211_X1 U18425 ( .C1(n14948), .C2(n16286), .A(n14947), .B(n14946), .ZN(
        n14970) );
  AND2_X1 U18426 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14951), .ZN(
        n15042) );
  NAND2_X1 U18427 ( .A1(n14949), .A2(n15042), .ZN(n15055) );
  NOR2_X1 U18428 ( .A1(n16245), .A2(n14950), .ZN(n16234) );
  AOI21_X1 U18429 ( .B1(n16234), .B2(n14951), .A(n15101), .ZN(n14953) );
  AOI211_X1 U18430 ( .C1(n15096), .C2(n15055), .A(n14953), .B(n14952), .ZN(
        n15056) );
  NOR2_X1 U18431 ( .A1(n14954), .A2(n15044), .ZN(n14956) );
  AOI21_X1 U18432 ( .B1(n15056), .B2(n14956), .A(n14955), .ZN(n16199) );
  NAND2_X1 U18433 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16204) );
  INV_X1 U18434 ( .A(n16204), .ZN(n14957) );
  NOR2_X1 U18435 ( .A1(n16270), .A2(n14957), .ZN(n14958) );
  NOR2_X1 U18436 ( .A1(n16199), .A2(n14958), .ZN(n16198) );
  OR2_X1 U18437 ( .A1(n15101), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14959) );
  NAND2_X1 U18438 ( .A1(n16198), .A2(n14959), .ZN(n15031) );
  INV_X1 U18439 ( .A(n15018), .ZN(n14960) );
  AND2_X1 U18440 ( .A1(n14961), .A2(n14960), .ZN(n14966) );
  NAND2_X1 U18441 ( .A1(n14963), .A2(n14962), .ZN(n14964) );
  OAI21_X1 U18442 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15101), .A(
        n14964), .ZN(n14965) );
  INV_X1 U18443 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15017) );
  OR3_X1 U18444 ( .A1(n15027), .A2(n15017), .A3(n15011), .ZN(n14967) );
  AOI21_X1 U18445 ( .B1(n10062), .B2(n14968), .A(n15007), .ZN(n14981) );
  OAI211_X1 U18446 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16270), .A(
        n14981), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14976) );
  NAND3_X1 U18447 ( .A1(n14976), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14968), .ZN(n14969) );
  OAI211_X1 U18448 ( .C1(n14971), .C2(n16222), .A(n14970), .B(n14969), .ZN(
        P1_U3000) );
  INV_X1 U18449 ( .A(n14972), .ZN(n14973) );
  AOI21_X1 U18450 ( .B1(n14974), .B2(n16286), .A(n14973), .ZN(n14979) );
  INV_X1 U18451 ( .A(n14975), .ZN(n14977) );
  OAI21_X1 U18452 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14977), .A(
        n14976), .ZN(n14978) );
  OAI211_X1 U18453 ( .C1(n14980), .C2(n16222), .A(n14979), .B(n14978), .ZN(
        P1_U3001) );
  INV_X1 U18454 ( .A(n14981), .ZN(n14989) );
  INV_X1 U18455 ( .A(n14982), .ZN(n14987) );
  NAND3_X1 U18456 ( .A1(n15003), .A2(n14984), .A3(n14983), .ZN(n14986) );
  OAI211_X1 U18457 ( .C1(n14987), .C2(n16239), .A(n14986), .B(n14985), .ZN(
        n14988) );
  AOI21_X1 U18458 ( .B1(n14989), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14988), .ZN(n14990) );
  OAI21_X1 U18459 ( .B1(n14991), .B2(n16222), .A(n14990), .ZN(P1_U3002) );
  INV_X1 U18460 ( .A(n14992), .ZN(n15000) );
  INV_X1 U18461 ( .A(n14993), .ZN(n14994) );
  NAND3_X1 U18462 ( .A1(n15003), .A2(n14994), .A3(n10062), .ZN(n14995) );
  OAI211_X1 U18463 ( .C1(n14997), .C2(n16239), .A(n14996), .B(n14995), .ZN(
        n14998) );
  AOI21_X1 U18464 ( .B1(n15007), .B2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14998), .ZN(n14999) );
  OAI21_X1 U18465 ( .B1(n15000), .B2(n16222), .A(n14999), .ZN(P1_U3003) );
  AOI21_X1 U18466 ( .B1(n15003), .B2(n15002), .A(n15001), .ZN(n15004) );
  OAI21_X1 U18467 ( .B1(n15005), .B2(n16239), .A(n15004), .ZN(n15006) );
  AOI21_X1 U18468 ( .B1(n15007), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15006), .ZN(n15008) );
  OAI21_X1 U18469 ( .B1(n15009), .B2(n16222), .A(n15008), .ZN(P1_U3004) );
  NAND3_X1 U18470 ( .A1(n14841), .A2(n15010), .A3(n16289), .ZN(n15022) );
  NAND2_X1 U18471 ( .A1(n15012), .A2(n15011), .ZN(n15014) );
  OAI21_X1 U18472 ( .B1(n15033), .B2(n15014), .A(n15013), .ZN(n15015) );
  AOI21_X1 U18473 ( .B1(n15016), .B2(n16286), .A(n15015), .ZN(n15021) );
  NAND2_X1 U18474 ( .A1(n15018), .A2(n15017), .ZN(n15019) );
  NOR2_X1 U18475 ( .A1(n15033), .A2(n15019), .ZN(n15026) );
  OAI21_X1 U18476 ( .B1(n15027), .B2(n15026), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15020) );
  NAND3_X1 U18477 ( .A1(n15022), .A2(n15021), .A3(n15020), .ZN(P1_U3005) );
  OAI21_X1 U18478 ( .B1(n15024), .B2(n16239), .A(n15023), .ZN(n15025) );
  AOI211_X1 U18479 ( .C1(n15027), .C2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15026), .B(n15025), .ZN(n15028) );
  OAI21_X1 U18480 ( .B1(n15029), .B2(n16222), .A(n15028), .ZN(P1_U3006) );
  AND2_X1 U18481 ( .A1(n15030), .A2(n16197), .ZN(n16189) );
  AOI21_X1 U18482 ( .B1(n16189), .B2(n15103), .A(n15031), .ZN(n15032) );
  INV_X1 U18483 ( .A(n15032), .ZN(n15038) );
  NOR3_X1 U18484 ( .A1(n15033), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n16197), .ZN(n15037) );
  OAI21_X1 U18485 ( .B1(n15035), .B2(n16239), .A(n15034), .ZN(n15036) );
  AOI211_X1 U18486 ( .C1(n15038), .C2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15037), .B(n15036), .ZN(n15039) );
  OAI21_X1 U18487 ( .B1(n15040), .B2(n16222), .A(n15039), .ZN(P1_U3007) );
  NAND2_X1 U18488 ( .A1(n15042), .A2(n15041), .ZN(n15054) );
  OAI21_X1 U18489 ( .B1(n15055), .B2(n15053), .A(n15054), .ZN(n15043) );
  NAND2_X1 U18490 ( .A1(n15043), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16032) );
  NOR2_X1 U18491 ( .A1(n16032), .A2(n15044), .ZN(n16205) );
  NAND2_X1 U18492 ( .A1(n16205), .A2(n15045), .ZN(n15047) );
  OAI211_X1 U18493 ( .C1(n16239), .C2(n16057), .A(n15047), .B(n15046), .ZN(
        n15048) );
  AOI21_X1 U18494 ( .B1(n16199), .B2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15048), .ZN(n15049) );
  OAI21_X1 U18495 ( .B1(n15050), .B2(n16222), .A(n15049), .ZN(P1_U3010) );
  XNOR2_X1 U18496 ( .A(n15065), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15051) );
  XNOR2_X1 U18497 ( .A(n15052), .B(n15051), .ZN(n16119) );
  AOI21_X1 U18498 ( .B1(n15054), .B2(n15053), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16027) );
  NAND2_X1 U18499 ( .A1(n15055), .A2(n15054), .ZN(n15060) );
  INV_X1 U18500 ( .A(n16066), .ZN(n15058) );
  INV_X1 U18501 ( .A(n15056), .ZN(n16026) );
  AOI22_X1 U18502 ( .A1(n16285), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16026), .ZN(n15057) );
  OAI21_X1 U18503 ( .B1(n15058), .B2(n16239), .A(n15057), .ZN(n15059) );
  AOI21_X1 U18504 ( .B1(n16027), .B2(n15060), .A(n15059), .ZN(n15061) );
  OAI21_X1 U18505 ( .B1(n16119), .B2(n16222), .A(n15061), .ZN(P1_U3012) );
  INV_X1 U18506 ( .A(n16130), .ZN(n15064) );
  INV_X1 U18507 ( .A(n15062), .ZN(n15063) );
  OAI21_X1 U18508 ( .B1(n14903), .B2(n15064), .A(n15063), .ZN(n15080) );
  NOR2_X1 U18509 ( .A1(n15065), .A2(n15084), .ZN(n16129) );
  NOR2_X1 U18510 ( .A1(n15080), .A2(n16129), .ZN(n15066) );
  NOR2_X1 U18511 ( .A1(n15066), .A2(n15072), .ZN(n15068) );
  OAI22_X1 U18512 ( .A1(n15068), .A2(n15067), .B1(n15066), .B2(n16132), .ZN(
        n16147) );
  OAI21_X1 U18513 ( .B1(n16245), .B2(n15069), .A(n15096), .ZN(n15071) );
  OAI211_X1 U18514 ( .C1(n16234), .C2(n15101), .A(n15071), .B(n15070), .ZN(
        n16230) );
  INV_X1 U18515 ( .A(n16230), .ZN(n16244) );
  OAI21_X1 U18516 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16270), .A(
        n16244), .ZN(n15083) );
  INV_X1 U18517 ( .A(n16190), .ZN(n16210) );
  NOR2_X1 U18518 ( .A1(n16233), .A2(n16210), .ZN(n16219) );
  NOR2_X1 U18519 ( .A1(n15072), .A2(n16220), .ZN(n15073) );
  AOI22_X1 U18520 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n15083), .B1(
        n16219), .B2(n15073), .ZN(n15076) );
  AOI22_X1 U18521 ( .A1(n15074), .A2(n16286), .B1(n16285), .B2(
        P1_REIP_REG_16__SCAN_IN), .ZN(n15075) );
  OAI211_X1 U18522 ( .C1(n16147), .C2(n16222), .A(n15076), .B(n15075), .ZN(
        P1_U3015) );
  INV_X1 U18523 ( .A(n15077), .ZN(n15078) );
  NOR2_X1 U18524 ( .A1(n16129), .A2(n15078), .ZN(n15079) );
  XNOR2_X1 U18525 ( .A(n15080), .B(n15079), .ZN(n16152) );
  OAI22_X1 U18526 ( .A1(n15081), .A2(n16239), .B1(n20848), .B2(n16238), .ZN(
        n15082) );
  AOI21_X1 U18527 ( .B1(n15083), .B2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15082), .ZN(n15086) );
  NAND2_X1 U18528 ( .A1(n16219), .A2(n15084), .ZN(n15085) );
  OAI211_X1 U18529 ( .C1(n16152), .C2(n16222), .A(n15086), .B(n15085), .ZN(
        P1_U3016) );
  OAI21_X1 U18530 ( .B1(n15089), .B2(n15088), .A(n15087), .ZN(n15090) );
  INV_X1 U18531 ( .A(n15090), .ZN(n16157) );
  INV_X1 U18532 ( .A(n15091), .ZN(n15094) );
  AOI21_X1 U18533 ( .B1(n16105), .B2(n16106), .A(n15092), .ZN(n15093) );
  NOR2_X1 U18534 ( .A1(n15094), .A2(n15093), .ZN(n16114) );
  AOI22_X1 U18535 ( .A1(n16114), .A2(n16286), .B1(n16285), .B2(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15109) );
  NOR2_X1 U18536 ( .A1(n15095), .A2(n16287), .ZN(n15106) );
  NOR2_X1 U18537 ( .A1(n15098), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16247) );
  INV_X1 U18538 ( .A(n15095), .ZN(n15102) );
  OAI21_X1 U18539 ( .B1(n15098), .B2(n15097), .A(n15096), .ZN(n15099) );
  OAI211_X1 U18540 ( .C1(n15102), .C2(n15101), .A(n15100), .B(n15099), .ZN(
        n16249) );
  AOI21_X1 U18541 ( .B1(n15103), .B2(n16247), .A(n16249), .ZN(n15104) );
  INV_X1 U18542 ( .A(n15104), .ZN(n15105) );
  MUX2_X1 U18543 ( .A(n15106), .B(n15105), .S(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n15107) );
  INV_X1 U18544 ( .A(n15107), .ZN(n15108) );
  OAI211_X1 U18545 ( .C1(n16157), .C2(n16222), .A(n15109), .B(n15108), .ZN(
        P1_U3019) );
  OAI22_X1 U18546 ( .A1(n15112), .A2(n20614), .B1(n15111), .B2(n15110), .ZN(
        n15113) );
  AOI21_X1 U18547 ( .B1(n20671), .B2(n20696), .A(n15113), .ZN(n15115) );
  NAND2_X1 U18548 ( .A1(n20549), .A2(n20746), .ZN(n20546) );
  NAND3_X1 U18549 ( .A1(n15115), .A2(n15114), .A3(n20546), .ZN(n15116) );
  MUX2_X1 U18550 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n15116), .S(
        n20372), .Z(P1_U3475) );
  INV_X1 U18551 ( .A(n15117), .ZN(n15119) );
  AOI211_X1 U18552 ( .C1(n20616), .C2(n15976), .A(n15119), .B(n15118), .ZN(
        n15978) );
  INV_X1 U18553 ( .A(n15120), .ZN(n15123) );
  AOI21_X1 U18554 ( .B1(n15123), .B2(n15122), .A(n15121), .ZN(n15124) );
  OAI21_X1 U18555 ( .B1(n15978), .B2(n20897), .A(n15124), .ZN(n15125) );
  MUX2_X1 U18556 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15125), .S(
        n20892), .Z(P1_U3473) );
  NAND2_X1 U18557 ( .A1(n15126), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n15134) );
  INV_X1 U18558 ( .A(n15127), .ZN(n15129) );
  AOI22_X1 U18559 ( .A1(n20796), .A2(n15129), .B1(n20794), .B2(n15128), .ZN(
        n15133) );
  NAND2_X1 U18560 ( .A1(n20788), .A2(n20797), .ZN(n15132) );
  NAND2_X1 U18561 ( .A1(n15130), .A2(n20688), .ZN(n15131) );
  NAND4_X1 U18562 ( .A1(n15134), .A2(n15133), .A3(n15132), .A4(n15131), .ZN(
        P1_U3152) );
  OAI211_X1 U18563 ( .C1(n15137), .C2(n15136), .A(n19342), .B(n15135), .ZN(
        n15139) );
  AOI22_X1 U18564 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(n19361), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19366), .ZN(n15138) );
  NAND2_X1 U18565 ( .A1(n15139), .A2(n15138), .ZN(n15140) );
  AOI21_X1 U18566 ( .B1(n19360), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15140), .ZN(n15150) );
  OAI21_X1 U18567 ( .B1(n15143), .B2(n15141), .A(n15142), .ZN(n16510) );
  INV_X1 U18568 ( .A(n16510), .ZN(n15148) );
  OR2_X1 U18569 ( .A1(n15145), .A2(n15144), .ZN(n15147) );
  AND2_X1 U18570 ( .A1(n15147), .A2(n15146), .ZN(n16508) );
  AOI22_X1 U18571 ( .A1(n15148), .A2(n19389), .B1(n19305), .B2(n16508), .ZN(
        n15149) );
  OAI211_X1 U18572 ( .C1(n15151), .C2(n19362), .A(n15150), .B(n15149), .ZN(
        P2_U2832) );
  OAI211_X1 U18573 ( .C1(n15449), .C2(n15153), .A(n19342), .B(n15152), .ZN(
        n15165) );
  NAND2_X1 U18574 ( .A1(n15154), .A2(n9807), .ZN(n15156) );
  INV_X1 U18575 ( .A(n15141), .ZN(n15155) );
  NAND2_X1 U18576 ( .A1(n15156), .A2(n15155), .ZN(n15621) );
  INV_X1 U18577 ( .A(n15621), .ZN(n16394) );
  INV_X1 U18578 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n16397) );
  OR2_X1 U18579 ( .A1(n15158), .A2(n15157), .ZN(n15160) );
  INV_X1 U18580 ( .A(n15144), .ZN(n15159) );
  NAND2_X1 U18581 ( .A1(n15160), .A2(n15159), .ZN(n15618) );
  INV_X1 U18582 ( .A(n15618), .ZN(n15348) );
  NAND2_X1 U18583 ( .A1(n19305), .A2(n15348), .ZN(n15162) );
  AOI22_X1 U18584 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19360), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19366), .ZN(n15161) );
  OAI211_X1 U18585 ( .C1(n16397), .C2(n19382), .A(n15162), .B(n15161), .ZN(
        n15163) );
  AOI21_X1 U18586 ( .B1(n16394), .B2(n19389), .A(n15163), .ZN(n15164) );
  OAI211_X1 U18587 ( .C1(n15166), .C2(n19362), .A(n15165), .B(n15164), .ZN(
        P2_U2833) );
  INV_X1 U18588 ( .A(n15167), .ZN(n15180) );
  NAND2_X1 U18589 ( .A1(n13243), .A2(n15168), .ZN(n15169) );
  INV_X1 U18590 ( .A(n15169), .ZN(n19222) );
  INV_X1 U18591 ( .A(n15471), .ZN(n15170) );
  AOI221_X1 U18592 ( .B1(n15471), .B2(n19222), .C1(n15170), .C2(n15169), .A(
        n20071), .ZN(n15173) );
  INV_X1 U18593 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n15282) );
  OAI22_X1 U18594 ( .A1(n15171), .A2(n19391), .B1(n15282), .B2(n19382), .ZN(
        n15172) );
  AOI211_X1 U18595 ( .C1(n19366), .C2(P2_REIP_REG_21__SCAN_IN), .A(n15173), 
        .B(n15172), .ZN(n15179) );
  OAI21_X1 U18596 ( .B1(n15174), .B2(n15175), .A(n9807), .ZN(n16042) );
  INV_X1 U18597 ( .A(n16042), .ZN(n15177) );
  AOI21_X1 U18598 ( .B1(n15176), .B2(n15366), .A(n15157), .ZN(n16040) );
  AOI22_X1 U18599 ( .A1(n15177), .A2(n19389), .B1(n19305), .B2(n16040), .ZN(
        n15178) );
  OAI211_X1 U18600 ( .C1(n15180), .C2(n19362), .A(n15179), .B(n15178), .ZN(
        P2_U2834) );
  INV_X1 U18601 ( .A(n15181), .ZN(n15192) );
  NAND2_X1 U18602 ( .A1(n13243), .A2(n15182), .ZN(n15183) );
  XNOR2_X1 U18603 ( .A(n16479), .B(n15183), .ZN(n15184) );
  NAND2_X1 U18604 ( .A1(n15184), .A2(n19342), .ZN(n15191) );
  INV_X1 U18605 ( .A(n15751), .ZN(n16481) );
  NOR2_X1 U18606 ( .A1(n19387), .A2(n15185), .ZN(n15189) );
  AOI21_X1 U18607 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19360), .A(
        n19517), .ZN(n15187) );
  NAND2_X1 U18608 ( .A1(n19361), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n15186) );
  OAI211_X1 U18609 ( .C1(n15752), .C2(n19381), .A(n15187), .B(n15186), .ZN(
        n15188) );
  AOI211_X1 U18610 ( .C1(n16481), .C2(n19389), .A(n15189), .B(n15188), .ZN(
        n15190) );
  OAI211_X1 U18611 ( .C1(n19362), .C2(n15192), .A(n15191), .B(n15190), .ZN(
        P2_U2846) );
  NAND2_X1 U18612 ( .A1(n19299), .A2(n15193), .ZN(n15194) );
  XNOR2_X1 U18613 ( .A(n16493), .B(n15194), .ZN(n15195) );
  NAND2_X1 U18614 ( .A1(n15195), .A2(n19342), .ZN(n15203) );
  OAI21_X1 U18615 ( .B1(n15196), .B2(n19382), .A(n19324), .ZN(n15198) );
  NOR2_X1 U18616 ( .A1(n19387), .A2(n10760), .ZN(n15197) );
  AOI211_X1 U18617 ( .C1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n19360), .A(
        n15198), .B(n15197), .ZN(n15199) );
  OAI21_X1 U18618 ( .B1(n15200), .B2(n19362), .A(n15199), .ZN(n15201) );
  AOI21_X1 U18619 ( .B1(n16572), .B2(n19305), .A(n15201), .ZN(n15202) );
  OAI211_X1 U18620 ( .C1(n16503), .C2(n19354), .A(n15203), .B(n15202), .ZN(
        P2_U2850) );
  INV_X1 U18621 ( .A(n19393), .ZN(n15238) );
  NAND2_X1 U18622 ( .A1(n19299), .A2(n15204), .ZN(n15205) );
  XNOR2_X1 U18623 ( .A(n15206), .B(n15205), .ZN(n15207) );
  NAND2_X1 U18624 ( .A1(n15207), .A2(n19342), .ZN(n15213) );
  AOI22_X1 U18625 ( .A1(n19305), .A2(n20153), .B1(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n19360), .ZN(n15208) );
  OAI21_X1 U18626 ( .B1(n15209), .B2(n19362), .A(n15208), .ZN(n15211) );
  OAI22_X1 U18627 ( .A1(n10862), .A2(n19382), .B1(n14034), .B2(n19387), .ZN(
        n15210) );
  AOI211_X1 U18628 ( .C1(n19389), .C2(n15817), .A(n15211), .B(n15210), .ZN(
        n15212) );
  OAI211_X1 U18629 ( .C1(n15819), .C2(n15238), .A(n15213), .B(n15212), .ZN(
        P2_U2852) );
  NAND2_X1 U18630 ( .A1(n19366), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n15215) );
  AOI22_X1 U18631 ( .A1(n19361), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19360), .ZN(n15214) );
  OAI211_X1 U18632 ( .C1(n19362), .C2(n15216), .A(n15215), .B(n15214), .ZN(
        n15217) );
  AOI21_X1 U18633 ( .B1(n20161), .B2(n19305), .A(n15217), .ZN(n15218) );
  OAI21_X1 U18634 ( .B1(n19541), .B2(n19354), .A(n15218), .ZN(n15224) );
  INV_X1 U18635 ( .A(n15221), .ZN(n15222) );
  NOR2_X1 U18636 ( .A1(n19372), .A2(n15219), .ZN(n15226) );
  INV_X1 U18637 ( .A(n15226), .ZN(n15220) );
  AOI221_X1 U18638 ( .B1(n15222), .B2(n15226), .C1(n15221), .C2(n15220), .A(
        n20071), .ZN(n15223) );
  AOI211_X1 U18639 ( .C1(n15796), .C2(n19393), .A(n15224), .B(n15223), .ZN(
        n15225) );
  INV_X1 U18640 ( .A(n15225), .ZN(P2_U2853) );
  OAI21_X1 U18641 ( .B1(n19398), .B2(n15227), .A(n15226), .ZN(n15779) );
  OAI21_X1 U18642 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19299), .A(
        n15779), .ZN(n15228) );
  NAND2_X1 U18643 ( .A1(n15228), .A2(n19342), .ZN(n15237) );
  NAND2_X1 U18644 ( .A1(n20171), .A2(n19305), .ZN(n15233) );
  OAI22_X1 U18645 ( .A1(n15230), .A2(n19382), .B1(n10673), .B2(n19387), .ZN(
        n15231) );
  AOI21_X1 U18646 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19360), .A(
        n15231), .ZN(n15232) );
  OAI211_X1 U18647 ( .C1(n19362), .C2(n15234), .A(n15233), .B(n15232), .ZN(
        n15235) );
  AOI21_X1 U18648 ( .B1(n19559), .B2(n19389), .A(n15235), .ZN(n15236) );
  OAI211_X1 U18649 ( .C1(n15238), .C2(n20166), .A(n15237), .B(n15236), .ZN(
        P2_U2854) );
  OR2_X1 U18650 ( .A1(n9786), .A2(n15239), .ZN(n15240) );
  NAND2_X1 U18651 ( .A1(n15241), .A2(n15240), .ZN(n16315) );
  INV_X1 U18652 ( .A(n15242), .ZN(n15292) );
  NAND2_X1 U18653 ( .A1(n15243), .A2(n15244), .ZN(n15291) );
  NAND3_X1 U18654 ( .A1(n15292), .A2(n19411), .A3(n15291), .ZN(n15246) );
  NAND2_X1 U18655 ( .A1(n16392), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15245) );
  OAI211_X1 U18656 ( .C1(n16392), .C2(n16315), .A(n15246), .B(n15245), .ZN(
        P2_U2858) );
  NAND2_X1 U18657 ( .A1(n15247), .A2(n15248), .ZN(n15250) );
  XNOR2_X1 U18658 ( .A(n15250), .B(n15249), .ZN(n15314) );
  AND2_X1 U18659 ( .A1(n15262), .A2(n15251), .ZN(n15252) );
  OR2_X1 U18660 ( .A1(n9786), .A2(n15252), .ZN(n16328) );
  NOR2_X1 U18661 ( .A1(n16328), .A2(n16392), .ZN(n15253) );
  AOI21_X1 U18662 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n16392), .A(n15253), .ZN(
        n15254) );
  OAI21_X1 U18663 ( .B1(n15314), .B2(n19403), .A(n15254), .ZN(P2_U2859) );
  AOI21_X1 U18664 ( .B1(n15255), .B2(n15257), .A(n15256), .ZN(n15258) );
  INV_X1 U18665 ( .A(n15258), .ZN(n15321) );
  OR2_X1 U18666 ( .A1(n15259), .A2(n15260), .ZN(n15261) );
  NAND2_X1 U18667 ( .A1(n15262), .A2(n15261), .ZN(n16339) );
  NOR2_X1 U18668 ( .A1(n16339), .A2(n16392), .ZN(n15263) );
  AOI21_X1 U18669 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n16392), .A(n15263), .ZN(
        n15264) );
  OAI21_X1 U18670 ( .B1(n15321), .B2(n19403), .A(n15264), .ZN(P2_U2860) );
  INV_X1 U18671 ( .A(n15259), .ZN(n15265) );
  OAI21_X1 U18672 ( .B1(n15277), .B2(n15266), .A(n15265), .ZN(n16349) );
  NAND2_X1 U18673 ( .A1(n15322), .A2(n19411), .ZN(n15271) );
  NAND2_X1 U18674 ( .A1(n16392), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15270) );
  OAI211_X1 U18675 ( .C1(n16349), .C2(n16392), .A(n15271), .B(n15270), .ZN(
        P2_U2861) );
  NAND2_X1 U18676 ( .A1(n15274), .A2(n15273), .ZN(n15343) );
  NAND2_X1 U18677 ( .A1(n16392), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n15279) );
  AND2_X1 U18678 ( .A1(n15430), .A2(n15275), .ZN(n15276) );
  NOR2_X1 U18679 ( .A1(n15277), .A2(n15276), .ZN(n16420) );
  NAND2_X1 U18680 ( .A1(n16420), .A2(n19406), .ZN(n15278) );
  OAI211_X1 U18681 ( .C1(n15343), .C2(n19403), .A(n15279), .B(n15278), .ZN(
        P2_U2862) );
  OAI21_X1 U18682 ( .B1(n9792), .B2(n15281), .A(n15280), .ZN(n15361) );
  MUX2_X1 U18683 ( .A(n15282), .B(n16042), .S(n19415), .Z(n15283) );
  OAI21_X1 U18684 ( .B1(n15361), .B2(n19403), .A(n15283), .ZN(P2_U2866) );
  NAND2_X1 U18685 ( .A1(n15285), .A2(n15286), .ZN(n15287) );
  NAND2_X1 U18686 ( .A1(n15284), .A2(n15287), .ZN(n19236) );
  NOR2_X1 U18687 ( .A1(n19236), .A2(n16392), .ZN(n15288) );
  AOI21_X1 U18688 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n16392), .A(n15288), .ZN(
        n15289) );
  OAI21_X1 U18689 ( .B1(n15290), .B2(n19403), .A(n15289), .ZN(P2_U2868) );
  NAND3_X1 U18690 ( .A1(n15292), .A2(n16413), .A3(n15291), .ZN(n15304) );
  INV_X1 U18691 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16739) );
  OR2_X1 U18692 ( .A1(n15293), .A2(n16739), .ZN(n15295) );
  NAND2_X1 U18693 ( .A1(n15293), .A2(BUF2_REG_13__SCAN_IN), .ZN(n15294) );
  NAND2_X1 U18694 ( .A1(n15295), .A2(n15294), .ZN(n19479) );
  NOR2_X1 U18695 ( .A1(n15296), .A2(n15297), .ZN(n15298) );
  INV_X1 U18696 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n15300) );
  OAI22_X1 U18697 ( .A1(n15338), .A2(n16314), .B1(n19428), .B2(n15300), .ZN(
        n15301) );
  AOI21_X1 U18698 ( .B1(n16412), .B2(n19479), .A(n15301), .ZN(n15303) );
  AOI22_X1 U18699 ( .A1(n19418), .A2(BUF2_REG_29__SCAN_IN), .B1(n19419), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n15302) );
  NAND3_X1 U18700 ( .A1(n15304), .A2(n15303), .A3(n15302), .ZN(P2_U2890) );
  INV_X1 U18701 ( .A(n15305), .ZN(n15317) );
  AND2_X1 U18702 ( .A1(n15317), .A2(n15306), .ZN(n15307) );
  INV_X1 U18703 ( .A(n16336), .ZN(n15311) );
  OAI22_X1 U18704 ( .A1(n15369), .A2(n15309), .B1(n19428), .B2(n15308), .ZN(
        n15310) );
  AOI21_X1 U18705 ( .B1(n19417), .B2(n15311), .A(n15310), .ZN(n15313) );
  AOI22_X1 U18706 ( .A1(n19418), .A2(BUF2_REG_28__SCAN_IN), .B1(n19419), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15312) );
  OAI211_X1 U18707 ( .C1(n15314), .C2(n15373), .A(n15313), .B(n15312), .ZN(
        P2_U2891) );
  NAND2_X1 U18708 ( .A1(n15326), .A2(n15315), .ZN(n15316) );
  NAND2_X1 U18709 ( .A1(n15317), .A2(n15316), .ZN(n16338) );
  OAI22_X1 U18710 ( .A1(n15338), .A2(n16338), .B1(n19428), .B2(n13404), .ZN(
        n15318) );
  AOI21_X1 U18711 ( .B1(n16412), .B2(n19429), .A(n15318), .ZN(n15320) );
  AOI22_X1 U18712 ( .A1(n19418), .A2(BUF2_REG_27__SCAN_IN), .B1(n19419), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15319) );
  OAI211_X1 U18713 ( .C1(n15321), .C2(n15373), .A(n15320), .B(n15319), .ZN(
        P2_U2892) );
  NAND2_X1 U18714 ( .A1(n15322), .A2(n16413), .ZN(n15331) );
  OR2_X1 U18715 ( .A1(n15335), .A2(n15324), .ZN(n15325) );
  AND2_X1 U18716 ( .A1(n15326), .A2(n15325), .ZN(n16350) );
  AOI22_X1 U18717 ( .A1(n19417), .A2(n16350), .B1(n19432), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15330) );
  AOI22_X1 U18718 ( .A1(n19418), .A2(BUF2_REG_26__SCAN_IN), .B1(n19419), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15329) );
  NAND2_X1 U18719 ( .A1(n16412), .A2(n15327), .ZN(n15328) );
  NAND4_X1 U18720 ( .A1(n15331), .A2(n15330), .A3(n15329), .A4(n15328), .ZN(
        P2_U2893) );
  AND2_X1 U18721 ( .A1(n15333), .A2(n15332), .ZN(n15334) );
  NOR2_X1 U18722 ( .A1(n15335), .A2(n15334), .ZN(n16360) );
  INV_X1 U18723 ( .A(n16360), .ZN(n15337) );
  OAI22_X1 U18724 ( .A1(n15338), .A2(n15337), .B1(n19428), .B2(n15336), .ZN(
        n15339) );
  AOI21_X1 U18725 ( .B1(n16412), .B2(n15340), .A(n15339), .ZN(n15342) );
  AOI22_X1 U18726 ( .A1(n19418), .A2(BUF2_REG_25__SCAN_IN), .B1(n19419), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15341) );
  OAI211_X1 U18727 ( .C1(n15343), .C2(n15373), .A(n15342), .B(n15341), .ZN(
        P2_U2894) );
  AOI21_X1 U18728 ( .B1(n15345), .B2(n15280), .A(n15344), .ZN(n16395) );
  INV_X1 U18729 ( .A(n16395), .ZN(n15351) );
  OAI22_X1 U18730 ( .A1(n15369), .A2(n19579), .B1(n15346), .B2(n19428), .ZN(
        n15347) );
  AOI21_X1 U18731 ( .B1(n19417), .B2(n15348), .A(n15347), .ZN(n15350) );
  AOI22_X1 U18732 ( .A1(n19418), .A2(BUF2_REG_22__SCAN_IN), .B1(n19419), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n15349) );
  OAI211_X1 U18733 ( .C1(n15351), .C2(n15373), .A(n15350), .B(n15349), .ZN(
        P2_U2897) );
  OAI22_X1 U18734 ( .A1(n15369), .A2(n15353), .B1(n15352), .B2(n19428), .ZN(
        n15359) );
  INV_X1 U18735 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n15356) );
  INV_X1 U18736 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n15354) );
  OAI22_X1 U18737 ( .A1(n15357), .A2(n15356), .B1(n15355), .B2(n15354), .ZN(
        n15358) );
  AOI211_X1 U18738 ( .C1(n19417), .C2(n16040), .A(n15359), .B(n15358), .ZN(
        n15360) );
  OAI21_X1 U18739 ( .B1(n15361), .B2(n15373), .A(n15360), .ZN(P2_U2898) );
  AOI21_X1 U18740 ( .B1(n15363), .B2(n15362), .A(n9792), .ZN(n16399) );
  INV_X1 U18741 ( .A(n16399), .ZN(n15374) );
  OR2_X1 U18742 ( .A1(n15365), .A2(n15364), .ZN(n15367) );
  AND2_X1 U18743 ( .A1(n15367), .A2(n15366), .ZN(n19215) );
  OAI22_X1 U18744 ( .A1(n15369), .A2(n19574), .B1(n15368), .B2(n19428), .ZN(
        n15370) );
  AOI21_X1 U18745 ( .B1(n19417), .B2(n19215), .A(n15370), .ZN(n15372) );
  AOI22_X1 U18746 ( .A1(n19418), .A2(BUF2_REG_20__SCAN_IN), .B1(n19419), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n15371) );
  OAI211_X1 U18747 ( .C1(n15374), .C2(n15373), .A(n15372), .B(n15371), .ZN(
        P2_U2899) );
  NAND2_X1 U18748 ( .A1(n15376), .A2(n15375), .ZN(n15378) );
  XOR2_X1 U18749 ( .A(n15378), .B(n15377), .Z(n15558) );
  NOR2_X1 U18750 ( .A1(n16315), .A2(n16436), .ZN(n15381) );
  NAND2_X1 U18751 ( .A1(n19517), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15552) );
  OAI21_X1 U18752 ( .B1(n16506), .B2(n15379), .A(n15552), .ZN(n15380) );
  AOI211_X1 U18753 ( .C1(n15382), .C2(n16494), .A(n15381), .B(n15380), .ZN(
        n15385) );
  AOI21_X1 U18754 ( .B1(n15550), .B2(n15399), .A(n15383), .ZN(n15555) );
  NAND2_X1 U18755 ( .A1(n15555), .A2(n19507), .ZN(n15384) );
  OAI211_X1 U18756 ( .C1(n15558), .C2(n19510), .A(n15385), .B(n15384), .ZN(
        P2_U2985) );
  INV_X1 U18757 ( .A(n15391), .ZN(n15386) );
  INV_X1 U18758 ( .A(n15388), .ZN(n15389) );
  NAND2_X1 U18759 ( .A1(n9782), .A2(n15389), .ZN(n15405) );
  INV_X1 U18760 ( .A(n15405), .ZN(n15390) );
  NOR2_X1 U18761 ( .A1(n15392), .A2(n15391), .ZN(n15394) );
  XNOR2_X1 U18762 ( .A(n15396), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15397) );
  XNOR2_X1 U18763 ( .A(n15398), .B(n15397), .ZN(n15569) );
  NAND2_X1 U18764 ( .A1(n15409), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15578) );
  INV_X1 U18765 ( .A(n15399), .ZN(n15400) );
  AOI21_X1 U18766 ( .B1(n12245), .B2(n15578), .A(n15400), .ZN(n15566) );
  NOR2_X1 U18767 ( .A1(n16333), .A2(n19501), .ZN(n15403) );
  NAND2_X1 U18768 ( .A1(n19517), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15562) );
  NAND2_X1 U18769 ( .A1(n19503), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15401) );
  OAI211_X1 U18770 ( .C1(n16328), .C2(n16436), .A(n15562), .B(n15401), .ZN(
        n15402) );
  AOI211_X1 U18771 ( .C1(n15566), .C2(n19507), .A(n15403), .B(n15402), .ZN(
        n15404) );
  OAI21_X1 U18772 ( .B1(n15569), .B2(n19510), .A(n15404), .ZN(P2_U2986) );
  NAND2_X1 U18773 ( .A1(n15405), .A2(n12246), .ZN(n15570) );
  NAND3_X1 U18774 ( .A1(n15571), .A2(n12279), .A3(n15570), .ZN(n15412) );
  NAND2_X1 U18775 ( .A1(n19517), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15574) );
  NAND2_X1 U18776 ( .A1(n19503), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15406) );
  OAI211_X1 U18777 ( .C1(n16339), .C2(n16436), .A(n15574), .B(n15406), .ZN(
        n15407) );
  AOI21_X1 U18778 ( .B1(n15408), .B2(n16494), .A(n15407), .ZN(n15411) );
  INV_X1 U18779 ( .A(n15409), .ZN(n15415) );
  NAND2_X1 U18780 ( .A1(n15415), .A2(n12246), .ZN(n15579) );
  NAND3_X1 U18781 ( .A1(n15579), .A2(n19507), .A3(n15578), .ZN(n15410) );
  NAND3_X1 U18782 ( .A1(n15412), .A2(n15411), .A3(n15410), .ZN(P2_U2987) );
  OAI21_X1 U18783 ( .B1(n15413), .B2(n15604), .A(n15588), .ZN(n15414) );
  NAND2_X1 U18784 ( .A1(n15415), .A2(n15414), .ZN(n15594) );
  NAND2_X1 U18785 ( .A1(n15416), .A2(n15595), .ZN(n15418) );
  MUX2_X1 U18786 ( .A(n15595), .B(n15418), .S(n15417), .Z(n15420) );
  AND2_X1 U18787 ( .A1(n15420), .A2(n15419), .ZN(n15591) );
  NOR2_X1 U18788 ( .A1(n19324), .A2(n20124), .ZN(n15583) );
  NOR2_X1 U18789 ( .A1(n16349), .A2(n16436), .ZN(n15421) );
  AOI211_X1 U18790 ( .C1(n19503), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15583), .B(n15421), .ZN(n15422) );
  OAI21_X1 U18791 ( .B1(n16354), .B2(n19501), .A(n15422), .ZN(n15423) );
  AOI21_X1 U18792 ( .B1(n15591), .B2(n12279), .A(n15423), .ZN(n15424) );
  OAI21_X1 U18793 ( .B1(n15594), .B2(n19495), .A(n15424), .ZN(P2_U2988) );
  OAI21_X1 U18794 ( .B1(n9727), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15413), .ZN(n15617) );
  XNOR2_X1 U18795 ( .A(n15425), .B(n15610), .ZN(n15426) );
  XNOR2_X1 U18796 ( .A(n15427), .B(n15426), .ZN(n15615) );
  OAI22_X1 U18797 ( .A1(n10820), .A2(n19324), .B1(n19501), .B2(n16371), .ZN(
        n15432) );
  NAND2_X1 U18798 ( .A1(n15142), .A2(n15428), .ZN(n15429) );
  NAND2_X1 U18799 ( .A1(n15430), .A2(n15429), .ZN(n16386) );
  OAI22_X1 U18800 ( .A1(n16386), .A2(n16436), .B1(n9967), .B2(n16506), .ZN(
        n15431) );
  AOI211_X1 U18801 ( .C1(n15615), .C2(n12279), .A(n15432), .B(n15431), .ZN(
        n15433) );
  OAI21_X1 U18802 ( .B1(n15617), .B2(n19495), .A(n15433), .ZN(P2_U2990) );
  XNOR2_X1 U18803 ( .A(n15434), .B(n15435), .ZN(n16511) );
  AOI21_X1 U18804 ( .B1(n15436), .B2(n15444), .A(n9727), .ZN(n16513) );
  NAND2_X1 U18805 ( .A1(n16513), .A2(n19507), .ZN(n15442) );
  OAI22_X1 U18806 ( .A1(n15437), .A2(n16506), .B1(n10662), .B2(n19324), .ZN(
        n15439) );
  NOR2_X1 U18807 ( .A1(n16510), .A2(n16436), .ZN(n15438) );
  AOI211_X1 U18808 ( .C1(n15440), .C2(n16494), .A(n15439), .B(n15438), .ZN(
        n15441) );
  OAI211_X1 U18809 ( .C1(n16511), .C2(n19510), .A(n15442), .B(n15441), .ZN(
        P2_U2991) );
  OAI21_X1 U18810 ( .B1(n15443), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15444), .ZN(n15627) );
  NAND2_X1 U18811 ( .A1(n15447), .A2(n15446), .ZN(n15448) );
  XNOR2_X1 U18812 ( .A(n15445), .B(n15448), .ZN(n15624) );
  OAI22_X1 U18813 ( .A1(n10816), .A2(n19324), .B1(n19501), .B2(n15449), .ZN(
        n15452) );
  INV_X1 U18814 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15450) );
  OAI22_X1 U18815 ( .A1(n15621), .A2(n16436), .B1(n16506), .B2(n15450), .ZN(
        n15451) );
  AOI211_X1 U18816 ( .C1(n15624), .C2(n12279), .A(n15452), .B(n15451), .ZN(
        n15453) );
  OAI21_X1 U18817 ( .B1(n15627), .B2(n19495), .A(n15453), .ZN(P2_U2992) );
  INV_X1 U18818 ( .A(n16449), .ZN(n15699) );
  OAI211_X1 U18819 ( .C1(n15699), .C2(n15455), .A(n15702), .B(n16448), .ZN(
        n15458) );
  INV_X1 U18820 ( .A(n15456), .ZN(n15457) );
  NAND2_X1 U18821 ( .A1(n15458), .A2(n15457), .ZN(n15460) );
  OAI21_X1 U18822 ( .B1(n15529), .B2(n15527), .A(n15461), .ZN(n15512) );
  NAND2_X1 U18823 ( .A1(n15463), .A2(n15462), .ZN(n15513) );
  AOI21_X1 U18824 ( .B1(n15478), .B2(n15482), .A(n15479), .ZN(n15468) );
  NAND2_X1 U18825 ( .A1(n15466), .A2(n15465), .ZN(n15467) );
  XNOR2_X1 U18826 ( .A(n15468), .B(n15467), .ZN(n16045) );
  INV_X1 U18827 ( .A(n16045), .ZN(n15475) );
  INV_X1 U18828 ( .A(n15469), .ZN(n15476) );
  AOI21_X1 U18829 ( .B1(n15470), .B2(n15476), .A(n15443), .ZN(n16041) );
  AOI22_X1 U18830 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n19503), .B1(
        n16494), .B2(n15471), .ZN(n15472) );
  NAND2_X1 U18831 ( .A1(P2_REIP_REG_21__SCAN_IN), .A2(n19517), .ZN(n16049) );
  OAI211_X1 U18832 ( .C1(n16042), .C2(n16436), .A(n15472), .B(n16049), .ZN(
        n15473) );
  AOI21_X1 U18833 ( .B1(n16041), .B2(n19507), .A(n15473), .ZN(n15474) );
  OAI21_X1 U18834 ( .B1(n15475), .B2(n19510), .A(n15474), .ZN(P2_U2993) );
  INV_X1 U18835 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16535) );
  AND2_X2 U18836 ( .A1(n16446), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15691) );
  INV_X1 U18837 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15652) );
  OAI21_X1 U18838 ( .B1(n15498), .B2(n15652), .A(n15636), .ZN(n15477) );
  NAND2_X1 U18839 ( .A1(n15477), .A2(n15476), .ZN(n15647) );
  INV_X1 U18840 ( .A(n15478), .ZN(n15480) );
  NOR2_X1 U18841 ( .A1(n15480), .A2(n15479), .ZN(n15481) );
  XNOR2_X1 U18842 ( .A(n15482), .B(n15481), .ZN(n15644) );
  AND2_X1 U18843 ( .A1(n19517), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15638) );
  AND2_X1 U18844 ( .A1(n15284), .A2(n15483), .ZN(n15484) );
  OR2_X1 U18845 ( .A1(n15484), .A2(n15174), .ZN(n19214) );
  NOR2_X1 U18846 ( .A1(n19214), .A2(n16436), .ZN(n15485) );
  AOI211_X1 U18847 ( .C1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n19503), .A(
        n15638), .B(n15485), .ZN(n15486) );
  OAI21_X1 U18848 ( .B1(n19226), .B2(n19501), .A(n15486), .ZN(n15487) );
  AOI21_X1 U18849 ( .B1(n15644), .B2(n12279), .A(n15487), .ZN(n15488) );
  OAI21_X1 U18850 ( .B1(n15647), .B2(n19495), .A(n15488), .ZN(P2_U2994) );
  XOR2_X1 U18851 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n15498), .Z(
        n15656) );
  NOR2_X1 U18852 ( .A1(n10039), .A2(n15490), .ZN(n15492) );
  XOR2_X1 U18853 ( .A(n15492), .B(n15491), .Z(n15654) );
  OAI22_X1 U18854 ( .A1(n16506), .A2(n19230), .B1(n15493), .B2(n19324), .ZN(
        n15494) );
  AOI21_X1 U18855 ( .B1(n19229), .B2(n16494), .A(n15494), .ZN(n15495) );
  OAI21_X1 U18856 ( .B1(n19236), .B2(n16436), .A(n15495), .ZN(n15496) );
  AOI21_X1 U18857 ( .B1(n15654), .B2(n12279), .A(n15496), .ZN(n15497) );
  OAI21_X1 U18858 ( .B1(n15656), .B2(n19495), .A(n15497), .ZN(P2_U2995) );
  NOR2_X1 U18859 ( .A1(n15668), .A2(n15679), .ZN(n15499) );
  OAI21_X1 U18860 ( .B1(n15499), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15498), .ZN(n15667) );
  NOR2_X1 U18861 ( .A1(n10038), .A2(n15501), .ZN(n15502) );
  XNOR2_X1 U18862 ( .A(n15503), .B(n15502), .ZN(n15662) );
  INV_X1 U18863 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20112) );
  OAI22_X1 U18864 ( .A1(n20112), .A2(n19324), .B1(n19501), .B2(n19246), .ZN(
        n15508) );
  OR2_X1 U18865 ( .A1(n15505), .A2(n15504), .ZN(n15506) );
  NAND2_X1 U18866 ( .A1(n15285), .A2(n15506), .ZN(n16402) );
  OAI22_X1 U18867 ( .A1(n16402), .A2(n16436), .B1(n16506), .B2(n9970), .ZN(
        n15507) );
  AOI211_X1 U18868 ( .C1(n15662), .C2(n12279), .A(n15508), .B(n15507), .ZN(
        n15509) );
  OAI21_X1 U18869 ( .B1(n15667), .B2(n19495), .A(n15509), .ZN(P2_U2996) );
  INV_X1 U18870 ( .A(n15510), .ZN(n15511) );
  AOI21_X1 U18871 ( .B1(n15513), .B2(n15512), .A(n15511), .ZN(n15674) );
  XNOR2_X1 U18872 ( .A(n15514), .B(n15679), .ZN(n15515) );
  NAND2_X1 U18873 ( .A1(n15515), .A2(n19507), .ZN(n15521) );
  OAI22_X1 U18874 ( .A1(n16506), .A2(n15516), .B1(n15672), .B2(n19324), .ZN(
        n15519) );
  INV_X1 U18875 ( .A(n15517), .ZN(n19258) );
  NOR2_X1 U18876 ( .A1(n19258), .A2(n19501), .ZN(n15518) );
  AOI211_X1 U18877 ( .C1(n19512), .C2(n19255), .A(n15519), .B(n15518), .ZN(
        n15520) );
  OAI211_X1 U18878 ( .C1(n15674), .C2(n19510), .A(n15521), .B(n15520), .ZN(
        P2_U2997) );
  XNOR2_X1 U18879 ( .A(n16435), .B(n15671), .ZN(n15532) );
  NAND2_X1 U18880 ( .A1(n14293), .A2(n15522), .ZN(n15523) );
  NAND2_X1 U18881 ( .A1(n15524), .A2(n15523), .ZN(n15683) );
  NOR2_X1 U18882 ( .A1(n15684), .A2(n19324), .ZN(n15526) );
  INV_X1 U18883 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n19264) );
  OAI22_X1 U18884 ( .A1(n19264), .A2(n16506), .B1(n19501), .B2(n19269), .ZN(
        n15525) );
  AOI211_X1 U18885 ( .C1(n19512), .C2(n19400), .A(n15526), .B(n15525), .ZN(
        n15531) );
  INV_X1 U18886 ( .A(n15527), .ZN(n15528) );
  XNOR2_X1 U18887 ( .A(n15529), .B(n15528), .ZN(n15687) );
  NAND2_X1 U18888 ( .A1(n15687), .A2(n12279), .ZN(n15530) );
  OAI211_X1 U18889 ( .C1(n15532), .C2(n19495), .A(n15531), .B(n15530), .ZN(
        P2_U2998) );
  OAI21_X1 U18890 ( .B1(n15535), .B2(n15534), .A(n15533), .ZN(n16566) );
  INV_X1 U18891 ( .A(n14344), .ZN(n15538) );
  OAI21_X1 U18892 ( .B1(n15538), .B2(n15537), .A(n15536), .ZN(n15759) );
  AOI21_X1 U18893 ( .B1(n15759), .B2(n15756), .A(n10032), .ZN(n15542) );
  NAND2_X1 U18894 ( .A1(n15540), .A2(n15539), .ZN(n15541) );
  XNOR2_X1 U18895 ( .A(n15542), .B(n15541), .ZN(n16570) );
  INV_X1 U18896 ( .A(n16570), .ZN(n15546) );
  OAI22_X1 U18897 ( .A1(n10767), .A2(n19350), .B1(n19501), .B2(n19339), .ZN(
        n15545) );
  OAI22_X1 U18898 ( .A1(n15543), .A2(n16436), .B1(n16506), .B2(n19334), .ZN(
        n15544) );
  AOI211_X1 U18899 ( .C1(n15546), .C2(n12279), .A(n15545), .B(n15544), .ZN(
        n15547) );
  OAI21_X1 U18900 ( .B1(n19495), .B2(n16566), .A(n15547), .ZN(P2_U3006) );
  INV_X1 U18901 ( .A(n15577), .ZN(n15548) );
  OAI21_X1 U18902 ( .B1(n15559), .B2(n15549), .A(n15548), .ZN(n15565) );
  NOR2_X1 U18903 ( .A1(n19554), .A2(n16314), .ZN(n15554) );
  INV_X1 U18904 ( .A(n15549), .ZN(n15572) );
  NAND3_X1 U18905 ( .A1(n15572), .A2(n15559), .A3(n15550), .ZN(n15551) );
  OAI211_X1 U18906 ( .C1(n16315), .C2(n19540), .A(n15552), .B(n15551), .ZN(
        n15553) );
  AOI211_X1 U18907 ( .C1(n15565), .C2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15554), .B(n15553), .ZN(n15557) );
  NAND2_X1 U18908 ( .A1(n15555), .A2(n16577), .ZN(n15556) );
  OAI211_X1 U18909 ( .C1(n15558), .C2(n16589), .A(n15557), .B(n15556), .ZN(
        P2_U3017) );
  NOR2_X1 U18910 ( .A1(n19554), .A2(n16336), .ZN(n15564) );
  INV_X1 U18911 ( .A(n15559), .ZN(n15560) );
  NAND3_X1 U18912 ( .A1(n15572), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15560), .ZN(n15561) );
  OAI211_X1 U18913 ( .C1(n16328), .C2(n19540), .A(n15562), .B(n15561), .ZN(
        n15563) );
  AOI211_X1 U18914 ( .C1(n15565), .C2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15564), .B(n15563), .ZN(n15568) );
  NAND2_X1 U18915 ( .A1(n15566), .A2(n16577), .ZN(n15567) );
  OAI211_X1 U18916 ( .C1(n15569), .C2(n16589), .A(n15568), .B(n15567), .ZN(
        P2_U3018) );
  NAND3_X1 U18917 ( .A1(n15571), .A2(n19551), .A3(n15570), .ZN(n15582) );
  NOR2_X1 U18918 ( .A1(n19554), .A2(n16338), .ZN(n15576) );
  NAND2_X1 U18919 ( .A1(n15572), .A2(n12246), .ZN(n15573) );
  OAI211_X1 U18920 ( .C1(n16339), .C2(n19540), .A(n15574), .B(n15573), .ZN(
        n15575) );
  AOI211_X1 U18921 ( .C1(n15577), .C2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15576), .B(n15575), .ZN(n15581) );
  NAND3_X1 U18922 ( .A1(n15579), .A2(n16577), .A3(n15578), .ZN(n15580) );
  NAND3_X1 U18923 ( .A1(n15582), .A2(n15581), .A3(n15580), .ZN(P2_U3019) );
  INV_X1 U18924 ( .A(n15583), .ZN(n15586) );
  NAND3_X1 U18925 ( .A1(n15584), .A2(n15588), .A3(n15587), .ZN(n15585) );
  OAI211_X1 U18926 ( .C1(n16349), .C2(n19540), .A(n15586), .B(n15585), .ZN(
        n15590) );
  NAND3_X1 U18927 ( .A1(n15604), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15587), .ZN(n15600) );
  AOI21_X1 U18928 ( .B1(n15605), .B2(n15600), .A(n15588), .ZN(n15589) );
  AOI211_X1 U18929 ( .C1(n19537), .C2(n16350), .A(n15590), .B(n15589), .ZN(
        n15593) );
  NAND2_X1 U18930 ( .A1(n15591), .A2(n19551), .ZN(n15592) );
  OAI211_X1 U18931 ( .C1(n15594), .C2(n19556), .A(n15593), .B(n15592), .ZN(
        P2_U3020) );
  XNOR2_X1 U18932 ( .A(n15413), .B(n15604), .ZN(n16419) );
  INV_X1 U18933 ( .A(n15595), .ZN(n15596) );
  NOR2_X1 U18934 ( .A1(n15597), .A2(n15596), .ZN(n15598) );
  XNOR2_X1 U18935 ( .A(n15599), .B(n15598), .ZN(n16421) );
  NAND2_X1 U18936 ( .A1(n19560), .A2(n16420), .ZN(n15601) );
  OAI211_X1 U18937 ( .C1(n19324), .C2(n20122), .A(n15601), .B(n15600), .ZN(
        n15602) );
  AOI21_X1 U18938 ( .B1(n19537), .B2(n16360), .A(n15602), .ZN(n15603) );
  OAI21_X1 U18939 ( .B1(n15605), .B2(n15604), .A(n15603), .ZN(n15606) );
  AOI21_X1 U18940 ( .B1(n16421), .B2(n19551), .A(n15606), .ZN(n15607) );
  OAI21_X1 U18941 ( .B1(n16419), .B2(n19556), .A(n15607), .ZN(P2_U3021) );
  NAND2_X1 U18942 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n19517), .ZN(n15608) );
  OAI221_X1 U18943 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15611), 
        .C1(n15610), .C2(n15609), .A(n15608), .ZN(n15614) );
  XNOR2_X1 U18944 ( .A(n15146), .B(n15612), .ZN(n16405) );
  OAI22_X1 U18945 ( .A1(n16405), .A2(n19554), .B1(n19540), .B2(n16386), .ZN(
        n15613) );
  AOI211_X1 U18946 ( .C1(n15615), .C2(n19551), .A(n15614), .B(n15613), .ZN(
        n15616) );
  OAI21_X1 U18947 ( .B1(n15617), .B2(n19556), .A(n15616), .ZN(P2_U3022) );
  NOR2_X1 U18948 ( .A1(n19554), .A2(n15618), .ZN(n15623) );
  AOI22_X1 U18949 ( .A1(n19517), .A2(P2_REIP_REG_22__SCAN_IN), .B1(n16515), 
        .B2(n15619), .ZN(n15620) );
  OAI21_X1 U18950 ( .B1(n19540), .B2(n15621), .A(n15620), .ZN(n15622) );
  AOI211_X1 U18951 ( .C1(n16509), .C2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15623), .B(n15622), .ZN(n15626) );
  NAND2_X1 U18952 ( .A1(n15624), .A2(n19551), .ZN(n15625) );
  OAI211_X1 U18953 ( .C1(n15627), .C2(n19556), .A(n15626), .B(n15625), .ZN(
        P2_U3024) );
  NAND2_X1 U18954 ( .A1(n15628), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15633) );
  NAND2_X1 U18955 ( .A1(n19549), .A2(n15633), .ZN(n15629) );
  NAND2_X1 U18956 ( .A1(n15748), .A2(n15629), .ZN(n15722) );
  INV_X1 U18957 ( .A(n15634), .ZN(n15630) );
  AND2_X1 U18958 ( .A1(n19549), .A2(n15630), .ZN(n15631) );
  AND2_X1 U18959 ( .A1(n19549), .A2(n15635), .ZN(n15632) );
  NOR2_X1 U18960 ( .A1(n16524), .A2(n15632), .ZN(n15663) );
  NAND2_X1 U18961 ( .A1(n16046), .A2(n15634), .ZN(n16522) );
  OR3_X1 U18962 ( .A1(n16522), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n15635), .ZN(n15650) );
  NAND2_X1 U18963 ( .A1(n15663), .A2(n15650), .ZN(n15643) );
  INV_X1 U18964 ( .A(n15635), .ZN(n15637) );
  NAND3_X1 U18965 ( .A1(n15637), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n15636), .ZN(n15641) );
  INV_X1 U18966 ( .A(n19214), .ZN(n16398) );
  AOI21_X1 U18967 ( .B1(n16398), .B2(n19560), .A(n15638), .ZN(n15640) );
  NAND2_X1 U18968 ( .A1(n19537), .A2(n19215), .ZN(n15639) );
  OAI211_X1 U18969 ( .C1(n16522), .C2(n15641), .A(n15640), .B(n15639), .ZN(
        n15642) );
  AOI21_X1 U18970 ( .B1(n15643), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15642), .ZN(n15646) );
  NAND2_X1 U18971 ( .A1(n15644), .A2(n19551), .ZN(n15645) );
  OAI211_X1 U18972 ( .C1(n15647), .C2(n19556), .A(n15646), .B(n15645), .ZN(
        P2_U3026) );
  NAND2_X1 U18973 ( .A1(P2_REIP_REG_19__SCAN_IN), .A2(n19517), .ZN(n15648) );
  OAI21_X1 U18974 ( .B1(n19236), .B2(n19540), .A(n15648), .ZN(n15649) );
  AOI21_X1 U18975 ( .B1(n19537), .B2(n19234), .A(n15649), .ZN(n15651) );
  OAI211_X1 U18976 ( .C1(n15663), .C2(n15652), .A(n15651), .B(n15650), .ZN(
        n15653) );
  AOI21_X1 U18977 ( .B1(n19551), .B2(n15654), .A(n15653), .ZN(n15655) );
  OAI21_X1 U18978 ( .B1(n15656), .B2(n19556), .A(n15655), .ZN(P2_U3027) );
  AOI22_X1 U18979 ( .A1(n19537), .A2(n15657), .B1(P2_REIP_REG_18__SCAN_IN), 
        .B2(n19517), .ZN(n15658) );
  OAI21_X1 U18980 ( .B1(n19540), .B2(n16402), .A(n15658), .ZN(n15661) );
  NOR3_X1 U18981 ( .A1(n16522), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15659), .ZN(n15660) );
  AOI211_X1 U18982 ( .C1(n15662), .C2(n19551), .A(n15661), .B(n15660), .ZN(
        n15666) );
  INV_X1 U18983 ( .A(n15663), .ZN(n15664) );
  NAND2_X1 U18984 ( .A1(n15664), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15665) );
  OAI211_X1 U18985 ( .C1(n15667), .C2(n19556), .A(n15666), .B(n15665), .ZN(
        P2_U3028) );
  INV_X1 U18986 ( .A(n16524), .ZN(n15669) );
  OAI211_X1 U18987 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n19533), .A(
        n15670), .B(n15669), .ZN(n15682) );
  AOI21_X1 U18988 ( .B1(n15671), .B2(n19549), .A(n15682), .ZN(n15680) );
  OAI22_X1 U18989 ( .A1(n15673), .A2(n19540), .B1(n15672), .B2(n19350), .ZN(
        n15676) );
  NOR2_X1 U18990 ( .A1(n15674), .A2(n16589), .ZN(n15675) );
  INV_X1 U18991 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16432) );
  OAI22_X1 U18992 ( .A1(n16435), .A2(n19556), .B1(n16432), .B2(n16522), .ZN(
        n15681) );
  NAND3_X1 U18993 ( .A1(n15681), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15679), .ZN(n15677) );
  OAI211_X1 U18994 ( .C1(n15680), .C2(n15679), .A(n15678), .B(n15677), .ZN(
        P2_U3029) );
  INV_X1 U18995 ( .A(n15681), .ZN(n15690) );
  NAND2_X1 U18996 ( .A1(n15682), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15689) );
  NOR2_X1 U18997 ( .A1(n19540), .A2(n15683), .ZN(n15686) );
  OAI22_X1 U18998 ( .A1(n19554), .A2(n19274), .B1(n15684), .B2(n19350), .ZN(
        n15685) );
  AOI211_X1 U18999 ( .C1(n15687), .C2(n19551), .A(n15686), .B(n15685), .ZN(
        n15688) );
  OAI211_X1 U19000 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15690), .A(
        n15689), .B(n15688), .ZN(P2_U3030) );
  INV_X1 U19001 ( .A(n15691), .ZN(n16433) );
  OAI21_X1 U19002 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16446), .A(
        n16433), .ZN(n16442) );
  OAI21_X1 U19003 ( .B1(n15693), .B2(n16531), .A(n15692), .ZN(n19424) );
  AND4_X1 U19004 ( .A1(n15696), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A4(n16046), .ZN(n15694) );
  AOI21_X1 U19005 ( .B1(n19517), .B2(P2_REIP_REG_14__SCAN_IN), .A(n15694), 
        .ZN(n15695) );
  OAI21_X1 U19006 ( .B1(n19554), .B2(n19424), .A(n15695), .ZN(n15698) );
  AOI21_X1 U19007 ( .B1(n16046), .B2(n16535), .A(n15722), .ZN(n16537) );
  NAND2_X1 U19008 ( .A1(n16046), .A2(n16536), .ZN(n16534) );
  AOI21_X1 U19009 ( .B1(n16537), .B2(n16534), .A(n15696), .ZN(n15697) );
  AOI211_X1 U19010 ( .C1(n19560), .C2(n19294), .A(n15698), .B(n15697), .ZN(
        n15707) );
  AOI21_X1 U19011 ( .B1(n15701), .B2(n15700), .A(n15699), .ZN(n15704) );
  INV_X1 U19012 ( .A(n15702), .ZN(n16429) );
  AND2_X1 U19013 ( .A1(n15704), .A2(n10165), .ZN(n16428) );
  NOR2_X1 U19014 ( .A1(n15704), .A2(n10165), .ZN(n15705) );
  NOR2_X1 U19015 ( .A1(n16428), .A2(n15705), .ZN(n16441) );
  OR2_X1 U19016 ( .A1(n16441), .A2(n16589), .ZN(n15706) );
  OAI211_X1 U19017 ( .C1(n16442), .C2(n19556), .A(n15707), .B(n15706), .ZN(
        P2_U3032) );
  INV_X1 U19018 ( .A(n15708), .ZN(n16469) );
  INV_X1 U19019 ( .A(n15709), .ZN(n16447) );
  OAI21_X1 U19020 ( .B1(n16469), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n16447), .ZN(n16459) );
  INV_X1 U19021 ( .A(n16046), .ZN(n15713) );
  INV_X1 U19022 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20104) );
  NOR2_X1 U19023 ( .A1(n20104), .A2(n19324), .ZN(n15711) );
  NOR2_X1 U19024 ( .A1(n19554), .A2(n19320), .ZN(n15710) );
  AOI211_X1 U19025 ( .C1(n19560), .C2(n19316), .A(n15711), .B(n15710), .ZN(
        n15712) );
  OAI21_X1 U19026 ( .B1(n15713), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15712), .ZN(n15721) );
  NAND2_X1 U19027 ( .A1(n15715), .A2(n15714), .ZN(n15719) );
  AND2_X1 U19028 ( .A1(n15717), .A2(n15716), .ZN(n15718) );
  XNOR2_X1 U19029 ( .A(n15719), .B(n15718), .ZN(n16458) );
  NOR2_X1 U19030 ( .A1(n16458), .A2(n16589), .ZN(n15720) );
  AOI211_X1 U19031 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n15722), .A(
        n15721), .B(n15720), .ZN(n15723) );
  OAI21_X1 U19032 ( .B1(n19556), .B2(n16459), .A(n15723), .ZN(P2_U3034) );
  XNOR2_X1 U19033 ( .A(n15724), .B(n15731), .ZN(n16475) );
  INV_X1 U19034 ( .A(n15725), .ZN(n15743) );
  OR2_X1 U19035 ( .A1(n9789), .A2(n15743), .ZN(n15729) );
  AND2_X1 U19036 ( .A1(n15727), .A2(n15726), .ZN(n15728) );
  XNOR2_X1 U19037 ( .A(n15729), .B(n15728), .ZN(n16474) );
  NOR2_X1 U19038 ( .A1(n15749), .A2(n15750), .ZN(n16552) );
  OAI21_X1 U19039 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15750), .A(
        n15748), .ZN(n16544) );
  NOR2_X1 U19040 ( .A1(n10777), .A2(n19324), .ZN(n15730) );
  AOI221_X1 U19041 ( .B1(n16552), .B2(n15731), .C1(n16544), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n15730), .ZN(n15739) );
  NAND2_X1 U19042 ( .A1(n15733), .A2(n15732), .ZN(n15734) );
  INV_X1 U19043 ( .A(n19407), .ZN(n15736) );
  OAI22_X1 U19044 ( .A1(n19554), .A2(n19333), .B1(n19540), .B2(n15736), .ZN(
        n15737) );
  INV_X1 U19045 ( .A(n15737), .ZN(n15738) );
  OAI211_X1 U19046 ( .C1(n16474), .C2(n16589), .A(n15739), .B(n15738), .ZN(
        n15740) );
  INV_X1 U19047 ( .A(n15740), .ZN(n15741) );
  OAI21_X1 U19048 ( .B1(n16475), .B2(n19556), .A(n15741), .ZN(P2_U3036) );
  OAI21_X1 U19049 ( .B1(n15742), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15724), .ZN(n16480) );
  NOR2_X1 U19050 ( .A1(n15744), .A2(n15743), .ZN(n15745) );
  XNOR2_X1 U19051 ( .A(n15746), .B(n15745), .ZN(n16482) );
  NAND2_X1 U19052 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19517), .ZN(n15747) );
  OAI221_X1 U19053 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15750), .C1(
        n15749), .C2(n15748), .A(n15747), .ZN(n15754) );
  OAI22_X1 U19054 ( .A1(n19554), .A2(n15752), .B1(n19540), .B2(n15751), .ZN(
        n15753) );
  AOI211_X1 U19055 ( .C1(n16482), .C2(n19551), .A(n15754), .B(n15753), .ZN(
        n15755) );
  OAI21_X1 U19056 ( .B1(n16480), .B2(n19556), .A(n15755), .ZN(P2_U3037) );
  NAND2_X1 U19057 ( .A1(n15757), .A2(n15756), .ZN(n15758) );
  XNOR2_X1 U19058 ( .A(n15759), .B(n15758), .ZN(n16489) );
  NAND2_X1 U19059 ( .A1(n16489), .A2(n19551), .ZN(n15770) );
  INV_X1 U19060 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20098) );
  NOR2_X1 U19061 ( .A1(n20098), .A2(n19324), .ZN(n15760) );
  AOI221_X1 U19062 ( .B1(n15761), .B2(n15763), .C1(n16565), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n15760), .ZN(n15769) );
  INV_X1 U19063 ( .A(n19353), .ZN(n16488) );
  AOI22_X1 U19064 ( .A1(n15762), .A2(n19537), .B1(n19560), .B2(n16488), .ZN(
        n15768) );
  XNOR2_X1 U19065 ( .A(n15764), .B(n15763), .ZN(n15765) );
  XNOR2_X1 U19066 ( .A(n15766), .B(n15765), .ZN(n16487) );
  NAND2_X1 U19067 ( .A1(n16487), .A2(n16577), .ZN(n15767) );
  NAND4_X1 U19068 ( .A1(n15770), .A2(n15769), .A3(n15768), .A4(n15767), .ZN(
        P2_U3039) );
  INV_X1 U19069 ( .A(n16634), .ZN(n15818) );
  INV_X1 U19070 ( .A(n15799), .ZN(n20148) );
  INV_X1 U19071 ( .A(n15795), .ZN(n15816) );
  INV_X1 U19072 ( .A(n12528), .ZN(n15772) );
  NAND2_X1 U19073 ( .A1(n15772), .A2(n15771), .ZN(n15782) );
  MUX2_X1 U19074 ( .A(n15782), .B(n15803), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15773) );
  AOI21_X1 U19075 ( .B1(n19513), .B2(n15816), .A(n15773), .ZN(n16596) );
  AOI22_X1 U19076 ( .A1(n19372), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n15774), .B2(n13243), .ZN(n15778) );
  INV_X1 U19077 ( .A(n15778), .ZN(n15775) );
  OAI222_X1 U19078 ( .A1(n15818), .A2(n13418), .B1(n20148), .B2(n16596), .C1(
        n15777), .C2(n15775), .ZN(n15776) );
  MUX2_X1 U19079 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n15776), .S(
        n15820), .Z(P2_U3601) );
  INV_X1 U19080 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n15777) );
  NOR2_X1 U19081 ( .A1(n15778), .A2(n15777), .ZN(n15797) );
  INV_X1 U19082 ( .A(n15797), .ZN(n15786) );
  OAI21_X1 U19083 ( .B1(n19299), .B2(n15780), .A(n15779), .ZN(n15798) );
  NAND2_X1 U19084 ( .A1(n19559), .A2(n15816), .ZN(n15785) );
  XNOR2_X1 U19085 ( .A(n10223), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15783) );
  AOI22_X1 U19086 ( .A1(n15803), .A2(n10223), .B1(n15783), .B2(n15782), .ZN(
        n15784) );
  AND2_X1 U19087 ( .A1(n15785), .A2(n15784), .ZN(n16597) );
  OAI222_X1 U19088 ( .A1(n20166), .A2(n15818), .B1(n15786), .B2(n15798), .C1(
        n20148), .C2(n16597), .ZN(n15787) );
  MUX2_X1 U19089 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15787), .S(
        n15820), .Z(P2_U3600) );
  NOR2_X1 U19090 ( .A1(n15788), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15810) );
  NOR2_X1 U19091 ( .A1(n15810), .A2(n10622), .ZN(n15793) );
  NAND2_X1 U19092 ( .A1(n10705), .A2(n15789), .ZN(n15805) );
  INV_X1 U19093 ( .A(n15803), .ZN(n15809) );
  NOR3_X1 U19094 ( .A1(n15809), .A2(n15790), .A3(n9694), .ZN(n15792) );
  NOR2_X1 U19095 ( .A1(n16607), .A2(n16613), .ZN(n15811) );
  NOR2_X1 U19096 ( .A1(n15811), .A2(n15793), .ZN(n15791) );
  AOI211_X1 U19097 ( .C1(n15793), .C2(n15805), .A(n15792), .B(n15791), .ZN(
        n15794) );
  OAI21_X1 U19098 ( .B1(n19541), .B2(n15795), .A(n15794), .ZN(n16601) );
  AOI222_X1 U19099 ( .A1(n16601), .A2(n15799), .B1(n15798), .B2(n15797), .C1(
        n16634), .C2(n15796), .ZN(n15802) );
  INV_X1 U19100 ( .A(n15820), .ZN(n15801) );
  NAND2_X1 U19101 ( .A1(n15801), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15800) );
  OAI21_X1 U19102 ( .B1(n15802), .B2(n15801), .A(n15800), .ZN(P2_U3599) );
  INV_X1 U19103 ( .A(n12269), .ZN(n15808) );
  AOI21_X1 U19104 ( .B1(n15803), .B2(n15808), .A(n15810), .ZN(n15807) );
  NAND2_X1 U19105 ( .A1(n15805), .A2(n15804), .ZN(n15806) );
  NAND2_X1 U19106 ( .A1(n15807), .A2(n15806), .ZN(n15813) );
  OAI22_X1 U19107 ( .A1(n15811), .A2(n15810), .B1(n15809), .B2(n15808), .ZN(
        n15812) );
  MUX2_X1 U19108 ( .A(n15813), .B(n15812), .S(n10283), .Z(n15814) );
  AOI211_X1 U19109 ( .C1(n15817), .C2(n15816), .A(n15815), .B(n15814), .ZN(
        n16595) );
  OAI22_X1 U19110 ( .A1(n15819), .A2(n15818), .B1(n16595), .B2(n20148), .ZN(
        n15821) );
  MUX2_X1 U19111 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15821), .S(
        n15820), .Z(P2_U3596) );
  INV_X1 U19112 ( .A(n19990), .ZN(n15822) );
  NAND2_X1 U19113 ( .A1(n15822), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n15824) );
  AOI22_X1 U19114 ( .A1(n20005), .A2(n20055), .B1(n20002), .B2(n19984), .ZN(
        n15823) );
  OAI211_X1 U19115 ( .C1(n15825), .C2(n19923), .A(n15824), .B(n15823), .ZN(
        n15826) );
  AOI21_X1 U19116 ( .B1(n20003), .B2(n19986), .A(n15826), .ZN(n15827) );
  INV_X1 U19117 ( .A(n15827), .ZN(P2_U3160) );
  AOI22_X1 U19118 ( .A1(n17431), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9685), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15829) );
  OAI21_X1 U19119 ( .B1(n12919), .B2(n17418), .A(n15829), .ZN(n15839) );
  AOI22_X1 U19120 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12952), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15837) );
  AOI22_X1 U19121 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17488), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15830) );
  OAI21_X1 U19122 ( .B1(n17485), .B2(n17413), .A(n15830), .ZN(n15835) );
  AOI22_X1 U19123 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15832) );
  AOI22_X1 U19124 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15831) );
  OAI211_X1 U19125 ( .C1(n12943), .C2(n15833), .A(n15832), .B(n15831), .ZN(
        n15834) );
  AOI211_X1 U19126 ( .C1(n17490), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n15835), .B(n15834), .ZN(n15836) );
  OAI211_X1 U19127 ( .C1(n12984), .C2(n18733), .A(n15837), .B(n15836), .ZN(
        n15838) );
  AOI211_X1 U19128 ( .C1(n15895), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n15839), .B(n15838), .ZN(n17245) );
  AOI22_X1 U19129 ( .A1(n17430), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15840) );
  OAI21_X1 U19130 ( .B1(n12959), .B2(n15841), .A(n15840), .ZN(n15850) );
  INV_X1 U19131 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18809) );
  AOI22_X1 U19132 ( .A1(n17467), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17288), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15848) );
  AOI22_X1 U19133 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15842) );
  OAI21_X1 U19134 ( .B1(n17485), .B2(n17452), .A(n15842), .ZN(n15846) );
  AOI22_X1 U19135 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15844) );
  AOI22_X1 U19136 ( .A1(n9685), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17448), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15843) );
  OAI211_X1 U19137 ( .C1(n12943), .C2(n17337), .A(n15844), .B(n15843), .ZN(
        n15845) );
  AOI211_X1 U19138 ( .C1(n17488), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n15846), .B(n15845), .ZN(n15847) );
  OAI211_X1 U19139 ( .C1(n17429), .C2(n18809), .A(n15848), .B(n15847), .ZN(
        n15849) );
  AOI211_X1 U19140 ( .C1(n15895), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n15850), .B(n15849), .ZN(n17255) );
  INV_X1 U19141 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17484) );
  AOI22_X1 U19142 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12952), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15851) );
  OAI21_X1 U19143 ( .B1(n12919), .B2(n17484), .A(n15851), .ZN(n15861) );
  INV_X1 U19144 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15859) );
  AOI22_X1 U19145 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17488), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15858) );
  OAI22_X1 U19146 ( .A1(n17429), .A2(n18802), .B1(n12984), .B2(n18722), .ZN(
        n15856) );
  AOI22_X1 U19147 ( .A1(n9685), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15854) );
  AOI22_X1 U19148 ( .A1(n17467), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15853) );
  AOI22_X1 U19149 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15852) );
  NAND3_X1 U19150 ( .A1(n15854), .A2(n15853), .A3(n15852), .ZN(n15855) );
  AOI211_X1 U19151 ( .C1(n17449), .C2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n15856), .B(n15855), .ZN(n15857) );
  OAI211_X1 U19152 ( .C1(n15864), .C2(n15859), .A(n15858), .B(n15857), .ZN(
        n15860) );
  AOI211_X1 U19153 ( .C1(n15895), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n15861), .B(n15860), .ZN(n17265) );
  INV_X1 U19154 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17382) );
  AOI22_X1 U19155 ( .A1(n17467), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15862) );
  OAI21_X1 U19156 ( .B1(n12919), .B2(n17382), .A(n15862), .ZN(n15873) );
  AOI22_X1 U19157 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15871) );
  INV_X1 U19158 ( .A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n15863) );
  OAI22_X1 U19159 ( .A1(n9682), .A2(n15863), .B1(n12943), .B2(n18825), .ZN(
        n15869) );
  AOI22_X1 U19160 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15867) );
  AOI22_X1 U19161 ( .A1(n9685), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9704), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15866) );
  AOI22_X1 U19162 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17488), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15865) );
  NAND3_X1 U19163 ( .A1(n15867), .A2(n15866), .A3(n15865), .ZN(n15868) );
  AOI211_X1 U19164 ( .C1(n17288), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n15869), .B(n15868), .ZN(n15870) );
  OAI211_X1 U19165 ( .C1(n17485), .C2(n18537), .A(n15871), .B(n15870), .ZN(
        n15872) );
  AOI211_X1 U19166 ( .C1(n9689), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n15873), .B(n15872), .ZN(n17266) );
  NOR2_X1 U19167 ( .A1(n17265), .A2(n17266), .ZN(n17264) );
  AOI22_X1 U19168 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17488), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15883) );
  AOI22_X1 U19169 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17430), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17448), .ZN(n15874) );
  OAI21_X1 U19170 ( .B1(n12951), .B2(n18501), .A(n15874), .ZN(n15881) );
  OAI22_X1 U19171 ( .A1(n17429), .A2(n18806), .B1(n17471), .B2(n17485), .ZN(
        n15875) );
  AOI21_X1 U19172 ( .B1(n9688), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n15875), .ZN(n15879) );
  AOI22_X1 U19173 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n15828), .B1(
        n17431), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15878) );
  AOI22_X1 U19174 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17482), .B1(
        n12970), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15877) );
  AOI22_X1 U19175 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17490), .B1(
        n17393), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15876) );
  NAND4_X1 U19176 ( .A1(n15879), .A2(n15878), .A3(n15877), .A4(n15876), .ZN(
        n15880) );
  AOI211_X1 U19177 ( .C1(n15895), .C2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n15881), .B(n15880), .ZN(n15882) );
  OAI211_X1 U19178 ( .C1(n17464), .C2(n12943), .A(n15883), .B(n15882), .ZN(
        n17260) );
  NAND2_X1 U19179 ( .A1(n17264), .A2(n17260), .ZN(n17259) );
  NOR2_X1 U19180 ( .A1(n17255), .A2(n17259), .ZN(n17254) );
  AOI22_X1 U19181 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15893) );
  AOI22_X1 U19182 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15892) );
  AOI22_X1 U19183 ( .A1(n17488), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15891) );
  OAI22_X1 U19184 ( .A1(n12951), .A2(n18512), .B1(n12984), .B2(n17315), .ZN(
        n15889) );
  AOI22_X1 U19185 ( .A1(n17467), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15887) );
  AOI22_X1 U19186 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15886) );
  AOI22_X1 U19187 ( .A1(n17490), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15885) );
  NAND2_X1 U19188 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n15884) );
  NAND4_X1 U19189 ( .A1(n15887), .A2(n15886), .A3(n15885), .A4(n15884), .ZN(
        n15888) );
  AOI211_X1 U19190 ( .C1(n17430), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n15889), .B(n15888), .ZN(n15890) );
  NAND4_X1 U19191 ( .A1(n15893), .A2(n15892), .A3(n15891), .A4(n15890), .ZN(
        n17250) );
  NAND2_X1 U19192 ( .A1(n17254), .A2(n17250), .ZN(n17249) );
  NOR2_X1 U19193 ( .A1(n17245), .A2(n17249), .ZN(n17244) );
  AOI22_X1 U19194 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15905) );
  INV_X1 U19195 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15916) );
  AOI22_X1 U19196 ( .A1(n17467), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9704), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15897) );
  AOI22_X1 U19197 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15896) );
  OAI211_X1 U19198 ( .C1(n17470), .C2(n15916), .A(n15897), .B(n15896), .ZN(
        n15903) );
  AOI22_X1 U19199 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15901) );
  AOI22_X1 U19200 ( .A1(n9685), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15900) );
  AOI22_X1 U19201 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15899) );
  NAND2_X1 U19202 ( .A1(n17490), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n15898) );
  NAND4_X1 U19203 ( .A1(n15901), .A2(n15900), .A3(n15899), .A4(n15898), .ZN(
        n15902) );
  AOI211_X1 U19204 ( .C1(n17393), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n15903), .B(n15902), .ZN(n15904) );
  OAI211_X1 U19205 ( .C1(n12984), .C2(n18736), .A(n15905), .B(n15904), .ZN(
        n15906) );
  NAND2_X1 U19206 ( .A1(n17244), .A2(n15906), .ZN(n17237) );
  OAI21_X1 U19207 ( .B1(n17244), .B2(n15906), .A(n17237), .ZN(n17552) );
  INV_X1 U19208 ( .A(n18957), .ZN(n15942) );
  NAND2_X1 U19209 ( .A1(n18533), .A2(n18514), .ZN(n15907) );
  INV_X1 U19210 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n17203) );
  INV_X1 U19211 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17202) );
  INV_X1 U19212 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16908) );
  INV_X1 U19213 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16928) );
  INV_X1 U19214 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16948) );
  INV_X1 U19215 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17341) );
  INV_X1 U19216 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n15910) );
  INV_X1 U19217 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17426) );
  NAND2_X1 U19218 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17521) );
  NOR2_X1 U19219 ( .A1(n17519), .A2(n17521), .ZN(n17512) );
  NAND3_X1 U19220 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17512), .ZN(n17421) );
  INV_X1 U19221 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17071) );
  INV_X1 U19222 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17442) );
  INV_X1 U19223 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17143) );
  NAND3_X1 U19224 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(P3_EBX_REG_6__SCAN_IN), .ZN(n17441) );
  NOR4_X1 U19225 ( .A1(n17071), .A2(n17442), .A3(n17143), .A4(n17441), .ZN(
        n15909) );
  NAND2_X1 U19226 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n15909), .ZN(n17422) );
  NOR3_X1 U19227 ( .A1(n17426), .A2(n17421), .A3(n17422), .ZN(n15923) );
  INV_X1 U19228 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17022) );
  INV_X1 U19229 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17408) );
  NOR3_X1 U19230 ( .A1(n17022), .A2(n17408), .A3(n17389), .ZN(n17368) );
  NAND3_X1 U19231 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n15923), .A3(n17368), 
        .ZN(n17340) );
  NAND2_X1 U19232 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17328), .ZN(n17326) );
  INV_X1 U19233 ( .A(n17326), .ZN(n17311) );
  NAND2_X1 U19234 ( .A1(n18533), .A2(n17285), .ZN(n17298) );
  NAND2_X1 U19235 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17270), .ZN(n17263) );
  NAND2_X1 U19236 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17269), .ZN(n17253) );
  NAND2_X1 U19237 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17258), .ZN(n17243) );
  NOR3_X1 U19238 ( .A1(n17203), .A2(n17202), .A3(n17243), .ZN(n17239) );
  NOR2_X1 U19239 ( .A1(n17530), .A2(n17239), .ZN(n17235) );
  NOR2_X1 U19240 ( .A1(n17202), .A2(n17243), .ZN(n17248) );
  AOI22_X1 U19241 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17235), .B1(n17248), 
        .B2(n17203), .ZN(n15911) );
  OAI21_X1 U19242 ( .B1(n17552), .B2(n17525), .A(n15911), .ZN(P3_U2675) );
  INV_X1 U19243 ( .A(n15923), .ZN(n15924) );
  NAND2_X1 U19244 ( .A1(n18533), .A2(n17533), .ZN(n17528) );
  INV_X1 U19245 ( .A(n17528), .ZN(n17529) );
  NAND2_X1 U19246 ( .A1(n17529), .A2(n17389), .ZN(n17407) );
  AOI22_X1 U19247 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15912) );
  OAI21_X1 U19248 ( .B1(n9756), .B2(n18736), .A(n15912), .ZN(n15922) );
  AOI22_X1 U19249 ( .A1(n9685), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15920) );
  AOI22_X1 U19250 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15913) );
  OAI21_X1 U19251 ( .B1(n17486), .B2(n18523), .A(n15913), .ZN(n15918) );
  AOI22_X1 U19252 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15915) );
  AOI22_X1 U19253 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17431), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15914) );
  OAI211_X1 U19254 ( .C1(n15864), .C2(n15916), .A(n15915), .B(n15914), .ZN(
        n15917) );
  AOI211_X1 U19255 ( .C1(n17488), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n15918), .B(n15917), .ZN(n15919) );
  OAI211_X1 U19256 ( .C1(n17485), .C2(n18933), .A(n15920), .B(n15919), .ZN(
        n15921) );
  AOI211_X1 U19257 ( .C1(n15828), .C2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n15922), .B(n15921), .ZN(n17627) );
  NAND2_X1 U19258 ( .A1(n17533), .A2(n15923), .ZN(n17385) );
  NAND2_X1 U19259 ( .A1(n17525), .A2(n17385), .ZN(n17406) );
  OAI222_X1 U19260 ( .A1(n15924), .A2(n17407), .B1(n17525), .B2(n17627), .C1(
        n17389), .C2(n17406), .ZN(P3_U2690) );
  NOR2_X1 U19261 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19125), .ZN(
        n18538) );
  NOR3_X1 U19262 ( .A1(n19134), .A2(n19174), .A3(n19183), .ZN(n15925) );
  NAND3_X1 U19263 ( .A1(n15945), .A2(n17485), .A3(n18963), .ZN(n18480) );
  INV_X1 U19264 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18481) );
  INV_X1 U19265 ( .A(n15925), .ZN(n19123) );
  NOR2_X1 U19266 ( .A1(n18481), .A2(n19123), .ZN(n15944) );
  AOI211_X1 U19267 ( .C1(n15925), .C2(n18480), .A(n18857), .B(n15944), .ZN(
        n15926) );
  NOR2_X1 U19268 ( .A1(n18538), .A2(n15926), .ZN(n15928) );
  INV_X1 U19269 ( .A(n15932), .ZN(n18855) );
  INV_X1 U19270 ( .A(n15926), .ZN(n18486) );
  INV_X1 U19271 ( .A(n18105), .ZN(n18048) );
  OAI22_X1 U19272 ( .A1(n19168), .A2(n18048), .B1(n18487), .B2(n19125), .ZN(
        n15931) );
  NAND3_X1 U19273 ( .A1(n18996), .A2(n18486), .A3(n15931), .ZN(n15927) );
  OAI221_X1 U19274 ( .B1(n18996), .B2(n15928), .C1(n18996), .C2(n18855), .A(
        n15927), .ZN(P3_U2864) );
  NAND2_X1 U19275 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18713) );
  NOR2_X1 U19276 ( .A1(n19168), .A2(n18048), .ZN(n15930) );
  INV_X1 U19277 ( .A(n15928), .ZN(n15929) );
  AOI221_X1 U19278 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18713), .C1(n15930), 
        .C2(n18713), .A(n15929), .ZN(n18485) );
  OAI221_X1 U19279 ( .B1(n15932), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n15932), .C2(n15931), .A(n18486), .ZN(n18483) );
  AOI22_X1 U19280 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18485), .B1(
        n18483), .B2(n19001), .ZN(P3_U2865) );
  INV_X1 U19281 ( .A(n18955), .ZN(n15951) );
  INV_X1 U19282 ( .A(n19165), .ZN(n19172) );
  NOR2_X1 U19283 ( .A1(n15951), .A2(n19172), .ZN(n15940) );
  INV_X1 U19284 ( .A(n15933), .ZN(n17729) );
  NAND2_X1 U19285 ( .A1(n18498), .A2(n17729), .ZN(n19014) );
  OAI21_X1 U19286 ( .B1(n15937), .B2(n15936), .A(n15935), .ZN(n15939) );
  NAND2_X1 U19287 ( .A1(n15939), .A2(n15938), .ZN(n15953) );
  AOI21_X1 U19288 ( .B1(n15940), .B2(n17688), .A(n15953), .ZN(n15941) );
  OAI211_X1 U19289 ( .C1(n15943), .C2(n15942), .A(n15941), .B(n16036), .ZN(
        n18987) );
  NOR2_X1 U19290 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19125), .ZN(n18492) );
  INV_X1 U19291 ( .A(n19152), .ZN(n19150) );
  AOI21_X1 U19292 ( .B1(n15945), .B2(n18963), .A(n9864), .ZN(n19011) );
  NAND3_X1 U19293 ( .A1(n19150), .A2(n19184), .A3(n19011), .ZN(n15946) );
  OAI21_X1 U19294 ( .B1(n19150), .B2(n18963), .A(n15946), .ZN(P3_U3284) );
  INV_X1 U19295 ( .A(n18958), .ZN(n15958) );
  OAI21_X1 U19296 ( .B1(n15948), .B2(n15947), .A(n18514), .ZN(n15955) );
  OAI21_X1 U19297 ( .B1(n18503), .B2(n19171), .A(n19038), .ZN(n15949) );
  OAI21_X1 U19298 ( .B1(n15950), .B2(n15949), .A(n19165), .ZN(n16813) );
  NOR3_X1 U19299 ( .A1(n15952), .A2(n15951), .A3(n16813), .ZN(n15954) );
  AOI211_X1 U19300 ( .C1(n18957), .C2(n15955), .A(n15954), .B(n15953), .ZN(
        n15957) );
  AOI221_X4 U19301 ( .B1(n15958), .B2(n15957), .C1(n15956), .C2(n15957), .A(
        n19020), .ZN(n18471) );
  NAND2_X1 U19302 ( .A1(n18953), .A2(n18471), .ZN(n18468) );
  INV_X1 U19303 ( .A(n16647), .ZN(n16658) );
  AND2_X1 U19304 ( .A1(n18155), .A2(n16658), .ZN(n16692) );
  NOR3_X1 U19305 ( .A1(n15962), .A2(n15963), .A3(n18460), .ZN(n18153) );
  NOR3_X1 U19306 ( .A1(n13040), .A2(n18427), .A3(n18432), .ZN(n18398) );
  NAND3_X1 U19307 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n18398), .ZN(n18382) );
  NOR2_X1 U19308 ( .A1(n18370), .A2(n18382), .ZN(n18311) );
  OAI21_X1 U19309 ( .B1(n19149), .B2(n13031), .A(n18443), .ZN(n18424) );
  NAND2_X1 U19310 ( .A1(n18311), .A2(n18424), .ZN(n18303) );
  NOR2_X1 U19311 ( .A1(n15959), .A2(n18303), .ZN(n18257) );
  INV_X1 U19312 ( .A(n18257), .ZN(n18214) );
  NOR2_X1 U19313 ( .A1(n18443), .A2(n13031), .ZN(n18254) );
  NAND2_X1 U19314 ( .A1(n18398), .A2(n18254), .ZN(n18384) );
  OR3_X1 U19315 ( .A1(n18400), .A2(n18399), .A3(n18384), .ZN(n18371) );
  NOR2_X1 U19316 ( .A1(n18370), .A2(n18371), .ZN(n18305) );
  NAND2_X1 U19317 ( .A1(n18256), .A2(n18305), .ZN(n18259) );
  INV_X1 U19318 ( .A(n18988), .ZN(n18306) );
  AOI21_X1 U19319 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18306), .A(
        n18972), .ZN(n18452) );
  OAI22_X1 U19320 ( .A1(n18983), .A2(n18214), .B1(n18259), .B2(n18452), .ZN(
        n18178) );
  INV_X1 U19321 ( .A(n18178), .ZN(n15960) );
  INV_X1 U19322 ( .A(n17872), .ZN(n18288) );
  INV_X1 U19323 ( .A(n16689), .ZN(n18959) );
  NOR2_X1 U19324 ( .A1(n18959), .A2(n16687), .ZN(n18217) );
  NAND2_X1 U19325 ( .A1(n18288), .A2(n18217), .ZN(n16695) );
  AOI21_X1 U19326 ( .B1(n15960), .B2(n16695), .A(n16647), .ZN(n15961) );
  AOI22_X1 U19327 ( .A1(n18476), .A2(n16692), .B1(n18153), .B2(n15961), .ZN(
        n16021) );
  INV_X1 U19328 ( .A(n18280), .ZN(n18385) );
  INV_X1 U19329 ( .A(n18359), .ZN(n18277) );
  INV_X1 U19330 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17821) );
  INV_X1 U19331 ( .A(n18972), .ZN(n18990) );
  NOR3_X1 U19332 ( .A1(n15962), .A2(n15963), .A3(n18259), .ZN(n15965) );
  AOI21_X1 U19333 ( .B1(n18179), .B2(n18257), .A(n18983), .ZN(n18181) );
  AOI211_X1 U19334 ( .C1(n18964), .C2(n15963), .A(n18181), .B(n18460), .ZN(
        n18161) );
  NOR2_X1 U19335 ( .A1(n19149), .A2(n18259), .ZN(n18279) );
  NAND2_X1 U19336 ( .A1(n16644), .A2(n18279), .ZN(n18156) );
  NAND2_X1 U19337 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18160) );
  NOR2_X1 U19338 ( .A1(n15963), .A2(n18160), .ZN(n16645) );
  NAND2_X1 U19339 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n16645), .ZN(
        n16696) );
  OAI21_X1 U19340 ( .B1(n18156), .B2(n16696), .A(n18306), .ZN(n15964) );
  OAI211_X1 U19341 ( .C1(n18990), .C2(n15965), .A(n18161), .B(n15964), .ZN(
        n16017) );
  AOI21_X1 U19342 ( .B1(n18277), .B2(n17821), .A(n16017), .ZN(n16691) );
  OAI21_X1 U19343 ( .B1(n18385), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16691), .ZN(n15968) );
  NAND2_X1 U19344 ( .A1(n16689), .A2(n18471), .ZN(n18458) );
  NOR2_X1 U19345 ( .A1(n16687), .A2(n18458), .ZN(n18322) );
  NAND2_X1 U19346 ( .A1(n18155), .A2(n15966), .ZN(n16662) );
  AOI22_X1 U19347 ( .A1(n18322), .A2(n16657), .B1(n18476), .B2(n16662), .ZN(
        n16018) );
  INV_X1 U19348 ( .A(n16018), .ZN(n15967) );
  AOI21_X1 U19349 ( .B1(n18375), .B2(n15968), .A(n15967), .ZN(n15973) );
  INV_X1 U19350 ( .A(n18375), .ZN(n18435) );
  NAND2_X1 U19351 ( .A1(n18057), .A2(n17803), .ZN(n16697) );
  INV_X1 U19352 ( .A(n16697), .ZN(n15969) );
  AOI21_X1 U19353 ( .B1(n16688), .B2(n15970), .A(n15969), .ZN(n15971) );
  XNOR2_X1 U19354 ( .A(n15971), .B(n16671), .ZN(n16669) );
  AOI22_X1 U19355 ( .A1(n18435), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n18391), 
        .B2(n16669), .ZN(n15972) );
  OAI221_X1 U19356 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16021), 
        .C1(n16671), .C2(n15973), .A(n15972), .ZN(P3_U2833) );
  INV_X1 U19357 ( .A(n15974), .ZN(n15975) );
  AOI22_X1 U19358 ( .A1(n11172), .A2(n15976), .B1(n15975), .B2(n10900), .ZN(
        n20891) );
  NAND2_X1 U19359 ( .A1(n15977), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n20896) );
  NAND3_X1 U19360 ( .A1(n20891), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(
        n20896), .ZN(n15981) );
  INV_X1 U19361 ( .A(n15978), .ZN(n15980) );
  OAI211_X1 U19362 ( .C1(n11726), .C2(n15981), .A(n15980), .B(n15979), .ZN(
        n15983) );
  NAND2_X1 U19363 ( .A1(n15981), .A2(n11726), .ZN(n15982) );
  NAND2_X1 U19364 ( .A1(n15983), .A2(n15982), .ZN(n15984) );
  AOI222_X1 U19365 ( .A1(n15985), .A2(n15984), .B1(n15985), .B2(n11729), .C1(
        n15984), .C2(n11729), .ZN(n15987) );
  AOI21_X1 U19366 ( .B1(n15987), .B2(n15986), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n15989) );
  NOR2_X1 U19367 ( .A1(n15987), .A2(n15986), .ZN(n15988) );
  OAI21_X1 U19368 ( .B1(n15989), .B2(n15988), .A(n11733), .ZN(n15998) );
  NOR2_X1 U19369 ( .A1(P1_MORE_REG_SCAN_IN), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(
        n15992) );
  OAI211_X1 U19370 ( .C1(n15993), .C2(n15992), .A(n15991), .B(n15990), .ZN(
        n15994) );
  NOR2_X1 U19371 ( .A1(n15995), .A2(n15994), .ZN(n15997) );
  NAND3_X1 U19372 ( .A1(n15998), .A2(n15997), .A3(n15996), .ZN(n16007) );
  NAND3_X1 U19373 ( .A1(n20906), .A2(n15999), .A3(n21095), .ZN(n16000) );
  OR2_X1 U19374 ( .A1(n16001), .A2(n16000), .ZN(n16004) );
  OAI21_X1 U19375 ( .B1(n20906), .B2(n16002), .A(n20804), .ZN(n16003) );
  INV_X1 U19376 ( .A(n16299), .ZN(n16005) );
  AOI221_X1 U19377 ( .B1(n20222), .B2(n13985), .C1(n16007), .C2(n13985), .A(
        n16005), .ZN(n16009) );
  NOR2_X1 U19378 ( .A1(n16009), .A2(n20222), .ZN(n20807) );
  OAI21_X1 U19379 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20906), .A(n20807), 
        .ZN(n16303) );
  AOI211_X1 U19380 ( .C1(n16008), .C2(n16007), .A(n16006), .B(n16303), .ZN(
        n16013) );
  AOI21_X1 U19381 ( .B1(n16010), .B2(n20911), .A(n16009), .ZN(n16011) );
  INV_X1 U19382 ( .A(n16011), .ZN(n16012) );
  AOI22_X1 U19383 ( .A1(n16013), .A2(n16300), .B1(n20222), .B2(n16012), .ZN(
        P1_U3161) );
  NAND2_X1 U19384 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16655), .ZN(
        n16646) );
  AOI21_X1 U19385 ( .B1(n16015), .B2(n16655), .A(n16014), .ZN(n16652) );
  OAI221_X1 U19386 ( .B1(n16017), .B2(n18280), .C1(n16017), .C2(n16016), .A(
        n18375), .ZN(n16675) );
  AOI21_X1 U19387 ( .B1(n16018), .B2(n16675), .A(n16655), .ZN(n16019) );
  AOI21_X1 U19388 ( .B1(n18391), .B2(n16652), .A(n16019), .ZN(n16020) );
  INV_X1 U19389 ( .A(n18375), .ZN(n18408) );
  NAND2_X1 U19390 ( .A1(n18408), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16648) );
  OAI211_X1 U19391 ( .C1(n16021), .C2(n16646), .A(n16020), .B(n16648), .ZN(
        P3_U2832) );
  INV_X1 U19392 ( .A(HOLD), .ZN(n20819) );
  NOR2_X1 U19393 ( .A1(n10997), .A2(n20819), .ZN(n20810) );
  AOI22_X1 U19394 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n16024) );
  NAND2_X1 U19395 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n16022), .ZN(n20808) );
  OAI211_X1 U19396 ( .C1(n20810), .C2(n16024), .A(n16023), .B(n20808), .ZN(
        P1_U3195) );
  AND2_X1 U19397 ( .A1(n20340), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  AOI221_X1 U19398 ( .B1(n16027), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), 
        .C1(n16026), .C2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n16025), .ZN(
        n16031) );
  AOI22_X1 U19399 ( .A1(n16029), .A2(n16289), .B1(n16286), .B2(n16028), .ZN(
        n16030) );
  OAI211_X1 U19400 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n16032), .A(
        n16031), .B(n16030), .ZN(P1_U3011) );
  NOR3_X1 U19401 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20201), .A3(n20202), 
        .ZN(n20061) );
  NOR4_X1 U19402 ( .A1(n16033), .A2(n16633), .A3(n16641), .A4(n20061), .ZN(
        P2_U3178) );
  INV_X1 U19403 ( .A(n16628), .ZN(n20186) );
  AOI221_X1 U19404 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16641), .C1(n20186), .C2(
        n16641), .A(n19995), .ZN(n20180) );
  INV_X1 U19405 ( .A(n20180), .ZN(n20181) );
  NOR2_X1 U19406 ( .A1(n16626), .A2(n20181), .ZN(P2_U3047) );
  NAND3_X1 U19407 ( .A1(n18493), .A2(n18498), .A3(n16034), .ZN(n16035) );
  INV_X1 U19408 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17759) );
  NOR2_X1 U19409 ( .A1(n16038), .A2(n17759), .ZN(n17681) );
  NAND2_X1 U19410 ( .A1(n18533), .A2(n17537), .ZN(n17673) );
  AOI22_X1 U19411 ( .A1(n17684), .A2(BUF2_REG_0__SCAN_IN), .B1(n17683), .B2(
        n18146), .ZN(n16039) );
  OAI221_X1 U19412 ( .B1(n17681), .B2(n17759), .C1(n17681), .C2(n17673), .A(
        n16039), .ZN(P3_U2735) );
  AOI22_X1 U19413 ( .A1(n16509), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n19537), .B2(n16040), .ZN(n16051) );
  INV_X1 U19414 ( .A(n16041), .ZN(n16043) );
  OAI22_X1 U19415 ( .A1(n16043), .A2(n19556), .B1(n16042), .B2(n19540), .ZN(
        n16044) );
  AOI21_X1 U19416 ( .B1(n16045), .B2(n19551), .A(n16044), .ZN(n16050) );
  NAND3_X1 U19417 ( .A1(n16047), .A2(n16046), .A3(n15470), .ZN(n16048) );
  NAND4_X1 U19418 ( .A1(n16050), .A2(n16051), .A3(n16049), .A4(n16048), .ZN(
        P2_U3025) );
  AOI22_X1 U19419 ( .A1(P1_EBX_REG_21__SCAN_IN), .A2(n20304), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(n16052), .ZN(n16056) );
  AOI22_X1 U19420 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n20306), .B1(
        n16054), .B2(n16053), .ZN(n16055) );
  OAI211_X1 U19421 ( .C1(n20274), .C2(n16057), .A(n16056), .B(n16055), .ZN(
        n16058) );
  AOI21_X1 U19422 ( .B1(n16059), .B2(n20268), .A(n16058), .ZN(n16060) );
  OAI21_X1 U19423 ( .B1(n16061), .B2(n20292), .A(n16060), .ZN(P1_U2819) );
  INV_X1 U19424 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20857) );
  OAI21_X1 U19425 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(P1_REIP_REG_18__SCAN_IN), 
        .A(n16062), .ZN(n16063) );
  OAI22_X1 U19426 ( .A1(n20857), .A2(n16080), .B1(n16064), .B2(n16063), .ZN(
        n16065) );
  AOI211_X1 U19427 ( .C1(n20306), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n20288), .B(n16065), .ZN(n16070) );
  INV_X1 U19428 ( .A(n16121), .ZN(n16068) );
  INV_X1 U19429 ( .A(n16125), .ZN(n16067) );
  AOI222_X1 U19430 ( .A1(n16068), .A2(n20268), .B1(n16067), .B2(n20307), .C1(
        n20303), .C2(n16066), .ZN(n16069) );
  OAI211_X1 U19431 ( .C1(n16071), .C2(n20289), .A(n16070), .B(n16069), .ZN(
        P1_U2821) );
  NOR2_X1 U19432 ( .A1(n20851), .A2(n20848), .ZN(n16073) );
  AOI21_X1 U19433 ( .B1(n16073), .B2(n16072), .A(P1_REIP_REG_17__SCAN_IN), 
        .ZN(n16081) );
  OAI22_X1 U19434 ( .A1(n16075), .A2(n20254), .B1(n16074), .B2(n20289), .ZN(
        n16076) );
  AOI211_X1 U19435 ( .C1(n20307), .C2(n16139), .A(n20288), .B(n16076), .ZN(
        n16079) );
  INV_X1 U19436 ( .A(n16221), .ZN(n16077) );
  AOI22_X1 U19437 ( .A1(n16140), .A2(n20268), .B1(n20303), .B2(n16077), .ZN(
        n16078) );
  OAI211_X1 U19438 ( .C1(n16081), .C2(n16080), .A(n16079), .B(n16078), .ZN(
        P1_U2823) );
  INV_X1 U19439 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20844) );
  NAND2_X1 U19440 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n16082), .ZN(n16109) );
  OAI21_X1 U19441 ( .B1(n16084), .B2(n16109), .A(n16083), .ZN(n16103) );
  NAND2_X1 U19442 ( .A1(n16085), .A2(n20844), .ZN(n16090) );
  OAI22_X1 U19443 ( .A1(n16086), .A2(n20289), .B1(n20274), .B2(n16240), .ZN(
        n16087) );
  NOR2_X1 U19444 ( .A1(n16087), .A2(n20288), .ZN(n16089) );
  NAND2_X1 U19445 ( .A1(n20306), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16088) );
  OAI211_X1 U19446 ( .C1(n20259), .C2(n16090), .A(n16089), .B(n16088), .ZN(
        n16091) );
  INV_X1 U19447 ( .A(n16091), .ZN(n16092) );
  OAI21_X1 U19448 ( .B1(n16094), .B2(n16093), .A(n16092), .ZN(n16095) );
  AOI21_X1 U19449 ( .B1(n16096), .B2(n20307), .A(n16095), .ZN(n16097) );
  OAI21_X1 U19450 ( .B1(n20844), .B2(n16103), .A(n16097), .ZN(P1_U2827) );
  AND2_X1 U19451 ( .A1(n20309), .A2(n16098), .ZN(n16111) );
  AOI21_X1 U19452 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n16111), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n16104) );
  OAI22_X1 U19453 ( .A1(n16099), .A2(n20254), .B1(n16116), .B2(n20289), .ZN(
        n16100) );
  AOI211_X1 U19454 ( .C1(n16114), .C2(n20303), .A(n20288), .B(n16100), .ZN(
        n16102) );
  AOI22_X1 U19455 ( .A1(n16154), .A2(n20307), .B1(n20268), .B2(n16153), .ZN(
        n16101) );
  OAI211_X1 U19456 ( .C1(n16104), .C2(n16103), .A(n16102), .B(n16101), .ZN(
        P1_U2828) );
  XOR2_X1 U19457 ( .A(n16106), .B(n16105), .Z(n16248) );
  AOI22_X1 U19458 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(n20304), .B1(n20303), 
        .B2(n16248), .ZN(n16107) );
  OAI211_X1 U19459 ( .C1(n20254), .C2(n11341), .A(n16107), .B(n20276), .ZN(
        n16108) );
  AOI21_X1 U19460 ( .B1(n20268), .B2(n16163), .A(n16108), .ZN(n16113) );
  OAI22_X1 U19461 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n16111), .B1(n16110), 
        .B2(n16109), .ZN(n16112) );
  OAI211_X1 U19462 ( .C1(n20292), .C2(n16166), .A(n16113), .B(n16112), .ZN(
        P1_U2829) );
  AOI22_X1 U19463 ( .A1(n16153), .A2(n11783), .B1(n20320), .B2(n16114), .ZN(
        n16115) );
  OAI21_X1 U19464 ( .B1(n20324), .B2(n16116), .A(n16115), .ZN(P1_U2860) );
  AOI22_X1 U19465 ( .A1(n16163), .A2(n11783), .B1(n20320), .B2(n16248), .ZN(
        n16117) );
  OAI21_X1 U19466 ( .B1(n20324), .B2(n16118), .A(n16117), .ZN(P1_U2861) );
  AOI22_X1 U19467 ( .A1(n16173), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n16285), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16124) );
  OAI22_X1 U19468 ( .A1(n16121), .A2(n16120), .B1(n16119), .B2(n20226), .ZN(
        n16122) );
  INV_X1 U19469 ( .A(n16122), .ZN(n16123) );
  OAI211_X1 U19470 ( .C1(n16180), .C2(n16125), .A(n16124), .B(n16123), .ZN(
        P1_U2980) );
  NAND2_X1 U19471 ( .A1(n16135), .A2(n16126), .ZN(n16136) );
  INV_X1 U19472 ( .A(n16127), .ZN(n16128) );
  AOI211_X1 U19473 ( .C1(n16131), .C2(n16130), .A(n16129), .B(n16128), .ZN(
        n16133) );
  NOR2_X1 U19474 ( .A1(n16133), .A2(n16132), .ZN(n16134) );
  MUX2_X1 U19475 ( .A(n16136), .B(n16135), .S(n16134), .Z(n16138) );
  XNOR2_X1 U19476 ( .A(n16138), .B(n16137), .ZN(n16223) );
  AOI22_X1 U19477 ( .A1(n16173), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n16285), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16142) );
  AOI22_X1 U19478 ( .A1(n16140), .A2(n14887), .B1(n16139), .B2(n16181), .ZN(
        n16141) );
  OAI211_X1 U19479 ( .C1(n16223), .C2(n20226), .A(n16142), .B(n16141), .ZN(
        P1_U2982) );
  AOI22_X1 U19480 ( .A1(n16173), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n16285), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16146) );
  AOI22_X1 U19481 ( .A1(n16144), .A2(n14887), .B1(n16181), .B2(n16143), .ZN(
        n16145) );
  OAI211_X1 U19482 ( .C1(n20226), .C2(n16147), .A(n16146), .B(n16145), .ZN(
        P1_U2983) );
  AOI22_X1 U19483 ( .A1(n16173), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n16285), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16151) );
  AOI22_X1 U19484 ( .A1(n16149), .A2(n14887), .B1(n16181), .B2(n16148), .ZN(
        n16150) );
  OAI211_X1 U19485 ( .C1(n16152), .C2(n20226), .A(n16151), .B(n16150), .ZN(
        P1_U2984) );
  AOI22_X1 U19486 ( .A1(n16173), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n16285), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16156) );
  AOI22_X1 U19487 ( .A1(n16181), .A2(n16154), .B1(n14887), .B2(n16153), .ZN(
        n16155) );
  OAI211_X1 U19488 ( .C1(n16157), .C2(n20226), .A(n16156), .B(n16155), .ZN(
        P1_U2987) );
  AOI22_X1 U19489 ( .A1(n16173), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16285), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16165) );
  NOR2_X1 U19490 ( .A1(n14927), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16160) );
  INV_X1 U19491 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16260) );
  NOR2_X1 U19492 ( .A1(n14903), .A2(n16260), .ZN(n16159) );
  MUX2_X1 U19493 ( .A(n16160), .B(n16159), .S(n16158), .Z(n16162) );
  XNOR2_X1 U19494 ( .A(n16162), .B(n16161), .ZN(n16250) );
  AOI22_X1 U19495 ( .A1(n16183), .A2(n16250), .B1(n14887), .B2(n16163), .ZN(
        n16164) );
  OAI211_X1 U19496 ( .C1(n16180), .C2(n16166), .A(n16165), .B(n16164), .ZN(
        P1_U2988) );
  AOI22_X1 U19497 ( .A1(n16173), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16285), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16172) );
  XNOR2_X1 U19498 ( .A(n16167), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16168) );
  XNOR2_X1 U19499 ( .A(n16169), .B(n16168), .ZN(n16278) );
  INV_X1 U19500 ( .A(n16170), .ZN(n20261) );
  AOI22_X1 U19501 ( .A1(n16278), .A2(n16183), .B1(n14887), .B2(n20261), .ZN(
        n16171) );
  OAI211_X1 U19502 ( .C1(n16180), .C2(n20264), .A(n16172), .B(n16171), .ZN(
        P1_U2992) );
  AOI22_X1 U19503 ( .A1(n16173), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n16285), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16179) );
  NAND2_X1 U19504 ( .A1(n16175), .A2(n16174), .ZN(n16176) );
  XNOR2_X1 U19505 ( .A(n16177), .B(n16176), .ZN(n16290) );
  AOI22_X1 U19506 ( .A1(n16290), .A2(n16183), .B1(n14887), .B2(n20321), .ZN(
        n16178) );
  OAI211_X1 U19507 ( .C1(n16180), .C2(n20272), .A(n16179), .B(n16178), .ZN(
        P1_U2993) );
  INV_X1 U19508 ( .A(n20282), .ZN(n16182) );
  AOI222_X1 U19509 ( .A1(n16184), .A2(n16183), .B1(n14887), .B2(n20280), .C1(
        n16182), .C2(n16181), .ZN(n16186) );
  OAI211_X1 U19510 ( .C1(n16188), .C2(n16187), .A(n16186), .B(n16185), .ZN(
        P1_U2994) );
  AOI22_X1 U19511 ( .A1(n16285), .A2(P1_REIP_REG_23__SCAN_IN), .B1(n16190), 
        .B2(n16189), .ZN(n16196) );
  INV_X1 U19512 ( .A(n16191), .ZN(n16194) );
  INV_X1 U19513 ( .A(n16192), .ZN(n16193) );
  AOI22_X1 U19514 ( .A1(n16194), .A2(n16289), .B1(n16286), .B2(n16193), .ZN(
        n16195) );
  OAI211_X1 U19515 ( .C1(n16198), .C2(n16197), .A(n16196), .B(n16195), .ZN(
        P1_U3008) );
  AOI22_X1 U19516 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n16199), .B1(
        n16285), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n16208) );
  INV_X1 U19517 ( .A(n16200), .ZN(n16203) );
  INV_X1 U19518 ( .A(n16201), .ZN(n16202) );
  AOI22_X1 U19519 ( .A1(n16203), .A2(n16289), .B1(n16286), .B2(n16202), .ZN(
        n16207) );
  OAI211_X1 U19520 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16205), .B(n16204), .ZN(
        n16206) );
  NAND3_X1 U19521 ( .A1(n16208), .A2(n16207), .A3(n16206), .ZN(P1_U3009) );
  AOI21_X1 U19522 ( .B1(n16209), .B2(n16211), .A(n16230), .ZN(n16227) );
  NOR3_X1 U19523 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16211), .A3(
        n16210), .ZN(n16212) );
  AOI21_X1 U19524 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n16285), .A(n16212), 
        .ZN(n16217) );
  INV_X1 U19525 ( .A(n16213), .ZN(n16215) );
  AOI22_X1 U19526 ( .A1(n16215), .A2(n16289), .B1(n16286), .B2(n16214), .ZN(
        n16216) );
  OAI211_X1 U19527 ( .C1(n16227), .C2(n16218), .A(n16217), .B(n16216), .ZN(
        P1_U3013) );
  AOI21_X1 U19528 ( .B1(n16220), .B2(n16219), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16226) );
  OAI22_X1 U19529 ( .A1(n16223), .A2(n16222), .B1(n16239), .B2(n16221), .ZN(
        n16224) );
  AOI21_X1 U19530 ( .B1(n16285), .B2(P1_REIP_REG_17__SCAN_IN), .A(n16224), 
        .ZN(n16225) );
  OAI21_X1 U19531 ( .B1(n16227), .B2(n16226), .A(n16225), .ZN(P1_U3014) );
  AOI21_X1 U19532 ( .B1(n16229), .B2(n16286), .A(n16228), .ZN(n16237) );
  AOI22_X1 U19533 ( .A1(n16231), .A2(n16289), .B1(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16230), .ZN(n16236) );
  NAND3_X1 U19534 ( .A1(n16234), .A2(n16233), .A3(n16232), .ZN(n16235) );
  NAND3_X1 U19535 ( .A1(n16237), .A2(n16236), .A3(n16235), .ZN(P1_U3017) );
  OAI22_X1 U19536 ( .A1(n16240), .A2(n16239), .B1(n20844), .B2(n16238), .ZN(
        n16241) );
  AOI21_X1 U19537 ( .B1(n16242), .B2(n16289), .A(n16241), .ZN(n16243) );
  OAI221_X1 U19538 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16246), 
        .C1(n16245), .C2(n16244), .A(n16243), .ZN(P1_U3018) );
  INV_X1 U19539 ( .A(n16247), .ZN(n16253) );
  AOI22_X1 U19540 ( .A1(n16248), .A2(n16286), .B1(n16285), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16252) );
  AOI22_X1 U19541 ( .A1(n16250), .A2(n16289), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16249), .ZN(n16251) );
  OAI211_X1 U19542 ( .C1(n16287), .C2(n16253), .A(n16252), .B(n16251), .ZN(
        P1_U3020) );
  AOI21_X1 U19543 ( .B1(n16255), .B2(n16286), .A(n16254), .ZN(n16263) );
  AOI22_X1 U19544 ( .A1(n16257), .A2(n16289), .B1(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16256), .ZN(n16262) );
  OAI221_X1 U19545 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n16260), .C2(n16259), .A(
        n16258), .ZN(n16261) );
  NAND3_X1 U19546 ( .A1(n16263), .A2(n16262), .A3(n16261), .ZN(P1_U3021) );
  AOI21_X1 U19547 ( .B1(n16265), .B2(n16286), .A(n16264), .ZN(n16275) );
  INV_X1 U19548 ( .A(n16266), .ZN(n16269) );
  AOI21_X1 U19549 ( .B1(n16269), .B2(n16268), .A(n16267), .ZN(n16294) );
  OAI21_X1 U19550 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16270), .A(
        n16294), .ZN(n16277) );
  AOI22_X1 U19551 ( .A1(n16271), .A2(n16289), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16277), .ZN(n16274) );
  NOR2_X1 U19552 ( .A1(n16293), .A2(n16287), .ZN(n16276) );
  OAI211_X1 U19553 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16276), .B(n16272), .ZN(n16273) );
  NAND3_X1 U19554 ( .A1(n16275), .A2(n16274), .A3(n16273), .ZN(P1_U3023) );
  INV_X1 U19555 ( .A(n16276), .ZN(n16281) );
  AOI22_X1 U19556 ( .A1(n20251), .A2(n16286), .B1(n16285), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16280) );
  AOI22_X1 U19557 ( .A1(n16278), .A2(n16289), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16277), .ZN(n16279) );
  OAI211_X1 U19558 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16281), .A(
        n16280), .B(n16279), .ZN(P1_U3024) );
  INV_X1 U19559 ( .A(n16282), .ZN(n16284) );
  AOI21_X1 U19560 ( .B1(n9830), .B2(n16284), .A(n16283), .ZN(n20319) );
  AOI22_X1 U19561 ( .A1(n20319), .A2(n16286), .B1(n16285), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16292) );
  INV_X1 U19562 ( .A(n16287), .ZN(n16288) );
  AOI22_X1 U19563 ( .A1(n16290), .A2(n16289), .B1(n16293), .B2(n16288), .ZN(
        n16291) );
  OAI211_X1 U19564 ( .C1(n16294), .C2(n16293), .A(n16292), .B(n16291), .ZN(
        P1_U3025) );
  OR4_X1 U19565 ( .A1(n20284), .A2(n20894), .A3(n20897), .A4(n13506), .ZN(
        n16295) );
  OAI21_X1 U19566 ( .B1(n20892), .B2(n16296), .A(n16295), .ZN(P1_U3468) );
  NAND4_X1 U19567 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20806), .A4(n20906), .ZN(n16297) );
  AND2_X1 U19568 ( .A1(n16298), .A2(n16297), .ZN(n20805) );
  AOI21_X1 U19569 ( .B1(n20805), .B2(n16304), .A(n16299), .ZN(n16302) );
  INV_X1 U19570 ( .A(n16300), .ZN(n16301) );
  AOI211_X1 U19571 ( .C1(n13985), .C2(n16303), .A(n16302), .B(n16301), .ZN(
        P1_U3162) );
  OAI22_X1 U19572 ( .A1(n20807), .A2(n20700), .B1(n20222), .B2(n16304), .ZN(
        P1_U3466) );
  INV_X1 U19573 ( .A(n16305), .ZN(n16307) );
  INV_X1 U19574 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16306) );
  OAI222_X1 U19575 ( .A1(n19387), .A2(n20135), .B1(n19362), .B2(n16307), .C1(
        n19382), .C2(n16306), .ZN(n16308) );
  AOI21_X1 U19576 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19360), .A(
        n16308), .ZN(n16311) );
  INV_X1 U19577 ( .A(n16309), .ZN(n19416) );
  AOI22_X1 U19578 ( .A1(n16379), .A2(n19389), .B1(n19305), .B2(n19416), .ZN(
        n16310) );
  OAI211_X1 U19579 ( .C1(n19397), .C2(n16312), .A(n16311), .B(n16310), .ZN(
        P2_U2824) );
  AOI22_X1 U19580 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n19361), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19366), .ZN(n16323) );
  AOI22_X1 U19581 ( .A1(n16313), .A2(n19385), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19360), .ZN(n16322) );
  OAI22_X1 U19582 ( .A1(n16315), .A2(n19354), .B1(n16314), .B2(n19381), .ZN(
        n16316) );
  INV_X1 U19583 ( .A(n16316), .ZN(n16321) );
  OAI211_X1 U19584 ( .C1(n16319), .C2(n16318), .A(n19342), .B(n16317), .ZN(
        n16320) );
  NAND4_X1 U19585 ( .A1(n16323), .A2(n16322), .A3(n16321), .A4(n16320), .ZN(
        P2_U2826) );
  INV_X1 U19586 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n16325) );
  INV_X1 U19587 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16324) );
  OAI22_X1 U19588 ( .A1(n19382), .A2(n16325), .B1(n16324), .B2(n19391), .ZN(
        n16326) );
  AOI21_X1 U19589 ( .B1(n19366), .B2(P2_REIP_REG_28__SCAN_IN), .A(n16326), 
        .ZN(n16327) );
  OAI21_X1 U19590 ( .B1(n16328), .B2(n19354), .A(n16327), .ZN(n16329) );
  AOI21_X1 U19591 ( .B1(n16330), .B2(n19385), .A(n16329), .ZN(n16335) );
  OAI211_X1 U19592 ( .C1(n16333), .C2(n16332), .A(n19342), .B(n16331), .ZN(
        n16334) );
  OAI211_X1 U19593 ( .C1(n19381), .C2(n16336), .A(n16335), .B(n16334), .ZN(
        P2_U2827) );
  AOI22_X1 U19594 ( .A1(P2_EBX_REG_27__SCAN_IN), .A2(n19361), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19366), .ZN(n16347) );
  AOI22_X1 U19595 ( .A1(n16337), .A2(n19385), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n19360), .ZN(n16346) );
  OAI22_X1 U19596 ( .A1(n16339), .A2(n19354), .B1(n16338), .B2(n19381), .ZN(
        n16340) );
  INV_X1 U19597 ( .A(n16340), .ZN(n16345) );
  OAI211_X1 U19598 ( .C1(n16343), .C2(n16342), .A(n19342), .B(n16341), .ZN(
        n16344) );
  NAND4_X1 U19599 ( .A1(n16347), .A2(n16346), .A3(n16345), .A4(n16344), .ZN(
        P2_U2828) );
  AOI22_X1 U19600 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n19361), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19366), .ZN(n16358) );
  AOI22_X1 U19601 ( .A1(n16348), .A2(n19385), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19360), .ZN(n16357) );
  INV_X1 U19602 ( .A(n16349), .ZN(n16351) );
  AOI22_X1 U19603 ( .A1(n16351), .A2(n19389), .B1(n16350), .B2(n19305), .ZN(
        n16356) );
  OAI211_X1 U19604 ( .C1(n16354), .C2(n16353), .A(n19342), .B(n16352), .ZN(
        n16355) );
  NAND4_X1 U19605 ( .A1(n16358), .A2(n16357), .A3(n16356), .A4(n16355), .ZN(
        P2_U2829) );
  AOI22_X1 U19606 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n19361), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19366), .ZN(n16367) );
  AOI22_X1 U19607 ( .A1(n16359), .A2(n19385), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19360), .ZN(n16366) );
  AOI22_X1 U19608 ( .A1(n16420), .A2(n19389), .B1(n16360), .B2(n19305), .ZN(
        n16365) );
  OAI211_X1 U19609 ( .C1(n16363), .C2(n16362), .A(n19342), .B(n16361), .ZN(
        n16364) );
  NAND4_X1 U19610 ( .A1(n16367), .A2(n16366), .A3(n16365), .A4(n16364), .ZN(
        P2_U2830) );
  OAI22_X1 U19611 ( .A1(n16386), .A2(n19354), .B1(n16405), .B2(n19381), .ZN(
        n16368) );
  INV_X1 U19612 ( .A(n16368), .ZN(n16378) );
  OAI211_X1 U19613 ( .C1(n16371), .C2(n16370), .A(n19342), .B(n16369), .ZN(
        n16376) );
  AOI22_X1 U19614 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19360), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19366), .ZN(n16375) );
  NAND2_X1 U19615 ( .A1(n19361), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n16374) );
  OR2_X1 U19616 ( .A1(n16372), .A2(n19362), .ZN(n16373) );
  AND4_X1 U19617 ( .A1(n16376), .A2(n16375), .A3(n16374), .A4(n16373), .ZN(
        n16377) );
  NAND2_X1 U19618 ( .A1(n16378), .A2(n16377), .ZN(P2_U2831) );
  OAI22_X1 U19619 ( .A1(n16392), .A2(n16379), .B1(P2_EBX_REG_31__SCAN_IN), 
        .B2(n19406), .ZN(n16380) );
  INV_X1 U19620 ( .A(n16380), .ZN(P2_U2856) );
  AOI21_X1 U19621 ( .B1(n16383), .B2(n16382), .A(n16381), .ZN(n16385) );
  XNOR2_X1 U19622 ( .A(n16385), .B(n16384), .ZN(n16407) );
  INV_X1 U19623 ( .A(n16386), .ZN(n16387) );
  AOI22_X1 U19624 ( .A1(n16407), .A2(n19411), .B1(n19415), .B2(n16387), .ZN(
        n16388) );
  OAI21_X1 U19625 ( .B1(n19415), .B2(n10879), .A(n16388), .ZN(P2_U2863) );
  AOI21_X1 U19626 ( .B1(n16389), .B2(n16391), .A(n16390), .ZN(n16414) );
  AOI22_X1 U19627 ( .A1(n16414), .A2(n19411), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n16392), .ZN(n16393) );
  OAI21_X1 U19628 ( .B1(n16392), .B2(n16510), .A(n16393), .ZN(P2_U2864) );
  AOI22_X1 U19629 ( .A1(n16395), .A2(n19411), .B1(n19406), .B2(n16394), .ZN(
        n16396) );
  OAI21_X1 U19630 ( .B1(n19406), .B2(n16397), .A(n16396), .ZN(P2_U2865) );
  AOI22_X1 U19631 ( .A1(n16399), .A2(n19411), .B1(n19415), .B2(n16398), .ZN(
        n16400) );
  OAI21_X1 U19632 ( .B1(n19415), .B2(n16401), .A(n16400), .ZN(P2_U2867) );
  INV_X1 U19633 ( .A(n16402), .ZN(n19247) );
  AOI22_X1 U19634 ( .A1(n16403), .A2(n19411), .B1(n19406), .B2(n19247), .ZN(
        n16404) );
  OAI21_X1 U19635 ( .B1(n19415), .B2(n19241), .A(n16404), .ZN(P2_U2869) );
  AOI22_X1 U19636 ( .A1(n16412), .A2(n19433), .B1(n19432), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n16410) );
  AOI22_X1 U19637 ( .A1(n19418), .A2(BUF2_REG_24__SCAN_IN), .B1(n19419), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n16409) );
  INV_X1 U19638 ( .A(n16405), .ZN(n16406) );
  AOI22_X1 U19639 ( .A1(n16407), .A2(n16413), .B1(n19417), .B2(n16406), .ZN(
        n16408) );
  NAND3_X1 U19640 ( .A1(n16410), .A2(n16409), .A3(n16408), .ZN(P2_U2895) );
  AOI22_X1 U19641 ( .A1(n16412), .A2(n16411), .B1(n19432), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16417) );
  AOI22_X1 U19642 ( .A1(n19418), .A2(BUF2_REG_23__SCAN_IN), .B1(n19419), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n16416) );
  AOI22_X1 U19643 ( .A1(n16414), .A2(n16413), .B1(n19417), .B2(n16508), .ZN(
        n16415) );
  NAND3_X1 U19644 ( .A1(n16417), .A2(n16416), .A3(n16415), .ZN(P2_U2896) );
  AOI22_X1 U19645 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19517), .B1(n16494), 
        .B2(n16418), .ZN(n16424) );
  INV_X1 U19646 ( .A(n16419), .ZN(n16422) );
  AOI222_X1 U19647 ( .A1(n16422), .A2(n19507), .B1(n12279), .B2(n16421), .C1(
        n19512), .C2(n16420), .ZN(n16423) );
  OAI211_X1 U19648 ( .C1(n16425), .C2(n16506), .A(n16424), .B(n16423), .ZN(
        P2_U2989) );
  AOI22_X1 U19649 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19517), .B1(n16494), 
        .B2(n19277), .ZN(n16440) );
  NOR2_X1 U19650 ( .A1(n16427), .A2(n16426), .ZN(n16431) );
  NOR2_X1 U19651 ( .A1(n16429), .A2(n16428), .ZN(n16430) );
  XNOR2_X1 U19652 ( .A(n16431), .B(n16430), .ZN(n16530) );
  INV_X1 U19653 ( .A(n16530), .ZN(n16438) );
  NAND2_X1 U19654 ( .A1(n16433), .A2(n16432), .ZN(n16434) );
  NAND2_X1 U19655 ( .A1(n16435), .A2(n16434), .ZN(n16525) );
  OAI22_X1 U19656 ( .A1(n16525), .A2(n19495), .B1(n16436), .B2(n16526), .ZN(
        n16437) );
  AOI21_X1 U19657 ( .B1(n16438), .B2(n12279), .A(n16437), .ZN(n16439) );
  OAI211_X1 U19658 ( .C1(n19279), .C2(n16506), .A(n16440), .B(n16439), .ZN(
        P2_U2999) );
  AOI22_X1 U19659 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19503), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19517), .ZN(n16445) );
  OAI22_X1 U19660 ( .A1(n16442), .A2(n19495), .B1(n16441), .B2(n19510), .ZN(
        n16443) );
  AOI21_X1 U19661 ( .B1(n19512), .B2(n19294), .A(n16443), .ZN(n16444) );
  OAI211_X1 U19662 ( .C1(n19501), .C2(n19292), .A(n16445), .B(n16444), .ZN(
        P2_U3000) );
  AOI22_X1 U19663 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19517), .B1(n16494), 
        .B2(n19301), .ZN(n16456) );
  AOI21_X1 U19664 ( .B1(n16536), .B2(n16447), .A(n16446), .ZN(n16540) );
  NAND2_X1 U19665 ( .A1(n16449), .A2(n16448), .ZN(n16453) );
  NOR2_X1 U19666 ( .A1(n16451), .A2(n16450), .ZN(n16452) );
  XOR2_X1 U19667 ( .A(n16453), .B(n16452), .Z(n16543) );
  INV_X1 U19668 ( .A(n16543), .ZN(n16454) );
  AOI222_X1 U19669 ( .A1(n19507), .A2(n16540), .B1(n16454), .B2(n12279), .C1(
        n19512), .C2(n19306), .ZN(n16455) );
  OAI211_X1 U19670 ( .C1(n16457), .C2(n16506), .A(n16456), .B(n16455), .ZN(
        P2_U3001) );
  AOI22_X1 U19671 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19503), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19517), .ZN(n16462) );
  OAI22_X1 U19672 ( .A1(n16459), .A2(n19495), .B1(n16458), .B2(n19510), .ZN(
        n16460) );
  AOI21_X1 U19673 ( .B1(n19512), .B2(n19316), .A(n16460), .ZN(n16461) );
  OAI211_X1 U19674 ( .C1(n19501), .C2(n19314), .A(n16462), .B(n16461), .ZN(
        P2_U3002) );
  AOI22_X1 U19675 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19517), .B1(n16494), 
        .B2(n16463), .ZN(n16472) );
  NAND2_X1 U19676 ( .A1(n9943), .A2(n10186), .ZN(n16467) );
  NAND2_X1 U19677 ( .A1(n12163), .A2(n16465), .ZN(n16466) );
  XNOR2_X1 U19678 ( .A(n16467), .B(n16466), .ZN(n16550) );
  INV_X1 U19679 ( .A(n15724), .ZN(n16468) );
  AOI21_X1 U19680 ( .B1(n16468), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16470) );
  NOR2_X1 U19681 ( .A1(n16470), .A2(n16469), .ZN(n16548) );
  AOI222_X1 U19682 ( .A1(n16550), .A2(n12279), .B1(n19512), .B2(n16549), .C1(
        n19507), .C2(n16548), .ZN(n16471) );
  OAI211_X1 U19683 ( .C1(n16473), .C2(n16506), .A(n16472), .B(n16471), .ZN(
        P2_U3003) );
  AOI22_X1 U19684 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19503), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19517), .ZN(n16478) );
  OAI22_X1 U19685 ( .A1(n16475), .A2(n19495), .B1(n16474), .B2(n19510), .ZN(
        n16476) );
  AOI21_X1 U19686 ( .B1(n19512), .B2(n19407), .A(n16476), .ZN(n16477) );
  OAI211_X1 U19687 ( .C1(n19501), .C2(n19328), .A(n16478), .B(n16477), .ZN(
        P2_U3004) );
  AOI22_X1 U19688 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19517), .B1(n16494), 
        .B2(n16479), .ZN(n16485) );
  INV_X1 U19689 ( .A(n16480), .ZN(n16483) );
  AOI222_X1 U19690 ( .A1(n16483), .A2(n19507), .B1(n12279), .B2(n16482), .C1(
        n19512), .C2(n16481), .ZN(n16484) );
  OAI211_X1 U19691 ( .C1(n16486), .C2(n16506), .A(n16485), .B(n16484), .ZN(
        P2_U3005) );
  AOI22_X1 U19692 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19517), .B1(n16494), 
        .B2(n19347), .ZN(n16491) );
  AOI222_X1 U19693 ( .A1(n16489), .A2(n12279), .B1(n19512), .B2(n16488), .C1(
        n19507), .C2(n16487), .ZN(n16490) );
  OAI211_X1 U19694 ( .C1(n16492), .C2(n16506), .A(n16491), .B(n16490), .ZN(
        P2_U3007) );
  AOI22_X1 U19695 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19517), .B1(n16494), 
        .B2(n16493), .ZN(n16505) );
  XOR2_X1 U19696 ( .A(n16496), .B(n16495), .Z(n16579) );
  INV_X1 U19697 ( .A(n16497), .ZN(n16502) );
  AOI21_X1 U19698 ( .B1(n16501), .B2(n16499), .A(n16498), .ZN(n16500) );
  AOI21_X1 U19699 ( .B1(n16502), .B2(n16501), .A(n16500), .ZN(n16578) );
  INV_X1 U19700 ( .A(n16503), .ZN(n16576) );
  AOI222_X1 U19701 ( .A1(n16579), .A2(n12279), .B1(n16578), .B2(n19507), .C1(
        n19512), .C2(n16576), .ZN(n16504) );
  OAI211_X1 U19702 ( .C1(n16507), .C2(n16506), .A(n16505), .B(n16504), .ZN(
        P2_U3009) );
  AOI22_X1 U19703 ( .A1(n16509), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n19537), .B2(n16508), .ZN(n16519) );
  OAI22_X1 U19704 ( .A1(n16511), .A2(n16589), .B1(n19540), .B2(n16510), .ZN(
        n16512) );
  AOI21_X1 U19705 ( .B1(n16513), .B2(n16577), .A(n16512), .ZN(n16518) );
  NAND2_X1 U19706 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19517), .ZN(n16517) );
  OAI211_X1 U19707 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n16515), .B(n16514), .ZN(
        n16516) );
  NAND4_X1 U19708 ( .A1(n16519), .A2(n16518), .A3(n16517), .A4(n16516), .ZN(
        P2_U3023) );
  NAND2_X1 U19709 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19517), .ZN(n16521) );
  NAND2_X1 U19710 ( .A1(n19537), .A2(n19283), .ZN(n16520) );
  OAI211_X1 U19711 ( .C1(n16522), .C2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16521), .B(n16520), .ZN(n16523) );
  AOI21_X1 U19712 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16524), .A(
        n16523), .ZN(n16529) );
  INV_X1 U19713 ( .A(n16525), .ZN(n16527) );
  INV_X1 U19714 ( .A(n16526), .ZN(n19284) );
  AOI22_X1 U19715 ( .A1(n16527), .A2(n16577), .B1(n19560), .B2(n19284), .ZN(
        n16528) );
  OAI211_X1 U19716 ( .C1(n16589), .C2(n16530), .A(n16529), .B(n16528), .ZN(
        P2_U3031) );
  AOI21_X1 U19717 ( .B1(n16533), .B2(n16532), .A(n16531), .ZN(n19425) );
  INV_X1 U19718 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n20106) );
  NOR2_X1 U19719 ( .A1(n19350), .A2(n20106), .ZN(n16539) );
  OAI22_X1 U19720 ( .A1(n16537), .A2(n16536), .B1(n16535), .B2(n16534), .ZN(
        n16538) );
  AOI211_X1 U19721 ( .C1(n19537), .C2(n19425), .A(n16539), .B(n16538), .ZN(
        n16542) );
  AOI22_X1 U19722 ( .A1(n16540), .A2(n16577), .B1(n19560), .B2(n19306), .ZN(
        n16541) );
  OAI211_X1 U19723 ( .C1(n16589), .C2(n16543), .A(n16542), .B(n16541), .ZN(
        P2_U3033) );
  INV_X1 U19724 ( .A(n16544), .ZN(n16545) );
  OAI22_X1 U19725 ( .A1(n19554), .A2(n19431), .B1(n16546), .B2(n16545), .ZN(
        n16547) );
  INV_X1 U19726 ( .A(n16547), .ZN(n16556) );
  AOI222_X1 U19727 ( .A1(n16550), .A2(n19551), .B1(n19560), .B2(n16549), .C1(
        n16577), .C2(n16548), .ZN(n16555) );
  NAND2_X1 U19728 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19517), .ZN(n16554) );
  OAI211_X1 U19729 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n16552), .B(n16551), .ZN(
        n16553) );
  NAND4_X1 U19730 ( .A1(n16556), .A2(n16555), .A3(n16554), .A4(n16553), .ZN(
        P2_U3035) );
  OR2_X1 U19731 ( .A1(n16558), .A2(n16557), .ZN(n16560) );
  NAND2_X1 U19732 ( .A1(n16560), .A2(n16559), .ZN(n19436) );
  OAI21_X1 U19733 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16561), .ZN(n16563) );
  NAND2_X1 U19734 ( .A1(n19517), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n16562) );
  OAI211_X1 U19735 ( .C1(n19554), .C2(n19436), .A(n16563), .B(n16562), .ZN(
        n16564) );
  AOI21_X1 U19736 ( .B1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16565), .A(
        n16564), .ZN(n16569) );
  INV_X1 U19737 ( .A(n16566), .ZN(n16567) );
  AOI22_X1 U19738 ( .A1(n16567), .A2(n16577), .B1(n19560), .B2(n19341), .ZN(
        n16568) );
  OAI211_X1 U19739 ( .C1(n16570), .C2(n16589), .A(n16569), .B(n16568), .ZN(
        P2_U3038) );
  AOI211_X1 U19740 ( .C1(n19520), .C2(n16582), .A(n16571), .B(n19521), .ZN(
        n16575) );
  NAND2_X1 U19741 ( .A1(n16572), .A2(n19537), .ZN(n16573) );
  OAI21_X1 U19742 ( .B1(n10760), .B2(n19350), .A(n16573), .ZN(n16574) );
  NOR2_X1 U19743 ( .A1(n16575), .A2(n16574), .ZN(n16581) );
  AOI222_X1 U19744 ( .A1(n16579), .A2(n19551), .B1(n16578), .B2(n16577), .C1(
        n19560), .C2(n16576), .ZN(n16580) );
  OAI211_X1 U19745 ( .C1(n19519), .C2(n16582), .A(n16581), .B(n16580), .ZN(
        P2_U3041) );
  AOI22_X1 U19746 ( .A1(n19552), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19537), .B2(n16583), .ZN(n16592) );
  NOR2_X1 U19747 ( .A1(n19324), .A2(n10313), .ZN(n19505) );
  OAI21_X1 U19748 ( .B1(n19384), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n16584), .ZN(n19509) );
  NAND2_X1 U19749 ( .A1(n16586), .A2(n16585), .ZN(n16587) );
  NAND2_X1 U19750 ( .A1(n16588), .A2(n16587), .ZN(n19504) );
  OAI22_X1 U19751 ( .A1(n16589), .A2(n19509), .B1(n19556), .B2(n19504), .ZN(
        n16590) );
  AOI211_X1 U19752 ( .C1(n19560), .C2(n19513), .A(n19505), .B(n16590), .ZN(
        n16591) );
  OAI211_X1 U19753 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n16593), .A(
        n16592), .B(n16591), .ZN(P2_U3046) );
  NAND2_X1 U19754 ( .A1(n16595), .A2(n16620), .ZN(n16594) );
  OAI21_X1 U19755 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n16620), .A(
        n16594), .ZN(n16622) );
  INV_X1 U19756 ( .A(n16595), .ZN(n16600) );
  INV_X1 U19757 ( .A(n16620), .ZN(n16602) );
  AOI21_X1 U19758 ( .B1(n16597), .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n16602), .ZN(n16599) );
  OAI211_X1 U19759 ( .C1(n16597), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16596), .ZN(n16598) );
  OAI211_X1 U19760 ( .C1(n16600), .C2(n20156), .A(n16599), .B(n16598), .ZN(
        n16603) );
  NAND2_X1 U19761 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16603), .ZN(
        n16605) );
  AOI22_X1 U19762 ( .A1(n16602), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n16601), .B2(n16620), .ZN(n16621) );
  OAI22_X1 U19763 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16603), .B1(
        n16621), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n16604) );
  NAND2_X1 U19764 ( .A1(n16605), .A2(n16604), .ZN(n16606) );
  OAI21_X1 U19765 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16622), .A(
        n16606), .ZN(n16625) );
  INV_X1 U19766 ( .A(n16607), .ZN(n16610) );
  INV_X1 U19767 ( .A(n10646), .ZN(n16609) );
  OAI22_X1 U19768 ( .A1(n16612), .A2(n16610), .B1(n16609), .B2(n16608), .ZN(
        n16611) );
  AOI21_X1 U19769 ( .B1(n16613), .B2(n16612), .A(n16611), .ZN(n20191) );
  AOI21_X1 U19770 ( .B1(n16616), .B2(n16615), .A(n16614), .ZN(n16619) );
  OAI21_X1 U19771 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n16617), .ZN(n16618) );
  NAND3_X1 U19772 ( .A1(n20191), .A2(n16619), .A3(n16618), .ZN(n16624) );
  OAI22_X1 U19773 ( .A1(n16622), .A2(n16621), .B1(n12270), .B2(n16620), .ZN(
        n16623) );
  AOI211_X1 U19774 ( .C1(n16626), .C2(n16625), .A(n16624), .B(n16623), .ZN(
        n16640) );
  AOI211_X1 U19775 ( .C1(n16628), .C2(n16641), .A(n16627), .B(n20061), .ZN(
        n16638) );
  INV_X1 U19776 ( .A(n16629), .ZN(n16630) );
  NAND3_X1 U19777 ( .A1(n10692), .A2(n20205), .A3(n16630), .ZN(n16632) );
  NOR2_X1 U19778 ( .A1(n16631), .A2(n20065), .ZN(n20194) );
  NAND2_X1 U19779 ( .A1(n16632), .A2(n20194), .ZN(n16635) );
  NOR2_X1 U19780 ( .A1(n16635), .A2(n20202), .ZN(n20063) );
  AOI21_X1 U19781 ( .B1(n16634), .B2(n16633), .A(n20063), .ZN(n16636) );
  AOI21_X1 U19782 ( .B1(n15777), .B2(n16640), .A(n20201), .ZN(n20060) );
  OR2_X1 U19783 ( .A1(n20060), .A2(n16635), .ZN(n20068) );
  NAND2_X1 U19784 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20068), .ZN(n16642) );
  OAI21_X1 U19785 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16636), .A(n16642), 
        .ZN(n16637) );
  OAI211_X1 U19786 ( .C1(n16640), .C2(n16639), .A(n16638), .B(n16637), .ZN(
        P2_U3176) );
  AOI21_X1 U19787 ( .B1(n16642), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n16641), 
        .ZN(n16643) );
  INV_X1 U19788 ( .A(n16643), .ZN(P2_U3593) );
  AOI22_X1 U19789 ( .A1(n18136), .A2(n16662), .B1(n18008), .B2(n16657), .ZN(
        n16656) );
  XOR2_X1 U19790 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n9827), .Z(n16854) );
  OAI22_X2 U19791 ( .A1(n18345), .A2(n18152), .B1(n9662), .B2(n18009), .ZN(
        n18041) );
  OAI221_X1 U19792 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16650), .C1(
        n9931), .C2(n16649), .A(n16648), .ZN(n16651) );
  AOI211_X1 U19793 ( .C1(n18004), .C2(n16854), .A(n9787), .B(n16651), .ZN(
        n16654) );
  NAND2_X1 U19794 ( .A1(n18058), .A2(n16652), .ZN(n16653) );
  OAI211_X1 U19795 ( .C1(n16656), .C2(n16655), .A(n16654), .B(n16653), .ZN(
        P3_U2800) );
  NAND2_X1 U19796 ( .A1(n18008), .A2(n16657), .ZN(n16672) );
  NAND2_X1 U19797 ( .A1(n16658), .A2(n17802), .ZN(n16693) );
  AOI22_X1 U19798 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16661), .B1(
        n16660), .B2(n16659), .ZN(n16667) );
  NAND2_X1 U19799 ( .A1(n18408), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16666) );
  OAI211_X1 U19800 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16692), .A(
        n18136), .B(n16662), .ZN(n16665) );
  AOI21_X1 U19801 ( .B1(n9928), .B2(n16830), .A(n9827), .ZN(n16863) );
  OAI21_X1 U19802 ( .B1(n16663), .B2(n18004), .A(n16863), .ZN(n16664) );
  NAND4_X1 U19803 ( .A1(n16667), .A2(n16666), .A3(n16665), .A4(n16664), .ZN(
        n16668) );
  AOI21_X1 U19804 ( .B1(n18058), .B2(n16669), .A(n16668), .ZN(n16670) );
  OAI221_X1 U19805 ( .B1(n16672), .B2(n16671), .C1(n16672), .C2(n16693), .A(
        n16670), .ZN(P3_U2801) );
  NOR2_X1 U19806 ( .A1(n18385), .A2(n18460), .ZN(n18465) );
  NAND2_X1 U19807 ( .A1(n18153), .A2(n18178), .ZN(n16673) );
  OAI22_X1 U19808 ( .A1(n19135), .A2(n16675), .B1(n16674), .B2(n16673), .ZN(
        n16676) );
  AOI211_X1 U19809 ( .C1(n16678), .C2(n18465), .A(n16677), .B(n16676), .ZN(
        n16684) );
  INV_X1 U19810 ( .A(n16679), .ZN(n16680) );
  AOI21_X1 U19811 ( .B1(n16682), .B2(n18391), .A(n16681), .ZN(n16683) );
  OAI211_X1 U19812 ( .C1(n16685), .C2(n18468), .A(n16684), .B(n16683), .ZN(
        P3_U2831) );
  INV_X1 U19813 ( .A(n18953), .ZN(n18326) );
  INV_X1 U19814 ( .A(n16686), .ZN(n16699) );
  AOI22_X1 U19815 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18057), .B1(
        n17968), .B2(n17803), .ZN(n17807) );
  NAND2_X1 U19816 ( .A1(n17808), .A2(n17807), .ZN(n17806) );
  NAND4_X1 U19817 ( .A1(n16689), .A2(n16688), .A3(n16687), .A4(n17806), .ZN(
        n16690) );
  OAI211_X1 U19818 ( .C1(n16692), .C2(n18326), .A(n16691), .B(n16690), .ZN(
        n16694) );
  OAI221_X1 U19819 ( .B1(n16694), .B2(n18217), .C1(n16694), .C2(n16693), .A(
        n18375), .ZN(n16702) );
  INV_X1 U19820 ( .A(n18287), .ZN(n17873) );
  OAI21_X1 U19821 ( .B1(n17873), .B2(n18326), .A(n16695), .ZN(n18255) );
  NOR2_X1 U19822 ( .A1(n18178), .A2(n18255), .ZN(n18229) );
  NOR2_X1 U19823 ( .A1(n18229), .A2(n18158), .ZN(n18225) );
  NAND2_X1 U19824 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18225), .ZN(
        n18208) );
  NOR2_X1 U19825 ( .A1(n18460), .A2(n18208), .ZN(n18204) );
  NOR2_X1 U19826 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16696), .ZN(
        n17805) );
  NOR3_X1 U19827 ( .A1(n18458), .A2(n16697), .A3(n17808), .ZN(n16698) );
  INV_X1 U19828 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19103) );
  NOR2_X1 U19829 ( .A1(n18375), .A2(n19103), .ZN(n17801) );
  AOI211_X1 U19830 ( .C1(n18204), .C2(n17805), .A(n16698), .B(n17801), .ZN(
        n16701) );
  OAI211_X1 U19831 ( .C1(n17803), .C2(n16702), .A(n16701), .B(n16700), .ZN(
        P3_U2834) );
  NOR3_X1 U19832 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16704) );
  NOR4_X1 U19833 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16703) );
  INV_X2 U19834 ( .A(n16801), .ZN(U215) );
  NAND4_X1 U19835 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16704), .A3(n16703), .A4(
        U215), .ZN(U213) );
  INV_X1 U19836 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19438) );
  INV_X2 U19837 ( .A(U214), .ZN(n16765) );
  NOR2_X1 U19838 ( .A1(n16765), .A2(n16705), .ZN(n16707) );
  INV_X1 U19839 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16803) );
  OAI222_X1 U19840 ( .A1(U212), .A2(n19438), .B1(n16767), .B2(n16706), .C1(
        U214), .C2(n16803), .ZN(U216) );
  AOI222_X1 U19841 ( .A1(n16764), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16707), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n16765), .C2(P1_DATAO_REG_30__SCAN_IN), 
        .ZN(n16708) );
  INV_X1 U19842 ( .A(n16708), .ZN(U217) );
  INV_X1 U19843 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n19444) );
  INV_X1 U19844 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n16709) );
  OAI222_X1 U19845 ( .A1(U212), .A2(n19444), .B1(n16767), .B2(n16710), .C1(
        U214), .C2(n16709), .ZN(U218) );
  AOI22_X1 U19846 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16764), .ZN(n16711) );
  OAI21_X1 U19847 ( .B1(n16712), .B2(n16767), .A(n16711), .ZN(U219) );
  INV_X1 U19848 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16714) );
  AOI22_X1 U19849 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16764), .ZN(n16713) );
  OAI21_X1 U19850 ( .B1(n16714), .B2(n16767), .A(n16713), .ZN(U220) );
  AOI22_X1 U19851 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16764), .ZN(n16715) );
  OAI21_X1 U19852 ( .B1(n16716), .B2(n16767), .A(n16715), .ZN(U221) );
  AOI22_X1 U19853 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16764), .ZN(n16717) );
  OAI21_X1 U19854 ( .B1(n16718), .B2(n16767), .A(n16717), .ZN(U222) );
  INV_X1 U19855 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16720) );
  AOI22_X1 U19856 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16764), .ZN(n16719) );
  OAI21_X1 U19857 ( .B1(n16720), .B2(n16767), .A(n16719), .ZN(U223) );
  AOI22_X1 U19858 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16764), .ZN(n16721) );
  OAI21_X1 U19859 ( .B1(n16722), .B2(n16767), .A(n16721), .ZN(U224) );
  AOI22_X1 U19860 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16764), .ZN(n16723) );
  OAI21_X1 U19861 ( .B1(n16724), .B2(n16767), .A(n16723), .ZN(U225) );
  AOI22_X1 U19862 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16764), .ZN(n16725) );
  OAI21_X1 U19863 ( .B1(n15354), .B2(n16767), .A(n16725), .ZN(U226) );
  INV_X1 U19864 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16727) );
  AOI22_X1 U19865 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16764), .ZN(n16726) );
  OAI21_X1 U19866 ( .B1(n16727), .B2(n16767), .A(n16726), .ZN(U227) );
  AOI22_X1 U19867 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16764), .ZN(n16728) );
  OAI21_X1 U19868 ( .B1(n16729), .B2(n16767), .A(n16728), .ZN(U228) );
  INV_X1 U19869 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16731) );
  AOI22_X1 U19870 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16764), .ZN(n16730) );
  OAI21_X1 U19871 ( .B1(n16731), .B2(n16767), .A(n16730), .ZN(U229) );
  AOI22_X1 U19872 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16764), .ZN(n16732) );
  OAI21_X1 U19873 ( .B1(n14370), .B2(n16767), .A(n16732), .ZN(U230) );
  AOI22_X1 U19874 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16764), .ZN(n16733) );
  OAI21_X1 U19875 ( .B1(n16734), .B2(n16767), .A(n16733), .ZN(U231) );
  AOI22_X1 U19876 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16764), .ZN(n16735) );
  OAI21_X1 U19877 ( .B1(n13474), .B2(n16767), .A(n16735), .ZN(U232) );
  AOI22_X1 U19878 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16764), .ZN(n16736) );
  OAI21_X1 U19879 ( .B1(n16737), .B2(n16767), .A(n16736), .ZN(U233) );
  AOI22_X1 U19880 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16764), .ZN(n16738) );
  OAI21_X1 U19881 ( .B1(n16739), .B2(n16767), .A(n16738), .ZN(U234) );
  INV_X1 U19882 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16741) );
  AOI22_X1 U19883 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16764), .ZN(n16740) );
  OAI21_X1 U19884 ( .B1(n16741), .B2(n16767), .A(n16740), .ZN(U235) );
  AOI22_X1 U19885 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16764), .ZN(n16742) );
  OAI21_X1 U19886 ( .B1(n16743), .B2(n16767), .A(n16742), .ZN(U236) );
  AOI22_X1 U19887 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16764), .ZN(n16744) );
  OAI21_X1 U19888 ( .B1(n16745), .B2(n16767), .A(n16744), .ZN(U237) );
  AOI22_X1 U19889 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16764), .ZN(n16746) );
  OAI21_X1 U19890 ( .B1(n16747), .B2(n16767), .A(n16746), .ZN(U238) );
  AOI22_X1 U19891 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16764), .ZN(n16748) );
  OAI21_X1 U19892 ( .B1(n16749), .B2(n16767), .A(n16748), .ZN(U239) );
  AOI22_X1 U19893 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16764), .ZN(n16750) );
  OAI21_X1 U19894 ( .B1(n16751), .B2(n16767), .A(n16750), .ZN(U240) );
  AOI22_X1 U19895 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16764), .ZN(n16752) );
  OAI21_X1 U19896 ( .B1(n16753), .B2(n16767), .A(n16752), .ZN(U241) );
  INV_X1 U19897 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16755) );
  AOI22_X1 U19898 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16764), .ZN(n16754) );
  OAI21_X1 U19899 ( .B1(n16755), .B2(n16767), .A(n16754), .ZN(U242) );
  AOI22_X1 U19900 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16764), .ZN(n16756) );
  OAI21_X1 U19901 ( .B1(n16757), .B2(n16767), .A(n16756), .ZN(U243) );
  AOI22_X1 U19902 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16764), .ZN(n16758) );
  OAI21_X1 U19903 ( .B1(n16759), .B2(n16767), .A(n16758), .ZN(U244) );
  AOI22_X1 U19904 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16764), .ZN(n16760) );
  OAI21_X1 U19905 ( .B1(n16761), .B2(n16767), .A(n16760), .ZN(U245) );
  AOI22_X1 U19906 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16764), .ZN(n16762) );
  OAI21_X1 U19907 ( .B1(n16763), .B2(n16767), .A(n16762), .ZN(U246) );
  AOI22_X1 U19908 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16765), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16764), .ZN(n16766) );
  OAI21_X1 U19909 ( .B1(n16768), .B2(n16767), .A(n16766), .ZN(U247) );
  OAI22_X1 U19910 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16801), .ZN(n16769) );
  INV_X1 U19911 ( .A(n16769), .ZN(U251) );
  OAI22_X1 U19912 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16797), .ZN(n16770) );
  INV_X1 U19913 ( .A(n16770), .ZN(U252) );
  INV_X1 U19914 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16771) );
  INV_X1 U19915 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18502) );
  AOI22_X1 U19916 ( .A1(n16801), .A2(n16771), .B1(n18502), .B2(U215), .ZN(U253) );
  INV_X1 U19917 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16772) );
  INV_X1 U19918 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18507) );
  AOI22_X1 U19919 ( .A1(n16801), .A2(n16772), .B1(n18507), .B2(U215), .ZN(U254) );
  INV_X1 U19920 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16773) );
  INV_X1 U19921 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18513) );
  AOI22_X1 U19922 ( .A1(n16801), .A2(n16773), .B1(n18513), .B2(U215), .ZN(U255) );
  INV_X1 U19923 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16774) );
  INV_X1 U19924 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18518) );
  AOI22_X1 U19925 ( .A1(n16801), .A2(n16774), .B1(n18518), .B2(U215), .ZN(U256) );
  INV_X1 U19926 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16775) );
  INV_X1 U19927 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18524) );
  AOI22_X1 U19928 ( .A1(n16801), .A2(n16775), .B1(n18524), .B2(U215), .ZN(U257) );
  INV_X1 U19929 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16776) );
  INV_X1 U19930 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18529) );
  AOI22_X1 U19931 ( .A1(n16797), .A2(n16776), .B1(n18529), .B2(U215), .ZN(U258) );
  INV_X1 U19932 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16777) );
  AOI22_X1 U19933 ( .A1(n16797), .A2(n16777), .B1(n17655), .B2(U215), .ZN(U259) );
  INV_X1 U19934 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16778) );
  INV_X1 U19935 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17650) );
  AOI22_X1 U19936 ( .A1(n16797), .A2(n16778), .B1(n17650), .B2(U215), .ZN(U260) );
  OAI22_X1 U19937 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16801), .ZN(n16779) );
  INV_X1 U19938 ( .A(n16779), .ZN(U261) );
  INV_X1 U19939 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16780) );
  INV_X1 U19940 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17639) );
  AOI22_X1 U19941 ( .A1(n16801), .A2(n16780), .B1(n17639), .B2(U215), .ZN(U262) );
  INV_X1 U19942 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16781) );
  INV_X1 U19943 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17635) );
  AOI22_X1 U19944 ( .A1(n16801), .A2(n16781), .B1(n17635), .B2(U215), .ZN(U263) );
  INV_X1 U19945 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16782) );
  INV_X1 U19946 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17630) );
  AOI22_X1 U19947 ( .A1(n16797), .A2(n16782), .B1(n17630), .B2(U215), .ZN(U264) );
  OAI22_X1 U19948 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16801), .ZN(n16783) );
  INV_X1 U19949 ( .A(n16783), .ZN(U265) );
  OAI22_X1 U19950 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16801), .ZN(n16784) );
  INV_X1 U19951 ( .A(n16784), .ZN(U266) );
  OAI22_X1 U19952 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16801), .ZN(n16785) );
  INV_X1 U19953 ( .A(n16785), .ZN(U267) );
  OAI22_X1 U19954 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16801), .ZN(n16786) );
  INV_X1 U19955 ( .A(n16786), .ZN(U268) );
  OAI22_X1 U19956 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16801), .ZN(n16787) );
  INV_X1 U19957 ( .A(n16787), .ZN(U269) );
  OAI22_X1 U19958 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16797), .ZN(n16788) );
  INV_X1 U19959 ( .A(n16788), .ZN(U270) );
  OAI22_X1 U19960 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16801), .ZN(n16789) );
  INV_X1 U19961 ( .A(n16789), .ZN(U271) );
  OAI22_X1 U19962 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16801), .ZN(n16790) );
  INV_X1 U19963 ( .A(n16790), .ZN(U272) );
  OAI22_X1 U19964 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16801), .ZN(n16791) );
  INV_X1 U19965 ( .A(n16791), .ZN(U273) );
  OAI22_X1 U19966 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16797), .ZN(n16792) );
  INV_X1 U19967 ( .A(n16792), .ZN(U274) );
  OAI22_X1 U19968 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16797), .ZN(n16793) );
  INV_X1 U19969 ( .A(n16793), .ZN(U275) );
  INV_X1 U19970 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n16794) );
  INV_X1 U19971 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18497) );
  AOI22_X1 U19972 ( .A1(n16801), .A2(n16794), .B1(n18497), .B2(U215), .ZN(U276) );
  OAI22_X1 U19973 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16797), .ZN(n16795) );
  INV_X1 U19974 ( .A(n16795), .ZN(U277) );
  INV_X1 U19975 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n16796) );
  INV_X1 U19976 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n18508) );
  AOI22_X1 U19977 ( .A1(n16801), .A2(n16796), .B1(n18508), .B2(U215), .ZN(U278) );
  OAI22_X1 U19978 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16797), .ZN(n16798) );
  INV_X1 U19979 ( .A(n16798), .ZN(U279) );
  INV_X1 U19980 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18519) );
  AOI22_X1 U19981 ( .A1(n16801), .A2(n19444), .B1(n18519), .B2(U215), .ZN(U280) );
  INV_X1 U19982 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19441) );
  INV_X1 U19983 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n16800) );
  AOI22_X1 U19984 ( .A1(n16801), .A2(n19441), .B1(n16800), .B2(U215), .ZN(U281) );
  INV_X1 U19985 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18531) );
  AOI22_X1 U19986 ( .A1(n16801), .A2(n19438), .B1(n18531), .B2(U215), .ZN(U282) );
  INV_X1 U19987 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16802) );
  AOI222_X1 U19988 ( .A1(n16803), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19438), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16802), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16804) );
  INV_X2 U19989 ( .A(n16806), .ZN(n16805) );
  INV_X1 U19990 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19066) );
  INV_X1 U19991 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20102) );
  AOI22_X1 U19992 ( .A1(n16805), .A2(n19066), .B1(n20102), .B2(n16806), .ZN(
        U347) );
  INV_X1 U19993 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19064) );
  INV_X1 U19994 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20101) );
  AOI22_X1 U19995 ( .A1(n16805), .A2(n19064), .B1(n20101), .B2(n16806), .ZN(
        U348) );
  INV_X1 U19996 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19062) );
  INV_X1 U19997 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20100) );
  AOI22_X1 U19998 ( .A1(n16805), .A2(n19062), .B1(n20100), .B2(n16806), .ZN(
        U349) );
  INV_X1 U19999 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19060) );
  INV_X1 U20000 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20099) );
  AOI22_X1 U20001 ( .A1(n16805), .A2(n19060), .B1(n20099), .B2(n16806), .ZN(
        U350) );
  INV_X1 U20002 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19058) );
  INV_X1 U20003 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20097) );
  AOI22_X1 U20004 ( .A1(n16805), .A2(n19058), .B1(n20097), .B2(n16806), .ZN(
        U351) );
  INV_X1 U20005 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19055) );
  INV_X1 U20006 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20095) );
  AOI22_X1 U20007 ( .A1(n16805), .A2(n19055), .B1(n20095), .B2(n16806), .ZN(
        U352) );
  INV_X1 U20008 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19054) );
  INV_X1 U20009 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20094) );
  AOI22_X1 U20010 ( .A1(n16805), .A2(n19054), .B1(n20094), .B2(n16806), .ZN(
        U353) );
  INV_X1 U20011 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19052) );
  AOI22_X1 U20012 ( .A1(n16805), .A2(n19052), .B1(n20093), .B2(n16806), .ZN(
        U354) );
  INV_X1 U20013 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19105) );
  INV_X1 U20014 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20130) );
  AOI22_X1 U20015 ( .A1(n16805), .A2(n19105), .B1(n20130), .B2(n16806), .ZN(
        U356) );
  INV_X1 U20016 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19102) );
  INV_X1 U20017 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20129) );
  AOI22_X1 U20018 ( .A1(n16805), .A2(n19102), .B1(n20129), .B2(n16806), .ZN(
        U357) );
  INV_X1 U20019 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19100) );
  INV_X1 U20020 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20126) );
  AOI22_X1 U20021 ( .A1(n16805), .A2(n19100), .B1(n20126), .B2(n16806), .ZN(
        U358) );
  INV_X1 U20022 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19098) );
  INV_X1 U20023 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20125) );
  AOI22_X1 U20024 ( .A1(n16805), .A2(n19098), .B1(n20125), .B2(n16806), .ZN(
        U359) );
  INV_X1 U20025 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19096) );
  INV_X1 U20026 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20123) );
  AOI22_X1 U20027 ( .A1(n16805), .A2(n19096), .B1(n20123), .B2(n16806), .ZN(
        U360) );
  INV_X1 U20028 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19094) );
  INV_X1 U20029 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20121) );
  AOI22_X1 U20030 ( .A1(n16805), .A2(n19094), .B1(n20121), .B2(n16806), .ZN(
        U361) );
  INV_X1 U20031 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19091) );
  INV_X1 U20032 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20120) );
  AOI22_X1 U20033 ( .A1(n16805), .A2(n19091), .B1(n20120), .B2(n16806), .ZN(
        U362) );
  INV_X1 U20034 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19090) );
  INV_X1 U20035 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20119) );
  AOI22_X1 U20036 ( .A1(n16805), .A2(n19090), .B1(n20119), .B2(n16806), .ZN(
        U363) );
  INV_X1 U20037 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19087) );
  INV_X1 U20038 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20118) );
  AOI22_X1 U20039 ( .A1(n16805), .A2(n19087), .B1(n20118), .B2(n16806), .ZN(
        U364) );
  INV_X1 U20040 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19050) );
  INV_X1 U20041 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20092) );
  AOI22_X1 U20042 ( .A1(n16805), .A2(n19050), .B1(n20092), .B2(n16806), .ZN(
        U365) );
  INV_X1 U20043 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19086) );
  INV_X1 U20044 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20116) );
  AOI22_X1 U20045 ( .A1(n16805), .A2(n19086), .B1(n20116), .B2(n16806), .ZN(
        U366) );
  INV_X1 U20046 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19083) );
  INV_X1 U20047 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20114) );
  AOI22_X1 U20048 ( .A1(n16805), .A2(n19083), .B1(n20114), .B2(n16806), .ZN(
        U367) );
  INV_X1 U20049 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19082) );
  INV_X1 U20050 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20113) );
  AOI22_X1 U20051 ( .A1(n16805), .A2(n19082), .B1(n20113), .B2(n16806), .ZN(
        U368) );
  INV_X1 U20052 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19080) );
  INV_X1 U20053 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20111) );
  AOI22_X1 U20054 ( .A1(n16805), .A2(n19080), .B1(n20111), .B2(n16806), .ZN(
        U369) );
  INV_X1 U20055 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19078) );
  INV_X1 U20056 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20110) );
  AOI22_X1 U20057 ( .A1(n16805), .A2(n19078), .B1(n20110), .B2(n16806), .ZN(
        U370) );
  INV_X1 U20058 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19076) );
  INV_X1 U20059 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20109) );
  AOI22_X1 U20060 ( .A1(n16805), .A2(n19076), .B1(n20109), .B2(n16806), .ZN(
        U371) );
  INV_X1 U20061 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19073) );
  INV_X1 U20062 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20108) );
  AOI22_X1 U20063 ( .A1(n16805), .A2(n19073), .B1(n20108), .B2(n16806), .ZN(
        U372) );
  INV_X1 U20064 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19072) );
  INV_X1 U20065 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20107) );
  AOI22_X1 U20066 ( .A1(n16805), .A2(n19072), .B1(n20107), .B2(n16806), .ZN(
        U373) );
  INV_X1 U20067 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19070) );
  INV_X1 U20068 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20105) );
  AOI22_X1 U20069 ( .A1(n16805), .A2(n19070), .B1(n20105), .B2(n16806), .ZN(
        U374) );
  INV_X1 U20070 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19068) );
  INV_X1 U20071 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20103) );
  AOI22_X1 U20072 ( .A1(n16805), .A2(n19068), .B1(n20103), .B2(n16806), .ZN(
        U375) );
  INV_X1 U20073 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19048) );
  INV_X1 U20074 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20091) );
  AOI22_X1 U20075 ( .A1(n16805), .A2(n19048), .B1(n20091), .B2(n16806), .ZN(
        U376) );
  INV_X1 U20076 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16807) );
  INV_X1 U20077 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19047) );
  NAND2_X1 U20078 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19047), .ZN(n19036) );
  AOI22_X1 U20079 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19036), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n19045), .ZN(n19122) );
  OAI21_X1 U20080 ( .B1(n19045), .B2(n16807), .A(n19119), .ZN(P3_U2633) );
  INV_X1 U20081 ( .A(n16814), .ZN(n16808) );
  OAI21_X1 U20082 ( .B1(n16808), .B2(n17727), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16809) );
  OAI21_X1 U20083 ( .B1(n16810), .B2(n19025), .A(n16809), .ZN(P3_U2634) );
  AOI21_X1 U20084 ( .B1(n19045), .B2(n19047), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16811) );
  AOI22_X1 U20085 ( .A1(n19116), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16811), 
        .B2(n19181), .ZN(P3_U2635) );
  NOR2_X1 U20086 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n19032) );
  OAI21_X1 U20087 ( .B1(n19032), .B2(BS16), .A(n19122), .ZN(n19120) );
  OAI21_X1 U20088 ( .B1(n19122), .B2(n16812), .A(n19120), .ZN(P3_U2636) );
  AND3_X1 U20089 ( .A1(n16814), .A2(n18955), .A3(n16813), .ZN(n18960) );
  NOR2_X1 U20090 ( .A1(n18960), .A2(n19020), .ZN(n19163) );
  OAI21_X1 U20091 ( .B1(n19163), .B2(n18481), .A(n16815), .ZN(P3_U2637) );
  NOR4_X1 U20092 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16819) );
  NOR4_X1 U20093 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16818) );
  NOR4_X1 U20094 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16817) );
  NOR4_X1 U20095 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16816) );
  NAND4_X1 U20096 ( .A1(n16819), .A2(n16818), .A3(n16817), .A4(n16816), .ZN(
        n16825) );
  NOR4_X1 U20097 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16823) );
  AOI211_X1 U20098 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16822) );
  NOR4_X1 U20099 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16821) );
  NOR4_X1 U20100 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16820) );
  NAND4_X1 U20101 ( .A1(n16823), .A2(n16822), .A3(n16821), .A4(n16820), .ZN(
        n16824) );
  NOR2_X1 U20102 ( .A1(n16825), .A2(n16824), .ZN(n19157) );
  INV_X1 U20103 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19114) );
  NOR3_X1 U20104 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16827) );
  OAI21_X1 U20105 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16827), .A(n19157), .ZN(
        n16826) );
  OAI21_X1 U20106 ( .B1(n19157), .B2(n19114), .A(n16826), .ZN(P3_U2638) );
  INV_X1 U20107 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19121) );
  AOI21_X1 U20108 ( .B1(n19153), .B2(n19121), .A(n16827), .ZN(n16828) );
  INV_X1 U20109 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19111) );
  INV_X1 U20110 ( .A(n19157), .ZN(n19160) );
  AOI22_X1 U20111 ( .A1(n19157), .A2(n16828), .B1(n19111), .B2(n19160), .ZN(
        P3_U2639) );
  INV_X1 U20112 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19108) );
  INV_X1 U20113 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19099) );
  INV_X1 U20114 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19097) );
  INV_X1 U20115 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19092) );
  INV_X1 U20116 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19088) );
  INV_X1 U20117 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19081) );
  INV_X1 U20118 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19074) );
  INV_X1 U20119 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19069) );
  INV_X1 U20120 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19056) );
  AND2_X1 U20121 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n17167), .ZN(n17164) );
  NAND2_X1 U20122 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17164), .ZN(n17065) );
  NOR2_X1 U20123 ( .A1(n19056), .A2(n17065), .ZN(n17043) );
  INV_X1 U20124 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19067) );
  INV_X1 U20125 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19063) );
  NAND3_X1 U20126 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(P3_REIP_REG_6__SCAN_IN), .ZN(n17079) );
  NOR2_X1 U20127 ( .A1(n19063), .A2(n17079), .ZN(n17081) );
  NAND2_X1 U20128 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n17081), .ZN(n17066) );
  NOR2_X1 U20129 ( .A1(n19067), .A2(n17066), .ZN(n17044) );
  NAND2_X1 U20130 ( .A1(n17043), .A2(n17044), .ZN(n17057) );
  NOR2_X1 U20131 ( .A1(n19069), .A2(n17057), .ZN(n17045) );
  NAND2_X1 U20132 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17045), .ZN(n16991) );
  NOR2_X1 U20133 ( .A1(n19074), .A2(n16991), .ZN(n17003) );
  NAND4_X1 U20134 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n17003), .A3(
        P3_REIP_REG_16__SCAN_IN), .A4(P3_REIP_REG_15__SCAN_IN), .ZN(n16976) );
  NOR2_X1 U20135 ( .A1(n19081), .A2(n16976), .ZN(n16972) );
  AND2_X1 U20136 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16972), .ZN(n16955) );
  NAND2_X1 U20137 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16955), .ZN(n16953) );
  INV_X1 U20138 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19089) );
  NOR4_X1 U20139 ( .A1(n19092), .A2(n19088), .A3(n16953), .A4(n19089), .ZN(
        n16915) );
  AND2_X1 U20140 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16915), .ZN(n16909) );
  NAND2_X1 U20141 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16909), .ZN(n16902) );
  NOR2_X1 U20142 ( .A1(n19097), .A2(n16902), .ZN(n16844) );
  NAND2_X1 U20143 ( .A1(n17155), .A2(n16844), .ZN(n16886) );
  NOR2_X1 U20144 ( .A1(n19099), .A2(n16886), .ZN(n16872) );
  NAND3_X1 U20145 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(n16872), .ZN(n16846) );
  NOR3_X1 U20146 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19108), .A3(n16846), 
        .ZN(n16829) );
  AOI21_X1 U20147 ( .B1(n17194), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16829), .ZN(
        n16851) );
  NAND2_X1 U20148 ( .A1(n17175), .A2(n17513), .ZN(n17174) );
  NOR2_X1 U20149 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17174), .ZN(n17153) );
  NAND2_X1 U20150 ( .A1(n17153), .A2(n17143), .ZN(n17142) );
  INV_X1 U20151 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17499) );
  NAND2_X1 U20152 ( .A1(n17120), .A2(n17499), .ZN(n17116) );
  NAND2_X1 U20153 ( .A1(n17088), .A2(n17442), .ZN(n17076) );
  NAND2_X1 U20154 ( .A1(n17075), .A2(n17071), .ZN(n17070) );
  NAND2_X1 U20155 ( .A1(n17053), .A2(n17389), .ZN(n17046) );
  NAND2_X1 U20156 ( .A1(n17027), .A2(n17022), .ZN(n17019) );
  NOR2_X1 U20157 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17019), .ZN(n17001) );
  INV_X1 U20158 ( .A(n17001), .ZN(n16994) );
  INV_X1 U20159 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16975) );
  NAND2_X1 U20160 ( .A1(n16987), .A2(n16975), .ZN(n16967) );
  NAND2_X1 U20161 ( .A1(n16958), .A2(n16948), .ZN(n16947) );
  NAND2_X1 U20162 ( .A1(n16933), .A2(n16928), .ZN(n16927) );
  NAND2_X1 U20163 ( .A1(n16916), .A2(n16908), .ZN(n16907) );
  NOR2_X1 U20164 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16907), .ZN(n16893) );
  NAND2_X1 U20165 ( .A1(n16893), .A2(n17202), .ZN(n16889) );
  NOR2_X1 U20166 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16889), .ZN(n16873) );
  INV_X1 U20167 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17242) );
  NAND2_X1 U20168 ( .A1(n16873), .A2(n17242), .ZN(n16852) );
  NOR2_X1 U20169 ( .A1(n17192), .A2(n16852), .ZN(n16858) );
  INV_X1 U20170 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17208) );
  INV_X1 U20171 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16885) );
  NOR2_X1 U20172 ( .A1(n16832), .A2(n16885), .ZN(n16831) );
  OAI21_X1 U20173 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16831), .A(
        n16830), .ZN(n17799) );
  INV_X1 U20174 ( .A(n17799), .ZN(n16876) );
  AOI21_X1 U20175 ( .B1(n16832), .B2(n16885), .A(n16831), .ZN(n17814) );
  NAND2_X1 U20176 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9820), .ZN(
        n17835) );
  NOR2_X1 U20177 ( .A1(n9923), .A2(n17835), .ZN(n16837) );
  INV_X1 U20178 ( .A(n16837), .ZN(n16836) );
  NOR2_X1 U20179 ( .A1(n17837), .A2(n16836), .ZN(n17794) );
  OAI21_X1 U20180 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17794), .A(
        n16832), .ZN(n16833) );
  INV_X1 U20181 ( .A(n16833), .ZN(n17830) );
  INV_X1 U20182 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17853) );
  NOR2_X1 U20183 ( .A1(n17853), .A2(n16836), .ZN(n16835) );
  INV_X1 U20184 ( .A(n17794), .ZN(n16834) );
  OAI21_X1 U20185 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16835), .A(
        n16834), .ZN(n17839) );
  INV_X1 U20186 ( .A(n17839), .ZN(n16905) );
  OAI22_X1 U20187 ( .A1(n17853), .A2(n16837), .B1(n16836), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17849) );
  AOI21_X1 U20188 ( .B1(n9923), .B2(n17835), .A(n16837), .ZN(n17861) );
  INV_X1 U20189 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17892) );
  OR2_X1 U20190 ( .A1(n18143), .A2(n17877), .ZN(n16840) );
  NOR2_X1 U20191 ( .A1(n17892), .A2(n16840), .ZN(n16838) );
  OAI21_X1 U20192 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n16838), .A(
        n17835), .ZN(n16839) );
  INV_X1 U20193 ( .A(n16839), .ZN(n17876) );
  XNOR2_X1 U20194 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n16840), .ZN(
        n17888) );
  NAND3_X1 U20195 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9797), .A3(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16988) );
  NOR2_X1 U20196 ( .A1(n17913), .A2(n16988), .ZN(n17874) );
  OAI21_X1 U20197 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17874), .A(
        n16840), .ZN(n16841) );
  INV_X1 U20198 ( .A(n16841), .ZN(n17904) );
  INV_X1 U20199 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17137) );
  NAND2_X1 U20200 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18086), .ZN(
        n17148) );
  NOR2_X1 U20201 ( .A1(n17137), .A2(n17148), .ZN(n17135) );
  NAND2_X1 U20202 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17135), .ZN(
        n17127) );
  NOR2_X1 U20203 ( .A1(n16842), .A2(n17127), .ZN(n17062) );
  NAND3_X1 U20204 ( .A1(n17984), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A3(
        n17062), .ZN(n17016) );
  INV_X1 U20205 ( .A(n17016), .ZN(n17944) );
  NAND2_X1 U20206 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17944), .ZN(
        n17015) );
  NOR2_X1 U20207 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17015), .ZN(
        n17005) );
  AND2_X1 U20208 ( .A1(n17005), .A2(n17874), .ZN(n16843) );
  NOR2_X1 U20209 ( .A1(n17904), .A2(n16957), .ZN(n16956) );
  NOR2_X1 U20210 ( .A1(n16956), .A2(n17182), .ZN(n16944) );
  NOR2_X1 U20211 ( .A1(n16943), .A2(n17182), .ZN(n16935) );
  NOR2_X1 U20212 ( .A1(n16934), .A2(n17182), .ZN(n16924) );
  NOR2_X1 U20213 ( .A1(n17861), .A2(n16924), .ZN(n16923) );
  NOR2_X1 U20214 ( .A1(n16923), .A2(n17182), .ZN(n16918) );
  NOR2_X1 U20215 ( .A1(n16917), .A2(n17182), .ZN(n16904) );
  NOR2_X1 U20216 ( .A1(n16905), .A2(n16904), .ZN(n16903) );
  NOR2_X1 U20217 ( .A1(n16903), .A2(n17182), .ZN(n16895) );
  NOR2_X1 U20218 ( .A1(n16894), .A2(n17182), .ZN(n16884) );
  NOR2_X1 U20219 ( .A1(n17814), .A2(n16884), .ZN(n16883) );
  NOR2_X1 U20220 ( .A1(n16883), .A2(n17182), .ZN(n16875) );
  NOR2_X1 U20221 ( .A1(n16874), .A2(n17182), .ZN(n16862) );
  NOR2_X1 U20222 ( .A1(n16861), .A2(n17182), .ZN(n16853) );
  NOR4_X1 U20223 ( .A1(n16854), .A2(n16853), .A3(n17182), .A4(n19028), .ZN(
        n16849) );
  NAND2_X1 U20224 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .ZN(n16845) );
  OR2_X1 U20225 ( .A1(n17187), .A2(n16844), .ZN(n16901) );
  NAND2_X1 U20226 ( .A1(n17196), .A2(n16901), .ZN(n16898) );
  AOI221_X1 U20227 ( .B1(n19099), .B2(n17155), .C1(n16845), .C2(n17155), .A(
        n16898), .ZN(n16871) );
  NOR2_X1 U20228 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16846), .ZN(n16856) );
  INV_X1 U20229 ( .A(n16856), .ZN(n16847) );
  AOI21_X1 U20230 ( .B1(n16871), .B2(n16847), .A(n19106), .ZN(n16848) );
  AOI211_X1 U20231 ( .C1(n16858), .C2(n17208), .A(n16849), .B(n16848), .ZN(
        n16850) );
  OAI211_X1 U20232 ( .C1(n9929), .C2(n17159), .A(n16851), .B(n16850), .ZN(
        P3_U2640) );
  NAND2_X1 U20233 ( .A1(n17193), .A2(n16852), .ZN(n16867) );
  XOR2_X1 U20234 ( .A(n16854), .B(n16853), .Z(n16857) );
  OAI22_X1 U20235 ( .A1(n16871), .A2(n19108), .B1(n9931), .B2(n17159), .ZN(
        n16855) );
  OAI21_X1 U20236 ( .B1(n17194), .B2(n16858), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16859) );
  INV_X1 U20237 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19104) );
  AOI211_X1 U20238 ( .C1(n16863), .C2(n16862), .A(n16861), .B(n19028), .ZN(
        n16866) );
  NAND2_X1 U20239 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n16872), .ZN(n16864) );
  OAI22_X1 U20240 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16864), .B1(n9928), 
        .B2(n17159), .ZN(n16865) );
  AOI211_X1 U20241 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n17194), .A(n16866), .B(
        n16865), .ZN(n16870) );
  INV_X1 U20242 ( .A(n16867), .ZN(n16868) );
  OAI21_X1 U20243 ( .B1(n16873), .B2(n17242), .A(n16868), .ZN(n16869) );
  OAI211_X1 U20244 ( .C1(n16871), .C2(n19104), .A(n16870), .B(n16869), .ZN(
        P3_U2642) );
  INV_X1 U20245 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16882) );
  AOI22_X1 U20246 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17194), .B1(n16872), 
        .B2(n19103), .ZN(n16881) );
  INV_X1 U20247 ( .A(n16898), .ZN(n16892) );
  OAI21_X1 U20248 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16886), .A(n16892), 
        .ZN(n16879) );
  AOI211_X1 U20249 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16889), .A(n16873), .B(
        n17192), .ZN(n16878) );
  AOI211_X1 U20250 ( .C1(n16876), .C2(n16875), .A(n16874), .B(n19028), .ZN(
        n16877) );
  AOI211_X1 U20251 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16879), .A(n16878), 
        .B(n16877), .ZN(n16880) );
  OAI211_X1 U20252 ( .C1(n16882), .C2(n17159), .A(n16881), .B(n16880), .ZN(
        P3_U2643) );
  AOI211_X1 U20253 ( .C1(n17814), .C2(n16884), .A(n16883), .B(n19028), .ZN(
        n16888) );
  OAI22_X1 U20254 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16886), .B1(n16885), 
        .B2(n17159), .ZN(n16887) );
  AOI211_X1 U20255 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n17194), .A(n16888), .B(
        n16887), .ZN(n16891) );
  OAI211_X1 U20256 ( .C1(n16893), .C2(n17202), .A(n17193), .B(n16889), .ZN(
        n16890) );
  OAI211_X1 U20257 ( .C1(n16892), .C2(n19099), .A(n16891), .B(n16890), .ZN(
        P3_U2644) );
  AOI22_X1 U20258 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17183), .B1(
        n17194), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16900) );
  AOI211_X1 U20259 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16907), .A(n16893), .B(
        n17192), .ZN(n16897) );
  AOI211_X1 U20260 ( .C1(n17830), .C2(n16895), .A(n16894), .B(n19028), .ZN(
        n16896) );
  AOI211_X1 U20261 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16898), .A(n16897), 
        .B(n16896), .ZN(n16899) );
  OAI211_X1 U20262 ( .C1(n16902), .C2(n16901), .A(n16900), .B(n16899), .ZN(
        P3_U2645) );
  AOI22_X1 U20263 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17183), .B1(
        n17194), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n16913) );
  OAI21_X1 U20264 ( .B1(n16915), .B2(n17187), .A(n17196), .ZN(n16926) );
  NOR2_X1 U20265 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17187), .ZN(n16914) );
  AOI211_X1 U20266 ( .C1(n16905), .C2(n16904), .A(n16903), .B(n19028), .ZN(
        n16906) );
  AOI221_X1 U20267 ( .B1(n16926), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n16914), 
        .C2(P3_REIP_REG_25__SCAN_IN), .A(n16906), .ZN(n16912) );
  OAI211_X1 U20268 ( .C1(n16916), .C2(n16908), .A(n17193), .B(n16907), .ZN(
        n16911) );
  INV_X1 U20269 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19095) );
  NAND3_X1 U20270 ( .A1(n17155), .A2(n16909), .A3(n19095), .ZN(n16910) );
  NAND4_X1 U20271 ( .A1(n16913), .A2(n16912), .A3(n16911), .A4(n16910), .ZN(
        P3_U2646) );
  AOI22_X1 U20272 ( .A1(n17194), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16915), 
        .B2(n16914), .ZN(n16922) );
  AOI211_X1 U20273 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16927), .A(n16916), .B(
        n17192), .ZN(n16920) );
  AOI211_X1 U20274 ( .C1(n17849), .C2(n16918), .A(n16917), .B(n19028), .ZN(
        n16919) );
  AOI211_X1 U20275 ( .C1(n16926), .C2(P3_REIP_REG_24__SCAN_IN), .A(n16920), 
        .B(n16919), .ZN(n16921) );
  OAI211_X1 U20276 ( .C1(n17853), .C2(n17159), .A(n16922), .B(n16921), .ZN(
        P3_U2647) );
  AOI22_X1 U20277 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17183), .B1(
        n17194), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n16932) );
  AOI211_X1 U20278 ( .C1(n17861), .C2(n16924), .A(n16923), .B(n19028), .ZN(
        n16925) );
  AOI21_X1 U20279 ( .B1(n16926), .B2(P3_REIP_REG_23__SCAN_IN), .A(n16925), 
        .ZN(n16931) );
  OAI211_X1 U20280 ( .C1(n16933), .C2(n16928), .A(n17193), .B(n16927), .ZN(
        n16930) );
  NOR2_X1 U20281 ( .A1(n17187), .A2(n16953), .ZN(n16939) );
  NAND4_X1 U20282 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .A3(n16939), .A4(n19092), .ZN(n16929) );
  NAND4_X1 U20283 ( .A1(n16932), .A2(n16931), .A3(n16930), .A4(n16929), .ZN(
        P3_U2648) );
  AOI22_X1 U20284 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17183), .B1(
        n17194), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16942) );
  AOI211_X1 U20285 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16947), .A(n16933), .B(
        n17192), .ZN(n16938) );
  AOI21_X1 U20286 ( .B1(n17155), .B2(n16953), .A(n17181), .ZN(n16963) );
  NAND2_X1 U20287 ( .A1(n16939), .A2(n19088), .ZN(n16950) );
  AOI21_X1 U20288 ( .B1(n16963), .B2(n16950), .A(n19089), .ZN(n16937) );
  AOI211_X1 U20289 ( .C1(n17876), .C2(n16935), .A(n16934), .B(n19028), .ZN(
        n16936) );
  NOR3_X1 U20290 ( .A1(n16938), .A2(n16937), .A3(n16936), .ZN(n16941) );
  NAND3_X1 U20291 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16939), .A3(n19089), 
        .ZN(n16940) );
  NAND3_X1 U20292 ( .A1(n16942), .A2(n16941), .A3(n16940), .ZN(P3_U2649) );
  AOI22_X1 U20293 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17183), .B1(
        n17194), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n16952) );
  INV_X1 U20294 ( .A(n16963), .ZN(n16946) );
  AOI211_X1 U20295 ( .C1(n17888), .C2(n16944), .A(n16943), .B(n19028), .ZN(
        n16945) );
  AOI21_X1 U20296 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16946), .A(n16945), 
        .ZN(n16951) );
  OAI211_X1 U20297 ( .C1(n16958), .C2(n16948), .A(n17193), .B(n16947), .ZN(
        n16949) );
  NAND4_X1 U20298 ( .A1(n16952), .A2(n16951), .A3(n16950), .A4(n16949), .ZN(
        P3_U2650) );
  INV_X1 U20299 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19085) );
  AND2_X1 U20300 ( .A1(n16953), .A2(n17155), .ZN(n16954) );
  AOI22_X1 U20301 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17183), .B1(
        n16955), .B2(n16954), .ZN(n16962) );
  AOI211_X1 U20302 ( .C1(n17904), .C2(n16957), .A(n16956), .B(n19028), .ZN(
        n16960) );
  AOI211_X1 U20303 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16967), .A(n16958), .B(
        n17192), .ZN(n16959) );
  AOI211_X1 U20304 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17194), .A(n16960), .B(
        n16959), .ZN(n16961) );
  OAI211_X1 U20305 ( .C1(n16963), .C2(n19085), .A(n16962), .B(n16961), .ZN(
        P3_U2651) );
  NOR2_X1 U20306 ( .A1(n17181), .A2(n16976), .ZN(n16992) );
  NOR2_X1 U20307 ( .A1(n17181), .A2(n17155), .ZN(n17123) );
  AOI21_X1 U20308 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16992), .A(n17123), 
        .ZN(n16984) );
  INV_X1 U20309 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16969) );
  INV_X1 U20310 ( .A(n16988), .ZN(n17911) );
  NAND2_X1 U20311 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17911), .ZN(
        n16977) );
  AOI21_X1 U20312 ( .B1(n16969), .B2(n16977), .A(n17874), .ZN(n16964) );
  INV_X1 U20313 ( .A(n16964), .ZN(n17916) );
  INV_X1 U20314 ( .A(n17005), .ZN(n16965) );
  OAI21_X1 U20315 ( .B1(n16977), .B2(n16965), .A(n9924), .ZN(n16980) );
  OAI21_X1 U20316 ( .B1(n17916), .B2(n16980), .A(n17173), .ZN(n16966) );
  AOI21_X1 U20317 ( .B1(n17916), .B2(n16980), .A(n16966), .ZN(n16971) );
  OAI211_X1 U20318 ( .C1(n16987), .C2(n16975), .A(n17193), .B(n16967), .ZN(
        n16968) );
  OAI211_X1 U20319 ( .C1(n16969), .C2(n17159), .A(n18375), .B(n16968), .ZN(
        n16970) );
  AOI211_X1 U20320 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n16984), .A(n16971), 
        .B(n16970), .ZN(n16974) );
  INV_X1 U20321 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19084) );
  NAND3_X1 U20322 ( .A1(n17155), .A2(n16972), .A3(n19084), .ZN(n16973) );
  OAI211_X1 U20323 ( .C1(n16975), .C2(n17136), .A(n16974), .B(n16973), .ZN(
        P3_U2652) );
  OAI21_X1 U20324 ( .B1(n16993), .B2(n17341), .A(n17193), .ZN(n16986) );
  OAI21_X1 U20325 ( .B1(n17187), .B2(n16976), .A(n19081), .ZN(n16983) );
  OAI21_X1 U20326 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17911), .A(
        n16977), .ZN(n17922) );
  OAI221_X1 U20327 ( .B1(n17922), .B2(n17911), .C1(n17922), .C2(n17005), .A(
        n17173), .ZN(n16978) );
  AOI22_X1 U20328 ( .A1(n17922), .A2(n16980), .B1(n16979), .B2(n16978), .ZN(
        n16982) );
  INV_X1 U20329 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17925) );
  OAI22_X1 U20330 ( .A1(n17925), .A2(n17159), .B1(n17136), .B2(n17341), .ZN(
        n16981) );
  AOI211_X1 U20331 ( .C1(n16984), .C2(n16983), .A(n16982), .B(n16981), .ZN(
        n16985) );
  OAI211_X1 U20332 ( .C1(n16987), .C2(n16986), .A(n16985), .B(n18375), .ZN(
        P3_U2653) );
  AND2_X1 U20333 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9797), .ZN(
        n17004) );
  OAI21_X1 U20334 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n17004), .A(
        n16988), .ZN(n17931) );
  AOI21_X1 U20335 ( .B1(n9797), .B2(n16989), .A(n17182), .ZN(n16990) );
  XOR2_X1 U20336 ( .A(n17931), .B(n16990), .Z(n17000) );
  AOI22_X1 U20337 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17183), .B1(
        n17194), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16999) );
  NAND2_X1 U20338 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n17008) );
  NOR2_X1 U20339 ( .A1(n17187), .A2(n16991), .ZN(n17029) );
  NAND2_X1 U20340 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n17029), .ZN(n17026) );
  NOR3_X1 U20341 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n17008), .A3(n17026), 
        .ZN(n16997) );
  INV_X1 U20342 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19079) );
  NOR3_X1 U20343 ( .A1(n17123), .A2(n16992), .A3(n19079), .ZN(n16996) );
  AOI211_X1 U20344 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n16994), .A(n16993), .B(
        n17192), .ZN(n16995) );
  NOR4_X1 U20345 ( .A1(n18369), .A2(n16997), .A3(n16996), .A4(n16995), .ZN(
        n16998) );
  OAI211_X1 U20346 ( .C1(n19028), .C2(n17000), .A(n16999), .B(n16998), .ZN(
        P3_U2654) );
  INV_X1 U20347 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17014) );
  AOI211_X1 U20348 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17019), .A(n17001), .B(
        n17192), .ZN(n17002) );
  AOI211_X1 U20349 ( .C1(n17194), .C2(P3_EBX_REG_16__SCAN_IN), .A(n18435), .B(
        n17002), .ZN(n17013) );
  OAI21_X1 U20350 ( .B1(n17003), .B2(n17187), .A(n17196), .ZN(n17028) );
  AOI21_X1 U20351 ( .B1(n17014), .B2(n17015), .A(n17004), .ZN(n17007) );
  NOR2_X1 U20352 ( .A1(n17005), .A2(n17182), .ZN(n17018) );
  INV_X1 U20353 ( .A(n17007), .ZN(n17950) );
  INV_X1 U20354 ( .A(n17018), .ZN(n17006) );
  AOI221_X1 U20355 ( .B1(n17007), .B2(n17018), .C1(n17950), .C2(n17006), .A(
        n19028), .ZN(n17011) );
  INV_X1 U20356 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19077) );
  INV_X1 U20357 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19075) );
  INV_X1 U20358 ( .A(n17008), .ZN(n17009) );
  AOI211_X1 U20359 ( .C1(n19077), .C2(n19075), .A(n17009), .B(n17026), .ZN(
        n17010) );
  AOI211_X1 U20360 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(n17028), .A(n17011), 
        .B(n17010), .ZN(n17012) );
  OAI211_X1 U20361 ( .C1(n17014), .C2(n17159), .A(n17013), .B(n17012), .ZN(
        P3_U2655) );
  NOR2_X1 U20362 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19028), .ZN(
        n17126) );
  NOR2_X1 U20363 ( .A1(n17125), .A2(n17126), .ZN(n17186) );
  OAI21_X1 U20364 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17944), .A(
        n17015), .ZN(n17959) );
  AOI211_X1 U20365 ( .C1(n9924), .C2(n17016), .A(n17186), .B(n17959), .ZN(
        n17017) );
  AOI21_X1 U20366 ( .B1(n17183), .B2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n17017), .ZN(n17025) );
  NAND3_X1 U20367 ( .A1(n17173), .A2(n17018), .A3(n17959), .ZN(n17021) );
  OAI211_X1 U20368 ( .C1(n17027), .C2(n17022), .A(n17193), .B(n17019), .ZN(
        n17020) );
  OAI211_X1 U20369 ( .C1(n17022), .C2(n17136), .A(n17021), .B(n17020), .ZN(
        n17023) );
  AOI211_X1 U20370 ( .C1(P3_REIP_REG_15__SCAN_IN), .C2(n17028), .A(n18435), 
        .B(n17023), .ZN(n17024) );
  OAI211_X1 U20371 ( .C1(P3_REIP_REG_15__SCAN_IN), .C2(n17026), .A(n17025), 
        .B(n17024), .ZN(P3_U2656) );
  NAND2_X1 U20372 ( .A1(n17984), .A2(n17062), .ZN(n17036) );
  OAI21_X1 U20373 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17036), .A(
        n9924), .ZN(n17037) );
  INV_X1 U20374 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17031) );
  AOI21_X1 U20375 ( .B1(n17031), .B2(n17036), .A(n17944), .ZN(n17977) );
  XOR2_X1 U20376 ( .A(n17037), .B(n17977), .Z(n17035) );
  AOI211_X1 U20377 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17046), .A(n17027), .B(
        n17192), .ZN(n17033) );
  OAI21_X1 U20378 ( .B1(P3_REIP_REG_14__SCAN_IN), .B2(n17029), .A(n17028), 
        .ZN(n17030) );
  OAI211_X1 U20379 ( .C1(n17031), .C2(n17159), .A(n18375), .B(n17030), .ZN(
        n17032) );
  AOI211_X1 U20380 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17194), .A(n17033), .B(
        n17032), .ZN(n17034) );
  OAI21_X1 U20381 ( .B1(n17035), .B2(n19028), .A(n17034), .ZN(P3_U2657) );
  INV_X1 U20382 ( .A(n17062), .ZN(n17988) );
  NOR2_X1 U20383 ( .A1(n18000), .A2(n17988), .ZN(n17051) );
  OAI21_X1 U20384 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17051), .A(
        n17036), .ZN(n17989) );
  INV_X1 U20385 ( .A(n17989), .ZN(n17038) );
  NOR3_X1 U20386 ( .A1(n17038), .A2(n19028), .A3(n17037), .ZN(n17042) );
  INV_X1 U20387 ( .A(n17051), .ZN(n17039) );
  AOI211_X1 U20388 ( .C1(n9924), .C2(n17039), .A(n17186), .B(n17989), .ZN(
        n17041) );
  OAI22_X1 U20389 ( .A1(n17991), .A2(n17159), .B1(n17136), .B2(n17389), .ZN(
        n17040) );
  NOR4_X1 U20390 ( .A1(n18369), .A2(n17042), .A3(n17041), .A4(n17040), .ZN(
        n17050) );
  NAND2_X1 U20391 ( .A1(n17043), .A2(n17196), .ZN(n17078) );
  INV_X1 U20392 ( .A(n17078), .ZN(n17122) );
  AOI21_X1 U20393 ( .B1(n17044), .B2(n17122), .A(n17123), .ZN(n17068) );
  NOR2_X1 U20394 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17187), .ZN(n17055) );
  OAI21_X1 U20395 ( .B1(n17068), .B2(n17055), .A(P3_REIP_REG_13__SCAN_IN), 
        .ZN(n17049) );
  INV_X1 U20396 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19071) );
  NAND3_X1 U20397 ( .A1(n17155), .A2(n17045), .A3(n19071), .ZN(n17048) );
  OAI211_X1 U20398 ( .C1(n17053), .C2(n17389), .A(n17193), .B(n17046), .ZN(
        n17047) );
  NAND4_X1 U20399 ( .A1(n17050), .A2(n17049), .A3(n17048), .A4(n17047), .ZN(
        P3_U2658) );
  AOI21_X1 U20400 ( .B1(n18000), .B2(n17988), .A(n17051), .ZN(n18003) );
  AOI21_X1 U20401 ( .B1(n17062), .B2(n17110), .A(n17182), .ZN(n17052) );
  XNOR2_X1 U20402 ( .A(n18003), .B(n17052), .ZN(n17061) );
  AOI211_X1 U20403 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17070), .A(n17053), .B(
        n17192), .ZN(n17054) );
  AOI21_X1 U20404 ( .B1(n17183), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n17054), .ZN(n17060) );
  INV_X1 U20405 ( .A(n17055), .ZN(n17056) );
  OAI22_X1 U20406 ( .A1(n17136), .A2(n17426), .B1(n17057), .B2(n17056), .ZN(
        n17058) );
  AOI211_X1 U20407 ( .C1(P3_REIP_REG_12__SCAN_IN), .C2(n17068), .A(n18435), 
        .B(n17058), .ZN(n17059) );
  OAI211_X1 U20408 ( .C1(n19028), .C2(n17061), .A(n17060), .B(n17059), .ZN(
        P3_U2659) );
  AOI22_X1 U20409 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n17183), .B1(
        n17194), .B2(P3_EBX_REG_11__SCAN_IN), .ZN(n17074) );
  INV_X1 U20410 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17063) );
  INV_X1 U20411 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17090) );
  NOR2_X1 U20412 ( .A1(n18065), .A2(n17127), .ZN(n17109) );
  NAND2_X1 U20413 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17109), .ZN(
        n17099) );
  NOR2_X1 U20414 ( .A1(n17090), .A2(n17099), .ZN(n17089) );
  NAND2_X1 U20415 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17089), .ZN(
        n17080) );
  AOI21_X1 U20416 ( .B1(n17063), .B2(n17080), .A(n17062), .ZN(n18016) );
  OAI21_X1 U20417 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17080), .A(
        n9924), .ZN(n17064) );
  XNOR2_X1 U20418 ( .A(n18016), .B(n17064), .ZN(n17069) );
  NOR2_X1 U20419 ( .A1(n17187), .A2(n17065), .ZN(n17141) );
  NAND2_X1 U20420 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n17141), .ZN(n17124) );
  OAI21_X1 U20421 ( .B1(n17066), .B2(n17124), .A(n19067), .ZN(n17067) );
  AOI22_X1 U20422 ( .A1(n17173), .A2(n17069), .B1(n17068), .B2(n17067), .ZN(
        n17073) );
  OAI211_X1 U20423 ( .C1(n17075), .C2(n17071), .A(n17193), .B(n17070), .ZN(
        n17072) );
  NAND4_X1 U20424 ( .A1(n17074), .A2(n17073), .A3(n18375), .A4(n17072), .ZN(
        P3_U2660) );
  INV_X1 U20425 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18012) );
  AOI211_X1 U20426 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17076), .A(n17075), .B(
        n17192), .ZN(n17077) );
  AOI211_X1 U20427 ( .C1(n17194), .C2(P3_EBX_REG_10__SCAN_IN), .A(n18435), .B(
        n17077), .ZN(n17086) );
  INV_X1 U20428 ( .A(n17123), .ZN(n17195) );
  OAI21_X1 U20429 ( .B1(n17079), .B2(n17078), .A(n17195), .ZN(n17108) );
  INV_X1 U20430 ( .A(n17108), .ZN(n17096) );
  NOR3_X1 U20431 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n17079), .A3(n17124), .ZN(
        n17087) );
  AOI21_X1 U20432 ( .B1(n17089), .B2(n17110), .A(n17182), .ZN(n17091) );
  OAI21_X1 U20433 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17089), .A(
        n17080), .ZN(n18032) );
  XOR2_X1 U20434 ( .A(n17091), .B(n18032), .Z(n17083) );
  INV_X1 U20435 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19065) );
  NAND2_X1 U20436 ( .A1(n17081), .A2(n19065), .ZN(n17082) );
  OAI22_X1 U20437 ( .A1(n19028), .A2(n17083), .B1(n17124), .B2(n17082), .ZN(
        n17084) );
  AOI221_X1 U20438 ( .B1(n17096), .B2(P3_REIP_REG_10__SCAN_IN), .C1(n17087), 
        .C2(P3_REIP_REG_10__SCAN_IN), .A(n17084), .ZN(n17085) );
  OAI211_X1 U20439 ( .C1(n18012), .C2(n17159), .A(n17086), .B(n17085), .ZN(
        P3_U2661) );
  AOI211_X1 U20440 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n17183), .A(
        n18408), .B(n17087), .ZN(n17098) );
  OR2_X1 U20441 ( .A1(n17192), .A2(n17088), .ZN(n17103) );
  AOI21_X1 U20442 ( .B1(n17193), .B2(n17088), .A(n17194), .ZN(n17094) );
  AOI21_X1 U20443 ( .B1(n17090), .B2(n17099), .A(n17089), .ZN(n18036) );
  AOI221_X1 U20444 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18036), .C1(
        n17099), .C2(n18036), .A(n19028), .ZN(n17092) );
  OAI22_X1 U20445 ( .A1(n17125), .A2(n17092), .B1(n18036), .B2(n17091), .ZN(
        n17093) );
  OAI221_X1 U20446 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17103), .C1(n17442), 
        .C2(n17094), .A(n17093), .ZN(n17095) );
  AOI21_X1 U20447 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n17096), .A(n17095), .ZN(
        n17097) );
  NAND2_X1 U20448 ( .A1(n17098), .A2(n17097), .ZN(P3_U2662) );
  INV_X1 U20449 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19061) );
  OAI21_X1 U20450 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17109), .A(
        n17099), .ZN(n18050) );
  OR2_X1 U20451 ( .A1(n18047), .A2(n18065), .ZN(n18046) );
  OAI21_X1 U20452 ( .B1(n18046), .B2(n17150), .A(n9924), .ZN(n17101) );
  OAI21_X1 U20453 ( .B1(n18050), .B2(n17101), .A(n17173), .ZN(n17100) );
  AOI21_X1 U20454 ( .B1(n18050), .B2(n17101), .A(n17100), .ZN(n17102) );
  AOI211_X1 U20455 ( .C1(n17194), .C2(P3_EBX_REG_8__SCAN_IN), .A(n18408), .B(
        n17102), .ZN(n17107) );
  INV_X1 U20456 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19059) );
  INV_X1 U20457 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19057) );
  NOR4_X1 U20458 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n19059), .A3(n19057), .A4(
        n17124), .ZN(n17105) );
  AOI21_X1 U20459 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17116), .A(n17103), .ZN(
        n17104) );
  AOI211_X1 U20460 ( .C1(n17183), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17105), .B(n17104), .ZN(n17106) );
  OAI211_X1 U20461 ( .C1(n19061), .C2(n17108), .A(n17107), .B(n17106), .ZN(
        P3_U2663) );
  AOI22_X1 U20462 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17183), .B1(
        n17194), .B2(P3_EBX_REG_7__SCAN_IN), .ZN(n17119) );
  NOR2_X1 U20463 ( .A1(n19057), .A2(n17124), .ZN(n17115) );
  OAI22_X1 U20464 ( .A1(n17123), .A2(n17122), .B1(P3_REIP_REG_6__SCAN_IN), 
        .B2(n17124), .ZN(n17114) );
  AOI21_X1 U20465 ( .B1(n18065), .B2(n17127), .A(n17109), .ZN(n18069) );
  INV_X1 U20466 ( .A(n17127), .ZN(n17111) );
  AOI21_X1 U20467 ( .B1(n17111), .B2(n17110), .A(n17182), .ZN(n17131) );
  OAI21_X1 U20468 ( .B1(n18069), .B2(n17131), .A(n17173), .ZN(n17112) );
  AOI21_X1 U20469 ( .B1(n18069), .B2(n17131), .A(n17112), .ZN(n17113) );
  AOI221_X1 U20470 ( .B1(n17115), .B2(n19059), .C1(n17114), .C2(
        P3_REIP_REG_7__SCAN_IN), .A(n17113), .ZN(n17118) );
  OAI211_X1 U20471 ( .C1(n17120), .C2(n17499), .A(n17193), .B(n17116), .ZN(
        n17117) );
  NAND4_X1 U20472 ( .A1(n17119), .A2(n17118), .A3(n18375), .A4(n17117), .ZN(
        P3_U2664) );
  AOI211_X1 U20473 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17142), .A(n17120), .B(
        n17192), .ZN(n17121) );
  AOI211_X1 U20474 ( .C1(n17194), .C2(P3_EBX_REG_6__SCAN_IN), .A(n18408), .B(
        n17121), .ZN(n17134) );
  NOR2_X1 U20475 ( .A1(n17123), .A2(n17122), .ZN(n17140) );
  INV_X1 U20476 ( .A(n17124), .ZN(n17130) );
  AOI21_X1 U20477 ( .B1(n17135), .B2(n17126), .A(n17125), .ZN(n17128) );
  OAI21_X1 U20478 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17135), .A(
        n17127), .ZN(n18084) );
  INV_X1 U20479 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18079) );
  OAI22_X1 U20480 ( .A1(n17128), .A2(n18084), .B1(n18079), .B2(n17159), .ZN(
        n17129) );
  AOI221_X1 U20481 ( .B1(n17140), .B2(P3_REIP_REG_6__SCAN_IN), .C1(n17130), 
        .C2(n19057), .A(n17129), .ZN(n17133) );
  NAND3_X1 U20482 ( .A1(n17173), .A2(n17131), .A3(n18084), .ZN(n17132) );
  NAND3_X1 U20483 ( .A1(n17134), .A2(n17133), .A3(n17132), .ZN(P3_U2665) );
  AOI21_X1 U20484 ( .B1(n17137), .B2(n17148), .A(n17135), .ZN(n18094) );
  OAI21_X1 U20485 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17148), .A(
        n9924), .ZN(n17147) );
  XNOR2_X1 U20486 ( .A(n18094), .B(n17147), .ZN(n17139) );
  OAI22_X1 U20487 ( .A1(n17137), .A2(n17159), .B1(n17136), .B2(n17143), .ZN(
        n17138) );
  AOI21_X1 U20488 ( .B1(n17173), .B2(n17139), .A(n17138), .ZN(n17146) );
  OAI21_X1 U20489 ( .B1(P3_REIP_REG_5__SCAN_IN), .B2(n17141), .A(n17140), .ZN(
        n17145) );
  OAI211_X1 U20490 ( .C1(n17153), .C2(n17143), .A(n17193), .B(n17142), .ZN(
        n17144) );
  NAND4_X1 U20491 ( .A1(n17146), .A2(n18375), .A3(n17145), .A4(n17144), .ZN(
        P3_U2666) );
  INV_X1 U20492 ( .A(n17147), .ZN(n17152) );
  NAND2_X1 U20493 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18106), .ZN(
        n17168) );
  INV_X1 U20494 ( .A(n17168), .ZN(n17149) );
  OAI21_X1 U20495 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17149), .A(
        n17148), .ZN(n18109) );
  INV_X1 U20496 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17158) );
  NAND2_X1 U20497 ( .A1(n18106), .A2(n17158), .ZN(n18100) );
  OAI22_X1 U20498 ( .A1(n9924), .A2(n18109), .B1(n17150), .B2(n18100), .ZN(
        n17151) );
  AOI21_X1 U20499 ( .B1(n17152), .B2(n18109), .A(n17151), .ZN(n17163) );
  AOI211_X1 U20500 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17174), .A(n17153), .B(
        n17192), .ZN(n17154) );
  AOI21_X1 U20501 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17194), .A(n17154), .ZN(
        n17162) );
  OAI21_X1 U20502 ( .B1(n17164), .B2(n17187), .A(n17196), .ZN(n17171) );
  INV_X1 U20503 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19053) );
  NAND3_X1 U20504 ( .A1(n17155), .A2(n17164), .A3(n19053), .ZN(n17157) );
  OAI21_X1 U20505 ( .B1(n17488), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n19188), .ZN(n17156) );
  OAI211_X1 U20506 ( .C1(n17159), .C2(n17158), .A(n17157), .B(n17156), .ZN(
        n17160) );
  AOI211_X1 U20507 ( .C1(P3_REIP_REG_4__SCAN_IN), .C2(n17171), .A(n18435), .B(
        n17160), .ZN(n17161) );
  OAI211_X1 U20508 ( .C1(n17163), .C2(n19028), .A(n17162), .B(n17161), .ZN(
        P3_U2667) );
  AOI22_X1 U20509 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n17183), .B1(
        n17194), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n17179) );
  NOR2_X1 U20510 ( .A1(n17164), .A2(n17187), .ZN(n17166) );
  OAI21_X1 U20511 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18970), .A(
        n17470), .ZN(n17165) );
  INV_X1 U20512 ( .A(n17165), .ZN(n19126) );
  AOI22_X1 U20513 ( .A1(n17167), .A2(n17166), .B1(n19188), .B2(n19126), .ZN(
        n17178) );
  NOR2_X1 U20514 ( .A1(n18143), .A2(n18133), .ZN(n17169) );
  OAI21_X1 U20515 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17169), .A(
        n17168), .ZN(n18123) );
  XNOR2_X1 U20516 ( .A(n17170), .B(n18123), .ZN(n17172) );
  AOI22_X1 U20517 ( .A1(n17173), .A2(n17172), .B1(P3_REIP_REG_3__SCAN_IN), 
        .B2(n17171), .ZN(n17177) );
  OAI211_X1 U20518 ( .C1(n17175), .C2(n17513), .A(n17193), .B(n17174), .ZN(
        n17176) );
  NAND4_X1 U20519 ( .A1(n17179), .A2(n17178), .A3(n17177), .A4(n17176), .ZN(
        P3_U2668) );
  OAI21_X1 U20520 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17521), .ZN(n17527) );
  NAND2_X1 U20521 ( .A1(n18974), .A2(n17180), .ZN(n18993) );
  INV_X1 U20522 ( .A(n18993), .ZN(n19143) );
  AOI22_X1 U20523 ( .A1(n17181), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n19143), 
        .B2(n19188), .ZN(n17191) );
  NOR2_X1 U20524 ( .A1(n17182), .A2(n19028), .ZN(n17184) );
  AOI211_X1 U20525 ( .C1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n17184), .A(
        n17183), .B(n18143), .ZN(n17185) );
  AOI21_X1 U20526 ( .B1(n17186), .B2(n18143), .A(n17185), .ZN(n17189) );
  NOR2_X1 U20527 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17187), .ZN(n17188) );
  AOI211_X1 U20528 ( .C1(P3_EBX_REG_1__SCAN_IN), .C2(n17194), .A(n17189), .B(
        n17188), .ZN(n17190) );
  OAI211_X1 U20529 ( .C1(n17192), .C2(n17527), .A(n17191), .B(n17190), .ZN(
        P3_U2670) );
  NOR2_X1 U20530 ( .A1(n17194), .A2(n17193), .ZN(n17200) );
  AOI22_X1 U20531 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n17195), .B1(n19188), 
        .B2(n12924), .ZN(n17199) );
  NAND3_X1 U20532 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17197), .A3(
        n17196), .ZN(n17198) );
  OAI211_X1 U20533 ( .C1(n17200), .C2(n17532), .A(n17199), .B(n17198), .ZN(
        P3_U2671) );
  NAND4_X1 U20534 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n17201)
         );
  NOR4_X1 U20535 ( .A1(n17242), .A2(n17203), .A3(n17202), .A4(n17201), .ZN(
        n17204) );
  NAND4_X1 U20536 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n17285), .A4(n17204), .ZN(n17207) );
  NOR2_X1 U20537 ( .A1(n17208), .A2(n17207), .ZN(n17234) );
  NAND2_X1 U20538 ( .A1(n17525), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17206) );
  NAND2_X1 U20539 ( .A1(n17234), .A2(n18533), .ZN(n17205) );
  OAI22_X1 U20540 ( .A1(n17234), .A2(n17206), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17205), .ZN(P3_U2672) );
  NAND2_X1 U20541 ( .A1(n17208), .A2(n17207), .ZN(n17209) );
  NAND2_X1 U20542 ( .A1(n17209), .A2(n17525), .ZN(n17233) );
  AOI22_X1 U20543 ( .A1(n17448), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17210) );
  OAI21_X1 U20544 ( .B1(n17373), .B2(n17402), .A(n17210), .ZN(n17220) );
  AOI22_X1 U20545 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17218) );
  INV_X1 U20546 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17211) );
  OAI22_X1 U20547 ( .A1(n12984), .A2(n18740), .B1(n9682), .B2(n17211), .ZN(
        n17216) );
  AOI22_X1 U20548 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17214) );
  AOI22_X1 U20549 ( .A1(n12970), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17213) );
  AOI22_X1 U20550 ( .A1(n17488), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17212) );
  NAND3_X1 U20551 ( .A1(n17214), .A2(n17213), .A3(n17212), .ZN(n17215) );
  AOI211_X1 U20552 ( .C1(n17393), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n17216), .B(n17215), .ZN(n17217) );
  OAI211_X1 U20553 ( .C1(n12951), .C2(n18528), .A(n17218), .B(n17217), .ZN(
        n17219) );
  AOI211_X1 U20554 ( .C1(n17431), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n17220), .B(n17219), .ZN(n17238) );
  NOR2_X1 U20555 ( .A1(n17238), .A2(n17237), .ZN(n17236) );
  AOI22_X1 U20556 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17231) );
  AOI22_X1 U20557 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U20558 ( .A1(n17431), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9685), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17221) );
  OAI211_X1 U20559 ( .C1(n12943), .C2(n17223), .A(n17222), .B(n17221), .ZN(
        n17229) );
  AOI22_X1 U20560 ( .A1(n17430), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17227) );
  AOI22_X1 U20561 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17226) );
  AOI22_X1 U20562 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17488), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17225) );
  NAND2_X1 U20563 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n17224) );
  NAND4_X1 U20564 ( .A1(n17227), .A2(n17226), .A3(n17225), .A4(n17224), .ZN(
        n17228) );
  AOI211_X1 U20565 ( .C1(n17490), .C2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n17229), .B(n17228), .ZN(n17230) );
  OAI211_X1 U20566 ( .C1(n17429), .C2(n18825), .A(n17231), .B(n17230), .ZN(
        n17232) );
  XNOR2_X1 U20567 ( .A(n17236), .B(n17232), .ZN(n17543) );
  OAI22_X1 U20568 ( .A1(n17234), .A2(n17233), .B1(n17543), .B2(n17525), .ZN(
        P3_U2673) );
  INV_X1 U20569 ( .A(n17235), .ZN(n17241) );
  AOI21_X1 U20570 ( .B1(n17238), .B2(n17237), .A(n17236), .ZN(n17544) );
  AOI22_X1 U20571 ( .A1(n17530), .A2(n17544), .B1(n17239), .B2(n17242), .ZN(
        n17240) );
  OAI21_X1 U20572 ( .B1(n17242), .B2(n17241), .A(n17240), .ZN(P3_U2674) );
  INV_X1 U20573 ( .A(n17243), .ZN(n17252) );
  AOI21_X1 U20574 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17525), .A(n17252), .ZN(
        n17247) );
  AOI21_X1 U20575 ( .B1(n17245), .B2(n17249), .A(n17244), .ZN(n17553) );
  INV_X1 U20576 ( .A(n17553), .ZN(n17246) );
  OAI22_X1 U20577 ( .A1(n17248), .A2(n17247), .B1(n17246), .B2(n17525), .ZN(
        P3_U2676) );
  AOI21_X1 U20578 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17525), .A(n17258), .ZN(
        n17251) );
  OAI21_X1 U20579 ( .B1(n17254), .B2(n17250), .A(n17249), .ZN(n17561) );
  OAI22_X1 U20580 ( .A1(n17252), .A2(n17251), .B1(n17561), .B2(n17525), .ZN(
        P3_U2677) );
  INV_X1 U20581 ( .A(n17253), .ZN(n17262) );
  AOI21_X1 U20582 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17525), .A(n17262), .ZN(
        n17257) );
  AOI21_X1 U20583 ( .B1(n17255), .B2(n17259), .A(n17254), .ZN(n17562) );
  INV_X1 U20584 ( .A(n17562), .ZN(n17256) );
  OAI22_X1 U20585 ( .A1(n17258), .A2(n17257), .B1(n17256), .B2(n17525), .ZN(
        P3_U2678) );
  AOI21_X1 U20586 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17525), .A(n17269), .ZN(
        n17261) );
  OAI21_X1 U20587 ( .B1(n17264), .B2(n17260), .A(n17259), .ZN(n17571) );
  OAI22_X1 U20588 ( .A1(n17262), .A2(n17261), .B1(n17571), .B2(n17525), .ZN(
        P3_U2679) );
  INV_X1 U20589 ( .A(n17263), .ZN(n17284) );
  AOI21_X1 U20590 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17525), .A(n17284), .ZN(
        n17268) );
  AOI21_X1 U20591 ( .B1(n17266), .B2(n17265), .A(n17264), .ZN(n17572) );
  INV_X1 U20592 ( .A(n17572), .ZN(n17267) );
  OAI22_X1 U20593 ( .A1(n17269), .A2(n17268), .B1(n17525), .B2(n17267), .ZN(
        P3_U2680) );
  AOI21_X1 U20594 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17525), .A(n17270), .ZN(
        n17283) );
  AOI22_X1 U20595 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17281) );
  INV_X1 U20596 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17273) );
  AOI22_X1 U20597 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12970), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17272) );
  AOI22_X1 U20598 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17271) );
  OAI211_X1 U20599 ( .C1(n17470), .C2(n17273), .A(n17272), .B(n17271), .ZN(
        n17279) );
  AOI22_X1 U20600 ( .A1(n17467), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17277) );
  AOI22_X1 U20601 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17276) );
  AOI22_X1 U20602 ( .A1(n9685), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17275) );
  NAND2_X1 U20603 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n17274) );
  NAND4_X1 U20604 ( .A1(n17277), .A2(n17276), .A3(n17275), .A4(n17274), .ZN(
        n17278) );
  AOI211_X1 U20605 ( .C1(n17490), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n17279), .B(n17278), .ZN(n17280) );
  OAI211_X1 U20606 ( .C1(n17485), .C2(n18528), .A(n17281), .B(n17280), .ZN(
        n17577) );
  INV_X1 U20607 ( .A(n17577), .ZN(n17282) );
  OAI22_X1 U20608 ( .A1(n17284), .A2(n17283), .B1(n17282), .B2(n17525), .ZN(
        P3_U2681) );
  NOR2_X1 U20609 ( .A1(n17530), .A2(n17285), .ZN(n17310) );
  AOI22_X1 U20610 ( .A1(n17490), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17488), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17296) );
  AOI22_X1 U20611 ( .A1(n12970), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17287) );
  AOI22_X1 U20612 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17286) );
  OAI211_X1 U20613 ( .C1(n12943), .C2(n9878), .A(n17287), .B(n17286), .ZN(
        n17294) );
  AOI22_X1 U20614 ( .A1(n9685), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9704), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17292) );
  AOI22_X1 U20615 ( .A1(n17431), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17291) );
  AOI22_X1 U20616 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17288), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17290) );
  NAND2_X1 U20617 ( .A1(n12952), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n17289) );
  NAND4_X1 U20618 ( .A1(n17292), .A2(n17291), .A3(n17290), .A4(n17289), .ZN(
        n17293) );
  AOI211_X1 U20619 ( .C1(n17393), .C2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n17294), .B(n17293), .ZN(n17295) );
  OAI211_X1 U20620 ( .C1(n17485), .C2(n18523), .A(n17296), .B(n17295), .ZN(
        n17584) );
  AOI22_X1 U20621 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17310), .B1(n17530), 
        .B2(n17584), .ZN(n17297) );
  OAI21_X1 U20622 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17298), .A(n17297), .ZN(
        P3_U2682) );
  AOI22_X1 U20623 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17309) );
  AOI22_X1 U20624 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17299) );
  OAI21_X1 U20625 ( .B1(n12977), .B2(n18733), .A(n17299), .ZN(n17307) );
  OAI22_X1 U20626 ( .A1(n12984), .A2(n17418), .B1(n17470), .B2(n17300), .ZN(
        n17301) );
  AOI21_X1 U20627 ( .B1(n17490), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n17301), .ZN(n17305) );
  AOI22_X1 U20628 ( .A1(n17430), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17304) );
  AOI22_X1 U20629 ( .A1(n9685), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17303) );
  AOI22_X1 U20630 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17302) );
  NAND4_X1 U20631 ( .A1(n17305), .A2(n17304), .A3(n17303), .A4(n17302), .ZN(
        n17306) );
  AOI211_X1 U20632 ( .C1(n15895), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n17307), .B(n17306), .ZN(n17308) );
  OAI211_X1 U20633 ( .C1(n17485), .C2(n18517), .A(n17309), .B(n17308), .ZN(
        n17588) );
  INV_X1 U20634 ( .A(n17588), .ZN(n17313) );
  OAI21_X1 U20635 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17311), .A(n17310), .ZN(
        n17312) );
  OAI21_X1 U20636 ( .B1(n17313), .B2(n17525), .A(n17312), .ZN(P3_U2683) );
  AOI22_X1 U20637 ( .A1(n9688), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17314) );
  OAI21_X1 U20638 ( .B1(n12977), .B2(n17315), .A(n17314), .ZN(n17325) );
  AOI22_X1 U20639 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17323) );
  OAI22_X1 U20640 ( .A1(n9682), .A2(n17316), .B1(n12943), .B2(n18812), .ZN(
        n17321) );
  AOI22_X1 U20641 ( .A1(n17430), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17319) );
  AOI22_X1 U20642 ( .A1(n9685), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17318) );
  AOI22_X1 U20643 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17488), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17317) );
  NAND3_X1 U20644 ( .A1(n17319), .A2(n17318), .A3(n17317), .ZN(n17320) );
  AOI211_X1 U20645 ( .C1(n17288), .C2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n17321), .B(n17320), .ZN(n17322) );
  OAI211_X1 U20646 ( .C1(n17485), .C2(n18512), .A(n17323), .B(n17322), .ZN(
        n17324) );
  AOI211_X1 U20647 ( .C1(n15895), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n17325), .B(n17324), .ZN(n17599) );
  OAI21_X1 U20648 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17328), .A(n17326), .ZN(
        n17327) );
  AOI22_X1 U20649 ( .A1(n17530), .A2(n17599), .B1(n17327), .B2(n17525), .ZN(
        P3_U2684) );
  OR2_X1 U20650 ( .A1(n17341), .A2(n17328), .ZN(n17343) );
  AOI22_X1 U20651 ( .A1(n9685), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17329) );
  OAI21_X1 U20652 ( .B1(n17429), .B2(n17447), .A(n17329), .ZN(n17339) );
  AOI22_X1 U20653 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17336) );
  AOI22_X1 U20654 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17488), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17330) );
  OAI21_X1 U20655 ( .B1(n12943), .B2(n18809), .A(n17330), .ZN(n17334) );
  AOI22_X1 U20656 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17332) );
  AOI22_X1 U20657 ( .A1(n17431), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12952), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17331) );
  OAI211_X1 U20658 ( .C1(n17486), .C2(n17452), .A(n17332), .B(n17331), .ZN(
        n17333) );
  AOI211_X1 U20659 ( .C1(n17490), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n17334), .B(n17333), .ZN(n17335) );
  OAI211_X1 U20660 ( .C1(n12959), .C2(n17337), .A(n17336), .B(n17335), .ZN(
        n17338) );
  AOI211_X1 U20661 ( .C1(n15895), .C2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n17339), .B(n17338), .ZN(n17604) );
  NOR2_X1 U20662 ( .A1(n17340), .A2(n17528), .ZN(n17370) );
  NAND3_X1 U20663 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17370), .A3(n17341), 
        .ZN(n17342) );
  OAI221_X1 U20664 ( .B1(n17530), .B2(n17343), .C1(n17525), .C2(n17604), .A(
        n17342), .ZN(P3_U2685) );
  INV_X1 U20665 ( .A(n17370), .ZN(n17356) );
  OAI22_X1 U20666 ( .A1(n17344), .A2(n12984), .B1(n12959), .B2(n17464), .ZN(
        n17354) );
  AOI22_X1 U20667 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9685), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17352) );
  AOI22_X1 U20668 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n15828), .B1(
        n17431), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17351) );
  OAI22_X1 U20669 ( .A1(n18806), .A2(n12943), .B1(n18501), .B2(n17485), .ZN(
        n17349) );
  AOI22_X1 U20670 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n12952), .ZN(n17347) );
  AOI22_X1 U20671 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17430), .B1(
        n12970), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17346) );
  AOI22_X1 U20672 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17488), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17345) );
  NAND3_X1 U20673 ( .A1(n17347), .A2(n17346), .A3(n17345), .ZN(n17348) );
  AOI211_X1 U20674 ( .C1(n17490), .C2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n17349), .B(n17348), .ZN(n17350) );
  NAND3_X1 U20675 ( .A1(n17352), .A2(n17351), .A3(n17350), .ZN(n17353) );
  AOI211_X1 U20676 ( .C1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .C2(n15894), .A(
        n17354), .B(n17353), .ZN(n17609) );
  NAND3_X1 U20677 ( .A1(n17356), .A2(P3_EBX_REG_17__SCAN_IN), .A3(n17525), 
        .ZN(n17355) );
  OAI221_X1 U20678 ( .B1(n17356), .B2(P3_EBX_REG_17__SCAN_IN), .C1(n17525), 
        .C2(n17609), .A(n17355), .ZN(P3_U2686) );
  OAI22_X1 U20679 ( .A1(n9756), .A2(n17357), .B1(n12984), .B2(n17484), .ZN(
        n17367) );
  AOI22_X1 U20680 ( .A1(n9704), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17365) );
  AOI22_X1 U20681 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17364) );
  OAI22_X1 U20682 ( .A1(n17485), .A2(n18496), .B1(n12943), .B2(n18802), .ZN(
        n17362) );
  AOI22_X1 U20683 ( .A1(n17431), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9685), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17360) );
  AOI22_X1 U20684 ( .A1(n17430), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12952), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17359) );
  AOI22_X1 U20685 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17358) );
  NAND3_X1 U20686 ( .A1(n17360), .A2(n17359), .A3(n17358), .ZN(n17361) );
  AOI211_X1 U20687 ( .C1(n17488), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n17362), .B(n17361), .ZN(n17363) );
  NAND3_X1 U20688 ( .A1(n17365), .A2(n17364), .A3(n17363), .ZN(n17366) );
  AOI211_X1 U20689 ( .C1(n17449), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n17367), .B(n17366), .ZN(n17615) );
  NOR2_X1 U20690 ( .A1(n17578), .A2(n17385), .ZN(n17403) );
  AND2_X1 U20691 ( .A1(n17368), .A2(n17403), .ZN(n17388) );
  AOI21_X1 U20692 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17525), .A(n17388), .ZN(
        n17369) );
  OAI22_X1 U20693 ( .A1(n17615), .A2(n17525), .B1(n17370), .B2(n17369), .ZN(
        P3_U2687) );
  AOI22_X1 U20694 ( .A1(n15828), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17371) );
  OAI21_X1 U20695 ( .B1(n17373), .B2(n17372), .A(n17371), .ZN(n17384) );
  AOI22_X1 U20696 ( .A1(n17431), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17381) );
  OAI22_X1 U20697 ( .A1(n17486), .A2(n18537), .B1(n17485), .B2(n17374), .ZN(
        n17379) );
  AOI22_X1 U20698 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9688), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17377) );
  AOI22_X1 U20699 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12970), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17376) );
  AOI22_X1 U20700 ( .A1(n17490), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17488), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17375) );
  NAND3_X1 U20701 ( .A1(n17377), .A2(n17376), .A3(n17375), .ZN(n17378) );
  AOI211_X1 U20702 ( .C1(n17489), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n17379), .B(n17378), .ZN(n17380) );
  OAI211_X1 U20703 ( .C1(n12984), .C2(n17382), .A(n17381), .B(n17380), .ZN(
        n17383) );
  AOI211_X1 U20704 ( .C1(n9685), .C2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n17384), .B(n17383), .ZN(n17619) );
  NOR3_X1 U20705 ( .A1(n17408), .A2(n17389), .A3(n17385), .ZN(n17386) );
  OAI21_X1 U20706 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17386), .A(n17525), .ZN(
        n17387) );
  OAI22_X1 U20707 ( .A1(n17619), .A2(n17525), .B1(n17388), .B2(n17387), .ZN(
        P3_U2688) );
  NOR2_X1 U20708 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17389), .ZN(n17404) );
  AOI22_X1 U20709 ( .A1(n9685), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9704), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17401) );
  INV_X1 U20710 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17392) );
  AOI22_X1 U20711 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17448), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17391) );
  AOI22_X1 U20712 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17431), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17390) );
  OAI211_X1 U20713 ( .C1(n17470), .C2(n17392), .A(n17391), .B(n17390), .ZN(
        n17399) );
  AOI22_X1 U20714 ( .A1(n15828), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17397) );
  AOI22_X1 U20715 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12952), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17396) );
  AOI22_X1 U20716 ( .A1(n17393), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17395) );
  NAND2_X1 U20717 ( .A1(n17489), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n17394) );
  NAND4_X1 U20718 ( .A1(n17397), .A2(n17396), .A3(n17395), .A4(n17394), .ZN(
        n17398) );
  AOI211_X1 U20719 ( .C1(n17490), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n17399), .B(n17398), .ZN(n17400) );
  OAI211_X1 U20720 ( .C1(n12984), .C2(n17402), .A(n17401), .B(n17400), .ZN(
        n17622) );
  AOI22_X1 U20721 ( .A1(n17404), .A2(n17403), .B1(n17530), .B2(n17622), .ZN(
        n17405) );
  OAI221_X1 U20722 ( .B1(n17408), .B2(n17407), .C1(n17408), .C2(n17406), .A(
        n17405), .ZN(P3_U2689) );
  AOI221_X1 U20723 ( .B1(n17421), .B2(n18533), .C1(n17422), .C2(n18533), .A(
        n17520), .ZN(n17443) );
  AOI22_X1 U20724 ( .A1(n9685), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17409) );
  OAI21_X1 U20725 ( .B1(n9756), .B2(n18733), .A(n17409), .ZN(n17420) );
  AOI22_X1 U20726 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17417) );
  AOI22_X1 U20727 ( .A1(n17490), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17410) );
  OAI21_X1 U20728 ( .B1(n17486), .B2(n18517), .A(n17410), .ZN(n17415) );
  AOI22_X1 U20729 ( .A1(n9688), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17448), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17412) );
  AOI22_X1 U20730 ( .A1(n17430), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12952), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17411) );
  OAI211_X1 U20731 ( .C1(n17470), .C2(n17413), .A(n17412), .B(n17411), .ZN(
        n17414) );
  AOI211_X1 U20732 ( .C1(n17489), .C2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A(
        n17415), .B(n17414), .ZN(n17416) );
  OAI211_X1 U20733 ( .C1(n12977), .C2(n17418), .A(n17417), .B(n17416), .ZN(
        n17419) );
  AOI211_X1 U20734 ( .C1(n9689), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n17420), .B(n17419), .ZN(n17632) );
  INV_X1 U20735 ( .A(n17632), .ZN(n17424) );
  NOR2_X1 U20736 ( .A1(n17520), .A2(n17421), .ZN(n17509) );
  NAND2_X1 U20737 ( .A1(n18533), .A2(n17509), .ZN(n17514) );
  NOR2_X1 U20738 ( .A1(n17422), .A2(n17514), .ZN(n17423) );
  AOI22_X1 U20739 ( .A1(n17530), .A2(n17424), .B1(n17423), .B2(n17426), .ZN(
        n17425) );
  OAI21_X1 U20740 ( .B1(n17426), .B2(n17443), .A(n17425), .ZN(P3_U2691) );
  AOI22_X1 U20741 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17427) );
  OAI21_X1 U20742 ( .B1(n17429), .B2(n17428), .A(n17427), .ZN(n17440) );
  AOI22_X1 U20743 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17438) );
  OAI22_X1 U20744 ( .A1(n17486), .A2(n18512), .B1(n17485), .B2(n18919), .ZN(
        n17436) );
  AOI22_X1 U20745 ( .A1(n17430), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17434) );
  AOI22_X1 U20746 ( .A1(n17431), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9685), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17433) );
  AOI22_X1 U20747 ( .A1(n17490), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17488), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17432) );
  NAND3_X1 U20748 ( .A1(n17434), .A2(n17433), .A3(n17432), .ZN(n17435) );
  AOI211_X1 U20749 ( .C1(n17489), .C2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n17436), .B(n17435), .ZN(n17437) );
  OAI211_X1 U20750 ( .C1(n12959), .C2(n18812), .A(n17438), .B(n17437), .ZN(
        n17439) );
  AOI211_X1 U20751 ( .C1(n15895), .C2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A(
        n17440), .B(n17439), .ZN(n17636) );
  NAND2_X1 U20752 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17509), .ZN(n17505) );
  NOR2_X1 U20753 ( .A1(n17441), .A2(n17505), .ZN(n17480) );
  INV_X1 U20754 ( .A(n17480), .ZN(n17500) );
  NOR2_X1 U20755 ( .A1(n17442), .A2(n17500), .ZN(n17461) );
  AOI21_X1 U20756 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17461), .A(
        P3_EBX_REG_11__SCAN_IN), .ZN(n17444) );
  OAI22_X1 U20757 ( .A1(n17636), .A2(n17525), .B1(n17444), .B2(n17443), .ZN(
        P3_U2692) );
  AOI22_X1 U20758 ( .A1(n9685), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17430), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17445) );
  OAI21_X1 U20759 ( .B1(n12959), .B2(n18809), .A(n17445), .ZN(n17459) );
  INV_X1 U20760 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17457) );
  AOI22_X1 U20761 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17456) );
  AOI22_X1 U20762 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17446) );
  OAI21_X1 U20763 ( .B1(n12943), .B2(n17447), .A(n17446), .ZN(n17454) );
  AOI22_X1 U20764 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17448), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17451) );
  AOI22_X1 U20765 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17450) );
  OAI211_X1 U20766 ( .C1(n17470), .C2(n17452), .A(n17451), .B(n17450), .ZN(
        n17453) );
  AOI211_X1 U20767 ( .C1(n17393), .C2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n17454), .B(n17453), .ZN(n17455) );
  OAI211_X1 U20768 ( .C1(n12977), .C2(n17457), .A(n17456), .B(n17455), .ZN(
        n17458) );
  AOI211_X1 U20769 ( .C1(n15895), .C2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n17459), .B(n17458), .ZN(n17644) );
  NOR2_X1 U20770 ( .A1(n17530), .A2(n17461), .ZN(n17479) );
  NOR2_X1 U20771 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17578), .ZN(n17460) );
  AOI22_X1 U20772 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17479), .B1(n17461), 
        .B2(n17460), .ZN(n17462) );
  OAI21_X1 U20773 ( .B1(n17644), .B2(n17525), .A(n17462), .ZN(P3_U2693) );
  AOI22_X1 U20774 ( .A1(n9689), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n12952), .ZN(n17463) );
  OAI21_X1 U20775 ( .B1(n17464), .B2(n9755), .A(n17463), .ZN(n17478) );
  INV_X1 U20776 ( .A(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17476) );
  AOI22_X1 U20777 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17430), .B1(
        n17449), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17475) );
  AOI22_X1 U20778 ( .A1(n17490), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17465), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17466) );
  OAI21_X1 U20779 ( .B1(n18501), .B2(n17486), .A(n17466), .ZN(n17473) );
  AOI22_X1 U20780 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n15828), .B1(
        n9685), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17469) );
  AOI22_X1 U20781 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17467), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n9704), .ZN(n17468) );
  OAI211_X1 U20782 ( .C1(n17471), .C2(n17470), .A(n17469), .B(n17468), .ZN(
        n17472) );
  AOI211_X1 U20783 ( .C1(n17489), .C2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n17473), .B(n17472), .ZN(n17474) );
  OAI211_X1 U20784 ( .C1(n17476), .C2(n12984), .A(n17475), .B(n17474), .ZN(
        n17477) );
  AOI211_X1 U20785 ( .C1(n15895), .C2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A(
        n17478), .B(n17477), .ZN(n17647) );
  OAI21_X1 U20786 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17480), .A(n17479), .ZN(
        n17481) );
  OAI21_X1 U20787 ( .B1(n17647), .B2(n17525), .A(n17481), .ZN(P3_U2694) );
  AOI22_X1 U20788 ( .A1(n17288), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17482), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17498) );
  AOI22_X1 U20789 ( .A1(n17449), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17483) );
  OAI21_X1 U20790 ( .B1(n12977), .B2(n17484), .A(n17483), .ZN(n17496) );
  OAI22_X1 U20791 ( .A1(n17486), .A2(n18496), .B1(n17485), .B2(n18900), .ZN(
        n17487) );
  AOI21_X1 U20792 ( .B1(n17488), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n17487), .ZN(n17494) );
  AOI22_X1 U20793 ( .A1(n17430), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15894), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17493) );
  AOI22_X1 U20794 ( .A1(n15895), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9685), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17492) );
  AOI22_X1 U20795 ( .A1(n17490), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17489), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17491) );
  NAND4_X1 U20796 ( .A1(n17494), .A2(n17493), .A3(n17492), .A4(n17491), .ZN(
        n17495) );
  AOI211_X1 U20797 ( .C1(n9689), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n17496), .B(n17495), .ZN(n17497) );
  OAI211_X1 U20798 ( .C1(n12959), .C2(n18802), .A(n17498), .B(n17497), .ZN(
        n17651) );
  INV_X1 U20799 ( .A(n17651), .ZN(n17502) );
  INV_X1 U20800 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17508) );
  NOR3_X1 U20801 ( .A1(n17499), .A2(n17508), .A3(n17505), .ZN(n17504) );
  OAI21_X1 U20802 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17504), .A(n17500), .ZN(
        n17501) );
  AOI22_X1 U20803 ( .A1(n17530), .A2(n17502), .B1(n17501), .B2(n17525), .ZN(
        P3_U2695) );
  NOR2_X1 U20804 ( .A1(n17578), .A2(n17505), .ZN(n17506) );
  AOI22_X1 U20805 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17525), .B1(
        P3_EBX_REG_6__SCAN_IN), .B2(n17506), .ZN(n17503) );
  OAI22_X1 U20806 ( .A1(n17504), .A2(n17503), .B1(n18537), .B2(n17525), .ZN(
        P3_U2696) );
  NAND2_X1 U20807 ( .A1(n17525), .A2(n17505), .ZN(n17510) );
  AOI22_X1 U20808 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17530), .B1(
        n17506), .B2(n17508), .ZN(n17507) );
  OAI21_X1 U20809 ( .B1(n17508), .B2(n17510), .A(n17507), .ZN(P3_U2697) );
  NOR2_X1 U20810 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17509), .ZN(n17511) );
  OAI22_X1 U20811 ( .A1(n17511), .A2(n17510), .B1(n18523), .B2(n17525), .ZN(
        P3_U2698) );
  NAND2_X1 U20812 ( .A1(n17512), .A2(n17529), .ZN(n17522) );
  NOR2_X1 U20813 ( .A1(n17513), .A2(n17522), .ZN(n17518) );
  OAI211_X1 U20814 ( .C1(n17518), .C2(P3_EBX_REG_4__SCAN_IN), .A(n17525), .B(
        n17514), .ZN(n17515) );
  OAI21_X1 U20815 ( .B1(n17525), .B2(n18517), .A(n17515), .ZN(P3_U2699) );
  INV_X1 U20816 ( .A(n17522), .ZN(n17516) );
  AOI21_X1 U20817 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17525), .A(n17516), .ZN(
        n17517) );
  OAI22_X1 U20818 ( .A1(n17518), .A2(n17517), .B1(n18512), .B2(n17525), .ZN(
        P3_U2700) );
  OAI221_X1 U20819 ( .B1(n17521), .B2(n17520), .C1(n18533), .C2(n17520), .A(
        n17519), .ZN(n17523) );
  OAI211_X1 U20820 ( .C1(n17525), .C2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n17523), .B(n17522), .ZN(n17524) );
  INV_X1 U20821 ( .A(n17524), .ZN(P3_U2701) );
  OAI222_X1 U20822 ( .A1(n17528), .A2(n17527), .B1(n17526), .B2(n17533), .C1(
        n18501), .C2(n17525), .ZN(P3_U2702) );
  AOI22_X1 U20823 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17530), .B1(
        n17529), .B2(n17532), .ZN(n17531) );
  OAI21_X1 U20824 ( .B1(n17533), .B2(n17532), .A(n17531), .ZN(P3_U2703) );
  INV_X1 U20825 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17753) );
  INV_X1 U20826 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17749) );
  INV_X1 U20827 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17793) );
  NAND2_X1 U20828 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n17674) );
  INV_X1 U20829 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17769) );
  INV_X1 U20830 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17767) );
  NAND4_X1 U20831 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17534) );
  NOR4_X1 U20832 ( .A1(n17674), .A2(n17769), .A3(n17767), .A4(n17534), .ZN(
        n17620) );
  NAND2_X1 U20833 ( .A1(n17537), .A2(n17620), .ZN(n17652) );
  NAND4_X1 U20834 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n17535)
         );
  NAND3_X1 U20835 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .ZN(n17579) );
  NAND3_X1 U20836 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_22__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .ZN(n17536) );
  NAND2_X1 U20837 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17557), .ZN(n17554) );
  NAND2_X1 U20838 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17548), .ZN(n17545) );
  NAND2_X1 U20839 ( .A1(n17540), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17539) );
  NOR2_X2 U20840 ( .A1(n17538), .A2(n17680), .ZN(n17611) );
  AOI22_X1 U20841 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17611), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17610), .ZN(n17542) );
  OAI211_X1 U20842 ( .C1(n17540), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17680), .B(
        n17539), .ZN(n17541) );
  OAI211_X1 U20843 ( .C1(n17543), .C2(n17676), .A(n17542), .B(n17541), .ZN(
        P3_U2705) );
  INV_X1 U20844 ( .A(n17610), .ZN(n17567) );
  AOI22_X1 U20845 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17611), .B1(n17683), .B2(
        n17544), .ZN(n17547) );
  OAI211_X1 U20846 ( .C1(n17548), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17680), .B(
        n17545), .ZN(n17546) );
  OAI211_X1 U20847 ( .C1(n17567), .C2(n18519), .A(n17547), .B(n17546), .ZN(
        P3_U2706) );
  AOI22_X1 U20848 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17611), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17610), .ZN(n17551) );
  AOI211_X1 U20849 ( .C1(n17753), .C2(n17554), .A(n17548), .B(n17641), .ZN(
        n17549) );
  INV_X1 U20850 ( .A(n17549), .ZN(n17550) );
  OAI211_X1 U20851 ( .C1(n17552), .C2(n17676), .A(n17551), .B(n17550), .ZN(
        P3_U2707) );
  AOI22_X1 U20852 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17611), .B1(n17683), .B2(
        n17553), .ZN(n17556) );
  OAI211_X1 U20853 ( .C1(n17557), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17680), .B(
        n17554), .ZN(n17555) );
  OAI211_X1 U20854 ( .C1(n17567), .C2(n18508), .A(n17556), .B(n17555), .ZN(
        P3_U2708) );
  AOI22_X1 U20855 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17611), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17610), .ZN(n17560) );
  AOI211_X1 U20856 ( .C1(n17749), .C2(n17563), .A(n17557), .B(n17641), .ZN(
        n17558) );
  INV_X1 U20857 ( .A(n17558), .ZN(n17559) );
  OAI211_X1 U20858 ( .C1(n17561), .C2(n17676), .A(n17560), .B(n17559), .ZN(
        P3_U2709) );
  AOI22_X1 U20859 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17611), .B1(n17683), .B2(
        n17562), .ZN(n17566) );
  OAI211_X1 U20860 ( .C1(n17564), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17680), .B(
        n17563), .ZN(n17565) );
  OAI211_X1 U20861 ( .C1(n17567), .C2(n18497), .A(n17566), .B(n17565), .ZN(
        P3_U2710) );
  AOI22_X1 U20862 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17611), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17610), .ZN(n17570) );
  OAI211_X1 U20863 ( .C1(n9806), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17680), .B(
        n17568), .ZN(n17569) );
  OAI211_X1 U20864 ( .C1(n17571), .C2(n17676), .A(n17570), .B(n17569), .ZN(
        P3_U2711) );
  INV_X1 U20865 ( .A(n17611), .ZN(n17593) );
  AOI22_X1 U20866 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n17610), .B1(n17683), .B2(
        n17572), .ZN(n17576) );
  OAI211_X1 U20867 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17574), .A(n17680), .B(
        n17573), .ZN(n17575) );
  OAI211_X1 U20868 ( .C1(n17593), .C2(n18529), .A(n17576), .B(n17575), .ZN(
        P3_U2712) );
  AOI22_X1 U20869 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17610), .B1(n17683), .B2(
        n17577), .ZN(n17583) );
  INV_X1 U20870 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17735) );
  NOR2_X1 U20871 ( .A1(n17578), .A2(n17612), .ZN(n17606) );
  NAND2_X1 U20872 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17606), .ZN(n17605) );
  NAND3_X1 U20873 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(n17600), .ZN(n17589) );
  NAND2_X1 U20874 ( .A1(n17680), .A2(n17589), .ZN(n17585) );
  OAI21_X1 U20875 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17673), .A(n17585), .ZN(
        n17581) );
  INV_X1 U20876 ( .A(n17600), .ZN(n17595) );
  NOR3_X1 U20877 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17579), .A3(n17595), .ZN(
        n17580) );
  AOI21_X1 U20878 ( .B1(P3_EAX_REG_22__SCAN_IN), .B2(n17581), .A(n17580), .ZN(
        n17582) );
  OAI211_X1 U20879 ( .C1(n18524), .C2(n17593), .A(n17583), .B(n17582), .ZN(
        P3_U2713) );
  AOI22_X1 U20880 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17610), .B1(n17683), .B2(
        n17584), .ZN(n17587) );
  INV_X1 U20881 ( .A(n17585), .ZN(n17590) );
  AOI22_X1 U20882 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17611), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n17590), .ZN(n17586) );
  OAI211_X1 U20883 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n17589), .A(n17587), .B(
        n17586), .ZN(P3_U2714) );
  AOI22_X1 U20884 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17610), .B1(n17683), .B2(
        n17588), .ZN(n17592) );
  INV_X1 U20885 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17737) );
  NOR2_X1 U20886 ( .A1(n17737), .A2(n17595), .ZN(n17594) );
  AOI22_X1 U20887 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17590), .B1(n17594), 
        .B2(n17589), .ZN(n17591) );
  OAI211_X1 U20888 ( .C1(n18513), .C2(n17593), .A(n17592), .B(n17591), .ZN(
        P3_U2715) );
  AOI22_X1 U20889 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17611), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17610), .ZN(n17598) );
  AOI211_X1 U20890 ( .C1(n17737), .C2(n17595), .A(n17594), .B(n17641), .ZN(
        n17596) );
  INV_X1 U20891 ( .A(n17596), .ZN(n17597) );
  OAI211_X1 U20892 ( .C1(n17599), .C2(n17676), .A(n17598), .B(n17597), .ZN(
        P3_U2716) );
  AOI22_X1 U20893 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17611), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17610), .ZN(n17603) );
  AOI211_X1 U20894 ( .C1(n17735), .C2(n17605), .A(n17600), .B(n17641), .ZN(
        n17601) );
  INV_X1 U20895 ( .A(n17601), .ZN(n17602) );
  OAI211_X1 U20896 ( .C1(n17604), .C2(n17676), .A(n17603), .B(n17602), .ZN(
        P3_U2717) );
  AOI22_X1 U20897 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17611), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17610), .ZN(n17608) );
  OAI211_X1 U20898 ( .C1(n17606), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17680), .B(
        n17605), .ZN(n17607) );
  OAI211_X1 U20899 ( .C1(n17609), .C2(n17676), .A(n17608), .B(n17607), .ZN(
        P3_U2718) );
  AOI22_X1 U20900 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17611), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17610), .ZN(n17614) );
  OAI211_X1 U20901 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17616), .A(n17680), .B(
        n17612), .ZN(n17613) );
  OAI211_X1 U20902 ( .C1(n17615), .C2(n17676), .A(n17614), .B(n17613), .ZN(
        P3_U2719) );
  AOI211_X1 U20903 ( .C1(n17793), .C2(n17623), .A(n17641), .B(n17616), .ZN(
        n17617) );
  AOI21_X1 U20904 ( .B1(n17684), .B2(BUF2_REG_15__SCAN_IN), .A(n17617), .ZN(
        n17618) );
  OAI21_X1 U20905 ( .B1(n17619), .B2(n17676), .A(n17618), .ZN(P3_U2720) );
  INV_X1 U20906 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17785) );
  INV_X1 U20907 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17779) );
  INV_X1 U20908 ( .A(n17620), .ZN(n17621) );
  NAND2_X1 U20909 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17646), .ZN(n17645) );
  NAND2_X1 U20910 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17640), .ZN(n17631) );
  NOR2_X1 U20911 ( .A1(n17785), .A2(n17631), .ZN(n17634) );
  NAND2_X1 U20912 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17634), .ZN(n17626) );
  AOI22_X1 U20913 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17684), .B1(n17683), .B2(
        n17622), .ZN(n17625) );
  NAND3_X1 U20914 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17680), .A3(n17623), 
        .ZN(n17624) );
  OAI211_X1 U20915 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17626), .A(n17625), .B(
        n17624), .ZN(P3_U2721) );
  INV_X1 U20916 ( .A(n17626), .ZN(n17629) );
  AOI21_X1 U20917 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17680), .A(n17634), .ZN(
        n17628) );
  OAI222_X1 U20918 ( .A1(n17679), .A2(n17630), .B1(n17629), .B2(n17628), .C1(
        n17676), .C2(n17627), .ZN(P3_U2722) );
  INV_X1 U20919 ( .A(n17631), .ZN(n17638) );
  AOI21_X1 U20920 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17680), .A(n17638), .ZN(
        n17633) );
  OAI222_X1 U20921 ( .A1(n17679), .A2(n17635), .B1(n17634), .B2(n17633), .C1(
        n17676), .C2(n17632), .ZN(P3_U2723) );
  AOI21_X1 U20922 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17680), .A(n17640), .ZN(
        n17637) );
  OAI222_X1 U20923 ( .A1(n17679), .A2(n17639), .B1(n17638), .B2(n17637), .C1(
        n17676), .C2(n17636), .ZN(P3_U2724) );
  AOI211_X1 U20924 ( .C1(n17779), .C2(n17645), .A(n17641), .B(n17640), .ZN(
        n17642) );
  AOI21_X1 U20925 ( .B1(n17684), .B2(BUF2_REG_10__SCAN_IN), .A(n17642), .ZN(
        n17643) );
  OAI21_X1 U20926 ( .B1(n17644), .B2(n17676), .A(n17643), .ZN(P3_U2725) );
  INV_X1 U20927 ( .A(n17645), .ZN(n17649) );
  AOI21_X1 U20928 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17680), .A(n17646), .ZN(
        n17648) );
  OAI222_X1 U20929 ( .A1(n17679), .A2(n17650), .B1(n17649), .B2(n17648), .C1(
        n17676), .C2(n17647), .ZN(P3_U2726) );
  INV_X1 U20930 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17775) );
  AOI22_X1 U20931 ( .A1(n17683), .A2(n17651), .B1(n17658), .B2(n17775), .ZN(
        n17654) );
  NAND3_X1 U20932 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17680), .A3(n17652), .ZN(
        n17653) );
  OAI211_X1 U20933 ( .C1(n17679), .C2(n17655), .A(n17654), .B(n17653), .ZN(
        P3_U2727) );
  INV_X1 U20934 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17771) );
  INV_X1 U20935 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17763) );
  NOR3_X1 U20936 ( .A1(n17674), .A2(n17763), .A3(n17673), .ZN(n17678) );
  NAND2_X1 U20937 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17678), .ZN(n17666) );
  NOR2_X1 U20938 ( .A1(n17767), .A2(n17666), .ZN(n17669) );
  NAND2_X1 U20939 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17669), .ZN(n17659) );
  NOR2_X1 U20940 ( .A1(n17771), .A2(n17659), .ZN(n17662) );
  AOI21_X1 U20941 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17680), .A(n17662), .ZN(
        n17657) );
  OAI222_X1 U20942 ( .A1(n17679), .A2(n18529), .B1(n17658), .B2(n17657), .C1(
        n17676), .C2(n17656), .ZN(P3_U2728) );
  INV_X1 U20943 ( .A(n17659), .ZN(n17665) );
  AOI21_X1 U20944 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17680), .A(n17665), .ZN(
        n17661) );
  OAI222_X1 U20945 ( .A1(n18524), .A2(n17679), .B1(n17662), .B2(n17661), .C1(
        n17676), .C2(n17660), .ZN(P3_U2729) );
  AOI21_X1 U20946 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17680), .A(n17669), .ZN(
        n17664) );
  OAI222_X1 U20947 ( .A1(n18518), .A2(n17679), .B1(n17665), .B2(n17664), .C1(
        n17676), .C2(n17663), .ZN(P3_U2730) );
  INV_X1 U20948 ( .A(n17666), .ZN(n17672) );
  AOI21_X1 U20949 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17680), .A(n17672), .ZN(
        n17668) );
  OAI222_X1 U20950 ( .A1(n18513), .A2(n17679), .B1(n17669), .B2(n17668), .C1(
        n17676), .C2(n17667), .ZN(P3_U2731) );
  AOI21_X1 U20951 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17680), .A(n17678), .ZN(
        n17671) );
  OAI222_X1 U20952 ( .A1(n18507), .A2(n17679), .B1(n17672), .B2(n17671), .C1(
        n17676), .C2(n17670), .ZN(P3_U2732) );
  NOR2_X1 U20953 ( .A1(n17674), .A2(n17673), .ZN(n17687) );
  AOI21_X1 U20954 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17680), .A(n17687), .ZN(
        n17677) );
  OAI222_X1 U20955 ( .A1(n18502), .A2(n17679), .B1(n17678), .B2(n17677), .C1(
        n17676), .C2(n17675), .ZN(P3_U2733) );
  OAI21_X1 U20956 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n17681), .A(n17680), .ZN(
        n17686) );
  AOI22_X1 U20957 ( .A1(n17684), .A2(BUF2_REG_1__SCAN_IN), .B1(n17683), .B2(
        n17682), .ZN(n17685) );
  OAI21_X1 U20958 ( .B1(n17687), .B2(n17686), .A(n17685), .ZN(P3_U2734) );
  AND2_X1 U20959 ( .A1(n17703), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20960 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17757) );
  AOI22_X1 U20961 ( .A1(n19166), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17723), .ZN(n17691) );
  OAI21_X1 U20962 ( .B1(n17757), .B2(n17707), .A(n17691), .ZN(P3_U2737) );
  INV_X1 U20963 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17755) );
  AOI22_X1 U20964 ( .A1(n19166), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17692) );
  OAI21_X1 U20965 ( .B1(n17755), .B2(n17707), .A(n17692), .ZN(P3_U2738) );
  AOI22_X1 U20966 ( .A1(n19166), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17703), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17693) );
  OAI21_X1 U20967 ( .B1(n17753), .B2(n17707), .A(n17693), .ZN(P3_U2739) );
  INV_X1 U20968 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17751) );
  AOI22_X1 U20969 ( .A1(n19166), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17703), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17694) );
  OAI21_X1 U20970 ( .B1(n17751), .B2(n17707), .A(n17694), .ZN(P3_U2740) );
  AOI22_X1 U20971 ( .A1(n19166), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17695) );
  OAI21_X1 U20972 ( .B1(n17749), .B2(n17707), .A(n17695), .ZN(P3_U2741) );
  INV_X1 U20973 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17747) );
  AOI22_X1 U20974 ( .A1(n19166), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17703), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17696) );
  OAI21_X1 U20975 ( .B1(n17747), .B2(n17707), .A(n17696), .ZN(P3_U2742) );
  AOI22_X1 U20976 ( .A1(n19166), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17703), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17697) );
  OAI21_X1 U20977 ( .B1(n9871), .B2(n17707), .A(n17697), .ZN(P3_U2743) );
  AOI22_X1 U20978 ( .A1(n17724), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17703), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17698) );
  OAI21_X1 U20979 ( .B1(n9870), .B2(n17707), .A(n17698), .ZN(P3_U2744) );
  INV_X1 U20980 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17743) );
  AOI22_X1 U20981 ( .A1(n17724), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17703), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17699) );
  OAI21_X1 U20982 ( .B1(n17743), .B2(n17707), .A(n17699), .ZN(P3_U2745) );
  INV_X1 U20983 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17741) );
  AOI22_X1 U20984 ( .A1(n17724), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17703), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17700) );
  OAI21_X1 U20985 ( .B1(n17741), .B2(n17707), .A(n17700), .ZN(P3_U2746) );
  INV_X1 U20986 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17739) );
  AOI22_X1 U20987 ( .A1(n17724), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17703), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17701) );
  OAI21_X1 U20988 ( .B1(n17739), .B2(n17707), .A(n17701), .ZN(P3_U2747) );
  AOI22_X1 U20989 ( .A1(n17724), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17703), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17702) );
  OAI21_X1 U20990 ( .B1(n17737), .B2(n17707), .A(n17702), .ZN(P3_U2748) );
  AOI22_X1 U20991 ( .A1(n17724), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17703), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17704) );
  OAI21_X1 U20992 ( .B1(n17735), .B2(n17707), .A(n17704), .ZN(P3_U2749) );
  INV_X1 U20993 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17733) );
  AOI22_X1 U20994 ( .A1(n17724), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17705) );
  OAI21_X1 U20995 ( .B1(n17733), .B2(n17707), .A(n17705), .ZN(P3_U2750) );
  INV_X1 U20996 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17731) );
  AOI22_X1 U20997 ( .A1(n17724), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17706) );
  OAI21_X1 U20998 ( .B1(n17731), .B2(n17707), .A(n17706), .ZN(P3_U2751) );
  AOI22_X1 U20999 ( .A1(n17724), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17708) );
  OAI21_X1 U21000 ( .B1(n17793), .B2(n17726), .A(n17708), .ZN(P3_U2752) );
  INV_X1 U21001 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17789) );
  AOI22_X1 U21002 ( .A1(n17724), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17709) );
  OAI21_X1 U21003 ( .B1(n17789), .B2(n17726), .A(n17709), .ZN(P3_U2753) );
  INV_X1 U21004 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17787) );
  AOI22_X1 U21005 ( .A1(n17724), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17710) );
  OAI21_X1 U21006 ( .B1(n17787), .B2(n17726), .A(n17710), .ZN(P3_U2754) );
  AOI22_X1 U21007 ( .A1(n17724), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17711) );
  OAI21_X1 U21008 ( .B1(n17785), .B2(n17726), .A(n17711), .ZN(P3_U2755) );
  INV_X1 U21009 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17781) );
  AOI22_X1 U21010 ( .A1(n17724), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17712) );
  OAI21_X1 U21011 ( .B1(n17781), .B2(n17726), .A(n17712), .ZN(P3_U2756) );
  AOI22_X1 U21012 ( .A1(n17724), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17713) );
  OAI21_X1 U21013 ( .B1(n17779), .B2(n17726), .A(n17713), .ZN(P3_U2757) );
  INV_X1 U21014 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17777) );
  AOI22_X1 U21015 ( .A1(n17724), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17714) );
  OAI21_X1 U21016 ( .B1(n17777), .B2(n17726), .A(n17714), .ZN(P3_U2758) );
  AOI22_X1 U21017 ( .A1(n17724), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17715) );
  OAI21_X1 U21018 ( .B1(n17775), .B2(n17726), .A(n17715), .ZN(P3_U2759) );
  INV_X1 U21019 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17773) );
  AOI22_X1 U21020 ( .A1(n17724), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17716) );
  OAI21_X1 U21021 ( .B1(n17773), .B2(n17726), .A(n17716), .ZN(P3_U2760) );
  AOI22_X1 U21022 ( .A1(n17724), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17717) );
  OAI21_X1 U21023 ( .B1(n17771), .B2(n17726), .A(n17717), .ZN(P3_U2761) );
  AOI22_X1 U21024 ( .A1(n17724), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17718) );
  OAI21_X1 U21025 ( .B1(n17769), .B2(n17726), .A(n17718), .ZN(P3_U2762) );
  AOI22_X1 U21026 ( .A1(n17724), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17719) );
  OAI21_X1 U21027 ( .B1(n17767), .B2(n17726), .A(n17719), .ZN(P3_U2763) );
  INV_X1 U21028 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17765) );
  AOI22_X1 U21029 ( .A1(n17724), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17720) );
  OAI21_X1 U21030 ( .B1(n17765), .B2(n17726), .A(n17720), .ZN(P3_U2764) );
  AOI22_X1 U21031 ( .A1(n17724), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17721) );
  OAI21_X1 U21032 ( .B1(n17763), .B2(n17726), .A(n17721), .ZN(P3_U2765) );
  INV_X1 U21033 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17761) );
  AOI22_X1 U21034 ( .A1(n17724), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17722) );
  OAI21_X1 U21035 ( .B1(n17761), .B2(n17726), .A(n17722), .ZN(P3_U2766) );
  AOI22_X1 U21036 ( .A1(n17724), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17723), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17725) );
  OAI21_X1 U21037 ( .B1(n17759), .B2(n17726), .A(n17725), .ZN(P3_U2767) );
  AOI22_X1 U21038 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17783), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17782), .ZN(n17730) );
  OAI21_X1 U21039 ( .B1(n17731), .B2(n17792), .A(n17730), .ZN(P3_U2768) );
  AOI22_X1 U21040 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17783), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17782), .ZN(n17732) );
  OAI21_X1 U21041 ( .B1(n17733), .B2(n17792), .A(n17732), .ZN(P3_U2769) );
  AOI22_X1 U21042 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17783), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17782), .ZN(n17734) );
  OAI21_X1 U21043 ( .B1(n17735), .B2(n17792), .A(n17734), .ZN(P3_U2770) );
  AOI22_X1 U21044 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n9723), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17782), .ZN(n17736) );
  OAI21_X1 U21045 ( .B1(n17737), .B2(n17792), .A(n17736), .ZN(P3_U2771) );
  AOI22_X1 U21046 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n9723), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17782), .ZN(n17738) );
  OAI21_X1 U21047 ( .B1(n17739), .B2(n17792), .A(n17738), .ZN(P3_U2772) );
  AOI22_X1 U21048 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n9723), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17782), .ZN(n17740) );
  OAI21_X1 U21049 ( .B1(n17741), .B2(n17792), .A(n17740), .ZN(P3_U2773) );
  AOI22_X1 U21050 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n9723), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17782), .ZN(n17742) );
  OAI21_X1 U21051 ( .B1(n17743), .B2(n17792), .A(n17742), .ZN(P3_U2774) );
  AOI22_X1 U21052 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n9723), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17782), .ZN(n17744) );
  OAI21_X1 U21053 ( .B1(n9870), .B2(n17792), .A(n17744), .ZN(P3_U2775) );
  AOI22_X1 U21054 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n9723), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17782), .ZN(n17745) );
  OAI21_X1 U21055 ( .B1(n9871), .B2(n17792), .A(n17745), .ZN(P3_U2776) );
  AOI22_X1 U21056 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n9723), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17782), .ZN(n17746) );
  OAI21_X1 U21057 ( .B1(n17747), .B2(n17792), .A(n17746), .ZN(P3_U2777) );
  AOI22_X1 U21058 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n9723), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17782), .ZN(n17748) );
  OAI21_X1 U21059 ( .B1(n17749), .B2(n17792), .A(n17748), .ZN(P3_U2778) );
  AOI22_X1 U21060 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n9723), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17782), .ZN(n17750) );
  OAI21_X1 U21061 ( .B1(n17751), .B2(n17792), .A(n17750), .ZN(P3_U2779) );
  AOI22_X1 U21062 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17783), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17782), .ZN(n17752) );
  OAI21_X1 U21063 ( .B1(n17753), .B2(n17792), .A(n17752), .ZN(P3_U2780) );
  AOI22_X1 U21064 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17783), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17782), .ZN(n17754) );
  OAI21_X1 U21065 ( .B1(n17755), .B2(n17792), .A(n17754), .ZN(P3_U2781) );
  AOI22_X1 U21066 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17783), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17782), .ZN(n17756) );
  OAI21_X1 U21067 ( .B1(n17757), .B2(n17792), .A(n17756), .ZN(P3_U2782) );
  AOI22_X1 U21068 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17783), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17782), .ZN(n17758) );
  OAI21_X1 U21069 ( .B1(n17759), .B2(n17792), .A(n17758), .ZN(P3_U2783) );
  AOI22_X1 U21070 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17783), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17782), .ZN(n17760) );
  OAI21_X1 U21071 ( .B1(n17761), .B2(n17792), .A(n17760), .ZN(P3_U2784) );
  AOI22_X1 U21072 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17783), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17782), .ZN(n17762) );
  OAI21_X1 U21073 ( .B1(n17763), .B2(n17792), .A(n17762), .ZN(P3_U2785) );
  AOI22_X1 U21074 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17783), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17782), .ZN(n17764) );
  OAI21_X1 U21075 ( .B1(n17765), .B2(n17792), .A(n17764), .ZN(P3_U2786) );
  AOI22_X1 U21076 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17783), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17790), .ZN(n17766) );
  OAI21_X1 U21077 ( .B1(n17767), .B2(n17792), .A(n17766), .ZN(P3_U2787) );
  AOI22_X1 U21078 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17783), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17790), .ZN(n17768) );
  OAI21_X1 U21079 ( .B1(n17769), .B2(n17792), .A(n17768), .ZN(P3_U2788) );
  AOI22_X1 U21080 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17783), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17790), .ZN(n17770) );
  OAI21_X1 U21081 ( .B1(n17771), .B2(n17792), .A(n17770), .ZN(P3_U2789) );
  AOI22_X1 U21082 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17783), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17790), .ZN(n17772) );
  OAI21_X1 U21083 ( .B1(n17773), .B2(n17792), .A(n17772), .ZN(P3_U2790) );
  AOI22_X1 U21084 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17783), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17790), .ZN(n17774) );
  OAI21_X1 U21085 ( .B1(n17775), .B2(n17792), .A(n17774), .ZN(P3_U2791) );
  AOI22_X1 U21086 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17783), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17790), .ZN(n17776) );
  OAI21_X1 U21087 ( .B1(n17777), .B2(n17792), .A(n17776), .ZN(P3_U2792) );
  AOI22_X1 U21088 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n9723), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17782), .ZN(n17778) );
  OAI21_X1 U21089 ( .B1(n17779), .B2(n17792), .A(n17778), .ZN(P3_U2793) );
  AOI22_X1 U21090 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17783), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17790), .ZN(n17780) );
  OAI21_X1 U21091 ( .B1(n17781), .B2(n17792), .A(n17780), .ZN(P3_U2794) );
  AOI22_X1 U21092 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n9723), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17782), .ZN(n17784) );
  OAI21_X1 U21093 ( .B1(n17785), .B2(n17792), .A(n17784), .ZN(P3_U2795) );
  AOI22_X1 U21094 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17783), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17790), .ZN(n17786) );
  OAI21_X1 U21095 ( .B1(n17787), .B2(n17792), .A(n17786), .ZN(P3_U2796) );
  AOI22_X1 U21096 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17783), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17790), .ZN(n17788) );
  OAI21_X1 U21097 ( .B1(n17789), .B2(n17792), .A(n17788), .ZN(P3_U2797) );
  AOI22_X1 U21098 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17783), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17790), .ZN(n17791) );
  OAI21_X1 U21099 ( .B1(n17793), .B2(n17792), .A(n17791), .ZN(P3_U2798) );
  OAI22_X1 U21100 ( .A1(n17796), .A2(n18105), .B1(n17794), .B2(n18148), .ZN(
        n17795) );
  NOR2_X1 U21101 ( .A1(n18118), .A2(n17795), .ZN(n17827) );
  OAI21_X1 U21102 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17899), .A(
        n17827), .ZN(n17815) );
  NAND2_X1 U21103 ( .A1(n17796), .A2(n17983), .ZN(n17817) );
  OAI21_X1 U21104 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17797), .ZN(n17798) );
  OAI22_X1 U21105 ( .A1(n17990), .A2(n17799), .B1(n17817), .B2(n17798), .ZN(
        n17800) );
  AOI211_X1 U21106 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17815), .A(
        n17801), .B(n17800), .ZN(n17811) );
  NOR2_X1 U21107 ( .A1(n18136), .A2(n18008), .ZN(n17905) );
  OAI22_X1 U21108 ( .A1(n18155), .A2(n18152), .B1(n17802), .B2(n9662), .ZN(
        n17831) );
  NOR2_X1 U21109 ( .A1(n17821), .A2(n17831), .ZN(n17822) );
  NOR3_X1 U21110 ( .A1(n17905), .A2(n17822), .A3(n17803), .ZN(n17804) );
  AOI21_X1 U21111 ( .B1(n17805), .B2(n9753), .A(n17804), .ZN(n17810) );
  OAI211_X1 U21112 ( .C1(n17808), .C2(n17807), .A(n18058), .B(n17806), .ZN(
        n17809) );
  NAND3_X1 U21113 ( .A1(n17811), .A2(n17810), .A3(n17809), .ZN(P3_U2802) );
  NOR2_X1 U21114 ( .A1(n17812), .A2(n16686), .ZN(n17813) );
  XNOR2_X1 U21115 ( .A(n17813), .B(n18057), .ZN(n18169) );
  AOI22_X1 U21116 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17815), .B1(
        n18004), .B2(n17814), .ZN(n17816) );
  NAND2_X1 U21117 ( .A1(n18408), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18170) );
  OAI211_X1 U21118 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17817), .A(
        n17816), .B(n18170), .ZN(n17818) );
  AOI21_X1 U21119 ( .B1(n18058), .B2(n18169), .A(n17818), .ZN(n17819) );
  OAI221_X1 U21120 ( .B1(n17822), .B2(n17821), .C1(n17822), .C2(n17820), .A(
        n17819), .ZN(P3_U2803) );
  AOI21_X1 U21121 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17824), .A(
        n17823), .ZN(n18177) );
  INV_X1 U21122 ( .A(n17899), .ZN(n17829) );
  AOI21_X1 U21123 ( .B1(n17825), .B2(n18891), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17826) );
  OAI22_X1 U21124 ( .A1(n17827), .A2(n17826), .B1(n18375), .B2(n19097), .ZN(
        n17828) );
  AOI221_X1 U21125 ( .B1(n18004), .B2(n17830), .C1(n17829), .C2(n17830), .A(
        n17828), .ZN(n17833) );
  NOR3_X1 U21126 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18180), .A3(
        n18160), .ZN(n18173) );
  AOI22_X1 U21127 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17831), .B1(
        n9753), .B2(n18173), .ZN(n17832) );
  OAI211_X1 U21128 ( .C1(n18177), .C2(n18044), .A(n17833), .B(n17832), .ZN(
        P3_U2804) );
  XNOR2_X1 U21129 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17834), .ZN(
        n18187) );
  AND2_X1 U21130 ( .A1(n17836), .A2(n18891), .ZN(n17862) );
  AOI211_X1 U21131 ( .C1(n17987), .C2(n17835), .A(n18118), .B(n17862), .ZN(
        n17864) );
  OAI21_X1 U21132 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17899), .A(
        n17864), .ZN(n17852) );
  INV_X1 U21133 ( .A(n17983), .ZN(n17946) );
  NOR2_X1 U21134 ( .A1(n17946), .A2(n17836), .ZN(n17854) );
  OAI211_X1 U21135 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17854), .B(n17837), .ZN(n17838) );
  NAND2_X1 U21136 ( .A1(n18408), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18182) );
  OAI211_X1 U21137 ( .C1(n17990), .C2(n17839), .A(n17838), .B(n18182), .ZN(
        n17845) );
  XNOR2_X1 U21138 ( .A(n17840), .B(n18180), .ZN(n18191) );
  OAI21_X1 U21139 ( .B1(n17968), .B2(n17842), .A(n17841), .ZN(n17843) );
  XNOR2_X1 U21140 ( .A(n17843), .B(n18180), .ZN(n18186) );
  OAI22_X1 U21141 ( .A1(n18152), .A2(n18191), .B1(n18044), .B2(n18186), .ZN(
        n17844) );
  AOI211_X1 U21142 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17852), .A(
        n17845), .B(n17844), .ZN(n17846) );
  OAI21_X1 U21143 ( .B1(n9662), .B2(n18187), .A(n17846), .ZN(P3_U2805) );
  AOI21_X1 U21144 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17848), .A(
        n17847), .ZN(n18207) );
  INV_X1 U21145 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19093) );
  INV_X1 U21146 ( .A(n17849), .ZN(n17850) );
  OAI22_X1 U21147 ( .A1(n18375), .A2(n19093), .B1(n17990), .B2(n17850), .ZN(
        n17851) );
  AOI221_X1 U21148 ( .B1(n17854), .B2(n17853), .C1(n17852), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17851), .ZN(n17857) );
  NOR2_X1 U21149 ( .A1(n17855), .A2(n17872), .ZN(n18193) );
  NOR2_X1 U21150 ( .A1(n17873), .A2(n17855), .ZN(n18192) );
  OAI22_X1 U21151 ( .A1(n18193), .A2(n9662), .B1(n18192), .B2(n18152), .ZN(
        n17866) );
  NOR2_X1 U21152 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18197), .ZN(
        n18203) );
  AOI22_X1 U21153 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17866), .B1(
        n9753), .B2(n18203), .ZN(n17856) );
  OAI211_X1 U21154 ( .C1(n18207), .C2(n18044), .A(n17857), .B(n17856), .ZN(
        P3_U2806) );
  AOI22_X1 U21155 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17968), .B1(
        n17858), .B2(n17870), .ZN(n17859) );
  NAND2_X1 U21156 ( .A1(n17897), .A2(n17859), .ZN(n17860) );
  XNOR2_X1 U21157 ( .A(n17860), .B(n18197), .ZN(n18213) );
  NAND2_X1 U21158 ( .A1(n17990), .A2(n17899), .ZN(n18139) );
  AOI22_X1 U21159 ( .A1(n9820), .A2(n17862), .B1(n17861), .B2(n18139), .ZN(
        n17863) );
  NAND2_X1 U21160 ( .A1(n18408), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18212) );
  OAI211_X1 U21161 ( .C1(n17864), .C2(n9923), .A(n17863), .B(n18212), .ZN(
        n17865) );
  AOI221_X1 U21162 ( .B1(n9753), .B2(n18197), .C1(n17866), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17865), .ZN(n17867) );
  OAI21_X1 U21163 ( .B1(n18044), .B2(n18213), .A(n17867), .ZN(P3_U2807) );
  INV_X1 U21164 ( .A(n17868), .ZN(n17942) );
  INV_X1 U21165 ( .A(n17897), .ZN(n17869) );
  AOI221_X1 U21166 ( .B1(n17942), .B2(n17870), .C1(n18158), .C2(n17870), .A(
        n17869), .ZN(n17871) );
  XNOR2_X1 U21167 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17871), .ZN(
        n18228) );
  NOR2_X1 U21168 ( .A1(n18158), .A2(n17954), .ZN(n17882) );
  INV_X1 U21169 ( .A(n18158), .ZN(n18218) );
  AOI22_X1 U21170 ( .A1(n18136), .A2(n17873), .B1(n18008), .B2(n17872), .ZN(
        n17953) );
  OAI21_X1 U21171 ( .B1(n18218), .B2(n17905), .A(n17953), .ZN(n17894) );
  OAI21_X1 U21172 ( .B1(n17874), .B2(n18148), .A(n18147), .ZN(n17875) );
  AOI21_X1 U21173 ( .B1(n18048), .B2(n17877), .A(n17875), .ZN(n17902) );
  OAI21_X1 U21174 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17899), .A(
        n17902), .ZN(n17891) );
  AOI22_X1 U21175 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17891), .B1(
        n18004), .B2(n17876), .ZN(n17880) );
  NOR2_X1 U21176 ( .A1(n17946), .A2(n17877), .ZN(n17893) );
  OAI211_X1 U21177 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17893), .B(n17878), .ZN(n17879) );
  OAI211_X1 U21178 ( .C1(n19089), .C2(n18375), .A(n17880), .B(n17879), .ZN(
        n17881) );
  AOI221_X1 U21179 ( .B1(n17882), .B2(n18157), .C1(n17894), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n17881), .ZN(n17883) );
  OAI21_X1 U21180 ( .B1(n18044), .B2(n18228), .A(n17883), .ZN(P3_U2808) );
  INV_X1 U21181 ( .A(n18221), .ZN(n18234) );
  NOR3_X1 U21182 ( .A1(n17921), .A2(n17968), .A3(n17884), .ZN(n17908) );
  INV_X1 U21183 ( .A(n17885), .ZN(n17909) );
  AOI22_X1 U21184 ( .A1(n18234), .A2(n17908), .B1(n17909), .B2(n17886), .ZN(
        n17887) );
  XNOR2_X1 U21185 ( .A(n17887), .B(n18220), .ZN(n18238) );
  AOI22_X1 U21186 ( .A1(n18435), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18004), 
        .B2(n17888), .ZN(n17889) );
  INV_X1 U21187 ( .A(n17889), .ZN(n17890) );
  AOI221_X1 U21188 ( .B1(n17893), .B2(n17892), .C1(n17891), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17890), .ZN(n17896) );
  NOR2_X1 U21189 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18221), .ZN(
        n18230) );
  NAND2_X1 U21190 ( .A1(n18261), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18231) );
  NOR2_X1 U21191 ( .A1(n17954), .A2(n18231), .ZN(n17919) );
  AOI22_X1 U21192 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17894), .B1(
        n18230), .B2(n17919), .ZN(n17895) );
  OAI211_X1 U21193 ( .C1(n18238), .C2(n18044), .A(n17896), .B(n17895), .ZN(
        P3_U2809) );
  OAI221_X1 U21194 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17927), 
        .C1(n18248), .C2(n17908), .A(n17897), .ZN(n17898) );
  XOR2_X1 U21195 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17898), .Z(
        n18247) );
  AOI21_X1 U21196 ( .B1(n17900), .B2(n18891), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17901) );
  OAI22_X1 U21197 ( .A1(n17902), .A2(n17901), .B1(n18375), .B2(n19085), .ZN(
        n17903) );
  AOI221_X1 U21198 ( .B1(n18004), .B2(n17904), .C1(n17829), .C2(n17904), .A(
        n17903), .ZN(n17907) );
  NOR2_X1 U21199 ( .A1(n18248), .A2(n18231), .ZN(n18243) );
  OAI21_X1 U21200 ( .B1(n17905), .B2(n18243), .A(n17953), .ZN(n17918) );
  NOR2_X1 U21201 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18248), .ZN(
        n18239) );
  AOI22_X1 U21202 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17918), .B1(
        n17919), .B2(n18239), .ZN(n17906) );
  OAI211_X1 U21203 ( .C1(n18044), .C2(n18247), .A(n17907), .B(n17906), .ZN(
        P3_U2810) );
  AOI21_X1 U21204 ( .B1(n17909), .B2(n17927), .A(n17908), .ZN(n17910) );
  XNOR2_X1 U21205 ( .A(n17910), .B(n18248), .ZN(n18253) );
  AOI21_X1 U21206 ( .B1(n18048), .B2(n17912), .A(n18118), .ZN(n17932) );
  OAI21_X1 U21207 ( .B1(n17911), .B2(n18148), .A(n17932), .ZN(n17924) );
  AOI22_X1 U21208 ( .A1(n18408), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17924), .ZN(n17915) );
  NOR2_X1 U21209 ( .A1(n17946), .A2(n17912), .ZN(n17926) );
  OAI211_X1 U21210 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17926), .B(n17913), .ZN(n17914) );
  OAI211_X1 U21211 ( .C1(n17990), .C2(n17916), .A(n17915), .B(n17914), .ZN(
        n17917) );
  AOI221_X1 U21212 ( .B1(n17919), .B2(n18248), .C1(n17918), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17917), .ZN(n17920) );
  OAI21_X1 U21213 ( .B1(n18253), .B2(n18044), .A(n17920), .ZN(P3_U2811) );
  NAND2_X1 U21214 ( .A1(n18261), .A2(n17921), .ZN(n18268) );
  OAI22_X1 U21215 ( .A1(n18375), .A2(n19081), .B1(n17990), .B2(n17922), .ZN(
        n17923) );
  AOI221_X1 U21216 ( .B1(n17926), .B2(n17925), .C1(n17924), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17923), .ZN(n17930) );
  OAI21_X1 U21217 ( .B1(n18261), .B2(n17954), .A(n17953), .ZN(n17938) );
  AOI21_X1 U21218 ( .B1(n18057), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17927), .ZN(n17928) );
  XNOR2_X1 U21219 ( .A(n17928), .B(n17885), .ZN(n18264) );
  AOI22_X1 U21220 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17938), .B1(
        n18058), .B2(n18264), .ZN(n17929) );
  OAI211_X1 U21221 ( .C1(n17954), .C2(n18268), .A(n17930), .B(n17929), .ZN(
        P3_U2812) );
  NAND2_X1 U21222 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18269), .ZN(
        n18275) );
  INV_X1 U21223 ( .A(n17931), .ZN(n17935) );
  AOI21_X1 U21224 ( .B1(n9797), .B2(n18891), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17933) );
  NAND2_X1 U21225 ( .A1(n18408), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18273) );
  OAI21_X1 U21226 ( .B1(n17933), .B2(n17932), .A(n18273), .ZN(n17934) );
  AOI21_X1 U21227 ( .B1(n17935), .B2(n18139), .A(n17934), .ZN(n17940) );
  OAI21_X1 U21228 ( .B1(n17937), .B2(n18269), .A(n17936), .ZN(n18272) );
  AOI22_X1 U21229 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17938), .B1(
        n18058), .B2(n18272), .ZN(n17939) );
  OAI211_X1 U21230 ( .C1(n17954), .C2(n18275), .A(n17940), .B(n17939), .ZN(
        P3_U2813) );
  AOI21_X1 U21231 ( .B1(n18057), .B2(n17942), .A(n17941), .ZN(n17943) );
  XNOR2_X1 U21232 ( .A(n17943), .B(n18285), .ZN(n18282) );
  AOI21_X1 U21233 ( .B1(n18048), .B2(n17945), .A(n18118), .ZN(n17972) );
  OAI21_X1 U21234 ( .B1(n17944), .B2(n18148), .A(n17972), .ZN(n17961) );
  AOI22_X1 U21235 ( .A1(n18435), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17961), .ZN(n17949) );
  NOR2_X1 U21236 ( .A1(n17946), .A2(n17945), .ZN(n17963) );
  OAI211_X1 U21237 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17963), .B(n17947), .ZN(n17948) );
  OAI211_X1 U21238 ( .C1(n17990), .C2(n17950), .A(n17949), .B(n17948), .ZN(
        n17951) );
  AOI21_X1 U21239 ( .B1(n18058), .B2(n18282), .A(n17951), .ZN(n17952) );
  OAI221_X1 U21240 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17954), 
        .C1(n18285), .C2(n17953), .A(n17952), .ZN(P3_U2814) );
  INV_X1 U21241 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18314) );
  OAI21_X1 U21242 ( .B1(n17956), .B2(n17979), .A(n17955), .ZN(n17957) );
  OAI221_X1 U21243 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18314), 
        .C1(n17997), .C2(n18057), .A(n17957), .ZN(n17958) );
  XOR2_X1 U21244 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17958), .Z(
        n18295) );
  INV_X1 U21245 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17962) );
  OAI22_X1 U21246 ( .A1(n18375), .A2(n19075), .B1(n17990), .B2(n17959), .ZN(
        n17960) );
  AOI221_X1 U21247 ( .B1(n17963), .B2(n17962), .C1(n17961), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17960), .ZN(n17967) );
  NOR2_X1 U21248 ( .A1(n18288), .A2(n9662), .ZN(n17965) );
  NAND2_X1 U21249 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18335), .ZN(
        n18307) );
  NOR2_X1 U21250 ( .A1(n18009), .A2(n18307), .ZN(n18328) );
  NAND3_X1 U21251 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n18328), .ZN(n17974) );
  NAND2_X1 U21252 ( .A1(n18302), .A2(n17974), .ZN(n18293) );
  NOR2_X1 U21253 ( .A1(n18287), .A2(n18152), .ZN(n17964) );
  NOR2_X1 U21254 ( .A1(n18345), .A2(n18307), .ZN(n18327) );
  NAND3_X1 U21255 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n18327), .ZN(n17973) );
  NAND2_X1 U21256 ( .A1(n18302), .A2(n17973), .ZN(n18298) );
  AOI22_X1 U21257 ( .A1(n17965), .A2(n18293), .B1(n17964), .B2(n18298), .ZN(
        n17966) );
  OAI211_X1 U21258 ( .C1(n18044), .C2(n18295), .A(n17967), .B(n17966), .ZN(
        P3_U2815) );
  NOR2_X1 U21259 ( .A1(n17981), .A2(n18307), .ZN(n18310) );
  NOR2_X1 U21260 ( .A1(n17968), .A2(n18009), .ZN(n18023) );
  AOI21_X1 U21261 ( .B1(n18310), .B2(n18023), .A(n17969), .ZN(n17970) );
  XOR2_X1 U21262 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17970), .Z(
        n18320) );
  AND2_X1 U21263 ( .A1(n17985), .A2(n18891), .ZN(n18014) );
  AOI21_X1 U21264 ( .B1(n17984), .B2(n18014), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17971) );
  OAI22_X1 U21265 ( .A1(n17972), .A2(n17971), .B1(n18375), .B2(n19074), .ZN(
        n17976) );
  OAI221_X1 U21266 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18327), .A(n17973), .ZN(
        n18315) );
  OAI221_X1 U21267 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18328), .A(n17974), .ZN(
        n18316) );
  OAI22_X1 U21268 ( .A1(n18152), .A2(n18315), .B1(n9662), .B2(n18316), .ZN(
        n17975) );
  AOI211_X1 U21269 ( .C1(n17977), .C2(n18139), .A(n17976), .B(n17975), .ZN(
        n17978) );
  OAI21_X1 U21270 ( .B1(n18320), .B2(n18044), .A(n17978), .ZN(P3_U2816) );
  OAI22_X1 U21271 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18057), .B1(
        n18307), .B2(n17979), .ZN(n17980) );
  OAI21_X1 U21272 ( .B1(n18057), .B2(n17996), .A(n17980), .ZN(n17982) );
  XNOR2_X1 U21273 ( .A(n17982), .B(n17981), .ZN(n18334) );
  NAND2_X1 U21274 ( .A1(n17985), .A2(n17983), .ZN(n18001) );
  AOI211_X1 U21275 ( .C1(n18000), .C2(n17991), .A(n17984), .B(n18001), .ZN(
        n17993) );
  NOR2_X1 U21276 ( .A1(n17985), .A2(n18105), .ZN(n17986) );
  AOI211_X1 U21277 ( .C1(n17988), .C2(n17987), .A(n18118), .B(n17986), .ZN(
        n17999) );
  OAI22_X1 U21278 ( .A1(n17991), .A2(n17999), .B1(n17990), .B2(n17989), .ZN(
        n17992) );
  AOI211_X1 U21279 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n18408), .A(n17993), 
        .B(n17992), .ZN(n17995) );
  OAI22_X1 U21280 ( .A1(n18328), .A2(n9662), .B1(n18327), .B2(n18152), .ZN(
        n18005) );
  NOR2_X1 U21281 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18307), .ZN(
        n18324) );
  AOI22_X1 U21282 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18005), .B1(
        n18324), .B2(n18041), .ZN(n17994) );
  OAI211_X1 U21283 ( .C1(n18044), .C2(n18334), .A(n17995), .B(n17994), .ZN(
        P3_U2817) );
  AOI21_X1 U21284 ( .B1(n18023), .B2(n18335), .A(n17996), .ZN(n17998) );
  XNOR2_X1 U21285 ( .A(n17998), .B(n17997), .ZN(n18341) );
  NAND2_X1 U21286 ( .A1(n18408), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18339) );
  OAI221_X1 U21287 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18001), .C1(
        n18000), .C2(n17999), .A(n18339), .ZN(n18002) );
  AOI21_X1 U21288 ( .B1(n18004), .B2(n18003), .A(n18002), .ZN(n18007) );
  OAI221_X1 U21289 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18041), 
        .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18335), .A(n18005), .ZN(
        n18006) );
  OAI211_X1 U21290 ( .C1(n18341), .C2(n18044), .A(n18007), .B(n18006), .ZN(
        P3_U2818) );
  AOI22_X1 U21291 ( .A1(n18009), .A2(n18008), .B1(n18136), .B2(n18345), .ZN(
        n18010) );
  INV_X1 U21292 ( .A(n18010), .ZN(n18042) );
  AOI21_X1 U21293 ( .B1(n18350), .B2(n18041), .A(n18042), .ZN(n18029) );
  NAND2_X1 U21294 ( .A1(n18011), .A2(n18891), .ZN(n18085) );
  NOR2_X1 U21295 ( .A1(n18079), .A2(n18085), .ZN(n18077) );
  NAND3_X1 U21296 ( .A1(n18045), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        n18077), .ZN(n18025) );
  NOR2_X1 U21297 ( .A1(n18012), .A2(n18025), .ZN(n18027) );
  AOI21_X1 U21298 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18078), .A(
        n18027), .ZN(n18013) );
  OAI22_X1 U21299 ( .A1(n18014), .A2(n18013), .B1(n18375), .B2(n19067), .ZN(
        n18015) );
  AOI21_X1 U21300 ( .B1(n18016), .B2(n18139), .A(n18015), .ZN(n18020) );
  INV_X1 U21301 ( .A(n18023), .ZN(n18034) );
  OAI21_X1 U21302 ( .B1(n18350), .B2(n18034), .A(n18017), .ZN(n18018) );
  XNOR2_X1 U21303 ( .A(n18018), .B(n18021), .ZN(n18354) );
  NOR2_X1 U21304 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18350), .ZN(
        n18353) );
  AOI22_X1 U21305 ( .A1(n18058), .A2(n18354), .B1(n18353), .B2(n18041), .ZN(
        n18019) );
  OAI211_X1 U21306 ( .C1(n18029), .C2(n18021), .A(n18020), .B(n18019), .ZN(
        P3_U2819) );
  AOI21_X1 U21307 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18023), .A(
        n18022), .ZN(n18024) );
  XNOR2_X1 U21308 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18024), .ZN(
        n18362) );
  AOI21_X1 U21309 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18041), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18028) );
  INV_X1 U21310 ( .A(n18025), .ZN(n18039) );
  AOI21_X1 U21311 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18078), .A(
        n18039), .ZN(n18026) );
  OAI22_X1 U21312 ( .A1(n18029), .A2(n18028), .B1(n18027), .B2(n18026), .ZN(
        n18030) );
  AOI21_X1 U21313 ( .B1(n18058), .B2(n18362), .A(n18030), .ZN(n18031) );
  NAND2_X1 U21314 ( .A1(n18408), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n18365) );
  OAI211_X1 U21315 ( .C1(n18130), .C2(n18032), .A(n18031), .B(n18365), .ZN(
        P3_U2820) );
  NAND2_X1 U21316 ( .A1(n18034), .A2(n18033), .ZN(n18035) );
  XNOR2_X1 U21317 ( .A(n18035), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n18381) );
  INV_X1 U21318 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18368) );
  AOI22_X1 U21319 ( .A1(n18045), .A2(n18077), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18078), .ZN(n18038) );
  AOI22_X1 U21320 ( .A1(n18435), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18036), 
        .B2(n18139), .ZN(n18037) );
  OAI21_X1 U21321 ( .B1(n18039), .B2(n18038), .A(n18037), .ZN(n18040) );
  AOI221_X1 U21322 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18042), .C1(
        n18368), .C2(n18041), .A(n18040), .ZN(n18043) );
  OAI21_X1 U21323 ( .B1(n18381), .B2(n18044), .A(n18043), .ZN(P3_U2821) );
  AOI211_X1 U21324 ( .C1(n18049), .C2(n18046), .A(n18045), .B(n18717), .ZN(
        n18052) );
  AOI21_X1 U21325 ( .B1(n18048), .B2(n18047), .A(n18118), .ZN(n18064) );
  OAI22_X1 U21326 ( .A1(n18130), .A2(n18050), .B1(n18049), .B2(n18064), .ZN(
        n18051) );
  AOI211_X1 U21327 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n18435), .A(n18052), .B(
        n18051), .ZN(n18060) );
  AOI21_X1 U21328 ( .B1(n18054), .B2(n18370), .A(n18053), .ZN(n18392) );
  OAI21_X1 U21329 ( .B1(n18057), .B2(n18056), .A(n18055), .ZN(n18390) );
  AOI22_X1 U21330 ( .A1(n18136), .A2(n18392), .B1(n18058), .B2(n18390), .ZN(
        n18059) );
  OAI211_X1 U21331 ( .C1(n9662), .C2(n18396), .A(n18060), .B(n18059), .ZN(
        P3_U2822) );
  NAND2_X1 U21332 ( .A1(n18062), .A2(n18061), .ZN(n18063) );
  XNOR2_X1 U21333 ( .A(n18063), .B(n18400), .ZN(n18406) );
  INV_X1 U21334 ( .A(n18064), .ZN(n18066) );
  NOR2_X1 U21335 ( .A1(n18375), .A2(n19059), .ZN(n18397) );
  AOI221_X1 U21336 ( .B1(n18066), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n18077), .C2(n18065), .A(n18397), .ZN(n18071) );
  AOI21_X1 U21337 ( .B1(n18400), .B2(n18068), .A(n18067), .ZN(n18403) );
  AOI22_X1 U21338 ( .A1(n18140), .A2(n18403), .B1(n18069), .B2(n18139), .ZN(
        n18070) );
  OAI211_X1 U21339 ( .C1(n18152), .C2(n18406), .A(n18071), .B(n18070), .ZN(
        P3_U2823) );
  AOI21_X1 U21340 ( .B1(n18074), .B2(n18073), .A(n18072), .ZN(n18410) );
  AOI22_X1 U21341 ( .A1(n18140), .A2(n18410), .B1(n18369), .B2(
        P3_REIP_REG_6__SCAN_IN), .ZN(n18083) );
  AOI21_X1 U21342 ( .B1(n18076), .B2(n18399), .A(n18075), .ZN(n18409) );
  INV_X1 U21343 ( .A(n18077), .ZN(n18081) );
  INV_X1 U21344 ( .A(n18078), .ZN(n18144) );
  OAI21_X1 U21345 ( .B1(n18144), .B2(n18079), .A(n18085), .ZN(n18080) );
  AOI22_X1 U21346 ( .A1(n18136), .A2(n18409), .B1(n18081), .B2(n18080), .ZN(
        n18082) );
  OAI211_X1 U21347 ( .C1(n18130), .C2(n18084), .A(n18083), .B(n18082), .ZN(
        P3_U2824) );
  OAI221_X1 U21348 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18086), .C1(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n18147), .A(n18085), .ZN(n18097) );
  OAI21_X1 U21349 ( .B1(n18089), .B2(n18088), .A(n18087), .ZN(n18090) );
  XNOR2_X1 U21350 ( .A(n18090), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18414) );
  AOI22_X1 U21351 ( .A1(n18140), .A2(n18414), .B1(n18369), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n18096) );
  AOI21_X1 U21352 ( .B1(n18093), .B2(n18092), .A(n18091), .ZN(n18415) );
  AOI22_X1 U21353 ( .A1(n18136), .A2(n18415), .B1(n18094), .B2(n18139), .ZN(
        n18095) );
  OAI211_X1 U21354 ( .C1(n18144), .C2(n18097), .A(n18096), .B(n18095), .ZN(
        P3_U2825) );
  AOI21_X1 U21355 ( .B1(n18432), .B2(n18099), .A(n18098), .ZN(n18429) );
  OAI22_X1 U21356 ( .A1(n18375), .A2(n19053), .B1(n18717), .B2(n18100), .ZN(
        n18101) );
  AOI21_X1 U21357 ( .B1(n18136), .B2(n18429), .A(n18101), .ZN(n18108) );
  AOI21_X1 U21358 ( .B1(n18104), .B2(n18103), .A(n18102), .ZN(n18425) );
  OAI21_X1 U21359 ( .B1(n18106), .B2(n18105), .A(n18147), .ZN(n18120) );
  AOI22_X1 U21360 ( .A1(n18140), .A2(n18425), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18120), .ZN(n18107) );
  OAI211_X1 U21361 ( .C1(n18130), .C2(n18109), .A(n18108), .B(n18107), .ZN(
        P3_U2826) );
  OAI21_X1 U21362 ( .B1(n18112), .B2(n18111), .A(n18110), .ZN(n18113) );
  XNOR2_X1 U21363 ( .A(n18113), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n18434) );
  AOI22_X1 U21364 ( .A1(n18140), .A2(n18434), .B1(n18369), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n18122) );
  AOI21_X1 U21365 ( .B1(n18116), .B2(n18115), .A(n18114), .ZN(n18436) );
  OAI21_X1 U21366 ( .B1(n18118), .B2(n18133), .A(n18117), .ZN(n18119) );
  AOI22_X1 U21367 ( .A1(n18136), .A2(n18436), .B1(n18120), .B2(n18119), .ZN(
        n18121) );
  OAI211_X1 U21368 ( .C1(n18130), .C2(n18123), .A(n18122), .B(n18121), .ZN(
        P3_U2827) );
  AOI21_X1 U21369 ( .B1(n18126), .B2(n18125), .A(n18124), .ZN(n18453) );
  NOR2_X1 U21370 ( .A1(n18375), .A2(n19049), .ZN(n18442) );
  XNOR2_X1 U21371 ( .A(n18128), .B(n18127), .ZN(n18457) );
  OAI22_X1 U21372 ( .A1(n18130), .A2(n18129), .B1(n18151), .B2(n18457), .ZN(
        n18131) );
  AOI211_X1 U21373 ( .C1(n18136), .C2(n18453), .A(n18442), .B(n18131), .ZN(
        n18132) );
  OAI221_X1 U21374 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18717), .C1(
        n18133), .C2(n18147), .A(n18132), .ZN(P3_U2828) );
  NOR2_X1 U21375 ( .A1(n18146), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18134) );
  XOR2_X1 U21376 ( .A(n18134), .B(n18138), .Z(n18469) );
  INV_X1 U21377 ( .A(n18469), .ZN(n18135) );
  AOI22_X1 U21378 ( .A1(n18136), .A2(n18135), .B1(n18369), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18142) );
  AOI21_X1 U21379 ( .B1(n18138), .B2(n18145), .A(n18137), .ZN(n18464) );
  AOI22_X1 U21380 ( .A1(n18140), .A2(n18464), .B1(n18143), .B2(n18139), .ZN(
        n18141) );
  OAI211_X1 U21381 ( .C1(n18144), .C2(n18143), .A(n18142), .B(n18141), .ZN(
        P3_U2829) );
  OAI21_X1 U21382 ( .B1(n18146), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18145), .ZN(n18475) );
  INV_X1 U21383 ( .A(n18475), .ZN(n18473) );
  NAND3_X1 U21384 ( .A1(n19134), .A2(n18148), .A3(n18147), .ZN(n18149) );
  AOI22_X1 U21385 ( .A1(n18435), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18149), .ZN(n18150) );
  OAI221_X1 U21386 ( .B1(n18473), .B2(n18152), .C1(n18475), .C2(n18151), .A(
        n18150), .ZN(P3_U2830) );
  INV_X1 U21387 ( .A(n18153), .ZN(n18154) );
  NOR2_X1 U21388 ( .A1(n18229), .A2(n18154), .ZN(n18167) );
  NOR2_X1 U21389 ( .A1(n18155), .A2(n18326), .ZN(n18164) );
  NOR2_X1 U21390 ( .A1(n18972), .A2(n18306), .ZN(n18445) );
  INV_X1 U21391 ( .A(n18445), .ZN(n18421) );
  OAI21_X1 U21392 ( .B1(n18157), .B2(n18306), .A(n18156), .ZN(n18222) );
  OAI21_X1 U21393 ( .B1(n18158), .B2(n18259), .A(n18972), .ZN(n18159) );
  OAI21_X1 U21394 ( .B1(n18445), .B2(n18222), .A(n18159), .ZN(n18195) );
  AOI21_X1 U21395 ( .B1(n18160), .B2(n18421), .A(n18195), .ZN(n18184) );
  OAI211_X1 U21396 ( .C1(n18162), .C2(n18445), .A(n18161), .B(n18184), .ZN(
        n18163) );
  AOI211_X1 U21397 ( .C1(n18217), .C2(n18165), .A(n18164), .B(n18163), .ZN(
        n18172) );
  INV_X1 U21398 ( .A(n18172), .ZN(n18166) );
  MUX2_X1 U21399 ( .A(n18167), .B(n18166), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n18168) );
  AOI22_X1 U21400 ( .A1(n18391), .A2(n18169), .B1(n18168), .B2(n18375), .ZN(
        n18171) );
  NAND2_X1 U21401 ( .A1(n18171), .A2(n18170), .ZN(P3_U2835) );
  NOR2_X1 U21402 ( .A1(n18369), .A2(n18172), .ZN(n18174) );
  AOI22_X1 U21403 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18174), .B1(
        n18204), .B2(n18173), .ZN(n18176) );
  NAND2_X1 U21404 ( .A1(n18408), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18175) );
  OAI211_X1 U21405 ( .C1(n18177), .C2(n18380), .A(n18176), .B(n18175), .ZN(
        P3_U2836) );
  OAI221_X1 U21406 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18179), 
        .C1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n18178), .A(n18471), .ZN(
        n18185) );
  NOR2_X1 U21407 ( .A1(n18181), .A2(n18180), .ZN(n18183) );
  OAI221_X1 U21408 ( .B1(n18185), .B2(n18184), .C1(n18185), .C2(n18183), .A(
        n18182), .ZN(n18189) );
  INV_X1 U21409 ( .A(n18322), .ZN(n18395) );
  OAI22_X1 U21410 ( .A1(n18395), .A2(n18187), .B1(n18380), .B2(n18186), .ZN(
        n18188) );
  AOI211_X1 U21411 ( .C1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n18470), .A(
        n18189), .B(n18188), .ZN(n18190) );
  OAI21_X1 U21412 ( .B1(n18468), .B2(n18191), .A(n18190), .ZN(P3_U2837) );
  INV_X1 U21413 ( .A(n18217), .ZN(n18347) );
  OAI22_X1 U21414 ( .A1(n18193), .A2(n18347), .B1(n18192), .B2(n18326), .ZN(
        n18194) );
  NOR3_X1 U21415 ( .A1(n18470), .A2(n18195), .A3(n18194), .ZN(n18201) );
  NAND3_X1 U21416 ( .A1(n18261), .A2(n18196), .A3(n18257), .ZN(n18198) );
  AOI21_X1 U21417 ( .B1(n18964), .B2(n18198), .A(n18197), .ZN(n18199) );
  AOI21_X1 U21418 ( .B1(n18201), .B2(n18199), .A(n18369), .ZN(n18209) );
  AOI21_X1 U21419 ( .B1(n18385), .B2(n18201), .A(n18200), .ZN(n18202) );
  AOI22_X1 U21420 ( .A1(n18204), .A2(n18203), .B1(n18209), .B2(n18202), .ZN(
        n18206) );
  NAND2_X1 U21421 ( .A1(n18408), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18205) );
  OAI211_X1 U21422 ( .C1(n18207), .C2(n18380), .A(n18206), .B(n18205), .ZN(
        P3_U2838) );
  NOR2_X1 U21423 ( .A1(n18470), .A2(n18208), .ZN(n18210) );
  OAI21_X1 U21424 ( .B1(n18210), .B2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n18209), .ZN(n18211) );
  OAI211_X1 U21425 ( .C1(n18213), .C2(n18380), .A(n18212), .B(n18211), .ZN(
        P3_U2839) );
  AOI22_X1 U21426 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18470), .B1(
        n18369), .B2(P3_REIP_REG_22__SCAN_IN), .ZN(n18227) );
  INV_X1 U21427 ( .A(n18259), .ZN(n18216) );
  OAI22_X1 U21428 ( .A1(n18287), .A2(n18326), .B1(n18288), .B2(n18347), .ZN(
        n18258) );
  AOI221_X1 U21429 ( .B1(n18214), .B2(n18964), .C1(n18231), .C2(n18964), .A(
        n18258), .ZN(n18215) );
  OAI221_X1 U21430 ( .B1(n18990), .B2(n18216), .C1(n18990), .C2(n18243), .A(
        n18215), .ZN(n18240) );
  NOR2_X1 U21431 ( .A1(n18953), .A2(n18217), .ZN(n18342) );
  OAI22_X1 U21432 ( .A1(n18990), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n18218), .B2(n18342), .ZN(n18219) );
  NOR2_X1 U21433 ( .A1(n18240), .A2(n18219), .ZN(n18233) );
  AOI22_X1 U21434 ( .A1(n18964), .A2(n18221), .B1(n18277), .B2(n18220), .ZN(
        n18223) );
  NAND3_X1 U21435 ( .A1(n18233), .A2(n18223), .A3(n18222), .ZN(n18224) );
  OAI211_X1 U21436 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n18225), .A(
        n18471), .B(n18224), .ZN(n18226) );
  OAI211_X1 U21437 ( .C1(n18228), .C2(n18380), .A(n18227), .B(n18226), .ZN(
        P3_U2840) );
  NOR3_X1 U21438 ( .A1(n18229), .A2(n18460), .A3(n18231), .ZN(n18249) );
  AOI22_X1 U21439 ( .A1(n18435), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18230), 
        .B2(n18249), .ZN(n18237) );
  INV_X1 U21440 ( .A(n18231), .ZN(n18232) );
  OAI221_X1 U21441 ( .B1(n18988), .B2(n18279), .C1(n18988), .C2(n18232), .A(
        n18471), .ZN(n18241) );
  NOR2_X1 U21442 ( .A1(n18964), .A2(n18306), .ZN(n18459) );
  OAI21_X1 U21443 ( .B1(n18234), .B2(n18459), .A(n18233), .ZN(n18235) );
  OAI211_X1 U21444 ( .C1(n18241), .C2(n18235), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18375), .ZN(n18236) );
  OAI211_X1 U21445 ( .C1(n18238), .C2(n18380), .A(n18237), .B(n18236), .ZN(
        P3_U2841) );
  AOI22_X1 U21446 ( .A1(n18435), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18249), 
        .B2(n18239), .ZN(n18246) );
  NOR2_X1 U21447 ( .A1(n18241), .A2(n18240), .ZN(n18242) );
  AOI221_X1 U21448 ( .B1(n18243), .B2(n18242), .C1(n18342), .C2(n18242), .A(
        n18408), .ZN(n18250) );
  NOR3_X1 U21449 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18459), .A3(
        n19183), .ZN(n18244) );
  OAI21_X1 U21450 ( .B1(n18250), .B2(n18244), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18245) );
  OAI211_X1 U21451 ( .C1(n18247), .C2(n18380), .A(n18246), .B(n18245), .ZN(
        P3_U2842) );
  AOI22_X1 U21452 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18250), .B1(
        n18249), .B2(n18248), .ZN(n18252) );
  NAND2_X1 U21453 ( .A1(n18408), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18251) );
  OAI211_X1 U21454 ( .C1(n18253), .C2(n18380), .A(n18252), .B(n18251), .ZN(
        P3_U2843) );
  INV_X1 U21455 ( .A(n18424), .ZN(n18448) );
  INV_X1 U21456 ( .A(n18254), .ZN(n18422) );
  OAI22_X1 U21457 ( .A1(n18448), .A2(n18983), .B1(n18422), .B2(n18452), .ZN(
        n18438) );
  NAND2_X1 U21458 ( .A1(n18471), .A2(n18438), .ZN(n18426) );
  INV_X1 U21459 ( .A(n18426), .ZN(n18417) );
  AOI22_X1 U21460 ( .A1(n18256), .A2(n18321), .B1(n18471), .B2(n18255), .ZN(
        n18286) );
  NAND2_X1 U21461 ( .A1(n18261), .A2(n18257), .ZN(n18263) );
  OR2_X1 U21462 ( .A1(n18460), .A2(n18258), .ZN(n18281) );
  NOR2_X1 U21463 ( .A1(n18988), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18447) );
  NOR3_X1 U21464 ( .A1(n18447), .A2(n18259), .A3(n18285), .ZN(n18260) );
  OAI22_X1 U21465 ( .A1(n18261), .A2(n18342), .B1(n18445), .B2(n18260), .ZN(
        n18262) );
  AOI211_X1 U21466 ( .C1(n18964), .C2(n18263), .A(n18281), .B(n18262), .ZN(
        n18270) );
  AOI221_X1 U21467 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18270), 
        .C1(n18445), .C2(n18270), .A(n18435), .ZN(n18265) );
  AOI22_X1 U21468 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18265), .B1(
        n18391), .B2(n18264), .ZN(n18267) );
  NAND2_X1 U21469 ( .A1(n18408), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18266) );
  OAI211_X1 U21470 ( .C1(n18286), .C2(n18268), .A(n18267), .B(n18266), .ZN(
        P3_U2844) );
  NOR3_X1 U21471 ( .A1(n18435), .A2(n18270), .A3(n18269), .ZN(n18271) );
  AOI21_X1 U21472 ( .B1(n18391), .B2(n18272), .A(n18271), .ZN(n18274) );
  OAI211_X1 U21473 ( .C1(n18286), .C2(n18275), .A(n18274), .B(n18273), .ZN(
        P3_U2845) );
  AND2_X1 U21474 ( .A1(n18303), .A2(n18964), .ZN(n18344) );
  OAI21_X1 U21475 ( .B1(n18370), .B2(n18371), .A(n18972), .ZN(n18358) );
  INV_X1 U21476 ( .A(n18358), .ZN(n18276) );
  AOI211_X1 U21477 ( .C1(n18277), .C2(n18290), .A(n18344), .B(n18276), .ZN(
        n18278) );
  OAI211_X1 U21478 ( .C1(n18279), .C2(n18988), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18278), .ZN(n18292) );
  OAI221_X1 U21479 ( .B1(n18281), .B2(n18280), .C1(n18281), .C2(n18292), .A(
        n18375), .ZN(n18284) );
  AOI22_X1 U21480 ( .A1(n18435), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18391), 
        .B2(n18282), .ZN(n18283) );
  OAI221_X1 U21481 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18286), 
        .C1(n18285), .C2(n18284), .A(n18283), .ZN(P3_U2846) );
  INV_X1 U21482 ( .A(n18470), .ZN(n18461) );
  NOR2_X1 U21483 ( .A1(n18287), .A2(n18468), .ZN(n18299) );
  NOR2_X1 U21484 ( .A1(n18288), .A2(n18347), .ZN(n18294) );
  NAND2_X1 U21485 ( .A1(n18311), .A2(n18438), .ZN(n18289) );
  OAI21_X1 U21486 ( .B1(n18290), .B2(n18289), .A(n18302), .ZN(n18291) );
  AOI22_X1 U21487 ( .A1(n18294), .A2(n18293), .B1(n18292), .B2(n18291), .ZN(
        n18296) );
  OAI22_X1 U21488 ( .A1(n18296), .A2(n18460), .B1(n18380), .B2(n18295), .ZN(
        n18297) );
  AOI21_X1 U21489 ( .B1(n18299), .B2(n18298), .A(n18297), .ZN(n18301) );
  NAND2_X1 U21490 ( .A1(n18408), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18300) );
  OAI211_X1 U21491 ( .C1(n18461), .C2(n18302), .A(n18301), .B(n18300), .ZN(
        P3_U2847) );
  OAI21_X1 U21492 ( .B1(n18303), .B2(n18307), .A(n18964), .ZN(n18304) );
  OAI211_X1 U21493 ( .C1(n18990), .C2(n18310), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18304), .ZN(n18309) );
  NAND2_X1 U21494 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18305), .ZN(
        n18343) );
  OAI21_X1 U21495 ( .B1(n18307), .B2(n18343), .A(n18306), .ZN(n18325) );
  OAI211_X1 U21496 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18459), .A(
        n18358), .B(n18325), .ZN(n18308) );
  OAI21_X1 U21497 ( .B1(n18309), .B2(n18308), .A(n18471), .ZN(n18313) );
  NAND3_X1 U21498 ( .A1(n18311), .A2(n18310), .A3(n18438), .ZN(n18312) );
  AOI222_X1 U21499 ( .A1(n18314), .A2(n18313), .B1(n18314), .B2(n18312), .C1(
        n18313), .C2(n18461), .ZN(n18318) );
  OAI22_X1 U21500 ( .A1(n18395), .A2(n18316), .B1(n18468), .B2(n18315), .ZN(
        n18317) );
  AOI211_X1 U21501 ( .C1(n18435), .C2(P3_REIP_REG_14__SCAN_IN), .A(n18318), 
        .B(n18317), .ZN(n18319) );
  OAI21_X1 U21502 ( .B1(n18320), .B2(n18380), .A(n18319), .ZN(P3_U2848) );
  AOI21_X1 U21503 ( .B1(n18322), .B2(n13224), .A(n18321), .ZN(n18323) );
  OAI21_X1 U21504 ( .B1(n18345), .B2(n18468), .A(n18323), .ZN(n18367) );
  AOI22_X1 U21505 ( .A1(n18435), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18324), 
        .B2(n18367), .ZN(n18333) );
  INV_X1 U21506 ( .A(n18325), .ZN(n18330) );
  OAI21_X1 U21507 ( .B1(n18359), .B2(n18335), .A(n18358), .ZN(n18352) );
  OAI22_X1 U21508 ( .A1(n18328), .A2(n18347), .B1(n18327), .B2(n18326), .ZN(
        n18329) );
  NOR4_X1 U21509 ( .A1(n18344), .A2(n18330), .A3(n18352), .A4(n18329), .ZN(
        n18337) );
  OAI211_X1 U21510 ( .C1(n18359), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18471), .B(n18337), .ZN(n18331) );
  NAND3_X1 U21511 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18375), .A3(
        n18331), .ZN(n18332) );
  OAI211_X1 U21512 ( .C1(n18334), .C2(n18380), .A(n18333), .B(n18332), .ZN(
        P3_U2849) );
  AOI22_X1 U21513 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18471), .B1(
        n18335), .B2(n18367), .ZN(n18336) );
  AOI21_X1 U21514 ( .B1(n18337), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18336), .ZN(n18338) );
  AOI21_X1 U21515 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18470), .A(
        n18338), .ZN(n18340) );
  OAI211_X1 U21516 ( .C1(n18341), .C2(n18380), .A(n18340), .B(n18339), .ZN(
        P3_U2850) );
  INV_X1 U21517 ( .A(n18342), .ZN(n18349) );
  INV_X1 U21518 ( .A(n18343), .ZN(n18374) );
  AOI21_X1 U21519 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18374), .A(
        n18988), .ZN(n18348) );
  AOI211_X1 U21520 ( .C1(n18345), .C2(n18953), .A(n18344), .B(n18460), .ZN(
        n18346) );
  OAI21_X1 U21521 ( .B1(n13224), .B2(n18347), .A(n18346), .ZN(n18377) );
  AOI211_X1 U21522 ( .C1(n18350), .C2(n18349), .A(n18348), .B(n18377), .ZN(
        n18357) );
  OAI21_X1 U21523 ( .B1(n18988), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18357), .ZN(n18351) );
  OAI21_X1 U21524 ( .B1(n18352), .B2(n18351), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18356) );
  AOI22_X1 U21525 ( .A1(n18391), .A2(n18354), .B1(n18353), .B2(n18367), .ZN(
        n18355) );
  OAI221_X1 U21526 ( .B1(n18435), .B2(n18356), .C1(n18375), .C2(n19067), .A(
        n18355), .ZN(P3_U2851) );
  NOR2_X1 U21527 ( .A1(n18369), .A2(n18363), .ZN(n18361) );
  OAI211_X1 U21528 ( .C1(n18359), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18358), .B(n18357), .ZN(n18360) );
  AOI22_X1 U21529 ( .A1(n18391), .A2(n18362), .B1(n18361), .B2(n18360), .ZN(
        n18366) );
  NAND3_X1 U21530 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18363), .A3(
        n18367), .ZN(n18364) );
  NAND3_X1 U21531 ( .A1(n18366), .A2(n18365), .A3(n18364), .ZN(P3_U2852) );
  AOI22_X1 U21532 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n18369), .B1(n18368), 
        .B2(n18367), .ZN(n18379) );
  NAND2_X1 U21533 ( .A1(n18972), .A2(n18370), .ZN(n18373) );
  NAND2_X1 U21534 ( .A1(n18972), .A2(n18371), .ZN(n18372) );
  OAI211_X1 U21535 ( .C1(n18374), .C2(n18988), .A(n18373), .B(n18372), .ZN(
        n18376) );
  OAI211_X1 U21536 ( .C1(n18377), .C2(n18376), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n18375), .ZN(n18378) );
  OAI211_X1 U21537 ( .C1(n18381), .C2(n18380), .A(n18379), .B(n18378), .ZN(
        P3_U2853) );
  NOR2_X1 U21538 ( .A1(n18382), .A2(n18426), .ZN(n18388) );
  AOI21_X1 U21539 ( .B1(n18398), .B2(n18424), .A(n18983), .ZN(n18383) );
  AOI211_X1 U21540 ( .C1(n18384), .C2(n18421), .A(n18383), .B(n18447), .ZN(
        n18407) );
  OAI211_X1 U21541 ( .C1(n18385), .C2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n18407), .ZN(n18402) );
  AOI21_X1 U21542 ( .B1(n18465), .B2(n18402), .A(n18470), .ZN(n18386) );
  INV_X1 U21543 ( .A(n18386), .ZN(n18387) );
  MUX2_X1 U21544 ( .A(n18388), .B(n18387), .S(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .Z(n18389) );
  AOI21_X1 U21545 ( .B1(n18408), .B2(P3_REIP_REG_8__SCAN_IN), .A(n18389), .ZN(
        n18394) );
  AOI22_X1 U21546 ( .A1(n18476), .A2(n18392), .B1(n18391), .B2(n18390), .ZN(
        n18393) );
  OAI211_X1 U21547 ( .C1(n18396), .C2(n18395), .A(n18394), .B(n18393), .ZN(
        P3_U2854) );
  AOI21_X1 U21548 ( .B1(n18470), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18397), .ZN(n18405) );
  NAND2_X1 U21549 ( .A1(n18398), .A2(n18417), .ZN(n18413) );
  OAI22_X1 U21550 ( .A1(n18400), .A2(n18460), .B1(n18399), .B2(n18413), .ZN(
        n18401) );
  AOI22_X1 U21551 ( .A1(n18474), .A2(n18403), .B1(n18402), .B2(n18401), .ZN(
        n18404) );
  OAI211_X1 U21552 ( .C1(n18468), .C2(n18406), .A(n18405), .B(n18404), .ZN(
        P3_U2855) );
  OAI21_X1 U21553 ( .B1(n18407), .B2(n18460), .A(n18461), .ZN(n18416) );
  AOI22_X1 U21554 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18416), .B1(
        n18408), .B2(P3_REIP_REG_6__SCAN_IN), .ZN(n18412) );
  AOI22_X1 U21555 ( .A1(n18474), .A2(n18410), .B1(n18476), .B2(n18409), .ZN(
        n18411) );
  OAI211_X1 U21556 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n18413), .A(
        n18412), .B(n18411), .ZN(P3_U2856) );
  AOI22_X1 U21557 ( .A1(n18435), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18474), 
        .B2(n18414), .ZN(n18420) );
  AOI22_X1 U21558 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18416), .B1(
        n18476), .B2(n18415), .ZN(n18419) );
  NAND4_X1 U21559 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n18417), .A4(n13040), .ZN(
        n18418) );
  NAND3_X1 U21560 ( .A1(n18420), .A2(n18419), .A3(n18418), .ZN(P3_U2857) );
  AOI211_X1 U21561 ( .C1(n18422), .C2(n18421), .A(n18447), .B(n18427), .ZN(
        n18423) );
  OAI21_X1 U21562 ( .B1(n18983), .B2(n18424), .A(n18423), .ZN(n18437) );
  AOI21_X1 U21563 ( .B1(n18465), .B2(n18437), .A(n18470), .ZN(n18433) );
  AOI22_X1 U21564 ( .A1(n18435), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18474), 
        .B2(n18425), .ZN(n18431) );
  NOR2_X1 U21565 ( .A1(n18427), .A2(n18426), .ZN(n18428) );
  AOI22_X1 U21566 ( .A1(n18429), .A2(n18476), .B1(n18428), .B2(n18432), .ZN(
        n18430) );
  OAI211_X1 U21567 ( .C1(n18433), .C2(n18432), .A(n18431), .B(n18430), .ZN(
        P3_U2858) );
  AOI22_X1 U21568 ( .A1(n18435), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18474), 
        .B2(n18434), .ZN(n18441) );
  AOI22_X1 U21569 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18470), .B1(
        n18476), .B2(n18436), .ZN(n18440) );
  OAI211_X1 U21570 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18438), .A(
        n18471), .B(n18437), .ZN(n18439) );
  NAND3_X1 U21571 ( .A1(n18441), .A2(n18440), .A3(n18439), .ZN(P3_U2859) );
  AOI21_X1 U21572 ( .B1(n18470), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n18442), .ZN(n18456) );
  NAND2_X1 U21573 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18443), .ZN(
        n18451) );
  NAND2_X1 U21574 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18444) );
  OAI22_X1 U21575 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18445), .B1(
        n18983), .B2(n18444), .ZN(n18446) );
  OAI21_X1 U21576 ( .B1(n18447), .B2(n18446), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18450) );
  NAND2_X1 U21577 ( .A1(n18964), .A2(n18448), .ZN(n18449) );
  OAI211_X1 U21578 ( .C1(n18452), .C2(n18451), .A(n18450), .B(n18449), .ZN(
        n18454) );
  AOI22_X1 U21579 ( .A1(n18471), .A2(n18454), .B1(n18476), .B2(n18453), .ZN(
        n18455) );
  OAI211_X1 U21580 ( .C1(n18458), .C2(n18457), .A(n18456), .B(n18455), .ZN(
        P3_U2860) );
  NOR2_X1 U21581 ( .A1(n18375), .A2(n19153), .ZN(n18463) );
  OR3_X1 U21582 ( .A1(n18460), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n18459), .ZN(n18477) );
  AOI21_X1 U21583 ( .B1(n18461), .B2(n18477), .A(n13031), .ZN(n18462) );
  AOI211_X1 U21584 ( .C1(n18464), .C2(n18474), .A(n18463), .B(n18462), .ZN(
        n18467) );
  OAI211_X1 U21585 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18972), .A(
        n18465), .B(n13031), .ZN(n18466) );
  OAI211_X1 U21586 ( .C1(n18469), .C2(n18468), .A(n18467), .B(n18466), .ZN(
        P3_U2861) );
  AOI21_X1 U21587 ( .B1(n18471), .B2(n18972), .A(n18470), .ZN(n18479) );
  INV_X1 U21588 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n19159) );
  NOR2_X1 U21589 ( .A1(n18375), .A2(n19159), .ZN(n18472) );
  AOI221_X1 U21590 ( .B1(n18476), .B2(n18475), .C1(n18474), .C2(n18473), .A(
        n18472), .ZN(n18478) );
  OAI211_X1 U21591 ( .C1(n18479), .C2(n19149), .A(n18478), .B(n18477), .ZN(
        P3_U2862) );
  AOI211_X1 U21592 ( .C1(n18481), .C2(n18480), .A(n19183), .B(n19134), .ZN(
        n19015) );
  OAI21_X1 U21593 ( .B1(n19015), .B2(n18538), .A(n18486), .ZN(n18482) );
  OAI221_X1 U21594 ( .B1(n18487), .B2(n19168), .C1(n18487), .C2(n18486), .A(
        n18482), .ZN(P3_U2863) );
  NOR2_X1 U21595 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19004), .ZN(
        n18771) );
  NOR2_X1 U21596 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19001), .ZN(
        n18668) );
  NOR2_X1 U21597 ( .A1(n18771), .A2(n18668), .ZN(n18484) );
  OAI22_X1 U21598 ( .A1(n18485), .A2(n19004), .B1(n18484), .B2(n18483), .ZN(
        P3_U2866) );
  NOR2_X1 U21599 ( .A1(n19005), .A2(n18486), .ZN(P3_U2867) );
  NAND2_X1 U21600 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18995) );
  NOR2_X1 U21601 ( .A1(n19001), .A2(n19004), .ZN(n18488) );
  INV_X1 U21602 ( .A(n18488), .ZN(n18489) );
  OR2_X1 U21603 ( .A1(n18995), .A2(n18489), .ZN(n18940) );
  INV_X1 U21604 ( .A(n18940), .ZN(n18946) );
  NAND2_X1 U21605 ( .A1(n18996), .A2(n18487), .ZN(n18997) );
  NAND2_X1 U21606 ( .A1(n19001), .A2(n19004), .ZN(n18621) );
  NOR2_X1 U21607 ( .A1(n18997), .A2(n18621), .ZN(n18581) );
  NOR2_X1 U21608 ( .A1(n18946), .A2(n18594), .ZN(n18557) );
  OAI21_X1 U21609 ( .B1(n18487), .B2(n19125), .A(n18857), .ZN(n18746) );
  NAND2_X1 U21610 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18487), .ZN(
        n18644) );
  NAND2_X1 U21611 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18996), .ZN(
        n18719) );
  NAND2_X1 U21612 ( .A1(n18644), .A2(n18719), .ZN(n18796) );
  NAND2_X1 U21613 ( .A1(n18488), .A2(n18796), .ZN(n18854) );
  OAI22_X1 U21614 ( .A1(n18557), .A2(n18746), .B1(n18717), .B2(n18854), .ZN(
        n18536) );
  NAND2_X1 U21615 ( .A1(n18488), .A2(n18996), .ZN(n18827) );
  INV_X1 U21616 ( .A(n18827), .ZN(n18890) );
  NAND2_X1 U21617 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18890), .ZN(
        n18952) );
  INV_X1 U21618 ( .A(n18952), .ZN(n18937) );
  NAND2_X1 U21619 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18891), .ZN(n18861) );
  INV_X1 U21620 ( .A(n18861), .ZN(n18895) );
  AND2_X1 U21621 ( .A1(n18857), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18894) );
  NOR2_X1 U21622 ( .A1(n19023), .A2(n18557), .ZN(n18530) );
  AOI22_X1 U21623 ( .A1(n18937), .A2(n18895), .B1(n18894), .B2(n18530), .ZN(
        n18495) );
  NOR2_X1 U21624 ( .A1(n18489), .A2(n18644), .ZN(n18884) );
  AND2_X1 U21625 ( .A1(n18891), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18897) );
  INV_X1 U21626 ( .A(n18490), .ZN(n18491) );
  NAND2_X1 U21627 ( .A1(n18492), .A2(n18491), .ZN(n18532) );
  NOR2_X2 U21628 ( .A1(n18493), .A2(n18532), .ZN(n18896) );
  AOI22_X1 U21629 ( .A1(n18877), .A2(n18897), .B1(n18896), .B2(n18594), .ZN(
        n18494) );
  OAI211_X1 U21630 ( .C1(n18496), .C2(n18536), .A(n18495), .B(n18494), .ZN(
        P3_U2868) );
  NAND2_X1 U21631 ( .A1(n18891), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18906) );
  AND2_X1 U21632 ( .A1(n18857), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18901) );
  AOI22_X1 U21633 ( .A1(n18884), .A2(n18803), .B1(n18901), .B2(n18530), .ZN(
        n18500) );
  NOR2_X2 U21634 ( .A1(n18497), .A2(n18717), .ZN(n18902) );
  NOR2_X1 U21635 ( .A1(n18498), .A2(n18532), .ZN(n18903) );
  AOI22_X1 U21636 ( .A1(n18937), .A2(n18902), .B1(n18903), .B2(n18594), .ZN(
        n18499) );
  OAI211_X1 U21637 ( .C1(n18501), .C2(n18536), .A(n18500), .B(n18499), .ZN(
        P3_U2869) );
  AND2_X1 U21638 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18891), .ZN(n18908) );
  INV_X1 U21639 ( .A(n18857), .ZN(n18798) );
  NOR2_X2 U21640 ( .A1(n18798), .A2(n18502), .ZN(n18907) );
  AOI22_X1 U21641 ( .A1(n18937), .A2(n18908), .B1(n18907), .B2(n18530), .ZN(
        n18505) );
  NAND2_X1 U21642 ( .A1(n18891), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18912) );
  INV_X1 U21643 ( .A(n18912), .ZN(n18833) );
  NOR2_X1 U21644 ( .A1(n18503), .A2(n18532), .ZN(n18909) );
  AOI22_X1 U21645 ( .A1(n18877), .A2(n18833), .B1(n18909), .B2(n18594), .ZN(
        n18504) );
  OAI211_X1 U21646 ( .C1(n18506), .C2(n18536), .A(n18505), .B(n18504), .ZN(
        P3_U2870) );
  NAND2_X1 U21647 ( .A1(n18891), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18868) );
  INV_X1 U21648 ( .A(n18868), .ZN(n18916) );
  NOR2_X2 U21649 ( .A1(n18798), .A2(n18507), .ZN(n18913) );
  AOI22_X1 U21650 ( .A1(n18884), .A2(n18916), .B1(n18913), .B2(n18530), .ZN(
        n18511) );
  NOR2_X2 U21651 ( .A1(n18508), .A2(n18717), .ZN(n18914) );
  NOR2_X1 U21652 ( .A1(n18509), .A2(n18532), .ZN(n18915) );
  AOI22_X1 U21653 ( .A1(n18937), .A2(n18914), .B1(n18915), .B2(n18581), .ZN(
        n18510) );
  OAI211_X1 U21654 ( .C1(n18512), .C2(n18536), .A(n18511), .B(n18510), .ZN(
        P3_U2871) );
  NAND2_X1 U21655 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18891), .ZN(n18872) );
  INV_X1 U21656 ( .A(n18872), .ZN(n18921) );
  NOR2_X2 U21657 ( .A1(n18798), .A2(n18513), .ZN(n18920) );
  AOI22_X1 U21658 ( .A1(n18937), .A2(n18921), .B1(n18920), .B2(n18530), .ZN(
        n18516) );
  NOR2_X1 U21659 ( .A1(n18514), .A2(n18532), .ZN(n18869) );
  AOI22_X1 U21660 ( .A1(n18884), .A2(n18922), .B1(n18869), .B2(n18581), .ZN(
        n18515) );
  OAI211_X1 U21661 ( .C1(n18517), .C2(n18536), .A(n18516), .B(n18515), .ZN(
        P3_U2872) );
  NAND2_X1 U21662 ( .A1(n18891), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18875) );
  INV_X1 U21663 ( .A(n18875), .ZN(n18929) );
  NOR2_X2 U21664 ( .A1(n18798), .A2(n18518), .ZN(n18926) );
  AOI22_X1 U21665 ( .A1(n18884), .A2(n18929), .B1(n18926), .B2(n18530), .ZN(
        n18522) );
  NOR2_X2 U21666 ( .A1(n18519), .A2(n18717), .ZN(n18927) );
  NOR2_X1 U21667 ( .A1(n18520), .A2(n18532), .ZN(n18928) );
  AOI22_X1 U21668 ( .A1(n18937), .A2(n18927), .B1(n18928), .B2(n18581), .ZN(
        n18521) );
  OAI211_X1 U21669 ( .C1(n18523), .C2(n18536), .A(n18522), .B(n18521), .ZN(
        P3_U2873) );
  NAND2_X1 U21670 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18891), .ZN(n18880) );
  NOR2_X2 U21671 ( .A1(n18798), .A2(n18524), .ZN(n18934) );
  AOI22_X1 U21672 ( .A1(n18937), .A2(n18935), .B1(n18934), .B2(n18530), .ZN(
        n18527) );
  AND2_X1 U21673 ( .A1(n18891), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18936) );
  NOR2_X1 U21674 ( .A1(n18525), .A2(n18532), .ZN(n18876) );
  AOI22_X1 U21675 ( .A1(n18877), .A2(n18936), .B1(n18876), .B2(n18581), .ZN(
        n18526) );
  OAI211_X1 U21676 ( .C1(n18528), .C2(n18536), .A(n18527), .B(n18526), .ZN(
        P3_U2874) );
  NAND2_X1 U21677 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18891), .ZN(n18951) );
  INV_X1 U21678 ( .A(n18951), .ZN(n18848) );
  NOR2_X2 U21679 ( .A1(n18529), .A2(n18798), .ZN(n18943) );
  AOI22_X1 U21680 ( .A1(n18884), .A2(n18848), .B1(n18943), .B2(n18530), .ZN(
        n18535) );
  NOR2_X2 U21681 ( .A1(n18717), .A2(n18531), .ZN(n18944) );
  NOR2_X1 U21682 ( .A1(n18533), .A2(n18532), .ZN(n18947) );
  AOI22_X1 U21683 ( .A1(n18937), .A2(n18944), .B1(n18947), .B2(n18581), .ZN(
        n18534) );
  OAI211_X1 U21684 ( .C1(n18537), .C2(n18536), .A(n18535), .B(n18534), .ZN(
        P3_U2875) );
  INV_X1 U21685 ( .A(n18896), .ZN(n18580) );
  NOR2_X2 U21686 ( .A1(n18719), .A2(n18621), .ZN(n18616) );
  NAND2_X1 U21687 ( .A1(n18996), .A2(n18893), .ZN(n18718) );
  NOR2_X1 U21688 ( .A1(n18621), .A2(n18718), .ZN(n18553) );
  AOI22_X1 U21689 ( .A1(n18884), .A2(n18895), .B1(n18894), .B2(n18553), .ZN(
        n18540) );
  NOR2_X1 U21690 ( .A1(n19004), .A2(n18713), .ZN(n18892) );
  INV_X1 U21691 ( .A(n18621), .ZN(n18577) );
  NOR2_X1 U21692 ( .A1(n18798), .A2(n18538), .ZN(n18889) );
  INV_X1 U21693 ( .A(n18889), .ZN(n18715) );
  NOR2_X1 U21694 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18715), .ZN(
        n18622) );
  AOI22_X1 U21695 ( .A1(n18891), .A2(n18892), .B1(n18577), .B2(n18622), .ZN(
        n18554) );
  AOI22_X1 U21696 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18554), .B1(
        n18897), .B2(n18946), .ZN(n18539) );
  OAI211_X1 U21697 ( .C1(n18580), .C2(n18615), .A(n18540), .B(n18539), .ZN(
        P3_U2876) );
  INV_X1 U21698 ( .A(n18903), .ZN(n18726) );
  AOI22_X1 U21699 ( .A1(n18884), .A2(n18902), .B1(n18901), .B2(n18553), .ZN(
        n18542) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18554), .B1(
        n18803), .B2(n18946), .ZN(n18541) );
  OAI211_X1 U21701 ( .C1(n18726), .C2(n18615), .A(n18542), .B(n18541), .ZN(
        P3_U2877) );
  AOI22_X1 U21702 ( .A1(n18833), .A2(n18946), .B1(n18907), .B2(n18553), .ZN(
        n18544) );
  AOI22_X1 U21703 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18554), .B1(
        n18877), .B2(n18908), .ZN(n18543) );
  OAI211_X1 U21704 ( .C1(n18836), .C2(n18615), .A(n18544), .B(n18543), .ZN(
        P3_U2878) );
  INV_X1 U21705 ( .A(n18915), .ZN(n18839) );
  AOI22_X1 U21706 ( .A1(n18884), .A2(n18914), .B1(n18913), .B2(n18553), .ZN(
        n18546) );
  AOI22_X1 U21707 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18554), .B1(
        n18916), .B2(n18946), .ZN(n18545) );
  OAI211_X1 U21708 ( .C1(n18839), .C2(n18615), .A(n18546), .B(n18545), .ZN(
        P3_U2879) );
  AOI22_X1 U21709 ( .A1(n18920), .A2(n18553), .B1(n18922), .B2(n18946), .ZN(
        n18548) );
  AOI22_X1 U21710 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18554), .B1(
        n18877), .B2(n18921), .ZN(n18547) );
  OAI211_X1 U21711 ( .C1(n18925), .C2(n18615), .A(n18548), .B(n18547), .ZN(
        P3_U2880) );
  INV_X1 U21712 ( .A(n18928), .ZN(n18786) );
  AOI22_X1 U21713 ( .A1(n18884), .A2(n18927), .B1(n18926), .B2(n18553), .ZN(
        n18550) );
  AOI22_X1 U21714 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18554), .B1(
        n18929), .B2(n18946), .ZN(n18549) );
  OAI211_X1 U21715 ( .C1(n18786), .C2(n18615), .A(n18550), .B(n18549), .ZN(
        P3_U2881) );
  AOI22_X1 U21716 ( .A1(n18934), .A2(n18553), .B1(n18936), .B2(n18946), .ZN(
        n18552) );
  AOI22_X1 U21717 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18554), .B1(
        n18877), .B2(n18935), .ZN(n18551) );
  OAI211_X1 U21718 ( .C1(n18941), .C2(n18615), .A(n18552), .B(n18551), .ZN(
        P3_U2882) );
  INV_X1 U21719 ( .A(n18947), .ZN(n18853) );
  AOI22_X1 U21720 ( .A1(n18884), .A2(n18944), .B1(n18943), .B2(n18553), .ZN(
        n18556) );
  AOI22_X1 U21721 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18554), .B1(
        n18848), .B2(n18946), .ZN(n18555) );
  OAI211_X1 U21722 ( .C1(n18853), .C2(n18615), .A(n18556), .B(n18555), .ZN(
        P3_U2883) );
  INV_X1 U21723 ( .A(n18644), .ZN(n18747) );
  NAND2_X1 U21724 ( .A1(n18747), .A2(n18577), .ZN(n18638) );
  NOR2_X1 U21725 ( .A1(n18616), .A2(n18640), .ZN(n18599) );
  NOR2_X1 U21726 ( .A1(n19023), .A2(n18599), .ZN(n18573) );
  AOI22_X1 U21727 ( .A1(n18897), .A2(n18594), .B1(n18894), .B2(n18573), .ZN(
        n18560) );
  AOI221_X1 U21728 ( .B1(n18599), .B2(n18855), .C1(n18599), .C2(n18557), .A(
        n18746), .ZN(n18558) );
  INV_X1 U21729 ( .A(n18558), .ZN(n18574) );
  AOI22_X1 U21730 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18574), .B1(
        n18895), .B2(n18946), .ZN(n18559) );
  OAI211_X1 U21731 ( .C1(n18580), .C2(n18638), .A(n18560), .B(n18559), .ZN(
        P3_U2884) );
  AOI22_X1 U21732 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18574), .B1(
        n18901), .B2(n18573), .ZN(n18562) );
  AOI22_X1 U21733 ( .A1(n18803), .A2(n18594), .B1(n18902), .B2(n18946), .ZN(
        n18561) );
  OAI211_X1 U21734 ( .C1(n18726), .C2(n18638), .A(n18562), .B(n18561), .ZN(
        P3_U2885) );
  AOI22_X1 U21735 ( .A1(n18833), .A2(n18594), .B1(n18907), .B2(n18573), .ZN(
        n18564) );
  AOI22_X1 U21736 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18574), .B1(
        n18908), .B2(n18946), .ZN(n18563) );
  OAI211_X1 U21737 ( .C1(n18836), .C2(n18638), .A(n18564), .B(n18563), .ZN(
        P3_U2886) );
  AOI22_X1 U21738 ( .A1(n18913), .A2(n18573), .B1(n18914), .B2(n18946), .ZN(
        n18566) );
  AOI22_X1 U21739 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18574), .B1(
        n18916), .B2(n18581), .ZN(n18565) );
  OAI211_X1 U21740 ( .C1(n18839), .C2(n18638), .A(n18566), .B(n18565), .ZN(
        P3_U2887) );
  AOI22_X1 U21741 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18574), .B1(
        n18920), .B2(n18573), .ZN(n18568) );
  AOI22_X1 U21742 ( .A1(n18921), .A2(n18946), .B1(n18922), .B2(n18581), .ZN(
        n18567) );
  OAI211_X1 U21743 ( .C1(n18925), .C2(n18638), .A(n18568), .B(n18567), .ZN(
        P3_U2888) );
  AOI22_X1 U21744 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18574), .B1(
        n18926), .B2(n18573), .ZN(n18570) );
  AOI22_X1 U21745 ( .A1(n18929), .A2(n18594), .B1(n18927), .B2(n18946), .ZN(
        n18569) );
  OAI211_X1 U21746 ( .C1(n18786), .C2(n18638), .A(n18570), .B(n18569), .ZN(
        P3_U2889) );
  AOI22_X1 U21747 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18574), .B1(
        n18934), .B2(n18573), .ZN(n18572) );
  AOI22_X1 U21748 ( .A1(n18935), .A2(n18946), .B1(n18936), .B2(n18581), .ZN(
        n18571) );
  OAI211_X1 U21749 ( .C1(n18941), .C2(n18638), .A(n18572), .B(n18571), .ZN(
        P3_U2890) );
  AOI22_X1 U21750 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18574), .B1(
        n18943), .B2(n18573), .ZN(n18576) );
  AOI22_X1 U21751 ( .A1(n18848), .A2(n18594), .B1(n18944), .B2(n18946), .ZN(
        n18575) );
  OAI211_X1 U21752 ( .C1(n18853), .C2(n18638), .A(n18576), .B(n18575), .ZN(
        P3_U2891) );
  INV_X1 U21753 ( .A(n18995), .ZN(n18772) );
  NAND2_X1 U21754 ( .A1(n18772), .A2(n18577), .ZN(n18649) );
  AOI22_X1 U21755 ( .A1(n18895), .A2(n18594), .B1(n18894), .B2(n18595), .ZN(
        n18579) );
  AOI21_X1 U21756 ( .B1(n18996), .B2(n18855), .A(n18715), .ZN(n18667) );
  NAND2_X1 U21757 ( .A1(n18577), .A2(n18667), .ZN(n18596) );
  AOI22_X1 U21758 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18596), .B1(
        n18897), .B2(n18616), .ZN(n18578) );
  OAI211_X1 U21759 ( .C1(n18580), .C2(n18649), .A(n18579), .B(n18578), .ZN(
        P3_U2892) );
  AOI22_X1 U21760 ( .A1(n18803), .A2(n18616), .B1(n18901), .B2(n18595), .ZN(
        n18583) );
  AOI22_X1 U21761 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18596), .B1(
        n18902), .B2(n18581), .ZN(n18582) );
  OAI211_X1 U21762 ( .C1(n18726), .C2(n18649), .A(n18583), .B(n18582), .ZN(
        P3_U2893) );
  AOI22_X1 U21763 ( .A1(n18907), .A2(n18595), .B1(n18908), .B2(n18594), .ZN(
        n18585) );
  AOI22_X1 U21764 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18596), .B1(
        n18833), .B2(n18616), .ZN(n18584) );
  OAI211_X1 U21765 ( .C1(n18836), .C2(n18649), .A(n18585), .B(n18584), .ZN(
        P3_U2894) );
  AOI22_X1 U21766 ( .A1(n18916), .A2(n18616), .B1(n18913), .B2(n18595), .ZN(
        n18587) );
  AOI22_X1 U21767 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18596), .B1(
        n18914), .B2(n18594), .ZN(n18586) );
  OAI211_X1 U21768 ( .C1(n18839), .C2(n18649), .A(n18587), .B(n18586), .ZN(
        P3_U2895) );
  AOI22_X1 U21769 ( .A1(n18921), .A2(n18594), .B1(n18920), .B2(n18595), .ZN(
        n18589) );
  AOI22_X1 U21770 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18596), .B1(
        n18922), .B2(n18616), .ZN(n18588) );
  OAI211_X1 U21771 ( .C1(n18925), .C2(n18649), .A(n18589), .B(n18588), .ZN(
        P3_U2896) );
  AOI22_X1 U21772 ( .A1(n18929), .A2(n18616), .B1(n18926), .B2(n18595), .ZN(
        n18591) );
  AOI22_X1 U21773 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18596), .B1(
        n18927), .B2(n18594), .ZN(n18590) );
  OAI211_X1 U21774 ( .C1(n18786), .C2(n18649), .A(n18591), .B(n18590), .ZN(
        P3_U2897) );
  AOI22_X1 U21775 ( .A1(n18935), .A2(n18594), .B1(n18934), .B2(n18595), .ZN(
        n18593) );
  AOI22_X1 U21776 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18596), .B1(
        n18936), .B2(n18616), .ZN(n18592) );
  OAI211_X1 U21777 ( .C1(n18941), .C2(n18649), .A(n18593), .B(n18592), .ZN(
        P3_U2898) );
  AOI22_X1 U21778 ( .A1(n18943), .A2(n18595), .B1(n18944), .B2(n18594), .ZN(
        n18598) );
  AOI22_X1 U21779 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18596), .B1(
        n18848), .B2(n18616), .ZN(n18597) );
  OAI211_X1 U21780 ( .C1(n18853), .C2(n18649), .A(n18598), .B(n18597), .ZN(
        P3_U2899) );
  INV_X1 U21781 ( .A(n18649), .ZN(n18663) );
  NOR2_X2 U21782 ( .A1(n18997), .A2(n18669), .ZN(n18686) );
  NOR2_X1 U21783 ( .A1(n18663), .A2(n18686), .ZN(n18645) );
  NOR2_X1 U21784 ( .A1(n19023), .A2(n18645), .ZN(n18617) );
  AOI22_X1 U21785 ( .A1(n18897), .A2(n18640), .B1(n18894), .B2(n18617), .ZN(
        n18602) );
  OAI21_X1 U21786 ( .B1(n18599), .B2(n18855), .A(n18645), .ZN(n18600) );
  OAI211_X1 U21787 ( .C1(n18686), .C2(n19125), .A(n18857), .B(n18600), .ZN(
        n18618) );
  AOI22_X1 U21788 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18618), .B1(
        n18896), .B2(n18686), .ZN(n18601) );
  OAI211_X1 U21789 ( .C1(n18861), .C2(n18615), .A(n18602), .B(n18601), .ZN(
        P3_U2900) );
  AOI22_X1 U21790 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18618), .B1(
        n18901), .B2(n18617), .ZN(n18604) );
  AOI22_X1 U21791 ( .A1(n18903), .A2(n18686), .B1(n18902), .B2(n18616), .ZN(
        n18603) );
  OAI211_X1 U21792 ( .C1(n18906), .C2(n18638), .A(n18604), .B(n18603), .ZN(
        P3_U2901) );
  AOI22_X1 U21793 ( .A1(n18907), .A2(n18617), .B1(n18908), .B2(n18616), .ZN(
        n18606) );
  AOI22_X1 U21794 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18618), .B1(
        n18909), .B2(n18686), .ZN(n18605) );
  OAI211_X1 U21795 ( .C1(n18912), .C2(n18638), .A(n18606), .B(n18605), .ZN(
        P3_U2902) );
  AOI22_X1 U21796 ( .A1(n18913), .A2(n18617), .B1(n18914), .B2(n18616), .ZN(
        n18608) );
  AOI22_X1 U21797 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18618), .B1(
        n18915), .B2(n18686), .ZN(n18607) );
  OAI211_X1 U21798 ( .C1(n18868), .C2(n18638), .A(n18608), .B(n18607), .ZN(
        P3_U2903) );
  INV_X1 U21799 ( .A(n18686), .ZN(n18684) );
  AOI22_X1 U21800 ( .A1(n18921), .A2(n18616), .B1(n18920), .B2(n18617), .ZN(
        n18610) );
  AOI22_X1 U21801 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18618), .B1(
        n18922), .B2(n18640), .ZN(n18609) );
  OAI211_X1 U21802 ( .C1(n18925), .C2(n18684), .A(n18610), .B(n18609), .ZN(
        P3_U2904) );
  AOI22_X1 U21803 ( .A1(n18927), .A2(n18616), .B1(n18926), .B2(n18617), .ZN(
        n18612) );
  AOI22_X1 U21804 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18618), .B1(
        n18928), .B2(n18686), .ZN(n18611) );
  OAI211_X1 U21805 ( .C1(n18875), .C2(n18638), .A(n18612), .B(n18611), .ZN(
        P3_U2905) );
  AOI22_X1 U21806 ( .A1(n18934), .A2(n18617), .B1(n18936), .B2(n18640), .ZN(
        n18614) );
  AOI22_X1 U21807 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18618), .B1(
        n18876), .B2(n18686), .ZN(n18613) );
  OAI211_X1 U21808 ( .C1(n18880), .C2(n18615), .A(n18614), .B(n18613), .ZN(
        P3_U2906) );
  AOI22_X1 U21809 ( .A1(n18943), .A2(n18617), .B1(n18944), .B2(n18616), .ZN(
        n18620) );
  AOI22_X1 U21810 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18618), .B1(
        n18947), .B2(n18686), .ZN(n18619) );
  OAI211_X1 U21811 ( .C1(n18951), .C2(n18638), .A(n18620), .B(n18619), .ZN(
        P3_U2907) );
  NOR2_X1 U21812 ( .A1(n18669), .A2(n18718), .ZN(n18639) );
  AOI22_X1 U21813 ( .A1(n18897), .A2(n18663), .B1(n18894), .B2(n18639), .ZN(
        n18625) );
  NOR2_X1 U21814 ( .A1(n18996), .A2(n18621), .ZN(n18623) );
  AOI22_X1 U21815 ( .A1(n18891), .A2(n18623), .B1(n18668), .B2(n18622), .ZN(
        n18641) );
  NOR2_X2 U21816 ( .A1(n18719), .A2(n18669), .ZN(n18707) );
  AOI22_X1 U21817 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18641), .B1(
        n18896), .B2(n18707), .ZN(n18624) );
  OAI211_X1 U21818 ( .C1(n18861), .C2(n18638), .A(n18625), .B(n18624), .ZN(
        P3_U2908) );
  AOI22_X1 U21819 ( .A1(n18803), .A2(n18663), .B1(n18901), .B2(n18639), .ZN(
        n18627) );
  AOI22_X1 U21820 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18641), .B1(
        n18902), .B2(n18640), .ZN(n18626) );
  OAI211_X1 U21821 ( .C1(n18726), .C2(n18694), .A(n18627), .B(n18626), .ZN(
        P3_U2909) );
  AOI22_X1 U21822 ( .A1(n18833), .A2(n18663), .B1(n18907), .B2(n18639), .ZN(
        n18629) );
  AOI22_X1 U21823 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18641), .B1(
        n18908), .B2(n18640), .ZN(n18628) );
  OAI211_X1 U21824 ( .C1(n18836), .C2(n18694), .A(n18629), .B(n18628), .ZN(
        P3_U2910) );
  AOI22_X1 U21825 ( .A1(n18916), .A2(n18663), .B1(n18913), .B2(n18639), .ZN(
        n18631) );
  AOI22_X1 U21826 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18641), .B1(
        n18914), .B2(n18640), .ZN(n18630) );
  OAI211_X1 U21827 ( .C1(n18839), .C2(n18694), .A(n18631), .B(n18630), .ZN(
        P3_U2911) );
  AOI22_X1 U21828 ( .A1(n18921), .A2(n18640), .B1(n18920), .B2(n18639), .ZN(
        n18633) );
  AOI22_X1 U21829 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18641), .B1(
        n18922), .B2(n18663), .ZN(n18632) );
  OAI211_X1 U21830 ( .C1(n18925), .C2(n18694), .A(n18633), .B(n18632), .ZN(
        P3_U2912) );
  AOI22_X1 U21831 ( .A1(n18929), .A2(n18663), .B1(n18926), .B2(n18639), .ZN(
        n18635) );
  AOI22_X1 U21832 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18641), .B1(
        n18927), .B2(n18640), .ZN(n18634) );
  OAI211_X1 U21833 ( .C1(n18786), .C2(n18694), .A(n18635), .B(n18634), .ZN(
        P3_U2913) );
  AOI22_X1 U21834 ( .A1(n18934), .A2(n18639), .B1(n18936), .B2(n18663), .ZN(
        n18637) );
  AOI22_X1 U21835 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18641), .B1(
        n18876), .B2(n18707), .ZN(n18636) );
  OAI211_X1 U21836 ( .C1(n18880), .C2(n18638), .A(n18637), .B(n18636), .ZN(
        P3_U2914) );
  AOI22_X1 U21837 ( .A1(n18848), .A2(n18663), .B1(n18943), .B2(n18639), .ZN(
        n18643) );
  AOI22_X1 U21838 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18641), .B1(
        n18944), .B2(n18640), .ZN(n18642) );
  OAI211_X1 U21839 ( .C1(n18853), .C2(n18694), .A(n18643), .B(n18642), .ZN(
        P3_U2915) );
  NOR2_X2 U21840 ( .A1(n18644), .A2(n18669), .ZN(n18741) );
  NOR2_X1 U21841 ( .A1(n18707), .A2(n18741), .ZN(n18690) );
  NOR2_X1 U21842 ( .A1(n19023), .A2(n18690), .ZN(n18662) );
  AOI22_X1 U21843 ( .A1(n18897), .A2(n18686), .B1(n18894), .B2(n18662), .ZN(
        n18648) );
  AOI221_X1 U21844 ( .B1(n18690), .B2(n18855), .C1(n18690), .C2(n18645), .A(
        n18746), .ZN(n18646) );
  INV_X1 U21845 ( .A(n18646), .ZN(n18664) );
  AOI22_X1 U21846 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18664), .B1(
        n18896), .B2(n18741), .ZN(n18647) );
  OAI211_X1 U21847 ( .C1(n18861), .C2(n18649), .A(n18648), .B(n18647), .ZN(
        P3_U2916) );
  AOI22_X1 U21848 ( .A1(n18901), .A2(n18662), .B1(n18902), .B2(n18663), .ZN(
        n18651) );
  AOI22_X1 U21849 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18664), .B1(
        n18903), .B2(n18741), .ZN(n18650) );
  OAI211_X1 U21850 ( .C1(n18906), .C2(n18684), .A(n18651), .B(n18650), .ZN(
        P3_U2917) );
  AOI22_X1 U21851 ( .A1(n18907), .A2(n18662), .B1(n18908), .B2(n18663), .ZN(
        n18653) );
  AOI22_X1 U21852 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18664), .B1(
        n18909), .B2(n18741), .ZN(n18652) );
  OAI211_X1 U21853 ( .C1(n18912), .C2(n18684), .A(n18653), .B(n18652), .ZN(
        P3_U2918) );
  AOI22_X1 U21854 ( .A1(n18913), .A2(n18662), .B1(n18914), .B2(n18663), .ZN(
        n18655) );
  AOI22_X1 U21855 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18664), .B1(
        n18915), .B2(n18741), .ZN(n18654) );
  OAI211_X1 U21856 ( .C1(n18868), .C2(n18684), .A(n18655), .B(n18654), .ZN(
        P3_U2919) );
  INV_X1 U21857 ( .A(n18741), .ZN(n18712) );
  AOI22_X1 U21858 ( .A1(n18921), .A2(n18663), .B1(n18920), .B2(n18662), .ZN(
        n18657) );
  AOI22_X1 U21859 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18664), .B1(
        n18922), .B2(n18686), .ZN(n18656) );
  OAI211_X1 U21860 ( .C1(n18925), .C2(n18712), .A(n18657), .B(n18656), .ZN(
        P3_U2920) );
  AOI22_X1 U21861 ( .A1(n18927), .A2(n18663), .B1(n18926), .B2(n18662), .ZN(
        n18659) );
  AOI22_X1 U21862 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18664), .B1(
        n18928), .B2(n18741), .ZN(n18658) );
  OAI211_X1 U21863 ( .C1(n18875), .C2(n18684), .A(n18659), .B(n18658), .ZN(
        P3_U2921) );
  AOI22_X1 U21864 ( .A1(n18935), .A2(n18663), .B1(n18934), .B2(n18662), .ZN(
        n18661) );
  AOI22_X1 U21865 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18664), .B1(
        n18936), .B2(n18686), .ZN(n18660) );
  OAI211_X1 U21866 ( .C1(n18941), .C2(n18712), .A(n18661), .B(n18660), .ZN(
        P3_U2922) );
  AOI22_X1 U21867 ( .A1(n18848), .A2(n18686), .B1(n18943), .B2(n18662), .ZN(
        n18666) );
  AOI22_X1 U21868 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18664), .B1(
        n18944), .B2(n18663), .ZN(n18665) );
  OAI211_X1 U21869 ( .C1(n18853), .C2(n18712), .A(n18666), .B(n18665), .ZN(
        P3_U2923) );
  AOI22_X1 U21870 ( .A1(n18897), .A2(n18707), .B1(n18894), .B2(n18685), .ZN(
        n18671) );
  NAND2_X1 U21871 ( .A1(n18668), .A2(n18667), .ZN(n18687) );
  NOR2_X2 U21872 ( .A1(n18995), .A2(n18669), .ZN(n18766) );
  AOI22_X1 U21873 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18687), .B1(
        n18896), .B2(n18766), .ZN(n18670) );
  OAI211_X1 U21874 ( .C1(n18861), .C2(n18684), .A(n18671), .B(n18670), .ZN(
        P3_U2924) );
  AOI22_X1 U21875 ( .A1(n18803), .A2(n18707), .B1(n18901), .B2(n18685), .ZN(
        n18673) );
  AOI22_X1 U21876 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18687), .B1(
        n18902), .B2(n18686), .ZN(n18672) );
  OAI211_X1 U21877 ( .C1(n18726), .C2(n18761), .A(n18673), .B(n18672), .ZN(
        P3_U2925) );
  AOI22_X1 U21878 ( .A1(n18907), .A2(n18685), .B1(n18908), .B2(n18686), .ZN(
        n18675) );
  AOI22_X1 U21879 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18687), .B1(
        n18909), .B2(n18766), .ZN(n18674) );
  OAI211_X1 U21880 ( .C1(n18912), .C2(n18694), .A(n18675), .B(n18674), .ZN(
        P3_U2926) );
  AOI22_X1 U21881 ( .A1(n18916), .A2(n18707), .B1(n18913), .B2(n18685), .ZN(
        n18677) );
  AOI22_X1 U21882 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18687), .B1(
        n18914), .B2(n18686), .ZN(n18676) );
  OAI211_X1 U21883 ( .C1(n18839), .C2(n18761), .A(n18677), .B(n18676), .ZN(
        P3_U2927) );
  AOI22_X1 U21884 ( .A1(n18921), .A2(n18686), .B1(n18920), .B2(n18685), .ZN(
        n18679) );
  AOI22_X1 U21885 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18687), .B1(
        n18922), .B2(n18707), .ZN(n18678) );
  OAI211_X1 U21886 ( .C1(n18925), .C2(n18761), .A(n18679), .B(n18678), .ZN(
        P3_U2928) );
  AOI22_X1 U21887 ( .A1(n18927), .A2(n18686), .B1(n18926), .B2(n18685), .ZN(
        n18681) );
  AOI22_X1 U21888 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18687), .B1(
        n18928), .B2(n18766), .ZN(n18680) );
  OAI211_X1 U21889 ( .C1(n18875), .C2(n18694), .A(n18681), .B(n18680), .ZN(
        P3_U2929) );
  AOI22_X1 U21890 ( .A1(n18934), .A2(n18685), .B1(n18936), .B2(n18707), .ZN(
        n18683) );
  AOI22_X1 U21891 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18687), .B1(
        n18876), .B2(n18766), .ZN(n18682) );
  OAI211_X1 U21892 ( .C1(n18880), .C2(n18684), .A(n18683), .B(n18682), .ZN(
        P3_U2930) );
  AOI22_X1 U21893 ( .A1(n18848), .A2(n18707), .B1(n18943), .B2(n18685), .ZN(
        n18689) );
  AOI22_X1 U21894 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18687), .B1(
        n18944), .B2(n18686), .ZN(n18688) );
  OAI211_X1 U21895 ( .C1(n18853), .C2(n18761), .A(n18689), .B(n18688), .ZN(
        P3_U2931) );
  INV_X1 U21896 ( .A(n18771), .ZN(n18794) );
  NOR2_X2 U21897 ( .A1(n18997), .A2(n18794), .ZN(n18790) );
  NOR2_X1 U21898 ( .A1(n18766), .A2(n18790), .ZN(n18748) );
  NOR2_X1 U21899 ( .A1(n19023), .A2(n18748), .ZN(n18708) );
  AOI22_X1 U21900 ( .A1(n18897), .A2(n18741), .B1(n18894), .B2(n18708), .ZN(
        n18693) );
  OAI21_X1 U21901 ( .B1(n18690), .B2(n18855), .A(n18748), .ZN(n18691) );
  OAI211_X1 U21902 ( .C1(n18790), .C2(n19125), .A(n18857), .B(n18691), .ZN(
        n18709) );
  AOI22_X1 U21903 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18709), .B1(
        n18896), .B2(n18790), .ZN(n18692) );
  OAI211_X1 U21904 ( .C1(n18861), .C2(n18694), .A(n18693), .B(n18692), .ZN(
        P3_U2932) );
  INV_X1 U21905 ( .A(n18790), .ZN(n18783) );
  AOI22_X1 U21906 ( .A1(n18803), .A2(n18741), .B1(n18901), .B2(n18708), .ZN(
        n18696) );
  AOI22_X1 U21907 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18709), .B1(
        n18902), .B2(n18707), .ZN(n18695) );
  OAI211_X1 U21908 ( .C1(n18726), .C2(n18783), .A(n18696), .B(n18695), .ZN(
        P3_U2933) );
  AOI22_X1 U21909 ( .A1(n18907), .A2(n18708), .B1(n18908), .B2(n18707), .ZN(
        n18698) );
  AOI22_X1 U21910 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18709), .B1(
        n18909), .B2(n18790), .ZN(n18697) );
  OAI211_X1 U21911 ( .C1(n18912), .C2(n18712), .A(n18698), .B(n18697), .ZN(
        P3_U2934) );
  AOI22_X1 U21912 ( .A1(n18913), .A2(n18708), .B1(n18914), .B2(n18707), .ZN(
        n18700) );
  AOI22_X1 U21913 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18709), .B1(
        n18915), .B2(n18790), .ZN(n18699) );
  OAI211_X1 U21914 ( .C1(n18868), .C2(n18712), .A(n18700), .B(n18699), .ZN(
        P3_U2935) );
  AOI22_X1 U21915 ( .A1(n18921), .A2(n18707), .B1(n18920), .B2(n18708), .ZN(
        n18702) );
  AOI22_X1 U21916 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18709), .B1(
        n18922), .B2(n18741), .ZN(n18701) );
  OAI211_X1 U21917 ( .C1(n18925), .C2(n18783), .A(n18702), .B(n18701), .ZN(
        P3_U2936) );
  AOI22_X1 U21918 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18709), .B1(
        n18926), .B2(n18708), .ZN(n18704) );
  AOI22_X1 U21919 ( .A1(n18928), .A2(n18790), .B1(n18927), .B2(n18707), .ZN(
        n18703) );
  OAI211_X1 U21920 ( .C1(n18875), .C2(n18712), .A(n18704), .B(n18703), .ZN(
        P3_U2937) );
  AOI22_X1 U21921 ( .A1(n18935), .A2(n18707), .B1(n18934), .B2(n18708), .ZN(
        n18706) );
  AOI22_X1 U21922 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18709), .B1(
        n18936), .B2(n18741), .ZN(n18705) );
  OAI211_X1 U21923 ( .C1(n18941), .C2(n18783), .A(n18706), .B(n18705), .ZN(
        P3_U2938) );
  AOI22_X1 U21924 ( .A1(n18943), .A2(n18708), .B1(n18944), .B2(n18707), .ZN(
        n18711) );
  AOI22_X1 U21925 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18709), .B1(
        n18947), .B2(n18790), .ZN(n18710) );
  OAI211_X1 U21926 ( .C1(n18951), .C2(n18712), .A(n18711), .B(n18710), .ZN(
        P3_U2939) );
  OR2_X1 U21927 ( .A1(n18713), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18716) );
  NAND2_X1 U21928 ( .A1(n18771), .A2(n18996), .ZN(n18714) );
  OAI22_X1 U21929 ( .A1(n18717), .A2(n18716), .B1(n18715), .B2(n18714), .ZN(
        n18739) );
  NOR2_X1 U21930 ( .A1(n18794), .A2(n18718), .ZN(n18742) );
  AOI22_X1 U21931 ( .A1(n18895), .A2(n18741), .B1(n18894), .B2(n18742), .ZN(
        n18721) );
  NOR2_X1 U21932 ( .A1(n18794), .A2(n18719), .ZN(n18723) );
  CLKBUF_X1 U21933 ( .A(n18723), .Z(n18822) );
  AOI22_X1 U21934 ( .A1(n18896), .A2(n18822), .B1(n18897), .B2(n18766), .ZN(
        n18720) );
  OAI211_X1 U21935 ( .C1(n18722), .C2(n18739), .A(n18721), .B(n18720), .ZN(
        P3_U2940) );
  INV_X1 U21936 ( .A(n18723), .ZN(n18820) );
  AOI22_X1 U21937 ( .A1(n18803), .A2(n18766), .B1(n18901), .B2(n18742), .ZN(
        n18725) );
  INV_X1 U21938 ( .A(n18739), .ZN(n18743) );
  AOI22_X1 U21939 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18743), .B1(
        n18902), .B2(n18741), .ZN(n18724) );
  OAI211_X1 U21940 ( .C1(n18726), .C2(n18820), .A(n18725), .B(n18724), .ZN(
        P3_U2941) );
  AOI22_X1 U21941 ( .A1(n18907), .A2(n18742), .B1(n18908), .B2(n18741), .ZN(
        n18728) );
  AOI22_X1 U21942 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18743), .B1(
        n18909), .B2(n18822), .ZN(n18727) );
  OAI211_X1 U21943 ( .C1(n18912), .C2(n18761), .A(n18728), .B(n18727), .ZN(
        P3_U2942) );
  AOI22_X1 U21944 ( .A1(n18913), .A2(n18742), .B1(n18914), .B2(n18741), .ZN(
        n18730) );
  AOI22_X1 U21945 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18743), .B1(
        n18915), .B2(n18822), .ZN(n18729) );
  OAI211_X1 U21946 ( .C1(n18868), .C2(n18761), .A(n18730), .B(n18729), .ZN(
        P3_U2943) );
  AOI22_X1 U21947 ( .A1(n18921), .A2(n18741), .B1(n18920), .B2(n18742), .ZN(
        n18732) );
  AOI22_X1 U21948 ( .A1(n18869), .A2(n18822), .B1(n18922), .B2(n18766), .ZN(
        n18731) );
  OAI211_X1 U21949 ( .C1(n18733), .C2(n18739), .A(n18732), .B(n18731), .ZN(
        P3_U2944) );
  AOI22_X1 U21950 ( .A1(n18929), .A2(n18766), .B1(n18926), .B2(n18742), .ZN(
        n18735) );
  AOI22_X1 U21951 ( .A1(n18928), .A2(n18822), .B1(n18927), .B2(n18741), .ZN(
        n18734) );
  OAI211_X1 U21952 ( .C1(n18736), .C2(n18739), .A(n18735), .B(n18734), .ZN(
        P3_U2945) );
  AOI22_X1 U21953 ( .A1(n18935), .A2(n18741), .B1(n18934), .B2(n18742), .ZN(
        n18738) );
  AOI22_X1 U21954 ( .A1(n18876), .A2(n18822), .B1(n18936), .B2(n18766), .ZN(
        n18737) );
  OAI211_X1 U21955 ( .C1(n18740), .C2(n18739), .A(n18738), .B(n18737), .ZN(
        P3_U2946) );
  AOI22_X1 U21956 ( .A1(n18943), .A2(n18742), .B1(n18944), .B2(n18741), .ZN(
        n18745) );
  AOI22_X1 U21957 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18743), .B1(
        n18947), .B2(n18822), .ZN(n18744) );
  OAI211_X1 U21958 ( .C1(n18951), .C2(n18761), .A(n18745), .B(n18744), .ZN(
        P3_U2947) );
  INV_X1 U21959 ( .A(n18746), .ZN(n18750) );
  NAND2_X1 U21960 ( .A1(n18747), .A2(n18771), .ZN(n18842) );
  OAI211_X1 U21961 ( .C1(n18748), .C2(n18855), .A(n18820), .B(n18842), .ZN(
        n18749) );
  NAND2_X1 U21962 ( .A1(n18750), .A2(n18749), .ZN(n18768) );
  AOI21_X1 U21963 ( .B1(n18820), .B2(n18842), .A(n19023), .ZN(n18767) );
  AOI22_X1 U21964 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18768), .B1(
        n18894), .B2(n18767), .ZN(n18752) );
  AOI22_X1 U21965 ( .A1(n18896), .A2(n18849), .B1(n18897), .B2(n18790), .ZN(
        n18751) );
  OAI211_X1 U21966 ( .C1(n18861), .C2(n18761), .A(n18752), .B(n18751), .ZN(
        P3_U2948) );
  AOI22_X1 U21967 ( .A1(n18901), .A2(n18767), .B1(n18902), .B2(n18766), .ZN(
        n18754) );
  AOI22_X1 U21968 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18768), .B1(
        n18903), .B2(n18849), .ZN(n18753) );
  OAI211_X1 U21969 ( .C1(n18906), .C2(n18783), .A(n18754), .B(n18753), .ZN(
        P3_U2949) );
  AOI22_X1 U21970 ( .A1(n18833), .A2(n18790), .B1(n18907), .B2(n18767), .ZN(
        n18756) );
  AOI22_X1 U21971 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18768), .B1(
        n18908), .B2(n18766), .ZN(n18755) );
  OAI211_X1 U21972 ( .C1(n18836), .C2(n18842), .A(n18756), .B(n18755), .ZN(
        P3_U2950) );
  AOI22_X1 U21973 ( .A1(n18916), .A2(n18790), .B1(n18913), .B2(n18767), .ZN(
        n18758) );
  AOI22_X1 U21974 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18768), .B1(
        n18914), .B2(n18766), .ZN(n18757) );
  OAI211_X1 U21975 ( .C1(n18839), .C2(n18842), .A(n18758), .B(n18757), .ZN(
        P3_U2951) );
  AOI22_X1 U21976 ( .A1(n18920), .A2(n18767), .B1(n18922), .B2(n18790), .ZN(
        n18760) );
  AOI22_X1 U21977 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18768), .B1(
        n18869), .B2(n18849), .ZN(n18759) );
  OAI211_X1 U21978 ( .C1(n18872), .C2(n18761), .A(n18760), .B(n18759), .ZN(
        P3_U2952) );
  AOI22_X1 U21979 ( .A1(n18929), .A2(n18790), .B1(n18926), .B2(n18767), .ZN(
        n18763) );
  AOI22_X1 U21980 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18768), .B1(
        n18927), .B2(n18766), .ZN(n18762) );
  OAI211_X1 U21981 ( .C1(n18786), .C2(n18842), .A(n18763), .B(n18762), .ZN(
        P3_U2953) );
  AOI22_X1 U21982 ( .A1(n18935), .A2(n18766), .B1(n18934), .B2(n18767), .ZN(
        n18765) );
  AOI22_X1 U21983 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18768), .B1(
        n18936), .B2(n18790), .ZN(n18764) );
  OAI211_X1 U21984 ( .C1(n18941), .C2(n18842), .A(n18765), .B(n18764), .ZN(
        P3_U2954) );
  AOI22_X1 U21985 ( .A1(n18943), .A2(n18767), .B1(n18944), .B2(n18766), .ZN(
        n18770) );
  AOI22_X1 U21986 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18768), .B1(
        n18947), .B2(n18849), .ZN(n18769) );
  OAI211_X1 U21987 ( .C1(n18951), .C2(n18783), .A(n18770), .B(n18769), .ZN(
        P3_U2955) );
  NOR2_X1 U21988 ( .A1(n18996), .A2(n18794), .ZN(n18828) );
  AND2_X1 U21989 ( .A1(n18893), .A2(n18828), .ZN(n18789) );
  AOI22_X1 U21990 ( .A1(n18897), .A2(n18822), .B1(n18894), .B2(n18789), .ZN(
        n18774) );
  OAI211_X1 U21991 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18891), .A(
        n18889), .B(n18771), .ZN(n18791) );
  NAND2_X1 U21992 ( .A1(n18772), .A2(n18771), .ZN(n18881) );
  INV_X1 U21993 ( .A(n18881), .ZN(n18883) );
  AOI22_X1 U21994 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18791), .B1(
        n18883), .B2(n18896), .ZN(n18773) );
  OAI211_X1 U21995 ( .C1(n18861), .C2(n18783), .A(n18774), .B(n18773), .ZN(
        P3_U2956) );
  AOI22_X1 U21996 ( .A1(n18901), .A2(n18789), .B1(n18902), .B2(n18790), .ZN(
        n18776) );
  AOI22_X1 U21997 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18791), .B1(
        n18883), .B2(n18903), .ZN(n18775) );
  OAI211_X1 U21998 ( .C1(n18906), .C2(n18820), .A(n18776), .B(n18775), .ZN(
        P3_U2957) );
  AOI22_X1 U21999 ( .A1(n18907), .A2(n18789), .B1(n18908), .B2(n18790), .ZN(
        n18778) );
  AOI22_X1 U22000 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18791), .B1(
        n18883), .B2(n18909), .ZN(n18777) );
  OAI211_X1 U22001 ( .C1(n18912), .C2(n18820), .A(n18778), .B(n18777), .ZN(
        P3_U2958) );
  AOI22_X1 U22002 ( .A1(n18916), .A2(n18822), .B1(n18913), .B2(n18789), .ZN(
        n18780) );
  AOI22_X1 U22003 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18791), .B1(
        n18914), .B2(n18790), .ZN(n18779) );
  OAI211_X1 U22004 ( .C1(n18881), .C2(n18839), .A(n18780), .B(n18779), .ZN(
        P3_U2959) );
  AOI22_X1 U22005 ( .A1(n18920), .A2(n18789), .B1(n18922), .B2(n18822), .ZN(
        n18782) );
  AOI22_X1 U22006 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18791), .B1(
        n18883), .B2(n18869), .ZN(n18781) );
  OAI211_X1 U22007 ( .C1(n18872), .C2(n18783), .A(n18782), .B(n18781), .ZN(
        P3_U2960) );
  AOI22_X1 U22008 ( .A1(n18929), .A2(n18822), .B1(n18926), .B2(n18789), .ZN(
        n18785) );
  AOI22_X1 U22009 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18791), .B1(
        n18927), .B2(n18790), .ZN(n18784) );
  OAI211_X1 U22010 ( .C1(n18881), .C2(n18786), .A(n18785), .B(n18784), .ZN(
        P3_U2961) );
  AOI22_X1 U22011 ( .A1(n18935), .A2(n18790), .B1(n18934), .B2(n18789), .ZN(
        n18788) );
  AOI22_X1 U22012 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18791), .B1(
        n18936), .B2(n18822), .ZN(n18787) );
  OAI211_X1 U22013 ( .C1(n18881), .C2(n18941), .A(n18788), .B(n18787), .ZN(
        P3_U2962) );
  AOI22_X1 U22014 ( .A1(n18848), .A2(n18822), .B1(n18943), .B2(n18789), .ZN(
        n18793) );
  AOI22_X1 U22015 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18791), .B1(
        n18944), .B2(n18790), .ZN(n18792) );
  OAI211_X1 U22016 ( .C1(n18881), .C2(n18853), .A(n18793), .B(n18792), .ZN(
        P3_U2963) );
  NOR2_X2 U22017 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18827), .ZN(
        n18945) );
  NOR2_X1 U22018 ( .A1(n18855), .A2(n18794), .ZN(n18797) );
  NOR2_X1 U22019 ( .A1(n18945), .A2(n18883), .ZN(n18856) );
  INV_X1 U22020 ( .A(n18856), .ZN(n18795) );
  AOI21_X1 U22021 ( .B1(n18797), .B2(n18796), .A(n18795), .ZN(n18799) );
  NOR2_X1 U22022 ( .A1(n19023), .A2(n18856), .ZN(n18821) );
  AOI22_X1 U22023 ( .A1(n18897), .A2(n18849), .B1(n18894), .B2(n18821), .ZN(
        n18801) );
  AOI22_X1 U22024 ( .A1(n18945), .A2(n18896), .B1(n18895), .B2(n18822), .ZN(
        n18800) );
  OAI211_X1 U22025 ( .C1(n18826), .C2(n18802), .A(n18801), .B(n18800), .ZN(
        P3_U2964) );
  AOI22_X1 U22026 ( .A1(n18803), .A2(n18849), .B1(n18901), .B2(n18821), .ZN(
        n18805) );
  AOI22_X1 U22027 ( .A1(n18945), .A2(n18903), .B1(n18902), .B2(n18822), .ZN(
        n18804) );
  OAI211_X1 U22028 ( .C1(n18826), .C2(n18806), .A(n18805), .B(n18804), .ZN(
        P3_U2965) );
  AOI22_X1 U22029 ( .A1(n18833), .A2(n18849), .B1(n18907), .B2(n18821), .ZN(
        n18808) );
  AOI22_X1 U22030 ( .A1(n18945), .A2(n18909), .B1(n18908), .B2(n18822), .ZN(
        n18807) );
  OAI211_X1 U22031 ( .C1(n18826), .C2(n18809), .A(n18808), .B(n18807), .ZN(
        P3_U2966) );
  AOI22_X1 U22032 ( .A1(n18916), .A2(n18849), .B1(n18913), .B2(n18821), .ZN(
        n18811) );
  AOI22_X1 U22033 ( .A1(n18945), .A2(n18915), .B1(n18914), .B2(n18822), .ZN(
        n18810) );
  OAI211_X1 U22034 ( .C1(n18826), .C2(n18812), .A(n18811), .B(n18810), .ZN(
        P3_U2967) );
  AOI22_X1 U22035 ( .A1(n18921), .A2(n18822), .B1(n18920), .B2(n18821), .ZN(
        n18814) );
  INV_X1 U22036 ( .A(n18826), .ZN(n18817) );
  AOI22_X1 U22037 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18817), .B1(
        n18922), .B2(n18849), .ZN(n18813) );
  OAI211_X1 U22038 ( .C1(n18888), .C2(n18925), .A(n18814), .B(n18813), .ZN(
        P3_U2968) );
  AOI22_X1 U22039 ( .A1(n18927), .A2(n18822), .B1(n18926), .B2(n18821), .ZN(
        n18816) );
  AOI22_X1 U22040 ( .A1(n18945), .A2(n18928), .B1(n18929), .B2(n18849), .ZN(
        n18815) );
  OAI211_X1 U22041 ( .C1(n18826), .C2(n9878), .A(n18816), .B(n18815), .ZN(
        P3_U2969) );
  AOI22_X1 U22042 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18817), .B1(
        n18934), .B2(n18821), .ZN(n18819) );
  AOI22_X1 U22043 ( .A1(n18945), .A2(n18876), .B1(n18936), .B2(n18849), .ZN(
        n18818) );
  OAI211_X1 U22044 ( .C1(n18880), .C2(n18820), .A(n18819), .B(n18818), .ZN(
        P3_U2970) );
  AOI22_X1 U22045 ( .A1(n18848), .A2(n18849), .B1(n18943), .B2(n18821), .ZN(
        n18824) );
  AOI22_X1 U22046 ( .A1(n18945), .A2(n18947), .B1(n18944), .B2(n18822), .ZN(
        n18823) );
  OAI211_X1 U22047 ( .C1(n18826), .C2(n18825), .A(n18824), .B(n18823), .ZN(
        P3_U2971) );
  NOR2_X1 U22048 ( .A1(n19023), .A2(n18827), .ZN(n18847) );
  AOI22_X1 U22049 ( .A1(n18883), .A2(n18897), .B1(n18894), .B2(n18847), .ZN(
        n18830) );
  AOI22_X1 U22050 ( .A1(n18891), .A2(n18828), .B1(n18890), .B2(n18889), .ZN(
        n18850) );
  AOI22_X1 U22051 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18850), .B1(
        n18937), .B2(n18896), .ZN(n18829) );
  OAI211_X1 U22052 ( .C1(n18861), .C2(n18842), .A(n18830), .B(n18829), .ZN(
        P3_U2972) );
  AOI22_X1 U22053 ( .A1(n18901), .A2(n18847), .B1(n18902), .B2(n18849), .ZN(
        n18832) );
  AOI22_X1 U22054 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18850), .B1(
        n18937), .B2(n18903), .ZN(n18831) );
  OAI211_X1 U22055 ( .C1(n18881), .C2(n18906), .A(n18832), .B(n18831), .ZN(
        P3_U2973) );
  AOI22_X1 U22056 ( .A1(n18883), .A2(n18833), .B1(n18907), .B2(n18847), .ZN(
        n18835) );
  AOI22_X1 U22057 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18850), .B1(
        n18908), .B2(n18849), .ZN(n18834) );
  OAI211_X1 U22058 ( .C1(n18952), .C2(n18836), .A(n18835), .B(n18834), .ZN(
        P3_U2974) );
  AOI22_X1 U22059 ( .A1(n18883), .A2(n18916), .B1(n18913), .B2(n18847), .ZN(
        n18838) );
  AOI22_X1 U22060 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18850), .B1(
        n18914), .B2(n18849), .ZN(n18837) );
  OAI211_X1 U22061 ( .C1(n18952), .C2(n18839), .A(n18838), .B(n18837), .ZN(
        P3_U2975) );
  AOI22_X1 U22062 ( .A1(n18883), .A2(n18922), .B1(n18920), .B2(n18847), .ZN(
        n18841) );
  AOI22_X1 U22063 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18850), .B1(
        n18937), .B2(n18869), .ZN(n18840) );
  OAI211_X1 U22064 ( .C1(n18872), .C2(n18842), .A(n18841), .B(n18840), .ZN(
        P3_U2976) );
  AOI22_X1 U22065 ( .A1(n18927), .A2(n18849), .B1(n18926), .B2(n18847), .ZN(
        n18844) );
  AOI22_X1 U22066 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18850), .B1(
        n18937), .B2(n18928), .ZN(n18843) );
  OAI211_X1 U22067 ( .C1(n18881), .C2(n18875), .A(n18844), .B(n18843), .ZN(
        P3_U2977) );
  AOI22_X1 U22068 ( .A1(n18935), .A2(n18849), .B1(n18934), .B2(n18847), .ZN(
        n18846) );
  AOI22_X1 U22069 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18850), .B1(
        n18883), .B2(n18936), .ZN(n18845) );
  OAI211_X1 U22070 ( .C1(n18952), .C2(n18941), .A(n18846), .B(n18845), .ZN(
        P3_U2978) );
  AOI22_X1 U22071 ( .A1(n18883), .A2(n18848), .B1(n18943), .B2(n18847), .ZN(
        n18852) );
  AOI22_X1 U22072 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18850), .B1(
        n18944), .B2(n18849), .ZN(n18851) );
  OAI211_X1 U22073 ( .C1(n18952), .C2(n18853), .A(n18852), .B(n18851), .ZN(
        P3_U2979) );
  NOR2_X1 U22074 ( .A1(n19023), .A2(n18854), .ZN(n18882) );
  AOI22_X1 U22075 ( .A1(n18945), .A2(n18897), .B1(n18894), .B2(n18882), .ZN(
        n18860) );
  AOI221_X1 U22076 ( .B1(n18856), .B2(n18952), .C1(n18855), .C2(n18952), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18858) );
  OAI21_X1 U22077 ( .B1(n18877), .B2(n18858), .A(n18857), .ZN(n18885) );
  AOI22_X1 U22078 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18885), .B1(
        n18877), .B2(n18896), .ZN(n18859) );
  OAI211_X1 U22079 ( .C1(n18881), .C2(n18861), .A(n18860), .B(n18859), .ZN(
        P3_U2980) );
  AOI22_X1 U22080 ( .A1(n18883), .A2(n18902), .B1(n18882), .B2(n18901), .ZN(
        n18863) );
  AOI22_X1 U22081 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18885), .B1(
        n18877), .B2(n18903), .ZN(n18862) );
  OAI211_X1 U22082 ( .C1(n18888), .C2(n18906), .A(n18863), .B(n18862), .ZN(
        P3_U2981) );
  AOI22_X1 U22083 ( .A1(n18883), .A2(n18908), .B1(n18882), .B2(n18907), .ZN(
        n18865) );
  AOI22_X1 U22084 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18885), .B1(
        n18877), .B2(n18909), .ZN(n18864) );
  OAI211_X1 U22085 ( .C1(n18888), .C2(n18912), .A(n18865), .B(n18864), .ZN(
        P3_U2982) );
  AOI22_X1 U22086 ( .A1(n18883), .A2(n18914), .B1(n18882), .B2(n18913), .ZN(
        n18867) );
  AOI22_X1 U22087 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18885), .B1(
        n18877), .B2(n18915), .ZN(n18866) );
  OAI211_X1 U22088 ( .C1(n18888), .C2(n18868), .A(n18867), .B(n18866), .ZN(
        P3_U2983) );
  AOI22_X1 U22089 ( .A1(n18945), .A2(n18922), .B1(n18882), .B2(n18920), .ZN(
        n18871) );
  AOI22_X1 U22090 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18885), .B1(
        n18877), .B2(n18869), .ZN(n18870) );
  OAI211_X1 U22091 ( .C1(n18881), .C2(n18872), .A(n18871), .B(n18870), .ZN(
        P3_U2984) );
  AOI22_X1 U22092 ( .A1(n18883), .A2(n18927), .B1(n18882), .B2(n18926), .ZN(
        n18874) );
  AOI22_X1 U22093 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18885), .B1(
        n18877), .B2(n18928), .ZN(n18873) );
  OAI211_X1 U22094 ( .C1(n18888), .C2(n18875), .A(n18874), .B(n18873), .ZN(
        P3_U2985) );
  AOI22_X1 U22095 ( .A1(n18945), .A2(n18936), .B1(n18882), .B2(n18934), .ZN(
        n18879) );
  AOI22_X1 U22096 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18885), .B1(
        n18877), .B2(n18876), .ZN(n18878) );
  OAI211_X1 U22097 ( .C1(n18881), .C2(n18880), .A(n18879), .B(n18878), .ZN(
        P3_U2986) );
  AOI22_X1 U22098 ( .A1(n18883), .A2(n18944), .B1(n18882), .B2(n18943), .ZN(
        n18887) );
  AOI22_X1 U22099 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18885), .B1(
        n18884), .B2(n18947), .ZN(n18886) );
  OAI211_X1 U22100 ( .C1(n18888), .C2(n18951), .A(n18887), .B(n18886), .ZN(
        P3_U2987) );
  AOI22_X1 U22101 ( .A1(n18891), .A2(n18890), .B1(n18889), .B2(n18892), .ZN(
        n18948) );
  INV_X1 U22102 ( .A(n18948), .ZN(n18932) );
  AND2_X1 U22103 ( .A1(n18893), .A2(n18892), .ZN(n18942) );
  AOI22_X1 U22104 ( .A1(n18945), .A2(n18895), .B1(n18894), .B2(n18942), .ZN(
        n18899) );
  AOI22_X1 U22105 ( .A1(n18937), .A2(n18897), .B1(n18896), .B2(n18946), .ZN(
        n18898) );
  OAI211_X1 U22106 ( .C1(n18900), .C2(n18932), .A(n18899), .B(n18898), .ZN(
        P3_U2988) );
  AOI22_X1 U22107 ( .A1(n18945), .A2(n18902), .B1(n18901), .B2(n18942), .ZN(
        n18905) );
  AOI22_X1 U22108 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18948), .B1(
        n18903), .B2(n18946), .ZN(n18904) );
  OAI211_X1 U22109 ( .C1(n18952), .C2(n18906), .A(n18905), .B(n18904), .ZN(
        P3_U2989) );
  AOI22_X1 U22110 ( .A1(n18945), .A2(n18908), .B1(n18907), .B2(n18942), .ZN(
        n18911) );
  AOI22_X1 U22111 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18948), .B1(
        n18909), .B2(n18946), .ZN(n18910) );
  OAI211_X1 U22112 ( .C1(n18952), .C2(n18912), .A(n18911), .B(n18910), .ZN(
        P3_U2990) );
  AOI22_X1 U22113 ( .A1(n18945), .A2(n18914), .B1(n18913), .B2(n18942), .ZN(
        n18918) );
  AOI22_X1 U22114 ( .A1(n18937), .A2(n18916), .B1(n18915), .B2(n18946), .ZN(
        n18917) );
  OAI211_X1 U22115 ( .C1(n18919), .C2(n18932), .A(n18918), .B(n18917), .ZN(
        P3_U2991) );
  AOI22_X1 U22116 ( .A1(n18945), .A2(n18921), .B1(n18920), .B2(n18942), .ZN(
        n18924) );
  AOI22_X1 U22117 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18948), .B1(
        n18937), .B2(n18922), .ZN(n18923) );
  OAI211_X1 U22118 ( .C1(n18925), .C2(n18940), .A(n18924), .B(n18923), .ZN(
        P3_U2992) );
  AOI22_X1 U22119 ( .A1(n18945), .A2(n18927), .B1(n18926), .B2(n18942), .ZN(
        n18931) );
  AOI22_X1 U22120 ( .A1(n18937), .A2(n18929), .B1(n18928), .B2(n18946), .ZN(
        n18930) );
  OAI211_X1 U22121 ( .C1(n18933), .C2(n18932), .A(n18931), .B(n18930), .ZN(
        P3_U2993) );
  AOI22_X1 U22122 ( .A1(n18945), .A2(n18935), .B1(n18934), .B2(n18942), .ZN(
        n18939) );
  AOI22_X1 U22123 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18948), .B1(
        n18937), .B2(n18936), .ZN(n18938) );
  OAI211_X1 U22124 ( .C1(n18941), .C2(n18940), .A(n18939), .B(n18938), .ZN(
        P3_U2994) );
  AOI22_X1 U22125 ( .A1(n18945), .A2(n18944), .B1(n18943), .B2(n18942), .ZN(
        n18950) );
  AOI22_X1 U22126 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18948), .B1(
        n18947), .B2(n18946), .ZN(n18949) );
  OAI211_X1 U22127 ( .C1(n18952), .C2(n18951), .A(n18950), .B(n18949), .ZN(
        P3_U2995) );
  NOR2_X1 U22128 ( .A1(n18964), .A2(n18953), .ZN(n18956) );
  OAI222_X1 U22129 ( .A1(n18959), .A2(n18958), .B1(n18957), .B2(n18956), .C1(
        n18955), .C2(n18954), .ZN(n19164) );
  OAI21_X1 U22130 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18960), .ZN(n18961) );
  OAI211_X1 U22131 ( .C1(n18963), .C2(n18987), .A(n18962), .B(n18961), .ZN(
        n19010) );
  NAND2_X1 U22132 ( .A1(n18990), .A2(n12924), .ZN(n18991) );
  NAND2_X1 U22133 ( .A1(n18974), .A2(n19139), .ZN(n18969) );
  AOI22_X1 U22134 ( .A1(n9904), .A2(n18991), .B1(n18964), .B2(n18969), .ZN(
        n18965) );
  NOR2_X1 U22135 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18965), .ZN(
        n19127) );
  AOI21_X1 U22136 ( .B1(n18968), .B2(n18967), .A(n18966), .ZN(n18975) );
  OAI21_X1 U22137 ( .B1(n18970), .B2(n18975), .A(n18969), .ZN(n18971) );
  AOI21_X1 U22138 ( .B1(n18977), .B2(n18972), .A(n18971), .ZN(n19128) );
  NAND2_X1 U22139 ( .A1(n18987), .A2(n19128), .ZN(n18973) );
  AOI22_X1 U22140 ( .A1(n18987), .A2(n19127), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18973), .ZN(n19008) );
  INV_X1 U22141 ( .A(n18987), .ZN(n18999) );
  AND2_X1 U22142 ( .A1(n18974), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n18986) );
  OAI21_X1 U22143 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18976), .A(
        n18975), .ZN(n18985) );
  OAI211_X1 U22144 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n18978), .B(n18977), .ZN(
        n18982) );
  NOR2_X1 U22145 ( .A1(n18988), .A2(n12924), .ZN(n18980) );
  OAI211_X1 U22146 ( .C1(n18980), .C2(n18979), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n19139), .ZN(n18981) );
  OAI211_X1 U22147 ( .C1(n19136), .C2(n18983), .A(n18982), .B(n18981), .ZN(
        n18984) );
  AOI21_X1 U22148 ( .B1(n18986), .B2(n18985), .A(n18984), .ZN(n19133) );
  AOI22_X1 U22149 ( .A1(n18999), .A2(n19139), .B1(n19133), .B2(n18987), .ZN(
        n19003) );
  AND2_X1 U22150 ( .A1(n18989), .A2(n18988), .ZN(n18994) );
  AOI22_X1 U22151 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18990), .B1(
        n18994), .B2(n12924), .ZN(n19148) );
  INV_X1 U22152 ( .A(n18991), .ZN(n18992) );
  OAI22_X1 U22153 ( .A1(n18994), .A2(n18993), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18992), .ZN(n19144) );
  AOI222_X1 U22154 ( .A1(n19148), .A2(n19144), .B1(n19148), .B2(n18996), .C1(
        n19144), .C2(n18995), .ZN(n18998) );
  OAI21_X1 U22155 ( .B1(n18999), .B2(n18998), .A(n18997), .ZN(n19002) );
  AND2_X1 U22156 ( .A1(n19003), .A2(n19002), .ZN(n19000) );
  OAI221_X1 U22157 ( .B1(n19003), .B2(n19002), .C1(n19001), .C2(n19000), .A(
        n19005), .ZN(n19007) );
  AOI21_X1 U22158 ( .B1(n19005), .B2(n19004), .A(n19003), .ZN(n19006) );
  AOI222_X1 U22159 ( .A1(n19008), .A2(n19007), .B1(n19008), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n19007), .C2(n19006), .ZN(
        n19009) );
  NOR4_X1 U22160 ( .A1(n19011), .A2(n19164), .A3(n19010), .A4(n19009), .ZN(
        n19021) );
  NOR2_X1 U22161 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19177) );
  AOI22_X1 U22162 ( .A1(n19147), .A2(n19177), .B1(n19172), .B2(n19166), .ZN(
        n19012) );
  INV_X1 U22163 ( .A(n19012), .ZN(n19017) );
  OAI211_X1 U22164 ( .C1(n19014), .C2(n19013), .A(n19169), .B(n19021), .ZN(
        n19124) );
  NAND2_X1 U22165 ( .A1(n19172), .A2(n19183), .ZN(n19022) );
  NAND2_X1 U22166 ( .A1(n19124), .A2(n19022), .ZN(n19024) );
  NOR2_X1 U22167 ( .A1(n19015), .A2(n19024), .ZN(n19016) );
  MUX2_X1 U22168 ( .A(n19017), .B(n19016), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n19019) );
  OAI211_X1 U22169 ( .C1(n19021), .C2(n19020), .A(n19019), .B(n19018), .ZN(
        P3_U2996) );
  NAND2_X1 U22170 ( .A1(n19172), .A2(n19166), .ZN(n19027) );
  OR3_X1 U22171 ( .A1(n19134), .A2(n19174), .A3(n19022), .ZN(n19029) );
  NAND4_X1 U22172 ( .A1(n19028), .A2(n19027), .A3(n19029), .A4(n19026), .ZN(
        P3_U2997) );
  INV_X1 U22173 ( .A(n19177), .ZN(n19031) );
  AND4_X1 U22174 ( .A1(n19031), .A2(n19030), .A3(n19029), .A4(n19123), .ZN(
        P3_U2998) );
  AND2_X1 U22175 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19119), .ZN(
        P3_U2999) );
  AND2_X1 U22176 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19119), .ZN(
        P3_U3000) );
  AND2_X1 U22177 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19119), .ZN(
        P3_U3001) );
  AND2_X1 U22178 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19119), .ZN(
        P3_U3002) );
  AND2_X1 U22179 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19119), .ZN(
        P3_U3003) );
  AND2_X1 U22180 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19119), .ZN(
        P3_U3004) );
  AND2_X1 U22181 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19119), .ZN(
        P3_U3005) );
  AND2_X1 U22182 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19119), .ZN(
        P3_U3006) );
  AND2_X1 U22183 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19119), .ZN(
        P3_U3007) );
  AND2_X1 U22184 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19119), .ZN(
        P3_U3008) );
  AND2_X1 U22185 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19119), .ZN(
        P3_U3009) );
  AND2_X1 U22186 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19119), .ZN(
        P3_U3010) );
  AND2_X1 U22187 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19119), .ZN(
        P3_U3011) );
  AND2_X1 U22188 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19119), .ZN(
        P3_U3012) );
  AND2_X1 U22189 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19119), .ZN(
        P3_U3013) );
  AND2_X1 U22190 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19119), .ZN(
        P3_U3014) );
  AND2_X1 U22191 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19119), .ZN(
        P3_U3015) );
  AND2_X1 U22192 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19119), .ZN(
        P3_U3016) );
  AND2_X1 U22193 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19119), .ZN(
        P3_U3017) );
  AND2_X1 U22194 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19119), .ZN(
        P3_U3018) );
  AND2_X1 U22195 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19119), .ZN(
        P3_U3019) );
  AND2_X1 U22196 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19119), .ZN(
        P3_U3020) );
  AND2_X1 U22197 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19119), .ZN(P3_U3021) );
  AND2_X1 U22198 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19119), .ZN(P3_U3022) );
  AND2_X1 U22199 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19119), .ZN(P3_U3023) );
  AND2_X1 U22200 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19119), .ZN(P3_U3024) );
  AND2_X1 U22201 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19119), .ZN(P3_U3025) );
  AND2_X1 U22202 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19119), .ZN(P3_U3026) );
  AND2_X1 U22203 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19119), .ZN(P3_U3027) );
  AND2_X1 U22204 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19119), .ZN(P3_U3028) );
  OAI21_X1 U22205 ( .B1(n19032), .B2(n20819), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19033) );
  AOI22_X1 U22206 ( .A1(n19045), .A2(n19047), .B1(n19181), .B2(n19033), .ZN(
        n19035) );
  INV_X1 U22207 ( .A(NA), .ZN(n21013) );
  OR3_X1 U22208 ( .A1(n21013), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n19034) );
  OAI211_X1 U22209 ( .C1(n19165), .C2(n19036), .A(n19035), .B(n19034), .ZN(
        P3_U3029) );
  INV_X1 U22210 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19179) );
  NOR2_X1 U22211 ( .A1(n19047), .A2(n20819), .ZN(n19043) );
  OAI22_X1 U22212 ( .A1(n19179), .A2(n19043), .B1(n20819), .B2(n19036), .ZN(
        n19037) );
  INV_X1 U22213 ( .A(n19037), .ZN(n19039) );
  NAND2_X1 U22214 ( .A1(n19172), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19041) );
  OAI211_X1 U22215 ( .C1(n19039), .C2(n19045), .A(n19041), .B(n19038), .ZN(
        P3_U3030) );
  INV_X1 U22216 ( .A(n19041), .ZN(n19040) );
  AOI221_X1 U22217 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n19045), .C1(n21013), 
        .C2(n19045), .A(n19040), .ZN(n19046) );
  OAI22_X1 U22218 ( .A1(NA), .A2(n19041), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19042) );
  OAI22_X1 U22219 ( .A1(n19043), .A2(n19042), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19044) );
  OAI22_X1 U22220 ( .A1(n19046), .A2(n19047), .B1(n19045), .B2(n19044), .ZN(
        P3_U3031) );
  OAI222_X1 U22221 ( .A1(n19153), .A2(n19109), .B1(n19048), .B2(n19116), .C1(
        n19049), .C2(n19101), .ZN(P3_U3032) );
  INV_X1 U22222 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19051) );
  OAI222_X1 U22223 ( .A1(n19101), .A2(n19051), .B1(n19050), .B2(n19116), .C1(
        n19049), .C2(n19109), .ZN(P3_U3033) );
  OAI222_X1 U22224 ( .A1(n19101), .A2(n19053), .B1(n19052), .B2(n19116), .C1(
        n19051), .C2(n19109), .ZN(P3_U3034) );
  OAI222_X1 U22225 ( .A1(n19101), .A2(n19056), .B1(n19054), .B2(n19116), .C1(
        n19053), .C2(n19109), .ZN(P3_U3035) );
  OAI222_X1 U22226 ( .A1(n19056), .A2(n19109), .B1(n19055), .B2(n19116), .C1(
        n19057), .C2(n19101), .ZN(P3_U3036) );
  OAI222_X1 U22227 ( .A1(n19101), .A2(n19059), .B1(n19058), .B2(n19116), .C1(
        n19057), .C2(n19109), .ZN(P3_U3037) );
  OAI222_X1 U22228 ( .A1(n19101), .A2(n19061), .B1(n19060), .B2(n19116), .C1(
        n19059), .C2(n19109), .ZN(P3_U3038) );
  OAI222_X1 U22229 ( .A1(n19101), .A2(n19063), .B1(n19062), .B2(n19116), .C1(
        n19061), .C2(n19109), .ZN(P3_U3039) );
  OAI222_X1 U22230 ( .A1(n19101), .A2(n19065), .B1(n19064), .B2(n19116), .C1(
        n19063), .C2(n19109), .ZN(P3_U3040) );
  OAI222_X1 U22231 ( .A1(n19101), .A2(n19067), .B1(n19066), .B2(n19116), .C1(
        n19065), .C2(n19109), .ZN(P3_U3041) );
  OAI222_X1 U22232 ( .A1(n19101), .A2(n19069), .B1(n19068), .B2(n19116), .C1(
        n19067), .C2(n19109), .ZN(P3_U3042) );
  OAI222_X1 U22233 ( .A1(n19101), .A2(n19071), .B1(n19070), .B2(n19116), .C1(
        n19069), .C2(n19109), .ZN(P3_U3043) );
  OAI222_X1 U22234 ( .A1(n19101), .A2(n19074), .B1(n19072), .B2(n19116), .C1(
        n19071), .C2(n19109), .ZN(P3_U3044) );
  OAI222_X1 U22235 ( .A1(n19074), .A2(n19109), .B1(n19073), .B2(n19116), .C1(
        n19075), .C2(n19101), .ZN(P3_U3045) );
  OAI222_X1 U22236 ( .A1(n19101), .A2(n19077), .B1(n19076), .B2(n19116), .C1(
        n19075), .C2(n19109), .ZN(P3_U3046) );
  OAI222_X1 U22237 ( .A1(n19101), .A2(n19079), .B1(n19078), .B2(n19116), .C1(
        n19077), .C2(n19109), .ZN(P3_U3047) );
  OAI222_X1 U22238 ( .A1(n19101), .A2(n19081), .B1(n19080), .B2(n19116), .C1(
        n19079), .C2(n19109), .ZN(P3_U3048) );
  OAI222_X1 U22239 ( .A1(n19101), .A2(n19084), .B1(n19082), .B2(n19116), .C1(
        n19081), .C2(n19109), .ZN(P3_U3049) );
  OAI222_X1 U22240 ( .A1(n19084), .A2(n19109), .B1(n19083), .B2(n19116), .C1(
        n19085), .C2(n19101), .ZN(P3_U3050) );
  OAI222_X1 U22241 ( .A1(n19101), .A2(n19088), .B1(n19086), .B2(n19116), .C1(
        n19085), .C2(n19109), .ZN(P3_U3051) );
  OAI222_X1 U22242 ( .A1(n19088), .A2(n19109), .B1(n19087), .B2(n19116), .C1(
        n19089), .C2(n19101), .ZN(P3_U3052) );
  OAI222_X1 U22243 ( .A1(n19101), .A2(n19092), .B1(n19090), .B2(n19116), .C1(
        n19089), .C2(n19109), .ZN(P3_U3053) );
  OAI222_X1 U22244 ( .A1(n19092), .A2(n19109), .B1(n19091), .B2(n19116), .C1(
        n19093), .C2(n19101), .ZN(P3_U3054) );
  OAI222_X1 U22245 ( .A1(n19101), .A2(n19095), .B1(n19094), .B2(n19116), .C1(
        n19093), .C2(n19109), .ZN(P3_U3055) );
  OAI222_X1 U22246 ( .A1(n19101), .A2(n19097), .B1(n19096), .B2(n19116), .C1(
        n19095), .C2(n19109), .ZN(P3_U3056) );
  OAI222_X1 U22247 ( .A1(n19101), .A2(n19099), .B1(n19098), .B2(n19116), .C1(
        n19097), .C2(n19109), .ZN(P3_U3057) );
  OAI222_X1 U22248 ( .A1(n19101), .A2(n19103), .B1(n19100), .B2(n19116), .C1(
        n19099), .C2(n19109), .ZN(P3_U3058) );
  OAI222_X1 U22249 ( .A1(n19103), .A2(n19109), .B1(n19102), .B2(n19116), .C1(
        n19104), .C2(n19101), .ZN(P3_U3059) );
  OAI222_X1 U22250 ( .A1(n19101), .A2(n19108), .B1(n19105), .B2(n19116), .C1(
        n19104), .C2(n19109), .ZN(P3_U3060) );
  INV_X1 U22251 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19107) );
  OAI222_X1 U22252 ( .A1(n19109), .A2(n19108), .B1(n19107), .B2(n19116), .C1(
        n19106), .C2(n19101), .ZN(P3_U3061) );
  INV_X1 U22253 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n19110) );
  AOI22_X1 U22254 ( .A1(n19116), .A2(n19111), .B1(n19110), .B2(n19181), .ZN(
        P3_U3274) );
  INV_X1 U22255 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19155) );
  INV_X1 U22256 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n19112) );
  AOI22_X1 U22257 ( .A1(n19116), .A2(n19155), .B1(n19112), .B2(n19181), .ZN(
        P3_U3275) );
  INV_X1 U22258 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n19113) );
  AOI22_X1 U22259 ( .A1(n19116), .A2(n19114), .B1(n19113), .B2(n19181), .ZN(
        P3_U3276) );
  INV_X1 U22260 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19161) );
  INV_X1 U22261 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n19115) );
  AOI22_X1 U22262 ( .A1(n19116), .A2(n19161), .B1(n19115), .B2(n19181), .ZN(
        P3_U3277) );
  INV_X1 U22263 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19118) );
  INV_X1 U22264 ( .A(n19120), .ZN(n19117) );
  AOI21_X1 U22265 ( .B1(n19119), .B2(n19118), .A(n19117), .ZN(P3_U3280) );
  OAI21_X1 U22266 ( .B1(n19122), .B2(n19121), .A(n19120), .ZN(P3_U3281) );
  OAI221_X1 U22267 ( .B1(n19125), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19125), 
        .C2(n19124), .A(n19123), .ZN(P3_U3282) );
  AOI22_X1 U22268 ( .A1(n19184), .A2(n19127), .B1(n19147), .B2(n19126), .ZN(
        n19132) );
  INV_X1 U22269 ( .A(n19128), .ZN(n19129) );
  AOI21_X1 U22270 ( .B1(n19184), .B2(n19129), .A(n19152), .ZN(n19131) );
  OAI22_X1 U22271 ( .A1(n19152), .A2(n19132), .B1(n19131), .B2(n19130), .ZN(
        P3_U3285) );
  INV_X1 U22272 ( .A(n19133), .ZN(n19137) );
  NOR2_X1 U22273 ( .A1(n19134), .A2(n19149), .ZN(n19141) );
  AOI22_X1 U22274 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13031), .B2(n19135), .ZN(
        n19140) );
  AOI222_X1 U22275 ( .A1(n19137), .A2(n19184), .B1(n19141), .B2(n19140), .C1(
        n19147), .C2(n19136), .ZN(n19138) );
  AOI22_X1 U22276 ( .A1(n19152), .A2(n19139), .B1(n19138), .B2(n19150), .ZN(
        P3_U3288) );
  INV_X1 U22277 ( .A(n19140), .ZN(n19142) );
  AOI222_X1 U22278 ( .A1(n19144), .A2(n19184), .B1(n19147), .B2(n19143), .C1(
        n19142), .C2(n19141), .ZN(n19145) );
  AOI22_X1 U22279 ( .A1(n19152), .A2(n19146), .B1(n19145), .B2(n19150), .ZN(
        P3_U3289) );
  AOI222_X1 U22280 ( .A1(n19149), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19184), 
        .B2(n19148), .C1(n12924), .C2(n19147), .ZN(n19151) );
  AOI22_X1 U22281 ( .A1(n19152), .A2(n12924), .B1(n19151), .B2(n19150), .ZN(
        P3_U3290) );
  AOI21_X1 U22282 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19154) );
  AOI22_X1 U22283 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19154), .B2(n19153), .ZN(n19156) );
  AOI22_X1 U22284 ( .A1(n19157), .A2(n19156), .B1(n19155), .B2(n19160), .ZN(
        P3_U3292) );
  NOR2_X1 U22285 ( .A1(n19160), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19158) );
  AOI22_X1 U22286 ( .A1(n19161), .A2(n19160), .B1(n19159), .B2(n19158), .ZN(
        P3_U3293) );
  INV_X1 U22287 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19162) );
  AOI22_X1 U22288 ( .A1(n19116), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19162), 
        .B2(n19181), .ZN(P3_U3294) );
  MUX2_X1 U22289 ( .A(P3_MORE_REG_SCAN_IN), .B(n19164), .S(n19163), .Z(
        P3_U3295) );
  AOI21_X1 U22290 ( .B1(n19166), .B2(n19165), .A(n19186), .ZN(n19167) );
  OAI21_X1 U22291 ( .B1(n19169), .B2(n19168), .A(n19167), .ZN(n19180) );
  OAI21_X1 U22292 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n19171), .A(n19170), 
        .ZN(n19173) );
  AOI211_X1 U22293 ( .C1(n19185), .C2(n19173), .A(n19172), .B(n19183), .ZN(
        n19175) );
  NOR2_X1 U22294 ( .A1(n19175), .A2(n19174), .ZN(n19176) );
  OAI21_X1 U22295 ( .B1(n19177), .B2(n19176), .A(n19180), .ZN(n19178) );
  OAI21_X1 U22296 ( .B1(n19180), .B2(n19179), .A(n19178), .ZN(P3_U3296) );
  INV_X1 U22297 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19189) );
  INV_X1 U22298 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n19182) );
  AOI22_X1 U22299 ( .A1(n19116), .A2(n19189), .B1(n19182), .B2(n19181), .ZN(
        P3_U3297) );
  AOI21_X1 U22300 ( .B1(n19184), .B2(n19183), .A(n19186), .ZN(n19190) );
  INV_X1 U22301 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n19187) );
  AOI22_X1 U22302 ( .A1(n19190), .A2(n19187), .B1(n19186), .B2(n19185), .ZN(
        P3_U3298) );
  AOI21_X1 U22303 ( .B1(n19190), .B2(n19189), .A(n19188), .ZN(P3_U3299) );
  INV_X1 U22304 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n19192) );
  INV_X1 U22305 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20090) );
  NAND2_X1 U22306 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20090), .ZN(n20081) );
  NOR2_X1 U22307 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n20078) );
  INV_X1 U22308 ( .A(n20078), .ZN(n19191) );
  OAI21_X1 U22309 ( .B1(n20074), .B2(n20081), .A(n19191), .ZN(n20146) );
  OAI21_X1 U22310 ( .B1(n20074), .B2(n19192), .A(n20073), .ZN(P2_U2815) );
  INV_X1 U22311 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19194) );
  OAI22_X1 U22312 ( .A1(n20198), .A2(n19194), .B1(n20201), .B2(n19193), .ZN(
        P2_U2816) );
  AOI22_X1 U22313 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(n20213), .B1(n19196), .B2(
        n20074), .ZN(n19195) );
  OAI21_X1 U22314 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n20213), .A(n19195), 
        .ZN(P2_U2817) );
  OAI21_X1 U22315 ( .B1(n19196), .B2(BS16), .A(n20146), .ZN(n20144) );
  OAI21_X1 U22316 ( .B1(n20146), .B2(n19595), .A(n20144), .ZN(P2_U2818) );
  NOR4_X1 U22317 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19200) );
  NOR4_X1 U22318 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19199) );
  NOR4_X1 U22319 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19198) );
  NOR4_X1 U22320 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19197) );
  NAND4_X1 U22321 ( .A1(n19200), .A2(n19199), .A3(n19198), .A4(n19197), .ZN(
        n19206) );
  NOR4_X1 U22322 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19204) );
  AOI211_X1 U22323 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19203) );
  NOR4_X1 U22324 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19202) );
  NOR4_X1 U22325 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19201) );
  NAND4_X1 U22326 ( .A1(n19204), .A2(n19203), .A3(n19202), .A4(n19201), .ZN(
        n19205) );
  NOR2_X1 U22327 ( .A1(n19206), .A2(n19205), .ZN(n19213) );
  INV_X1 U22328 ( .A(n19213), .ZN(n19212) );
  NOR2_X1 U22329 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19212), .ZN(n19207) );
  INV_X1 U22330 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20142) );
  AOI22_X1 U22331 ( .A1(n19207), .A2(n10313), .B1(n19212), .B2(n20142), .ZN(
        P2_U2820) );
  OR3_X1 U22332 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19211) );
  INV_X1 U22333 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20140) );
  AOI22_X1 U22334 ( .A1(n19207), .A2(n19211), .B1(n19212), .B2(n20140), .ZN(
        P2_U2821) );
  INV_X1 U22335 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20145) );
  NAND2_X1 U22336 ( .A1(n19207), .A2(n20145), .ZN(n19210) );
  OAI21_X1 U22337 ( .B1(n10313), .B2(n10673), .A(n19213), .ZN(n19208) );
  OAI21_X1 U22338 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19213), .A(n19208), 
        .ZN(n19209) );
  OAI221_X1 U22339 ( .B1(n19210), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19210), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19209), .ZN(P2_U2822) );
  INV_X1 U22340 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20138) );
  OAI221_X1 U22341 ( .B1(n19213), .B2(n20138), .C1(n19212), .C2(n19211), .A(
        n19210), .ZN(P2_U2823) );
  NOR2_X1 U22342 ( .A1(n19214), .A2(n19354), .ZN(n19220) );
  INV_X1 U22343 ( .A(n19215), .ZN(n19218) );
  AOI22_X1 U22344 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n19361), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19366), .ZN(n19217) );
  NAND2_X1 U22345 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19360), .ZN(
        n19216) );
  OAI211_X1 U22346 ( .C1(n19381), .C2(n19218), .A(n19217), .B(n19216), .ZN(
        n19219) );
  AOI211_X1 U22347 ( .C1(n19221), .C2(n19385), .A(n19220), .B(n19219), .ZN(
        n19225) );
  OAI211_X1 U22348 ( .C1(n19223), .C2(n19226), .A(n19342), .B(n19222), .ZN(
        n19224) );
  OAI211_X1 U22349 ( .C1(n19390), .C2(n19226), .A(n19225), .B(n19224), .ZN(
        P2_U2835) );
  NAND2_X1 U22350 ( .A1(n13243), .A2(n19227), .ZN(n19228) );
  XOR2_X1 U22351 ( .A(n19229), .B(n19228), .Z(n19240) );
  OAI222_X1 U22352 ( .A1(n19362), .A2(n19232), .B1(n19382), .B2(n19231), .C1(
        n19391), .C2(n19230), .ZN(n19233) );
  AOI211_X1 U22353 ( .C1(P2_REIP_REG_19__SCAN_IN), .C2(n19366), .A(n19517), 
        .B(n19233), .ZN(n19239) );
  INV_X1 U22354 ( .A(n19234), .ZN(n19235) );
  OAI22_X1 U22355 ( .A1(n19236), .A2(n19354), .B1(n19235), .B2(n19381), .ZN(
        n19237) );
  INV_X1 U22356 ( .A(n19237), .ZN(n19238) );
  OAI211_X1 U22357 ( .C1(n20071), .C2(n19240), .A(n19239), .B(n19238), .ZN(
        P2_U2836) );
  OAI21_X1 U22358 ( .B1(n20112), .B2(n19387), .A(n19350), .ZN(n19244) );
  OAI22_X1 U22359 ( .A1(n19242), .A2(n19362), .B1(n19241), .B2(n19382), .ZN(
        n19243) );
  AOI211_X1 U22360 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19360), .A(
        n19244), .B(n19243), .ZN(n19250) );
  NOR2_X1 U22361 ( .A1(n19372), .A2(n19245), .ZN(n19257) );
  XNOR2_X1 U22362 ( .A(n19257), .B(n19246), .ZN(n19248) );
  AOI22_X1 U22363 ( .A1(n19248), .A2(n19342), .B1(n19247), .B2(n19389), .ZN(
        n19249) );
  OAI211_X1 U22364 ( .C1(n19251), .C2(n19381), .A(n19250), .B(n19249), .ZN(
        P2_U2837) );
  AOI22_X1 U22365 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19360), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19366), .ZN(n19263) );
  OAI22_X1 U22366 ( .A1(n19252), .A2(n19362), .B1(n19258), .B2(n19390), .ZN(
        n19253) );
  AOI211_X1 U22367 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19361), .A(n19517), .B(
        n19253), .ZN(n19262) );
  AOI22_X1 U22368 ( .A1(n19255), .A2(n19389), .B1(n19254), .B2(n19305), .ZN(
        n19261) );
  INV_X1 U22369 ( .A(n19256), .ZN(n19259) );
  OAI211_X1 U22370 ( .C1(n19259), .C2(n19258), .A(n19342), .B(n19257), .ZN(
        n19260) );
  NAND4_X1 U22371 ( .A1(n19263), .A2(n19262), .A3(n19261), .A4(n19260), .ZN(
        P2_U2838) );
  OAI21_X1 U22372 ( .B1(n12181), .B2(n19382), .A(n19350), .ZN(n19267) );
  OAI22_X1 U22373 ( .A1(n19265), .A2(n19362), .B1(n19264), .B2(n19391), .ZN(
        n19266) );
  AOI211_X1 U22374 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n19366), .A(n19267), 
        .B(n19266), .ZN(n19273) );
  NOR2_X1 U22375 ( .A1(n19372), .A2(n19268), .ZN(n19270) );
  XNOR2_X1 U22376 ( .A(n19270), .B(n19269), .ZN(n19271) );
  AOI22_X1 U22377 ( .A1(n19271), .A2(n19342), .B1(n19400), .B2(n19389), .ZN(
        n19272) );
  OAI211_X1 U22378 ( .C1(n19274), .C2(n19381), .A(n19273), .B(n19272), .ZN(
        P2_U2839) );
  NAND2_X1 U22379 ( .A1(n19299), .A2(n19275), .ZN(n19276) );
  XOR2_X1 U22380 ( .A(n19277), .B(n19276), .Z(n19287) );
  OAI21_X1 U22381 ( .B1(n19278), .B2(n19382), .A(n19324), .ZN(n19282) );
  OAI22_X1 U22382 ( .A1(n19280), .A2(n19362), .B1(n19279), .B2(n19391), .ZN(
        n19281) );
  AOI211_X1 U22383 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n19366), .A(n19282), 
        .B(n19281), .ZN(n19286) );
  AOI22_X1 U22384 ( .A1(n19284), .A2(n19389), .B1(n19305), .B2(n19283), .ZN(
        n19285) );
  OAI211_X1 U22385 ( .C1(n20071), .C2(n19287), .A(n19286), .B(n19285), .ZN(
        P2_U2840) );
  AOI22_X1 U22386 ( .A1(n19361), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19360), .ZN(n19288) );
  OAI21_X1 U22387 ( .B1(n19289), .B2(n19362), .A(n19288), .ZN(n19290) );
  AOI211_X1 U22388 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19366), .A(n19517), 
        .B(n19290), .ZN(n19297) );
  NOR2_X1 U22389 ( .A1(n19372), .A2(n19291), .ZN(n19293) );
  XNOR2_X1 U22390 ( .A(n19293), .B(n19292), .ZN(n19295) );
  AOI22_X1 U22391 ( .A1(n19295), .A2(n19342), .B1(n19294), .B2(n19389), .ZN(
        n19296) );
  OAI211_X1 U22392 ( .C1(n19424), .C2(n19381), .A(n19297), .B(n19296), .ZN(
        P2_U2841) );
  NAND2_X1 U22393 ( .A1(n19299), .A2(n19298), .ZN(n19300) );
  XOR2_X1 U22394 ( .A(n19301), .B(n19300), .Z(n19309) );
  AOI22_X1 U22395 ( .A1(n19302), .A2(n19385), .B1(n19360), .B2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n19303) );
  OAI211_X1 U22396 ( .C1(n10790), .C2(n19382), .A(n19303), .B(n19324), .ZN(
        n19304) );
  AOI21_X1 U22397 ( .B1(P2_REIP_REG_13__SCAN_IN), .B2(n19366), .A(n19304), 
        .ZN(n19308) );
  AOI22_X1 U22398 ( .A1(n19306), .A2(n19389), .B1(n19305), .B2(n19425), .ZN(
        n19307) );
  OAI211_X1 U22399 ( .C1(n20071), .C2(n19309), .A(n19308), .B(n19307), .ZN(
        P2_U2842) );
  AOI222_X1 U22400 ( .A1(n19310), .A2(n19385), .B1(P2_EBX_REG_12__SCAN_IN), 
        .B2(n19361), .C1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n19360), .ZN(
        n19311) );
  INV_X1 U22401 ( .A(n19311), .ZN(n19312) );
  AOI211_X1 U22402 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19366), .A(n19517), 
        .B(n19312), .ZN(n19319) );
  NOR2_X1 U22403 ( .A1(n19372), .A2(n19313), .ZN(n19315) );
  XNOR2_X1 U22404 ( .A(n19315), .B(n19314), .ZN(n19317) );
  AOI22_X1 U22405 ( .A1(n19317), .A2(n19342), .B1(n19316), .B2(n19389), .ZN(
        n19318) );
  OAI211_X1 U22406 ( .C1(n19320), .C2(n19381), .A(n19319), .B(n19318), .ZN(
        P2_U2843) );
  INV_X1 U22407 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n19321) );
  OAI22_X1 U22408 ( .A1(n19322), .A2(n19362), .B1(n19321), .B2(n19391), .ZN(
        n19323) );
  INV_X1 U22409 ( .A(n19323), .ZN(n19325) );
  OAI211_X1 U22410 ( .C1(n19410), .C2(n19382), .A(n19325), .B(n19324), .ZN(
        n19326) );
  AOI21_X1 U22411 ( .B1(P2_REIP_REG_10__SCAN_IN), .B2(n19366), .A(n19326), 
        .ZN(n19332) );
  NOR2_X1 U22412 ( .A1(n19372), .A2(n19327), .ZN(n19329) );
  XNOR2_X1 U22413 ( .A(n19329), .B(n19328), .ZN(n19330) );
  AOI22_X1 U22414 ( .A1(n19330), .A2(n19342), .B1(n19407), .B2(n19389), .ZN(
        n19331) );
  OAI211_X1 U22415 ( .C1(n19333), .C2(n19381), .A(n19332), .B(n19331), .ZN(
        P2_U2845) );
  OAI222_X1 U22416 ( .A1(n19336), .A2(n19362), .B1(n19382), .B2(n19335), .C1(
        n19334), .C2(n19391), .ZN(n19337) );
  AOI211_X1 U22417 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n19366), .A(n19517), .B(
        n19337), .ZN(n19345) );
  NOR2_X1 U22418 ( .A1(n19372), .A2(n19338), .ZN(n19340) );
  XNOR2_X1 U22419 ( .A(n19340), .B(n19339), .ZN(n19343) );
  AOI22_X1 U22420 ( .A1(n19343), .A2(n19342), .B1(n19389), .B2(n19341), .ZN(
        n19344) );
  OAI211_X1 U22421 ( .C1(n19381), .C2(n19436), .A(n19345), .B(n19344), .ZN(
        P2_U2847) );
  NAND2_X1 U22422 ( .A1(n13243), .A2(n19346), .ZN(n19348) );
  XOR2_X1 U22423 ( .A(n19348), .B(n19347), .Z(n19359) );
  AOI22_X1 U22424 ( .A1(n19349), .A2(n19385), .B1(n19366), .B2(
        P2_REIP_REG_7__SCAN_IN), .ZN(n19351) );
  OAI211_X1 U22425 ( .C1(n19352), .C2(n19382), .A(n19351), .B(n19350), .ZN(
        n19357) );
  OAI22_X1 U22426 ( .A1(n19355), .A2(n19381), .B1(n19354), .B2(n19353), .ZN(
        n19356) );
  AOI211_X1 U22427 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19360), .A(
        n19357), .B(n19356), .ZN(n19358) );
  OAI21_X1 U22428 ( .B1(n19359), .B2(n20071), .A(n19358), .ZN(P2_U2848) );
  AOI22_X1 U22429 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19361), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19360), .ZN(n19379) );
  INV_X1 U22430 ( .A(n19524), .ZN(n19364) );
  OAI22_X1 U22431 ( .A1(n19364), .A2(n19381), .B1(n19363), .B2(n19362), .ZN(
        n19365) );
  AOI211_X1 U22432 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19366), .A(n19517), .B(
        n19365), .ZN(n19378) );
  INV_X1 U22433 ( .A(n19367), .ZN(n19412) );
  NAND2_X1 U22434 ( .A1(n19369), .A2(n19368), .ZN(n19370) );
  AOI22_X1 U22435 ( .A1(n19412), .A2(n19393), .B1(n19389), .B2(n19523), .ZN(
        n19377) );
  INV_X1 U22436 ( .A(n19500), .ZN(n19375) );
  NOR2_X1 U22437 ( .A1(n19372), .A2(n19371), .ZN(n19374) );
  AOI21_X1 U22438 ( .B1(n19375), .B2(n19374), .A(n20071), .ZN(n19373) );
  OAI21_X1 U22439 ( .B1(n19375), .B2(n19374), .A(n19373), .ZN(n19376) );
  NAND4_X1 U22440 ( .A1(n19379), .A2(n19378), .A3(n19377), .A4(n19376), .ZN(
        P2_U2851) );
  OAI22_X1 U22441 ( .A1(n19382), .A2(n10858), .B1(n19381), .B2(n19380), .ZN(
        n19383) );
  AOI21_X1 U22442 ( .B1(n19385), .B2(n19384), .A(n19383), .ZN(n19386) );
  OAI21_X1 U22443 ( .B1(n10313), .B2(n19387), .A(n19386), .ZN(n19388) );
  AOI21_X1 U22444 ( .B1(n19513), .B2(n19389), .A(n19388), .ZN(n19396) );
  AOI21_X1 U22445 ( .B1(n19391), .B2(n19390), .A(n19515), .ZN(n19392) );
  AOI21_X1 U22446 ( .B1(n19394), .B2(n19393), .A(n19392), .ZN(n19395) );
  OAI211_X1 U22447 ( .C1(n19398), .C2(n19397), .A(n19396), .B(n19395), .ZN(
        P2_U2855) );
  INV_X1 U22448 ( .A(n19399), .ZN(n19401) );
  AOI22_X1 U22449 ( .A1(n19401), .A2(n19411), .B1(n19406), .B2(n19400), .ZN(
        n19402) );
  OAI21_X1 U22450 ( .B1(n19415), .B2(n12181), .A(n19402), .ZN(P2_U2871) );
  AOI21_X1 U22451 ( .B1(n19405), .B2(n19404), .A(n19403), .ZN(n19408) );
  AOI22_X1 U22452 ( .A1(n19408), .A2(n13923), .B1(n19407), .B2(n19406), .ZN(
        n19409) );
  OAI21_X1 U22453 ( .B1(n19415), .B2(n19410), .A(n19409), .ZN(P2_U2877) );
  AOI22_X1 U22454 ( .A1(n19412), .A2(n19411), .B1(n19415), .B2(n19523), .ZN(
        n19413) );
  OAI21_X1 U22455 ( .B1(n19415), .B2(n19414), .A(n19413), .ZN(P2_U2883) );
  AOI22_X1 U22456 ( .A1(n19418), .A2(BUF2_REG_31__SCAN_IN), .B1(n19417), .B2(
        n19416), .ZN(n19421) );
  AOI22_X1 U22457 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19419), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19432), .ZN(n19420) );
  NAND2_X1 U22458 ( .A1(n19421), .A2(n19420), .ZN(P2_U2888) );
  INV_X1 U22459 ( .A(n19422), .ZN(n19481) );
  AOI22_X1 U22460 ( .A1(n19434), .A2(n19481), .B1(n19432), .B2(
        P2_EAX_REG_14__SCAN_IN), .ZN(n19423) );
  OAI21_X1 U22461 ( .B1(n19437), .B2(n19424), .A(n19423), .ZN(P2_U2905) );
  INV_X1 U22462 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19450) );
  INV_X1 U22463 ( .A(n19437), .ZN(n19426) );
  AOI22_X1 U22464 ( .A1(n19426), .A2(n19425), .B1(n19434), .B2(n19479), .ZN(
        n19427) );
  OAI21_X1 U22465 ( .B1(n19428), .B2(n19450), .A(n19427), .ZN(P2_U2906) );
  AOI22_X1 U22466 ( .A1(n19434), .A2(n19429), .B1(n19432), .B2(
        P2_EAX_REG_11__SCAN_IN), .ZN(n19430) );
  OAI21_X1 U22467 ( .B1(n19437), .B2(n19431), .A(n19430), .ZN(P2_U2908) );
  AOI22_X1 U22468 ( .A1(n19434), .A2(n19433), .B1(n19432), .B2(
        P2_EAX_REG_8__SCAN_IN), .ZN(n19435) );
  OAI21_X1 U22469 ( .B1(n19437), .B2(n19436), .A(n19435), .ZN(P2_U2911) );
  NOR2_X1 U22470 ( .A1(n19445), .A2(n19438), .ZN(P2_U2920) );
  INV_X1 U22471 ( .A(n19439), .ZN(n19442) );
  AOI22_X1 U22472 ( .A1(n19442), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n19475), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19440) );
  OAI21_X1 U22473 ( .B1(n19441), .B2(n19445), .A(n19440), .ZN(P2_U2921) );
  AOI22_X1 U22474 ( .A1(n19442), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n19475), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n19443) );
  OAI21_X1 U22475 ( .B1(n19445), .B2(n19444), .A(n19443), .ZN(P2_U2922) );
  AOI22_X1 U22476 ( .A1(n19475), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19446) );
  OAI21_X1 U22477 ( .B1(n14046), .B2(n19477), .A(n19446), .ZN(P2_U2936) );
  INV_X1 U22478 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19448) );
  AOI22_X1 U22479 ( .A1(n19475), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19447) );
  OAI21_X1 U22480 ( .B1(n19448), .B2(n19477), .A(n19447), .ZN(P2_U2937) );
  AOI22_X1 U22481 ( .A1(n19475), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19449) );
  OAI21_X1 U22482 ( .B1(n19450), .B2(n19477), .A(n19449), .ZN(P2_U2938) );
  AOI22_X1 U22483 ( .A1(n19475), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19451) );
  OAI21_X1 U22484 ( .B1(n19452), .B2(n19477), .A(n19451), .ZN(P2_U2939) );
  AOI22_X1 U22485 ( .A1(n19475), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19453) );
  OAI21_X1 U22486 ( .B1(n19454), .B2(n19477), .A(n19453), .ZN(P2_U2940) );
  AOI22_X1 U22487 ( .A1(n19475), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19455) );
  OAI21_X1 U22488 ( .B1(n19456), .B2(n19477), .A(n19455), .ZN(P2_U2941) );
  INV_X1 U22489 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19458) );
  AOI22_X1 U22490 ( .A1(n19475), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19457) );
  OAI21_X1 U22491 ( .B1(n19458), .B2(n19477), .A(n19457), .ZN(P2_U2942) );
  AOI22_X1 U22492 ( .A1(n19475), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19459) );
  OAI21_X1 U22493 ( .B1(n19460), .B2(n19477), .A(n19459), .ZN(P2_U2943) );
  AOI22_X1 U22494 ( .A1(n19475), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19461) );
  OAI21_X1 U22495 ( .B1(n19462), .B2(n19477), .A(n19461), .ZN(P2_U2944) );
  AOI22_X1 U22496 ( .A1(n19475), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19463) );
  OAI21_X1 U22497 ( .B1(n13444), .B2(n19477), .A(n19463), .ZN(P2_U2945) );
  INV_X1 U22498 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19465) );
  AOI22_X1 U22499 ( .A1(n19475), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19464) );
  OAI21_X1 U22500 ( .B1(n19465), .B2(n19477), .A(n19464), .ZN(P2_U2946) );
  INV_X1 U22501 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19467) );
  AOI22_X1 U22502 ( .A1(n19475), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19466) );
  OAI21_X1 U22503 ( .B1(n19467), .B2(n19477), .A(n19466), .ZN(P2_U2947) );
  INV_X1 U22504 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19469) );
  AOI22_X1 U22505 ( .A1(n19475), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19468) );
  OAI21_X1 U22506 ( .B1(n19469), .B2(n19477), .A(n19468), .ZN(P2_U2948) );
  INV_X1 U22507 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19471) );
  AOI22_X1 U22508 ( .A1(n19475), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19470) );
  OAI21_X1 U22509 ( .B1(n19471), .B2(n19477), .A(n19470), .ZN(P2_U2949) );
  INV_X1 U22510 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19473) );
  AOI22_X1 U22511 ( .A1(n19475), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19472) );
  OAI21_X1 U22512 ( .B1(n19473), .B2(n19477), .A(n19472), .ZN(P2_U2950) );
  AOI22_X1 U22513 ( .A1(n19475), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19474), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19476) );
  OAI21_X1 U22514 ( .B1(n19478), .B2(n19477), .A(n19476), .ZN(P2_U2951) );
  AOI22_X1 U22515 ( .A1(n19487), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n19480) );
  NAND2_X1 U22516 ( .A1(n19482), .A2(n19479), .ZN(n19484) );
  NAND2_X1 U22517 ( .A1(n19480), .A2(n19484), .ZN(P2_U2965) );
  AOI22_X1 U22518 ( .A1(n19487), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n19486), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19483) );
  NAND2_X1 U22519 ( .A1(n19482), .A2(n19481), .ZN(n19488) );
  NAND2_X1 U22520 ( .A1(n19483), .A2(n19488), .ZN(P2_U2966) );
  AOI22_X1 U22521 ( .A1(n19487), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n19486), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n19485) );
  NAND2_X1 U22522 ( .A1(n19485), .A2(n19484), .ZN(P2_U2980) );
  AOI22_X1 U22523 ( .A1(n19487), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n19486), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19489) );
  NAND2_X1 U22524 ( .A1(n19489), .A2(n19488), .ZN(P2_U2981) );
  AOI22_X1 U22525 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19503), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19517), .ZN(n19499) );
  INV_X1 U22526 ( .A(n19490), .ZN(n19491) );
  XNOR2_X1 U22527 ( .A(n19492), .B(n19491), .ZN(n19528) );
  INV_X1 U22528 ( .A(n19528), .ZN(n19496) );
  XNOR2_X1 U22529 ( .A(n9696), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19494) );
  XNOR2_X1 U22530 ( .A(n19494), .B(n19493), .ZN(n19530) );
  OAI22_X1 U22531 ( .A1(n19496), .A2(n19510), .B1(n19495), .B2(n19530), .ZN(
        n19497) );
  AOI21_X1 U22532 ( .B1(n19512), .B2(n19523), .A(n19497), .ZN(n19498) );
  OAI211_X1 U22533 ( .C1(n19501), .C2(n19500), .A(n19499), .B(n19498), .ZN(
        P2_U3010) );
  NOR2_X1 U22534 ( .A1(n19503), .A2(n19502), .ZN(n19516) );
  INV_X1 U22535 ( .A(n19504), .ZN(n19506) );
  AOI21_X1 U22536 ( .B1(n19507), .B2(n19506), .A(n19505), .ZN(n19508) );
  OAI21_X1 U22537 ( .B1(n19510), .B2(n19509), .A(n19508), .ZN(n19511) );
  AOI21_X1 U22538 ( .B1(n19513), .B2(n19512), .A(n19511), .ZN(n19514) );
  OAI21_X1 U22539 ( .B1(n19516), .B2(n19515), .A(n19514), .ZN(P2_U3014) );
  NAND2_X1 U22540 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19517), .ZN(n19518) );
  OAI221_X1 U22541 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19521), .C1(
        n19520), .C2(n19519), .A(n19518), .ZN(n19522) );
  INV_X1 U22542 ( .A(n19522), .ZN(n19526) );
  AOI22_X1 U22543 ( .A1(n19524), .A2(n19537), .B1(n19560), .B2(n19523), .ZN(
        n19525) );
  NAND2_X1 U22544 ( .A1(n19526), .A2(n19525), .ZN(n19527) );
  AOI21_X1 U22545 ( .B1(n19528), .B2(n19551), .A(n19527), .ZN(n19529) );
  OAI21_X1 U22546 ( .B1(n19556), .B2(n19530), .A(n19529), .ZN(P2_U3042) );
  NOR2_X1 U22547 ( .A1(n19532), .A2(n19531), .ZN(n19544) );
  INV_X1 U22548 ( .A(n19533), .ZN(n19543) );
  INV_X1 U22549 ( .A(n19544), .ZN(n19534) );
  AOI22_X1 U22550 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19552), .B1(
        n19535), .B2(n19534), .ZN(n19539) );
  AOI21_X1 U22551 ( .B1(n19537), .B2(n20161), .A(n19536), .ZN(n19538) );
  OAI211_X1 U22552 ( .C1(n19541), .C2(n19540), .A(n19539), .B(n19538), .ZN(
        n19542) );
  AOI21_X1 U22553 ( .B1(n19544), .B2(n19543), .A(n19542), .ZN(n19547) );
  NAND2_X1 U22554 ( .A1(n19551), .A2(n19545), .ZN(n19546) );
  OAI211_X1 U22555 ( .C1(n19548), .C2(n19556), .A(n19547), .B(n19546), .ZN(
        P2_U3044) );
  OAI21_X1 U22556 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n19549), .ZN(n19563) );
  AOI22_X1 U22557 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19552), .B1(
        n19551), .B2(n19550), .ZN(n19562) );
  OAI22_X1 U22558 ( .A1(n19556), .A2(n19555), .B1(n19554), .B2(n19553), .ZN(
        n19557) );
  AOI211_X1 U22559 ( .C1(n19560), .C2(n19559), .A(n19558), .B(n19557), .ZN(
        n19561) );
  OAI211_X1 U22560 ( .C1(n19564), .C2(n19563), .A(n19562), .B(n19561), .ZN(
        P2_U3045) );
  INV_X1 U22561 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19569) );
  AOI22_X1 U22562 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19588), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19587), .ZN(n19929) );
  NOR2_X2 U22563 ( .A1(n19565), .A2(n19583), .ZN(n20016) );
  AOI22_X1 U22564 ( .A1(n20019), .A2(n20053), .B1(n19585), .B2(n20016), .ZN(
        n19568) );
  NOR2_X2 U22565 ( .A1(n19566), .A2(n19915), .ZN(n20017) );
  AOI22_X1 U22566 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19588), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19587), .ZN(n19888) );
  INV_X1 U22567 ( .A(n19888), .ZN(n20018) );
  AOI22_X1 U22568 ( .A1(n20017), .A2(n19589), .B1(n19619), .B2(n20018), .ZN(
        n19567) );
  OAI211_X1 U22569 ( .C1(n19593), .C2(n19569), .A(n19568), .B(n19567), .ZN(
        P2_U3050) );
  AOI22_X1 U22570 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19588), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19587), .ZN(n19932) );
  NOR2_X2 U22571 ( .A1(n9853), .A2(n19583), .ZN(n20023) );
  AOI22_X1 U22572 ( .A1(n20026), .A2(n20053), .B1(n19585), .B2(n20023), .ZN(
        n19572) );
  NOR2_X2 U22573 ( .A1(n19570), .A2(n19915), .ZN(n20024) );
  AOI22_X1 U22574 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19588), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19587), .ZN(n19891) );
  INV_X1 U22575 ( .A(n19891), .ZN(n20025) );
  AOI22_X1 U22576 ( .A1(n20024), .A2(n19589), .B1(n19619), .B2(n20025), .ZN(
        n19571) );
  OAI211_X1 U22577 ( .C1(n19593), .C2(n19573), .A(n19572), .B(n19571), .ZN(
        P2_U3051) );
  INV_X1 U22578 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19577) );
  AOI22_X1 U22579 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19588), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19587), .ZN(n19935) );
  AOI22_X1 U22580 ( .A1(n20032), .A2(n20053), .B1(n19585), .B2(n9671), .ZN(
        n19576) );
  NOR2_X2 U22581 ( .A1(n19574), .A2(n19915), .ZN(n20030) );
  AOI22_X1 U22582 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19588), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19587), .ZN(n19894) );
  INV_X1 U22583 ( .A(n19894), .ZN(n20031) );
  AOI22_X1 U22584 ( .A1(n20030), .A2(n19589), .B1(n19619), .B2(n20031), .ZN(
        n19575) );
  OAI211_X1 U22585 ( .C1(n19593), .C2(n19577), .A(n19576), .B(n19575), .ZN(
        P2_U3052) );
  AOI22_X1 U22586 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19587), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19588), .ZN(n19941) );
  NOR2_X2 U22587 ( .A1(n19578), .A2(n19583), .ZN(n20042) );
  AOI22_X1 U22588 ( .A1(n20045), .A2(n20053), .B1(n19585), .B2(n20042), .ZN(
        n19581) );
  NOR2_X2 U22589 ( .A1(n19579), .A2(n19915), .ZN(n20043) );
  AOI22_X1 U22590 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19588), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19587), .ZN(n19901) );
  INV_X1 U22591 ( .A(n19901), .ZN(n20044) );
  AOI22_X1 U22592 ( .A1(n20043), .A2(n19589), .B1(n19619), .B2(n20044), .ZN(
        n19580) );
  OAI211_X1 U22593 ( .C1(n19593), .C2(n19582), .A(n19581), .B(n19580), .ZN(
        P2_U3054) );
  AOI22_X1 U22594 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19588), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19587), .ZN(n19948) );
  NOR2_X2 U22595 ( .A1(n19584), .A2(n19583), .ZN(n20048) );
  AOI22_X1 U22596 ( .A1(n20054), .A2(n20053), .B1(n19585), .B2(n20048), .ZN(
        n19591) );
  NOR2_X2 U22597 ( .A1(n19586), .A2(n19915), .ZN(n20050) );
  AOI22_X1 U22598 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19588), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19587), .ZN(n19882) );
  INV_X1 U22599 ( .A(n19882), .ZN(n20052) );
  AOI22_X1 U22600 ( .A1(n20050), .A2(n19589), .B1(n19619), .B2(n20052), .ZN(
        n19590) );
  OAI211_X1 U22601 ( .C1(n19593), .C2(n19592), .A(n19591), .B(n19590), .ZN(
        P2_U3055) );
  INV_X1 U22602 ( .A(n20067), .ZN(n19758) );
  NOR2_X1 U22603 ( .A1(n19819), .A2(n19644), .ZN(n19617) );
  NOR3_X1 U22604 ( .A1(n19594), .A2(n19617), .A3(n20065), .ZN(n19598) );
  AOI211_X2 U22605 ( .C1(n19599), .C2(n20065), .A(n19758), .B(n19598), .ZN(
        n19618) );
  AOI22_X1 U22606 ( .A1(n19618), .A2(n20003), .B1(n20002), .B2(n19617), .ZN(
        n19603) );
  OR2_X1 U22607 ( .A1(n20154), .A2(n19595), .ZN(n19761) );
  INV_X1 U22608 ( .A(n19761), .ZN(n19597) );
  NAND2_X1 U22609 ( .A1(n19597), .A2(n19596), .ZN(n19600) );
  AOI21_X1 U22610 ( .B1(n19600), .B2(n19599), .A(n19598), .ZN(n19601) );
  OAI211_X1 U22611 ( .C1(n19617), .C2(n19920), .A(n19601), .B(n19995), .ZN(
        n19620) );
  AOI22_X1 U22612 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19620), .B1(
        n19619), .B2(n20004), .ZN(n19602) );
  OAI211_X1 U22613 ( .C1(n19831), .C2(n19623), .A(n19603), .B(n19602), .ZN(
        P2_U3056) );
  AOI22_X1 U22614 ( .A1(n19618), .A2(n20010), .B1(n20009), .B2(n19617), .ZN(
        n19605) );
  AOI22_X1 U22615 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19620), .B1(
        n19619), .B2(n20012), .ZN(n19604) );
  OAI211_X1 U22616 ( .C1(n19864), .C2(n19623), .A(n19605), .B(n19604), .ZN(
        P2_U3057) );
  AOI22_X1 U22617 ( .A1(n19618), .A2(n20017), .B1(n20016), .B2(n19617), .ZN(
        n19607) );
  AOI22_X1 U22618 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19620), .B1(
        n19619), .B2(n20019), .ZN(n19606) );
  OAI211_X1 U22619 ( .C1(n19888), .C2(n19623), .A(n19607), .B(n19606), .ZN(
        P2_U3058) );
  AOI22_X1 U22620 ( .A1(n19618), .A2(n20024), .B1(n20023), .B2(n19617), .ZN(
        n19609) );
  AOI22_X1 U22621 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19620), .B1(
        n19619), .B2(n20026), .ZN(n19608) );
  OAI211_X1 U22622 ( .C1(n19891), .C2(n19623), .A(n19609), .B(n19608), .ZN(
        P2_U3059) );
  AOI22_X1 U22623 ( .A1(n19618), .A2(n20030), .B1(n9671), .B2(n19617), .ZN(
        n19611) );
  AOI22_X1 U22624 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19620), .B1(
        n19619), .B2(n20032), .ZN(n19610) );
  OAI211_X1 U22625 ( .C1(n19894), .C2(n19623), .A(n19611), .B(n19610), .ZN(
        P2_U3060) );
  AOI22_X1 U22626 ( .A1(n19618), .A2(n20037), .B1(n20036), .B2(n19617), .ZN(
        n19614) );
  AOI22_X1 U22627 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19620), .B1(
        n19619), .B2(n20039), .ZN(n19613) );
  OAI211_X1 U22628 ( .C1(n19897), .C2(n19623), .A(n19614), .B(n19613), .ZN(
        P2_U3061) );
  AOI22_X1 U22629 ( .A1(n19618), .A2(n20043), .B1(n20042), .B2(n19617), .ZN(
        n19616) );
  AOI22_X1 U22630 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19620), .B1(
        n19619), .B2(n20045), .ZN(n19615) );
  OAI211_X1 U22631 ( .C1(n19901), .C2(n19623), .A(n19616), .B(n19615), .ZN(
        P2_U3062) );
  AOI22_X1 U22632 ( .A1(n19618), .A2(n20050), .B1(n20048), .B2(n19617), .ZN(
        n19622) );
  AOI22_X1 U22633 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19620), .B1(
        n19619), .B2(n20054), .ZN(n19621) );
  OAI211_X1 U22634 ( .C1(n19882), .C2(n19623), .A(n19622), .B(n19621), .ZN(
        P2_U3063) );
  AOI22_X1 U22635 ( .A1(n19638), .A2(n20010), .B1(n20009), .B2(n19637), .ZN(
        n19626) );
  INV_X1 U22636 ( .A(n19624), .ZN(n19640) );
  AOI22_X1 U22637 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n20012), .ZN(n19625) );
  OAI211_X1 U22638 ( .C1(n19864), .C2(n19664), .A(n19626), .B(n19625), .ZN(
        P2_U3065) );
  AOI22_X1 U22639 ( .A1(n19638), .A2(n20017), .B1(n20016), .B2(n19637), .ZN(
        n19628) );
  AOI22_X1 U22640 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n20019), .ZN(n19627) );
  OAI211_X1 U22641 ( .C1(n19888), .C2(n19664), .A(n19628), .B(n19627), .ZN(
        P2_U3066) );
  AOI22_X1 U22642 ( .A1(n19638), .A2(n20024), .B1(n20023), .B2(n19637), .ZN(
        n19630) );
  AOI22_X1 U22643 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n20026), .ZN(n19629) );
  OAI211_X1 U22644 ( .C1(n19891), .C2(n19664), .A(n19630), .B(n19629), .ZN(
        P2_U3067) );
  AOI22_X1 U22645 ( .A1(n19638), .A2(n20030), .B1(n9671), .B2(n19637), .ZN(
        n19632) );
  AOI22_X1 U22646 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n20032), .ZN(n19631) );
  OAI211_X1 U22647 ( .C1(n19894), .C2(n19664), .A(n19632), .B(n19631), .ZN(
        P2_U3068) );
  AOI22_X1 U22648 ( .A1(n19638), .A2(n20037), .B1(n20036), .B2(n19637), .ZN(
        n19634) );
  AOI22_X1 U22649 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n20039), .ZN(n19633) );
  OAI211_X1 U22650 ( .C1(n19897), .C2(n19664), .A(n19634), .B(n19633), .ZN(
        P2_U3069) );
  AOI22_X1 U22651 ( .A1(n19638), .A2(n20043), .B1(n20042), .B2(n19637), .ZN(
        n19636) );
  AOI22_X1 U22652 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n20045), .ZN(n19635) );
  OAI211_X1 U22653 ( .C1(n19901), .C2(n19664), .A(n19636), .B(n19635), .ZN(
        P2_U3070) );
  AOI22_X1 U22654 ( .A1(n19638), .A2(n20050), .B1(n20048), .B2(n19637), .ZN(
        n19642) );
  AOI22_X1 U22655 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19640), .B1(
        n19639), .B2(n20054), .ZN(n19641) );
  OAI211_X1 U22656 ( .C1(n19882), .C2(n19664), .A(n19642), .B(n19641), .ZN(
        P2_U3071) );
  NOR2_X1 U22657 ( .A1(n19755), .A2(n19644), .ZN(n19667) );
  AOI22_X1 U22658 ( .A1(n20004), .A2(n19668), .B1(n20002), .B2(n19667), .ZN(
        n19653) );
  OAI21_X1 U22659 ( .B1(n19761), .B2(n19643), .A(n20157), .ZN(n19651) );
  NOR2_X1 U22660 ( .A1(n10356), .A2(n19644), .ZN(n19647) );
  INV_X1 U22661 ( .A(n19667), .ZN(n19645) );
  OAI211_X1 U22662 ( .C1(n12021), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20150), 
        .B(n19645), .ZN(n19646) );
  OAI211_X1 U22663 ( .C1(n19651), .C2(n19647), .A(n19995), .B(n19646), .ZN(
        n19670) );
  INV_X1 U22664 ( .A(n19647), .ZN(n19650) );
  OAI21_X1 U22665 ( .B1(n19648), .B2(n19667), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19649) );
  OAI21_X1 U22666 ( .B1(n19651), .B2(n19650), .A(n19649), .ZN(n19669) );
  AOI22_X1 U22667 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19670), .B1(
        n20003), .B2(n19669), .ZN(n19652) );
  OAI211_X1 U22668 ( .C1(n19831), .C2(n19686), .A(n19653), .B(n19652), .ZN(
        P2_U3072) );
  AOI22_X1 U22669 ( .A1(n19668), .A2(n20012), .B1(n20009), .B2(n19667), .ZN(
        n19655) );
  AOI22_X1 U22670 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19670), .B1(
        n20010), .B2(n19669), .ZN(n19654) );
  OAI211_X1 U22671 ( .C1(n19864), .C2(n19686), .A(n19655), .B(n19654), .ZN(
        P2_U3073) );
  AOI22_X1 U22672 ( .A1(n19668), .A2(n20019), .B1(n19667), .B2(n20016), .ZN(
        n19657) );
  AOI22_X1 U22673 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19670), .B1(
        n20017), .B2(n19669), .ZN(n19656) );
  OAI211_X1 U22674 ( .C1(n19888), .C2(n19686), .A(n19657), .B(n19656), .ZN(
        P2_U3074) );
  AOI22_X1 U22675 ( .A1(n20025), .A2(n19691), .B1(n19667), .B2(n20023), .ZN(
        n19659) );
  AOI22_X1 U22676 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19670), .B1(
        n20024), .B2(n19669), .ZN(n19658) );
  OAI211_X1 U22677 ( .C1(n19932), .C2(n19664), .A(n19659), .B(n19658), .ZN(
        P2_U3075) );
  AOI22_X1 U22678 ( .A1(n20031), .A2(n19691), .B1(n19667), .B2(n9671), .ZN(
        n19661) );
  AOI22_X1 U22679 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19670), .B1(
        n20030), .B2(n19669), .ZN(n19660) );
  OAI211_X1 U22680 ( .C1(n19935), .C2(n19664), .A(n19661), .B(n19660), .ZN(
        P2_U3076) );
  INV_X1 U22681 ( .A(n19897), .ZN(n20038) );
  AOI22_X1 U22682 ( .A1(n20038), .A2(n19691), .B1(n20036), .B2(n19667), .ZN(
        n19663) );
  AOI22_X1 U22683 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19670), .B1(
        n20037), .B2(n19669), .ZN(n19662) );
  OAI211_X1 U22684 ( .C1(n19938), .C2(n19664), .A(n19663), .B(n19662), .ZN(
        P2_U3077) );
  AOI22_X1 U22685 ( .A1(n19668), .A2(n20045), .B1(n19667), .B2(n20042), .ZN(
        n19666) );
  AOI22_X1 U22686 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19670), .B1(
        n20043), .B2(n19669), .ZN(n19665) );
  OAI211_X1 U22687 ( .C1(n19901), .C2(n19686), .A(n19666), .B(n19665), .ZN(
        P2_U3078) );
  AOI22_X1 U22688 ( .A1(n19668), .A2(n20054), .B1(n19667), .B2(n20048), .ZN(
        n19672) );
  AOI22_X1 U22689 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19670), .B1(
        n20050), .B2(n19669), .ZN(n19671) );
  OAI211_X1 U22690 ( .C1(n19882), .C2(n19686), .A(n19672), .B(n19671), .ZN(
        P2_U3079) );
  INV_X1 U22691 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n19675) );
  AOI22_X1 U22692 ( .A1(n19690), .A2(n20003), .B1(n20002), .B2(n19689), .ZN(
        n19674) );
  AOI22_X1 U22693 ( .A1(n19713), .A2(n20005), .B1(n19691), .B2(n20004), .ZN(
        n19673) );
  OAI211_X1 U22694 ( .C1(n19679), .C2(n19675), .A(n19674), .B(n19673), .ZN(
        P2_U3080) );
  INV_X1 U22695 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n19678) );
  AOI22_X1 U22696 ( .A1(n19690), .A2(n20017), .B1(n20016), .B2(n19689), .ZN(
        n19677) );
  AOI22_X1 U22697 ( .A1(n19691), .A2(n20019), .B1(n19713), .B2(n20018), .ZN(
        n19676) );
  OAI211_X1 U22698 ( .C1(n19679), .C2(n19678), .A(n19677), .B(n19676), .ZN(
        P2_U3082) );
  AOI22_X1 U22699 ( .A1(n19690), .A2(n20024), .B1(n20023), .B2(n19689), .ZN(
        n19681) );
  AOI22_X1 U22700 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19692), .B1(
        n19713), .B2(n20025), .ZN(n19680) );
  OAI211_X1 U22701 ( .C1(n19932), .C2(n19686), .A(n19681), .B(n19680), .ZN(
        P2_U3083) );
  AOI22_X1 U22702 ( .A1(n19690), .A2(n20030), .B1(n9671), .B2(n19689), .ZN(
        n19683) );
  AOI22_X1 U22703 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19692), .B1(
        n19713), .B2(n20031), .ZN(n19682) );
  OAI211_X1 U22704 ( .C1(n19935), .C2(n19686), .A(n19683), .B(n19682), .ZN(
        P2_U3084) );
  AOI22_X1 U22705 ( .A1(n19690), .A2(n20037), .B1(n20036), .B2(n19689), .ZN(
        n19685) );
  AOI22_X1 U22706 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19692), .B1(
        n19713), .B2(n20038), .ZN(n19684) );
  OAI211_X1 U22707 ( .C1(n19938), .C2(n19686), .A(n19685), .B(n19684), .ZN(
        P2_U3085) );
  AOI22_X1 U22708 ( .A1(n19690), .A2(n20043), .B1(n20042), .B2(n19689), .ZN(
        n19688) );
  AOI22_X1 U22709 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19692), .B1(
        n19691), .B2(n20045), .ZN(n19687) );
  OAI211_X1 U22710 ( .C1(n19901), .C2(n19724), .A(n19688), .B(n19687), .ZN(
        P2_U3086) );
  AOI22_X1 U22711 ( .A1(n19690), .A2(n20050), .B1(n20048), .B2(n19689), .ZN(
        n19694) );
  AOI22_X1 U22712 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19692), .B1(
        n19691), .B2(n20054), .ZN(n19693) );
  OAI211_X1 U22713 ( .C1(n19882), .C2(n19724), .A(n19694), .B(n19693), .ZN(
        P2_U3087) );
  NOR2_X2 U22714 ( .A1(n19695), .A2(n19696), .ZN(n19749) );
  NOR2_X1 U22715 ( .A1(n19819), .A2(n19754), .ZN(n19728) );
  AOI22_X1 U22716 ( .A1(n20005), .A2(n19749), .B1(n20002), .B2(n19728), .ZN(
        n19706) );
  OAI21_X1 U22717 ( .B1(n19761), .B2(n19696), .A(n20157), .ZN(n19704) );
  NOR2_X1 U22718 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19754), .ZN(
        n19700) );
  OAI21_X1 U22719 ( .B1(n19701), .B2(n20065), .A(n19920), .ZN(n19698) );
  INV_X1 U22720 ( .A(n19728), .ZN(n19697) );
  AOI21_X1 U22721 ( .B1(n19698), .B2(n19697), .A(n19915), .ZN(n19699) );
  OAI21_X1 U22722 ( .B1(n19704), .B2(n19700), .A(n19699), .ZN(n19721) );
  INV_X1 U22723 ( .A(n19700), .ZN(n19703) );
  OAI21_X1 U22724 ( .B1(n19701), .B2(n19728), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19702) );
  OAI21_X1 U22725 ( .B1(n19704), .B2(n19703), .A(n19702), .ZN(n19720) );
  AOI22_X1 U22726 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19721), .B1(
        n20003), .B2(n19720), .ZN(n19705) );
  OAI211_X1 U22727 ( .C1(n19923), .C2(n19724), .A(n19706), .B(n19705), .ZN(
        P2_U3088) );
  AOI22_X1 U22728 ( .A1(n20011), .A2(n19749), .B1(n20009), .B2(n19728), .ZN(
        n19708) );
  AOI22_X1 U22729 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19721), .B1(
        n20010), .B2(n19720), .ZN(n19707) );
  OAI211_X1 U22730 ( .C1(n19926), .C2(n19724), .A(n19708), .B(n19707), .ZN(
        P2_U3089) );
  AOI22_X1 U22731 ( .A1(n20018), .A2(n19749), .B1(n19728), .B2(n20016), .ZN(
        n19710) );
  AOI22_X1 U22732 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19721), .B1(
        n20017), .B2(n19720), .ZN(n19709) );
  OAI211_X1 U22733 ( .C1(n19929), .C2(n19724), .A(n19710), .B(n19709), .ZN(
        P2_U3090) );
  AOI22_X1 U22734 ( .A1(n20025), .A2(n19749), .B1(n19728), .B2(n20023), .ZN(
        n19712) );
  AOI22_X1 U22735 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19721), .B1(
        n20024), .B2(n19720), .ZN(n19711) );
  OAI211_X1 U22736 ( .C1(n19932), .C2(n19724), .A(n19712), .B(n19711), .ZN(
        P2_U3091) );
  INV_X1 U22737 ( .A(n19749), .ZN(n19734) );
  AOI22_X1 U22738 ( .A1(n20032), .A2(n19713), .B1(n9671), .B2(n19728), .ZN(
        n19715) );
  AOI22_X1 U22739 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19721), .B1(
        n20030), .B2(n19720), .ZN(n19714) );
  OAI211_X1 U22740 ( .C1(n19894), .C2(n19734), .A(n19715), .B(n19714), .ZN(
        P2_U3092) );
  AOI22_X1 U22741 ( .A1(n20038), .A2(n19749), .B1(n20036), .B2(n19728), .ZN(
        n19717) );
  AOI22_X1 U22742 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19721), .B1(
        n20037), .B2(n19720), .ZN(n19716) );
  OAI211_X1 U22743 ( .C1(n19938), .C2(n19724), .A(n19717), .B(n19716), .ZN(
        P2_U3093) );
  AOI22_X1 U22744 ( .A1(n20044), .A2(n19749), .B1(n19728), .B2(n20042), .ZN(
        n19719) );
  AOI22_X1 U22745 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19721), .B1(
        n20043), .B2(n19720), .ZN(n19718) );
  OAI211_X1 U22746 ( .C1(n19941), .C2(n19724), .A(n19719), .B(n19718), .ZN(
        P2_U3094) );
  AOI22_X1 U22747 ( .A1(n20052), .A2(n19749), .B1(n19728), .B2(n20048), .ZN(
        n19723) );
  AOI22_X1 U22748 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19721), .B1(
        n20050), .B2(n19720), .ZN(n19722) );
  OAI211_X1 U22749 ( .C1(n19948), .C2(n19724), .A(n19723), .B(n19722), .ZN(
        P2_U3095) );
  NOR2_X1 U22750 ( .A1(n19850), .A2(n19754), .ZN(n19747) );
  OAI21_X1 U22751 ( .B1(n19725), .B2(n19747), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19726) );
  OAI21_X1 U22752 ( .B1(n19754), .B2(n19853), .A(n19726), .ZN(n19748) );
  AOI22_X1 U22753 ( .A1(n19748), .A2(n20003), .B1(n20002), .B2(n19747), .ZN(
        n19733) );
  AOI221_X1 U22754 ( .B1(n19749), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19782), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19728), .ZN(n19729) );
  AOI211_X1 U22755 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19730), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19729), .ZN(n19731) );
  AOI22_X1 U22756 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19750), .B1(
        n19782), .B2(n20005), .ZN(n19732) );
  OAI211_X1 U22757 ( .C1(n19923), .C2(n19734), .A(n19733), .B(n19732), .ZN(
        P2_U3096) );
  AOI22_X1 U22758 ( .A1(n19748), .A2(n20010), .B1(n20009), .B2(n19747), .ZN(
        n19736) );
  AOI22_X1 U22759 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19750), .B1(
        n19749), .B2(n20012), .ZN(n19735) );
  OAI211_X1 U22760 ( .C1(n19864), .C2(n19780), .A(n19736), .B(n19735), .ZN(
        P2_U3097) );
  AOI22_X1 U22761 ( .A1(n19748), .A2(n20017), .B1(n20016), .B2(n19747), .ZN(
        n19738) );
  AOI22_X1 U22762 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19750), .B1(
        n19749), .B2(n20019), .ZN(n19737) );
  OAI211_X1 U22763 ( .C1(n19888), .C2(n19780), .A(n19738), .B(n19737), .ZN(
        P2_U3098) );
  AOI22_X1 U22764 ( .A1(n19748), .A2(n20024), .B1(n20023), .B2(n19747), .ZN(
        n19740) );
  AOI22_X1 U22765 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19750), .B1(
        n19749), .B2(n20026), .ZN(n19739) );
  OAI211_X1 U22766 ( .C1(n19891), .C2(n19780), .A(n19740), .B(n19739), .ZN(
        P2_U3099) );
  AOI22_X1 U22767 ( .A1(n19748), .A2(n20030), .B1(n9671), .B2(n19747), .ZN(
        n19742) );
  AOI22_X1 U22768 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19750), .B1(
        n19749), .B2(n20032), .ZN(n19741) );
  OAI211_X1 U22769 ( .C1(n19894), .C2(n19780), .A(n19742), .B(n19741), .ZN(
        P2_U3100) );
  AOI22_X1 U22770 ( .A1(n19748), .A2(n20037), .B1(n20036), .B2(n19747), .ZN(
        n19744) );
  AOI22_X1 U22771 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19750), .B1(
        n19749), .B2(n20039), .ZN(n19743) );
  OAI211_X1 U22772 ( .C1(n19897), .C2(n19780), .A(n19744), .B(n19743), .ZN(
        P2_U3101) );
  AOI22_X1 U22773 ( .A1(n19748), .A2(n20043), .B1(n20042), .B2(n19747), .ZN(
        n19746) );
  AOI22_X1 U22774 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19750), .B1(
        n19749), .B2(n20045), .ZN(n19745) );
  OAI211_X1 U22775 ( .C1(n19901), .C2(n19780), .A(n19746), .B(n19745), .ZN(
        P2_U3102) );
  AOI22_X1 U22776 ( .A1(n19748), .A2(n20050), .B1(n20048), .B2(n19747), .ZN(
        n19752) );
  AOI22_X1 U22777 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19750), .B1(
        n19749), .B2(n20054), .ZN(n19751) );
  OAI211_X1 U22778 ( .C1(n19882), .C2(n19780), .A(n19752), .B(n19751), .ZN(
        P2_U3103) );
  NOR2_X1 U22779 ( .A1(n19991), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19765) );
  INV_X1 U22780 ( .A(n19765), .ZN(n19759) );
  NOR2_X1 U22781 ( .A1(n19755), .A2(n19754), .ZN(n19791) );
  NOR2_X1 U22782 ( .A1(n19791), .A2(n20065), .ZN(n19756) );
  AND2_X1 U22783 ( .A1(n19757), .A2(n19756), .ZN(n19763) );
  AOI211_X2 U22784 ( .C1(n19759), .C2(n20065), .A(n19758), .B(n19763), .ZN(
        n19781) );
  AOI22_X1 U22785 ( .A1(n19781), .A2(n20003), .B1(n20002), .B2(n19791), .ZN(
        n19767) );
  NOR2_X1 U22786 ( .A1(n19761), .A2(n19760), .ZN(n20152) );
  OAI21_X1 U22787 ( .B1(n19791), .B2(n19920), .A(n19995), .ZN(n19762) );
  NOR2_X1 U22788 ( .A1(n19763), .A2(n19762), .ZN(n19764) );
  OAI21_X1 U22789 ( .B1(n20152), .B2(n19765), .A(n19764), .ZN(n19783) );
  AOI22_X1 U22790 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19783), .B1(
        n19782), .B2(n20004), .ZN(n19766) );
  OAI211_X1 U22791 ( .C1(n19831), .C2(n19799), .A(n19767), .B(n19766), .ZN(
        P2_U3104) );
  AOI22_X1 U22792 ( .A1(n19781), .A2(n20010), .B1(n20009), .B2(n19791), .ZN(
        n19769) );
  AOI22_X1 U22793 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19783), .B1(
        n19782), .B2(n20012), .ZN(n19768) );
  OAI211_X1 U22794 ( .C1(n19864), .C2(n19799), .A(n19769), .B(n19768), .ZN(
        P2_U3105) );
  AOI22_X1 U22795 ( .A1(n19781), .A2(n20017), .B1(n19791), .B2(n20016), .ZN(
        n19771) );
  AOI22_X1 U22796 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19783), .B1(
        n19813), .B2(n20018), .ZN(n19770) );
  OAI211_X1 U22797 ( .C1(n19929), .C2(n19780), .A(n19771), .B(n19770), .ZN(
        P2_U3106) );
  AOI22_X1 U22798 ( .A1(n19781), .A2(n20024), .B1(n19791), .B2(n20023), .ZN(
        n19773) );
  AOI22_X1 U22799 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19783), .B1(
        n19782), .B2(n20026), .ZN(n19772) );
  OAI211_X1 U22800 ( .C1(n19891), .C2(n19799), .A(n19773), .B(n19772), .ZN(
        P2_U3107) );
  AOI22_X1 U22801 ( .A1(n19781), .A2(n20030), .B1(n19791), .B2(n9671), .ZN(
        n19775) );
  AOI22_X1 U22802 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19783), .B1(
        n19813), .B2(n20031), .ZN(n19774) );
  OAI211_X1 U22803 ( .C1(n19935), .C2(n19780), .A(n19775), .B(n19774), .ZN(
        P2_U3108) );
  AOI22_X1 U22804 ( .A1(n19781), .A2(n20037), .B1(n20036), .B2(n19791), .ZN(
        n19777) );
  AOI22_X1 U22805 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19783), .B1(
        n19782), .B2(n20039), .ZN(n19776) );
  OAI211_X1 U22806 ( .C1(n19897), .C2(n19799), .A(n19777), .B(n19776), .ZN(
        P2_U3109) );
  AOI22_X1 U22807 ( .A1(n19781), .A2(n20043), .B1(n19791), .B2(n20042), .ZN(
        n19779) );
  AOI22_X1 U22808 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19783), .B1(
        n19813), .B2(n20044), .ZN(n19778) );
  OAI211_X1 U22809 ( .C1(n19941), .C2(n19780), .A(n19779), .B(n19778), .ZN(
        P2_U3110) );
  AOI22_X1 U22810 ( .A1(n19781), .A2(n20050), .B1(n19791), .B2(n20048), .ZN(
        n19785) );
  AOI22_X1 U22811 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19783), .B1(
        n19782), .B2(n20054), .ZN(n19784) );
  OAI211_X1 U22812 ( .C1(n19882), .C2(n19799), .A(n19785), .B(n19784), .ZN(
        P2_U3111) );
  NAND2_X1 U22813 ( .A1(n19787), .A2(n10356), .ZN(n19827) );
  NOR2_X1 U22814 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19827), .ZN(
        n19812) );
  AOI22_X1 U22815 ( .A1(n20005), .A2(n19845), .B1(n20002), .B2(n19812), .ZN(
        n19798) );
  OAI21_X1 U22816 ( .B1(n19813), .B2(n19845), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19788) );
  NAND2_X1 U22817 ( .A1(n19788), .A2(n20157), .ZN(n19796) );
  NOR2_X1 U22818 ( .A1(n19791), .A2(n19796), .ZN(n19789) );
  NOR2_X1 U22819 ( .A1(n19791), .A2(n19812), .ZN(n19795) );
  INV_X1 U22820 ( .A(n19792), .ZN(n19793) );
  OAI21_X1 U22821 ( .B1(n19793), .B2(n19812), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19794) );
  AOI22_X1 U22822 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19815), .B1(
        n20003), .B2(n19814), .ZN(n19797) );
  OAI211_X1 U22823 ( .C1(n19923), .C2(n19799), .A(n19798), .B(n19797), .ZN(
        P2_U3112) );
  AOI22_X1 U22824 ( .A1(n19813), .A2(n20012), .B1(n20009), .B2(n19812), .ZN(
        n19801) );
  AOI22_X1 U22825 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n20010), .ZN(n19800) );
  OAI211_X1 U22826 ( .C1(n19864), .C2(n19844), .A(n19801), .B(n19800), .ZN(
        P2_U3113) );
  AOI22_X1 U22827 ( .A1(n19813), .A2(n20019), .B1(n20016), .B2(n19812), .ZN(
        n19803) );
  AOI22_X1 U22828 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n20017), .ZN(n19802) );
  OAI211_X1 U22829 ( .C1(n19888), .C2(n19844), .A(n19803), .B(n19802), .ZN(
        P2_U3114) );
  AOI22_X1 U22830 ( .A1(n20026), .A2(n19813), .B1(n19812), .B2(n20023), .ZN(
        n19805) );
  AOI22_X1 U22831 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n20024), .ZN(n19804) );
  OAI211_X1 U22832 ( .C1(n19891), .C2(n19844), .A(n19805), .B(n19804), .ZN(
        P2_U3115) );
  AOI22_X1 U22833 ( .A1(n20032), .A2(n19813), .B1(n9671), .B2(n19812), .ZN(
        n19807) );
  AOI22_X1 U22834 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n20030), .ZN(n19806) );
  OAI211_X1 U22835 ( .C1(n19894), .C2(n19844), .A(n19807), .B(n19806), .ZN(
        P2_U3116) );
  AOI22_X1 U22836 ( .A1(n20039), .A2(n19813), .B1(n20036), .B2(n19812), .ZN(
        n19809) );
  AOI22_X1 U22837 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n20037), .ZN(n19808) );
  OAI211_X1 U22838 ( .C1(n19897), .C2(n19844), .A(n19809), .B(n19808), .ZN(
        P2_U3117) );
  AOI22_X1 U22839 ( .A1(n19813), .A2(n20045), .B1(n20042), .B2(n19812), .ZN(
        n19811) );
  AOI22_X1 U22840 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n20043), .ZN(n19810) );
  OAI211_X1 U22841 ( .C1(n19901), .C2(n19844), .A(n19811), .B(n19810), .ZN(
        P2_U3118) );
  AOI22_X1 U22842 ( .A1(n19813), .A2(n20054), .B1(n20048), .B2(n19812), .ZN(
        n19817) );
  AOI22_X1 U22843 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19815), .B1(
        n19814), .B2(n20050), .ZN(n19816) );
  OAI211_X1 U22844 ( .C1(n19882), .C2(n19844), .A(n19817), .B(n19816), .ZN(
        P2_U3119) );
  NOR2_X2 U22845 ( .A1(n19820), .A2(n19818), .ZN(n19877) );
  INV_X1 U22846 ( .A(n19877), .ZN(n19861) );
  NOR2_X1 U22847 ( .A1(n19819), .A2(n19854), .ZN(n19855) );
  AOI22_X1 U22848 ( .A1(n20004), .A2(n19845), .B1(n20002), .B2(n19855), .ZN(
        n19830) );
  INV_X1 U22849 ( .A(n19992), .ZN(n19821) );
  OAI21_X1 U22850 ( .B1(n19821), .B2(n19820), .A(n20157), .ZN(n19828) );
  INV_X1 U22851 ( .A(n19828), .ZN(n19824) );
  INV_X1 U22852 ( .A(n19822), .ZN(n19823) );
  NOR2_X1 U22853 ( .A1(n19823), .A2(n19855), .ZN(n19826) );
  AOI22_X1 U22854 ( .A1(n19824), .A2(n19827), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19826), .ZN(n19825) );
  OAI211_X1 U22855 ( .C1(n19855), .C2(n19920), .A(n19825), .B(n19995), .ZN(
        n19847) );
  OAI22_X1 U22856 ( .A1(n19828), .A2(n19827), .B1(n19826), .B2(n20065), .ZN(
        n19846) );
  AOI22_X1 U22857 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19847), .B1(
        n20003), .B2(n19846), .ZN(n19829) );
  OAI211_X1 U22858 ( .C1(n19831), .C2(n19861), .A(n19830), .B(n19829), .ZN(
        P2_U3120) );
  AOI22_X1 U22859 ( .A1(n20011), .A2(n19877), .B1(n20009), .B2(n19855), .ZN(
        n19833) );
  AOI22_X1 U22860 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19847), .B1(
        n20010), .B2(n19846), .ZN(n19832) );
  OAI211_X1 U22861 ( .C1(n19926), .C2(n19844), .A(n19833), .B(n19832), .ZN(
        P2_U3121) );
  AOI22_X1 U22862 ( .A1(n20018), .A2(n19877), .B1(n20016), .B2(n19855), .ZN(
        n19835) );
  AOI22_X1 U22863 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19847), .B1(
        n20017), .B2(n19846), .ZN(n19834) );
  OAI211_X1 U22864 ( .C1(n19929), .C2(n19844), .A(n19835), .B(n19834), .ZN(
        P2_U3122) );
  AOI22_X1 U22865 ( .A1(n20025), .A2(n19877), .B1(n20023), .B2(n19855), .ZN(
        n19837) );
  AOI22_X1 U22866 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19847), .B1(
        n20024), .B2(n19846), .ZN(n19836) );
  OAI211_X1 U22867 ( .C1(n19932), .C2(n19844), .A(n19837), .B(n19836), .ZN(
        P2_U3123) );
  AOI22_X1 U22868 ( .A1(n20031), .A2(n19877), .B1(n9671), .B2(n19855), .ZN(
        n19839) );
  AOI22_X1 U22869 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19847), .B1(
        n20030), .B2(n19846), .ZN(n19838) );
  OAI211_X1 U22870 ( .C1(n19935), .C2(n19844), .A(n19839), .B(n19838), .ZN(
        P2_U3124) );
  AOI22_X1 U22871 ( .A1(n20038), .A2(n19877), .B1(n20036), .B2(n19855), .ZN(
        n19841) );
  AOI22_X1 U22872 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19847), .B1(
        n20037), .B2(n19846), .ZN(n19840) );
  OAI211_X1 U22873 ( .C1(n19938), .C2(n19844), .A(n19841), .B(n19840), .ZN(
        P2_U3125) );
  AOI22_X1 U22874 ( .A1(n20044), .A2(n19877), .B1(n20042), .B2(n19855), .ZN(
        n19843) );
  AOI22_X1 U22875 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19847), .B1(
        n20043), .B2(n19846), .ZN(n19842) );
  OAI211_X1 U22876 ( .C1(n19941), .C2(n19844), .A(n19843), .B(n19842), .ZN(
        P2_U3126) );
  AOI22_X1 U22877 ( .A1(n19845), .A2(n20054), .B1(n20048), .B2(n19855), .ZN(
        n19849) );
  AOI22_X1 U22878 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19847), .B1(
        n20050), .B2(n19846), .ZN(n19848) );
  OAI211_X1 U22879 ( .C1(n19882), .C2(n19861), .A(n19849), .B(n19848), .ZN(
        P2_U3127) );
  NOR2_X1 U22880 ( .A1(n19850), .A2(n19854), .ZN(n19875) );
  OAI21_X1 U22881 ( .B1(n19851), .B2(n19875), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19852) );
  OAI21_X1 U22882 ( .B1(n19854), .B2(n19853), .A(n19852), .ZN(n19876) );
  AOI22_X1 U22883 ( .A1(n19876), .A2(n20003), .B1(n20002), .B2(n19875), .ZN(
        n19860) );
  AOI221_X1 U22884 ( .B1(n19877), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19904), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19855), .ZN(n19856) );
  AOI211_X1 U22885 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19857), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19856), .ZN(n19858) );
  AOI22_X1 U22886 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19878), .B1(
        n19904), .B2(n20005), .ZN(n19859) );
  OAI211_X1 U22887 ( .C1(n19923), .C2(n19861), .A(n19860), .B(n19859), .ZN(
        P2_U3128) );
  AOI22_X1 U22888 ( .A1(n19876), .A2(n20010), .B1(n20009), .B2(n19875), .ZN(
        n19863) );
  AOI22_X1 U22889 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19878), .B1(
        n19877), .B2(n20012), .ZN(n19862) );
  OAI211_X1 U22890 ( .C1(n19864), .C2(n19881), .A(n19863), .B(n19862), .ZN(
        P2_U3129) );
  AOI22_X1 U22891 ( .A1(n19876), .A2(n20017), .B1(n20016), .B2(n19875), .ZN(
        n19866) );
  AOI22_X1 U22892 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19878), .B1(
        n19877), .B2(n20019), .ZN(n19865) );
  OAI211_X1 U22893 ( .C1(n19888), .C2(n19881), .A(n19866), .B(n19865), .ZN(
        P2_U3130) );
  AOI22_X1 U22894 ( .A1(n19876), .A2(n20024), .B1(n20023), .B2(n19875), .ZN(
        n19868) );
  AOI22_X1 U22895 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19878), .B1(
        n19877), .B2(n20026), .ZN(n19867) );
  OAI211_X1 U22896 ( .C1(n19891), .C2(n19881), .A(n19868), .B(n19867), .ZN(
        P2_U3131) );
  AOI22_X1 U22897 ( .A1(n19876), .A2(n20030), .B1(n9671), .B2(n19875), .ZN(
        n19870) );
  AOI22_X1 U22898 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19878), .B1(
        n19877), .B2(n20032), .ZN(n19869) );
  OAI211_X1 U22899 ( .C1(n19894), .C2(n19881), .A(n19870), .B(n19869), .ZN(
        P2_U3132) );
  AOI22_X1 U22900 ( .A1(n19876), .A2(n20037), .B1(n20036), .B2(n19875), .ZN(
        n19872) );
  AOI22_X1 U22901 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19878), .B1(
        n19877), .B2(n20039), .ZN(n19871) );
  OAI211_X1 U22902 ( .C1(n19897), .C2(n19881), .A(n19872), .B(n19871), .ZN(
        P2_U3133) );
  AOI22_X1 U22903 ( .A1(n19876), .A2(n20043), .B1(n20042), .B2(n19875), .ZN(
        n19874) );
  AOI22_X1 U22904 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19878), .B1(
        n19877), .B2(n20045), .ZN(n19873) );
  OAI211_X1 U22905 ( .C1(n19901), .C2(n19881), .A(n19874), .B(n19873), .ZN(
        P2_U3134) );
  AOI22_X1 U22906 ( .A1(n19876), .A2(n20050), .B1(n20048), .B2(n19875), .ZN(
        n19880) );
  AOI22_X1 U22907 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19878), .B1(
        n19877), .B2(n20054), .ZN(n19879) );
  OAI211_X1 U22908 ( .C1(n19882), .C2(n19881), .A(n19880), .B(n19879), .ZN(
        P2_U3135) );
  INV_X1 U22909 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n19885) );
  AOI22_X1 U22910 ( .A1(n19903), .A2(n20003), .B1(n20002), .B2(n19902), .ZN(
        n19884) );
  AOI22_X1 U22911 ( .A1(n19914), .A2(n20005), .B1(n19904), .B2(n20004), .ZN(
        n19883) );
  OAI211_X1 U22912 ( .C1(n19908), .C2(n19885), .A(n19884), .B(n19883), .ZN(
        P2_U3136) );
  AOI22_X1 U22913 ( .A1(n19903), .A2(n20017), .B1(n19902), .B2(n20016), .ZN(
        n19887) );
  AOI22_X1 U22914 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19898), .B1(
        n19904), .B2(n20019), .ZN(n19886) );
  OAI211_X1 U22915 ( .C1(n19888), .C2(n19947), .A(n19887), .B(n19886), .ZN(
        P2_U3138) );
  AOI22_X1 U22916 ( .A1(n19903), .A2(n20024), .B1(n19902), .B2(n20023), .ZN(
        n19890) );
  AOI22_X1 U22917 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19898), .B1(
        n19904), .B2(n20026), .ZN(n19889) );
  OAI211_X1 U22918 ( .C1(n19891), .C2(n19947), .A(n19890), .B(n19889), .ZN(
        P2_U3139) );
  AOI22_X1 U22919 ( .A1(n19903), .A2(n20030), .B1(n19902), .B2(n9671), .ZN(
        n19893) );
  AOI22_X1 U22920 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19898), .B1(
        n19904), .B2(n20032), .ZN(n19892) );
  OAI211_X1 U22921 ( .C1(n19894), .C2(n19947), .A(n19893), .B(n19892), .ZN(
        P2_U3140) );
  AOI22_X1 U22922 ( .A1(n19903), .A2(n20037), .B1(n19902), .B2(n20036), .ZN(
        n19896) );
  AOI22_X1 U22923 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19898), .B1(
        n19904), .B2(n20039), .ZN(n19895) );
  OAI211_X1 U22924 ( .C1(n19897), .C2(n19947), .A(n19896), .B(n19895), .ZN(
        P2_U3141) );
  AOI22_X1 U22925 ( .A1(n19903), .A2(n20043), .B1(n19902), .B2(n20042), .ZN(
        n19900) );
  AOI22_X1 U22926 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19898), .B1(
        n19904), .B2(n20045), .ZN(n19899) );
  OAI211_X1 U22927 ( .C1(n19901), .C2(n19947), .A(n19900), .B(n19899), .ZN(
        P2_U3142) );
  INV_X1 U22928 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n19907) );
  AOI22_X1 U22929 ( .A1(n19903), .A2(n20050), .B1(n19902), .B2(n20048), .ZN(
        n19906) );
  AOI22_X1 U22930 ( .A1(n19904), .A2(n20054), .B1(n19914), .B2(n20052), .ZN(
        n19905) );
  OAI211_X1 U22931 ( .C1(n19908), .C2(n19907), .A(n19906), .B(n19905), .ZN(
        P2_U3143) );
  NAND2_X1 U22932 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19909), .ZN(
        n19917) );
  OR2_X1 U22933 ( .A1(n19917), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19913) );
  INV_X1 U22934 ( .A(n19910), .ZN(n19912) );
  NOR2_X1 U22935 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19911), .ZN(
        n19942) );
  NOR3_X1 U22936 ( .A1(n19912), .A2(n19942), .A3(n20065), .ZN(n19916) );
  AOI21_X1 U22937 ( .B1(n20065), .B2(n19913), .A(n19916), .ZN(n19943) );
  AOI22_X1 U22938 ( .A1(n19943), .A2(n20003), .B1(n20002), .B2(n19942), .ZN(
        n19922) );
  OAI21_X1 U22939 ( .B1(n19914), .B2(n19966), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19918) );
  AOI211_X1 U22940 ( .C1(n19918), .C2(n19917), .A(n19916), .B(n19915), .ZN(
        n19919) );
  AOI22_X1 U22941 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19944), .B1(
        n19966), .B2(n20005), .ZN(n19921) );
  OAI211_X1 U22942 ( .C1(n19923), .C2(n19947), .A(n19922), .B(n19921), .ZN(
        P2_U3144) );
  AOI22_X1 U22943 ( .A1(n19943), .A2(n20010), .B1(n20009), .B2(n19942), .ZN(
        n19925) );
  AOI22_X1 U22944 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19944), .B1(
        n19966), .B2(n20011), .ZN(n19924) );
  OAI211_X1 U22945 ( .C1(n19926), .C2(n19947), .A(n19925), .B(n19924), .ZN(
        P2_U3145) );
  AOI22_X1 U22946 ( .A1(n19943), .A2(n20017), .B1(n20016), .B2(n19942), .ZN(
        n19928) );
  AOI22_X1 U22947 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19944), .B1(
        n19966), .B2(n20018), .ZN(n19927) );
  OAI211_X1 U22948 ( .C1(n19929), .C2(n19947), .A(n19928), .B(n19927), .ZN(
        P2_U3146) );
  AOI22_X1 U22949 ( .A1(n19943), .A2(n20024), .B1(n20023), .B2(n19942), .ZN(
        n19931) );
  AOI22_X1 U22950 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19944), .B1(
        n19966), .B2(n20025), .ZN(n19930) );
  OAI211_X1 U22951 ( .C1(n19932), .C2(n19947), .A(n19931), .B(n19930), .ZN(
        P2_U3147) );
  AOI22_X1 U22952 ( .A1(n19943), .A2(n20030), .B1(n9671), .B2(n19942), .ZN(
        n19934) );
  AOI22_X1 U22953 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19944), .B1(
        n19966), .B2(n20031), .ZN(n19933) );
  OAI211_X1 U22954 ( .C1(n19935), .C2(n19947), .A(n19934), .B(n19933), .ZN(
        P2_U3148) );
  AOI22_X1 U22955 ( .A1(n19943), .A2(n20037), .B1(n20036), .B2(n19942), .ZN(
        n19937) );
  AOI22_X1 U22956 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19944), .B1(
        n19966), .B2(n20038), .ZN(n19936) );
  OAI211_X1 U22957 ( .C1(n19938), .C2(n19947), .A(n19937), .B(n19936), .ZN(
        P2_U3149) );
  AOI22_X1 U22958 ( .A1(n19943), .A2(n20043), .B1(n20042), .B2(n19942), .ZN(
        n19940) );
  AOI22_X1 U22959 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19944), .B1(
        n19966), .B2(n20044), .ZN(n19939) );
  OAI211_X1 U22960 ( .C1(n19941), .C2(n19947), .A(n19940), .B(n19939), .ZN(
        P2_U3150) );
  AOI22_X1 U22961 ( .A1(n19943), .A2(n20050), .B1(n20048), .B2(n19942), .ZN(
        n19946) );
  AOI22_X1 U22962 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19944), .B1(
        n19966), .B2(n20052), .ZN(n19945) );
  OAI211_X1 U22963 ( .C1(n19948), .C2(n19947), .A(n19946), .B(n19945), .ZN(
        P2_U3151) );
  INV_X1 U22964 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n19951) );
  AOI22_X1 U22965 ( .A1(n19965), .A2(n20010), .B1(n19964), .B2(n20009), .ZN(
        n19950) );
  AOI22_X1 U22966 ( .A1(n19966), .A2(n20012), .B1(n19985), .B2(n20011), .ZN(
        n19949) );
  OAI211_X1 U22967 ( .C1(n19970), .C2(n19951), .A(n19950), .B(n19949), .ZN(
        P2_U3153) );
  INV_X1 U22968 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n19954) );
  AOI22_X1 U22969 ( .A1(n19965), .A2(n20017), .B1(n19964), .B2(n20016), .ZN(
        n19953) );
  AOI22_X1 U22970 ( .A1(n19966), .A2(n20019), .B1(n19985), .B2(n20018), .ZN(
        n19952) );
  OAI211_X1 U22971 ( .C1(n19970), .C2(n19954), .A(n19953), .B(n19952), .ZN(
        P2_U3154) );
  AOI22_X1 U22972 ( .A1(n19965), .A2(n20024), .B1(n19964), .B2(n20023), .ZN(
        n19956) );
  AOI22_X1 U22973 ( .A1(n19966), .A2(n20026), .B1(n19985), .B2(n20025), .ZN(
        n19955) );
  OAI211_X1 U22974 ( .C1(n19970), .C2(n12006), .A(n19956), .B(n19955), .ZN(
        P2_U3155) );
  INV_X1 U22975 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n19959) );
  AOI22_X1 U22976 ( .A1(n19965), .A2(n20030), .B1(n19964), .B2(n9671), .ZN(
        n19958) );
  AOI22_X1 U22977 ( .A1(n19966), .A2(n20032), .B1(n19985), .B2(n20031), .ZN(
        n19957) );
  OAI211_X1 U22978 ( .C1(n19970), .C2(n19959), .A(n19958), .B(n19957), .ZN(
        P2_U3156) );
  AOI22_X1 U22979 ( .A1(n19965), .A2(n20037), .B1(n19964), .B2(n20036), .ZN(
        n19961) );
  AOI22_X1 U22980 ( .A1(n19966), .A2(n20039), .B1(n19985), .B2(n20038), .ZN(
        n19960) );
  OAI211_X1 U22981 ( .C1(n19970), .C2(n12636), .A(n19961), .B(n19960), .ZN(
        P2_U3157) );
  AOI22_X1 U22982 ( .A1(n19965), .A2(n20043), .B1(n19964), .B2(n20042), .ZN(
        n19963) );
  AOI22_X1 U22983 ( .A1(n19966), .A2(n20045), .B1(n19985), .B2(n20044), .ZN(
        n19962) );
  OAI211_X1 U22984 ( .C1(n19970), .C2(n12073), .A(n19963), .B(n19962), .ZN(
        P2_U3158) );
  INV_X1 U22985 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n19969) );
  AOI22_X1 U22986 ( .A1(n19965), .A2(n20050), .B1(n19964), .B2(n20048), .ZN(
        n19968) );
  AOI22_X1 U22987 ( .A1(n19966), .A2(n20054), .B1(n19985), .B2(n20052), .ZN(
        n19967) );
  OAI211_X1 U22988 ( .C1(n19970), .C2(n19969), .A(n19968), .B(n19967), .ZN(
        P2_U3159) );
  INV_X1 U22989 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n19973) );
  AOI22_X1 U22990 ( .A1(n20011), .A2(n20055), .B1(n20009), .B2(n19984), .ZN(
        n19972) );
  AOI22_X1 U22991 ( .A1(n20010), .A2(n19986), .B1(n19985), .B2(n20012), .ZN(
        n19971) );
  OAI211_X1 U22992 ( .C1(n19990), .C2(n19973), .A(n19972), .B(n19971), .ZN(
        P2_U3161) );
  INV_X1 U22993 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n19976) );
  AOI22_X1 U22994 ( .A1(n20019), .A2(n19985), .B1(n19984), .B2(n20016), .ZN(
        n19975) );
  AOI22_X1 U22995 ( .A1(n20017), .A2(n19986), .B1(n20055), .B2(n20018), .ZN(
        n19974) );
  OAI211_X1 U22996 ( .C1(n19990), .C2(n19976), .A(n19975), .B(n19974), .ZN(
        P2_U3162) );
  AOI22_X1 U22997 ( .A1(n20025), .A2(n20055), .B1(n19984), .B2(n20023), .ZN(
        n19978) );
  AOI22_X1 U22998 ( .A1(n20024), .A2(n19986), .B1(n19985), .B2(n20026), .ZN(
        n19977) );
  OAI211_X1 U22999 ( .C1(n19990), .C2(n12002), .A(n19978), .B(n19977), .ZN(
        P2_U3163) );
  INV_X1 U23000 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n19981) );
  AOI22_X1 U23001 ( .A1(n20032), .A2(n19985), .B1(n19984), .B2(n9671), .ZN(
        n19980) );
  AOI22_X1 U23002 ( .A1(n20030), .A2(n19986), .B1(n20055), .B2(n20031), .ZN(
        n19979) );
  OAI211_X1 U23003 ( .C1(n19990), .C2(n19981), .A(n19980), .B(n19979), .ZN(
        P2_U3164) );
  AOI22_X1 U23004 ( .A1(n20045), .A2(n19985), .B1(n19984), .B2(n20042), .ZN(
        n19983) );
  AOI22_X1 U23005 ( .A1(n20043), .A2(n19986), .B1(n20055), .B2(n20044), .ZN(
        n19982) );
  OAI211_X1 U23006 ( .C1(n19990), .C2(n12061), .A(n19983), .B(n19982), .ZN(
        P2_U3166) );
  INV_X1 U23007 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n19989) );
  AOI22_X1 U23008 ( .A1(n20052), .A2(n20055), .B1(n19984), .B2(n20048), .ZN(
        n19988) );
  AOI22_X1 U23009 ( .A1(n20050), .A2(n19986), .B1(n19985), .B2(n20054), .ZN(
        n19987) );
  OAI211_X1 U23010 ( .C1(n19990), .C2(n19989), .A(n19988), .B(n19987), .ZN(
        P2_U3167) );
  NOR2_X1 U23011 ( .A1(n20156), .A2(n19991), .ZN(n19998) );
  AOI21_X1 U23012 ( .B1(n19992), .B2(n20151), .A(n19998), .ZN(n19997) );
  INV_X1 U23013 ( .A(n19993), .ZN(n20049) );
  AND2_X1 U23014 ( .A1(n19993), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19994) );
  NAND2_X1 U23015 ( .A1(n12009), .A2(n19994), .ZN(n20001) );
  OAI211_X1 U23016 ( .C1(n20049), .C2(n19920), .A(n20001), .B(n19995), .ZN(
        n19996) );
  INV_X1 U23017 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n20008) );
  INV_X1 U23018 ( .A(n19998), .ZN(n19999) );
  OAI21_X1 U23019 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19999), .A(n20065), 
        .ZN(n20000) );
  AND2_X1 U23020 ( .A1(n20001), .A2(n20000), .ZN(n20051) );
  AOI22_X1 U23021 ( .A1(n20051), .A2(n20003), .B1(n20049), .B2(n20002), .ZN(
        n20007) );
  AOI22_X1 U23022 ( .A1(n20053), .A2(n20005), .B1(n20055), .B2(n20004), .ZN(
        n20006) );
  OAI211_X1 U23023 ( .C1(n20059), .C2(n20008), .A(n20007), .B(n20006), .ZN(
        P2_U3168) );
  INV_X1 U23024 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n20015) );
  AOI22_X1 U23025 ( .A1(n20051), .A2(n20010), .B1(n20049), .B2(n20009), .ZN(
        n20014) );
  AOI22_X1 U23026 ( .A1(n20055), .A2(n20012), .B1(n20053), .B2(n20011), .ZN(
        n20013) );
  OAI211_X1 U23027 ( .C1(n20059), .C2(n20015), .A(n20014), .B(n20013), .ZN(
        P2_U3169) );
  INV_X1 U23028 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n20022) );
  AOI22_X1 U23029 ( .A1(n20051), .A2(n20017), .B1(n20049), .B2(n20016), .ZN(
        n20021) );
  AOI22_X1 U23030 ( .A1(n20055), .A2(n20019), .B1(n20053), .B2(n20018), .ZN(
        n20020) );
  OAI211_X1 U23031 ( .C1(n20059), .C2(n20022), .A(n20021), .B(n20020), .ZN(
        P2_U3170) );
  AOI22_X1 U23032 ( .A1(n20051), .A2(n20024), .B1(n20049), .B2(n20023), .ZN(
        n20028) );
  AOI22_X1 U23033 ( .A1(n20055), .A2(n20026), .B1(n20053), .B2(n20025), .ZN(
        n20027) );
  OAI211_X1 U23034 ( .C1(n20059), .C2(n12008), .A(n20028), .B(n20027), .ZN(
        P2_U3171) );
  AOI22_X1 U23035 ( .A1(n20051), .A2(n20030), .B1(n20049), .B2(n9671), .ZN(
        n20034) );
  AOI22_X1 U23036 ( .A1(n20055), .A2(n20032), .B1(n20053), .B2(n20031), .ZN(
        n20033) );
  OAI211_X1 U23037 ( .C1(n20059), .C2(n20035), .A(n20034), .B(n20033), .ZN(
        P2_U3172) );
  AOI22_X1 U23038 ( .A1(n20051), .A2(n20037), .B1(n20049), .B2(n20036), .ZN(
        n20041) );
  AOI22_X1 U23039 ( .A1(n20055), .A2(n20039), .B1(n20053), .B2(n20038), .ZN(
        n20040) );
  OAI211_X1 U23040 ( .C1(n20059), .C2(n12634), .A(n20041), .B(n20040), .ZN(
        P2_U3173) );
  AOI22_X1 U23041 ( .A1(n20051), .A2(n20043), .B1(n20049), .B2(n20042), .ZN(
        n20047) );
  AOI22_X1 U23042 ( .A1(n20055), .A2(n20045), .B1(n20053), .B2(n20044), .ZN(
        n20046) );
  OAI211_X1 U23043 ( .C1(n20059), .C2(n12070), .A(n20047), .B(n20046), .ZN(
        P2_U3174) );
  INV_X1 U23044 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n20058) );
  AOI22_X1 U23045 ( .A1(n20051), .A2(n20050), .B1(n20049), .B2(n20048), .ZN(
        n20057) );
  AOI22_X1 U23046 ( .A1(n20055), .A2(n20054), .B1(n20053), .B2(n20052), .ZN(
        n20056) );
  OAI211_X1 U23047 ( .C1(n20059), .C2(n20058), .A(n20057), .B(n20056), .ZN(
        P2_U3175) );
  INV_X1 U23048 ( .A(n20060), .ZN(n20062) );
  AOI21_X1 U23049 ( .B1(n20063), .B2(n20062), .A(n20061), .ZN(n20072) );
  INV_X1 U23050 ( .A(n20064), .ZN(n20069) );
  NAND2_X1 U23051 ( .A1(n20196), .A2(n20065), .ZN(n20066) );
  NAND4_X1 U23052 ( .A1(n20069), .A2(n20068), .A3(n20067), .A4(n20066), .ZN(
        n20070) );
  OAI211_X1 U23053 ( .C1(n20072), .C2(n15777), .A(n20071), .B(n20070), .ZN(
        P2_U3177) );
  AND2_X1 U23054 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20073), .ZN(
        P2_U3179) );
  AND2_X1 U23055 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20073), .ZN(
        P2_U3180) );
  AND2_X1 U23056 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20073), .ZN(
        P2_U3181) );
  AND2_X1 U23057 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20073), .ZN(
        P2_U3182) );
  AND2_X1 U23058 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20073), .ZN(
        P2_U3183) );
  AND2_X1 U23059 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20073), .ZN(
        P2_U3184) );
  AND2_X1 U23060 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20073), .ZN(
        P2_U3185) );
  AND2_X1 U23061 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20073), .ZN(
        P2_U3186) );
  AND2_X1 U23062 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20073), .ZN(
        P2_U3187) );
  AND2_X1 U23063 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20073), .ZN(
        P2_U3188) );
  AND2_X1 U23064 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20073), .ZN(
        P2_U3189) );
  AND2_X1 U23065 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20073), .ZN(
        P2_U3190) );
  AND2_X1 U23066 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20073), .ZN(
        P2_U3191) );
  AND2_X1 U23067 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20073), .ZN(
        P2_U3192) );
  AND2_X1 U23068 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20073), .ZN(
        P2_U3193) );
  AND2_X1 U23069 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20073), .ZN(
        P2_U3194) );
  AND2_X1 U23070 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20073), .ZN(
        P2_U3195) );
  AND2_X1 U23071 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20073), .ZN(
        P2_U3196) );
  AND2_X1 U23072 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20073), .ZN(
        P2_U3197) );
  AND2_X1 U23073 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20073), .ZN(
        P2_U3198) );
  AND2_X1 U23074 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20073), .ZN(
        P2_U3199) );
  AND2_X1 U23075 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20073), .ZN(
        P2_U3200) );
  AND2_X1 U23076 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20073), .ZN(P2_U3201) );
  AND2_X1 U23077 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20073), .ZN(P2_U3202) );
  AND2_X1 U23078 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20073), .ZN(P2_U3203) );
  AND2_X1 U23079 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20073), .ZN(P2_U3204) );
  AND2_X1 U23080 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20073), .ZN(P2_U3205) );
  AND2_X1 U23081 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20073), .ZN(P2_U3206) );
  AND2_X1 U23082 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20073), .ZN(P2_U3207) );
  AND2_X1 U23083 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20073), .ZN(P2_U3208) );
  NAND2_X1 U23084 ( .A1(n20196), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20082) );
  INV_X1 U23085 ( .A(n20082), .ZN(n20087) );
  INV_X1 U23086 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20077) );
  NOR3_X1 U23087 ( .A1(n20087), .A2(n20077), .A3(n20074), .ZN(n20076) );
  OAI211_X1 U23088 ( .C1(HOLD), .C2(n20077), .A(n20213), .B(n20083), .ZN(
        n20075) );
  NAND2_X1 U23089 ( .A1(NA), .A2(n20078), .ZN(n20085) );
  OAI211_X1 U23090 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n20076), .A(n20075), 
        .B(n20085), .ZN(P2_U3209) );
  NAND2_X1 U23091 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20819), .ZN(n20086) );
  AOI211_X1 U23092 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n20086), .A(n20078), 
        .B(n20077), .ZN(n20079) );
  NOR3_X1 U23093 ( .A1(n20208), .A2(n20087), .A3(n20079), .ZN(n20080) );
  OAI21_X1 U23094 ( .B1(n20819), .B2(n20081), .A(n20080), .ZN(P2_U3210) );
  OAI22_X1 U23095 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n20083), .B1(NA), 
        .B2(n20082), .ZN(n20084) );
  OAI211_X1 U23096 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20084), .ZN(n20089) );
  OAI211_X1 U23097 ( .C1(n20087), .C2(n20086), .A(P2_STATE_REG_2__SCAN_IN), 
        .B(n20085), .ZN(n20088) );
  NAND2_X1 U23098 ( .A1(n20089), .A2(n20088), .ZN(P2_U3211) );
  NAND2_X1 U23099 ( .A1(n20216), .A2(n20090), .ZN(n20136) );
  OAI222_X1 U23100 ( .A1(n20131), .A2(n10734), .B1(n20091), .B2(n20216), .C1(
        n10673), .C2(n20132), .ZN(P2_U3212) );
  OAI222_X1 U23101 ( .A1(n20132), .A2(n10734), .B1(n20092), .B2(n20216), .C1(
        n14034), .C2(n20131), .ZN(P2_U3213) );
  OAI222_X1 U23102 ( .A1(n20132), .A2(n14034), .B1(n20093), .B2(n20216), .C1(
        n10753), .C2(n20131), .ZN(P2_U3214) );
  OAI222_X1 U23103 ( .A1(n20136), .A2(n10760), .B1(n20094), .B2(n20216), .C1(
        n10753), .C2(n20132), .ZN(P2_U3215) );
  OAI222_X1 U23104 ( .A1(n20136), .A2(n20096), .B1(n20095), .B2(n20216), .C1(
        n10760), .C2(n20132), .ZN(P2_U3216) );
  OAI222_X1 U23105 ( .A1(n20136), .A2(n20098), .B1(n20097), .B2(n20216), .C1(
        n20096), .C2(n20132), .ZN(P2_U3217) );
  OAI222_X1 U23106 ( .A1(n20136), .A2(n10767), .B1(n20099), .B2(n20216), .C1(
        n20098), .C2(n20132), .ZN(P2_U3218) );
  OAI222_X1 U23107 ( .A1(n20136), .A2(n15185), .B1(n20100), .B2(n20216), .C1(
        n10767), .C2(n20132), .ZN(P2_U3219) );
  OAI222_X1 U23108 ( .A1(n20131), .A2(n10777), .B1(n20101), .B2(n20216), .C1(
        n15185), .C2(n20132), .ZN(P2_U3220) );
  OAI222_X1 U23109 ( .A1(n20131), .A2(n10783), .B1(n20102), .B2(n20216), .C1(
        n10777), .C2(n20132), .ZN(P2_U3221) );
  OAI222_X1 U23110 ( .A1(n20131), .A2(n20104), .B1(n20103), .B2(n20216), .C1(
        n10783), .C2(n20132), .ZN(P2_U3222) );
  OAI222_X1 U23111 ( .A1(n20131), .A2(n20106), .B1(n20105), .B2(n20216), .C1(
        n20104), .C2(n20132), .ZN(P2_U3223) );
  OAI222_X1 U23112 ( .A1(n20131), .A2(n10793), .B1(n20107), .B2(n20216), .C1(
        n20106), .C2(n20132), .ZN(P2_U3224) );
  OAI222_X1 U23113 ( .A1(n20131), .A2(n10668), .B1(n20108), .B2(n20216), .C1(
        n10793), .C2(n20132), .ZN(P2_U3225) );
  OAI222_X1 U23114 ( .A1(n20136), .A2(n15684), .B1(n20109), .B2(n20216), .C1(
        n10668), .C2(n20132), .ZN(P2_U3226) );
  OAI222_X1 U23115 ( .A1(n20136), .A2(n15672), .B1(n20110), .B2(n20216), .C1(
        n15684), .C2(n20132), .ZN(P2_U3227) );
  OAI222_X1 U23116 ( .A1(n20136), .A2(n20112), .B1(n20111), .B2(n20216), .C1(
        n15672), .C2(n20132), .ZN(P2_U3228) );
  OAI222_X1 U23117 ( .A1(n20136), .A2(n15493), .B1(n20113), .B2(n20216), .C1(
        n20112), .C2(n20132), .ZN(P2_U3229) );
  OAI222_X1 U23118 ( .A1(n20136), .A2(n20115), .B1(n20114), .B2(n20216), .C1(
        n15493), .C2(n20132), .ZN(P2_U3230) );
  INV_X1 U23119 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20117) );
  OAI222_X1 U23120 ( .A1(n20136), .A2(n20117), .B1(n20116), .B2(n20216), .C1(
        n20115), .C2(n20132), .ZN(P2_U3231) );
  OAI222_X1 U23121 ( .A1(n20131), .A2(n10816), .B1(n20118), .B2(n20216), .C1(
        n20117), .C2(n20132), .ZN(P2_U3232) );
  OAI222_X1 U23122 ( .A1(n20131), .A2(n10662), .B1(n20119), .B2(n20216), .C1(
        n10816), .C2(n20132), .ZN(P2_U3233) );
  OAI222_X1 U23123 ( .A1(n20131), .A2(n10820), .B1(n20120), .B2(n20216), .C1(
        n10662), .C2(n20132), .ZN(P2_U3234) );
  OAI222_X1 U23124 ( .A1(n20131), .A2(n20122), .B1(n20121), .B2(n20216), .C1(
        n10820), .C2(n20132), .ZN(P2_U3235) );
  OAI222_X1 U23125 ( .A1(n20131), .A2(n20124), .B1(n20123), .B2(n20216), .C1(
        n20122), .C2(n20132), .ZN(P2_U3236) );
  INV_X1 U23126 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20127) );
  OAI222_X1 U23127 ( .A1(n20131), .A2(n20127), .B1(n20125), .B2(n20216), .C1(
        n20124), .C2(n20132), .ZN(P2_U3237) );
  OAI222_X1 U23128 ( .A1(n20132), .A2(n20127), .B1(n20126), .B2(n20216), .C1(
        n20128), .C2(n20131), .ZN(P2_U3238) );
  OAI222_X1 U23129 ( .A1(n20131), .A2(n10841), .B1(n20129), .B2(n20216), .C1(
        n20128), .C2(n20132), .ZN(P2_U3239) );
  OAI222_X1 U23130 ( .A1(n20131), .A2(n20133), .B1(n20130), .B2(n20216), .C1(
        n10841), .C2(n20132), .ZN(P2_U3240) );
  INV_X1 U23131 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20134) );
  OAI222_X1 U23132 ( .A1(n20136), .A2(n20135), .B1(n20134), .B2(n20216), .C1(
        n20133), .C2(n20132), .ZN(P2_U3241) );
  INV_X1 U23133 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20137) );
  AOI22_X1 U23134 ( .A1(n20216), .A2(n20138), .B1(n20137), .B2(n20213), .ZN(
        P2_U3585) );
  MUX2_X1 U23135 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20216), .Z(P2_U3586) );
  INV_X1 U23136 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20139) );
  AOI22_X1 U23137 ( .A1(n20216), .A2(n20140), .B1(n20139), .B2(n20213), .ZN(
        P2_U3587) );
  INV_X1 U23138 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20141) );
  AOI22_X1 U23139 ( .A1(n20216), .A2(n20142), .B1(n20141), .B2(n20213), .ZN(
        P2_U3588) );
  OAI21_X1 U23140 ( .B1(n20146), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20144), 
        .ZN(n20143) );
  INV_X1 U23141 ( .A(n20143), .ZN(P2_U3591) );
  OAI21_X1 U23142 ( .B1(n20146), .B2(n20145), .A(n20144), .ZN(P2_U3592) );
  INV_X1 U23143 ( .A(n20147), .ZN(n20149) );
  OAI211_X1 U23144 ( .C1(n20151), .C2(n20150), .A(n20149), .B(n20148), .ZN(
        n20160) );
  AOI222_X1 U23145 ( .A1(n20160), .A2(n20154), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20153), .C1(n20157), .C2(n20152), .ZN(n20155) );
  AOI22_X1 U23146 ( .A1(n20180), .A2(n20156), .B1(n20155), .B2(n20181), .ZN(
        P2_U3602) );
  NAND2_X1 U23147 ( .A1(n20157), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20168) );
  OAI21_X1 U23148 ( .B1(n20166), .B2(n20168), .A(n20158), .ZN(n20159) );
  AOI22_X1 U23149 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20161), .B1(n20160), 
        .B2(n20159), .ZN(n20162) );
  AOI22_X1 U23150 ( .A1(n20180), .A2(n20163), .B1(n20162), .B2(n20181), .ZN(
        P2_U3603) );
  INV_X1 U23151 ( .A(n20164), .ZN(n20176) );
  OR3_X1 U23152 ( .A1(n20166), .A2(n20176), .A3(n20165), .ZN(n20167) );
  OAI21_X1 U23153 ( .B1(n20169), .B2(n20168), .A(n20167), .ZN(n20170) );
  AOI21_X1 U23154 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20171), .A(n20170), 
        .ZN(n20172) );
  AOI22_X1 U23155 ( .A1(n20180), .A2(n10356), .B1(n20172), .B2(n20181), .ZN(
        P2_U3604) );
  INV_X1 U23156 ( .A(n20173), .ZN(n20175) );
  OAI22_X1 U23157 ( .A1(n20177), .A2(n20176), .B1(n20175), .B2(n20174), .ZN(
        n20178) );
  AOI21_X1 U23158 ( .B1(n20182), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20178), 
        .ZN(n20179) );
  OAI22_X1 U23159 ( .A1(n20182), .A2(n20181), .B1(n20180), .B2(n20179), .ZN(
        P2_U3605) );
  INV_X1 U23160 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20183) );
  AOI22_X1 U23161 ( .A1(n20216), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20183), 
        .B2(n20213), .ZN(P2_U3608) );
  NAND2_X1 U23162 ( .A1(n20185), .A2(n20184), .ZN(n20188) );
  AOI22_X1 U23163 ( .A1(n20189), .A2(n20188), .B1(n20187), .B2(n20186), .ZN(
        n20190) );
  NAND2_X1 U23164 ( .A1(n20191), .A2(n20190), .ZN(n20193) );
  MUX2_X1 U23165 ( .A(P2_MORE_REG_SCAN_IN), .B(n20193), .S(n20192), .Z(
        P2_U3609) );
  OAI22_X1 U23166 ( .A1(n20196), .A2(n20195), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20194), .ZN(n20197) );
  NOR2_X1 U23167 ( .A1(n20198), .A2(n20197), .ZN(n20212) );
  NAND3_X1 U23168 ( .A1(n20199), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10648), 
        .ZN(n20207) );
  AOI21_X1 U23169 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n20208), .A(n20201), 
        .ZN(n20204) );
  AOI22_X1 U23170 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20202), .B1(n20201), 
        .B2(n20200), .ZN(n20203) );
  AOI21_X1 U23171 ( .B1(n20205), .B2(n20204), .A(n20203), .ZN(n20206) );
  OAI21_X1 U23172 ( .B1(n20208), .B2(n20207), .A(n20206), .ZN(n20209) );
  INV_X1 U23173 ( .A(n20209), .ZN(n20211) );
  NAND2_X1 U23174 ( .A1(n20212), .A2(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20210) );
  OAI21_X1 U23175 ( .B1(n20212), .B2(n20211), .A(n20210), .ZN(P2_U3610) );
  INV_X1 U23176 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n20214) );
  AOI22_X1 U23177 ( .A1(n20216), .A2(n20215), .B1(n20214), .B2(n20213), .ZN(
        P2_U3611) );
  AOI21_X1 U23178 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n10997), .A(n20814), 
        .ZN(n20817) );
  INV_X1 U23179 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20217) );
  NAND2_X1 U23180 ( .A1(n20814), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20916) );
  AOI21_X1 U23181 ( .B1(n20817), .B2(n20217), .A(n20875), .ZN(P1_U2802) );
  INV_X1 U23182 ( .A(n20218), .ZN(n20220) );
  OAI21_X1 U23183 ( .B1(n20220), .B2(n20219), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20221) );
  OAI21_X1 U23184 ( .B1(n20223), .B2(n20222), .A(n20221), .ZN(P1_U2803) );
  INV_X1 U23185 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n21061) );
  NOR2_X1 U23186 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20225) );
  NOR2_X1 U23187 ( .A1(n20875), .A2(n20225), .ZN(n20224) );
  AOI22_X1 U23188 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n20875), .B1(n21061), 
        .B2(n20224), .ZN(P1_U2804) );
  OAI21_X1 U23189 ( .B1(BS16), .B2(n20225), .A(n20884), .ZN(n20882) );
  OAI21_X1 U23190 ( .B1(n20884), .B2(n21095), .A(n20882), .ZN(P1_U2805) );
  OAI21_X1 U23191 ( .B1(n20227), .B2(n20957), .A(n20226), .ZN(P1_U2806) );
  NOR4_X1 U23192 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20231) );
  NOR4_X1 U23193 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20230) );
  NOR4_X1 U23194 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20229) );
  NOR4_X1 U23195 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20228) );
  NAND4_X1 U23196 ( .A1(n20231), .A2(n20230), .A3(n20229), .A4(n20228), .ZN(
        n20237) );
  NOR4_X1 U23197 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20235) );
  AOI211_X1 U23198 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20234) );
  NOR4_X1 U23199 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20233) );
  NOR4_X1 U23200 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20232) );
  NAND4_X1 U23201 ( .A1(n20235), .A2(n20234), .A3(n20233), .A4(n20232), .ZN(
        n20236) );
  NOR2_X1 U23202 ( .A1(n20237), .A2(n20236), .ZN(n20903) );
  INV_X1 U23203 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20877) );
  NOR3_X1 U23204 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20239) );
  OAI21_X1 U23205 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20239), .A(n20903), .ZN(
        n20238) );
  OAI21_X1 U23206 ( .B1(n20903), .B2(n20877), .A(n20238), .ZN(P1_U2807) );
  INV_X1 U23207 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20883) );
  AOI21_X1 U23208 ( .B1(n20898), .B2(n20883), .A(n20239), .ZN(n20240) );
  INV_X1 U23209 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20969) );
  INV_X1 U23210 ( .A(n20903), .ZN(n20900) );
  AOI22_X1 U23211 ( .A1(n20903), .A2(n20240), .B1(n20969), .B2(n20900), .ZN(
        P1_U2808) );
  AOI21_X1 U23212 ( .B1(n20306), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n20288), .ZN(n20243) );
  NAND3_X1 U23213 ( .A1(n20309), .A2(n20241), .A3(n20837), .ZN(n20242) );
  OAI211_X1 U23214 ( .C1(n20244), .C2(n20274), .A(n20243), .B(n20242), .ZN(
        n20245) );
  AOI21_X1 U23215 ( .B1(P1_EBX_REG_9__SCAN_IN), .B2(n20304), .A(n20245), .ZN(
        n20249) );
  AOI22_X1 U23216 ( .A1(n20247), .A2(n20268), .B1(n20307), .B2(n20246), .ZN(
        n20248) );
  OAI211_X1 U23217 ( .C1(n20250), .C2(n20837), .A(n20249), .B(n20248), .ZN(
        P1_U2831) );
  NAND2_X1 U23218 ( .A1(n20309), .A2(n20258), .ZN(n20275) );
  NAND2_X1 U23219 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20257) );
  NOR3_X1 U23220 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20275), .A3(n20257), .ZN(
        n20256) );
  AOI22_X1 U23221 ( .A1(P1_EBX_REG_7__SCAN_IN), .A2(n20304), .B1(n20303), .B2(
        n20251), .ZN(n20252) );
  OAI211_X1 U23222 ( .C1(n20254), .C2(n20253), .A(n20252), .B(n20276), .ZN(
        n20255) );
  NOR2_X1 U23223 ( .A1(n20256), .A2(n20255), .ZN(n20263) );
  INV_X1 U23224 ( .A(n20257), .ZN(n20260) );
  NOR2_X1 U23225 ( .A1(n20258), .A2(n20259), .ZN(n20283) );
  NOR2_X1 U23226 ( .A1(n20301), .A2(n20283), .ZN(n20291) );
  OAI21_X1 U23227 ( .B1(n20260), .B2(n20259), .A(n20291), .ZN(n20269) );
  AOI22_X1 U23228 ( .A1(n20268), .A2(n20261), .B1(n20269), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n20262) );
  OAI211_X1 U23229 ( .C1(n20264), .C2(n20292), .A(n20263), .B(n20262), .ZN(
        P1_U2833) );
  NOR2_X1 U23230 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20275), .ZN(n20265) );
  AOI22_X1 U23231 ( .A1(n20303), .A2(n20319), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n20265), .ZN(n20266) );
  OAI21_X1 U23232 ( .B1(n20323), .B2(n20289), .A(n20266), .ZN(n20267) );
  AOI211_X1 U23233 ( .C1(n20306), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20288), .B(n20267), .ZN(n20271) );
  AOI22_X1 U23234 ( .A1(n20269), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n20268), 
        .B2(n20321), .ZN(n20270) );
  OAI211_X1 U23235 ( .C1(n20272), .C2(n20292), .A(n20271), .B(n20270), .ZN(
        P1_U2834) );
  OAI22_X1 U23236 ( .A1(n20275), .A2(P1_REIP_REG_5__SCAN_IN), .B1(n20274), 
        .B2(n20273), .ZN(n20279) );
  INV_X1 U23237 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20830) );
  AOI22_X1 U23238 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20306), .B1(
        P1_EBX_REG_5__SCAN_IN), .B2(n20304), .ZN(n20277) );
  OAI211_X1 U23239 ( .C1(n20291), .C2(n20830), .A(n20277), .B(n20276), .ZN(
        n20278) );
  AOI211_X1 U23240 ( .C1(n20280), .C2(n20314), .A(n20279), .B(n20278), .ZN(
        n20281) );
  OAI21_X1 U23241 ( .B1(n20282), .B2(n20292), .A(n20281), .ZN(P1_U2835) );
  INV_X1 U23242 ( .A(n20283), .ZN(n20285) );
  OAI22_X1 U23243 ( .A1(n20286), .A2(n20285), .B1(n20284), .B2(n20312), .ZN(
        n20287) );
  AOI211_X1 U23244 ( .C1(n20306), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20288), .B(n20287), .ZN(n20300) );
  OAI22_X1 U23245 ( .A1(n20291), .A2(n20827), .B1(n20290), .B2(n20289), .ZN(
        n20297) );
  OAI22_X1 U23246 ( .A1(n20295), .A2(n20294), .B1(n20293), .B2(n20292), .ZN(
        n20296) );
  AOI211_X1 U23247 ( .C1(n20303), .C2(n20298), .A(n20297), .B(n20296), .ZN(
        n20299) );
  NAND2_X1 U23248 ( .A1(n20300), .A2(n20299), .ZN(P1_U2836) );
  AOI21_X1 U23249 ( .B1(n20309), .B2(n20898), .A(n20301), .ZN(n20318) );
  AOI22_X1 U23250 ( .A1(P1_EBX_REG_2__SCAN_IN), .A2(n20304), .B1(n20303), .B2(
        n20302), .ZN(n20317) );
  INV_X1 U23251 ( .A(n20305), .ZN(n20308) );
  AOI22_X1 U23252 ( .A1(n20308), .A2(n20307), .B1(n20306), .B2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20311) );
  NAND3_X1 U23253 ( .A1(n20309), .A2(P1_REIP_REG_1__SCAN_IN), .A3(n20824), 
        .ZN(n20310) );
  OAI211_X1 U23254 ( .C1(n13496), .C2(n20312), .A(n20311), .B(n20310), .ZN(
        n20313) );
  AOI21_X1 U23255 ( .B1(n20315), .B2(n20314), .A(n20313), .ZN(n20316) );
  OAI211_X1 U23256 ( .C1(n20318), .C2(n20824), .A(n20317), .B(n20316), .ZN(
        P1_U2838) );
  AOI22_X1 U23257 ( .A1(n20321), .A2(n11783), .B1(n20320), .B2(n20319), .ZN(
        n20322) );
  OAI21_X1 U23258 ( .B1(n20324), .B2(n20323), .A(n20322), .ZN(P1_U2866) );
  AOI22_X1 U23259 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20328), .B1(n20340), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20325) );
  OAI21_X1 U23260 ( .B1(n20327), .B2(n20326), .A(n20325), .ZN(P1_U2921) );
  INV_X1 U23261 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20330) );
  AOI22_X1 U23262 ( .A1(n20907), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20329) );
  OAI21_X1 U23263 ( .B1(n20330), .B2(n20356), .A(n20329), .ZN(P1_U2922) );
  INV_X1 U23264 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20332) );
  AOI22_X1 U23265 ( .A1(n20907), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20331) );
  OAI21_X1 U23266 ( .B1(n20332), .B2(n20356), .A(n20331), .ZN(P1_U2923) );
  AOI22_X1 U23267 ( .A1(n20907), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20333) );
  OAI21_X1 U23268 ( .B1(n14488), .B2(n20356), .A(n20333), .ZN(P1_U2924) );
  INV_X1 U23269 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20335) );
  AOI22_X1 U23270 ( .A1(n20907), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20334) );
  OAI21_X1 U23271 ( .B1(n20335), .B2(n20356), .A(n20334), .ZN(P1_U2925) );
  INV_X1 U23272 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20337) );
  AOI22_X1 U23273 ( .A1(n20907), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20336) );
  OAI21_X1 U23274 ( .B1(n20337), .B2(n20356), .A(n20336), .ZN(P1_U2926) );
  INV_X1 U23275 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20339) );
  AOI22_X1 U23276 ( .A1(n20907), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20338) );
  OAI21_X1 U23277 ( .B1(n20339), .B2(n20356), .A(n20338), .ZN(P1_U2927) );
  AOI22_X1 U23278 ( .A1(n20907), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20341) );
  OAI21_X1 U23279 ( .B1(n20342), .B2(n20356), .A(n20341), .ZN(P1_U2928) );
  AOI22_X1 U23280 ( .A1(n20907), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20343) );
  OAI21_X1 U23281 ( .B1(n20344), .B2(n20356), .A(n20343), .ZN(P1_U2929) );
  AOI22_X1 U23282 ( .A1(n20907), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20345) );
  OAI21_X1 U23283 ( .B1(n14138), .B2(n20356), .A(n20345), .ZN(P1_U2930) );
  AOI22_X1 U23284 ( .A1(n20907), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20346) );
  OAI21_X1 U23285 ( .B1(n11259), .B2(n20356), .A(n20346), .ZN(P1_U2931) );
  AOI22_X1 U23286 ( .A1(n20907), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20347) );
  OAI21_X1 U23287 ( .B1(n20348), .B2(n20356), .A(n20347), .ZN(P1_U2932) );
  AOI22_X1 U23288 ( .A1(n20907), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20349) );
  OAI21_X1 U23289 ( .B1(n20350), .B2(n20356), .A(n20349), .ZN(P1_U2933) );
  AOI22_X1 U23290 ( .A1(n20907), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20351) );
  OAI21_X1 U23291 ( .B1(n20352), .B2(n20356), .A(n20351), .ZN(P1_U2934) );
  AOI22_X1 U23292 ( .A1(n20907), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20353) );
  OAI21_X1 U23293 ( .B1(n20354), .B2(n20356), .A(n20353), .ZN(P1_U2935) );
  AOI22_X1 U23294 ( .A1(n20907), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20340), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20355) );
  OAI21_X1 U23295 ( .B1(n20357), .B2(n20356), .A(n20355), .ZN(P1_U2936) );
  AOI22_X1 U23296 ( .A1(n20369), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20368), .ZN(n20359) );
  NAND2_X1 U23297 ( .A1(n20359), .A2(n20358), .ZN(P1_U2961) );
  AOI22_X1 U23298 ( .A1(n20369), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20368), .ZN(n20361) );
  NAND2_X1 U23299 ( .A1(n20361), .A2(n20360), .ZN(P1_U2962) );
  AOI22_X1 U23300 ( .A1(n20369), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20368), .ZN(n20363) );
  NAND2_X1 U23301 ( .A1(n20363), .A2(n20362), .ZN(P1_U2963) );
  AOI22_X1 U23302 ( .A1(n20369), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20368), .ZN(n20365) );
  NAND2_X1 U23303 ( .A1(n20365), .A2(n20364), .ZN(P1_U2964) );
  AOI22_X1 U23304 ( .A1(n20369), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20368), .ZN(n20367) );
  NAND2_X1 U23305 ( .A1(n20367), .A2(n20366), .ZN(P1_U2965) );
  AOI22_X1 U23306 ( .A1(n20369), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20368), .ZN(n20371) );
  NAND2_X1 U23307 ( .A1(n20371), .A2(n20370), .ZN(P1_U2966) );
  NOR2_X1 U23308 ( .A1(n11733), .A2(n20372), .ZN(P1_U3032) );
  AOI22_X1 U23309 ( .A1(n20798), .A2(n20373), .B1(n20392), .B2(n20745), .ZN(
        n20375) );
  AOI22_X1 U23310 ( .A1(n20393), .A2(n20744), .B1(n20751), .B2(n20409), .ZN(
        n20374) );
  OAI211_X1 U23311 ( .C1(n20397), .C2(n20376), .A(n20375), .B(n20374), .ZN(
        P1_U3033) );
  AOI22_X1 U23312 ( .A1(n20798), .A2(n20757), .B1(n20756), .B2(n20392), .ZN(
        n20378) );
  AOI22_X1 U23313 ( .A1(n20393), .A2(n20755), .B1(n20409), .B2(n20711), .ZN(
        n20377) );
  OAI211_X1 U23314 ( .C1(n20397), .C2(n20379), .A(n20378), .B(n20377), .ZN(
        P1_U3034) );
  AOI22_X1 U23315 ( .A1(n20798), .A2(n20497), .B1(n20762), .B2(n20392), .ZN(
        n20381) );
  AOI22_X1 U23316 ( .A1(n20393), .A2(n20761), .B1(n20409), .B2(n20763), .ZN(
        n20380) );
  OAI211_X1 U23317 ( .C1(n20397), .C2(n20382), .A(n20381), .B(n20380), .ZN(
        P1_U3035) );
  INV_X1 U23318 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20385) );
  AOI22_X1 U23319 ( .A1(n20798), .A2(n20769), .B1(n20392), .B2(n20768), .ZN(
        n20384) );
  AOI22_X1 U23320 ( .A1(n20393), .A2(n20767), .B1(n20717), .B2(n20409), .ZN(
        n20383) );
  OAI211_X1 U23321 ( .C1(n20397), .C2(n20385), .A(n20384), .B(n20383), .ZN(
        P1_U3036) );
  AOI22_X1 U23322 ( .A1(n20798), .A2(n20775), .B1(n20774), .B2(n20392), .ZN(
        n20387) );
  AOI22_X1 U23323 ( .A1(n20393), .A2(n20773), .B1(n20409), .B2(n20721), .ZN(
        n20386) );
  OAI211_X1 U23324 ( .C1(n20397), .C2(n20388), .A(n20387), .B(n20386), .ZN(
        P1_U3037) );
  AOI22_X1 U23325 ( .A1(n20798), .A2(n20787), .B1(n20392), .B2(n20786), .ZN(
        n20390) );
  AOI22_X1 U23326 ( .A1(n20393), .A2(n20785), .B1(n20727), .B2(n20409), .ZN(
        n20389) );
  OAI211_X1 U23327 ( .C1(n20397), .C2(n20391), .A(n20390), .B(n20389), .ZN(
        P1_U3039) );
  AOI22_X1 U23328 ( .A1(n20798), .A2(n20688), .B1(n20794), .B2(n20392), .ZN(
        n20395) );
  AOI22_X1 U23329 ( .A1(n20393), .A2(n20796), .B1(n20409), .B2(n20797), .ZN(
        n20394) );
  OAI211_X1 U23330 ( .C1(n20397), .C2(n20396), .A(n20395), .B(n20394), .ZN(
        P1_U3040) );
  INV_X1 U23331 ( .A(n20398), .ZN(n20408) );
  AOI22_X1 U23332 ( .A1(n20408), .A2(n20761), .B1(n20762), .B2(n20407), .ZN(
        n20400) );
  AOI22_X1 U23333 ( .A1(n20410), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n20497), .B2(n20409), .ZN(n20399) );
  OAI211_X1 U23334 ( .C1(n20635), .C2(n20442), .A(n20400), .B(n20399), .ZN(
        P1_U3043) );
  AOI22_X1 U23335 ( .A1(n20408), .A2(n20767), .B1(n20768), .B2(n20407), .ZN(
        n20402) );
  AOI22_X1 U23336 ( .A1(n20410), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n20409), .B2(n20769), .ZN(n20401) );
  OAI211_X1 U23337 ( .C1(n20772), .C2(n20442), .A(n20402), .B(n20401), .ZN(
        P1_U3044) );
  AOI22_X1 U23338 ( .A1(n20408), .A2(n20779), .B1(n20780), .B2(n20407), .ZN(
        n20404) );
  AOI22_X1 U23339 ( .A1(n20410), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n20560), .B2(n20409), .ZN(n20403) );
  OAI211_X1 U23340 ( .C1(n20648), .C2(n20442), .A(n20404), .B(n20403), .ZN(
        P1_U3046) );
  AOI22_X1 U23341 ( .A1(n20408), .A2(n20785), .B1(n20786), .B2(n20407), .ZN(
        n20406) );
  AOI22_X1 U23342 ( .A1(n20410), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n20409), .B2(n20787), .ZN(n20405) );
  OAI211_X1 U23343 ( .C1(n20792), .C2(n20442), .A(n20406), .B(n20405), .ZN(
        P1_U3047) );
  AOI22_X1 U23344 ( .A1(n20408), .A2(n20796), .B1(n20794), .B2(n20407), .ZN(
        n20412) );
  AOI22_X1 U23345 ( .A1(n20410), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n20688), .B2(n20409), .ZN(n20411) );
  OAI211_X1 U23346 ( .C1(n20693), .C2(n20442), .A(n20412), .B(n20411), .ZN(
        P1_U3048) );
  NAND3_X1 U23347 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20661), .A3(
        n11729), .ZN(n20455) );
  OR2_X1 U23348 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20455), .ZN(
        n20441) );
  OAI22_X1 U23349 ( .A1(n20479), .A2(n20612), .B1(n20611), .B2(n20441), .ZN(
        n20414) );
  INV_X1 U23350 ( .A(n20414), .ZN(n20422) );
  AOI21_X1 U23351 ( .B1(n20442), .B2(n20479), .A(n21095), .ZN(n20415) );
  NOR2_X1 U23352 ( .A1(n20415), .A2(n20743), .ZN(n20417) );
  NAND2_X1 U23353 ( .A1(n20452), .A2(n20616), .ZN(n20419) );
  AOI22_X1 U23354 ( .A1(n20417), .A2(n20419), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20441), .ZN(n20416) );
  OAI21_X1 U23355 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20574), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20514) );
  NAND3_X1 U23356 ( .A1(n20619), .A2(n20416), .A3(n20514), .ZN(n20445) );
  INV_X1 U23357 ( .A(n20417), .ZN(n20420) );
  INV_X1 U23358 ( .A(n20574), .ZN(n20418) );
  NAND2_X1 U23359 ( .A1(n20418), .A2(n20661), .ZN(n20518) );
  AOI22_X1 U23360 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20445), .B1(
        n20744), .B2(n20444), .ZN(n20421) );
  OAI211_X1 U23361 ( .C1(n20754), .C2(n20442), .A(n20422), .B(n20421), .ZN(
        P1_U3049) );
  OAI22_X1 U23362 ( .A1(n20442), .A2(n20714), .B1(n20627), .B2(n20441), .ZN(
        n20423) );
  INV_X1 U23363 ( .A(n20423), .ZN(n20425) );
  AOI22_X1 U23364 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20445), .B1(
        n20755), .B2(n20444), .ZN(n20424) );
  OAI211_X1 U23365 ( .C1(n20760), .C2(n20479), .A(n20425), .B(n20424), .ZN(
        P1_U3050) );
  OAI22_X1 U23366 ( .A1(n20442), .A2(n20766), .B1(n20631), .B2(n20441), .ZN(
        n20426) );
  INV_X1 U23367 ( .A(n20426), .ZN(n20428) );
  AOI22_X1 U23368 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20445), .B1(
        n20761), .B2(n20444), .ZN(n20427) );
  OAI211_X1 U23369 ( .C1(n20635), .C2(n20479), .A(n20428), .B(n20427), .ZN(
        P1_U3051) );
  OAI22_X1 U23370 ( .A1(n20479), .A2(n20772), .B1(n20636), .B2(n20441), .ZN(
        n20429) );
  INV_X1 U23371 ( .A(n20429), .ZN(n20431) );
  AOI22_X1 U23372 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20445), .B1(
        n20767), .B2(n20444), .ZN(n20430) );
  OAI211_X1 U23373 ( .C1(n20720), .C2(n20442), .A(n20431), .B(n20430), .ZN(
        P1_U3052) );
  OAI22_X1 U23374 ( .A1(n20442), .A2(n20724), .B1(n20640), .B2(n20441), .ZN(
        n20432) );
  INV_X1 U23375 ( .A(n20432), .ZN(n20434) );
  AOI22_X1 U23376 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20445), .B1(
        n20773), .B2(n20444), .ZN(n20433) );
  OAI211_X1 U23377 ( .C1(n20778), .C2(n20479), .A(n20434), .B(n20433), .ZN(
        P1_U3053) );
  OAI22_X1 U23378 ( .A1(n20442), .A2(n20784), .B1(n20644), .B2(n20441), .ZN(
        n20435) );
  INV_X1 U23379 ( .A(n20435), .ZN(n20437) );
  AOI22_X1 U23380 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20445), .B1(
        n20779), .B2(n20444), .ZN(n20436) );
  OAI211_X1 U23381 ( .C1(n20648), .C2(n20479), .A(n20437), .B(n20436), .ZN(
        P1_U3054) );
  OAI22_X1 U23382 ( .A1(n20479), .A2(n20792), .B1(n20649), .B2(n20441), .ZN(
        n20438) );
  INV_X1 U23383 ( .A(n20438), .ZN(n20440) );
  AOI22_X1 U23384 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20445), .B1(
        n20785), .B2(n20444), .ZN(n20439) );
  OAI211_X1 U23385 ( .C1(n20730), .C2(n20442), .A(n20440), .B(n20439), .ZN(
        P1_U3055) );
  OAI22_X1 U23386 ( .A1(n20442), .A2(n20803), .B1(n20654), .B2(n20441), .ZN(
        n20443) );
  INV_X1 U23387 ( .A(n20443), .ZN(n20447) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20445), .B1(
        n20796), .B2(n20444), .ZN(n20446) );
  OAI211_X1 U23389 ( .C1(n20693), .C2(n20479), .A(n20447), .B(n20446), .ZN(
        P1_U3056) );
  OR2_X1 U23390 ( .A1(n20662), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20478) );
  OAI22_X1 U23391 ( .A1(n20495), .A2(n20612), .B1(n20611), .B2(n20478), .ZN(
        n20448) );
  INV_X1 U23392 ( .A(n20448), .ZN(n20459) );
  AOI21_X1 U23393 ( .B1(n20449), .B2(n20696), .A(n20666), .ZN(n20456) );
  AND2_X1 U23394 ( .A1(n20450), .A2(n11172), .ZN(n20738) );
  INV_X1 U23395 ( .A(n20478), .ZN(n20451) );
  AOI21_X1 U23396 ( .B1(n20452), .B2(n20738), .A(n20451), .ZN(n20457) );
  INV_X1 U23397 ( .A(n20457), .ZN(n20454) );
  NAND2_X1 U23398 ( .A1(n20743), .A2(n20455), .ZN(n20453) );
  OAI211_X1 U23399 ( .C1(n20456), .C2(n20454), .A(n20748), .B(n20453), .ZN(
        n20482) );
  OAI22_X1 U23400 ( .A1(n20457), .A2(n20456), .B1(n20806), .B2(n20455), .ZN(
        n20481) );
  AOI22_X1 U23401 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20482), .B1(
        n20744), .B2(n20481), .ZN(n20458) );
  OAI211_X1 U23402 ( .C1(n20754), .C2(n20479), .A(n20459), .B(n20458), .ZN(
        P1_U3057) );
  OAI22_X1 U23403 ( .A1(n20479), .A2(n20714), .B1(n20627), .B2(n20478), .ZN(
        n20460) );
  INV_X1 U23404 ( .A(n20460), .ZN(n20462) );
  AOI22_X1 U23405 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20482), .B1(
        n20755), .B2(n20481), .ZN(n20461) );
  OAI211_X1 U23406 ( .C1(n20760), .C2(n20495), .A(n20462), .B(n20461), .ZN(
        P1_U3058) );
  OAI22_X1 U23407 ( .A1(n20479), .A2(n20766), .B1(n20631), .B2(n20478), .ZN(
        n20463) );
  INV_X1 U23408 ( .A(n20463), .ZN(n20465) );
  AOI22_X1 U23409 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20482), .B1(
        n20761), .B2(n20481), .ZN(n20464) );
  OAI211_X1 U23410 ( .C1(n20635), .C2(n20495), .A(n20465), .B(n20464), .ZN(
        P1_U3059) );
  OAI22_X1 U23411 ( .A1(n20479), .A2(n20720), .B1(n20478), .B2(n20636), .ZN(
        n20466) );
  INV_X1 U23412 ( .A(n20466), .ZN(n20468) );
  AOI22_X1 U23413 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20482), .B1(
        n20767), .B2(n20481), .ZN(n20467) );
  OAI211_X1 U23414 ( .C1(n20772), .C2(n20495), .A(n20468), .B(n20467), .ZN(
        P1_U3060) );
  OAI22_X1 U23415 ( .A1(n20495), .A2(n20778), .B1(n20478), .B2(n20640), .ZN(
        n20469) );
  INV_X1 U23416 ( .A(n20469), .ZN(n20471) );
  AOI22_X1 U23417 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20482), .B1(
        n20773), .B2(n20481), .ZN(n20470) );
  OAI211_X1 U23418 ( .C1(n20724), .C2(n20479), .A(n20471), .B(n20470), .ZN(
        P1_U3061) );
  OAI22_X1 U23419 ( .A1(n20495), .A2(n20648), .B1(n20478), .B2(n20644), .ZN(
        n20472) );
  INV_X1 U23420 ( .A(n20472), .ZN(n20474) );
  AOI22_X1 U23421 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20482), .B1(
        n20779), .B2(n20481), .ZN(n20473) );
  OAI211_X1 U23422 ( .C1(n20784), .C2(n20479), .A(n20474), .B(n20473), .ZN(
        P1_U3062) );
  OAI22_X1 U23423 ( .A1(n20479), .A2(n20730), .B1(n20478), .B2(n20649), .ZN(
        n20475) );
  INV_X1 U23424 ( .A(n20475), .ZN(n20477) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20482), .B1(
        n20785), .B2(n20481), .ZN(n20476) );
  OAI211_X1 U23426 ( .C1(n20792), .C2(n20495), .A(n20477), .B(n20476), .ZN(
        P1_U3063) );
  OAI22_X1 U23427 ( .A1(n20479), .A2(n20803), .B1(n20654), .B2(n20478), .ZN(
        n20480) );
  INV_X1 U23428 ( .A(n20480), .ZN(n20484) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20482), .B1(
        n20796), .B2(n20481), .ZN(n20483) );
  OAI211_X1 U23430 ( .C1(n20693), .C2(n20495), .A(n20484), .B(n20483), .ZN(
        P1_U3064) );
  INV_X1 U23431 ( .A(n20485), .ZN(n20490) );
  AOI22_X1 U23432 ( .A1(n20745), .A2(n20491), .B1(n20744), .B2(n20490), .ZN(
        n20487) );
  AOI22_X1 U23433 ( .A1(n20492), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n20751), .B2(n20508), .ZN(n20486) );
  OAI211_X1 U23434 ( .C1(n20754), .C2(n20495), .A(n20487), .B(n20486), .ZN(
        P1_U3065) );
  AOI22_X1 U23435 ( .A1(n20768), .A2(n20491), .B1(n20767), .B2(n20490), .ZN(
        n20489) );
  AOI22_X1 U23436 ( .A1(n20492), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n20717), .B2(n20508), .ZN(n20488) );
  OAI211_X1 U23437 ( .C1(n20720), .C2(n20495), .A(n20489), .B(n20488), .ZN(
        P1_U3068) );
  AOI22_X1 U23438 ( .A1(n20786), .A2(n20491), .B1(n20785), .B2(n20490), .ZN(
        n20494) );
  AOI22_X1 U23439 ( .A1(n20492), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n20727), .B2(n20508), .ZN(n20493) );
  OAI211_X1 U23440 ( .C1(n20730), .C2(n20495), .A(n20494), .B(n20493), .ZN(
        P1_U3071) );
  INV_X1 U23441 ( .A(n20496), .ZN(n20507) );
  AOI22_X1 U23442 ( .A1(n20761), .A2(n20507), .B1(n20762), .B2(n20506), .ZN(
        n20499) );
  AOI22_X1 U23443 ( .A1(n20509), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n20497), .B2(n20508), .ZN(n20498) );
  OAI211_X1 U23444 ( .C1(n20635), .C2(n20531), .A(n20499), .B(n20498), .ZN(
        P1_U3075) );
  AOI22_X1 U23445 ( .A1(n20767), .A2(n20507), .B1(n20768), .B2(n20506), .ZN(
        n20501) );
  AOI22_X1 U23446 ( .A1(n20509), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n20508), .B2(n20769), .ZN(n20500) );
  OAI211_X1 U23447 ( .C1(n20772), .C2(n20531), .A(n20501), .B(n20500), .ZN(
        P1_U3076) );
  AOI22_X1 U23448 ( .A1(n20773), .A2(n20507), .B1(n20774), .B2(n20506), .ZN(
        n20503) );
  AOI22_X1 U23449 ( .A1(n20509), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n20775), .B2(n20508), .ZN(n20502) );
  OAI211_X1 U23450 ( .C1(n20778), .C2(n20531), .A(n20503), .B(n20502), .ZN(
        P1_U3077) );
  AOI22_X1 U23451 ( .A1(n20779), .A2(n20507), .B1(n20780), .B2(n20506), .ZN(
        n20505) );
  AOI22_X1 U23452 ( .A1(n20509), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n20560), .B2(n20508), .ZN(n20504) );
  OAI211_X1 U23453 ( .C1(n20648), .C2(n20531), .A(n20505), .B(n20504), .ZN(
        P1_U3078) );
  AOI22_X1 U23454 ( .A1(n20785), .A2(n20507), .B1(n20786), .B2(n20506), .ZN(
        n20511) );
  AOI22_X1 U23455 ( .A1(n20509), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n20508), .B2(n20787), .ZN(n20510) );
  OAI211_X1 U23456 ( .C1(n20792), .C2(n20531), .A(n20511), .B(n20510), .ZN(
        P1_U3079) );
  NOR2_X1 U23457 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20547), .ZN(
        n20536) );
  AOI22_X1 U23458 ( .A1(n20561), .A2(n20751), .B1(n20745), .B2(n20536), .ZN(
        n20522) );
  NAND2_X1 U23459 ( .A1(n20531), .A2(n20571), .ZN(n20512) );
  AOI21_X1 U23460 ( .B1(n20512), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20743), 
        .ZN(n20517) );
  NAND2_X1 U23461 ( .A1(n20543), .A2(n20616), .ZN(n20519) );
  INV_X1 U23462 ( .A(n20536), .ZN(n20513) );
  AOI22_X1 U23463 ( .A1(n20517), .A2(n20519), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20513), .ZN(n20515) );
  NAND3_X1 U23464 ( .A1(n20516), .A2(n20515), .A3(n20514), .ZN(n20539) );
  INV_X1 U23465 ( .A(n20517), .ZN(n20520) );
  AOI22_X1 U23466 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20539), .B1(
        n20744), .B2(n20538), .ZN(n20521) );
  OAI211_X1 U23467 ( .C1(n20754), .C2(n20531), .A(n20522), .B(n20521), .ZN(
        P1_U3081) );
  AOI22_X1 U23468 ( .A1(n20561), .A2(n20711), .B1(n20536), .B2(n20756), .ZN(
        n20524) );
  AOI22_X1 U23469 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20539), .B1(
        n20755), .B2(n20538), .ZN(n20523) );
  OAI211_X1 U23470 ( .C1(n20714), .C2(n20531), .A(n20524), .B(n20523), .ZN(
        P1_U3082) );
  AOI22_X1 U23471 ( .A1(n20561), .A2(n20763), .B1(n20536), .B2(n20762), .ZN(
        n20526) );
  AOI22_X1 U23472 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20539), .B1(
        n20761), .B2(n20538), .ZN(n20525) );
  OAI211_X1 U23473 ( .C1(n20766), .C2(n20531), .A(n20526), .B(n20525), .ZN(
        P1_U3083) );
  INV_X1 U23474 ( .A(n20531), .ZN(n20537) );
  AOI22_X1 U23475 ( .A1(n20537), .A2(n20769), .B1(n20536), .B2(n20768), .ZN(
        n20528) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20539), .B1(
        n20767), .B2(n20538), .ZN(n20527) );
  OAI211_X1 U23477 ( .C1(n20772), .C2(n20571), .A(n20528), .B(n20527), .ZN(
        P1_U3084) );
  AOI22_X1 U23478 ( .A1(n20561), .A2(n20721), .B1(n20536), .B2(n20774), .ZN(
        n20530) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20539), .B1(
        n20773), .B2(n20538), .ZN(n20529) );
  OAI211_X1 U23480 ( .C1(n20724), .C2(n20531), .A(n20530), .B(n20529), .ZN(
        P1_U3085) );
  AOI22_X1 U23481 ( .A1(n20537), .A2(n20560), .B1(n20780), .B2(n20536), .ZN(
        n20533) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20539), .B1(
        n20779), .B2(n20538), .ZN(n20532) );
  OAI211_X1 U23483 ( .C1(n20648), .C2(n20571), .A(n20533), .B(n20532), .ZN(
        P1_U3086) );
  AOI22_X1 U23484 ( .A1(n20537), .A2(n20787), .B1(n20536), .B2(n20786), .ZN(
        n20535) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20539), .B1(
        n20785), .B2(n20538), .ZN(n20534) );
  OAI211_X1 U23486 ( .C1(n20792), .C2(n20571), .A(n20535), .B(n20534), .ZN(
        P1_U3087) );
  AOI22_X1 U23487 ( .A1(n20537), .A2(n20688), .B1(n20794), .B2(n20536), .ZN(
        n20541) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20539), .B1(
        n20796), .B2(n20538), .ZN(n20540) );
  OAI211_X1 U23489 ( .C1(n20693), .C2(n20571), .A(n20541), .B(n20540), .ZN(
        P1_U3088) );
  INV_X1 U23490 ( .A(n20542), .ZN(n20566) );
  AOI21_X1 U23491 ( .B1(n20543), .B2(n20738), .A(n20566), .ZN(n20544) );
  OAI22_X1 U23492 ( .A1(n20544), .A2(n20743), .B1(n20547), .B2(n20806), .ZN(
        n20567) );
  AOI22_X1 U23493 ( .A1(n20745), .A2(n20566), .B1(n20744), .B2(n20567), .ZN(
        n20551) );
  AOI21_X1 U23494 ( .B1(n20547), .B2(n20546), .A(n20545), .ZN(n20548) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20568), .B1(
        n20576), .B2(n20751), .ZN(n20550) );
  OAI211_X1 U23496 ( .C1(n20754), .C2(n20571), .A(n20551), .B(n20550), .ZN(
        P1_U3089) );
  AOI22_X1 U23497 ( .A1(n20756), .A2(n20566), .B1(n20755), .B2(n20567), .ZN(
        n20553) );
  AOI22_X1 U23498 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20568), .B1(
        n20561), .B2(n20757), .ZN(n20552) );
  OAI211_X1 U23499 ( .C1(n20760), .C2(n20599), .A(n20553), .B(n20552), .ZN(
        P1_U3090) );
  AOI22_X1 U23500 ( .A1(n20762), .A2(n20566), .B1(n20761), .B2(n20567), .ZN(
        n20555) );
  AOI22_X1 U23501 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20568), .B1(
        n20576), .B2(n20763), .ZN(n20554) );
  OAI211_X1 U23502 ( .C1(n20766), .C2(n20571), .A(n20555), .B(n20554), .ZN(
        P1_U3091) );
  AOI22_X1 U23503 ( .A1(n20768), .A2(n20566), .B1(n20767), .B2(n20567), .ZN(
        n20557) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20568), .B1(
        n20576), .B2(n20717), .ZN(n20556) );
  OAI211_X1 U23505 ( .C1(n20720), .C2(n20571), .A(n20557), .B(n20556), .ZN(
        P1_U3092) );
  AOI22_X1 U23506 ( .A1(n20774), .A2(n20566), .B1(n20773), .B2(n20567), .ZN(
        n20559) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20568), .B1(
        n20576), .B2(n20721), .ZN(n20558) );
  OAI211_X1 U23508 ( .C1(n20724), .C2(n20571), .A(n20559), .B(n20558), .ZN(
        P1_U3093) );
  AOI22_X1 U23509 ( .A1(n20780), .A2(n20566), .B1(n20779), .B2(n20567), .ZN(
        n20563) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20568), .B1(
        n20561), .B2(n20560), .ZN(n20562) );
  OAI211_X1 U23511 ( .C1(n20648), .C2(n20599), .A(n20563), .B(n20562), .ZN(
        P1_U3094) );
  AOI22_X1 U23512 ( .A1(n20786), .A2(n20566), .B1(n20785), .B2(n20567), .ZN(
        n20565) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20568), .B1(
        n20576), .B2(n20727), .ZN(n20564) );
  OAI211_X1 U23514 ( .C1(n20730), .C2(n20571), .A(n20565), .B(n20564), .ZN(
        P1_U3095) );
  AOI22_X1 U23515 ( .A1(n20796), .A2(n20567), .B1(n20794), .B2(n20566), .ZN(
        n20570) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20568), .B1(
        n20576), .B2(n20797), .ZN(n20569) );
  OAI211_X1 U23517 ( .C1(n20803), .C2(n20571), .A(n20570), .B(n20569), .ZN(
        P1_U3096) );
  NOR2_X1 U23518 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20572), .ZN(
        n20594) );
  AOI21_X1 U23519 ( .B1(n20663), .B2(n20698), .A(n20594), .ZN(n20577) );
  INV_X1 U23520 ( .A(n20573), .ZN(n20575) );
  NAND2_X1 U23521 ( .A1(n20575), .A2(n20574), .ZN(n20705) );
  OAI22_X1 U23522 ( .A1(n20577), .A2(n20743), .B1(n20621), .B2(n20705), .ZN(
        n20595) );
  AOI22_X1 U23523 ( .A1(n20745), .A2(n20594), .B1(n20744), .B2(n20595), .ZN(
        n20581) );
  OAI21_X1 U23524 ( .B1(n20606), .B2(n20576), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20578) );
  NAND2_X1 U23525 ( .A1(n20578), .A2(n20577), .ZN(n20579) );
  AOI22_X1 U23526 ( .A1(n20596), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n20751), .B2(n20606), .ZN(n20580) );
  OAI211_X1 U23527 ( .C1(n20754), .C2(n20599), .A(n20581), .B(n20580), .ZN(
        P1_U3097) );
  AOI22_X1 U23528 ( .A1(n20756), .A2(n20594), .B1(n20755), .B2(n20595), .ZN(
        n20583) );
  AOI22_X1 U23529 ( .A1(n20596), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n20606), .B2(n20711), .ZN(n20582) );
  OAI211_X1 U23530 ( .C1(n20714), .C2(n20599), .A(n20583), .B(n20582), .ZN(
        P1_U3098) );
  AOI22_X1 U23531 ( .A1(n20762), .A2(n20594), .B1(n20761), .B2(n20595), .ZN(
        n20585) );
  AOI22_X1 U23532 ( .A1(n20596), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n20606), .B2(n20763), .ZN(n20584) );
  OAI211_X1 U23533 ( .C1(n20766), .C2(n20599), .A(n20585), .B(n20584), .ZN(
        P1_U3099) );
  AOI22_X1 U23534 ( .A1(n20768), .A2(n20594), .B1(n20767), .B2(n20595), .ZN(
        n20587) );
  AOI22_X1 U23535 ( .A1(n20596), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n20717), .B2(n20606), .ZN(n20586) );
  OAI211_X1 U23536 ( .C1(n20720), .C2(n20599), .A(n20587), .B(n20586), .ZN(
        P1_U3100) );
  AOI22_X1 U23537 ( .A1(n20774), .A2(n20594), .B1(n20773), .B2(n20595), .ZN(
        n20589) );
  AOI22_X1 U23538 ( .A1(n20596), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n20606), .B2(n20721), .ZN(n20588) );
  OAI211_X1 U23539 ( .C1(n20724), .C2(n20599), .A(n20589), .B(n20588), .ZN(
        P1_U3101) );
  AOI22_X1 U23540 ( .A1(n20780), .A2(n20594), .B1(n20779), .B2(n20595), .ZN(
        n20591) );
  AOI22_X1 U23541 ( .A1(n20596), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n20606), .B2(n20781), .ZN(n20590) );
  OAI211_X1 U23542 ( .C1(n20784), .C2(n20599), .A(n20591), .B(n20590), .ZN(
        P1_U3102) );
  AOI22_X1 U23543 ( .A1(n20786), .A2(n20594), .B1(n20785), .B2(n20595), .ZN(
        n20593) );
  AOI22_X1 U23544 ( .A1(n20596), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n20727), .B2(n20606), .ZN(n20592) );
  OAI211_X1 U23545 ( .C1(n20730), .C2(n20599), .A(n20593), .B(n20592), .ZN(
        P1_U3103) );
  AOI22_X1 U23546 ( .A1(n20796), .A2(n20595), .B1(n20794), .B2(n20594), .ZN(
        n20598) );
  AOI22_X1 U23547 ( .A1(n20596), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n20606), .B2(n20797), .ZN(n20597) );
  OAI211_X1 U23548 ( .C1(n20803), .C2(n20599), .A(n20598), .B(n20597), .ZN(
        P1_U3104) );
  AOI22_X1 U23549 ( .A1(n20756), .A2(n20605), .B1(n20755), .B2(n20604), .ZN(
        n20601) );
  AOI22_X1 U23550 ( .A1(n20607), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n20757), .B2(n20606), .ZN(n20600) );
  OAI211_X1 U23551 ( .C1(n20760), .C2(n20655), .A(n20601), .B(n20600), .ZN(
        P1_U3106) );
  AOI22_X1 U23552 ( .A1(n20774), .A2(n20605), .B1(n20773), .B2(n20604), .ZN(
        n20603) );
  AOI22_X1 U23553 ( .A1(n20607), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n20775), .B2(n20606), .ZN(n20602) );
  OAI211_X1 U23554 ( .C1(n20778), .C2(n20655), .A(n20603), .B(n20602), .ZN(
        P1_U3109) );
  AOI22_X1 U23555 ( .A1(n20786), .A2(n20605), .B1(n20785), .B2(n20604), .ZN(
        n20609) );
  AOI22_X1 U23556 ( .A1(n20607), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n20606), .B2(n20787), .ZN(n20608) );
  OAI211_X1 U23557 ( .C1(n20792), .C2(n20655), .A(n20609), .B(n20608), .ZN(
        P1_U3111) );
  NAND3_X1 U23558 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n11729), .ZN(n20664) );
  OR2_X1 U23559 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20664), .ZN(
        n20653) );
  OAI22_X1 U23560 ( .A1(n20684), .A2(n20612), .B1(n20611), .B2(n20653), .ZN(
        n20613) );
  INV_X1 U23561 ( .A(n20613), .ZN(n20626) );
  NAND3_X1 U23562 ( .A1(n20655), .A2(n20684), .A3(n20696), .ZN(n20615) );
  NAND2_X1 U23563 ( .A1(n20615), .A2(n20614), .ZN(n20620) );
  NAND2_X1 U23564 ( .A1(n20663), .A2(n20616), .ZN(n20623) );
  AOI22_X1 U23565 ( .A1(n20620), .A2(n20623), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20653), .ZN(n20618) );
  NAND3_X1 U23566 ( .A1(n20619), .A2(n20618), .A3(n20617), .ZN(n20658) );
  INV_X1 U23567 ( .A(n20620), .ZN(n20624) );
  AOI22_X1 U23568 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20658), .B1(
        n20744), .B2(n20657), .ZN(n20625) );
  OAI211_X1 U23569 ( .C1(n20754), .C2(n20655), .A(n20626), .B(n20625), .ZN(
        P1_U3113) );
  OAI22_X1 U23570 ( .A1(n20655), .A2(n20714), .B1(n20627), .B2(n20653), .ZN(
        n20628) );
  INV_X1 U23571 ( .A(n20628), .ZN(n20630) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20658), .B1(
        n20755), .B2(n20657), .ZN(n20629) );
  OAI211_X1 U23573 ( .C1(n20760), .C2(n20684), .A(n20630), .B(n20629), .ZN(
        P1_U3114) );
  OAI22_X1 U23574 ( .A1(n20655), .A2(n20766), .B1(n20631), .B2(n20653), .ZN(
        n20632) );
  INV_X1 U23575 ( .A(n20632), .ZN(n20634) );
  AOI22_X1 U23576 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20658), .B1(
        n20761), .B2(n20657), .ZN(n20633) );
  OAI211_X1 U23577 ( .C1(n20635), .C2(n20684), .A(n20634), .B(n20633), .ZN(
        P1_U3115) );
  OAI22_X1 U23578 ( .A1(n20684), .A2(n20772), .B1(n20636), .B2(n20653), .ZN(
        n20637) );
  INV_X1 U23579 ( .A(n20637), .ZN(n20639) );
  AOI22_X1 U23580 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20658), .B1(
        n20767), .B2(n20657), .ZN(n20638) );
  OAI211_X1 U23581 ( .C1(n20720), .C2(n20655), .A(n20639), .B(n20638), .ZN(
        P1_U3116) );
  OAI22_X1 U23582 ( .A1(n20684), .A2(n20778), .B1(n20653), .B2(n20640), .ZN(
        n20641) );
  INV_X1 U23583 ( .A(n20641), .ZN(n20643) );
  AOI22_X1 U23584 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20658), .B1(
        n20773), .B2(n20657), .ZN(n20642) );
  OAI211_X1 U23585 ( .C1(n20724), .C2(n20655), .A(n20643), .B(n20642), .ZN(
        P1_U3117) );
  OAI22_X1 U23586 ( .A1(n20655), .A2(n20784), .B1(n20644), .B2(n20653), .ZN(
        n20645) );
  INV_X1 U23587 ( .A(n20645), .ZN(n20647) );
  AOI22_X1 U23588 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20658), .B1(
        n20779), .B2(n20657), .ZN(n20646) );
  OAI211_X1 U23589 ( .C1(n20648), .C2(n20684), .A(n20647), .B(n20646), .ZN(
        P1_U3118) );
  OAI22_X1 U23590 ( .A1(n20655), .A2(n20730), .B1(n20653), .B2(n20649), .ZN(
        n20650) );
  INV_X1 U23591 ( .A(n20650), .ZN(n20652) );
  AOI22_X1 U23592 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20658), .B1(
        n20785), .B2(n20657), .ZN(n20651) );
  OAI211_X1 U23593 ( .C1(n20792), .C2(n20684), .A(n20652), .B(n20651), .ZN(
        P1_U3119) );
  OAI22_X1 U23594 ( .A1(n20655), .A2(n20803), .B1(n20654), .B2(n20653), .ZN(
        n20656) );
  INV_X1 U23595 ( .A(n20656), .ZN(n20660) );
  AOI22_X1 U23596 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20658), .B1(
        n20796), .B2(n20657), .ZN(n20659) );
  OAI211_X1 U23597 ( .C1(n20693), .C2(n20684), .A(n20660), .B(n20659), .ZN(
        P1_U3120) );
  AOI21_X1 U23598 ( .B1(n20663), .B2(n20738), .A(n10179), .ZN(n20665) );
  OAI22_X1 U23599 ( .A1(n20665), .A2(n20743), .B1(n20664), .B2(n20806), .ZN(
        n20687) );
  AOI22_X1 U23600 ( .A1(n20745), .A2(n10179), .B1(n20744), .B2(n20687), .ZN(
        n20673) );
  INV_X1 U23601 ( .A(n20664), .ZN(n20669) );
  NOR2_X1 U23602 ( .A1(n20671), .A2(n20743), .ZN(n20667) );
  OAI21_X1 U23603 ( .B1(n20667), .B2(n20666), .A(n20665), .ZN(n20668) );
  OAI211_X1 U23604 ( .C1(n20696), .C2(n20669), .A(n20748), .B(n20668), .ZN(
        n20690) );
  AOI22_X1 U23605 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20690), .B1(
        n20695), .B2(n20751), .ZN(n20672) );
  OAI211_X1 U23606 ( .C1(n20754), .C2(n20684), .A(n20673), .B(n20672), .ZN(
        P1_U3121) );
  AOI22_X1 U23607 ( .A1(n20756), .A2(n10179), .B1(n20755), .B2(n20687), .ZN(
        n20675) );
  INV_X1 U23608 ( .A(n20684), .ZN(n20689) );
  AOI22_X1 U23609 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20690), .B1(
        n20689), .B2(n20757), .ZN(n20674) );
  OAI211_X1 U23610 ( .C1(n20760), .C2(n20737), .A(n20675), .B(n20674), .ZN(
        P1_U3122) );
  AOI22_X1 U23611 ( .A1(n20762), .A2(n10179), .B1(n20761), .B2(n20687), .ZN(
        n20677) );
  AOI22_X1 U23612 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20690), .B1(
        n20695), .B2(n20763), .ZN(n20676) );
  OAI211_X1 U23613 ( .C1(n20766), .C2(n20684), .A(n20677), .B(n20676), .ZN(
        P1_U3123) );
  AOI22_X1 U23614 ( .A1(n20768), .A2(n10179), .B1(n20767), .B2(n20687), .ZN(
        n20679) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20690), .B1(
        n20695), .B2(n20717), .ZN(n20678) );
  OAI211_X1 U23616 ( .C1(n20720), .C2(n20684), .A(n20679), .B(n20678), .ZN(
        P1_U3124) );
  AOI22_X1 U23617 ( .A1(n20774), .A2(n10179), .B1(n20773), .B2(n20687), .ZN(
        n20681) );
  AOI22_X1 U23618 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20690), .B1(
        n20695), .B2(n20721), .ZN(n20680) );
  OAI211_X1 U23619 ( .C1(n20724), .C2(n20684), .A(n20681), .B(n20680), .ZN(
        P1_U3125) );
  AOI22_X1 U23620 ( .A1(n20780), .A2(n10179), .B1(n20779), .B2(n20687), .ZN(
        n20683) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20690), .B1(
        n20695), .B2(n20781), .ZN(n20682) );
  OAI211_X1 U23622 ( .C1(n20784), .C2(n20684), .A(n20683), .B(n20682), .ZN(
        P1_U3126) );
  AOI22_X1 U23623 ( .A1(n20786), .A2(n10179), .B1(n20785), .B2(n20687), .ZN(
        n20686) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20690), .B1(
        n20689), .B2(n20787), .ZN(n20685) );
  OAI211_X1 U23625 ( .C1(n20792), .C2(n20737), .A(n20686), .B(n20685), .ZN(
        P1_U3127) );
  AOI22_X1 U23626 ( .A1(n20796), .A2(n20687), .B1(n20794), .B2(n10179), .ZN(
        n20692) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20690), .B1(
        n20689), .B2(n20688), .ZN(n20691) );
  OAI211_X1 U23628 ( .C1(n20693), .C2(n20737), .A(n20692), .B(n20691), .ZN(
        P1_U3128) );
  NOR2_X1 U23629 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20694), .ZN(
        n20731) );
  AOI22_X1 U23630 ( .A1(n20732), .A2(n20751), .B1(n20745), .B2(n20731), .ZN(
        n20710) );
  OAI21_X1 U23631 ( .B1(n20695), .B2(n20732), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20697) );
  NAND2_X1 U23632 ( .A1(n20697), .A2(n20696), .ZN(n20708) );
  NAND2_X1 U23633 ( .A1(n20699), .A2(n20698), .ZN(n20707) );
  INV_X1 U23634 ( .A(n20707), .ZN(n20701) );
  OAI22_X1 U23635 ( .A1(n20708), .A2(n20701), .B1(n20731), .B2(n20700), .ZN(
        n20702) );
  AOI211_X1 U23636 ( .C1(n20705), .C2(P1_STATE2_REG_2__SCAN_IN), .A(n20703), 
        .B(n20702), .ZN(n20704) );
  AOI22_X1 U23637 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20734), .B1(
        n20744), .B2(n20733), .ZN(n20709) );
  OAI211_X1 U23638 ( .C1(n20754), .C2(n20737), .A(n20710), .B(n20709), .ZN(
        P1_U3129) );
  AOI22_X1 U23639 ( .A1(n20732), .A2(n20711), .B1(n20731), .B2(n20756), .ZN(
        n20713) );
  AOI22_X1 U23640 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20734), .B1(
        n20755), .B2(n20733), .ZN(n20712) );
  OAI211_X1 U23641 ( .C1(n20714), .C2(n20737), .A(n20713), .B(n20712), .ZN(
        P1_U3130) );
  AOI22_X1 U23642 ( .A1(n20732), .A2(n20763), .B1(n20731), .B2(n20762), .ZN(
        n20716) );
  AOI22_X1 U23643 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20734), .B1(
        n20761), .B2(n20733), .ZN(n20715) );
  OAI211_X1 U23644 ( .C1(n20766), .C2(n20737), .A(n20716), .B(n20715), .ZN(
        P1_U3131) );
  AOI22_X1 U23645 ( .A1(n20732), .A2(n20717), .B1(n20768), .B2(n20731), .ZN(
        n20719) );
  AOI22_X1 U23646 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20734), .B1(
        n20767), .B2(n20733), .ZN(n20718) );
  OAI211_X1 U23647 ( .C1(n20720), .C2(n20737), .A(n20719), .B(n20718), .ZN(
        P1_U3132) );
  AOI22_X1 U23648 ( .A1(n20732), .A2(n20721), .B1(n20731), .B2(n20774), .ZN(
        n20723) );
  AOI22_X1 U23649 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20734), .B1(
        n20773), .B2(n20733), .ZN(n20722) );
  OAI211_X1 U23650 ( .C1(n20724), .C2(n20737), .A(n20723), .B(n20722), .ZN(
        P1_U3133) );
  AOI22_X1 U23651 ( .A1(n20732), .A2(n20781), .B1(n20731), .B2(n20780), .ZN(
        n20726) );
  AOI22_X1 U23652 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20734), .B1(
        n20779), .B2(n20733), .ZN(n20725) );
  OAI211_X1 U23653 ( .C1(n20784), .C2(n20737), .A(n20726), .B(n20725), .ZN(
        P1_U3134) );
  AOI22_X1 U23654 ( .A1(n20732), .A2(n20727), .B1(n20786), .B2(n20731), .ZN(
        n20729) );
  AOI22_X1 U23655 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20734), .B1(
        n20785), .B2(n20733), .ZN(n20728) );
  OAI211_X1 U23656 ( .C1(n20730), .C2(n20737), .A(n20729), .B(n20728), .ZN(
        P1_U3135) );
  AOI22_X1 U23657 ( .A1(n20732), .A2(n20797), .B1(n20731), .B2(n20794), .ZN(
        n20736) );
  AOI22_X1 U23658 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20734), .B1(
        n20796), .B2(n20733), .ZN(n20735) );
  OAI211_X1 U23659 ( .C1(n20803), .C2(n20737), .A(n20736), .B(n20735), .ZN(
        P1_U3136) );
  INV_X1 U23660 ( .A(n20742), .ZN(n20793) );
  INV_X1 U23661 ( .A(n20738), .ZN(n20739) );
  OAI222_X1 U23662 ( .A1(n20743), .A2(n20742), .B1(n20806), .B2(n20741), .C1(
        n20740), .C2(n20739), .ZN(n20795) );
  AOI22_X1 U23663 ( .A1(n20745), .A2(n20793), .B1(n20795), .B2(n20744), .ZN(
        n20753) );
  AND2_X1 U23664 ( .A1(n20747), .A2(n20746), .ZN(n20750) );
  AOI22_X1 U23665 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20799), .B1(
        n20798), .B2(n20751), .ZN(n20752) );
  OAI211_X1 U23666 ( .C1(n20754), .C2(n20802), .A(n20753), .B(n20752), .ZN(
        P1_U3153) );
  AOI22_X1 U23667 ( .A1(n20756), .A2(n20793), .B1(n20795), .B2(n20755), .ZN(
        n20759) );
  AOI22_X1 U23668 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20799), .B1(
        n20788), .B2(n20757), .ZN(n20758) );
  OAI211_X1 U23669 ( .C1(n20760), .C2(n20791), .A(n20759), .B(n20758), .ZN(
        P1_U3154) );
  AOI22_X1 U23670 ( .A1(n20762), .A2(n20793), .B1(n20795), .B2(n20761), .ZN(
        n20765) );
  AOI22_X1 U23671 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20799), .B1(
        n20798), .B2(n20763), .ZN(n20764) );
  OAI211_X1 U23672 ( .C1(n20766), .C2(n20802), .A(n20765), .B(n20764), .ZN(
        P1_U3155) );
  AOI22_X1 U23673 ( .A1(n20768), .A2(n20793), .B1(n20795), .B2(n20767), .ZN(
        n20771) );
  AOI22_X1 U23674 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20799), .B1(
        n20788), .B2(n20769), .ZN(n20770) );
  OAI211_X1 U23675 ( .C1(n20772), .C2(n20791), .A(n20771), .B(n20770), .ZN(
        P1_U3156) );
  AOI22_X1 U23676 ( .A1(n20774), .A2(n20793), .B1(n20795), .B2(n20773), .ZN(
        n20777) );
  AOI22_X1 U23677 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20799), .B1(
        n20788), .B2(n20775), .ZN(n20776) );
  OAI211_X1 U23678 ( .C1(n20778), .C2(n20791), .A(n20777), .B(n20776), .ZN(
        P1_U3157) );
  AOI22_X1 U23679 ( .A1(n20780), .A2(n20793), .B1(n20795), .B2(n20779), .ZN(
        n20783) );
  AOI22_X1 U23680 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20799), .B1(
        n20798), .B2(n20781), .ZN(n20782) );
  OAI211_X1 U23681 ( .C1(n20784), .C2(n20802), .A(n20783), .B(n20782), .ZN(
        P1_U3158) );
  AOI22_X1 U23682 ( .A1(n20786), .A2(n20793), .B1(n20795), .B2(n20785), .ZN(
        n20790) );
  AOI22_X1 U23683 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20799), .B1(
        n20788), .B2(n20787), .ZN(n20789) );
  OAI211_X1 U23684 ( .C1(n20792), .C2(n20791), .A(n20790), .B(n20789), .ZN(
        P1_U3159) );
  AOI22_X1 U23685 ( .A1(n20796), .A2(n20795), .B1(n20794), .B2(n20793), .ZN(
        n20801) );
  AOI22_X1 U23686 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20799), .B1(
        n20798), .B2(n20797), .ZN(n20800) );
  OAI211_X1 U23687 ( .C1(n20803), .C2(n20802), .A(n20801), .B(n20800), .ZN(
        P1_U3160) );
  OAI211_X1 U23688 ( .C1(n20807), .C2(n20806), .A(n20805), .B(n20804), .ZN(
        P1_U3163) );
  INV_X1 U23689 ( .A(n20884), .ZN(n20880) );
  AND2_X1 U23690 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20880), .ZN(
        P1_U3164) );
  AND2_X1 U23691 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20880), .ZN(
        P1_U3165) );
  AND2_X1 U23692 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20880), .ZN(
        P1_U3166) );
  AND2_X1 U23693 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20880), .ZN(
        P1_U3167) );
  AND2_X1 U23694 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20880), .ZN(
        P1_U3168) );
  AND2_X1 U23695 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20880), .ZN(
        P1_U3169) );
  AND2_X1 U23696 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20880), .ZN(
        P1_U3170) );
  AND2_X1 U23697 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20880), .ZN(
        P1_U3171) );
  AND2_X1 U23698 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20880), .ZN(
        P1_U3172) );
  AND2_X1 U23699 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20880), .ZN(
        P1_U3173) );
  AND2_X1 U23700 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20880), .ZN(
        P1_U3174) );
  AND2_X1 U23701 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20880), .ZN(
        P1_U3175) );
  AND2_X1 U23702 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20880), .ZN(
        P1_U3176) );
  AND2_X1 U23703 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20880), .ZN(
        P1_U3177) );
  AND2_X1 U23704 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20880), .ZN(
        P1_U3178) );
  AND2_X1 U23705 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20880), .ZN(
        P1_U3179) );
  AND2_X1 U23706 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20880), .ZN(
        P1_U3180) );
  AND2_X1 U23707 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20880), .ZN(
        P1_U3181) );
  AND2_X1 U23708 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20880), .ZN(
        P1_U3182) );
  AND2_X1 U23709 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20880), .ZN(
        P1_U3183) );
  AND2_X1 U23710 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20880), .ZN(
        P1_U3184) );
  AND2_X1 U23711 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20880), .ZN(
        P1_U3185) );
  AND2_X1 U23712 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20880), .ZN(P1_U3186) );
  AND2_X1 U23713 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20880), .ZN(P1_U3187) );
  AND2_X1 U23714 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20880), .ZN(P1_U3188) );
  AND2_X1 U23715 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20880), .ZN(P1_U3189) );
  AND2_X1 U23716 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20880), .ZN(P1_U3190) );
  AND2_X1 U23717 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20880), .ZN(P1_U3191) );
  AND2_X1 U23718 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20880), .ZN(P1_U3192) );
  AND2_X1 U23719 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20880), .ZN(P1_U3193) );
  AND2_X1 U23720 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20808), .ZN(n20821) );
  OAI21_X1 U23721 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n21013), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20809) );
  AOI211_X1 U23722 ( .C1(HOLD), .C2(P1_STATE_REG_1__SCAN_IN), .A(n20810), .B(
        n20809), .ZN(n20811) );
  OAI22_X1 U23723 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20821), .B1(n20875), 
        .B2(n20811), .ZN(P1_U3194) );
  AND2_X1 U23724 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20813) );
  INV_X1 U23725 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20815) );
  NOR2_X1 U23726 ( .A1(n20814), .A2(n20815), .ZN(n20812) );
  OAI22_X1 U23727 ( .A1(n20813), .A2(n21013), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20812), .ZN(n20820) );
  NOR3_X1 U23728 ( .A1(NA), .A2(n20814), .A3(n20906), .ZN(n20816) );
  OAI22_X1 U23729 ( .A1(n20817), .A2(n20816), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20815), .ZN(n20818) );
  OAI22_X1 U23730 ( .A1(n20821), .A2(n20820), .B1(n20819), .B2(n20818), .ZN(
        P1_U3196) );
  INV_X1 U23731 ( .A(n20849), .ZN(n20870) );
  INV_X1 U23732 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20822) );
  NAND2_X1 U23733 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20875), .ZN(n20872) );
  OAI222_X1 U23734 ( .A1(n20870), .A2(n20824), .B1(n20822), .B2(n20875), .C1(
        n20898), .C2(n20868), .ZN(P1_U3197) );
  AOI22_X1 U23735 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20916), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n20849), .ZN(n20823) );
  OAI21_X1 U23736 ( .B1(n20824), .B2(n20868), .A(n20823), .ZN(P1_U3198) );
  INV_X1 U23737 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20826) );
  OAI222_X1 U23738 ( .A1(n20868), .A2(n20826), .B1(n20825), .B2(n20875), .C1(
        n20827), .C2(n20870), .ZN(P1_U3199) );
  INV_X1 U23739 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20828) );
  OAI222_X1 U23740 ( .A1(n20870), .A2(n20830), .B1(n20828), .B2(n20875), .C1(
        n20827), .C2(n20868), .ZN(P1_U3200) );
  AOI22_X1 U23741 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n20916), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n20849), .ZN(n20829) );
  OAI21_X1 U23742 ( .B1(n20830), .B2(n20868), .A(n20829), .ZN(P1_U3201) );
  INV_X1 U23743 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20832) );
  AOI22_X1 U23744 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20916), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20849), .ZN(n20831) );
  OAI21_X1 U23745 ( .B1(n20832), .B2(n20868), .A(n20831), .ZN(P1_U3202) );
  AOI22_X1 U23746 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20916), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20852), .ZN(n20833) );
  OAI21_X1 U23747 ( .B1(n20835), .B2(n20870), .A(n20833), .ZN(P1_U3203) );
  INV_X1 U23748 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20834) );
  OAI222_X1 U23749 ( .A1(n20872), .A2(n20835), .B1(n20834), .B2(n20875), .C1(
        n20837), .C2(n20870), .ZN(P1_U3204) );
  INV_X1 U23750 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20836) );
  OAI222_X1 U23751 ( .A1(n20872), .A2(n20837), .B1(n20836), .B2(n20875), .C1(
        n20840), .C2(n20870), .ZN(P1_U3205) );
  INV_X1 U23752 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20839) );
  OAI222_X1 U23753 ( .A1(n20868), .A2(n20840), .B1(n20839), .B2(n20875), .C1(
        n20838), .C2(n20870), .ZN(P1_U3206) );
  AOI222_X1 U23754 ( .A1(n20849), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20852), .ZN(n20841) );
  INV_X1 U23755 ( .A(n20841), .ZN(P1_U3207) );
  AOI222_X1 U23756 ( .A1(n20852), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20916), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20849), .ZN(n20842) );
  INV_X1 U23757 ( .A(n20842), .ZN(P1_U3208) );
  INV_X1 U23758 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20843) );
  OAI222_X1 U23759 ( .A1(n20868), .A2(n20844), .B1(n20843), .B2(n20875), .C1(
        n20845), .C2(n20870), .ZN(P1_U3209) );
  INV_X1 U23760 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20846) );
  OAI222_X1 U23761 ( .A1(n20870), .A2(n20848), .B1(n20846), .B2(n20875), .C1(
        n20845), .C2(n20868), .ZN(P1_U3210) );
  INV_X1 U23762 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20847) );
  OAI222_X1 U23763 ( .A1(n20868), .A2(n20848), .B1(n20847), .B2(n20875), .C1(
        n20851), .C2(n20870), .ZN(P1_U3211) );
  AOI22_X1 U23764 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20916), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20849), .ZN(n20850) );
  OAI21_X1 U23765 ( .B1(n20851), .B2(n20868), .A(n20850), .ZN(P1_U3212) );
  AOI22_X1 U23766 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20916), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20852), .ZN(n20853) );
  OAI21_X1 U23767 ( .B1(n20855), .B2(n20870), .A(n20853), .ZN(P1_U3213) );
  INV_X1 U23768 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20854) );
  OAI222_X1 U23769 ( .A1(n20868), .A2(n20855), .B1(n20854), .B2(n20875), .C1(
        n20857), .C2(n20870), .ZN(P1_U3214) );
  INV_X1 U23770 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n20856) );
  OAI222_X1 U23771 ( .A1(n20868), .A2(n20857), .B1(n20856), .B2(n20875), .C1(
        n21119), .C2(n20870), .ZN(P1_U3215) );
  INV_X1 U23772 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20858) );
  INV_X1 U23773 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21042) );
  OAI222_X1 U23774 ( .A1(n20872), .A2(n21119), .B1(n20858), .B2(n20875), .C1(
        n21042), .C2(n20870), .ZN(P1_U3216) );
  INV_X1 U23775 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20859) );
  OAI222_X1 U23776 ( .A1(n20872), .A2(n21042), .B1(n20859), .B2(n20875), .C1(
        n21098), .C2(n20870), .ZN(P1_U3217) );
  INV_X1 U23777 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20860) );
  OAI222_X1 U23778 ( .A1(n20872), .A2(n21098), .B1(n20860), .B2(n20875), .C1(
        n21058), .C2(n20870), .ZN(P1_U3218) );
  INV_X1 U23779 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20861) );
  INV_X1 U23780 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21026) );
  OAI222_X1 U23781 ( .A1(n20872), .A2(n21058), .B1(n20861), .B2(n20875), .C1(
        n21026), .C2(n20870), .ZN(P1_U3219) );
  INV_X1 U23782 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20990) );
  INV_X1 U23783 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20862) );
  OAI222_X1 U23784 ( .A1(n20870), .A2(n20990), .B1(n20862), .B2(n20875), .C1(
        n21026), .C2(n20868), .ZN(P1_U3220) );
  INV_X1 U23785 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20863) );
  INV_X1 U23786 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21007) );
  OAI222_X1 U23787 ( .A1(n20872), .A2(n20990), .B1(n20863), .B2(n20875), .C1(
        n21007), .C2(n20870), .ZN(P1_U3221) );
  INV_X1 U23788 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20864) );
  OAI222_X1 U23789 ( .A1(n20872), .A2(n21007), .B1(n20864), .B2(n20875), .C1(
        n20866), .C2(n20870), .ZN(P1_U3222) );
  INV_X1 U23790 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20865) );
  INV_X1 U23791 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21023) );
  OAI222_X1 U23792 ( .A1(n20868), .A2(n20866), .B1(n20865), .B2(n20875), .C1(
        n21023), .C2(n20870), .ZN(P1_U3223) );
  INV_X1 U23793 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20867) );
  OAI222_X1 U23794 ( .A1(n20868), .A2(n21023), .B1(n20867), .B2(n20875), .C1(
        n21040), .C2(n20870), .ZN(P1_U3224) );
  INV_X1 U23795 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n20959) );
  INV_X1 U23796 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20869) );
  OAI222_X1 U23797 ( .A1(n20870), .A2(n20959), .B1(n20869), .B2(n20875), .C1(
        n21040), .C2(n20868), .ZN(P1_U3225) );
  INV_X1 U23798 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20871) );
  OAI222_X1 U23799 ( .A1(n20872), .A2(n20959), .B1(n20871), .B2(n20875), .C1(
        n21032), .C2(n20870), .ZN(P1_U3226) );
  INV_X1 U23800 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20873) );
  AOI22_X1 U23801 ( .A1(n20875), .A2(n20969), .B1(n20873), .B2(n20916), .ZN(
        P1_U3458) );
  INV_X1 U23802 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21016) );
  INV_X1 U23803 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20874) );
  AOI22_X1 U23804 ( .A1(n20875), .A2(n21016), .B1(n20874), .B2(n20916), .ZN(
        P1_U3459) );
  INV_X1 U23805 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20876) );
  AOI22_X1 U23806 ( .A1(n20875), .A2(n20877), .B1(n20876), .B2(n20916), .ZN(
        P1_U3460) );
  INV_X1 U23807 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21027) );
  INV_X1 U23808 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20878) );
  AOI22_X1 U23809 ( .A1(n20875), .A2(n21027), .B1(n20878), .B2(n20916), .ZN(
        P1_U3461) );
  INV_X1 U23810 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20881) );
  INV_X1 U23811 ( .A(n20882), .ZN(n20879) );
  AOI21_X1 U23812 ( .B1(n20881), .B2(n20880), .A(n20879), .ZN(P1_U3464) );
  OAI21_X1 U23813 ( .B1(n20884), .B2(n20883), .A(n20882), .ZN(P1_U3465) );
  OAI22_X1 U23814 ( .A1(n20886), .A2(n20897), .B1(n20888), .B2(n20885), .ZN(
        n20887) );
  MUX2_X1 U23815 ( .A(n20887), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n20894), .Z(P1_U3469) );
  OAI22_X1 U23816 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20888), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13985), .ZN(n20889) );
  INV_X1 U23817 ( .A(n20889), .ZN(n20890) );
  OAI21_X1 U23818 ( .B1(n20891), .B2(n20897), .A(n20890), .ZN(n20893) );
  AOI22_X1 U23819 ( .A1(n20894), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20893), .B2(n20892), .ZN(n20895) );
  OAI21_X1 U23820 ( .B1(n20897), .B2(n20896), .A(n20895), .ZN(P1_U3474) );
  AOI21_X1 U23821 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20899) );
  AOI22_X1 U23822 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20899), .B2(n20898), .ZN(n20901) );
  AOI22_X1 U23823 ( .A1(n20903), .A2(n20901), .B1(n21016), .B2(n20900), .ZN(
        P1_U3481) );
  OAI21_X1 U23824 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20903), .ZN(n20902) );
  OAI21_X1 U23825 ( .B1(n20903), .B2(n21027), .A(n20902), .ZN(P1_U3482) );
  AOI22_X1 U23826 ( .A1(n20875), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20994), 
        .B2(n20916), .ZN(P1_U3483) );
  AOI211_X1 U23827 ( .C1(n20907), .C2(n20906), .A(n20905), .B(n20904), .ZN(
        n20915) );
  INV_X1 U23828 ( .A(n20908), .ZN(n20909) );
  OAI211_X1 U23829 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20910), .A(n20909), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20912) );
  AOI21_X1 U23830 ( .B1(n20912), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20911), 
        .ZN(n20914) );
  NAND2_X1 U23831 ( .A1(n20915), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20913) );
  OAI21_X1 U23832 ( .B1(n20915), .B2(n20914), .A(n20913), .ZN(P1_U3485) );
  AOI22_X1 U23833 ( .A1(n20875), .A2(n21011), .B1(n20967), .B2(n20916), .ZN(
        P1_U3486) );
  AOI22_X1 U23834 ( .A1(DATAI_19_), .A2(keyinput_f13), .B1(DATAI_26_), .B2(
        keyinput_f6), .ZN(n20917) );
  OAI221_X1 U23835 ( .B1(DATAI_19_), .B2(keyinput_f13), .C1(DATAI_26_), .C2(
        keyinput_f6), .A(n20917), .ZN(n20924) );
  AOI22_X1 U23836 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_f43), 
        .B1(DATAI_12_), .B2(keyinput_f20), .ZN(n20918) );
  OAI221_X1 U23837 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_f43), 
        .C1(DATAI_12_), .C2(keyinput_f20), .A(n20918), .ZN(n20923) );
  AOI22_X1 U23838 ( .A1(DATAI_9_), .A2(keyinput_f23), .B1(
        P1_REIP_REG_28__SCAN_IN), .B2(keyinput_f55), .ZN(n20919) );
  OAI221_X1 U23839 ( .B1(DATAI_9_), .B2(keyinput_f23), .C1(
        P1_REIP_REG_28__SCAN_IN), .C2(keyinput_f55), .A(n20919), .ZN(n20922)
         );
  AOI22_X1 U23840 ( .A1(DATAI_17_), .A2(keyinput_f15), .B1(
        P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_f44), .ZN(n20920) );
  OAI221_X1 U23841 ( .B1(DATAI_17_), .B2(keyinput_f15), .C1(
        P1_STATEBS16_REG_SCAN_IN), .C2(keyinput_f44), .A(n20920), .ZN(n20921)
         );
  NOR4_X1 U23842 ( .A1(n20924), .A2(n20923), .A3(n20922), .A4(n20921), .ZN(
        n20952) );
  XNOR2_X1 U23843 ( .A(P1_REIP_REG_21__SCAN_IN), .B(keyinput_f62), .ZN(n20932)
         );
  AOI22_X1 U23844 ( .A1(DATAI_27_), .A2(keyinput_f5), .B1(n20926), .B2(
        keyinput_f3), .ZN(n20925) );
  OAI221_X1 U23845 ( .B1(DATAI_27_), .B2(keyinput_f5), .C1(n20926), .C2(
        keyinput_f3), .A(n20925), .ZN(n20931) );
  AOI22_X1 U23846 ( .A1(READY2), .A2(keyinput_f37), .B1(
        P1_REIP_REG_27__SCAN_IN), .B2(keyinput_f56), .ZN(n20927) );
  OAI221_X1 U23847 ( .B1(READY2), .B2(keyinput_f37), .C1(
        P1_REIP_REG_27__SCAN_IN), .C2(keyinput_f56), .A(n20927), .ZN(n20930)
         );
  AOI22_X1 U23848 ( .A1(keyinput_f42), .A2(P1_D_C_N_REG_SCAN_IN), .B1(
        keyinput_f34), .B2(NA), .ZN(n20928) );
  OAI221_X1 U23849 ( .B1(keyinput_f42), .B2(P1_D_C_N_REG_SCAN_IN), .C1(
        keyinput_f34), .C2(NA), .A(n20928), .ZN(n20929) );
  NOR4_X1 U23850 ( .A1(n20932), .A2(n20931), .A3(n20930), .A4(n20929), .ZN(
        n20951) );
  AOI22_X1 U23851 ( .A1(keyinput_f39), .A2(P1_ADS_N_REG_SCAN_IN), .B1(DATAI_6_), .B2(keyinput_f26), .ZN(n20933) );
  OAI221_X1 U23852 ( .B1(keyinput_f39), .B2(P1_ADS_N_REG_SCAN_IN), .C1(
        DATAI_6_), .C2(keyinput_f26), .A(n20933), .ZN(n20940) );
  AOI22_X1 U23853 ( .A1(DATAI_30_), .A2(keyinput_f2), .B1(
        P1_REIP_REG_26__SCAN_IN), .B2(keyinput_f57), .ZN(n20934) );
  OAI221_X1 U23854 ( .B1(DATAI_30_), .B2(keyinput_f2), .C1(
        P1_REIP_REG_26__SCAN_IN), .C2(keyinput_f57), .A(n20934), .ZN(n20939)
         );
  AOI22_X1 U23855 ( .A1(n21098), .A2(keyinput_f61), .B1(keyinput_f0), .B2(
        n21011), .ZN(n20935) );
  OAI221_X1 U23856 ( .B1(n21098), .B2(keyinput_f61), .C1(n21011), .C2(
        keyinput_f0), .A(n20935), .ZN(n20938) );
  AOI22_X1 U23857 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(keyinput_f38), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(keyinput_f59), .ZN(n20936) );
  OAI221_X1 U23858 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_f38), .C1(
        P1_REIP_REG_24__SCAN_IN), .C2(keyinput_f59), .A(n20936), .ZN(n20937)
         );
  NOR4_X1 U23859 ( .A1(n20940), .A2(n20939), .A3(n20938), .A4(n20937), .ZN(
        n20950) );
  AOI22_X1 U23860 ( .A1(keyinput_f49), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        DATAI_31_), .B2(keyinput_f1), .ZN(n20941) );
  OAI221_X1 U23861 ( .B1(keyinput_f49), .B2(P1_BYTEENABLE_REG_1__SCAN_IN), 
        .C1(DATAI_31_), .C2(keyinput_f1), .A(n20941), .ZN(n20948) );
  AOI22_X1 U23862 ( .A1(DATAI_23_), .A2(keyinput_f9), .B1(DATAI_28_), .B2(
        keyinput_f4), .ZN(n20942) );
  OAI221_X1 U23863 ( .B1(DATAI_23_), .B2(keyinput_f9), .C1(DATAI_28_), .C2(
        keyinput_f4), .A(n20942), .ZN(n20947) );
  AOI22_X1 U23864 ( .A1(DATAI_2_), .A2(keyinput_f30), .B1(DATAI_5_), .B2(
        keyinput_f27), .ZN(n20943) );
  OAI221_X1 U23865 ( .B1(DATAI_2_), .B2(keyinput_f30), .C1(DATAI_5_), .C2(
        keyinput_f27), .A(n20943), .ZN(n20946) );
  AOI22_X1 U23866 ( .A1(keyinput_f33), .A2(HOLD), .B1(READY1), .B2(
        keyinput_f36), .ZN(n20944) );
  OAI221_X1 U23867 ( .B1(keyinput_f33), .B2(HOLD), .C1(READY1), .C2(
        keyinput_f36), .A(n20944), .ZN(n20945) );
  NOR4_X1 U23868 ( .A1(n20948), .A2(n20947), .A3(n20946), .A4(n20945), .ZN(
        n20949) );
  NAND4_X1 U23869 ( .A1(n20952), .A2(n20951), .A3(n20950), .A4(n20949), .ZN(
        n21004) );
  INV_X1 U23870 ( .A(DATAI_20_), .ZN(n20955) );
  INV_X1 U23871 ( .A(DATAI_14_), .ZN(n20954) );
  AOI22_X1 U23872 ( .A1(n20955), .A2(keyinput_f12), .B1(n20954), .B2(
        keyinput_f18), .ZN(n20953) );
  OAI221_X1 U23873 ( .B1(n20955), .B2(keyinput_f12), .C1(n20954), .C2(
        keyinput_f18), .A(n20953), .ZN(n20965) );
  AOI22_X1 U23874 ( .A1(n20957), .A2(keyinput_f46), .B1(n21040), .B2(
        keyinput_f54), .ZN(n20956) );
  OAI221_X1 U23875 ( .B1(n20957), .B2(keyinput_f46), .C1(n21040), .C2(
        keyinput_f54), .A(n20956), .ZN(n20964) );
  AOI22_X1 U23876 ( .A1(n21043), .A2(keyinput_f10), .B1(n20959), .B2(
        keyinput_f53), .ZN(n20958) );
  OAI221_X1 U23877 ( .B1(n21043), .B2(keyinput_f10), .C1(n20959), .C2(
        keyinput_f53), .A(n20958), .ZN(n20963) );
  INV_X1 U23878 ( .A(DATAI_8_), .ZN(n20961) );
  AOI22_X1 U23879 ( .A1(n21048), .A2(keyinput_f25), .B1(n20961), .B2(
        keyinput_f24), .ZN(n20960) );
  OAI221_X1 U23880 ( .B1(n21048), .B2(keyinput_f25), .C1(n20961), .C2(
        keyinput_f24), .A(n20960), .ZN(n20962) );
  NOR4_X1 U23881 ( .A1(n20965), .A2(n20964), .A3(n20963), .A4(n20962), .ZN(
        n21002) );
  AOI22_X1 U23882 ( .A1(n21032), .A2(keyinput_f52), .B1(keyinput_f41), .B2(
        n20967), .ZN(n20966) );
  OAI221_X1 U23883 ( .B1(n21032), .B2(keyinput_f52), .C1(n20967), .C2(
        keyinput_f41), .A(n20966), .ZN(n20977) );
  INV_X1 U23884 ( .A(DATAI_21_), .ZN(n20970) );
  AOI22_X1 U23885 ( .A1(n20970), .A2(keyinput_f11), .B1(keyinput_f51), .B2(
        n20969), .ZN(n20968) );
  OAI221_X1 U23886 ( .B1(n20970), .B2(keyinput_f11), .C1(n20969), .C2(
        keyinput_f51), .A(n20968), .ZN(n20976) );
  INV_X1 U23887 ( .A(DATAI_18_), .ZN(n20972) );
  INV_X1 U23888 ( .A(BS16), .ZN(n21064) );
  AOI22_X1 U23889 ( .A1(n20972), .A2(keyinput_f14), .B1(keyinput_f35), .B2(
        n21064), .ZN(n20971) );
  OAI221_X1 U23890 ( .B1(n20972), .B2(keyinput_f14), .C1(n21064), .C2(
        keyinput_f35), .A(n20971), .ZN(n20975) );
  INV_X1 U23891 ( .A(DATAI_15_), .ZN(n21030) );
  INV_X1 U23892 ( .A(DATAI_4_), .ZN(n21094) );
  AOI22_X1 U23893 ( .A1(n21030), .A2(keyinput_f17), .B1(n21094), .B2(
        keyinput_f28), .ZN(n20973) );
  OAI221_X1 U23894 ( .B1(n21030), .B2(keyinput_f17), .C1(n21094), .C2(
        keyinput_f28), .A(n20973), .ZN(n20974) );
  NOR4_X1 U23895 ( .A1(n20977), .A2(n20976), .A3(n20975), .A4(n20974), .ZN(
        n21001) );
  INV_X1 U23896 ( .A(DATAI_11_), .ZN(n21082) );
  AOI22_X1 U23897 ( .A1(n21082), .A2(keyinput_f21), .B1(keyinput_f50), .B2(
        n21016), .ZN(n20978) );
  OAI221_X1 U23898 ( .B1(n21082), .B2(keyinput_f21), .C1(n21016), .C2(
        keyinput_f50), .A(n20978), .ZN(n20986) );
  INV_X1 U23899 ( .A(DATAI_13_), .ZN(n20980) );
  AOI22_X1 U23900 ( .A1(n21058), .A2(keyinput_f60), .B1(keyinput_f19), .B2(
        n20980), .ZN(n20979) );
  OAI221_X1 U23901 ( .B1(n21058), .B2(keyinput_f60), .C1(n20980), .C2(
        keyinput_f19), .A(n20979), .ZN(n20985) );
  INV_X1 U23902 ( .A(DATAI_0_), .ZN(n21033) );
  AOI22_X1 U23903 ( .A1(n21033), .A2(keyinput_f32), .B1(n21091), .B2(
        keyinput_f7), .ZN(n20981) );
  OAI221_X1 U23904 ( .B1(n21033), .B2(keyinput_f32), .C1(n21091), .C2(
        keyinput_f7), .A(n20981), .ZN(n20984) );
  INV_X1 U23905 ( .A(DATAI_24_), .ZN(n21063) );
  INV_X1 U23906 ( .A(DATAI_3_), .ZN(n21024) );
  AOI22_X1 U23907 ( .A1(n21063), .A2(keyinput_f8), .B1(keyinput_f29), .B2(
        n21024), .ZN(n20982) );
  OAI221_X1 U23908 ( .B1(n21063), .B2(keyinput_f8), .C1(n21024), .C2(
        keyinput_f29), .A(n20982), .ZN(n20983) );
  NOR4_X1 U23909 ( .A1(n20986), .A2(n20985), .A3(n20984), .A4(n20983), .ZN(
        n21000) );
  INV_X1 U23910 ( .A(DATAI_10_), .ZN(n20988) );
  AOI22_X1 U23911 ( .A1(n20988), .A2(keyinput_f22), .B1(keyinput_f16), .B2(
        n21029), .ZN(n20987) );
  OAI221_X1 U23912 ( .B1(n20988), .B2(keyinput_f22), .C1(n21029), .C2(
        keyinput_f16), .A(n20987), .ZN(n20998) );
  AOI22_X1 U23913 ( .A1(n20990), .A2(keyinput_f58), .B1(keyinput_f48), .B2(
        n21027), .ZN(n20989) );
  OAI221_X1 U23914 ( .B1(n20990), .B2(keyinput_f58), .C1(n21027), .C2(
        keyinput_f48), .A(n20989), .ZN(n20997) );
  INV_X1 U23915 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n20992) );
  AOI22_X1 U23916 ( .A1(n21056), .A2(keyinput_f45), .B1(keyinput_f40), .B2(
        n20992), .ZN(n20991) );
  OAI221_X1 U23917 ( .B1(n21056), .B2(keyinput_f45), .C1(n20992), .C2(
        keyinput_f40), .A(n20991), .ZN(n20996) );
  INV_X1 U23918 ( .A(DATAI_1_), .ZN(n21010) );
  AOI22_X1 U23919 ( .A1(n21010), .A2(keyinput_f31), .B1(keyinput_f47), .B2(
        n20994), .ZN(n20993) );
  OAI221_X1 U23920 ( .B1(n21010), .B2(keyinput_f31), .C1(n20994), .C2(
        keyinput_f47), .A(n20993), .ZN(n20995) );
  NOR4_X1 U23921 ( .A1(n20998), .A2(n20997), .A3(n20996), .A4(n20995), .ZN(
        n20999) );
  NAND4_X1 U23922 ( .A1(n21002), .A2(n21001), .A3(n21000), .A4(n20999), .ZN(
        n21003) );
  OAI22_X1 U23923 ( .A1(n21004), .A2(n21003), .B1(keyinput_f63), .B2(
        P1_REIP_REG_20__SCAN_IN), .ZN(n21005) );
  AOI21_X1 U23924 ( .B1(keyinput_f63), .B2(P1_REIP_REG_20__SCAN_IN), .A(n21005), .ZN(n21118) );
  AOI22_X1 U23925 ( .A1(n21008), .A2(keyinput_g6), .B1(n21007), .B2(
        keyinput_g57), .ZN(n21006) );
  OAI221_X1 U23926 ( .B1(n21008), .B2(keyinput_g6), .C1(n21007), .C2(
        keyinput_g57), .A(n21006), .ZN(n21021) );
  AOI22_X1 U23927 ( .A1(n21011), .A2(keyinput_g0), .B1(n21010), .B2(
        keyinput_g31), .ZN(n21009) );
  OAI221_X1 U23928 ( .B1(n21011), .B2(keyinput_g0), .C1(n21010), .C2(
        keyinput_g31), .A(n21009), .ZN(n21020) );
  AOI22_X1 U23929 ( .A1(n21014), .A2(keyinput_g13), .B1(keyinput_g34), .B2(
        n21013), .ZN(n21012) );
  OAI221_X1 U23930 ( .B1(n21014), .B2(keyinput_g13), .C1(n21013), .C2(
        keyinput_g34), .A(n21012), .ZN(n21019) );
  INV_X1 U23931 ( .A(DATAI_30_), .ZN(n21017) );
  AOI22_X1 U23932 ( .A1(n21017), .A2(keyinput_g2), .B1(keyinput_g50), .B2(
        n21016), .ZN(n21015) );
  OAI221_X1 U23933 ( .B1(n21017), .B2(keyinput_g2), .C1(n21016), .C2(
        keyinput_g50), .A(n21015), .ZN(n21018) );
  NOR4_X1 U23934 ( .A1(n21021), .A2(n21020), .A3(n21019), .A4(n21018), .ZN(
        n21072) );
  AOI22_X1 U23935 ( .A1(n21024), .A2(keyinput_g29), .B1(n21023), .B2(
        keyinput_g55), .ZN(n21022) );
  OAI221_X1 U23936 ( .B1(n21024), .B2(keyinput_g29), .C1(n21023), .C2(
        keyinput_g55), .A(n21022), .ZN(n21037) );
  AOI22_X1 U23937 ( .A1(n21027), .A2(keyinput_g48), .B1(n21026), .B2(
        keyinput_g59), .ZN(n21025) );
  OAI221_X1 U23938 ( .B1(n21027), .B2(keyinput_g48), .C1(n21026), .C2(
        keyinput_g59), .A(n21025), .ZN(n21036) );
  AOI22_X1 U23939 ( .A1(n21030), .A2(keyinput_g17), .B1(n21029), .B2(
        keyinput_g16), .ZN(n21028) );
  OAI221_X1 U23940 ( .B1(n21030), .B2(keyinput_g17), .C1(n21029), .C2(
        keyinput_g16), .A(n21028), .ZN(n21035) );
  AOI22_X1 U23941 ( .A1(n21033), .A2(keyinput_g32), .B1(n21032), .B2(
        keyinput_g52), .ZN(n21031) );
  OAI221_X1 U23942 ( .B1(n21033), .B2(keyinput_g32), .C1(n21032), .C2(
        keyinput_g52), .A(n21031), .ZN(n21034) );
  NOR4_X1 U23943 ( .A1(n21037), .A2(n21036), .A3(n21035), .A4(n21034), .ZN(
        n21071) );
  INV_X1 U23944 ( .A(DATAI_6_), .ZN(n21039) );
  AOI22_X1 U23945 ( .A1(n21040), .A2(keyinput_g54), .B1(keyinput_g26), .B2(
        n21039), .ZN(n21038) );
  OAI221_X1 U23946 ( .B1(n21040), .B2(keyinput_g54), .C1(n21039), .C2(
        keyinput_g26), .A(n21038), .ZN(n21053) );
  AOI22_X1 U23947 ( .A1(n21043), .A2(keyinput_g10), .B1(n21042), .B2(
        keyinput_g62), .ZN(n21041) );
  OAI221_X1 U23948 ( .B1(n21043), .B2(keyinput_g10), .C1(n21042), .C2(
        keyinput_g62), .A(n21041), .ZN(n21052) );
  INV_X1 U23949 ( .A(DATAI_9_), .ZN(n21046) );
  INV_X1 U23950 ( .A(DATAI_17_), .ZN(n21045) );
  AOI22_X1 U23951 ( .A1(n21046), .A2(keyinput_g23), .B1(keyinput_g15), .B2(
        n21045), .ZN(n21044) );
  OAI221_X1 U23952 ( .B1(n21046), .B2(keyinput_g23), .C1(n21045), .C2(
        keyinput_g15), .A(n21044), .ZN(n21051) );
  AOI22_X1 U23953 ( .A1(n21049), .A2(keyinput_g1), .B1(keyinput_g25), .B2(
        n21048), .ZN(n21047) );
  OAI221_X1 U23954 ( .B1(n21049), .B2(keyinput_g1), .C1(n21048), .C2(
        keyinput_g25), .A(n21047), .ZN(n21050) );
  NOR4_X1 U23955 ( .A1(n21053), .A2(n21052), .A3(n21051), .A4(n21050), .ZN(
        n21070) );
  INV_X1 U23956 ( .A(DATAI_27_), .ZN(n21055) );
  AOI22_X1 U23957 ( .A1(n21056), .A2(keyinput_g45), .B1(n21055), .B2(
        keyinput_g5), .ZN(n21054) );
  OAI221_X1 U23958 ( .B1(n21056), .B2(keyinput_g45), .C1(n21055), .C2(
        keyinput_g5), .A(n21054), .ZN(n21068) );
  AOI22_X1 U23959 ( .A1(n21058), .A2(keyinput_g60), .B1(keyinput_g9), .B2(
        n14768), .ZN(n21057) );
  OAI221_X1 U23960 ( .B1(n21058), .B2(keyinput_g60), .C1(n14768), .C2(
        keyinput_g9), .A(n21057), .ZN(n21067) );
  INV_X1 U23961 ( .A(DATAI_2_), .ZN(n21060) );
  AOI22_X1 U23962 ( .A1(n21061), .A2(keyinput_g42), .B1(n21060), .B2(
        keyinput_g30), .ZN(n21059) );
  OAI221_X1 U23963 ( .B1(n21061), .B2(keyinput_g42), .C1(n21060), .C2(
        keyinput_g30), .A(n21059), .ZN(n21066) );
  AOI22_X1 U23964 ( .A1(n21064), .A2(keyinput_g35), .B1(n21063), .B2(
        keyinput_g8), .ZN(n21062) );
  OAI221_X1 U23965 ( .B1(n21064), .B2(keyinput_g35), .C1(n21063), .C2(
        keyinput_g8), .A(n21062), .ZN(n21065) );
  NOR4_X1 U23966 ( .A1(n21068), .A2(n21067), .A3(n21066), .A4(n21065), .ZN(
        n21069) );
  NAND4_X1 U23967 ( .A1(n21072), .A2(n21071), .A3(n21070), .A4(n21069), .ZN(
        n21116) );
  AOI22_X1 U23968 ( .A1(DATAI_13_), .A2(keyinput_g19), .B1(DATAI_29_), .B2(
        keyinput_g3), .ZN(n21073) );
  OAI221_X1 U23969 ( .B1(DATAI_13_), .B2(keyinput_g19), .C1(DATAI_29_), .C2(
        keyinput_g3), .A(n21073), .ZN(n21080) );
  AOI22_X1 U23970 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(keyinput_g40), .B1(
        DATAI_21_), .B2(keyinput_g11), .ZN(n21074) );
  OAI221_X1 U23971 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_g40), .C1(
        DATAI_21_), .C2(keyinput_g11), .A(n21074), .ZN(n21079) );
  AOI22_X1 U23972 ( .A1(DATAI_12_), .A2(keyinput_g20), .B1(
        P1_REIP_REG_27__SCAN_IN), .B2(keyinput_g56), .ZN(n21075) );
  OAI221_X1 U23973 ( .B1(DATAI_12_), .B2(keyinput_g20), .C1(
        P1_REIP_REG_27__SCAN_IN), .C2(keyinput_g56), .A(n21075), .ZN(n21078)
         );
  AOI22_X1 U23974 ( .A1(HOLD), .A2(keyinput_g33), .B1(
        P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_g38), .ZN(n21076) );
  OAI221_X1 U23975 ( .B1(HOLD), .B2(keyinput_g33), .C1(
        P1_READREQUEST_REG_SCAN_IN), .C2(keyinput_g38), .A(n21076), .ZN(n21077) );
  NOR4_X1 U23976 ( .A1(n21080), .A2(n21079), .A3(n21078), .A4(n21077), .ZN(
        n21114) );
  XNOR2_X1 U23977 ( .A(DATAI_18_), .B(keyinput_g14), .ZN(n21088) );
  AOI22_X1 U23978 ( .A1(DATAI_8_), .A2(keyinput_g24), .B1(n21082), .B2(
        keyinput_g21), .ZN(n21081) );
  OAI221_X1 U23979 ( .B1(DATAI_8_), .B2(keyinput_g24), .C1(n21082), .C2(
        keyinput_g21), .A(n21081), .ZN(n21087) );
  AOI22_X1 U23980 ( .A1(P1_M_IO_N_REG_SCAN_IN), .A2(keyinput_g41), .B1(
        P1_ADS_N_REG_SCAN_IN), .B2(keyinput_g39), .ZN(n21083) );
  OAI221_X1 U23981 ( .B1(P1_M_IO_N_REG_SCAN_IN), .B2(keyinput_g41), .C1(
        P1_ADS_N_REG_SCAN_IN), .C2(keyinput_g39), .A(n21083), .ZN(n21086) );
  AOI22_X1 U23982 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(keyinput_g46), .B1(
        DATAI_20_), .B2(keyinput_g12), .ZN(n21084) );
  OAI221_X1 U23983 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(keyinput_g46), .C1(
        DATAI_20_), .C2(keyinput_g12), .A(n21084), .ZN(n21085) );
  NOR4_X1 U23984 ( .A1(n21088), .A2(n21087), .A3(n21086), .A4(n21085), .ZN(
        n21113) );
  INV_X1 U23985 ( .A(READY1), .ZN(n21090) );
  AOI22_X1 U23986 ( .A1(n21091), .A2(keyinput_g7), .B1(n21090), .B2(
        keyinput_g36), .ZN(n21089) );
  OAI221_X1 U23987 ( .B1(n21091), .B2(keyinput_g7), .C1(n21090), .C2(
        keyinput_g36), .A(n21089), .ZN(n21102) );
  AOI22_X1 U23988 ( .A1(P1_W_R_N_REG_SCAN_IN), .A2(keyinput_g47), .B1(DATAI_5_), .B2(keyinput_g27), .ZN(n21092) );
  OAI221_X1 U23989 ( .B1(P1_W_R_N_REG_SCAN_IN), .B2(keyinput_g47), .C1(
        DATAI_5_), .C2(keyinput_g27), .A(n21092), .ZN(n21101) );
  AOI22_X1 U23990 ( .A1(n21095), .A2(keyinput_g44), .B1(keyinput_g28), .B2(
        n21094), .ZN(n21093) );
  OAI221_X1 U23991 ( .B1(n21095), .B2(keyinput_g44), .C1(n21094), .C2(
        keyinput_g28), .A(n21093), .ZN(n21100) );
  AOI22_X1 U23992 ( .A1(n21098), .A2(keyinput_g61), .B1(keyinput_g4), .B2(
        n21097), .ZN(n21096) );
  OAI221_X1 U23993 ( .B1(n21098), .B2(keyinput_g61), .C1(n21097), .C2(
        keyinput_g4), .A(n21096), .ZN(n21099) );
  NOR4_X1 U23994 ( .A1(n21102), .A2(n21101), .A3(n21100), .A4(n21099), .ZN(
        n21112) );
  AOI22_X1 U23995 ( .A1(READY2), .A2(keyinput_g37), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(keyinput_g53), .ZN(n21103) );
  OAI221_X1 U23996 ( .B1(READY2), .B2(keyinput_g37), .C1(
        P1_REIP_REG_30__SCAN_IN), .C2(keyinput_g53), .A(n21103), .ZN(n21110)
         );
  AOI22_X1 U23997 ( .A1(DATAI_10_), .A2(keyinput_g22), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(keyinput_g58), .ZN(n21104) );
  OAI221_X1 U23998 ( .B1(DATAI_10_), .B2(keyinput_g22), .C1(
        P1_REIP_REG_25__SCAN_IN), .C2(keyinput_g58), .A(n21104), .ZN(n21109)
         );
  AOI22_X1 U23999 ( .A1(P1_BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_g49), .B1(
        DATAI_14_), .B2(keyinput_g18), .ZN(n21105) );
  OAI221_X1 U24000 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_g49), 
        .C1(DATAI_14_), .C2(keyinput_g18), .A(n21105), .ZN(n21108) );
  AOI22_X1 U24001 ( .A1(P1_BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_g51), .B1(
        P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_g43), .ZN(n21106) );
  OAI221_X1 U24002 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_g51), 
        .C1(P1_REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_g43), .A(n21106), 
        .ZN(n21107) );
  NOR4_X1 U24003 ( .A1(n21110), .A2(n21109), .A3(n21108), .A4(n21107), .ZN(
        n21111) );
  NAND4_X1 U24004 ( .A1(n21114), .A2(n21113), .A3(n21112), .A4(n21111), .ZN(
        n21115) );
  OAI22_X1 U24005 ( .A1(keyinput_g63), .A2(n21119), .B1(n21116), .B2(n21115), 
        .ZN(n21117) );
  AOI211_X1 U24006 ( .C1(keyinput_g63), .C2(n21119), .A(n21118), .B(n21117), 
        .ZN(n21121) );
  AOI22_X1 U24007 ( .A1(n16804), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16806), .ZN(n21120) );
  XNOR2_X1 U24008 ( .A(n21121), .B(n21120), .ZN(U355) );
  AND2_X1 U11480 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14062) );
  AND2_X1 U11219 ( .A1(n14064), .A2(n10907), .ZN(n10933) );
  OR2_X1 U16042 ( .A1(n14980), .A2(n20226), .ZN(n12917) );
  NAND2_X2 U11145 ( .A1(n9657), .A2(n9658), .ZN(n16615) );
  CLKBUF_X1 U11138 ( .A(n10998), .Z(n11050) );
  CLKBUF_X1 U11143 ( .A(n11807), .Z(n11797) );
  CLKBUF_X1 U11160 ( .A(n11943), .Z(n11940) );
  NAND2_X2 U11172 ( .A1(n9684), .A2(n11808), .ZN(n11892) );
  NOR2_X2 U11173 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10908) );
  CLKBUF_X1 U11179 ( .A(n10845), .Z(n10838) );
  CLKBUF_X1 U11184 ( .A(n12446), .Z(n12537) );
  NAND2_X1 U11185 ( .A1(n12574), .A2(n12551), .ZN(n13950) );
  BUF_X1 U11191 ( .A(n10642), .Z(n12504) );
  NAND2_X2 U11223 ( .A1(n13508), .A2(n14062), .ZN(n14059) );
  CLKBUF_X1 U11246 ( .A(n10692), .Z(n10654) );
  CLKBUF_X1 U11376 ( .A(n12556), .Z(n19559) );
  NOR2_X1 U11387 ( .A1(n9716), .A2(n9669), .ZN(n21122) );
  OR2_X1 U11440 ( .A1(n10657), .A2(n19583), .ZN(n21123) );
  CLKBUF_X1 U11443 ( .A(n19166), .Z(n17724) );
endmodule

