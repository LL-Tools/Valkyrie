

module b15_C_SARLock_k_64_7 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690;

  INV_X1 U3405 ( .A(n6057), .ZN(n6041) );
  CLKBUF_X2 U3406 ( .A(n4106), .Z(n4215) );
  INV_X1 U3407 ( .A(n4169), .ZN(n3289) );
  INV_X1 U3408 ( .A(n3538), .ZN(n3559) );
  INV_X4 U3409 ( .A(n4993), .ZN(n4332) );
  OR2_X1 U3410 ( .A1(n3099), .A2(n3098), .ZN(n3219) );
  INV_X1 U3411 ( .A(n3218), .ZN(n3210) );
  AND2_X1 U3412 ( .A1(n4447), .A2(n4528), .ZN(n4106) );
  AND2_X1 U3413 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4548) );
  CLKBUF_X2 U3414 ( .A(n3183), .Z(n4195) );
  AND2_X1 U3415 ( .A1(n4439), .A2(n3083), .ZN(n3316) );
  NAND2_X1 U3416 ( .A1(n5561), .A2(n4998), .ZN(n3705) );
  INV_X2 U3417 ( .A(n3705), .ZN(n3001) );
  NAND2_X1 U3418 ( .A1(n3066), .A2(n3063), .ZN(n5423) );
  INV_X1 U3419 ( .A(n6024), .ZN(n6038) );
  NAND2_X2 U3422 ( .A1(n3283), .A2(n3281), .ZN(n3304) );
  NAND2_X2 U3423 ( .A1(n6147), .A2(n6146), .ZN(n6145) );
  NAND2_X2 U3424 ( .A1(n4596), .A2(n3441), .ZN(n6147) );
  XNOR2_X1 U3425 ( .A(n3369), .B(n3370), .ZN(n4562) );
  NOR2_X2 U3426 ( .A1(n4490), .A2(n4501), .ZN(n4493) );
  NOR2_X1 U3428 ( .A1(n5835), .A2(n5836), .ZN(n5834) );
  OAI21_X1 U3429 ( .B1(n3204), .B2(n3203), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3229) );
  INV_X2 U3430 ( .A(n5561), .ZN(n3617) );
  AND2_X1 U3433 ( .A1(n2973), .A2(n3148), .ZN(n3712) );
  AND4_X1 U3434 ( .A1(n3188), .A2(n3187), .A3(n3186), .A4(n3185), .ZN(n3189)
         );
  CLKBUF_X2 U3435 ( .A(n3267), .Z(n4532) );
  BUF_X2 U3436 ( .A(n3266), .Z(n4174) );
  CLKBUF_X2 U3437 ( .A(n3172), .Z(n4173) );
  CLKBUF_X2 U3438 ( .A(n3174), .Z(n4208) );
  BUF_X2 U3439 ( .A(n3316), .Z(n3261) );
  CLKBUF_X2 U3440 ( .A(n4517), .Z(n6521) );
  CLKBUF_X2 U3441 ( .A(n3184), .Z(n4210) );
  AND2_X2 U3442 ( .A1(n3000), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4444)
         );
  AND2_X1 U3443 ( .A1(n4237), .A2(n4236), .ZN(n5608) );
  AOI211_X1 U3444 ( .C1(n5728), .C2(n5629), .A(n5628), .B(n5627), .ZN(n5630)
         );
  XNOR2_X1 U34450 ( .A(n2992), .B(n4282), .ZN(n4306) );
  NAND2_X1 U34460 ( .A1(n3514), .A2(n3074), .ZN(n3515) );
  INV_X1 U34470 ( .A(n2993), .ZN(n4272) );
  OAI21_X1 U34480 ( .B1(n5436), .B2(n5438), .A(n5437), .ZN(n5626) );
  CLKBUF_X1 U3449 ( .A(n3512), .Z(n3513) );
  NAND2_X1 U3450 ( .A1(n5677), .A2(n5646), .ZN(n3030) );
  OAI21_X1 U34510 ( .B1(n4697), .B2(n2970), .A(n5017), .ZN(n2997) );
  XNOR2_X1 U34520 ( .A(n3480), .B(n3479), .ZN(n4697) );
  AOI21_X1 U34530 ( .B1(n3802), .B2(n3916), .A(n3801), .ZN(n4587) );
  AND2_X1 U3454 ( .A1(n3368), .A2(n3076), .ZN(n6154) );
  XNOR2_X1 U34550 ( .A(n3485), .B(n3472), .ZN(n3802) );
  NAND2_X1 U34560 ( .A1(n2999), .A2(n3458), .ZN(n3485) );
  OR2_X1 U3457 ( .A1(n3764), .A2(n4484), .ZN(n4396) );
  AND2_X1 U3458 ( .A1(n4482), .A2(n4481), .ZN(n4484) );
  OR2_X1 U34590 ( .A1(n6163), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3076)
         );
  NAND2_X1 U34600 ( .A1(n2998), .A2(n3370), .ZN(n3400) );
  NAND2_X1 U34610 ( .A1(n3391), .A2(n3390), .ZN(n4706) );
  CLKBUF_X1 U34620 ( .A(n4559), .Z(n5098) );
  NAND2_X1 U34630 ( .A1(n3329), .A2(n3328), .ZN(n3332) );
  NAND2_X1 U34640 ( .A1(n3344), .A2(n3343), .ZN(n4559) );
  AND2_X1 U34650 ( .A1(n3229), .A2(n3226), .ZN(n3225) );
  OR2_X1 U3466 ( .A1(n3229), .A2(n3228), .ZN(n3230) );
  NOR2_X1 U3467 ( .A1(n4331), .A2(n3209), .ZN(n3203) );
  AND3_X1 U34680 ( .A1(n3197), .A2(n3215), .A3(n3214), .ZN(n3587) );
  AND2_X1 U34690 ( .A1(n3222), .A2(n4420), .ZN(n3239) );
  OR2_X1 U34700 ( .A1(n3601), .A2(n3520), .ZN(n3596) );
  AND2_X1 U34710 ( .A1(n4240), .A2(n3333), .ZN(n3241) );
  INV_X1 U34720 ( .A(n4998), .ZN(n2956) );
  NAND2_X1 U34730 ( .A1(n3193), .A2(n3218), .ZN(n4391) );
  AND2_X2 U34740 ( .A1(n3605), .A2(n4993), .ZN(n4241) );
  INV_X1 U3475 ( .A(n3220), .ZN(n4325) );
  AND2_X1 U3476 ( .A1(n3192), .A2(n3220), .ZN(n4327) );
  CLKBUF_X3 U3477 ( .A(n4631), .Z(n2958) );
  NAND2_X1 U3478 ( .A1(n3712), .A2(n3219), .ZN(n3714) );
  INV_X1 U3479 ( .A(n3712), .ZN(n4621) );
  BUF_X2 U3480 ( .A(n3170), .Z(n3220) );
  NAND4_X1 U3481 ( .A1(n3139), .A2(n3138), .A3(n3137), .A4(n3136), .ZN(n4631)
         );
  OR2_X1 U3482 ( .A1(n3169), .A2(n3168), .ZN(n3170) );
  AND4_X1 U3483 ( .A1(n3135), .A2(n3134), .A3(n3133), .A4(n3132), .ZN(n3136)
         );
  AND4_X1 U3484 ( .A1(n3087), .A2(n3086), .A3(n3085), .A4(n3084), .ZN(n3088)
         );
  AND4_X1 U3485 ( .A1(n3147), .A2(n3146), .A3(n3145), .A4(n3144), .ZN(n3148)
         );
  AND4_X1 U3486 ( .A1(n3131), .A2(n3130), .A3(n3129), .A4(n3128), .ZN(n3137)
         );
  AND4_X1 U3487 ( .A1(n3082), .A2(n3081), .A3(n3080), .A4(n3079), .ZN(n3089)
         );
  AND4_X1 U3488 ( .A1(n3103), .A2(n3102), .A3(n3101), .A4(n3100), .ZN(n3119)
         );
  AND4_X1 U3489 ( .A1(n3127), .A2(n3126), .A3(n3125), .A4(n3124), .ZN(n3138)
         );
  AND4_X1 U3490 ( .A1(n3123), .A2(n3122), .A3(n3121), .A4(n3120), .ZN(n3139)
         );
  AND4_X1 U3491 ( .A1(n3153), .A2(n3152), .A3(n3151), .A4(n3150), .ZN(n3159)
         );
  AND4_X1 U3492 ( .A1(n3157), .A2(n3156), .A3(n3155), .A4(n3154), .ZN(n3158)
         );
  AND4_X1 U3493 ( .A1(n3178), .A2(n3177), .A3(n3176), .A4(n3175), .ZN(n3190)
         );
  BUF_X2 U3494 ( .A(n3247), .Z(n4216) );
  BUF_X2 U3495 ( .A(n3284), .Z(n3803) );
  BUF_X1 U3496 ( .A(n3179), .Z(n3253) );
  BUF_X2 U3497 ( .A(n3173), .Z(n4209) );
  BUF_X2 U3498 ( .A(n3182), .Z(n3290) );
  AND2_X2 U3499 ( .A1(n4444), .A2(n4530), .ZN(n3183) );
  AND2_X2 U3500 ( .A1(n3048), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4530)
         );
  NAND2_X1 U3501 ( .A1(n5611), .A2(n2990), .ZN(n2993) );
  INV_X1 U3502 ( .A(n3369), .ZN(n2998) );
  OAI21_X1 U3503 ( .B1(n4307), .B2(n4309), .A(n4308), .ZN(n5587) );
  AND2_X1 U3504 ( .A1(n3218), .A2(n4631), .ZN(n3333) );
  AND2_X4 U3505 ( .A1(n4439), .A2(n4548), .ZN(n3181) );
  OR2_X2 U3506 ( .A1(n4988), .A2(n4986), .ZN(n6024) );
  AND2_X1 U3507 ( .A1(n4439), .A2(n3083), .ZN(n2959) );
  INV_X1 U3508 ( .A(n3253), .ZN(n2960) );
  AND2_X4 U3509 ( .A1(n4447), .A2(n3083), .ZN(n3179) );
  XNOR2_X1 U3510 ( .A(n4410), .B(n4603), .ZN(n4527) );
  AND2_X1 U3511 ( .A1(n4447), .A2(n4528), .ZN(n2962) );
  NAND2_X2 U3512 ( .A1(n5690), .A2(n3505), .ZN(n5710) );
  NOR2_X2 U3513 ( .A1(n5442), .A2(n5425), .ZN(n5426) );
  XNOR2_X2 U3514 ( .A(n3400), .B(n4706), .ZN(n3767) );
  BUF_X2 U3515 ( .A(n4563), .Z(n2963) );
  AND2_X4 U3516 ( .A1(n4993), .A2(n2958), .ZN(n4998) );
  NOR2_X1 U3517 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6614), .ZN(n3531)
         );
  INV_X1 U3518 ( .A(n3460), .ZN(n2999) );
  OR2_X1 U3519 ( .A1(n3273), .A2(n3272), .ZN(n3481) );
  NAND2_X1 U3520 ( .A1(n5554), .A2(n3060), .ZN(n3059) );
  INV_X1 U3521 ( .A(n3061), .ZN(n3060) );
  NOR2_X1 U3522 ( .A1(n2970), .A2(n3038), .ZN(n3036) );
  INV_X1 U3523 ( .A(n4494), .ZN(n3051) );
  NOR2_X2 U3524 ( .A1(n3192), .A2(n5069), .ZN(n3916) );
  NOR2_X1 U3525 ( .A1(n4993), .A2(n2958), .ZN(n3198) );
  AND2_X1 U3526 ( .A1(n3201), .A2(n3206), .ZN(n3518) );
  XNOR2_X1 U3527 ( .A(n3611), .B(n4361), .ZN(n4452) );
  INV_X1 U3528 ( .A(n5710), .ZN(n3506) );
  OR2_X1 U3529 ( .A1(n3028), .A2(n5647), .ZN(n3025) );
  INV_X1 U3530 ( .A(n3496), .ZN(n3492) );
  AND2_X1 U3531 ( .A1(n3611), .A2(n5199), .ZN(n3009) );
  INV_X1 U3532 ( .A(n3199), .ZN(n4240) );
  NAND2_X1 U3533 ( .A1(n3569), .A2(n3568), .ZN(n5401) );
  INV_X1 U3534 ( .A(n6198), .ZN(n6237) );
  BUF_X1 U3535 ( .A(n3819), .Z(n4150) );
  NAND2_X1 U3536 ( .A1(n3420), .A2(n3447), .ZN(n3460) );
  AND2_X2 U3537 ( .A1(n3078), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3083)
         );
  OR2_X1 U3538 ( .A1(n4438), .A2(n4400), .ZN(n3723) );
  NOR2_X1 U3539 ( .A1(n3064), .A2(n3069), .ZN(n3063) );
  INV_X1 U3540 ( .A(n5438), .ZN(n3069) );
  INV_X1 U3541 ( .A(n3755), .ZN(n3984) );
  INV_X1 U3542 ( .A(n3984), .ZN(n4227) );
  NAND2_X1 U3543 ( .A1(n5069), .A2(n6424), .ZN(n4233) );
  INV_X1 U3544 ( .A(n5453), .ZN(n3017) );
  NOR2_X1 U3545 ( .A1(n3483), .A2(n3482), .ZN(n3484) );
  AND2_X1 U3546 ( .A1(n4422), .A2(n3722), .ZN(n4239) );
  OR2_X1 U3547 ( .A1(n6010), .A2(n3005), .ZN(n3004) );
  AND2_X1 U3548 ( .A1(n4998), .A2(n3617), .ZN(n3690) );
  NOR2_X1 U3549 ( .A1(n3723), .A2(n5401), .ZN(n4238) );
  AOI21_X1 U3550 ( .B1(n3532), .B2(n3528), .A(n3531), .ZN(n3575) );
  OAI21_X1 U3551 ( .B1(n3307), .B2(n3306), .A(n3305), .ZN(n3371) );
  NAND2_X1 U3552 ( .A1(n3315), .A2(n3314), .ZN(n3372) );
  AND4_X1 U3553 ( .A1(n3107), .A2(n3106), .A3(n3105), .A4(n3104), .ZN(n3118)
         );
  AND2_X1 U3554 ( .A1(n4526), .A2(n4525), .ZN(n6397) );
  AND2_X1 U3555 ( .A1(n5396), .A2(n4330), .ZN(n5404) );
  OR2_X1 U3556 ( .A1(n6518), .A2(n4985), .ZN(n5378) );
  NAND2_X1 U3557 ( .A1(n5378), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5375) );
  NOR2_X1 U3558 ( .A1(n2971), .A2(n5330), .ZN(n5317) );
  NOR2_X1 U3559 ( .A1(n4589), .A2(n4590), .ZN(n4802) );
  NOR2_X1 U3560 ( .A1(n3220), .A2(n5069), .ZN(n3755) );
  INV_X1 U3561 ( .A(n3883), .ZN(n4288) );
  NAND2_X1 U3562 ( .A1(n4207), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4293)
         );
  INV_X1 U3563 ( .A(n4206), .ZN(n4207) );
  BUF_X1 U3564 ( .A(n4234), .Z(n4308) );
  NAND2_X1 U3565 ( .A1(n4039), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4085)
         );
  NAND2_X1 U3566 ( .A1(n3058), .A2(n4057), .ZN(n3057) );
  INV_X1 U3567 ( .A(n3059), .ZN(n3058) );
  OAI21_X1 U3568 ( .B1(n5710), .B2(n3044), .A(n3042), .ZN(n5684) );
  INV_X1 U3569 ( .A(n2997), .ZN(n3037) );
  NAND2_X1 U3570 ( .A1(n6145), .A2(n3036), .ZN(n3035) );
  NAND2_X1 U3571 ( .A1(n3796), .A2(n4643), .ZN(n3050) );
  NAND2_X1 U3572 ( .A1(n3051), .A2(n3796), .ZN(n4588) );
  OR2_X1 U3573 ( .A1(n4352), .A2(n3759), .ZN(n4353) );
  NAND2_X1 U3574 ( .A1(n5540), .A2(n3015), .ZN(n5442) );
  AND2_X1 U3575 ( .A1(n2983), .A2(n3016), .ZN(n3015) );
  INV_X1 U3576 ( .A(n5440), .ZN(n3016) );
  AND2_X1 U3577 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  AND2_X1 U3578 ( .A1(n2980), .A2(n5778), .ZN(n3024) );
  INV_X1 U3579 ( .A(n3025), .ZN(n3023) );
  AOI21_X1 U3580 ( .B1(n3025), .B2(n3022), .A(n3021), .ZN(n3020) );
  NAND2_X1 U3581 ( .A1(n5648), .A2(n2987), .ZN(n3021) );
  INV_X1 U3582 ( .A(n3026), .ZN(n3022) );
  NOR2_X1 U3583 ( .A1(n5647), .A2(n3027), .ZN(n3026) );
  INV_X1 U3584 ( .A(n5646), .ZN(n3027) );
  NOR2_X1 U3585 ( .A1(n3031), .A2(n3029), .ZN(n3028) );
  INV_X1 U3586 ( .A(n5671), .ZN(n3029) );
  NOR2_X1 U3587 ( .A1(n2977), .A2(n2996), .ZN(n2995) );
  INV_X1 U3588 ( .A(n3500), .ZN(n2996) );
  AND3_X1 U3589 ( .A1(n3010), .A2(n3009), .A3(n3008), .ZN(n6043) );
  INV_X1 U3590 ( .A(n6045), .ZN(n3008) );
  NAND2_X1 U3591 ( .A1(n3001), .A2(n3604), .ZN(n3608) );
  AND2_X1 U3592 ( .A1(n3730), .A2(n5346), .ZN(n5332) );
  AND2_X1 U3593 ( .A1(n3587), .A2(n4332), .ZN(n5396) );
  XNOR2_X1 U3594 ( .A(n3711), .B(n3710), .ZN(n5529) );
  AND2_X1 U3595 ( .A1(n5581), .A2(n4327), .ZN(n6081) );
  AND2_X1 U3596 ( .A1(n5581), .A2(n5580), .ZN(n6085) );
  AND2_X1 U3597 ( .A1(n3210), .A2(n3220), .ZN(n5580) );
  AND2_X1 U3598 ( .A1(n5581), .A2(n4393), .ZN(n5357) );
  CLKBUF_X1 U3599 ( .A(n6130), .Z(n6126) );
  INV_X1 U3600 ( .A(n3040), .ZN(n3039) );
  OAI21_X1 U3601 ( .B1(n3043), .B2(n3041), .A(n5683), .ZN(n3040) );
  INV_X1 U3602 ( .A(n3042), .ZN(n3041) );
  INV_X1 U3603 ( .A(n5725), .ZN(n6161) );
  INV_X1 U3604 ( .A(n6144), .ZN(n6165) );
  OR2_X1 U3605 ( .A1(n6380), .A2(n6418), .ZN(n6144) );
  NAND2_X1 U3606 ( .A1(n2993), .A2(n4271), .ZN(n2992) );
  INV_X1 U3607 ( .A(n5271), .ZN(n5831) );
  NAND2_X1 U3608 ( .A1(n3725), .A2(n3603), .ZN(n6198) );
  AND2_X1 U3609 ( .A1(n6404), .A2(n6403), .ZN(n6419) );
  NAND3_X1 U3610 ( .A1(n2998), .A2(n4706), .A3(n3370), .ZN(n3442) );
  OR2_X1 U3611 ( .A1(n3410), .A2(n3409), .ZN(n3462) );
  OR2_X1 U3612 ( .A1(n3259), .A2(n3258), .ZN(n3359) );
  AND2_X1 U3613 ( .A1(n3571), .A2(n3576), .ZN(n3563) );
  NAND2_X1 U3614 ( .A1(n4332), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3379) );
  INV_X1 U3615 ( .A(n4296), .ZN(n3313) );
  INV_X1 U3616 ( .A(n3192), .ZN(n3193) );
  AOI22_X1 U3617 ( .A1(n3180), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3147) );
  AOI22_X1 U3618 ( .A1(n3284), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3144) );
  OR2_X1 U3619 ( .A1(n3389), .A2(n3388), .ZN(n3413) );
  INV_X1 U3620 ( .A(n5537), .ZN(n3065) );
  NOR2_X1 U3621 ( .A1(n5450), .A2(n3068), .ZN(n3067) );
  INV_X1 U3622 ( .A(n5463), .ZN(n3068) );
  NAND2_X1 U3623 ( .A1(n4022), .A2(n3062), .ZN(n3061) );
  NAND2_X1 U3624 ( .A1(n5648), .A2(n3727), .ZN(n3045) );
  NOR2_X1 U3625 ( .A1(n3071), .A2(n3054), .ZN(n3053) );
  INV_X1 U3626 ( .A(n5515), .ZN(n3054) );
  AND2_X1 U3627 ( .A1(n2981), .A2(n3849), .ZN(n3052) );
  NAND2_X1 U3628 ( .A1(n3851), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3866)
         );
  INV_X1 U3629 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3865) );
  NAND2_X1 U3630 ( .A1(n3478), .A2(n3477), .ZN(n3480) );
  XNOR2_X1 U3631 ( .A(n3434), .B(n3444), .ZN(n3784) );
  NAND2_X1 U3632 ( .A1(n3420), .A2(n3443), .ZN(n3434) );
  NAND2_X1 U3633 ( .A1(n3766), .A2(n3765), .ZN(n4394) );
  INV_X1 U3634 ( .A(n3170), .ZN(n3171) );
  INV_X1 U3635 ( .A(n3278), .ZN(n3276) );
  OR2_X1 U3636 ( .A1(n3199), .A2(n6421), .ZN(n3378) );
  INV_X1 U3637 ( .A(n3245), .ZN(n3246) );
  NOR2_X1 U3638 ( .A1(n3538), .A2(n3533), .ZN(n3567) );
  NAND2_X1 U3639 ( .A1(n3379), .A2(n3378), .ZN(n3548) );
  INV_X1 U3640 ( .A(n5857), .ZN(n5023) );
  AOI21_X1 U3641 ( .B1(n6430), .B2(n4557), .A(n5363), .ZN(n4606) );
  INV_X1 U3642 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6394) );
  AND2_X1 U3643 ( .A1(n3577), .A2(n3576), .ZN(n5395) );
  AND2_X1 U3644 ( .A1(n4239), .A2(n3724), .ZN(n5392) );
  AND2_X1 U3645 ( .A1(n3693), .A2(n3692), .ZN(n5465) );
  NAND2_X1 U3646 ( .A1(n5540), .A2(n5465), .ZN(n5464) );
  AND3_X1 U3647 ( .A1(n3915), .A2(n3914), .A3(n3913), .ZN(n5353) );
  NAND2_X1 U3648 ( .A1(n3220), .A2(n4391), .ZN(n4392) );
  AND2_X1 U3649 ( .A1(n4339), .A2(n4338), .ZN(n6088) );
  NOR2_X1 U3650 ( .A1(n4120), .A2(n5637), .ZN(n4121) );
  OR2_X1 U3651 ( .A1(n4086), .A2(n5869), .ZN(n4120) );
  NOR2_X1 U3652 ( .A1(n5474), .A2(n5537), .ZN(n5462) );
  AND2_X1 U3653 ( .A1(n4038), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4039)
         );
  OR2_X1 U3654 ( .A1(n5882), .A2(n4233), .ZN(n4056) );
  NAND2_X1 U3655 ( .A1(n3492), .A2(n2986), .ZN(n3042) );
  NAND2_X1 U3656 ( .A1(n3969), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4005)
         );
  INV_X1 U3657 ( .A(n5566), .ZN(n3987) );
  NAND2_X1 U3658 ( .A1(n3951), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3968)
         );
  OR2_X1 U3659 ( .A1(n3927), .A2(n3928), .ZN(n3936) );
  AND2_X1 U3660 ( .A1(n3880), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3881)
         );
  NAND2_X1 U3661 ( .A1(n3881), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3927)
         );
  NOR2_X1 U3662 ( .A1(n3866), .A2(n3865), .ZN(n3880) );
  NOR2_X1 U3663 ( .A1(n3834), .A2(n6018), .ZN(n3851) );
  INV_X1 U3664 ( .A(n3469), .ZN(n3038) );
  AND2_X1 U3665 ( .A1(n3797), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3818)
         );
  AOI21_X1 U3666 ( .B1(n3795), .B2(n3916), .A(n3794), .ZN(n4576) );
  CLKBUF_X1 U3667 ( .A(n4494), .Z(n4495) );
  INV_X1 U3668 ( .A(n3777), .ZN(n3778) );
  NAND2_X1 U3669 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3778), .ZN(n3790)
         );
  NOR2_X1 U3670 ( .A1(n6591), .A2(n6623), .ZN(n3768) );
  AND2_X1 U3671 ( .A1(n2968), .A2(n2991), .ZN(n2990) );
  NAND2_X1 U3672 ( .A1(n4260), .A2(n4259), .ZN(n4271) );
  NAND2_X1 U3673 ( .A1(n5540), .A2(n2983), .ZN(n5455) );
  NOR2_X1 U3674 ( .A1(n5551), .A2(n5480), .ZN(n5539) );
  AND2_X1 U3675 ( .A1(n3682), .A2(n3681), .ZN(n5549) );
  OR2_X1 U3676 ( .A1(n5548), .A2(n5549), .ZN(n5551) );
  AND2_X1 U3677 ( .A1(n5834), .A2(n3006), .ZN(n5556) );
  AND2_X1 U3678 ( .A1(n3007), .A2(n2964), .ZN(n3006) );
  INV_X1 U3679 ( .A(n3677), .ZN(n3007) );
  AND2_X1 U3680 ( .A1(n3668), .A2(n3667), .ZN(n5507) );
  AND2_X1 U3681 ( .A1(n5834), .A2(n5516), .ZN(n5518) );
  NAND2_X1 U3682 ( .A1(n3506), .A2(n2979), .ZN(n5696) );
  INV_X1 U3683 ( .A(n5719), .ZN(n3504) );
  NAND2_X1 U3684 ( .A1(n3003), .A2(n5287), .ZN(n3002) );
  INV_X1 U3685 ( .A(n3004), .ZN(n3003) );
  NOR3_X1 U3686 ( .A1(n6009), .A2(n5222), .A3(n3004), .ZN(n5286) );
  NAND2_X1 U3687 ( .A1(n5016), .A2(n3491), .ZN(n2989) );
  NOR2_X1 U3688 ( .A1(n4504), .A2(n4497), .ZN(n4581) );
  NAND2_X1 U3689 ( .A1(n6043), .A2(n4503), .ZN(n4504) );
  NAND2_X1 U3690 ( .A1(n6236), .A2(n4683), .ZN(n4688) );
  AND2_X1 U3691 ( .A1(n5270), .A2(n4364), .ZN(n4685) );
  AND2_X1 U3692 ( .A1(n3610), .A2(n3609), .ZN(n4361) );
  NAND2_X1 U3693 ( .A1(n3698), .A2(n3617), .ZN(n4359) );
  CLKBUF_X1 U3694 ( .A(n4417), .Z(n4418) );
  NAND2_X1 U3695 ( .A1(n3373), .A2(n3372), .ZN(n4410) );
  AND3_X1 U3696 ( .A1(n4408), .A2(n4407), .A3(n4406), .ZN(n4544) );
  NOR2_X1 U3697 ( .A1(n4765), .A2(n2963), .ZN(n4803) );
  NOR2_X1 U3698 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4606), .ZN(n4872) );
  AND2_X1 U3699 ( .A1(n5857), .A2(n4564), .ZN(n4825) );
  INV_X1 U3700 ( .A(n5098), .ZN(n6250) );
  AND2_X1 U3701 ( .A1(n5857), .A2(n4707), .ZN(n4955) );
  NAND2_X1 U3702 ( .A1(n5389), .A2(n5390), .ZN(n6518) );
  NAND2_X1 U3703 ( .A1(n5385), .A2(n5386), .ZN(n3013) );
  INV_X1 U3704 ( .A(n6046), .ZN(n6035) );
  OR2_X1 U3705 ( .A1(n5375), .A2(n4995), .ZN(n6016) );
  AND2_X1 U3706 ( .A1(n5378), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U3707 ( .A1(n4324), .A2(n6119), .ZN(n5581) );
  INV_X1 U3708 ( .A(n4460), .ZN(n6129) );
  OAI21_X1 U3709 ( .B1(n3335), .B2(n6520), .A(n4369), .ZN(n6130) );
  INV_X1 U3710 ( .A(n6119), .ZN(n6131) );
  INV_X1 U3711 ( .A(n6129), .ZN(n4480) );
  XNOR2_X1 U3712 ( .A(n4295), .B(n4294), .ZN(n4988) );
  INV_X1 U3713 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5678) );
  INV_X1 U3714 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5685) );
  INV_X1 U3715 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5703) );
  OR2_X1 U3716 ( .A1(n6420), .A2(n6425), .ZN(n6196) );
  NOR2_X1 U3717 ( .A1(n4588), .A2(n4587), .ZN(n4644) );
  INV_X1 U3718 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6623) );
  INV_X1 U3719 ( .A(n6170), .ZN(n5728) );
  OR2_X1 U3720 ( .A1(n4484), .A2(n4483), .ZN(n5152) );
  NAND2_X1 U3721 ( .A1(n6144), .A2(n4297), .ZN(n5725) );
  OR2_X1 U3722 ( .A1(n5427), .A2(n5426), .ZN(n5732) );
  NAND2_X1 U3723 ( .A1(n5611), .A2(n2968), .ZN(n5623) );
  AND2_X1 U3724 ( .A1(n5779), .A2(n3744), .ZN(n5758) );
  AND2_X1 U3725 ( .A1(n5776), .A2(n3738), .ZN(n5767) );
  OAI21_X1 U3726 ( .B1(n5677), .B2(n3023), .A(n3020), .ZN(n3032) );
  NAND2_X1 U3727 ( .A1(n3030), .A2(n3024), .ZN(n3018) );
  NAND2_X1 U3728 ( .A1(n3019), .A2(n3025), .ZN(n5665) );
  NAND2_X1 U3729 ( .A1(n5677), .A2(n3026), .ZN(n3019) );
  NAND2_X1 U3730 ( .A1(n5834), .A2(n2964), .ZN(n5560) );
  NAND2_X1 U3731 ( .A1(n5342), .A2(n6230), .ZN(n6179) );
  NAND2_X1 U3732 ( .A1(n5262), .A2(n5261), .ZN(n6135) );
  NAND2_X1 U3733 ( .A1(n3010), .A2(n3009), .ZN(n6044) );
  NAND2_X1 U3734 ( .A1(n4688), .A2(n4689), .ZN(n6230) );
  INV_X1 U3735 ( .A(n4684), .ZN(n6236) );
  AND2_X1 U3736 ( .A1(n3010), .A2(n3611), .ZN(n5198) );
  NOR2_X1 U3737 ( .A1(n5332), .A2(n4456), .ZN(n6244) );
  AND2_X1 U3738 ( .A1(n5346), .A2(n4431), .ZN(n4456) );
  NAND2_X1 U3739 ( .A1(n3725), .A2(n6389), .ZN(n5346) );
  INV_X1 U3740 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6388) );
  CLKBUF_X1 U3741 ( .A(n4437), .Z(n5854) );
  INV_X1 U3742 ( .A(n6310), .ZN(n6297) );
  INV_X1 U3743 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5362) );
  AND2_X1 U3744 ( .A1(n5396), .A2(n2958), .ZN(n6389) );
  AND2_X1 U3745 ( .A1(n5401), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5363) );
  INV_X1 U3746 ( .A(n5035), .ZN(n5058) );
  INV_X1 U3747 ( .A(n6291), .ZN(n4635) );
  INV_X1 U3748 ( .A(n6295), .ZN(n6346) );
  OR2_X1 U3749 ( .A1(n6251), .A2(n5098), .ZN(n6302) );
  OAI211_X1 U3750 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n5069), .A(n5227), .B(n4772), .ZN(n4795) );
  AND2_X1 U3751 ( .A1(n4825), .A2(n5098), .ZN(n4913) );
  NAND2_X1 U3752 ( .A1(n3072), .A2(n3220), .ZN(n4838) );
  INV_X1 U3753 ( .A(n4847), .ZN(n6304) );
  INV_X1 U3754 ( .A(n6315), .ZN(n6256) );
  INV_X1 U3755 ( .A(n6319), .ZN(n6359) );
  INV_X1 U3756 ( .A(n4857), .ZN(n6321) );
  INV_X1 U3757 ( .A(n6325), .ZN(n6270) );
  INV_X1 U3758 ( .A(n4828), .ZN(n6364) );
  INV_X1 U3759 ( .A(n6329), .ZN(n6365) );
  INV_X1 U3760 ( .A(n6335), .ZN(n6277) );
  INV_X1 U3761 ( .A(n4844), .ZN(n6372) );
  INV_X1 U3762 ( .A(n6339), .ZN(n6374) );
  INV_X1 U3763 ( .A(n4835), .ZN(n6341) );
  INV_X1 U3764 ( .A(n6345), .ZN(n6284) );
  AND2_X1 U3765 ( .A1(n4955), .A2(n5098), .ZN(n4977) );
  AND2_X1 U3766 ( .A1(n4955), .A2(n6250), .ZN(n5035) );
  INV_X1 U3767 ( .A(n6355), .ZN(n6290) );
  AND2_X1 U3768 ( .A1(n6412), .A2(n6411), .ZN(n6429) );
  INV_X1 U3769 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6421) );
  INV_X1 U3770 ( .A(n6524), .ZN(n6430) );
  INV_X1 U3771 ( .A(n6429), .ZN(n6507) );
  NAND2_X1 U3772 ( .A1(n3014), .A2(n3011), .ZN(U2796) );
  OR2_X1 U3773 ( .A1(n5529), .A2(n5988), .ZN(n3014) );
  AOI21_X1 U3774 ( .B1(n5388), .B2(n6038), .A(n3012), .ZN(n3011) );
  OR2_X1 U3775 ( .A1(n5387), .A2(n3013), .ZN(n3012) );
  AOI21_X1 U3776 ( .B1(n4256), .B2(n4255), .A(n4254), .ZN(n4257) );
  NOR2_X1 U3777 ( .A1(n4253), .A2(n6076), .ZN(n4254) );
  INV_X1 U3778 ( .A(n4314), .ZN(n4315) );
  OAI21_X1 U3779 ( .B1(n5587), .B2(n6139), .A(n4313), .ZN(n4314) );
  AND2_X1 U3780 ( .A1(n3746), .A2(n3745), .ZN(n3747) );
  AND2_X1 U3781 ( .A1(n4269), .A2(n4268), .ZN(n4270) );
  AND2_X1 U3782 ( .A1(n4284), .A2(n4283), .ZN(n4285) );
  AND2_X1 U3783 ( .A1(n2969), .A2(n2985), .ZN(n2964) );
  NAND2_X1 U3784 ( .A1(n2994), .A2(n2976), .ZN(n5690) );
  NAND2_X1 U3785 ( .A1(n5308), .A2(n5313), .ZN(n3055) );
  OR2_X1 U3786 ( .A1(n5488), .A2(n3059), .ZN(n2965) );
  OR2_X1 U3787 ( .A1(n5488), .A2(n5487), .ZN(n2966) );
  AND2_X1 U3788 ( .A1(n5315), .A2(n3056), .ZN(n5355) );
  OR2_X1 U3789 ( .A1(n5648), .A2(n6638), .ZN(n2967) );
  AND2_X1 U3790 ( .A1(n5648), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n2968)
         );
  AND2_X1 U3791 ( .A1(n5507), .A2(n5516), .ZN(n2969) );
  INV_X2 U3792 ( .A(n5544), .ZN(n6076) );
  AND2_X1 U3793 ( .A1(n3480), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n2970)
         );
  OR3_X1 U3794 ( .A1(n6009), .A2(n5222), .A3(n3002), .ZN(n2971) );
  NAND2_X1 U3795 ( .A1(n5462), .A2(n5463), .ZN(n5449) );
  NAND2_X1 U3796 ( .A1(n5315), .A2(n3053), .ZN(n5504) );
  AND2_X2 U3797 ( .A1(n4528), .A2(n4424), .ZN(n3182) );
  NAND2_X1 U3798 ( .A1(n3485), .A2(n3484), .ZN(n3496) );
  NOR2_X1 U3799 ( .A1(n5488), .A2(n3061), .ZN(n2972) );
  AND4_X1 U3800 ( .A1(n3143), .A2(n3142), .A3(n3141), .A4(n3140), .ZN(n2973)
         );
  NAND2_X1 U3801 ( .A1(n5648), .A2(n3495), .ZN(n2974) );
  NOR2_X1 U3802 ( .A1(n5423), .A2(n5424), .ZN(n4307) );
  NAND2_X1 U3803 ( .A1(n2994), .A2(n3503), .ZN(n5717) );
  NAND2_X1 U3804 ( .A1(n3030), .A2(n3028), .ZN(n2975) );
  AND2_X1 U3805 ( .A1(n3504), .A2(n3503), .ZN(n2976) );
  AND2_X1 U3806 ( .A1(n5648), .A2(n3502), .ZN(n2977) );
  INV_X1 U3807 ( .A(n3513), .ZN(n3514) );
  AND2_X1 U3808 ( .A1(n2974), .A2(n5261), .ZN(n2978) );
  NAND2_X1 U3809 ( .A1(n5648), .A2(n5934), .ZN(n2979) );
  NAND2_X1 U3810 ( .A1(n5834), .A2(n2969), .ZN(n5493) );
  NOR2_X1 U3811 ( .A1(n5138), .A2(n5218), .ZN(n5219) );
  NAND2_X1 U3812 ( .A1(n3049), .A2(n3051), .ZN(n4642) );
  NAND2_X1 U3813 ( .A1(n3850), .A2(n3849), .ZN(n5138) );
  NAND2_X1 U3814 ( .A1(n3493), .A2(n5182), .ZN(n5262) );
  NAND2_X1 U3815 ( .A1(n3501), .A2(n3500), .ZN(n5723) );
  AND2_X1 U3816 ( .A1(n3028), .A2(n5664), .ZN(n2980) );
  INV_X1 U3817 ( .A(n3864), .ZN(n5218) );
  INV_X1 U3818 ( .A(n3044), .ZN(n3043) );
  NAND2_X1 U3819 ( .A1(n2979), .A2(n3045), .ZN(n3044) );
  AND2_X1 U3820 ( .A1(n5282), .A2(n3864), .ZN(n2981) );
  AND2_X1 U3821 ( .A1(n3053), .A2(n3070), .ZN(n2982) );
  NAND2_X1 U3822 ( .A1(n3067), .A2(n3065), .ZN(n3064) );
  INV_X1 U3823 ( .A(n2967), .ZN(n3031) );
  INV_X1 U3824 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3048) );
  NOR2_X1 U3825 ( .A1(n5544), .A2(n4325), .ZN(n6073) );
  AND2_X1 U3826 ( .A1(n5465), .A2(n3017), .ZN(n2983) );
  INV_X1 U3827 ( .A(n5487), .ZN(n3062) );
  OR2_X1 U3828 ( .A1(n6009), .A2(n3004), .ZN(n2984) );
  INV_X1 U3829 ( .A(n3071), .ZN(n3056) );
  OR2_X1 U3830 ( .A1(n4452), .A2(n3709), .ZN(n3010) );
  NAND2_X1 U3831 ( .A1(n3670), .A2(n3669), .ZN(n2985) );
  INV_X1 U3832 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3000) );
  NAND2_X1 U3833 ( .A1(n4291), .A2(n6310), .ZN(n6139) );
  NAND3_X1 U3834 ( .A1(n5934), .A2(n5824), .A3(n5829), .ZN(n2986) );
  INV_X1 U3835 ( .A(n5735), .ZN(n2991) );
  AND2_X1 U3836 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n2987) );
  OAI33_X1 U3837 ( .A1(n4713), .A2(n6263), .A3(n5103), .B1(n6252), .B2(n6297), 
        .B3(n6052), .ZN(n2988) );
  INV_X1 U3838 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6263) );
  INV_X1 U3839 ( .A(n2961), .ZN(n6052) );
  NOR2_X4 U3840 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4528) );
  AND2_X2 U3841 ( .A1(n4439), .A2(n4528), .ZN(n3173) );
  NOR2_X4 U3842 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4439) );
  NAND2_X1 U3843 ( .A1(n2989), .A2(n5181), .ZN(n3493) );
  XNOR2_X1 U3844 ( .A(n2989), .B(n5183), .ZN(n6190) );
  NAND2_X1 U3845 ( .A1(n3501), .A2(n2995), .ZN(n2994) );
  XNOR2_X2 U3846 ( .A(n3332), .B(n3331), .ZN(n3370) );
  AOI21_X2 U3847 ( .B1(n5684), .B2(n3510), .A(n3509), .ZN(n5640) );
  NAND2_X1 U3848 ( .A1(n3001), .A2(n5496), .ZN(n3669) );
  NAND2_X1 U3849 ( .A1(n3001), .A2(n5534), .ZN(n3696) );
  NAND2_X1 U3850 ( .A1(n3001), .A2(n5532), .ZN(n3701) );
  NAND2_X1 U3851 ( .A1(n3001), .A2(n6075), .ZN(n3613) );
  NAND2_X1 U3852 ( .A1(n3001), .A2(n3620), .ZN(n3623) );
  NAND2_X1 U3853 ( .A1(n3001), .A2(n6537), .ZN(n3629) );
  NAND2_X1 U3854 ( .A1(n3001), .A2(n5191), .ZN(n3637) );
  NAND2_X1 U3855 ( .A1(n3001), .A2(n3642), .ZN(n3645) );
  NAND2_X1 U3856 ( .A1(n3001), .A2(n3648), .ZN(n3651) );
  NAND2_X1 U3857 ( .A1(n3001), .A2(n3655), .ZN(n3659) );
  NAND2_X1 U3858 ( .A1(n3001), .A2(n5552), .ZN(n3681) );
  NOR2_X1 U3859 ( .A1(n6009), .A2(n6010), .ZN(n6011) );
  INV_X1 U3860 ( .A(n5142), .ZN(n3005) );
  NAND2_X1 U3861 ( .A1(n3030), .A2(n2980), .ZN(n5655) );
  AND2_X1 U3862 ( .A1(n3030), .A2(n2967), .ZN(n5670) );
  NAND2_X1 U3863 ( .A1(n3032), .A2(n3018), .ZN(n5649) );
  OAI21_X1 U3864 ( .B1(n3034), .B2(n6145), .A(n3033), .ZN(n5018) );
  AOI21_X1 U3865 ( .B1(n4697), .B2(n3038), .A(n2970), .ZN(n3033) );
  INV_X1 U3866 ( .A(n4697), .ZN(n3034) );
  NAND2_X1 U3867 ( .A1(n3037), .A2(n3035), .ZN(n5016) );
  NAND2_X1 U3868 ( .A1(n4698), .A2(n4697), .ZN(n4696) );
  NAND2_X1 U3869 ( .A1(n6145), .A2(n3469), .ZN(n4698) );
  NAND2_X1 U3870 ( .A1(n3221), .A2(n3220), .ZN(n3582) );
  NAND3_X1 U3871 ( .A1(n3201), .A2(n3206), .A3(n4993), .ZN(n4331) );
  NAND2_X1 U3872 ( .A1(n5262), .A2(n2978), .ZN(n3499) );
  OAI21_X1 U3873 ( .B1(n3506), .B2(n3041), .A(n3039), .ZN(n5654) );
  NAND2_X1 U3874 ( .A1(n3046), .A2(n3223), .ZN(n3308) );
  NAND2_X1 U3875 ( .A1(n3047), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3046) );
  NAND4_X1 U3876 ( .A1(n3240), .A2(n3239), .A3(n3212), .A4(n3243), .ZN(n3047)
         );
  NAND2_X1 U3877 ( .A1(n3217), .A2(n4332), .ZN(n3240) );
  AND2_X2 U3878 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4424) );
  AND2_X2 U3879 ( .A1(n4530), .A2(n4424), .ZN(n3172) );
  NOR2_X1 U3880 ( .A1(n4587), .A2(n3050), .ZN(n3049) );
  NAND2_X1 U3881 ( .A1(n3850), .A2(n3052), .ZN(n3887) );
  NAND2_X1 U3882 ( .A1(n3887), .A2(n3886), .ZN(n3888) );
  NAND2_X1 U3883 ( .A1(n3055), .A2(n2982), .ZN(n5505) );
  OR2_X2 U3884 ( .A1(n5488), .A2(n3057), .ZN(n5475) );
  INV_X1 U3885 ( .A(n5474), .ZN(n3066) );
  NOR2_X1 U3886 ( .A1(n5474), .A2(n3064), .ZN(n5436) );
  XNOR2_X1 U3887 ( .A(n4263), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5610)
         );
  NAND2_X1 U3888 ( .A1(n4262), .A2(n4261), .ZN(n4263) );
  XNOR2_X1 U3889 ( .A(n4290), .B(n4289), .ZN(n5388) );
  NAND2_X2 U3890 ( .A1(n3587), .A2(n5402), .ZN(n3598) );
  NAND2_X1 U3891 ( .A1(n5388), .A2(n4326), .ZN(n4329) );
  NAND2_X1 U3892 ( .A1(n3338), .A2(n3337), .ZN(n6163) );
  CLKBUF_X1 U3893 ( .A(n5505), .Z(n5567) );
  NOR2_X2 U3894 ( .A1(n4234), .A2(n4235), .ZN(n4290) );
  NAND2_X1 U3895 ( .A1(n4307), .A2(n4309), .ZN(n4234) );
  CLKBUF_X1 U3896 ( .A(n4562), .Z(n5857) );
  AOI21_X1 U3897 ( .B1(n3211), .B2(n3210), .A(n3714), .ZN(n3212) );
  NOR2_X1 U3898 ( .A1(n3714), .A2(n3199), .ZN(n3201) );
  AND2_X1 U3899 ( .A1(n3967), .A2(n3966), .ZN(n3070) );
  NAND2_X1 U3900 ( .A1(n3934), .A2(n5314), .ZN(n3071) );
  NOR3_X2 U3901 ( .A1(n6508), .A2(STATE2_REG_0__SCAN_IN), .A3(n4606), .ZN(
        n3072) );
  AND2_X1 U3902 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3073) );
  INV_X1 U3903 ( .A(n5578), .ZN(n4255) );
  AND3_X1 U3904 ( .A1(n4259), .A2(n4266), .A3(n4282), .ZN(n3074) );
  INV_X1 U3905 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3928) );
  INV_X1 U3906 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6614) );
  INV_X1 U3907 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U3908 ( .A1(n5648), .A2(n5612), .ZN(n3511) );
  AOI21_X1 U3909 ( .B1(n6388), .B2(STATE2_REG_3__SCAN_IN), .A(n4911), .ZN(
        n6309) );
  INV_X1 U3910 ( .A(n6309), .ZN(n5065) );
  INV_X1 U3911 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3526) );
  NOR2_X1 U3912 ( .A1(n6253), .A2(n4871), .ZN(n3075) );
  OAI21_X1 U3913 ( .B1(n5301), .B2(n5297), .A(n5298), .ZN(n5337) );
  AND4_X1 U3914 ( .A1(n3239), .A2(n3238), .A3(n3237), .A4(n4538), .ZN(n3077)
         );
  AOI21_X1 U3915 ( .B1(n3536), .B2(n4607), .A(n5402), .ZN(n3545) );
  AND2_X1 U3916 ( .A1(n6388), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3540)
         );
  INV_X1 U3917 ( .A(n3443), .ZN(n3446) );
  NOR2_X1 U3918 ( .A1(n3446), .A2(n3445), .ZN(n3447) );
  OR2_X1 U3919 ( .A1(n3431), .A2(n3430), .ZN(n3461) );
  NAND2_X1 U3920 ( .A1(n3525), .A2(n3524), .ZN(n3530) );
  OR2_X1 U3921 ( .A1(n3326), .A2(n3325), .ZN(n3334) );
  OR2_X1 U3922 ( .A1(n3457), .A2(n3456), .ZN(n3474) );
  INV_X1 U3923 ( .A(n3241), .ZN(n3483) );
  AOI21_X1 U3924 ( .B1(n3530), .B2(n3529), .A(n3527), .ZN(n3532) );
  NAND3_X1 U3925 ( .A1(n3199), .A2(n4993), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3538) );
  INV_X1 U3926 ( .A(n5140), .ZN(n3849) );
  OR2_X1 U3927 ( .A1(n4105), .A2(n4104), .ZN(n4125) );
  OR2_X1 U3928 ( .A1(n4438), .A2(n6421), .ZN(n4230) );
  INV_X1 U3929 ( .A(n3481), .ZN(n3486) );
  OR2_X1 U3930 ( .A1(n3296), .A2(n3295), .ZN(n3360) );
  AND2_X1 U3931 ( .A1(n4161), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4162)
         );
  INV_X1 U3932 ( .A(n5476), .ZN(n4083) );
  NAND2_X1 U3933 ( .A1(n3753), .A2(n4559), .ZN(n3754) );
  OR2_X1 U3934 ( .A1(n4085), .A2(n5658), .ZN(n4086) );
  INV_X1 U3935 ( .A(n4233), .ZN(n3792) );
  INV_X1 U3936 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3935) );
  INV_X1 U3937 ( .A(n2957), .ZN(n3533) );
  NAND2_X1 U3938 ( .A1(n3377), .A2(n3376), .ZN(n4603) );
  NAND2_X1 U3939 ( .A1(n3342), .A2(n3341), .ZN(n3343) );
  NAND2_X1 U3940 ( .A1(n3316), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3105) );
  OR2_X1 U3941 ( .A1(n6420), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4296) );
  NAND2_X1 U3942 ( .A1(n4162), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4206)
         );
  OR2_X1 U3943 ( .A1(n4005), .A2(n5685), .ZN(n4006) );
  NOR2_X1 U3944 ( .A1(n3968), .A2(n5703), .ZN(n3969) );
  OR2_X1 U3945 ( .A1(n4293), .A2(n4292), .ZN(n4295) );
  OR2_X1 U3946 ( .A1(n5375), .A2(n4999), .ZN(n5988) );
  INV_X1 U3947 ( .A(n4998), .ZN(n3709) );
  AND3_X1 U3948 ( .A1(n3680), .A2(n3679), .A3(n3678), .ZN(n5555) );
  NAND2_X1 U3949 ( .A1(n4408), .A2(n4244), .ZN(n4245) );
  AND2_X1 U3950 ( .A1(n4337), .A2(n6408), .ZN(n4338) );
  NAND2_X1 U3951 ( .A1(n4121), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4160)
         );
  NOR2_X1 U3952 ( .A1(n3936), .A2(n3935), .ZN(n3951) );
  NAND2_X1 U3953 ( .A1(n3818), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3834)
         );
  INV_X1 U3954 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6591) );
  OR2_X1 U3955 ( .A1(n4271), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4261)
         );
  AND2_X1 U3956 ( .A1(n5648), .A2(n6549), .ZN(n5647) );
  NAND2_X1 U3957 ( .A1(n3725), .A2(n5392), .ZN(n4684) );
  NAND2_X1 U3958 ( .A1(n3592), .A2(n6422), .ZN(n3729) );
  INV_X1 U3959 ( .A(n3767), .ZN(n5025) );
  AND2_X1 U3960 ( .A1(n5857), .A2(n4602), .ZN(n4608) );
  INV_X1 U3961 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5030) );
  INV_X1 U3962 ( .A(n4913), .ZN(n4939) );
  AND2_X1 U3963 ( .A1(n5362), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3591) );
  NOR2_X1 U3964 ( .A1(n5889), .A2(n5372), .ZN(n5878) );
  NOR2_X1 U3965 ( .A1(n4006), .A2(n5678), .ZN(n4038) );
  INV_X1 U3966 ( .A(n6029), .ZN(n6048) );
  INV_X1 U3967 ( .A(n6033), .ZN(n6020) );
  INV_X1 U3968 ( .A(n5988), .ZN(n6047) );
  AND2_X1 U3969 ( .A1(n4988), .A2(n4987), .ZN(n6057) );
  NOR2_X1 U3970 ( .A1(n4279), .A2(n4278), .ZN(n5530) );
  NAND2_X1 U3971 ( .A1(n4245), .A2(n6422), .ZN(n5544) );
  OAI21_X1 U3972 ( .B1(n4401), .B2(n4323), .A(n6422), .ZN(n4324) );
  NOR2_X1 U3973 ( .A1(n4557), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4517) );
  AND2_X1 U3974 ( .A1(n5401), .A2(n6422), .ZN(n4337) );
  AND2_X1 U3975 ( .A1(n5308), .A2(n5311), .ZN(n5994) );
  NOR2_X1 U3976 ( .A1(n3790), .A2(n3789), .ZN(n3797) );
  NAND2_X1 U3977 ( .A1(n3768), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3777)
         );
  AND2_X1 U3978 ( .A1(n5784), .A2(n5786), .ZN(n5779) );
  NOR2_X1 U3979 ( .A1(n5933), .A2(n3743), .ZN(n5784) );
  AND2_X1 U3980 ( .A1(n5571), .A2(n5570), .ZN(n5972) );
  INV_X1 U3981 ( .A(n6184), .ZN(n6242) );
  INV_X1 U3982 ( .A(n3729), .ZN(n3725) );
  INV_X1 U3983 ( .A(n4872), .ZN(n4911) );
  OAI21_X1 U3984 ( .B1(n5064), .B2(n5034), .A(n5033), .ZN(n5057) );
  OAI21_X1 U3985 ( .B1(n4654), .B2(n4653), .A(n4652), .ZN(n4677) );
  OAI21_X1 U3986 ( .B1(n4612), .B2(n4611), .A(n4610), .ZN(n4638) );
  AND2_X1 U3987 ( .A1(n4608), .A2(n6250), .ZN(n6291) );
  INV_X1 U3988 ( .A(n6302), .ZN(n6350) );
  OR2_X1 U3989 ( .A1(n5105), .A2(n5104), .ZN(n5134) );
  INV_X1 U3990 ( .A(n4773), .ZN(n4867) );
  AND2_X1 U3991 ( .A1(n4741), .A2(n2961), .ZN(n4768) );
  INV_X1 U3992 ( .A(n4946), .ZN(n6369) );
  NAND2_X1 U3993 ( .A1(n3767), .A2(n5023), .ZN(n4765) );
  AND2_X1 U3994 ( .A1(n4825), .A2(n6250), .ZN(n4853) );
  INV_X1 U3995 ( .A(n4850), .ZN(n6358) );
  INV_X1 U3996 ( .A(n4841), .ZN(n6331) );
  INV_X1 U3997 ( .A(n4838), .ZN(n6349) );
  AND2_X1 U3998 ( .A1(n3591), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6422) );
  NAND2_X1 U3999 ( .A1(n5403), .A2(n4337), .ZN(n5390) );
  INV_X1 U4000 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6424) );
  OR2_X1 U4001 ( .A1(n5375), .A2(n4992), .ZN(n6029) );
  AOI21_X1 U4002 ( .B1(n5402), .B2(n5144), .A(n6038), .ZN(n6053) );
  INV_X1 U4003 ( .A(n6073), .ZN(n5579) );
  INV_X1 U4004 ( .A(n5994), .ZN(n5331) );
  INV_X1 U4005 ( .A(n5357), .ZN(n4705) );
  INV_X1 U4006 ( .A(n6088), .ZN(n6115) );
  NAND3_X1 U4007 ( .A1(n4403), .A2(n4337), .A3(n6520), .ZN(n6119) );
  OR2_X1 U4008 ( .A1(n5390), .A2(n2958), .ZN(n4460) );
  AOI21_X1 U4009 ( .B1(n5608), .B2(n5681), .A(n5607), .ZN(n5609) );
  OAI21_X1 U4010 ( .B1(n3062), .B2(n5489), .A(n2966), .ZN(n5921) );
  NAND2_X1 U4011 ( .A1(n5725), .A2(n4300), .ZN(n6170) );
  OR2_X1 U4012 ( .A1(n6179), .A2(n3742), .ZN(n5933) );
  NAND2_X1 U4013 ( .A1(n3725), .A2(n3600), .ZN(n6184) );
  NAND2_X1 U4014 ( .A1(n5026), .A2(n5098), .ZN(n5092) );
  INV_X1 U4015 ( .A(n5229), .ZN(n5260) );
  AOI22_X1 U4016 ( .A1(n4651), .A2(n4653), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4650), .ZN(n4682) );
  OR2_X1 U4017 ( .A1(n4655), .A2(n5098), .ZN(n4906) );
  OR2_X1 U4018 ( .A1(n6251), .A2(n6250), .ZN(n6295) );
  NAND2_X1 U4019 ( .A1(n4803), .A2(n5098), .ZN(n5137) );
  OR2_X1 U4020 ( .A1(n4765), .A2(n4747), .ZN(n6378) );
  OR2_X1 U4021 ( .A1(n4765), .A2(n4748), .ZN(n4946) );
  INV_X1 U4022 ( .A(n4711), .ZN(n4740) );
  INV_X1 U4023 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6508) );
  INV_X1 U4024 ( .A(READY_N), .ZN(n6520) );
  INV_X1 U4025 ( .A(n6495), .ZN(n6494) );
  NAND2_X1 U4026 ( .A1(n4258), .A2(n4257), .ZN(U2829) );
  AND2_X2 U4027 ( .A1(n4444), .A2(n4528), .ZN(n3174) );
  AND2_X4 U4028 ( .A1(n5367), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4447)
         );
  AOI22_X1 U4029 ( .A1(n3174), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3082) );
  INV_X1 U4030 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3078) );
  AND2_X4 U4031 ( .A1(n3083), .A2(n4444), .ZN(n3819) );
  AOI22_X1 U4032 ( .A1(n3819), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3081) );
  AND2_X2 U4033 ( .A1(n4530), .A2(n4439), .ZN(n3266) );
  AND2_X2 U4034 ( .A1(n3083), .A2(n4424), .ZN(n3267) );
  AOI22_X1 U4035 ( .A1(n3266), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3080) );
  AND2_X2 U4036 ( .A1(n4548), .A2(n4424), .ZN(n3184) );
  AOI22_X1 U4037 ( .A1(n3181), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3079) );
  AND2_X2 U4038 ( .A1(n4530), .A2(n4447), .ZN(n3180) );
  AOI22_X1 U4039 ( .A1(n3183), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3087) );
  AND2_X2 U4040 ( .A1(n4444), .A2(n4548), .ZN(n3247) );
  AOI22_X1 U4041 ( .A1(n3247), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3086) );
  AND2_X2 U4042 ( .A1(n4447), .A2(n4548), .ZN(n3284) );
  AOI22_X1 U4043 ( .A1(n3284), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3085) );
  AOI22_X1 U4044 ( .A1(n2959), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3084) );
  NAND2_X2 U4045 ( .A1(n3089), .A2(n3088), .ZN(n3218) );
  AOI22_X1 U4046 ( .A1(n3819), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3093) );
  AOI22_X1 U4047 ( .A1(n3180), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3092) );
  AOI22_X1 U4048 ( .A1(n3316), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3091) );
  AOI22_X1 U4049 ( .A1(n3284), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3090) );
  NAND4_X1 U4050 ( .A1(n3093), .A2(n3092), .A3(n3091), .A4(n3090), .ZN(n3099)
         );
  AOI22_X1 U4051 ( .A1(n3247), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3097) );
  AOI22_X1 U4052 ( .A1(n3174), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3096) );
  AOI22_X1 U4053 ( .A1(n3266), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3181), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3095) );
  AOI22_X1 U4054 ( .A1(n3183), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3094) );
  NAND4_X1 U4055 ( .A1(n3097), .A2(n3096), .A3(n3095), .A4(n3094), .ZN(n3098)
         );
  NOR2_X1 U4056 ( .A1(n4607), .A2(n3219), .ZN(n3149) );
  NAND2_X1 U4057 ( .A1(n3819), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3103) );
  NAND2_X1 U4058 ( .A1(n3247), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3102)
         );
  NAND2_X1 U4059 ( .A1(n3266), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3101) );
  NAND2_X1 U4060 ( .A1(n3172), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3100)
         );
  NAND2_X1 U4061 ( .A1(n4106), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3107) );
  NAND2_X1 U4062 ( .A1(n3174), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3106) );
  NAND2_X1 U4063 ( .A1(n3173), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3104) );
  NAND2_X1 U4064 ( .A1(n3180), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3111)
         );
  NAND2_X1 U4065 ( .A1(n3179), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3110) );
  NAND2_X1 U4066 ( .A1(n3267), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3109) );
  NAND2_X1 U4067 ( .A1(n3181), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3108)
         );
  AND4_X1 U4068 ( .A1(n3111), .A2(n3110), .A3(n3109), .A4(n3108), .ZN(n3117)
         );
  NAND2_X1 U4069 ( .A1(n3183), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3115) );
  NAND2_X1 U4070 ( .A1(n3284), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3114)
         );
  NAND2_X1 U4071 ( .A1(n3182), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3113) );
  NAND2_X1 U4072 ( .A1(n3184), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3112)
         );
  AND4_X1 U4073 ( .A1(n3115), .A2(n3114), .A3(n3113), .A4(n3112), .ZN(n3116)
         );
  NAND4_X4 U4074 ( .A1(n3119), .A2(n3118), .A3(n3117), .A4(n3116), .ZN(n4993)
         );
  NAND2_X1 U4075 ( .A1(n3174), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3123) );
  NAND2_X1 U4076 ( .A1(n3819), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3122) );
  NAND2_X1 U4077 ( .A1(n3247), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3121)
         );
  NAND2_X1 U4078 ( .A1(n2959), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3120) );
  NAND2_X1 U4079 ( .A1(n3183), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3127) );
  NAND2_X1 U4080 ( .A1(n3172), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3126)
         );
  NAND2_X1 U4081 ( .A1(n3267), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3125) );
  NAND2_X1 U4082 ( .A1(n3184), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3124)
         );
  NAND2_X1 U4083 ( .A1(n3266), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3131) );
  NAND2_X1 U4084 ( .A1(n3179), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3130) );
  NAND2_X1 U4085 ( .A1(n2962), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3129) );
  NAND2_X1 U4086 ( .A1(n3173), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3128) );
  NAND2_X1 U4087 ( .A1(n3180), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3135)
         );
  NAND2_X1 U4088 ( .A1(n3284), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3134)
         );
  NAND2_X1 U4089 ( .A1(n3181), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3133)
         );
  NAND2_X1 U4090 ( .A1(n3182), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3132) );
  AOI22_X1 U4091 ( .A1(n3819), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3143) );
  AOI22_X1 U4092 ( .A1(n3266), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3142) );
  AOI22_X1 U4093 ( .A1(n3174), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n2959), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3141) );
  AOI22_X1 U4094 ( .A1(n2962), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3140) );
  INV_X1 U4095 ( .A(n3180), .ZN(n3252) );
  AOI22_X1 U4096 ( .A1(n3267), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3181), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3146) );
  AOI22_X1 U4097 ( .A1(n3183), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3145) );
  NAND3_X1 U4098 ( .A1(n3149), .A2(n3198), .A3(n3712), .ZN(n3601) );
  AOI22_X1 U4099 ( .A1(n3819), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3153) );
  AOI22_X1 U4100 ( .A1(n3266), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3152) );
  AOI22_X1 U4101 ( .A1(n2962), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U4102 ( .A1(n3174), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n2959), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3150) );
  AOI22_X1 U4103 ( .A1(n3180), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3157) );
  AOI22_X1 U4104 ( .A1(n3267), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3181), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3156) );
  AOI22_X1 U4105 ( .A1(n3183), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3155) );
  AOI22_X1 U4106 ( .A1(n3284), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3154) );
  NAND2_X2 U4107 ( .A1(n3159), .A2(n3158), .ZN(n3192) );
  AOI22_X1 U4108 ( .A1(n3819), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3163) );
  AOI22_X1 U4109 ( .A1(n3266), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3162) );
  AOI22_X1 U4110 ( .A1(n3174), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3161) );
  AOI22_X1 U4111 ( .A1(n4106), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3160) );
  NAND4_X1 U4112 ( .A1(n3163), .A2(n3162), .A3(n3161), .A4(n3160), .ZN(n3169)
         );
  AOI22_X1 U4113 ( .A1(n3180), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3167) );
  AOI22_X1 U4114 ( .A1(n3267), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3181), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3166) );
  AOI22_X1 U4115 ( .A1(n3183), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3165) );
  AOI22_X1 U4116 ( .A1(n3284), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3164) );
  NAND4_X1 U4117 ( .A1(n3167), .A2(n3166), .A3(n3165), .A4(n3164), .ZN(n3168)
         );
  INV_X1 U4118 ( .A(n4327), .ZN(n3520) );
  NOR2_X2 U4119 ( .A1(n3192), .A2(n3171), .ZN(n3753) );
  INV_X1 U4120 ( .A(n3753), .ZN(n3191) );
  AOI22_X1 U4121 ( .A1(n3819), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3178) );
  AOI22_X1 U4122 ( .A1(n3266), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3172), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3177) );
  AOI22_X1 U4123 ( .A1(n4106), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3176) );
  AOI22_X1 U4124 ( .A1(n3174), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3175) );
  AOI22_X1 U4125 ( .A1(n3180), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3188) );
  AOI22_X1 U4126 ( .A1(n3267), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3181), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3187) );
  AOI22_X1 U4127 ( .A1(n3183), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3186) );
  AOI22_X1 U4128 ( .A1(n3284), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3185) );
  NAND2_X2 U4129 ( .A1(n3190), .A2(n3189), .ZN(n3199) );
  AOI21_X2 U4130 ( .B1(n3192), .B2(n3210), .A(n3199), .ZN(n3221) );
  NAND2_X1 U4131 ( .A1(n3191), .A2(n3221), .ZN(n3213) );
  INV_X1 U4132 ( .A(n3213), .ZN(n3197) );
  AOI21_X2 U4133 ( .B1(n4391), .B2(n3219), .A(n4325), .ZN(n3215) );
  NAND2_X1 U4134 ( .A1(n3192), .A2(n3218), .ZN(n3195) );
  NAND2_X1 U4135 ( .A1(n4240), .A2(n3193), .ZN(n3194) );
  NAND2_X1 U4136 ( .A1(n3195), .A2(n3194), .ZN(n3196) );
  NAND2_X1 U4137 ( .A1(n3196), .A2(n3712), .ZN(n3214) );
  NAND2_X1 U4138 ( .A1(n3596), .A2(n3598), .ZN(n3204) );
  NAND2_X1 U4139 ( .A1(n3753), .A2(n3199), .ZN(n3235) );
  NAND2_X1 U4140 ( .A1(n3753), .A2(n3210), .ZN(n3200) );
  NAND2_X1 U4141 ( .A1(n3235), .A2(n3200), .ZN(n3206) );
  NAND2_X1 U4142 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6434) );
  OAI21_X1 U4143 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6434), .ZN(n3519) );
  INV_X1 U4144 ( .A(n3519), .ZN(n3202) );
  NOR2_X1 U4145 ( .A1(n2958), .A2(n3202), .ZN(n3209) );
  NAND2_X1 U4146 ( .A1(n6508), .A2(n5362), .ZN(n6420) );
  XNOR2_X1 U4147 ( .A(n6388), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6253)
         );
  INV_X1 U4148 ( .A(n3591), .ZN(n3312) );
  AND2_X1 U4149 ( .A1(n3312), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3205)
         );
  AOI21_X1 U4150 ( .B1(n3313), .B2(n6253), .A(n3205), .ZN(n3226) );
  INV_X1 U4151 ( .A(n3206), .ZN(n3208) );
  NAND2_X1 U4152 ( .A1(n4327), .A2(n4607), .ZN(n3207) );
  NAND2_X1 U4153 ( .A1(n3208), .A2(n3207), .ZN(n3243) );
  INV_X1 U4154 ( .A(n3209), .ZN(n3211) );
  NAND2_X1 U4155 ( .A1(n3213), .A2(n4621), .ZN(n3216) );
  NAND4_X1 U4156 ( .A1(n3216), .A2(n3215), .A3(n3214), .A4(n3536), .ZN(n3217)
         );
  NAND2_X1 U4157 ( .A1(n3241), .A2(n3219), .ZN(n4420) );
  INV_X2 U4158 ( .A(n2958), .ZN(n3536) );
  AND2_X4 U4159 ( .A1(n3536), .A2(n4993), .ZN(n3335) );
  NAND2_X1 U4160 ( .A1(n3582), .A2(n3335), .ZN(n3222) );
  NAND2_X1 U4161 ( .A1(n4391), .A2(n3559), .ZN(n3223) );
  NAND2_X1 U4162 ( .A1(n3308), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3224) );
  NAND2_X1 U4163 ( .A1(n3225), .A2(n3224), .ZN(n3305) );
  INV_X1 U4164 ( .A(n3226), .ZN(n3227) );
  NOR2_X1 U4165 ( .A1(n3227), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3228)
         );
  NAND2_X1 U4166 ( .A1(n3305), .A2(n3230), .ZN(n3306) );
  NAND2_X1 U4167 ( .A1(n3308), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3233) );
  MUX2_X1 U4168 ( .A(n3312), .B(n3313), .S(n6388), .Z(n3231) );
  INV_X1 U4169 ( .A(n3231), .ZN(n3232) );
  NAND2_X1 U4170 ( .A1(n3233), .A2(n3232), .ZN(n3283) );
  INV_X1 U4171 ( .A(n4391), .ZN(n3583) );
  OR2_X1 U4172 ( .A1(n6420), .A2(n6421), .ZN(n3234) );
  AOI21_X1 U4173 ( .B1(n3583), .B2(n3335), .A(n3234), .ZN(n3238) );
  NAND2_X1 U4174 ( .A1(n3714), .A2(n4993), .ZN(n3237) );
  INV_X1 U4175 ( .A(n3235), .ZN(n3581) );
  NOR2_X1 U4176 ( .A1(n4621), .A2(n3219), .ZN(n3236) );
  NAND2_X1 U4177 ( .A1(n3581), .A2(n3236), .ZN(n4538) );
  INV_X1 U4178 ( .A(n3240), .ZN(n3242) );
  NAND2_X1 U4179 ( .A1(n3242), .A2(n3483), .ZN(n3719) );
  INV_X1 U4180 ( .A(n3219), .ZN(n3605) );
  AOI21_X1 U4181 ( .B1(n4391), .B2(n3199), .A(n3605), .ZN(n3244) );
  AOI21_X1 U4182 ( .B1(n3243), .B2(n3244), .A(n3536), .ZN(n3245) );
  NAND3_X1 U4183 ( .A1(n3077), .A2(n3719), .A3(n3246), .ZN(n3281) );
  XNOR2_X1 U4184 ( .A(n3306), .B(n3304), .ZN(n4437) );
  INV_X1 U4185 ( .A(n3378), .ZN(n3327) );
  AOI22_X1 U4186 ( .A1(n4215), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3251) );
  AOI22_X1 U4187 ( .A1(n3174), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3250) );
  AOI22_X1 U4188 ( .A1(n3183), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4532), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3249) );
  AOI22_X1 U4189 ( .A1(n3803), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3248) );
  NAND4_X1 U4190 ( .A1(n3251), .A2(n3250), .A3(n3249), .A4(n3248), .ZN(n3259)
         );
  AOI22_X1 U4191 ( .A1(n4174), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3257) );
  INV_X2 U4192 ( .A(n3252), .ZN(n3425) );
  AOI22_X1 U4193 ( .A1(n3425), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3256) );
  AOI22_X1 U4194 ( .A1(n3819), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3255) );
  INV_X1 U4195 ( .A(n3181), .ZN(n4169) );
  AOI22_X1 U4196 ( .A1(n3289), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3254) );
  NAND4_X1 U4197 ( .A1(n3257), .A2(n3256), .A3(n3255), .A4(n3254), .ZN(n3258)
         );
  NAND2_X1 U4198 ( .A1(n3327), .A2(n3359), .ZN(n3260) );
  OAI21_X2 U4199 ( .B1(n4437), .B2(STATE2_REG_0__SCAN_IN), .A(n3260), .ZN(
        n3279) );
  INV_X1 U4200 ( .A(n3279), .ZN(n3277) );
  AOI22_X1 U4201 ( .A1(n3174), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3265) );
  AOI22_X1 U4202 ( .A1(n4173), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3264) );
  AOI22_X1 U4203 ( .A1(n4215), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3316), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U4204 ( .A1(n3289), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3262) );
  NAND4_X1 U4205 ( .A1(n3265), .A2(n3264), .A3(n3263), .A4(n3262), .ZN(n3273)
         );
  AOI22_X1 U4206 ( .A1(n3266), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3271) );
  AOI22_X1 U4207 ( .A1(n4195), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4532), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3270) );
  AOI22_X1 U4208 ( .A1(n3819), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3269) );
  AOI22_X1 U4209 ( .A1(n3803), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3268) );
  NAND4_X1 U4210 ( .A1(n3271), .A2(n3270), .A3(n3269), .A4(n3268), .ZN(n3272)
         );
  NAND2_X1 U4211 ( .A1(n3559), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3275) );
  INV_X1 U4212 ( .A(n3379), .ZN(n3330) );
  NAND2_X1 U4213 ( .A1(n3330), .A2(n3359), .ZN(n3274) );
  OAI211_X1 U4214 ( .C1(n3378), .C2(n3481), .A(n3275), .B(n3274), .ZN(n3278)
         );
  NAND2_X1 U4215 ( .A1(n3277), .A2(n3276), .ZN(n3303) );
  NAND2_X1 U4216 ( .A1(n3279), .A2(n3278), .ZN(n3280) );
  AND2_X2 U4217 ( .A1(n3303), .A2(n3280), .ZN(n3353) );
  INV_X1 U4218 ( .A(n3281), .ZN(n3282) );
  XNOR2_X2 U4219 ( .A(n3283), .B(n3282), .ZN(n5361) );
  NAND2_X1 U4220 ( .A1(n5361), .A2(n6421), .ZN(n3298) );
  AOI22_X1 U4221 ( .A1(n3174), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3288) );
  AOI22_X1 U4222 ( .A1(n4174), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4223 ( .A1(n3253), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3803), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4224 ( .A1(n4215), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3285) );
  NAND4_X1 U4225 ( .A1(n3288), .A2(n3287), .A3(n3286), .A4(n3285), .ZN(n3296)
         );
  AOI22_X1 U4226 ( .A1(n3819), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n2959), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3294) );
  AOI22_X1 U4227 ( .A1(n3425), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3267), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3293) );
  AOI22_X1 U4228 ( .A1(n3183), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U4229 ( .A1(n3290), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3291) );
  NAND4_X1 U4230 ( .A1(n3294), .A2(n3293), .A3(n3292), .A4(n3291), .ZN(n3295)
         );
  XNOR2_X1 U4231 ( .A(n3486), .B(n3360), .ZN(n3297) );
  NAND2_X1 U4232 ( .A1(n3297), .A2(n3327), .ZN(n3341) );
  NAND2_X1 U4233 ( .A1(n3298), .A2(n3341), .ZN(n3339) );
  INV_X1 U4234 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3301) );
  AOI21_X1 U4235 ( .B1(n4240), .B2(n3481), .A(n6421), .ZN(n3300) );
  NAND2_X1 U4236 ( .A1(n4332), .A2(n3360), .ZN(n3299) );
  OAI211_X1 U4237 ( .C1(n3538), .C2(n3301), .A(n3300), .B(n3299), .ZN(n3340)
         );
  NOR2_X1 U4238 ( .A1(n3486), .A2(n3378), .ZN(n3302) );
  AOI21_X1 U4239 ( .B1(n3339), .B2(n3340), .A(n3302), .ZN(n3354) );
  NAND2_X1 U4240 ( .A1(n3353), .A2(n3354), .ZN(n3358) );
  NAND2_X1 U4241 ( .A1(n3358), .A2(n3303), .ZN(n3369) );
  INV_X1 U4242 ( .A(n3304), .ZN(n3307) );
  NAND2_X1 U4243 ( .A1(n3308), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3315) );
  AND2_X1 U4244 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3309) );
  NAND2_X1 U4245 ( .A1(n3309), .A2(n5030), .ZN(n4742) );
  INV_X1 U4246 ( .A(n3309), .ZN(n3310) );
  NAND2_X1 U4247 ( .A1(n3310), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3311) );
  NAND2_X1 U4248 ( .A1(n4742), .A2(n3311), .ZN(n4712) );
  AOI22_X1 U4249 ( .A1(n3313), .A2(n4712), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3312), .ZN(n3314) );
  XNOR2_X1 U4250 ( .A(n3371), .B(n3372), .ZN(n4417) );
  NAND2_X1 U4251 ( .A1(n4417), .A2(n6421), .ZN(n3329) );
  AOI22_X1 U4252 ( .A1(n3819), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3247), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4253 ( .A1(n4174), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3319) );
  AOI22_X1 U4254 ( .A1(n4208), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4255 ( .A1(n4215), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3317) );
  NAND4_X1 U4256 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n3326)
         );
  AOI22_X1 U4257 ( .A1(n3425), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4258 ( .A1(n4532), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3323) );
  AOI22_X1 U4259 ( .A1(n4195), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3322) );
  AOI22_X1 U4260 ( .A1(n3803), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3321) );
  NAND4_X1 U4261 ( .A1(n3324), .A2(n3323), .A3(n3322), .A4(n3321), .ZN(n3325)
         );
  NAND2_X1 U4262 ( .A1(n3327), .A2(n3334), .ZN(n3328) );
  AOI22_X1 U4263 ( .A1(n3559), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3330), 
        .B2(n3334), .ZN(n3331) );
  NAND2_X1 U4264 ( .A1(n4562), .A2(n2957), .ZN(n3338) );
  NAND2_X1 U4265 ( .A1(n3359), .A2(n3360), .ZN(n3393) );
  INV_X1 U4266 ( .A(n3334), .ZN(n3392) );
  XNOR2_X1 U4267 ( .A(n3393), .B(n3392), .ZN(n3336) );
  AND2_X1 U4268 ( .A1(n4332), .A2(n3219), .ZN(n3345) );
  AOI21_X1 U4269 ( .B1(n3336), .B2(n3335), .A(n3345), .ZN(n3337) );
  NAND2_X1 U4270 ( .A1(n6163), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3367)
         );
  NAND2_X1 U4271 ( .A1(n3339), .A2(n3340), .ZN(n3344) );
  INV_X1 U4272 ( .A(n3340), .ZN(n3342) );
  OR2_X1 U4273 ( .A1(n4559), .A2(n3533), .ZN(n3349) );
  INV_X1 U4274 ( .A(n3335), .ZN(n6523) );
  INV_X1 U4275 ( .A(n3345), .ZN(n3346) );
  OAI21_X1 U4276 ( .B1(n6523), .B2(n3360), .A(n3346), .ZN(n3347) );
  INV_X1 U4277 ( .A(n3347), .ZN(n3348) );
  NAND2_X1 U4278 ( .A1(n3349), .A2(n3348), .ZN(n4350) );
  NAND2_X1 U4279 ( .A1(n4350), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3350)
         );
  INV_X1 U4280 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4453) );
  NAND2_X1 U4281 ( .A1(n3350), .A2(n4453), .ZN(n3352) );
  AND2_X1 U4282 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3351) );
  NAND2_X1 U4283 ( .A1(n4350), .A2(n3351), .ZN(n3365) );
  AND2_X1 U4284 ( .A1(n3352), .A2(n3365), .ZN(n4451) );
  INV_X1 U4285 ( .A(n3353), .ZN(n3356) );
  INV_X1 U4286 ( .A(n3354), .ZN(n3355) );
  NAND2_X1 U4287 ( .A1(n3356), .A2(n3355), .ZN(n3357) );
  NAND2_X1 U4288 ( .A1(n3358), .A2(n3357), .ZN(n4563) );
  NAND2_X1 U4289 ( .A1(n2963), .A2(n2957), .ZN(n3364) );
  OAI21_X1 U4290 ( .B1(n3360), .B2(n3359), .A(n3393), .ZN(n3361) );
  INV_X1 U4291 ( .A(n3714), .ZN(n3585) );
  OAI211_X1 U4292 ( .C1(n3361), .C2(n6523), .A(n3585), .B(n4607), .ZN(n3362)
         );
  INV_X1 U4293 ( .A(n3362), .ZN(n3363) );
  NAND2_X1 U4294 ( .A1(n3364), .A2(n3363), .ZN(n4450) );
  INV_X1 U4295 ( .A(n3365), .ZN(n3366) );
  AOI21_X2 U4296 ( .B1(n4451), .B2(n4450), .A(n3366), .ZN(n6162) );
  NAND2_X1 U4297 ( .A1(n3367), .A2(n6162), .ZN(n3368) );
  INV_X1 U4298 ( .A(n3371), .ZN(n3373) );
  NAND2_X1 U4299 ( .A1(n3308), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3377) );
  NOR3_X1 U4300 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5030), .A3(n6394), 
        .ZN(n6311) );
  NAND2_X1 U4301 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6311), .ZN(n6301) );
  NAND2_X1 U4302 ( .A1(n6263), .A2(n6301), .ZN(n3374) );
  NOR3_X1 U4303 ( .A1(n6263), .A2(n5030), .A3(n6394), .ZN(n4950) );
  NAND2_X1 U4304 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4950), .ZN(n4947) );
  NAND2_X1 U4305 ( .A1(n3374), .A2(n4947), .ZN(n4908) );
  OAI22_X1 U4306 ( .A1(n4296), .A2(n4908), .B1(n3591), .B2(n6263), .ZN(n3375)
         );
  INV_X1 U4307 ( .A(n3375), .ZN(n3376) );
  NAND2_X1 U4308 ( .A1(n4527), .A2(n6421), .ZN(n3391) );
  AOI22_X1 U4309 ( .A1(n3819), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4310 ( .A1(n4174), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4311 ( .A1(n4208), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4312 ( .A1(n4215), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3380) );
  NAND4_X1 U4313 ( .A1(n3383), .A2(n3382), .A3(n3381), .A4(n3380), .ZN(n3389)
         );
  AOI22_X1 U4314 ( .A1(n3425), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3387) );
  AOI22_X1 U4315 ( .A1(n4532), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4316 ( .A1(n4195), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3385) );
  INV_X1 U4317 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U4318 ( .A1(n3803), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3384) );
  NAND4_X1 U4319 ( .A1(n3387), .A2(n3386), .A3(n3385), .A4(n3384), .ZN(n3388)
         );
  AOI22_X1 U4320 ( .A1(n3548), .A2(n3413), .B1(n3559), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3390) );
  NAND2_X1 U4321 ( .A1(n3767), .A2(n2957), .ZN(n3397) );
  NAND2_X1 U4322 ( .A1(n3393), .A2(n3392), .ZN(n3414) );
  INV_X1 U4323 ( .A(n3413), .ZN(n3394) );
  XNOR2_X1 U4324 ( .A(n3414), .B(n3394), .ZN(n3395) );
  NAND2_X1 U4325 ( .A1(n3395), .A2(n3335), .ZN(n3396) );
  NAND2_X1 U4326 ( .A1(n3397), .A2(n3396), .ZN(n3398) );
  INV_X1 U4327 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6233) );
  XNOR2_X1 U4328 ( .A(n3398), .B(n6233), .ZN(n6153) );
  NAND2_X1 U4329 ( .A1(n6154), .A2(n6153), .ZN(n6156) );
  NAND2_X1 U4330 ( .A1(n3398), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3399)
         );
  NAND2_X1 U4331 ( .A1(n6156), .A2(n3399), .ZN(n4571) );
  AOI22_X1 U4332 ( .A1(n4150), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4333 ( .A1(n4174), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4334 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n4208), .B1(n3261), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3402) );
  AOI22_X1 U4335 ( .A1(n4215), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3401) );
  NAND4_X1 U4336 ( .A1(n3404), .A2(n3403), .A3(n3402), .A4(n3401), .ZN(n3410)
         );
  AOI22_X1 U4337 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3425), .B1(n3253), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3408) );
  AOI22_X1 U4338 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4532), .B1(n3289), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3407) );
  AOI22_X1 U4339 ( .A1(n4195), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3406) );
  AOI22_X1 U4340 ( .A1(n3803), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3405) );
  NAND4_X1 U4341 ( .A1(n3408), .A2(n3407), .A3(n3406), .A4(n3405), .ZN(n3409)
         );
  NAND2_X1 U4342 ( .A1(n3548), .A2(n3462), .ZN(n3412) );
  NAND2_X1 U4343 ( .A1(n3559), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3411) );
  NAND2_X1 U4344 ( .A1(n3412), .A2(n3411), .ZN(n3443) );
  XNOR2_X1 U4345 ( .A(n3442), .B(n3443), .ZN(n3783) );
  NAND2_X1 U4346 ( .A1(n3783), .A2(n2957), .ZN(n3417) );
  NAND2_X1 U4347 ( .A1(n3414), .A2(n3413), .ZN(n3464) );
  XNOR2_X1 U4348 ( .A(n3464), .B(n3462), .ZN(n3415) );
  NAND2_X1 U4349 ( .A1(n3415), .A2(n3335), .ZN(n3416) );
  NAND2_X1 U4350 ( .A1(n3417), .A2(n3416), .ZN(n3418) );
  INV_X1 U4351 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6227) );
  XNOR2_X1 U4352 ( .A(n3418), .B(n6227), .ZN(n4568) );
  NAND2_X1 U4353 ( .A1(n4571), .A2(n4568), .ZN(n4569) );
  NAND2_X1 U4354 ( .A1(n3418), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3419)
         );
  NAND2_X1 U4355 ( .A1(n4569), .A2(n3419), .ZN(n4597) );
  INV_X1 U4356 ( .A(n3442), .ZN(n3420) );
  AOI22_X1 U4357 ( .A1(n3819), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3424) );
  AOI22_X1 U4358 ( .A1(n4174), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3423) );
  AOI22_X1 U4359 ( .A1(n4208), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3422) );
  AOI22_X1 U4360 ( .A1(n4215), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3421) );
  NAND4_X1 U4361 ( .A1(n3424), .A2(n3423), .A3(n3422), .A4(n3421), .ZN(n3431)
         );
  AOI22_X1 U4362 ( .A1(n3425), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4363 ( .A1(n4532), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4364 ( .A1(n4195), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3427) );
  INV_X1 U4365 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U4366 ( .A1(n3803), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3426) );
  NAND4_X1 U4367 ( .A1(n3429), .A2(n3428), .A3(n3427), .A4(n3426), .ZN(n3430)
         );
  NAND2_X1 U4368 ( .A1(n3548), .A2(n3461), .ZN(n3433) );
  NAND2_X1 U4369 ( .A1(n3559), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3432) );
  NAND2_X1 U4370 ( .A1(n3433), .A2(n3432), .ZN(n3444) );
  NAND2_X1 U4371 ( .A1(n3784), .A2(n2957), .ZN(n3439) );
  INV_X1 U4372 ( .A(n3462), .ZN(n3435) );
  OR2_X1 U4373 ( .A1(n3464), .A2(n3435), .ZN(n3436) );
  XNOR2_X1 U4374 ( .A(n3436), .B(n3461), .ZN(n3437) );
  NAND2_X1 U4375 ( .A1(n3437), .A2(n3335), .ZN(n3438) );
  NAND2_X1 U4376 ( .A1(n3439), .A2(n3438), .ZN(n3440) );
  INV_X1 U4377 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4687) );
  XNOR2_X1 U4378 ( .A(n3440), .B(n4687), .ZN(n4595) );
  NAND2_X1 U4379 ( .A1(n4597), .A2(n4595), .ZN(n4596) );
  NAND2_X1 U4380 ( .A1(n3440), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3441)
         );
  INV_X1 U4381 ( .A(n3444), .ZN(n3445) );
  AOI22_X1 U4382 ( .A1(n4150), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4383 ( .A1(n4174), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4384 ( .A1(n4208), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4385 ( .A1(n4215), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3448) );
  NAND4_X1 U4386 ( .A1(n3451), .A2(n3450), .A3(n3449), .A4(n3448), .ZN(n3457)
         );
  AOI22_X1 U4387 ( .A1(n3425), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4388 ( .A1(n4532), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4389 ( .A1(n4195), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4390 ( .A1(n3803), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3452) );
  NAND4_X1 U4391 ( .A1(n3455), .A2(n3454), .A3(n3453), .A4(n3452), .ZN(n3456)
         );
  AOI22_X1 U4392 ( .A1(n3548), .A2(n3474), .B1(n3559), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3459) );
  INV_X1 U4393 ( .A(n3459), .ZN(n3458) );
  NAND2_X1 U4394 ( .A1(n3460), .A2(n3459), .ZN(n3795) );
  NAND3_X1 U4395 ( .A1(n3485), .A2(n2957), .A3(n3795), .ZN(n3467) );
  NAND2_X1 U4396 ( .A1(n3462), .A2(n3461), .ZN(n3463) );
  OR2_X1 U4397 ( .A1(n3464), .A2(n3463), .ZN(n3473) );
  XNOR2_X1 U4398 ( .A(n3473), .B(n3474), .ZN(n3465) );
  NAND2_X1 U4399 ( .A1(n3465), .A2(n3335), .ZN(n3466) );
  NAND2_X1 U4400 ( .A1(n3467), .A2(n3466), .ZN(n3468) );
  INV_X1 U4401 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6219) );
  XNOR2_X1 U4402 ( .A(n3468), .B(n6219), .ZN(n6146) );
  NAND2_X1 U4403 ( .A1(n3468), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3469)
         );
  INV_X1 U4404 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3471) );
  NAND2_X1 U4405 ( .A1(n3548), .A2(n3481), .ZN(n3470) );
  OAI21_X1 U4406 ( .B1(n3471), .B2(n3538), .A(n3470), .ZN(n3472) );
  NAND2_X1 U4407 ( .A1(n3802), .A2(n2957), .ZN(n3478) );
  INV_X1 U4408 ( .A(n3473), .ZN(n3475) );
  NAND2_X1 U4409 ( .A1(n3475), .A2(n3474), .ZN(n3487) );
  XNOR2_X1 U4410 ( .A(n3487), .B(n3481), .ZN(n3476) );
  NAND2_X1 U4411 ( .A1(n3476), .A2(n3335), .ZN(n3477) );
  INV_X1 U4412 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3479) );
  NAND2_X1 U4413 ( .A1(n3481), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3482) );
  OR3_X1 U4414 ( .A1(n3487), .A2(n3486), .A3(n6523), .ZN(n3488) );
  NAND2_X1 U4415 ( .A1(n3496), .A2(n3488), .ZN(n3490) );
  INV_X1 U4416 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3489) );
  XNOR2_X1 U4417 ( .A(n3490), .B(n3489), .ZN(n5017) );
  NAND2_X1 U4418 ( .A1(n3490), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3491)
         );
  INV_X4 U4419 ( .A(n3492), .ZN(n5648) );
  INV_X1 U4420 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6193) );
  NAND2_X1 U4421 ( .A1(n5648), .A2(n6193), .ZN(n5181) );
  NAND2_X1 U4422 ( .A1(n3492), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5182)
         );
  INV_X1 U4423 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3494) );
  NAND2_X1 U4424 ( .A1(n5648), .A2(n3494), .ZN(n5261) );
  INV_X1 U4425 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3495) );
  NAND2_X1 U4426 ( .A1(n3492), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U4427 ( .A1(n3492), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3497) );
  AND2_X1 U4428 ( .A1(n6134), .A2(n3497), .ZN(n3498) );
  NAND2_X1 U4429 ( .A1(n3499), .A2(n3498), .ZN(n5301) );
  INV_X1 U4430 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6177) );
  NOR2_X1 U4431 ( .A1(n5648), .A2(n6177), .ZN(n5297) );
  NAND2_X1 U4432 ( .A1(n5648), .A2(n6177), .ZN(n5298) );
  XNOR2_X1 U4433 ( .A(n5648), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5338)
         );
  NAND2_X1 U4434 ( .A1(n5337), .A2(n5338), .ZN(n3501) );
  NAND2_X1 U4435 ( .A1(n5648), .A2(n3726), .ZN(n3500) );
  INV_X1 U4436 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3502) );
  NAND2_X1 U4437 ( .A1(n3492), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3503) );
  INV_X1 U4438 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6570) );
  XNOR2_X1 U4439 ( .A(n5648), .B(n6570), .ZN(n5719) );
  NAND2_X1 U4440 ( .A1(n5648), .A2(n6570), .ZN(n3505) );
  INV_X1 U4441 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5934) );
  INV_X1 U4442 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5824) );
  INV_X1 U4443 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5829) );
  NAND2_X1 U4444 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3727) );
  AND2_X1 U4445 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5786) );
  AND2_X1 U4446 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5808) );
  AND2_X1 U4447 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3744) );
  NAND3_X1 U4448 ( .A1(n5786), .A2(n5808), .A3(n3744), .ZN(n3507) );
  NAND2_X1 U4449 ( .A1(n5648), .A2(n3507), .ZN(n3510) );
  NOR2_X1 U4450 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5807) );
  NOR2_X1 U4451 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5785) );
  INV_X1 U4452 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5778) );
  INV_X1 U4453 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3685) );
  AND4_X1 U4454 ( .A1(n5807), .A2(n5785), .A3(n5778), .A4(n3685), .ZN(n3508)
         );
  NOR2_X1 U4455 ( .A1(n5648), .A2(n3508), .ZN(n3509) );
  XNOR2_X1 U4456 ( .A(n5648), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5641)
         );
  NAND2_X1 U4457 ( .A1(n5640), .A2(n5641), .ZN(n3512) );
  INV_X1 U4458 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5612) );
  AND2_X2 U4459 ( .A1(n3512), .A2(n3511), .ZN(n5611) );
  NAND2_X1 U4460 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U4461 ( .A1(n4272), .A2(n3073), .ZN(n3516) );
  OR2_X1 U4462 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5736) );
  NOR3_X1 U4463 ( .A1(n5648), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n5736), 
        .ZN(n4259) );
  INV_X1 U4464 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4266) );
  INV_X1 U4465 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4282) );
  NAND2_X1 U4466 ( .A1(n3516), .A2(n3515), .ZN(n3517) );
  XNOR2_X1 U4467 ( .A(n3517), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4305)
         );
  OR2_X1 U4468 ( .A1(n3519), .A2(STATE_REG_0__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U4469 ( .A1(n3536), .A2(n6440), .ZN(n4994) );
  NAND3_X1 U4470 ( .A1(n3518), .A2(n4994), .A3(n6520), .ZN(n3521) );
  NAND3_X1 U4471 ( .A1(n3521), .A2(n4993), .A3(n3520), .ZN(n3570) );
  XNOR2_X1 U4472 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3539) );
  NAND2_X1 U4473 ( .A1(n3540), .A2(n3539), .ZN(n3523) );
  NAND2_X1 U4474 ( .A1(n6394), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3522) );
  NAND2_X1 U4475 ( .A1(n3523), .A2(n3522), .ZN(n3535) );
  XNOR2_X1 U4476 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3534) );
  NAND2_X1 U4477 ( .A1(n3535), .A2(n3534), .ZN(n3525) );
  NAND2_X1 U4478 ( .A1(n5030), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3524) );
  XNOR2_X1 U4479 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3529) );
  NOR2_X1 U4480 ( .A1(n3526), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3527)
         );
  NAND2_X1 U4481 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6614), .ZN(n3528) );
  NAND2_X1 U4482 ( .A1(n3548), .A2(n3575), .ZN(n3566) );
  XOR2_X1 U4483 ( .A(n3530), .B(n3529), .Z(n3571) );
  NAND2_X1 U4484 ( .A1(n3532), .A2(n3531), .ZN(n3576) );
  INV_X1 U4485 ( .A(n3567), .ZN(n3562) );
  XOR2_X1 U4486 ( .A(n3535), .B(n3534), .Z(n3572) );
  NAND2_X1 U4487 ( .A1(n3572), .A2(n3548), .ZN(n3537) );
  INV_X1 U4488 ( .A(n3537), .ZN(n3558) );
  INV_X1 U4489 ( .A(n3545), .ZN(n3557) );
  OAI211_X1 U4490 ( .C1(n3572), .C2(n3538), .A(n3545), .B(n3537), .ZN(n3556)
         );
  AOI21_X1 U4491 ( .B1(n3548), .B2(n2958), .A(n3210), .ZN(n3554) );
  XOR2_X1 U4492 ( .A(n3540), .B(n3539), .Z(n3573) );
  NAND2_X1 U4493 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n3573), .ZN(n3553) );
  INV_X1 U4494 ( .A(n3573), .ZN(n3546) );
  NAND2_X1 U4495 ( .A1(n4240), .A2(n4607), .ZN(n3594) );
  INV_X1 U4496 ( .A(n3594), .ZN(n3543) );
  INV_X1 U4497 ( .A(n3540), .ZN(n3542) );
  INV_X2 U4498 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U4499 ( .A1(n5367), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3541) );
  NAND2_X1 U4500 ( .A1(n3542), .A2(n3541), .ZN(n3547) );
  OAI21_X1 U4501 ( .B1(n3543), .B2(n3547), .A(n4993), .ZN(n3544) );
  AOI22_X1 U4502 ( .A1(n3545), .A2(n3544), .B1(n3554), .B2(n3553), .ZN(n3549)
         );
  OAI21_X1 U4503 ( .B1(n3546), .B2(n3549), .A(n3567), .ZN(n3552) );
  INV_X1 U4504 ( .A(n3547), .ZN(n3550) );
  NAND3_X1 U4505 ( .A1(n3550), .A2(n3549), .A3(n3548), .ZN(n3551) );
  OAI211_X1 U4506 ( .C1(n3554), .C2(n3553), .A(n3552), .B(n3551), .ZN(n3555)
         );
  AOI22_X1 U4507 ( .A1(n3558), .A2(n3557), .B1(n3556), .B2(n3555), .ZN(n3561)
         );
  NOR2_X1 U4508 ( .A1(n3559), .A2(n3563), .ZN(n3560) );
  OAI22_X1 U4509 ( .A1(n3563), .A2(n3562), .B1(n3561), .B2(n3560), .ZN(n3564)
         );
  AOI21_X1 U4510 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6421), .A(n3564), 
        .ZN(n3565) );
  NAND2_X1 U4511 ( .A1(n3566), .A2(n3565), .ZN(n3569) );
  NAND2_X1 U4512 ( .A1(n3567), .A2(n3575), .ZN(n3568) );
  NAND2_X1 U4513 ( .A1(n3570), .A2(n5401), .ZN(n3580) );
  NAND2_X1 U4514 ( .A1(n2958), .A2(n6440), .ZN(n3578) );
  AND3_X1 U4515 ( .A1(n3573), .A2(n3572), .A3(n3571), .ZN(n3574) );
  OR2_X1 U4516 ( .A1(n3575), .A2(n3574), .ZN(n3577) );
  NOR2_X1 U4517 ( .A1(n5395), .A2(READY_N), .ZN(n4318) );
  NAND2_X1 U4518 ( .A1(n3578), .A2(n4318), .ZN(n3579) );
  MUX2_X1 U4519 ( .A(n3580), .B(n3579), .S(n4621), .Z(n3590) );
  NAND2_X1 U4520 ( .A1(n3581), .A2(n4607), .ZN(n4438) );
  AND2_X1 U4521 ( .A1(n3712), .A2(n2958), .ZN(n4242) );
  INV_X1 U4522 ( .A(n4242), .ZN(n4400) );
  INV_X1 U4523 ( .A(n4238), .ZN(n3589) );
  AND2_X1 U4524 ( .A1(n3582), .A2(n4993), .ZN(n3584) );
  MUX2_X1 U4525 ( .A(n3584), .B(n3335), .S(n3583), .Z(n3717) );
  NAND2_X1 U4526 ( .A1(n4438), .A2(n4332), .ZN(n3586) );
  NAND3_X1 U4527 ( .A1(n3243), .A2(n3586), .A3(n3585), .ZN(n3595) );
  INV_X1 U4528 ( .A(n5396), .ZN(n3588) );
  OAI21_X1 U4529 ( .B1(n3717), .B2(n3595), .A(n3588), .ZN(n4399) );
  NAND3_X1 U4530 ( .A1(n3590), .A2(n3589), .A3(n4399), .ZN(n3592) );
  INV_X1 U4531 ( .A(n5402), .ZN(n3593) );
  NOR2_X1 U4532 ( .A1(n3595), .A2(n3593), .ZN(n4317) );
  INV_X1 U4533 ( .A(n4317), .ZN(n5394) );
  NOR2_X1 U4534 ( .A1(n3595), .A2(n3594), .ZN(n4287) );
  INV_X1 U4535 ( .A(n4287), .ZN(n5393) );
  AND2_X1 U4536 ( .A1(n3518), .A2(n4998), .ZN(n4403) );
  NOR2_X1 U4537 ( .A1(n3596), .A2(n4240), .ZN(n3597) );
  NOR2_X1 U4538 ( .A1(n4403), .A2(n3597), .ZN(n3599) );
  NAND4_X1 U4539 ( .A1(n5394), .A2(n5393), .A3(n3599), .A4(n3598), .ZN(n3600)
         );
  NAND2_X1 U4540 ( .A1(n4327), .A2(n4240), .ZN(n3602) );
  NAND2_X1 U4541 ( .A1(n3518), .A2(n3335), .ZN(n4336) );
  OAI21_X1 U4542 ( .B1(n3601), .B2(n3602), .A(n4336), .ZN(n3603) );
  AND2_X2 U4543 ( .A1(n3219), .A2(n2958), .ZN(n5561) );
  INV_X1 U4544 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3604) );
  NAND2_X1 U4545 ( .A1(n4241), .A2(n2956), .ZN(n3657) );
  NAND2_X1 U4546 ( .A1(n4241), .A2(EBX_REG_1__SCAN_IN), .ZN(n3607) );
  NAND2_X1 U4547 ( .A1(n2956), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3606)
         );
  NAND4_X1 U4548 ( .A1(n3608), .A2(n3657), .A3(n3607), .A4(n3606), .ZN(n3611)
         );
  INV_X1 U4549 ( .A(EBX_REG_0__SCAN_IN), .ZN(n6626) );
  NAND2_X1 U4550 ( .A1(n3617), .A2(n6626), .ZN(n3610) );
  INV_X2 U4551 ( .A(n4241), .ZN(n3698) );
  NAND2_X1 U4552 ( .A1(n3698), .A2(EBX_REG_0__SCAN_IN), .ZN(n3609) );
  INV_X1 U4553 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U4554 ( .A1(n4998), .A2(n6075), .ZN(n3612) );
  OAI211_X1 U4555 ( .C1(n4241), .C2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(n3612), 
        .B(n3617), .ZN(n3614) );
  NAND2_X1 U4556 ( .A1(n3614), .A2(n3613), .ZN(n5199) );
  INV_X1 U4557 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U4558 ( .A1(n4998), .A2(n6071), .ZN(n3616) );
  NAND2_X1 U4559 ( .A1(n3617), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3615)
         );
  NAND3_X1 U4560 ( .A1(n3698), .A2(n3616), .A3(n3615), .ZN(n3619) );
  NAND2_X1 U4561 ( .A1(n3690), .A2(n6071), .ZN(n3618) );
  NAND2_X1 U4562 ( .A1(n3619), .A2(n3618), .ZN(n6045) );
  INV_X1 U4563 ( .A(EBX_REG_4__SCAN_IN), .ZN(n3620) );
  NAND2_X1 U4564 ( .A1(n4241), .A2(EBX_REG_4__SCAN_IN), .ZN(n3622) );
  NAND2_X1 U4565 ( .A1(n3709), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3621)
         );
  NAND4_X1 U4566 ( .A1(n3623), .A2(n3657), .A3(n3622), .A4(n3621), .ZN(n4503)
         );
  INV_X1 U4567 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4498) );
  NAND2_X1 U4568 ( .A1(n4998), .A2(n4498), .ZN(n3625) );
  NAND2_X1 U4569 ( .A1(n3617), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3624)
         );
  NAND3_X1 U4570 ( .A1(n3698), .A2(n3625), .A3(n3624), .ZN(n3627) );
  NAND2_X1 U4571 ( .A1(n3690), .A2(n4498), .ZN(n3626) );
  NAND2_X1 U4572 ( .A1(n3627), .A2(n3626), .ZN(n4497) );
  INV_X1 U4573 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U4574 ( .A1(n4998), .A2(n6537), .ZN(n3628) );
  OAI211_X1 U4575 ( .C1(n4241), .C2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n3628), 
        .B(n3617), .ZN(n3630) );
  NAND2_X1 U4576 ( .A1(n3630), .A2(n3629), .ZN(n4582) );
  NAND2_X1 U4577 ( .A1(n4581), .A2(n4582), .ZN(n4589) );
  INV_X1 U4578 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5007) );
  NAND2_X1 U4579 ( .A1(n4998), .A2(n5007), .ZN(n3632) );
  NAND2_X1 U4580 ( .A1(n3617), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3631)
         );
  NAND3_X1 U4581 ( .A1(n3698), .A2(n3632), .A3(n3631), .ZN(n3634) );
  NAND2_X1 U4582 ( .A1(n3690), .A2(n5007), .ZN(n3633) );
  NAND2_X1 U4583 ( .A1(n3634), .A2(n3633), .ZN(n4590) );
  INV_X1 U4584 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5191) );
  NAND2_X1 U4585 ( .A1(n4241), .A2(EBX_REG_8__SCAN_IN), .ZN(n3636) );
  NAND2_X1 U4586 ( .A1(n3709), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3635)
         );
  NAND4_X1 U4587 ( .A1(n3637), .A2(n3657), .A3(n3636), .A4(n3635), .ZN(n4801)
         );
  NAND2_X1 U4588 ( .A1(n4802), .A2(n4801), .ZN(n6009) );
  INV_X1 U4589 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6576) );
  NAND2_X1 U4590 ( .A1(n4998), .A2(n6576), .ZN(n3639) );
  NAND2_X1 U4591 ( .A1(n3617), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3638)
         );
  NAND3_X1 U4592 ( .A1(n3698), .A2(n3639), .A3(n3638), .ZN(n3641) );
  NAND2_X1 U4593 ( .A1(n3690), .A2(n6576), .ZN(n3640) );
  NAND2_X1 U4594 ( .A1(n3641), .A2(n3640), .ZN(n6010) );
  INV_X1 U4595 ( .A(EBX_REG_10__SCAN_IN), .ZN(n3642) );
  NAND2_X1 U4596 ( .A1(n4241), .A2(EBX_REG_10__SCAN_IN), .ZN(n3644) );
  NAND2_X1 U4597 ( .A1(n3709), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3643) );
  NAND4_X1 U4598 ( .A1(n3645), .A2(n3657), .A3(n3644), .A4(n3643), .ZN(n5142)
         );
  INV_X1 U4599 ( .A(n3690), .ZN(n3700) );
  NAND2_X1 U4600 ( .A1(EBX_REG_11__SCAN_IN), .A2(n5561), .ZN(n3647) );
  INV_X1 U4601 ( .A(n4359), .ZN(n3704) );
  NAND2_X1 U4602 ( .A1(n3704), .A2(n3495), .ZN(n3646) );
  OAI211_X1 U4603 ( .C1(EBX_REG_11__SCAN_IN), .C2(n3700), .A(n3647), .B(n3646), 
        .ZN(n5222) );
  INV_X1 U4604 ( .A(EBX_REG_12__SCAN_IN), .ZN(n3648) );
  NAND2_X1 U4605 ( .A1(n4241), .A2(EBX_REG_12__SCAN_IN), .ZN(n3650) );
  NAND2_X1 U4606 ( .A1(n3709), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3649) );
  NAND4_X1 U4607 ( .A1(n3651), .A2(n3657), .A3(n3650), .A4(n3649), .ZN(n5287)
         );
  NAND2_X1 U4608 ( .A1(n5561), .A2(EBX_REG_13__SCAN_IN), .ZN(n3654) );
  INV_X1 U4609 ( .A(EBX_REG_13__SCAN_IN), .ZN(n3652) );
  NAND2_X1 U4610 ( .A1(n3690), .A2(n3652), .ZN(n3653) );
  OAI211_X1 U4611 ( .C1(n4359), .C2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n3654), .B(n3653), .ZN(n5330) );
  INV_X1 U4612 ( .A(EBX_REG_14__SCAN_IN), .ZN(n3655) );
  NAND2_X1 U4613 ( .A1(n4241), .A2(EBX_REG_14__SCAN_IN), .ZN(n3658) );
  NAND2_X1 U4614 ( .A1(n3709), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3656) );
  NAND4_X1 U4615 ( .A1(n3659), .A2(n3658), .A3(n3657), .A4(n3656), .ZN(n5318)
         );
  NAND2_X1 U4616 ( .A1(n5317), .A2(n5318), .ZN(n5835) );
  INV_X1 U4617 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U4618 ( .A1(n4998), .A2(n6064), .ZN(n3661) );
  NAND2_X1 U4619 ( .A1(n3617), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3660) );
  NAND3_X1 U4620 ( .A1(n3698), .A2(n3661), .A3(n3660), .ZN(n3663) );
  NAND2_X1 U4621 ( .A1(n3690), .A2(n6064), .ZN(n3662) );
  NAND2_X1 U4622 ( .A1(n3663), .A2(n3662), .ZN(n5836) );
  NAND2_X1 U4623 ( .A1(n3709), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3665) );
  NAND2_X1 U4624 ( .A1(n4241), .A2(EBX_REG_16__SCAN_IN), .ZN(n3664) );
  OAI211_X1 U4625 ( .C1(n3705), .C2(EBX_REG_16__SCAN_IN), .A(n3665), .B(n3664), 
        .ZN(n5516) );
  INV_X1 U4626 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6639) );
  NAND2_X1 U4627 ( .A1(n3690), .A2(n6639), .ZN(n3668) );
  NAND2_X1 U4628 ( .A1(n3617), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3666) );
  OAI211_X1 U4629 ( .C1(n3709), .C2(EBX_REG_17__SCAN_IN), .A(n3698), .B(n3666), 
        .ZN(n3667) );
  AOI22_X1 U4630 ( .A1(n4241), .A2(EBX_REG_19__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n3709), .ZN(n3670) );
  INV_X1 U4631 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5496) );
  OR2_X1 U4632 ( .A1(n4359), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3673)
         );
  INV_X1 U4633 ( .A(EBX_REG_20__SCAN_IN), .ZN(n3671) );
  NAND2_X1 U4634 ( .A1(n4998), .A2(n3671), .ZN(n3672) );
  AND2_X1 U4635 ( .A1(n3673), .A2(n3672), .ZN(n5563) );
  OR2_X1 U4636 ( .A1(n4359), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3674)
         );
  INV_X1 U4637 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U4638 ( .A1(n4998), .A2(n5573), .ZN(n5491) );
  NAND2_X1 U4639 ( .A1(n3674), .A2(n5491), .ZN(n5490) );
  NAND2_X1 U4640 ( .A1(n5561), .A2(EBX_REG_20__SCAN_IN), .ZN(n3676) );
  NAND2_X1 U4641 ( .A1(n5490), .A2(n3617), .ZN(n3675) );
  OAI211_X1 U4642 ( .C1(n5563), .C2(n5490), .A(n3676), .B(n3675), .ZN(n3677)
         );
  OR2_X1 U4643 ( .A1(n4359), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3680)
         );
  INV_X1 U4644 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U4645 ( .A1(n3690), .A2(n5558), .ZN(n3679) );
  NAND2_X1 U4646 ( .A1(n5561), .A2(EBX_REG_21__SCAN_IN), .ZN(n3678) );
  NAND2_X1 U4647 ( .A1(n5556), .A2(n5555), .ZN(n5548) );
  AOI22_X1 U4648 ( .A1(n4241), .A2(EBX_REG_22__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n3709), .ZN(n3682) );
  INV_X1 U4649 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U4650 ( .A1(n3617), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3683) );
  OAI211_X1 U4651 ( .C1(n3709), .C2(EBX_REG_23__SCAN_IN), .A(n3698), .B(n3683), 
        .ZN(n3684) );
  OAI21_X1 U4652 ( .B1(n3700), .B2(EBX_REG_23__SCAN_IN), .A(n3684), .ZN(n5480)
         );
  NAND2_X1 U4653 ( .A1(n3698), .A2(n3685), .ZN(n3687) );
  INV_X1 U4654 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U4655 ( .A1(n4998), .A2(n5881), .ZN(n3686) );
  NAND3_X1 U4656 ( .A1(n3687), .A2(n3617), .A3(n3686), .ZN(n3688) );
  OAI21_X1 U4657 ( .B1(n3705), .B2(EBX_REG_24__SCAN_IN), .A(n3688), .ZN(n5538)
         );
  INV_X1 U4658 ( .A(EBX_REG_25__SCAN_IN), .ZN(n3689) );
  NAND2_X1 U4659 ( .A1(n3690), .A2(n3689), .ZN(n3693) );
  NAND2_X1 U4660 ( .A1(n3617), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3691) );
  OAI211_X1 U4661 ( .C1(n3709), .C2(EBX_REG_25__SCAN_IN), .A(n3698), .B(n3691), 
        .ZN(n3692) );
  INV_X1 U4662 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5534) );
  INV_X1 U4663 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U4664 ( .A1(n3698), .A2(n5614), .ZN(n3694) );
  OAI211_X1 U4665 ( .C1(EBX_REG_26__SCAN_IN), .C2(n3709), .A(n3694), .B(n3617), 
        .ZN(n3695) );
  AND2_X1 U4666 ( .A1(n3696), .A2(n3695), .ZN(n5453) );
  NAND2_X1 U4667 ( .A1(n3617), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3697) );
  OAI211_X1 U4668 ( .C1(n3709), .C2(EBX_REG_27__SCAN_IN), .A(n3698), .B(n3697), 
        .ZN(n3699) );
  OAI21_X1 U4669 ( .B1(n3700), .B2(EBX_REG_27__SCAN_IN), .A(n3699), .ZN(n5440)
         );
  AOI22_X1 U4670 ( .A1(n4241), .A2(EBX_REG_28__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n3709), .ZN(n3702) );
  INV_X1 U4671 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5532) );
  AND2_X1 U4672 ( .A1(n3702), .A2(n3701), .ZN(n5425) );
  NOR2_X1 U4673 ( .A1(n3709), .A2(EBX_REG_29__SCAN_IN), .ZN(n3703) );
  AOI21_X1 U4674 ( .B1(n3704), .B2(n4282), .A(n3703), .ZN(n4273) );
  NAND2_X1 U4675 ( .A1(n5426), .A2(n4273), .ZN(n4250) );
  NOR2_X1 U4676 ( .A1(n3705), .A2(EBX_REG_29__SCAN_IN), .ZN(n4274) );
  NAND2_X1 U4677 ( .A1(n5426), .A2(n4274), .ZN(n3706) );
  OAI21_X1 U4678 ( .B1(n4250), .B2(n5561), .A(n3706), .ZN(n4279) );
  AND2_X1 U4679 ( .A1(n3709), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3707)
         );
  AOI21_X1 U4680 ( .B1(n4359), .B2(EBX_REG_30__SCAN_IN), .A(n3707), .ZN(n4249)
         );
  NAND2_X1 U4681 ( .A1(n4279), .A2(n4249), .ZN(n3708) );
  NAND2_X1 U4682 ( .A1(n4250), .A2(n3617), .ZN(n4248) );
  NAND2_X1 U4683 ( .A1(n3708), .A2(n4248), .ZN(n3711) );
  OAI22_X1 U4684 ( .A1(n4359), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n3709), .ZN(n3710) );
  INV_X1 U4685 ( .A(n5529), .ZN(n3741) );
  OR2_X1 U4686 ( .A1(n4242), .A2(n4359), .ZN(n3715) );
  AOI21_X1 U4687 ( .B1(n4327), .B2(n4332), .A(n3712), .ZN(n3713) );
  AOI21_X1 U4688 ( .B1(n3715), .B2(n3714), .A(n3713), .ZN(n3716) );
  OAI21_X1 U4689 ( .B1(n3243), .B2(n3617), .A(n3716), .ZN(n3718) );
  NOR2_X1 U4690 ( .A1(n3718), .A2(n3717), .ZN(n3720) );
  AND2_X1 U4691 ( .A1(n3720), .A2(n3719), .ZN(n4422) );
  OAI21_X1 U4692 ( .B1(n4420), .B2(n4993), .A(n4538), .ZN(n3721) );
  INV_X1 U4693 ( .A(n3721), .ZN(n3722) );
  NOR2_X1 U4694 ( .A1(n3729), .A2(n4239), .ZN(n5341) );
  INV_X1 U4695 ( .A(n5341), .ZN(n3730) );
  INV_X1 U4696 ( .A(n3723), .ZN(n3724) );
  NAND2_X1 U4697 ( .A1(n5332), .A2(n4684), .ZN(n5271) );
  AND2_X1 U4698 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5752) );
  INV_X1 U4699 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3726) );
  NAND2_X1 U4700 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6173) );
  NOR2_X1 U4701 ( .A1(n3726), .A2(n6173), .ZN(n5843) );
  NAND2_X1 U4702 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5843), .ZN(n5833) );
  NOR2_X1 U4703 ( .A1(n6570), .A2(n5833), .ZN(n5935) );
  NAND2_X1 U4704 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n5935), .ZN(n3742) );
  INV_X1 U4705 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6643) );
  NOR2_X1 U4706 ( .A1(n6643), .A2(n4453), .ZN(n5339) );
  NAND2_X1 U4707 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6224) );
  NOR2_X1 U4708 ( .A1(n4687), .A2(n6224), .ZN(n6214) );
  NAND2_X1 U4709 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6214), .ZN(n5269)
         );
  NAND2_X1 U4710 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U4711 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5273) );
  NOR3_X1 U4712 ( .A1(n5269), .A2(n6195), .A3(n5273), .ZN(n5342) );
  NAND2_X1 U4713 ( .A1(n5339), .A2(n5342), .ZN(n5345) );
  OR2_X1 U4714 ( .A1(n3742), .A2(n5345), .ZN(n5799) );
  INV_X1 U4715 ( .A(n3727), .ZN(n5805) );
  AND2_X1 U4716 ( .A1(n5805), .A2(n5808), .ZN(n3731) );
  INV_X1 U4717 ( .A(n3731), .ZN(n3743) );
  NOR2_X1 U4718 ( .A1(n5799), .A2(n3743), .ZN(n3728) );
  OR2_X1 U4719 ( .A1(n5332), .A2(n3728), .ZN(n3734) );
  INV_X1 U4720 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4431) );
  OAI21_X1 U4721 ( .B1(n4453), .B2(n4431), .A(n6643), .ZN(n4683) );
  INV_X1 U4722 ( .A(n4688), .ZN(n5340) );
  NAND2_X1 U4723 ( .A1(n5340), .A2(n5342), .ZN(n5333) );
  NOR2_X1 U4724 ( .A1(n3742), .A2(n5333), .ZN(n5798) );
  INV_X2 U4725 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n5069) );
  NAND2_X1 U4726 ( .A1(n6421), .A2(n5069), .ZN(n6425) );
  NAND2_X1 U4727 ( .A1(n3729), .A2(n6196), .ZN(n5270) );
  NAND2_X1 U4728 ( .A1(n3730), .A2(n4684), .ZN(n5335) );
  NAND2_X1 U4729 ( .A1(n4431), .A2(n5335), .ZN(n4364) );
  NAND2_X1 U4730 ( .A1(n4684), .A2(n4685), .ZN(n5334) );
  INV_X1 U4731 ( .A(n5334), .ZN(n5802) );
  AOI21_X1 U4732 ( .B1(n3731), .B2(n5798), .A(n5802), .ZN(n3732) );
  INV_X1 U4733 ( .A(n3732), .ZN(n3733) );
  AND2_X1 U4734 ( .A1(n3734), .A2(n3733), .ZN(n5782) );
  INV_X1 U4735 ( .A(n5786), .ZN(n3735) );
  NAND2_X1 U4736 ( .A1(n5271), .A2(n3735), .ZN(n3736) );
  AND2_X1 U4737 ( .A1(n5782), .A2(n3736), .ZN(n5776) );
  INV_X1 U4738 ( .A(n3744), .ZN(n3737) );
  OAI21_X1 U4739 ( .B1(n6244), .B2(n6236), .A(n3737), .ZN(n3738) );
  OAI21_X1 U4740 ( .B1(n5752), .B2(n5831), .A(n5767), .ZN(n5746) );
  AOI21_X1 U4741 ( .B1(n5735), .B2(n5271), .A(n5746), .ZN(n4280) );
  OAI21_X1 U4742 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5831), .A(n4280), 
        .ZN(n4265) );
  AOI21_X1 U4743 ( .B1(n4266), .B2(n5271), .A(n4265), .ZN(n3739) );
  INV_X1 U4744 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4432) );
  INV_X2 U4745 ( .A(n6196), .ZN(n6240) );
  NAND2_X1 U4746 ( .A1(n6240), .A2(REIP_REG_31__SCAN_IN), .ZN(n4302) );
  OAI21_X1 U4747 ( .B1(n3739), .B2(n4432), .A(n4302), .ZN(n3740) );
  AOI21_X1 U4748 ( .B1(n6237), .B2(n3741), .A(n3740), .ZN(n3746) );
  NAND2_X1 U4749 ( .A1(n5339), .A2(n6244), .ZN(n4689) );
  NAND2_X1 U4750 ( .A1(n5758), .A2(n5752), .ZN(n5743) );
  NOR3_X1 U4751 ( .A1(n5743), .A2(n4282), .A3(n5735), .ZN(n4267) );
  NAND3_X1 U4752 ( .A1(n4267), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n4432), .ZN(n3745) );
  OAI21_X1 U4753 ( .B1(n4305), .B2(n6184), .A(n3747), .ZN(U2987) );
  NAND2_X1 U4754 ( .A1(n4562), .A2(n3916), .ZN(n3748) );
  NAND2_X1 U4755 ( .A1(n5069), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3883) );
  NAND2_X1 U4756 ( .A1(n3748), .A2(n3883), .ZN(n3764) );
  NAND2_X1 U4757 ( .A1(n4563), .A2(n3916), .ZN(n3752) );
  AOI22_X1 U4758 ( .A1(n4227), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n5069), .ZN(n3750) );
  AND2_X1 U4759 ( .A1(n4327), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3775) );
  NAND2_X1 U4760 ( .A1(n3775), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3749) );
  AND2_X1 U4761 ( .A1(n3750), .A2(n3749), .ZN(n3751) );
  NAND2_X1 U4762 ( .A1(n3752), .A2(n3751), .ZN(n4482) );
  NAND2_X1 U4763 ( .A1(n3754), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4352) );
  INV_X1 U4764 ( .A(n3775), .ZN(n3771) );
  NAND2_X1 U4765 ( .A1(n3755), .A2(EAX_REG_0__SCAN_IN), .ZN(n3757) );
  NAND2_X1 U4766 ( .A1(n5069), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3756)
         );
  OAI211_X1 U4767 ( .C1(n3771), .C2(n5367), .A(n3757), .B(n3756), .ZN(n3758)
         );
  AOI21_X1 U4768 ( .B1(n5361), .B2(n3916), .A(n3758), .ZN(n3759) );
  INV_X1 U4769 ( .A(n3759), .ZN(n4354) );
  OR2_X1 U4770 ( .A1(n4354), .A2(n4233), .ZN(n3760) );
  NAND2_X1 U4771 ( .A1(n4353), .A2(n3760), .ZN(n4481) );
  INV_X1 U4772 ( .A(n3768), .ZN(n3761) );
  OAI21_X1 U4773 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3761), .ZN(n6169) );
  AOI22_X1 U4774 ( .A1(n3792), .A2(n6169), .B1(n4288), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3763) );
  NAND2_X1 U4775 ( .A1(n4227), .A2(EAX_REG_2__SCAN_IN), .ZN(n3762) );
  OAI211_X1 U4776 ( .C1(n3771), .C2(n3048), .A(n3763), .B(n3762), .ZN(n4397)
         );
  NAND2_X1 U4777 ( .A1(n4396), .A2(n4397), .ZN(n3766) );
  NAND2_X1 U4778 ( .A1(n3764), .A2(n4484), .ZN(n3765) );
  NAND2_X1 U4779 ( .A1(n3767), .A2(n3916), .ZN(n3774) );
  OAI21_X1 U4780 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3768), .A(n3777), 
        .ZN(n6160) );
  AOI22_X1 U4781 ( .A1(n3792), .A2(n6160), .B1(n4288), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3770) );
  NAND2_X1 U4782 ( .A1(n4227), .A2(EAX_REG_3__SCAN_IN), .ZN(n3769) );
  OAI211_X1 U4783 ( .C1(n3771), .C2(n3526), .A(n3770), .B(n3769), .ZN(n3772)
         );
  INV_X1 U4784 ( .A(n3772), .ZN(n3773) );
  NAND2_X1 U4785 ( .A1(n3774), .A2(n3773), .ZN(n4491) );
  NAND2_X1 U4786 ( .A1(n4394), .A2(n4491), .ZN(n4490) );
  NAND2_X1 U4787 ( .A1(n3775), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3781) );
  INV_X1 U4788 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6536) );
  AOI21_X1 U4789 ( .B1(n6536), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3776) );
  AOI21_X1 U4790 ( .B1(n4227), .B2(EAX_REG_4__SCAN_IN), .A(n3776), .ZN(n3780)
         );
  OAI21_X1 U4791 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3778), .A(n3790), 
        .ZN(n5164) );
  NOR2_X1 U4792 ( .A1(n5164), .A2(n4233), .ZN(n3779) );
  AOI21_X1 U4793 ( .B1(n3781), .B2(n3780), .A(n3779), .ZN(n3782) );
  AOI21_X1 U4794 ( .B1(n3783), .B2(n3916), .A(n3782), .ZN(n4501) );
  NAND2_X1 U4795 ( .A1(n3784), .A2(n3916), .ZN(n3787) );
  XNOR2_X1 U4796 ( .A(n3790), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5161) );
  INV_X1 U4797 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4598) );
  OAI22_X1 U4798 ( .A1(n5161), .A2(n4233), .B1(n3883), .B2(n4598), .ZN(n3785)
         );
  AOI21_X1 U4799 ( .B1(n4227), .B2(EAX_REG_5__SCAN_IN), .A(n3785), .ZN(n3786)
         );
  NAND2_X1 U4800 ( .A1(n3787), .A2(n3786), .ZN(n4496) );
  NAND2_X1 U4801 ( .A1(n4493), .A2(n4496), .ZN(n4494) );
  INV_X1 U4802 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4579) );
  INV_X1 U4803 ( .A(n3790), .ZN(n3788) );
  AOI21_X1 U4804 ( .B1(n3788), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3791) );
  NAND2_X1 U4805 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3789) );
  OR2_X1 U4806 ( .A1(n3791), .A2(n3797), .ZN(n6152) );
  AOI22_X1 U4807 ( .A1(n6152), .A2(n3792), .B1(n4288), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3793) );
  OAI21_X1 U4808 ( .B1(n3984), .B2(n4579), .A(n3793), .ZN(n3794) );
  INV_X1 U4809 ( .A(n4576), .ZN(n3796) );
  INV_X1 U4810 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4703) );
  NOR2_X1 U4811 ( .A1(n3797), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3798)
         );
  OR2_X1 U4812 ( .A1(n3818), .A2(n3798), .ZN(n4989) );
  INV_X1 U4813 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6628) );
  NOR2_X1 U4814 ( .A1(n3883), .A2(n6628), .ZN(n3799) );
  AOI21_X1 U4815 ( .B1(n4989), .B2(n3792), .A(n3799), .ZN(n3800) );
  OAI21_X1 U4816 ( .B1(n3984), .B2(n4703), .A(n3800), .ZN(n3801) );
  AOI22_X1 U4817 ( .A1(n4173), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4818 ( .A1(n3253), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4532), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4819 ( .A1(n4215), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4820 ( .A1(n3803), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3804) );
  NAND4_X1 U4821 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3813)
         );
  AOI22_X1 U4822 ( .A1(n4208), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4823 ( .A1(n4150), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4824 ( .A1(n3425), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4825 ( .A1(n4195), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3808) );
  NAND4_X1 U4826 ( .A1(n3811), .A2(n3810), .A3(n3809), .A4(n3808), .ZN(n3812)
         );
  OAI21_X1 U4827 ( .B1(n3813), .B2(n3812), .A(n3916), .ZN(n3817) );
  NAND2_X1 U4828 ( .A1(n4227), .A2(EAX_REG_8__SCAN_IN), .ZN(n3816) );
  NAND2_X1 U4829 ( .A1(n4288), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3815)
         );
  XNOR2_X1 U4830 ( .A(n3818), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U4831 ( .A1(n5192), .A2(n3792), .ZN(n3814) );
  NAND4_X1 U4832 ( .A1(n3817), .A2(n3816), .A3(n3815), .A4(n3814), .ZN(n4643)
         );
  INV_X1 U4833 ( .A(n4642), .ZN(n3833) );
  XOR2_X1 U4834 ( .A(n6018), .B(n3834), .Z(n6022) );
  AOI22_X1 U4835 ( .A1(n4227), .A2(EAX_REG_9__SCAN_IN), .B1(n4288), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4836 ( .A1(n4208), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4837 ( .A1(n4215), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4838 ( .A1(n3253), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4839 ( .A1(n3803), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3820) );
  NAND4_X1 U4840 ( .A1(n3823), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3829)
         );
  AOI22_X1 U4841 ( .A1(n4174), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4842 ( .A1(n3425), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4532), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4843 ( .A1(n4216), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4844 ( .A1(n4195), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3824) );
  NAND4_X1 U4845 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3828)
         );
  OAI21_X1 U4846 ( .B1(n3829), .B2(n3828), .A(n3916), .ZN(n3830) );
  OAI211_X1 U4847 ( .C1(n6022), .C2(n4233), .A(n3831), .B(n3830), .ZN(n3832)
         );
  INV_X1 U4848 ( .A(n3832), .ZN(n5013) );
  NAND2_X1 U4849 ( .A1(n3833), .A2(n3832), .ZN(n5012) );
  INV_X1 U4850 ( .A(n5012), .ZN(n3850) );
  XNOR2_X1 U4851 ( .A(n3851), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5265)
         );
  AOI22_X1 U4852 ( .A1(n4150), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4853 ( .A1(n4208), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4854 ( .A1(n4195), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4855 ( .A1(n3803), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3835) );
  NAND4_X1 U4856 ( .A1(n3838), .A2(n3837), .A3(n3836), .A4(n3835), .ZN(n3844)
         );
  AOI22_X1 U4857 ( .A1(n4174), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4858 ( .A1(n3425), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4859 ( .A1(n4215), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4860 ( .A1(n4532), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3839) );
  NAND4_X1 U4861 ( .A1(n3842), .A2(n3841), .A3(n3840), .A4(n3839), .ZN(n3843)
         );
  OAI21_X1 U4862 ( .B1(n3844), .B2(n3843), .A(n3916), .ZN(n3847) );
  NAND2_X1 U4863 ( .A1(n4227), .A2(EAX_REG_10__SCAN_IN), .ZN(n3846) );
  NAND2_X1 U4864 ( .A1(n4288), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3845)
         );
  NAND3_X1 U4865 ( .A1(n3847), .A2(n3846), .A3(n3845), .ZN(n3848) );
  AOI21_X1 U4866 ( .B1(n5265), .B2(n3792), .A(n3848), .ZN(n5140) );
  XOR2_X1 U4867 ( .A(n3865), .B(n3866), .Z(n5999) );
  AOI22_X1 U4868 ( .A1(n4227), .A2(EAX_REG_11__SCAN_IN), .B1(n4288), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4869 ( .A1(n4174), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4870 ( .A1(n4216), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4871 ( .A1(n4215), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4872 ( .A1(n3803), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3852) );
  NAND4_X1 U4873 ( .A1(n3855), .A2(n3854), .A3(n3853), .A4(n3852), .ZN(n3861)
         );
  AOI22_X1 U4874 ( .A1(n4208), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4875 ( .A1(n4173), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4876 ( .A1(n4195), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4532), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4877 ( .A1(n3290), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3856) );
  NAND4_X1 U4878 ( .A1(n3859), .A2(n3858), .A3(n3857), .A4(n3856), .ZN(n3860)
         );
  OAI21_X1 U4879 ( .B1(n3861), .B2(n3860), .A(n3916), .ZN(n3862) );
  OAI211_X1 U4880 ( .C1(n5999), .C2(n4233), .A(n3863), .B(n3862), .ZN(n3864)
         );
  AOI22_X1 U4881 ( .A1(n4227), .A2(EAX_REG_12__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n5069), .ZN(n3879) );
  XNOR2_X1 U4882 ( .A(n3880), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5303)
         );
  NAND2_X1 U4883 ( .A1(n5303), .A2(n3792), .ZN(n3878) );
  AOI22_X1 U4884 ( .A1(n4215), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4885 ( .A1(n4150), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4886 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n3253), .B1(n4532), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4887 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n3803), .B1(n3290), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3867) );
  NAND4_X1 U4888 ( .A1(n3870), .A2(n3869), .A3(n3868), .A4(n3867), .ZN(n3876)
         );
  AOI22_X1 U4889 ( .A1(n4216), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4890 ( .A1(n4208), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4891 ( .A1(n3425), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4892 ( .A1(n4195), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3871) );
  NAND4_X1 U4893 ( .A1(n3874), .A2(n3873), .A3(n3872), .A4(n3871), .ZN(n3875)
         );
  OAI21_X1 U4894 ( .B1(n3876), .B2(n3875), .A(n3916), .ZN(n3877) );
  OAI211_X1 U4895 ( .C1(n3792), .C2(n3879), .A(n3878), .B(n3877), .ZN(n5282)
         );
  INV_X1 U4896 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3884) );
  OAI21_X1 U4897 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3881), .A(n3927), 
        .ZN(n5998) );
  NAND2_X1 U4898 ( .A1(n5998), .A2(n3792), .ZN(n3882) );
  OAI21_X1 U4899 ( .B1(n3884), .B2(n3883), .A(n3882), .ZN(n3885) );
  AOI21_X1 U4900 ( .B1(n4227), .B2(EAX_REG_13__SCAN_IN), .A(n3885), .ZN(n3886)
         );
  OR2_X2 U4901 ( .A1(n3887), .A2(n3886), .ZN(n5313) );
  NAND2_X1 U4902 ( .A1(n5313), .A2(n3888), .ZN(n5310) );
  INV_X1 U4903 ( .A(n5310), .ZN(n3901) );
  AOI22_X1 U4904 ( .A1(n4208), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4905 ( .A1(n4173), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4906 ( .A1(n4195), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4907 ( .A1(n3803), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3889) );
  NAND4_X1 U4908 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(n3898)
         );
  AOI22_X1 U4909 ( .A1(n4174), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4910 ( .A1(n4150), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4911 ( .A1(n4215), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4912 ( .A1(n4532), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3893) );
  NAND4_X1 U4913 ( .A1(n3896), .A2(n3895), .A3(n3894), .A4(n3893), .ZN(n3897)
         );
  OR2_X1 U4914 ( .A1(n3898), .A2(n3897), .ZN(n3899) );
  NAND2_X1 U4915 ( .A1(n3916), .A2(n3899), .ZN(n5309) );
  INV_X1 U4916 ( .A(n5309), .ZN(n3900) );
  NAND2_X1 U4917 ( .A1(n3901), .A2(n3900), .ZN(n5308) );
  AOI22_X1 U4918 ( .A1(n4216), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4919 ( .A1(n4150), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4920 ( .A1(n4195), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3803), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4921 ( .A1(n4532), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3902) );
  NAND4_X1 U4922 ( .A1(n3905), .A2(n3904), .A3(n3903), .A4(n3902), .ZN(n3911)
         );
  AOI22_X1 U4923 ( .A1(n4208), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4924 ( .A1(n3425), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4925 ( .A1(n4215), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4926 ( .A1(n3290), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3906) );
  NAND4_X1 U4927 ( .A1(n3909), .A2(n3908), .A3(n3907), .A4(n3906), .ZN(n3910)
         );
  OAI21_X1 U4928 ( .B1(n3911), .B2(n3910), .A(n3916), .ZN(n3915) );
  INV_X1 U4929 ( .A(n3936), .ZN(n3912) );
  XNOR2_X1 U4930 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3912), .ZN(n5982)
         );
  AOI22_X1 U4931 ( .A1(n3792), .A2(n5982), .B1(n4288), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3914) );
  NAND2_X1 U4932 ( .A1(n4227), .A2(EAX_REG_15__SCAN_IN), .ZN(n3913) );
  INV_X1 U4933 ( .A(n5353), .ZN(n3934) );
  INV_X1 U4934 ( .A(n3916), .ZN(n3933) );
  AOI22_X1 U4935 ( .A1(n4174), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4936 ( .A1(n3425), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4937 ( .A1(n3261), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4938 ( .A1(n4195), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3917) );
  NAND4_X1 U4939 ( .A1(n3920), .A2(n3919), .A3(n3918), .A4(n3917), .ZN(n3926)
         );
  AOI22_X1 U4940 ( .A1(n4150), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4941 ( .A1(n4208), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4215), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4942 ( .A1(n4532), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4943 ( .A1(n3803), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3921) );
  NAND4_X1 U4944 ( .A1(n3924), .A2(n3923), .A3(n3922), .A4(n3921), .ZN(n3925)
         );
  NOR2_X1 U4945 ( .A1(n3926), .A2(n3925), .ZN(n3932) );
  XOR2_X1 U4946 ( .A(n3928), .B(n3927), .Z(n5727) );
  INV_X1 U4947 ( .A(n5727), .ZN(n3929) );
  AOI22_X1 U4948 ( .A1(n4288), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n3792), 
        .B2(n3929), .ZN(n3931) );
  NAND2_X1 U4949 ( .A1(n4227), .A2(EAX_REG_14__SCAN_IN), .ZN(n3930) );
  OAI211_X1 U4950 ( .C1(n3933), .C2(n3932), .A(n3931), .B(n3930), .ZN(n5314)
         );
  XOR2_X1 U4951 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3951), .Z(n5715) );
  AOI22_X1 U4952 ( .A1(n4208), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4953 ( .A1(n4150), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4954 ( .A1(n4195), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4532), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3938) );
  AOI22_X1 U4955 ( .A1(n3803), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3937) );
  NAND4_X1 U4956 ( .A1(n3940), .A2(n3939), .A3(n3938), .A4(n3937), .ZN(n3946)
         );
  AOI22_X1 U4957 ( .A1(n4174), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4958 ( .A1(n4173), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4959 ( .A1(n4215), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4960 ( .A1(n3289), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3941) );
  NAND4_X1 U4961 ( .A1(n3944), .A2(n3943), .A3(n3942), .A4(n3941), .ZN(n3945)
         );
  NOR2_X1 U4962 ( .A1(n3946), .A2(n3945), .ZN(n3948) );
  AOI22_X1 U4963 ( .A1(n4227), .A2(EAX_REG_16__SCAN_IN), .B1(n4288), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3947) );
  OAI21_X1 U4964 ( .B1(n4230), .B2(n3948), .A(n3947), .ZN(n3949) );
  INV_X1 U4965 ( .A(n3949), .ZN(n3950) );
  OAI21_X1 U4966 ( .B1(n5715), .B2(n4233), .A(n3950), .ZN(n5515) );
  XNOR2_X1 U4967 ( .A(n3968), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5705)
         );
  NAND2_X1 U4968 ( .A1(n5705), .A2(n3792), .ZN(n3967) );
  AOI22_X1 U4969 ( .A1(n4173), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4215), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4970 ( .A1(n4195), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4971 ( .A1(n3425), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3803), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4972 ( .A1(n3261), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3952) );
  NAND4_X1 U4973 ( .A1(n3955), .A2(n3954), .A3(n3953), .A4(n3952), .ZN(n3963)
         );
  AOI22_X1 U4974 ( .A1(n4216), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4532), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3961) );
  NAND2_X1 U4975 ( .A1(n4208), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3957) );
  NAND2_X1 U4976 ( .A1(n3290), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3956) );
  AND3_X1 U4977 ( .A1(n3957), .A2(n4233), .A3(n3956), .ZN(n3960) );
  AOI22_X1 U4978 ( .A1(n4174), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4979 ( .A1(n3179), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3181), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3958) );
  NAND4_X1 U4980 ( .A1(n3961), .A2(n3960), .A3(n3959), .A4(n3958), .ZN(n3962)
         );
  NAND2_X1 U4981 ( .A1(n4230), .A2(n4233), .ZN(n4033) );
  OAI21_X1 U4982 ( .B1(n3963), .B2(n3962), .A(n4033), .ZN(n3965) );
  AOI22_X1 U4983 ( .A1(n4227), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n5069), .ZN(n3964) );
  NAND2_X1 U4984 ( .A1(n3965), .A2(n3964), .ZN(n3966) );
  INV_X1 U4985 ( .A(n5505), .ZN(n3988) );
  OR2_X1 U4986 ( .A1(n3969), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3970)
         );
  NAND2_X1 U4987 ( .A1(n4005), .A2(n3970), .ZN(n5975) );
  AOI22_X1 U4988 ( .A1(n4208), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4150), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4989 ( .A1(n4173), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4990 ( .A1(n3261), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4991 ( .A1(n4532), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3971) );
  NAND4_X1 U4992 ( .A1(n3974), .A2(n3973), .A3(n3972), .A4(n3971), .ZN(n3980)
         );
  AOI22_X1 U4993 ( .A1(n4174), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4994 ( .A1(n4216), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4215), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4995 ( .A1(n4195), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3181), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4996 ( .A1(n3803), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3975) );
  NAND4_X1 U4997 ( .A1(n3978), .A2(n3977), .A3(n3976), .A4(n3975), .ZN(n3979)
         );
  NOR2_X1 U4998 ( .A1(n3980), .A2(n3979), .ZN(n3981) );
  NOR2_X1 U4999 ( .A1(n4230), .A2(n3981), .ZN(n3986) );
  INV_X1 U5000 ( .A(EAX_REG_18__SCAN_IN), .ZN(n3983) );
  NAND2_X1 U5001 ( .A1(n5069), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3982)
         );
  OAI211_X1 U5002 ( .C1(n3984), .C2(n3983), .A(n4233), .B(n3982), .ZN(n3985)
         );
  OAI22_X1 U5003 ( .A1(n5975), .A2(n4233), .B1(n3986), .B2(n3985), .ZN(n5566)
         );
  NAND2_X1 U5004 ( .A1(n3988), .A2(n3987), .ZN(n5488) );
  XNOR2_X1 U5005 ( .A(n4005), .B(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5687)
         );
  NAND2_X1 U5006 ( .A1(n5687), .A2(n3792), .ZN(n4004) );
  AOI22_X1 U5007 ( .A1(n4208), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U5008 ( .A1(n4150), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4532), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U5009 ( .A1(n3179), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3803), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U5010 ( .A1(n4215), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3989) );
  NAND4_X1 U5011 ( .A1(n3992), .A2(n3991), .A3(n3990), .A4(n3989), .ZN(n4000)
         );
  AOI22_X1 U5012 ( .A1(n4195), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3998) );
  NAND2_X1 U5013 ( .A1(n4216), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3994) );
  NAND2_X1 U5014 ( .A1(n4210), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3993) );
  AND3_X1 U5015 ( .A1(n3994), .A2(n4233), .A3(n3993), .ZN(n3997) );
  AOI22_X1 U5016 ( .A1(n4173), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U5017 ( .A1(n3425), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3995) );
  NAND4_X1 U5018 ( .A1(n3998), .A2(n3997), .A3(n3996), .A4(n3995), .ZN(n3999)
         );
  OAI21_X1 U5019 ( .B1(n4000), .B2(n3999), .A(n4033), .ZN(n4002) );
  AOI22_X1 U5020 ( .A1(n4227), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n5069), .ZN(n4001) );
  NAND2_X1 U5021 ( .A1(n4002), .A2(n4001), .ZN(n4003) );
  NAND2_X1 U5022 ( .A1(n4004), .A2(n4003), .ZN(n5487) );
  AND2_X1 U5023 ( .A1(n4006), .A2(n5678), .ZN(n4007) );
  OR2_X1 U5024 ( .A1(n4007), .A2(n4038), .ZN(n5910) );
  AOI22_X1 U5025 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n4216), .B1(n3253), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U5026 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n4195), .B1(n3425), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U5027 ( .A1(n4208), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U5028 ( .A1(n4215), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4008) );
  NAND4_X1 U5029 ( .A1(n4011), .A2(n4010), .A3(n4009), .A4(n4008), .ZN(n4017)
         );
  AOI22_X1 U5030 ( .A1(n4150), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U5031 ( .A1(n4174), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4532), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U5032 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3290), .B1(n3289), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U5033 ( .A1(n3803), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4012) );
  NAND4_X1 U5034 ( .A1(n4015), .A2(n4014), .A3(n4013), .A4(n4012), .ZN(n4016)
         );
  NOR2_X1 U5035 ( .A1(n4017), .A2(n4016), .ZN(n4020) );
  OAI21_X1 U5036 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6424), .A(n5069), 
        .ZN(n4019) );
  NAND2_X1 U5037 ( .A1(n4227), .A2(EAX_REG_20__SCAN_IN), .ZN(n4018) );
  OAI211_X1 U5038 ( .C1(n4230), .C2(n4020), .A(n4019), .B(n4018), .ZN(n4021)
         );
  OAI21_X1 U5039 ( .B1(n5910), .B2(n4233), .A(n4021), .ZN(n5559) );
  INV_X1 U5040 ( .A(n5559), .ZN(n4022) );
  INV_X1 U5041 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5672) );
  XNOR2_X1 U5042 ( .A(n4038), .B(n5672), .ZN(n5894) );
  AOI22_X1 U5043 ( .A1(n4227), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n5069), .ZN(n4037) );
  AOI22_X1 U5044 ( .A1(n4195), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3803), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U5045 ( .A1(n4150), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3181), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U5046 ( .A1(n3425), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U5047 ( .A1(n4215), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4023) );
  NAND4_X1 U5048 ( .A1(n4026), .A2(n4025), .A3(n4024), .A4(n4023), .ZN(n4035)
         );
  NAND2_X1 U5049 ( .A1(n4174), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4028)
         );
  NAND2_X1 U5050 ( .A1(n4532), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4027)
         );
  AND3_X1 U5051 ( .A1(n4028), .A2(n4027), .A3(n4233), .ZN(n4032) );
  AOI22_X1 U5052 ( .A1(n4216), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U5053 ( .A1(n4173), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U5054 ( .A1(n4208), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4029) );
  NAND4_X1 U5055 ( .A1(n4032), .A2(n4031), .A3(n4030), .A4(n4029), .ZN(n4034)
         );
  OAI21_X1 U5056 ( .B1(n4035), .B2(n4034), .A(n4033), .ZN(n4036) );
  AOI22_X1 U5057 ( .A1(n5894), .A2(n3792), .B1(n4037), .B2(n4036), .ZN(n5554)
         );
  OR2_X1 U5058 ( .A1(n4039), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4040)
         );
  NAND2_X1 U5059 ( .A1(n4085), .A2(n4040), .ZN(n5882) );
  AOI22_X1 U5060 ( .A1(n4208), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U5061 ( .A1(n4173), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5062 ( .A1(n4215), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U5063 ( .A1(n3803), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4041) );
  NAND4_X1 U5064 ( .A1(n4044), .A2(n4043), .A3(n4042), .A4(n4041), .ZN(n4050)
         );
  AOI22_X1 U5065 ( .A1(n4174), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U5066 ( .A1(n3819), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U5067 ( .A1(n4532), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3181), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U5068 ( .A1(n3183), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4045) );
  NAND4_X1 U5069 ( .A1(n4048), .A2(n4047), .A3(n4046), .A4(n4045), .ZN(n4049)
         );
  NOR2_X1 U5070 ( .A1(n4050), .A2(n4049), .ZN(n4054) );
  NAND2_X1 U5071 ( .A1(n5069), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4051)
         );
  NAND2_X1 U5072 ( .A1(n4233), .A2(n4051), .ZN(n4052) );
  AOI21_X1 U5073 ( .B1(n4227), .B2(EAX_REG_22__SCAN_IN), .A(n4052), .ZN(n4053)
         );
  OAI21_X1 U5074 ( .B1(n4230), .B2(n4054), .A(n4053), .ZN(n4055) );
  NAND2_X1 U5075 ( .A1(n4056), .A2(n4055), .ZN(n5547) );
  INV_X1 U5076 ( .A(n5547), .ZN(n4057) );
  XNOR2_X1 U5078 ( .A(n4085), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5662)
         );
  NAND2_X1 U5079 ( .A1(n5662), .A2(n3792), .ZN(n4082) );
  AOI22_X1 U5080 ( .A1(n4150), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U5081 ( .A1(n4174), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5082 ( .A1(n4208), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U5083 ( .A1(n4215), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4058) );
  NAND4_X1 U5084 ( .A1(n4061), .A2(n4060), .A3(n4059), .A4(n4058), .ZN(n4067)
         );
  AOI22_X1 U5085 ( .A1(n3425), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U5086 ( .A1(n4532), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5087 ( .A1(n4195), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U5088 ( .A1(n3803), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4062) );
  NAND4_X1 U5089 ( .A1(n4065), .A2(n4064), .A3(n4063), .A4(n4062), .ZN(n4066)
         );
  NOR2_X1 U5090 ( .A1(n4067), .A2(n4066), .ZN(n4089) );
  AOI22_X1 U5091 ( .A1(n3425), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U5092 ( .A1(n4174), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4215), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U5093 ( .A1(n4195), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U5094 ( .A1(n3290), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4068) );
  NAND4_X1 U5095 ( .A1(n4071), .A2(n4070), .A3(n4069), .A4(n4068), .ZN(n4077)
         );
  AOI22_X1 U5096 ( .A1(n4208), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4075) );
  AOI22_X1 U5097 ( .A1(n4150), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4074) );
  AOI22_X1 U5098 ( .A1(n4532), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3803), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U5099 ( .A1(n3261), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4072) );
  NAND4_X1 U5100 ( .A1(n4075), .A2(n4074), .A3(n4073), .A4(n4072), .ZN(n4076)
         );
  NOR2_X1 U5101 ( .A1(n4077), .A2(n4076), .ZN(n4088) );
  XNOR2_X1 U5102 ( .A(n4089), .B(n4088), .ZN(n4080) );
  INV_X1 U5103 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5658) );
  AOI21_X1 U5104 ( .B1(n5658), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4078) );
  AOI21_X1 U5105 ( .B1(n4227), .B2(EAX_REG_23__SCAN_IN), .A(n4078), .ZN(n4079)
         );
  OAI21_X1 U5106 ( .B1(n4230), .B2(n4080), .A(n4079), .ZN(n4081) );
  NAND2_X1 U5107 ( .A1(n4082), .A2(n4081), .ZN(n5476) );
  NAND2_X1 U5108 ( .A1(n5546), .A2(n4083), .ZN(n5474) );
  INV_X1 U5109 ( .A(n4086), .ZN(n4087) );
  INV_X1 U5110 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5869) );
  OAI21_X1 U5111 ( .B1(n4087), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n4120), 
        .ZN(n5868) );
  OR2_X1 U5112 ( .A1(n4089), .A2(n4088), .ZN(n4105) );
  AOI22_X1 U5113 ( .A1(n4174), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4093) );
  AOI22_X1 U5114 ( .A1(n4215), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4092) );
  AOI22_X1 U5115 ( .A1(n3819), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U5116 ( .A1(n4216), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4090) );
  NAND4_X1 U5117 ( .A1(n4093), .A2(n4092), .A3(n4091), .A4(n4090), .ZN(n4099)
         );
  AOI22_X1 U5118 ( .A1(n4195), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4097) );
  AOI22_X1 U5119 ( .A1(n4208), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3803), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4096) );
  AOI22_X1 U5120 ( .A1(n3425), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4095) );
  AOI22_X1 U5121 ( .A1(n4532), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4094) );
  NAND4_X1 U5122 ( .A1(n4097), .A2(n4096), .A3(n4095), .A4(n4094), .ZN(n4098)
         );
  NOR2_X1 U5123 ( .A1(n4099), .A2(n4098), .ZN(n4104) );
  XNOR2_X1 U5124 ( .A(n4105), .B(n4104), .ZN(n4101) );
  AOI22_X1 U5125 ( .A1(n4227), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n4288), .ZN(n4100) );
  OAI21_X1 U5126 ( .B1(n4230), .B2(n4101), .A(n4100), .ZN(n4102) );
  AOI21_X1 U5127 ( .B1(n5868), .B2(n3792), .A(n4102), .ZN(n5537) );
  XNOR2_X1 U5128 ( .A(n4120), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5639)
         );
  INV_X1 U5129 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5637) );
  NOR2_X1 U5130 ( .A1(n5637), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4103) );
  AOI211_X1 U5131 ( .C1(n3755), .C2(EAX_REG_25__SCAN_IN), .A(n3792), .B(n4103), 
        .ZN(n4119) );
  AOI22_X1 U5132 ( .A1(n4173), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4110) );
  AOI22_X1 U5133 ( .A1(n4208), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4215), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5134 ( .A1(n4532), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U5135 ( .A1(n3290), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4107) );
  NAND4_X1 U5136 ( .A1(n4110), .A2(n4109), .A3(n4108), .A4(n4107), .ZN(n4116)
         );
  AOI22_X1 U5137 ( .A1(n4150), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4114) );
  AOI22_X1 U5138 ( .A1(n4174), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U5139 ( .A1(n4195), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3803), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4112) );
  AOI22_X1 U5140 ( .A1(n3261), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4111) );
  NAND4_X1 U5141 ( .A1(n4114), .A2(n4113), .A3(n4112), .A4(n4111), .ZN(n4115)
         );
  NOR2_X1 U5142 ( .A1(n4116), .A2(n4115), .ZN(n4126) );
  XOR2_X1 U5143 ( .A(n4125), .B(n4126), .Z(n4117) );
  INV_X1 U5144 ( .A(n4230), .ZN(n4202) );
  NAND2_X1 U5145 ( .A1(n4117), .A2(n4202), .ZN(n4118) );
  AOI22_X1 U5146 ( .A1(n5639), .A2(n3792), .B1(n4119), .B2(n4118), .ZN(n5463)
         );
  INV_X1 U5147 ( .A(n4121), .ZN(n4123) );
  INV_X1 U5148 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4122) );
  NAND2_X1 U5149 ( .A1(n4123), .A2(n4122), .ZN(n4124) );
  NAND2_X1 U5150 ( .A1(n4160), .A2(n4124), .ZN(n5633) );
  NOR2_X1 U5151 ( .A1(n4126), .A2(n4125), .ZN(n4145) );
  NOR2_X1 U5152 ( .A1(n4169), .A2(n4127), .ZN(n4130) );
  INV_X1 U5153 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4728) );
  INV_X1 U5154 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4128) );
  OAI22_X1 U5155 ( .A1(n3252), .A2(n4728), .B1(n2960), .B2(n4128), .ZN(n4129)
         );
  AOI211_X1 U5156 ( .C1(INSTQUEUE_REG_11__3__SCAN_IN), .C2(n4532), .A(n4130), 
        .B(n4129), .ZN(n4138) );
  AOI22_X1 U5157 ( .A1(n4150), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U5158 ( .A1(n4174), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U5159 ( .A1(n4208), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U5160 ( .A1(n4215), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4131) );
  AND4_X1 U5161 ( .A1(n4134), .A2(n4133), .A3(n4132), .A4(n4131), .ZN(n4137)
         );
  AOI22_X1 U5162 ( .A1(n4195), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U5163 ( .A1(n3803), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4135) );
  NAND4_X1 U5164 ( .A1(n4138), .A2(n4137), .A3(n4136), .A4(n4135), .ZN(n4144)
         );
  XNOR2_X1 U5165 ( .A(n4145), .B(n4144), .ZN(n4141) );
  AOI21_X1 U5166 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n5069), .A(n3792), 
        .ZN(n4140) );
  NAND2_X1 U5167 ( .A1(n4227), .A2(EAX_REG_26__SCAN_IN), .ZN(n4139) );
  OAI211_X1 U5168 ( .C1(n4141), .C2(n4230), .A(n4140), .B(n4139), .ZN(n4142)
         );
  OAI21_X1 U5169 ( .B1(n5633), .B2(n4233), .A(n4142), .ZN(n5450) );
  XNOR2_X1 U5170 ( .A(n4160), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5629)
         );
  INV_X1 U5171 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5625) );
  NOR2_X1 U5172 ( .A1(n5625), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4143) );
  AOI211_X1 U5173 ( .C1(n3755), .C2(EAX_REG_27__SCAN_IN), .A(n3792), .B(n4143), 
        .ZN(n4159) );
  NAND2_X1 U5174 ( .A1(n4145), .A2(n4144), .ZN(n4166) );
  AOI22_X1 U5175 ( .A1(n4174), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U5176 ( .A1(n4215), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U5177 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4532), .B1(n3289), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4147) );
  AOI22_X1 U5178 ( .A1(n3803), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4146) );
  NAND4_X1 U5179 ( .A1(n4149), .A2(n4148), .A3(n4147), .A4(n4146), .ZN(n4156)
         );
  AOI22_X1 U5180 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4216), .B1(n4150), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5181 ( .A1(n4173), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U5182 ( .A1(n4208), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4152) );
  AOI22_X1 U5183 ( .A1(n4195), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4151) );
  NAND4_X1 U5184 ( .A1(n4154), .A2(n4153), .A3(n4152), .A4(n4151), .ZN(n4155)
         );
  NOR2_X1 U5185 ( .A1(n4156), .A2(n4155), .ZN(n4167) );
  XOR2_X1 U5186 ( .A(n4166), .B(n4167), .Z(n4157) );
  NAND2_X1 U5187 ( .A1(n4157), .A2(n4202), .ZN(n4158) );
  AOI22_X1 U5188 ( .A1(n5629), .A2(n3792), .B1(n4159), .B2(n4158), .ZN(n5438)
         );
  INV_X1 U5189 ( .A(n4160), .ZN(n4161) );
  INV_X1 U5190 ( .A(n4162), .ZN(n4164) );
  INV_X1 U5191 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4163) );
  NAND2_X1 U5192 ( .A1(n4164), .A2(n4163), .ZN(n4165) );
  NAND2_X1 U5193 ( .A1(n4206), .A2(n4165), .ZN(n5618) );
  NOR2_X1 U5194 ( .A1(n4167), .A2(n4166), .ZN(n4190) );
  NOR2_X1 U5195 ( .A1(n4169), .A2(n4168), .ZN(n4172) );
  INV_X1 U5196 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4719) );
  INV_X1 U5197 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4170) );
  OAI22_X1 U5198 ( .A1(n3252), .A2(n4719), .B1(n2960), .B2(n4170), .ZN(n4171)
         );
  AOI211_X1 U5199 ( .C1(INSTQUEUE_REG_11__5__SCAN_IN), .C2(n4532), .A(n4172), 
        .B(n4171), .ZN(n4182) );
  AOI22_X1 U5200 ( .A1(n4150), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4178) );
  AOI22_X1 U5201 ( .A1(n4174), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4177) );
  AOI22_X1 U5202 ( .A1(n4208), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4176) );
  AOI22_X1 U5203 ( .A1(n4215), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4175) );
  AND4_X1 U5204 ( .A1(n4178), .A2(n4177), .A3(n4176), .A4(n4175), .ZN(n4181)
         );
  AOI22_X1 U5205 ( .A1(n4195), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4180) );
  AOI22_X1 U5206 ( .A1(n3803), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4179) );
  NAND4_X1 U5207 ( .A1(n4182), .A2(n4181), .A3(n4180), .A4(n4179), .ZN(n4189)
         );
  XNOR2_X1 U5208 ( .A(n4190), .B(n4189), .ZN(n4185) );
  AOI21_X1 U5209 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n5069), .A(n3792), 
        .ZN(n4184) );
  NAND2_X1 U5210 ( .A1(n4227), .A2(EAX_REG_28__SCAN_IN), .ZN(n4183) );
  OAI211_X1 U5211 ( .C1(n4185), .C2(n4230), .A(n4184), .B(n4183), .ZN(n4186)
         );
  OAI21_X1 U5212 ( .B1(n5618), .B2(n4233), .A(n4186), .ZN(n5424) );
  XNOR2_X1 U5213 ( .A(n4206), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5420)
         );
  INV_X1 U5214 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4187) );
  AOI21_X1 U5215 ( .B1(n4187), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4188) );
  AOI21_X1 U5216 ( .B1(n3755), .B2(EAX_REG_29__SCAN_IN), .A(n4188), .ZN(n4205)
         );
  NAND2_X1 U5217 ( .A1(n4190), .A2(n4189), .ZN(n4223) );
  AOI22_X1 U5218 ( .A1(n4174), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3253), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4194) );
  AOI22_X1 U5219 ( .A1(n4173), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4193) );
  AOI22_X1 U5220 ( .A1(n4532), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3181), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4192) );
  AOI22_X1 U5221 ( .A1(n3803), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4191) );
  NAND4_X1 U5222 ( .A1(n4194), .A2(n4193), .A3(n4192), .A4(n4191), .ZN(n4201)
         );
  AOI22_X1 U5223 ( .A1(n4208), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4216), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4199) );
  AOI22_X1 U5224 ( .A1(n4150), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4198) );
  AOI22_X1 U5225 ( .A1(n4215), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3261), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4197) );
  AOI22_X1 U5226 ( .A1(n4195), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4196) );
  NAND4_X1 U5227 ( .A1(n4199), .A2(n4198), .A3(n4197), .A4(n4196), .ZN(n4200)
         );
  NOR2_X1 U5228 ( .A1(n4201), .A2(n4200), .ZN(n4224) );
  XOR2_X1 U5229 ( .A(n4223), .B(n4224), .Z(n4203) );
  NAND2_X1 U5230 ( .A1(n4203), .A2(n4202), .ZN(n4204) );
  AOI22_X1 U5231 ( .A1(n5420), .A2(n3792), .B1(n4205), .B2(n4204), .ZN(n4309)
         );
  XOR2_X1 U5232 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .B(n4293), .Z(n5606) );
  AOI22_X1 U5233 ( .A1(n4208), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4173), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4214) );
  AOI22_X1 U5234 ( .A1(n3425), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3179), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4213) );
  AOI22_X1 U5235 ( .A1(n3261), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4209), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4212) );
  AOI22_X1 U5236 ( .A1(n3183), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4210), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4211) );
  NAND4_X1 U5237 ( .A1(n4214), .A2(n4213), .A3(n4212), .A4(n4211), .ZN(n4222)
         );
  AOI22_X1 U5238 ( .A1(n3819), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4174), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U5239 ( .A1(n4216), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4215), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4219) );
  AOI22_X1 U5240 ( .A1(n4532), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3181), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4218) );
  AOI22_X1 U5241 ( .A1(n3803), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4217) );
  NAND4_X1 U5242 ( .A1(n4220), .A2(n4219), .A3(n4218), .A4(n4217), .ZN(n4221)
         );
  NOR2_X1 U5243 ( .A1(n4222), .A2(n4221), .ZN(n4226) );
  NOR2_X1 U5244 ( .A1(n4224), .A2(n4223), .ZN(n4225) );
  XOR2_X1 U5245 ( .A(n4226), .B(n4225), .Z(n4231) );
  AOI21_X1 U5246 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n5069), .A(n3792), 
        .ZN(n4229) );
  NAND2_X1 U5247 ( .A1(n4227), .A2(EAX_REG_30__SCAN_IN), .ZN(n4228) );
  OAI211_X1 U5248 ( .C1(n4231), .C2(n4230), .A(n4229), .B(n4228), .ZN(n4232)
         );
  OAI21_X1 U5249 ( .B1(n5606), .B2(n4233), .A(n4232), .ZN(n4235) );
  INV_X1 U5250 ( .A(n4290), .ZN(n4237) );
  NAND2_X1 U5251 ( .A1(n4308), .A2(n4235), .ZN(n4236) );
  NAND2_X1 U5252 ( .A1(n4239), .A2(n4238), .ZN(n4408) );
  NAND4_X1 U5253 ( .A1(n4325), .A2(n4240), .A3(n3210), .A4(n3192), .ZN(n4322)
         );
  INV_X1 U5254 ( .A(n4322), .ZN(n4243) );
  NAND3_X1 U5255 ( .A1(n4243), .A2(n4242), .A3(n4241), .ZN(n4244) );
  NAND2_X1 U5256 ( .A1(n5608), .A2(n6073), .ZN(n4258) );
  NAND2_X1 U5257 ( .A1(n4250), .A2(n5426), .ZN(n4247) );
  INV_X1 U5258 ( .A(n4249), .ZN(n4246) );
  NAND3_X1 U5259 ( .A1(n4248), .A2(n4247), .A3(n4246), .ZN(n4252) );
  OAI211_X1 U5260 ( .C1(n5426), .C2(n3617), .A(n4250), .B(n4249), .ZN(n4251)
         );
  NAND2_X1 U5261 ( .A1(n4252), .A2(n4251), .ZN(n5410) );
  INV_X1 U5262 ( .A(n5410), .ZN(n4256) );
  NAND2_X1 U5263 ( .A1(n4325), .A2(n6076), .ZN(n5578) );
  INV_X1 U5264 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4253) );
  NAND2_X1 U5265 ( .A1(n4272), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4262) );
  INV_X1 U5266 ( .A(n5611), .ZN(n4260) );
  INV_X1 U5267 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6498) );
  NOR2_X1 U5268 ( .A1(n6196), .A2(n6498), .ZN(n5604) );
  NOR2_X1 U5269 ( .A1(n5410), .A2(n6198), .ZN(n4264) );
  AOI211_X1 U5270 ( .C1(n4265), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5604), .B(n4264), .ZN(n4269) );
  NAND2_X1 U5271 ( .A1(n4267), .A2(n4266), .ZN(n4268) );
  OAI21_X1 U5272 ( .B1(n5610), .B2(n6184), .A(n4270), .ZN(U2988) );
  NAND2_X1 U5273 ( .A1(n4306), .A2(n6242), .ZN(n4286) );
  NAND2_X1 U5274 ( .A1(n4273), .A2(n3617), .ZN(n4276) );
  INV_X1 U5275 ( .A(n4274), .ZN(n4275) );
  NAND2_X1 U5276 ( .A1(n4276), .A2(n4275), .ZN(n4277) );
  NOR2_X1 U5277 ( .A1(n5426), .A2(n4277), .ZN(n4278) );
  INV_X1 U5278 ( .A(REIP_REG_29__SCAN_IN), .ZN(n5418) );
  NOR2_X1 U5279 ( .A1(n6196), .A2(n5418), .ZN(n4312) );
  NOR2_X1 U5280 ( .A1(n4280), .A2(n4282), .ZN(n4281) );
  AOI211_X1 U5281 ( .C1(n6237), .C2(n5530), .A(n4312), .B(n4281), .ZN(n4284)
         );
  INV_X1 U5282 ( .A(n5743), .ZN(n5737) );
  NAND3_X1 U5283 ( .A1(n5737), .A2(n2991), .A3(n4282), .ZN(n4283) );
  NAND2_X1 U5284 ( .A1(n4286), .A2(n4285), .ZN(U2989) );
  NAND2_X1 U5285 ( .A1(n4287), .A2(n5401), .ZN(n6380) );
  INV_X1 U5286 ( .A(n6422), .ZN(n6418) );
  AOI22_X1 U5287 ( .A1(n3755), .A2(EAX_REG_31__SCAN_IN), .B1(n4288), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4289) );
  NAND3_X1 U5288 ( .A1(n6421), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6431) );
  INV_X1 U5289 ( .A(n6431), .ZN(n4291) );
  NOR2_X2 U5290 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6310) );
  INV_X2 U5291 ( .A(n6139), .ZN(n5681) );
  INV_X1 U5292 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4292) );
  INV_X1 U5293 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4294) );
  NAND2_X1 U5294 ( .A1(n6297), .A2(n4296), .ZN(n6519) );
  NAND2_X1 U5295 ( .A1(n6519), .A2(n6421), .ZN(n4297) );
  NAND2_X1 U5296 ( .A1(n6421), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4299) );
  NAND2_X1 U5297 ( .A1(n6424), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4298) );
  AND2_X1 U5298 ( .A1(n4299), .A2(n4298), .ZN(n4351) );
  INV_X1 U5299 ( .A(n4351), .ZN(n4300) );
  NAND2_X1 U5300 ( .A1(n6161), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4301)
         );
  OAI211_X1 U5301 ( .C1(n4988), .C2(n6170), .A(n4302), .B(n4301), .ZN(n4303)
         );
  AOI21_X1 U5302 ( .B1(n5388), .B2(n5681), .A(n4303), .ZN(n4304) );
  OAI21_X1 U5303 ( .B1(n6144), .B2(n4305), .A(n4304), .ZN(U2955) );
  NAND2_X1 U5304 ( .A1(n4306), .A2(n6165), .ZN(n4316) );
  INV_X1 U5305 ( .A(n5420), .ZN(n4310) );
  NOR2_X1 U5306 ( .A1(n4310), .A2(n6170), .ZN(n4311) );
  AOI211_X1 U5307 ( .C1(n6161), .C2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n4312), 
        .B(n4311), .ZN(n4313) );
  NAND2_X1 U5308 ( .A1(n4316), .A2(n4315), .ZN(U2957) );
  NAND2_X1 U5309 ( .A1(n4317), .A2(n5401), .ZN(n4321) );
  INV_X1 U5310 ( .A(n4318), .ZN(n4319) );
  OR2_X1 U5311 ( .A1(n3598), .A2(n4319), .ZN(n4320) );
  NAND2_X1 U5312 ( .A1(n4321), .A2(n4320), .ZN(n4401) );
  NOR2_X1 U5313 ( .A1(n3601), .A2(n4322), .ZN(n4323) );
  AND2_X1 U5314 ( .A1(n5581), .A2(n4325), .ZN(n4326) );
  INV_X2 U5315 ( .A(n5581), .ZN(n6084) );
  AOI22_X1 U5316 ( .A1(n6081), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6084), .ZN(n4328) );
  NAND2_X1 U5317 ( .A1(n4329), .A2(n4328), .ZN(U2860) );
  INV_X1 U5318 ( .A(n5395), .ZN(n4330) );
  NAND2_X1 U5319 ( .A1(n5404), .A2(n6422), .ZN(n5389) );
  INV_X1 U5320 ( .A(n4331), .ZN(n5403) );
  INV_X1 U5321 ( .A(n6518), .ZN(n4335) );
  NAND2_X1 U5322 ( .A1(n4332), .A2(n2958), .ZN(n5145) );
  INV_X1 U5323 ( .A(n5145), .ZN(n4333) );
  OR2_X1 U5324 ( .A1(n3335), .A2(n4333), .ZN(n5405) );
  NAND2_X1 U5325 ( .A1(n6310), .A2(n5362), .ZN(n5947) );
  INV_X1 U5326 ( .A(n5947), .ZN(n5001) );
  OAI21_X1 U5327 ( .B1(n5001), .B2(READREQUEST_REG_SCAN_IN), .A(n4335), .ZN(
        n4334) );
  OAI21_X1 U5328 ( .B1(n4335), .B2(n5405), .A(n4334), .ZN(U3474) );
  INV_X1 U5329 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4381) );
  INV_X1 U5330 ( .A(n4336), .ZN(n6410) );
  OR2_X1 U5331 ( .A1(n6389), .A2(n6410), .ZN(n4339) );
  INV_X1 U5332 ( .A(n6440), .ZN(n6408) );
  NAND2_X1 U5333 ( .A1(n6088), .A2(n4993), .ZN(n4519) );
  NAND2_X1 U5334 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4557) );
  NOR2_X4 U5335 ( .A1(n6521), .A2(n6088), .ZN(n5867) );
  AOI22_X1 U5336 ( .A1(n6521), .A2(UWORD_REG_3__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4340) );
  OAI21_X1 U5337 ( .B1(n4381), .B2(n4519), .A(n4340), .ZN(U2904) );
  AOI22_X1 U5338 ( .A1(n6521), .A2(UWORD_REG_2__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4341) );
  OAI21_X1 U5339 ( .B1(n3983), .B2(n4519), .A(n4341), .ZN(U2905) );
  INV_X1 U5340 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4383) );
  AOI22_X1 U5341 ( .A1(n6521), .A2(UWORD_REG_4__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4342) );
  OAI21_X1 U5342 ( .B1(n4383), .B2(n4519), .A(n4342), .ZN(U2903) );
  INV_X1 U5343 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4467) );
  AOI22_X1 U5344 ( .A1(n4517), .A2(UWORD_REG_7__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4343) );
  OAI21_X1 U5345 ( .B1(n4467), .B2(n4519), .A(n4343), .ZN(U2900) );
  INV_X1 U5346 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6599) );
  AOI22_X1 U5347 ( .A1(n4517), .A2(UWORD_REG_9__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4344) );
  OAI21_X1 U5348 ( .B1(n6599), .B2(n4519), .A(n4344), .ZN(U2898) );
  INV_X1 U5349 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4376) );
  AOI22_X1 U5350 ( .A1(n4517), .A2(UWORD_REG_5__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4345) );
  OAI21_X1 U5351 ( .B1(n4376), .B2(n4519), .A(n4345), .ZN(U2902) );
  INV_X1 U5352 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4472) );
  AOI22_X1 U5353 ( .A1(n4517), .A2(UWORD_REG_8__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4346) );
  OAI21_X1 U5354 ( .B1(n4472), .B2(n4519), .A(n4346), .ZN(U2899) );
  INV_X1 U5355 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4465) );
  AOI22_X1 U5356 ( .A1(n4517), .A2(UWORD_REG_6__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4347) );
  OAI21_X1 U5357 ( .B1(n4465), .B2(n4519), .A(n4347), .ZN(U2901) );
  INV_X1 U5358 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4372) );
  AOI22_X1 U5359 ( .A1(n4517), .A2(UWORD_REG_12__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4348) );
  OAI21_X1 U5360 ( .B1(n4372), .B2(n4519), .A(n4348), .ZN(U2895) );
  INV_X1 U5361 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4469) );
  AOI22_X1 U5362 ( .A1(n4517), .A2(UWORD_REG_11__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4349) );
  OAI21_X1 U5363 ( .B1(n4469), .B2(n4519), .A(n4349), .ZN(U2896) );
  XNOR2_X1 U5364 ( .A(n4350), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4368)
         );
  NAND2_X1 U5365 ( .A1(n4351), .A2(n5725), .ZN(n4357) );
  AND2_X1 U5366 ( .A1(n6240), .A2(REIP_REG_0__SCAN_IN), .ZN(n4362) );
  INV_X1 U5367 ( .A(n4352), .ZN(n4355) );
  OAI21_X1 U5368 ( .B1(n4355), .B2(n4354), .A(n4353), .ZN(n5180) );
  NOR2_X1 U5369 ( .A1(n5180), .A2(n6139), .ZN(n4356) );
  AOI211_X1 U5370 ( .C1(PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n4357), .A(n4362), 
        .B(n4356), .ZN(n4358) );
  OAI21_X1 U5371 ( .B1(n4368), .B2(n6144), .A(n4358), .ZN(U2986) );
  NOR2_X1 U5372 ( .A1(n4359), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4360)
         );
  OR2_X1 U5373 ( .A1(n4361), .A2(n4360), .ZN(n5175) );
  INV_X1 U5374 ( .A(n4362), .ZN(n4363) );
  OAI211_X1 U5375 ( .C1(n6198), .C2(n5175), .A(n4364), .B(n4363), .ZN(n4366)
         );
  AOI21_X1 U5376 ( .B1(n5346), .B2(n5270), .A(n4431), .ZN(n4365) );
  NOR2_X1 U5377 ( .A1(n4366), .A2(n4365), .ZN(n4367) );
  OAI21_X1 U5378 ( .B1(n4368), .B2(n6184), .A(n4367), .ZN(U3018) );
  INV_X1 U5379 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6116) );
  INV_X1 U5380 ( .A(n5390), .ZN(n4369) );
  NAND2_X1 U5381 ( .A1(n6126), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4370) );
  NAND2_X1 U5382 ( .A1(n6131), .A2(DATAI_0_), .ZN(n4377) );
  OAI211_X1 U5383 ( .C1(n6116), .C2(n4460), .A(n4370), .B(n4377), .ZN(U2939)
         );
  NAND2_X1 U5384 ( .A1(n6126), .A2(UWORD_REG_12__SCAN_IN), .ZN(n4371) );
  NAND2_X1 U5385 ( .A1(n6131), .A2(DATAI_12_), .ZN(n4386) );
  OAI211_X1 U5386 ( .C1(n4372), .C2(n4460), .A(n4371), .B(n4386), .ZN(U2936)
         );
  INV_X1 U5387 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U5388 ( .A1(n6126), .A2(LWORD_REG_3__SCAN_IN), .ZN(n4373) );
  NAND2_X1 U5389 ( .A1(n6131), .A2(DATAI_3_), .ZN(n4379) );
  OAI211_X1 U5390 ( .C1(n6608), .C2(n4460), .A(n4373), .B(n4379), .ZN(U2942)
         );
  INV_X1 U5391 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U5392 ( .A1(n6126), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4374) );
  NAND2_X1 U5393 ( .A1(n6131), .A2(DATAI_10_), .ZN(n4476) );
  OAI211_X1 U5394 ( .C1(n6641), .C2(n4460), .A(n4374), .B(n4476), .ZN(U2949)
         );
  NAND2_X1 U5395 ( .A1(n6126), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4375) );
  NAND2_X1 U5396 ( .A1(n6131), .A2(DATAI_5_), .ZN(n4478) );
  OAI211_X1 U5397 ( .C1(n4376), .C2(n4460), .A(n4375), .B(n4478), .ZN(U2929)
         );
  INV_X1 U5398 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4510) );
  NAND2_X1 U5399 ( .A1(n6126), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4378) );
  OAI211_X1 U5400 ( .C1(n4510), .C2(n4460), .A(n4378), .B(n4377), .ZN(U2924)
         );
  NAND2_X1 U5401 ( .A1(n6126), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4380) );
  OAI211_X1 U5402 ( .C1(n4381), .C2(n4460), .A(n4380), .B(n4379), .ZN(U2927)
         );
  NAND2_X1 U5403 ( .A1(n6126), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4382) );
  NAND2_X1 U5404 ( .A1(n6131), .A2(DATAI_4_), .ZN(n4384) );
  OAI211_X1 U5405 ( .C1(n4460), .C2(n4383), .A(n4382), .B(n4384), .ZN(U2928)
         );
  INV_X1 U5406 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U5407 ( .A1(n6126), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4385) );
  OAI211_X1 U5408 ( .C1(n4460), .C2(n6108), .A(n4385), .B(n4384), .ZN(U2943)
         );
  INV_X1 U5409 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U5410 ( .A1(n6126), .A2(LWORD_REG_12__SCAN_IN), .ZN(n4387) );
  OAI211_X1 U5411 ( .C1(n6598), .C2(n4460), .A(n4387), .B(n4386), .ZN(U2951)
         );
  INV_X1 U5412 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U5413 ( .A1(n6126), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4388) );
  NAND2_X1 U5414 ( .A1(n6131), .A2(DATAI_1_), .ZN(n4389) );
  OAI211_X1 U5415 ( .C1(n6113), .C2(n4460), .A(n4388), .B(n4389), .ZN(U2940)
         );
  INV_X1 U5416 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4512) );
  NAND2_X1 U5417 ( .A1(n6126), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4390) );
  OAI211_X1 U5418 ( .C1(n4512), .C2(n4460), .A(n4390), .B(n4389), .ZN(U2925)
         );
  NAND2_X2 U5419 ( .A1(n5581), .A2(n4392), .ZN(n5911) );
  INV_X1 U5420 ( .A(n4392), .ZN(n4393) );
  INV_X1 U5421 ( .A(DATAI_0_), .ZN(n6562) );
  OAI222_X1 U5422 ( .A1(n5180), .A2(n5911), .B1(n4705), .B2(n6562), .C1(n5581), 
        .C2(n6116), .ZN(U2891) );
  INV_X1 U5423 ( .A(n4394), .ZN(n4395) );
  OAI21_X1 U5424 ( .B1(n4397), .B2(n4396), .A(n4395), .ZN(n6072) );
  AOI22_X1 U5425 ( .A1(n5357), .A2(DATAI_2_), .B1(n6084), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n4398) );
  OAI21_X1 U5426 ( .B1(n6072), .B2(n5911), .A(n4398), .ZN(U2889) );
  OAI21_X1 U5427 ( .B1(n4400), .B2(n4993), .A(n4399), .ZN(n4402) );
  NOR2_X1 U5428 ( .A1(n4402), .A2(n4401), .ZN(n4407) );
  INV_X1 U5429 ( .A(n4403), .ZN(n4404) );
  AOI21_X1 U5430 ( .B1(n4404), .B2(n6440), .A(READY_N), .ZN(n4405) );
  OAI211_X1 U5431 ( .C1(n6389), .C2(n3518), .A(n4405), .B(n5401), .ZN(n4406)
         );
  INV_X1 U5432 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6577) );
  NOR2_X1 U5433 ( .A1(n6421), .A2(n4557), .ZN(n4555) );
  INV_X1 U5434 ( .A(n4555), .ZN(n6506) );
  OAI22_X1 U5435 ( .A1(n4544), .A2(n6418), .B1(n6577), .B2(n6506), .ZN(n4414)
         );
  AOI21_X1 U5436 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6421), .A(n4414), .ZN(
        n5369) );
  INV_X1 U5437 ( .A(n5369), .ZN(n5865) );
  INV_X1 U5438 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4416) );
  INV_X1 U5439 ( .A(n6420), .ZN(n5366) );
  INV_X1 U5440 ( .A(n3598), .ZN(n4413) );
  INV_X1 U5441 ( .A(n4603), .ZN(n4409) );
  OR2_X1 U5442 ( .A1(n4410), .A2(n4409), .ZN(n4411) );
  XNOR2_X1 U5443 ( .A(n4411), .B(n4416), .ZN(n5170) );
  INV_X1 U5444 ( .A(n5170), .ZN(n4412) );
  NAND4_X1 U5445 ( .A1(n4414), .A2(n5366), .A3(n4413), .A4(n4412), .ZN(n4415)
         );
  OAI21_X1 U5446 ( .B1(n5865), .B2(n4416), .A(n4415), .ZN(U3455) );
  INV_X1 U5447 ( .A(n3518), .ZN(n4419) );
  AND4_X1 U5448 ( .A1(n4420), .A2(n3598), .A3(n4419), .A4(n3601), .ZN(n4421)
         );
  NAND2_X1 U5449 ( .A1(n4422), .A2(n4421), .ZN(n5360) );
  NAND2_X1 U5450 ( .A1(n4418), .A2(n5360), .ZN(n4430) );
  INV_X1 U5451 ( .A(n5392), .ZN(n4423) );
  NAND2_X1 U5452 ( .A1(n4423), .A2(n5394), .ZN(n4541) );
  XNOR2_X1 U5453 ( .A(n4424), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4428)
         );
  XNOR2_X1 U5454 ( .A(n3000), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4425)
         );
  NAND2_X1 U5455 ( .A1(n6389), .A2(n4425), .ZN(n4426) );
  OAI21_X1 U5456 ( .B1(n4428), .B2(n4538), .A(n4426), .ZN(n4427) );
  AOI21_X1 U5457 ( .B1(n4541), .B2(n4428), .A(n4427), .ZN(n4429) );
  NAND2_X1 U5458 ( .A1(n4430), .A2(n4429), .ZN(n4524) );
  NOR2_X1 U5459 ( .A1(n5362), .A2(n4431), .ZN(n4446) );
  INV_X1 U5460 ( .A(n4446), .ZN(n5364) );
  AOI22_X1 U5461 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4432), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4453), .ZN(n4445) );
  NOR2_X1 U5462 ( .A1(n5364), .A2(n4445), .ZN(n4434) );
  INV_X1 U5463 ( .A(n5363), .ZN(n6415) );
  INV_X1 U5464 ( .A(n4424), .ZN(n4440) );
  NOR3_X1 U5465 ( .A1(n6415), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n4440), 
        .ZN(n4433) );
  AOI211_X1 U5466 ( .C1(n4524), .C2(n5366), .A(n4434), .B(n4433), .ZN(n4436)
         );
  AOI21_X1 U5467 ( .B1(n5363), .B2(n4440), .A(n5369), .ZN(n4435) );
  OAI22_X1 U5468 ( .A1(n4436), .A2(n5369), .B1(n4435), .B2(n3048), .ZN(U3459)
         );
  INV_X1 U5469 ( .A(n6389), .ZN(n4443) );
  INV_X1 U5470 ( .A(n5854), .ZN(n4806) );
  NAND2_X1 U5471 ( .A1(n4806), .A2(n5360), .ZN(n4442) );
  INV_X1 U5472 ( .A(n4438), .ZN(n5359) );
  INV_X1 U5473 ( .A(n4439), .ZN(n4552) );
  NAND3_X1 U5474 ( .A1(n5359), .A2(n4552), .A3(n4440), .ZN(n4441) );
  OAI211_X1 U5475 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n4443), .A(n4442), .B(n4441), .ZN(n6386) );
  AOI222_X1 U5476 ( .A1(n6386), .A2(n5366), .B1(n4446), .B2(n4445), .C1(n4444), 
        .C2(n5363), .ZN(n4449) );
  AOI22_X1 U5477 ( .A1(n5363), .A2(n4447), .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n5369), .ZN(n4448) );
  OAI21_X1 U5478 ( .B1(n4449), .B2(n5369), .A(n4448), .ZN(U3460) );
  XOR2_X1 U5479 ( .A(n4451), .B(n4450), .Z(n4485) );
  INV_X1 U5480 ( .A(n4485), .ZN(n4459) );
  XNOR2_X1 U5481 ( .A(n4452), .B(n4998), .ZN(n5147) );
  INV_X1 U5482 ( .A(n5147), .ZN(n4455) );
  INV_X1 U5483 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6509) );
  NOR2_X1 U5484 ( .A1(n6196), .A2(n6509), .ZN(n4487) );
  NOR2_X1 U5485 ( .A1(n4453), .A2(n4685), .ZN(n4454) );
  AOI211_X1 U5486 ( .C1(n6237), .C2(n4455), .A(n4487), .B(n4454), .ZN(n4458)
         );
  OR3_X1 U5487 ( .A1(n5831), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4456), 
        .ZN(n4457) );
  OAI211_X1 U5488 ( .C1(n4459), .C2(n6184), .A(n4458), .B(n4457), .ZN(U3017)
         );
  INV_X1 U5489 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4514) );
  AOI22_X1 U5490 ( .A1(n6130), .A2(UWORD_REG_13__SCAN_IN), .B1(n6131), .B2(
        DATAI_13_), .ZN(n4461) );
  OAI21_X1 U5491 ( .B1(n4514), .B2(n4480), .A(n4461), .ZN(U2937) );
  INV_X1 U5492 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6090) );
  AOI22_X1 U5493 ( .A1(n6130), .A2(LWORD_REG_15__SCAN_IN), .B1(n6131), .B2(
        DATAI_15_), .ZN(n4462) );
  OAI21_X1 U5494 ( .B1(n6090), .B2(n4480), .A(n4462), .ZN(U2954) );
  AOI22_X1 U5495 ( .A1(n6130), .A2(UWORD_REG_9__SCAN_IN), .B1(n6131), .B2(
        DATAI_9_), .ZN(n4463) );
  OAI21_X1 U5496 ( .B1(n6599), .B2(n4480), .A(n4463), .ZN(U2933) );
  AOI22_X1 U5497 ( .A1(n6126), .A2(UWORD_REG_6__SCAN_IN), .B1(n6131), .B2(
        DATAI_6_), .ZN(n4464) );
  OAI21_X1 U5498 ( .B1(n4465), .B2(n4480), .A(n4464), .ZN(U2930) );
  AOI22_X1 U5499 ( .A1(n6126), .A2(UWORD_REG_7__SCAN_IN), .B1(n6131), .B2(
        DATAI_7_), .ZN(n4466) );
  OAI21_X1 U5500 ( .B1(n4467), .B2(n4480), .A(n4466), .ZN(U2931) );
  AOI22_X1 U5501 ( .A1(n6130), .A2(UWORD_REG_11__SCAN_IN), .B1(n6131), .B2(
        DATAI_11_), .ZN(n4468) );
  OAI21_X1 U5502 ( .B1(n4469), .B2(n4480), .A(n4468), .ZN(U2935) );
  INV_X1 U5503 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4520) );
  AOI22_X1 U5504 ( .A1(n6130), .A2(UWORD_REG_14__SCAN_IN), .B1(n6131), .B2(
        DATAI_14_), .ZN(n4470) );
  OAI21_X1 U5505 ( .B1(n4520), .B2(n4480), .A(n4470), .ZN(U2938) );
  AOI22_X1 U5506 ( .A1(n6126), .A2(UWORD_REG_8__SCAN_IN), .B1(n6131), .B2(
        DATAI_8_), .ZN(n4471) );
  OAI21_X1 U5507 ( .B1(n4472), .B2(n4480), .A(n4471), .ZN(U2932) );
  INV_X1 U5508 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U5509 ( .A1(n6126), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4473) );
  NAND2_X1 U5510 ( .A1(n6131), .A2(DATAI_2_), .ZN(n4474) );
  OAI211_X1 U5511 ( .C1(n6111), .C2(n4480), .A(n4473), .B(n4474), .ZN(U2941)
         );
  NAND2_X1 U5512 ( .A1(n6126), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4475) );
  OAI211_X1 U5513 ( .C1(n3983), .C2(n4480), .A(n4475), .B(n4474), .ZN(U2926)
         );
  INV_X1 U5514 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4516) );
  NAND2_X1 U5515 ( .A1(n6126), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4477) );
  OAI211_X1 U5516 ( .C1(n4516), .C2(n4480), .A(n4477), .B(n4476), .ZN(U2934)
         );
  INV_X1 U5517 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U5518 ( .A1(n6126), .A2(LWORD_REG_5__SCAN_IN), .ZN(n4479) );
  OAI211_X1 U5519 ( .C1(n6106), .C2(n4480), .A(n4479), .B(n4478), .ZN(U2944)
         );
  NOR2_X1 U5520 ( .A1(n4482), .A2(n4481), .ZN(n4483) );
  NAND2_X1 U5521 ( .A1(n4485), .A2(n6165), .ZN(n4489) );
  NOR2_X1 U5522 ( .A1(n5725), .A2(n6623), .ZN(n4486) );
  AOI211_X1 U5523 ( .C1(n5728), .C2(n6623), .A(n4487), .B(n4486), .ZN(n4488)
         );
  OAI211_X1 U5524 ( .C1(n5152), .C2(n6139), .A(n4489), .B(n4488), .ZN(U2985)
         );
  OAI21_X1 U5525 ( .B1(n4394), .B2(n4491), .A(n4490), .ZN(n6069) );
  AOI22_X1 U5526 ( .A1(n5357), .A2(DATAI_3_), .B1(n6084), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n4492) );
  OAI21_X1 U5527 ( .B1(n6069), .B2(n5911), .A(n4492), .ZN(U2888) );
  OAI21_X1 U5528 ( .B1(n4493), .B2(n4496), .A(n4495), .ZN(n5163) );
  XNOR2_X1 U5529 ( .A(n4497), .B(n4504), .ZN(n5155) );
  OAI22_X1 U5530 ( .A1(n5578), .A2(n5155), .B1(n6076), .B2(n4498), .ZN(n4499)
         );
  INV_X1 U5531 ( .A(n4499), .ZN(n4500) );
  OAI21_X1 U5532 ( .B1(n5163), .B2(n5579), .A(n4500), .ZN(U2854) );
  AND2_X1 U5533 ( .A1(n4490), .A2(n4501), .ZN(n4502) );
  OR2_X1 U5534 ( .A1(n4502), .A2(n4493), .ZN(n5174) );
  OR2_X1 U5535 ( .A1(n4503), .A2(n6043), .ZN(n4505) );
  AND2_X1 U5536 ( .A1(n4505), .A2(n4504), .ZN(n6223) );
  INV_X1 U5537 ( .A(n6223), .ZN(n4506) );
  OAI222_X1 U5538 ( .A1(n5174), .A2(n5579), .B1(n6076), .B2(n3620), .C1(n4506), 
        .C2(n5578), .ZN(U2855) );
  INV_X1 U5539 ( .A(DATAI_4_), .ZN(n4507) );
  OAI222_X1 U5540 ( .A1(n5174), .A2(n5911), .B1(n4705), .B2(n4507), .C1(n6108), 
        .C2(n5581), .ZN(U2887) );
  INV_X1 U5541 ( .A(DATAI_1_), .ZN(n4508) );
  OAI222_X1 U5542 ( .A1(n5152), .A2(n5911), .B1(n4705), .B2(n4508), .C1(n5581), 
        .C2(n6113), .ZN(U2890) );
  AOI22_X1 U5543 ( .A1(n6521), .A2(UWORD_REG_0__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4509) );
  OAI21_X1 U5544 ( .B1(n4510), .B2(n4519), .A(n4509), .ZN(U2907) );
  AOI22_X1 U5545 ( .A1(n6521), .A2(UWORD_REG_1__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4511) );
  OAI21_X1 U5546 ( .B1(n4512), .B2(n4519), .A(n4511), .ZN(U2906) );
  AOI22_X1 U5547 ( .A1(n4517), .A2(UWORD_REG_13__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4513) );
  OAI21_X1 U5548 ( .B1(n4514), .B2(n4519), .A(n4513), .ZN(U2894) );
  AOI22_X1 U5549 ( .A1(n4517), .A2(UWORD_REG_10__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4515) );
  OAI21_X1 U5550 ( .B1(n4516), .B2(n4519), .A(n4515), .ZN(U2897) );
  AOI22_X1 U5551 ( .A1(n4517), .A2(UWORD_REG_14__SCAN_IN), .B1(
        DATAO_REG_30__SCAN_IN), .B2(n5867), .ZN(n4518) );
  OAI21_X1 U5552 ( .B1(n4520), .B2(n4519), .A(n4518), .ZN(U2893) );
  INV_X1 U5553 ( .A(DATAI_5_), .ZN(n6565) );
  OAI222_X1 U5554 ( .A1(n5163), .A2(n5911), .B1(n4705), .B2(n6565), .C1(n5581), 
        .C2(n6106), .ZN(U2886) );
  NOR2_X1 U5555 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6524) );
  OR3_X1 U5556 ( .A1(n5170), .A2(STATE2_REG_1__SCAN_IN), .A3(n3598), .ZN(n4523) );
  MUX2_X1 U5557 ( .A(n4544), .B(n6577), .S(STATE2_REG_1__SCAN_IN), .Z(n4521)
         );
  NAND2_X1 U5558 ( .A1(n4521), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4522) );
  NAND2_X1 U5559 ( .A1(n4523), .A2(n4522), .ZN(n4553) );
  INV_X1 U5560 ( .A(n4544), .ZN(n6387) );
  NAND2_X1 U5561 ( .A1(n4524), .A2(n6387), .ZN(n4526) );
  NAND2_X1 U5562 ( .A1(n4544), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4525) );
  NAND2_X1 U5563 ( .A1(n2961), .A2(n5360), .ZN(n4543) );
  MUX2_X1 U5564 ( .A(n4528), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4424), 
        .Z(n4529) );
  NOR2_X1 U5565 ( .A1(n4529), .A2(n4548), .ZN(n4540) );
  INV_X1 U5566 ( .A(n4530), .ZN(n4531) );
  OAI21_X1 U5567 ( .B1(n4424), .B2(n3526), .A(n4531), .ZN(n4533) );
  NOR2_X1 U5568 ( .A1(n4533), .A2(n4532), .ZN(n5863) );
  AND2_X1 U5569 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4535) );
  INV_X1 U5570 ( .A(n4535), .ZN(n4534) );
  MUX2_X1 U5571 ( .A(n4535), .B(n4534), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4536) );
  NAND2_X1 U5572 ( .A1(n6389), .A2(n4536), .ZN(n4537) );
  OAI21_X1 U5573 ( .B1(n5863), .B2(n4538), .A(n4537), .ZN(n4539) );
  AOI21_X1 U5574 ( .B1(n4541), .B2(n4540), .A(n4539), .ZN(n4542) );
  NAND2_X1 U5575 ( .A1(n4543), .A2(n4542), .ZN(n5862) );
  OR2_X1 U5576 ( .A1(n5862), .A2(n4544), .ZN(n4546) );
  NAND2_X1 U5577 ( .A1(n4544), .A2(n3526), .ZN(n4545) );
  NAND2_X1 U5578 ( .A1(n4546), .A2(n4545), .ZN(n6401) );
  OR3_X1 U5579 ( .A1(n6397), .A2(n6401), .A3(STATE2_REG_1__SCAN_IN), .ZN(n4551) );
  NOR2_X1 U5580 ( .A1(FLUSH_REG_SCAN_IN), .A2(n5362), .ZN(n4547) );
  AND2_X1 U5581 ( .A1(n4548), .A2(n4547), .ZN(n4549) );
  NOR2_X1 U5582 ( .A1(n4553), .A2(n4549), .ZN(n4550) );
  NAND2_X1 U5583 ( .A1(n4551), .A2(n4550), .ZN(n6385) );
  OAI21_X1 U5584 ( .B1(n4553), .B2(n4552), .A(n6385), .ZN(n4554) );
  INV_X1 U5585 ( .A(n4554), .ZN(n4558) );
  OAI21_X1 U5586 ( .B1(n4558), .B2(FLUSH_REG_SCAN_IN), .A(n4555), .ZN(n4556)
         );
  NAND2_X1 U5587 ( .A1(n4911), .A2(n4556), .ZN(n6249) );
  NOR2_X1 U5588 ( .A1(n4558), .A2(n4557), .ZN(n6414) );
  INV_X1 U5589 ( .A(n5361), .ZN(n6299) );
  AND2_X1 U5590 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6508), .ZN(n5858) );
  OAI22_X1 U5591 ( .A1(n5098), .A2(n6297), .B1(n6299), .B2(n5858), .ZN(n4560)
         );
  OAI21_X1 U5592 ( .B1(n6414), .B2(n4560), .A(n6249), .ZN(n4561) );
  OAI21_X1 U5593 ( .B1(n6249), .B2(n6388), .A(n4561), .ZN(U3465) );
  NAND2_X1 U5594 ( .A1(n2963), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5852) );
  NOR3_X1 U5595 ( .A1(n5023), .A2(n4706), .A3(n5852), .ZN(n6298) );
  INV_X1 U5596 ( .A(n4765), .ZN(n4804) );
  NOR2_X1 U5597 ( .A1(n6298), .A2(n4804), .ZN(n4565) );
  INV_X1 U5598 ( .A(n4706), .ZN(n5096) );
  NOR2_X1 U5599 ( .A1(n2963), .A2(n5096), .ZN(n4564) );
  NAND2_X1 U5600 ( .A1(n4825), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4818) );
  AOI21_X1 U5601 ( .B1(n4565), .B2(n4818), .A(n6297), .ZN(n4647) );
  AND2_X1 U5602 ( .A1(n6310), .A2(n6424), .ZN(n5028) );
  INV_X1 U5603 ( .A(n5028), .ZN(n5225) );
  OAI22_X1 U5604 ( .A1(n5025), .A2(n5225), .B1(n6052), .B2(n5858), .ZN(n4566)
         );
  OAI21_X1 U5605 ( .B1(n4647), .B2(n4566), .A(n6249), .ZN(n4567) );
  OAI21_X1 U5606 ( .B1(n6249), .B2(n6263), .A(n4567), .ZN(U3462) );
  OAI222_X1 U5607 ( .A1(n5147), .A2(n5578), .B1(n6076), .B2(n3604), .C1(n5152), 
        .C2(n5579), .ZN(U2858) );
  CLKBUF_X1 U5608 ( .A(n4569), .Z(n4570) );
  OAI21_X1 U5609 ( .B1(n4571), .B2(n4568), .A(n4570), .ZN(n6221) );
  INV_X1 U5610 ( .A(n5174), .ZN(n4574) );
  AOI22_X1 U5611 ( .A1(n6161), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6240), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n4572) );
  OAI21_X1 U5612 ( .B1(n5164), .B2(n6170), .A(n4572), .ZN(n4573) );
  AOI21_X1 U5613 ( .B1(n4574), .B2(n5681), .A(n4573), .ZN(n4575) );
  OAI21_X1 U5614 ( .B1(n6144), .B2(n6221), .A(n4575), .ZN(U2982) );
  OAI222_X1 U5615 ( .A1(n5175), .A2(n5578), .B1(n6626), .B2(n6076), .C1(n5180), 
        .C2(n5579), .ZN(U2859) );
  NAND2_X1 U5616 ( .A1(n4495), .A2(n4576), .ZN(n4577) );
  AND2_X1 U5617 ( .A1(n4588), .A2(n4577), .ZN(n6149) );
  INV_X1 U5618 ( .A(n6149), .ZN(n4580) );
  INV_X1 U5619 ( .A(DATAI_6_), .ZN(n4578) );
  OAI222_X1 U5620 ( .A1(n4580), .A2(n5911), .B1(n5581), .B2(n4579), .C1(n4705), 
        .C2(n4578), .ZN(U2885) );
  OR2_X1 U5621 ( .A1(n4582), .A2(n4581), .ZN(n4583) );
  AND2_X1 U5622 ( .A1(n4583), .A2(n4589), .ZN(n6216) );
  INV_X1 U5623 ( .A(n6216), .ZN(n4584) );
  OAI22_X1 U5624 ( .A1(n5578), .A2(n4584), .B1(n6076), .B2(n6537), .ZN(n4585)
         );
  AOI21_X1 U5625 ( .B1(n6149), .B2(n6073), .A(n4585), .ZN(n4586) );
  INV_X1 U5626 ( .A(n4586), .ZN(U2853) );
  XOR2_X1 U5627 ( .A(n4587), .B(n4588), .Z(n4702) );
  NAND2_X1 U5628 ( .A1(n4590), .A2(n4589), .ZN(n4592) );
  INV_X1 U5629 ( .A(n4802), .ZN(n4591) );
  NAND2_X1 U5630 ( .A1(n4592), .A2(n4591), .ZN(n5000) );
  OAI22_X1 U5631 ( .A1(n5578), .A2(n5000), .B1(n6076), .B2(n5007), .ZN(n4593)
         );
  AOI21_X1 U5632 ( .B1(n4702), .B2(n6073), .A(n4593), .ZN(n4594) );
  INV_X1 U5633 ( .A(n4594), .ZN(U2852) );
  OAI21_X1 U5634 ( .B1(n4597), .B2(n4595), .A(n4596), .ZN(n4695) );
  NAND2_X1 U5635 ( .A1(n6240), .A2(REIP_REG_5__SCAN_IN), .ZN(n4690) );
  OAI21_X1 U5636 ( .B1(n5725), .B2(n4598), .A(n4690), .ZN(n4600) );
  NOR2_X1 U5637 ( .A1(n5163), .A2(n6139), .ZN(n4599) );
  AOI211_X1 U5638 ( .C1(n5728), .C2(n5161), .A(n4600), .B(n4599), .ZN(n4601)
         );
  OAI21_X1 U5639 ( .B1(n6144), .B2(n4695), .A(n4601), .ZN(U2981) );
  NOR2_X1 U5640 ( .A1(n2963), .A2(n4706), .ZN(n4602) );
  AOI21_X1 U5641 ( .B1(n4608), .B2(STATEBS16_REG_SCAN_IN), .A(n6297), .ZN(
        n4875) );
  NAND2_X1 U5642 ( .A1(n4418), .A2(n5854), .ZN(n4915) );
  OR2_X1 U5643 ( .A1(n4915), .A2(n4603), .ZN(n4874) );
  NAND2_X1 U5644 ( .A1(n6394), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4822) );
  INV_X1 U5645 ( .A(n4822), .ZN(n4815) );
  NAND2_X1 U5646 ( .A1(n4815), .A2(n6263), .ZN(n4870) );
  NOR2_X1 U5647 ( .A1(n6388), .A2(n4870), .ZN(n4637) );
  INV_X1 U5648 ( .A(n4637), .ZN(n4604) );
  OAI21_X1 U5649 ( .B1(n4874), .B2(n6299), .A(n4604), .ZN(n4611) );
  INV_X1 U5650 ( .A(n4870), .ZN(n4605) );
  AOI22_X1 U5651 ( .A1(n4875), .A2(n4611), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4605), .ZN(n4641) );
  NAND2_X1 U5652 ( .A1(DATAI_5_), .A2(n4872), .ZN(n6339) );
  NAND2_X1 U5653 ( .A1(n3072), .A2(n4607), .ZN(n4844) );
  NAND2_X1 U5654 ( .A1(n5681), .A2(DATAI_21_), .ZN(n6283) );
  NAND2_X1 U5655 ( .A1(n5681), .A2(DATAI_29_), .ZN(n6379) );
  NAND2_X1 U5656 ( .A1(n4608), .A2(n5098), .ZN(n4900) );
  OAI22_X1 U5657 ( .A1(n4635), .A2(n6283), .B1(n6379), .B2(n4900), .ZN(n4609)
         );
  AOI21_X1 U5658 ( .B1(n6372), .B2(n4637), .A(n4609), .ZN(n4614) );
  INV_X1 U5659 ( .A(n4875), .ZN(n4612) );
  AOI21_X1 U5660 ( .B1(n4870), .B2(n6297), .A(n5065), .ZN(n4610) );
  NAND2_X1 U5661 ( .A1(n4638), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4613) );
  OAI211_X1 U5662 ( .C1(n4641), .C2(n6339), .A(n4614), .B(n4613), .ZN(U3065)
         );
  NAND2_X1 U5663 ( .A1(DATAI_4_), .A2(n4872), .ZN(n6335) );
  NAND2_X1 U5664 ( .A1(n3072), .A2(n3199), .ZN(n4841) );
  NAND2_X1 U5665 ( .A1(n5681), .A2(DATAI_20_), .ZN(n6280) );
  AND2_X1 U5666 ( .A1(n5681), .A2(DATAI_28_), .ZN(n6330) );
  INV_X1 U5667 ( .A(n6330), .ZN(n5130) );
  OAI22_X1 U5668 ( .A1(n4635), .A2(n6280), .B1(n5130), .B2(n4900), .ZN(n4615)
         );
  AOI21_X1 U5669 ( .B1(n6331), .B2(n4637), .A(n4615), .ZN(n4617) );
  NAND2_X1 U5670 ( .A1(n4638), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4616) );
  OAI211_X1 U5671 ( .C1(n4641), .C2(n6335), .A(n4617), .B(n4616), .ZN(U3064)
         );
  NAND2_X1 U5672 ( .A1(DATAI_3_), .A2(n4872), .ZN(n6329) );
  NAND2_X1 U5673 ( .A1(n3072), .A2(n3219), .ZN(n4828) );
  NAND2_X1 U5674 ( .A1(n5681), .A2(DATAI_19_), .ZN(n6276) );
  AND2_X1 U5675 ( .A1(n5681), .A2(DATAI_27_), .ZN(n6326) );
  INV_X1 U5676 ( .A(n6326), .ZN(n6368) );
  OAI22_X1 U5677 ( .A1(n4635), .A2(n6276), .B1(n6368), .B2(n4900), .ZN(n4618)
         );
  AOI21_X1 U5678 ( .B1(n6364), .B2(n4637), .A(n4618), .ZN(n4620) );
  NAND2_X1 U5679 ( .A1(n4638), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4619) );
  OAI211_X1 U5680 ( .C1(n4641), .C2(n6329), .A(n4620), .B(n4619), .ZN(U3063)
         );
  NAND2_X1 U5681 ( .A1(DATAI_2_), .A2(n4872), .ZN(n6325) );
  NAND2_X1 U5682 ( .A1(n3072), .A2(n4621), .ZN(n4857) );
  NAND2_X1 U5683 ( .A1(n5681), .A2(DATAI_18_), .ZN(n6273) );
  AND2_X1 U5684 ( .A1(n5681), .A2(DATAI_26_), .ZN(n6320) );
  INV_X1 U5685 ( .A(n6320), .ZN(n5126) );
  OAI22_X1 U5686 ( .A1(n4635), .A2(n6273), .B1(n5126), .B2(n4900), .ZN(n4622)
         );
  AOI21_X1 U5687 ( .B1(n6321), .B2(n4637), .A(n4622), .ZN(n4624) );
  NAND2_X1 U5688 ( .A1(n4638), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4623) );
  OAI211_X1 U5689 ( .C1(n4641), .C2(n6325), .A(n4624), .B(n4623), .ZN(U3062)
         );
  NAND2_X1 U5690 ( .A1(DATAI_6_), .A2(n4872), .ZN(n6345) );
  NAND2_X1 U5691 ( .A1(n3072), .A2(n3192), .ZN(n4835) );
  NAND2_X1 U5692 ( .A1(n5681), .A2(DATAI_22_), .ZN(n6287) );
  AND2_X1 U5693 ( .A1(n5681), .A2(DATAI_30_), .ZN(n6340) );
  INV_X1 U5694 ( .A(n6340), .ZN(n5108) );
  OAI22_X1 U5695 ( .A1(n4635), .A2(n6287), .B1(n5108), .B2(n4900), .ZN(n4625)
         );
  AOI21_X1 U5696 ( .B1(n6341), .B2(n4637), .A(n4625), .ZN(n4627) );
  NAND2_X1 U5697 ( .A1(n4638), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4626) );
  OAI211_X1 U5698 ( .C1(n4641), .C2(n6345), .A(n4627), .B(n4626), .ZN(U3066)
         );
  NAND2_X1 U5699 ( .A1(DATAI_7_), .A2(n4872), .ZN(n6355) );
  NAND2_X1 U5700 ( .A1(n5681), .A2(DATAI_23_), .ZN(n6296) );
  AND2_X1 U5701 ( .A1(n5681), .A2(DATAI_31_), .ZN(n6347) );
  INV_X1 U5702 ( .A(n6347), .ZN(n5122) );
  OAI22_X1 U5703 ( .A1(n4635), .A2(n6296), .B1(n5122), .B2(n4900), .ZN(n4628)
         );
  AOI21_X1 U5704 ( .B1(n6349), .B2(n4637), .A(n4628), .ZN(n4630) );
  NAND2_X1 U5705 ( .A1(n4638), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4629) );
  OAI211_X1 U5706 ( .C1(n4641), .C2(n6355), .A(n4630), .B(n4629), .ZN(U3067)
         );
  NAND2_X1 U5707 ( .A1(DATAI_1_), .A2(n4872), .ZN(n6319) );
  NAND2_X1 U5708 ( .A1(n3072), .A2(n2958), .ZN(n4850) );
  NAND2_X1 U5709 ( .A1(n5681), .A2(DATAI_17_), .ZN(n6269) );
  NAND2_X1 U5710 ( .A1(n5681), .A2(DATAI_25_), .ZN(n6362) );
  OAI22_X1 U5711 ( .A1(n4635), .A2(n6269), .B1(n6362), .B2(n4900), .ZN(n4632)
         );
  AOI21_X1 U5712 ( .B1(n6358), .B2(n4637), .A(n4632), .ZN(n4634) );
  NAND2_X1 U5713 ( .A1(n4638), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4633) );
  OAI211_X1 U5714 ( .C1(n4641), .C2(n6319), .A(n4634), .B(n4633), .ZN(U3061)
         );
  NAND2_X1 U5715 ( .A1(DATAI_0_), .A2(n4872), .ZN(n6315) );
  NAND2_X1 U5716 ( .A1(n3072), .A2(n4993), .ZN(n4847) );
  NAND2_X1 U5717 ( .A1(n5681), .A2(DATAI_16_), .ZN(n6266) );
  AND2_X1 U5718 ( .A1(n5681), .A2(DATAI_24_), .ZN(n6312) );
  INV_X1 U5719 ( .A(n6312), .ZN(n5118) );
  OAI22_X1 U5720 ( .A1(n4635), .A2(n6266), .B1(n5118), .B2(n4900), .ZN(n4636)
         );
  AOI21_X1 U5721 ( .B1(n6304), .B2(n4637), .A(n4636), .ZN(n4640) );
  NAND2_X1 U5722 ( .A1(n4638), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4639) );
  OAI211_X1 U5723 ( .C1(n4641), .C2(n6315), .A(n4640), .B(n4639), .ZN(U3060)
         );
  OAI21_X1 U5724 ( .B1(n4644), .B2(n4643), .A(n4642), .ZN(n5197) );
  AOI22_X1 U5725 ( .A1(n5357), .A2(DATAI_8_), .B1(n6084), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4645) );
  OAI21_X1 U5726 ( .B1(n5197), .B2(n5911), .A(n4645), .ZN(U2883) );
  INV_X1 U5727 ( .A(n5852), .ZN(n5856) );
  AOI21_X1 U5728 ( .B1(n5023), .B2(n5856), .A(n6297), .ZN(n4646) );
  NOR2_X1 U5729 ( .A1(n4647), .A2(n4646), .ZN(n4654) );
  INV_X1 U5730 ( .A(n4654), .ZN(n4651) );
  NOR2_X1 U5731 ( .A1(n4418), .A2(n5854), .ZN(n4741) );
  NAND2_X1 U5732 ( .A1(n6052), .A2(n4741), .ZN(n5231) );
  OR2_X1 U5733 ( .A1(n5231), .A2(n6299), .ZN(n4649) );
  INV_X1 U5734 ( .A(n4742), .ZN(n4648) );
  NAND2_X1 U5735 ( .A1(n4648), .A2(n6263), .ZN(n4678) );
  NAND2_X1 U5736 ( .A1(n4649), .A2(n4678), .ZN(n4653) );
  NAND3_X1 U5737 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6263), .A3(n5030), .ZN(n5224) );
  INV_X1 U5738 ( .A(n5224), .ZN(n4650) );
  AOI21_X1 U5739 ( .B1(n6297), .B2(n5224), .A(n5065), .ZN(n4652) );
  NAND2_X1 U5740 ( .A1(n4677), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4658) );
  NAND3_X1 U5741 ( .A1(n5025), .A2(n5023), .A3(n2963), .ZN(n4655) );
  NOR2_X2 U5742 ( .A1(n4655), .A2(n6250), .ZN(n5255) );
  OAI22_X1 U5743 ( .A1(n4857), .A2(n4678), .B1(n6273), .B2(n4906), .ZN(n4656)
         );
  AOI21_X1 U5744 ( .B1(n6320), .B2(n5255), .A(n4656), .ZN(n4657) );
  OAI211_X1 U5745 ( .C1(n4682), .C2(n6325), .A(n4658), .B(n4657), .ZN(U3046)
         );
  NAND2_X1 U5746 ( .A1(n4677), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4661) );
  OAI22_X1 U5747 ( .A1(n4847), .A2(n4678), .B1(n6266), .B2(n4906), .ZN(n4659)
         );
  AOI21_X1 U5748 ( .B1(n6312), .B2(n5255), .A(n4659), .ZN(n4660) );
  OAI211_X1 U5749 ( .C1(n4682), .C2(n6315), .A(n4661), .B(n4660), .ZN(U3044)
         );
  NAND2_X1 U5750 ( .A1(n4677), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4664) );
  OAI22_X1 U5751 ( .A1(n4841), .A2(n4678), .B1(n6280), .B2(n4906), .ZN(n4662)
         );
  AOI21_X1 U5752 ( .B1(n6330), .B2(n5255), .A(n4662), .ZN(n4663) );
  OAI211_X1 U5753 ( .C1(n4682), .C2(n6335), .A(n4664), .B(n4663), .ZN(U3048)
         );
  NAND2_X1 U5754 ( .A1(n4677), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4667) );
  OAI22_X1 U5755 ( .A1(n4828), .A2(n4678), .B1(n6276), .B2(n4906), .ZN(n4665)
         );
  AOI21_X1 U5756 ( .B1(n6326), .B2(n5255), .A(n4665), .ZN(n4666) );
  OAI211_X1 U5757 ( .C1(n4682), .C2(n6329), .A(n4667), .B(n4666), .ZN(U3047)
         );
  NAND2_X1 U5758 ( .A1(n4677), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4670) );
  OAI22_X1 U5759 ( .A1(n4838), .A2(n4678), .B1(n6296), .B2(n4906), .ZN(n4668)
         );
  AOI21_X1 U5760 ( .B1(n6347), .B2(n5255), .A(n4668), .ZN(n4669) );
  OAI211_X1 U5761 ( .C1(n4682), .C2(n6355), .A(n4670), .B(n4669), .ZN(U3051)
         );
  NAND2_X1 U5762 ( .A1(n4677), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4673) );
  OAI22_X1 U5763 ( .A1(n4835), .A2(n4678), .B1(n6287), .B2(n4906), .ZN(n4671)
         );
  AOI21_X1 U5764 ( .B1(n6340), .B2(n5255), .A(n4671), .ZN(n4672) );
  OAI211_X1 U5765 ( .C1(n4682), .C2(n6345), .A(n4673), .B(n4672), .ZN(U3050)
         );
  NAND2_X1 U5766 ( .A1(n4677), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4676) );
  INV_X1 U5767 ( .A(n6379), .ZN(n6336) );
  OAI22_X1 U5768 ( .A1(n4844), .A2(n4678), .B1(n6283), .B2(n4906), .ZN(n4674)
         );
  AOI21_X1 U5769 ( .B1(n6336), .B2(n5255), .A(n4674), .ZN(n4675) );
  OAI211_X1 U5770 ( .C1(n4682), .C2(n6339), .A(n4676), .B(n4675), .ZN(U3049)
         );
  NAND2_X1 U5771 ( .A1(n4677), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4681) );
  INV_X1 U5772 ( .A(n6362), .ZN(n6316) );
  OAI22_X1 U5773 ( .A1(n4850), .A2(n4678), .B1(n6269), .B2(n4906), .ZN(n4679)
         );
  AOI21_X1 U5774 ( .B1(n6316), .B2(n5255), .A(n4679), .ZN(n4680) );
  OAI211_X1 U5775 ( .C1(n4682), .C2(n6319), .A(n4681), .B(n4680), .ZN(U3045)
         );
  NOR2_X1 U5776 ( .A1(n4684), .A2(n4683), .ZN(n6239) );
  OAI22_X1 U5777 ( .A1(n6236), .A2(n4685), .B1(n5339), .B2(n5332), .ZN(n6243)
         );
  NOR2_X1 U5778 ( .A1(n6239), .A2(n6243), .ZN(n6234) );
  OAI21_X1 U5779 ( .B1(n6214), .B2(n5831), .A(n6234), .ZN(n4686) );
  INV_X1 U5780 ( .A(n4686), .ZN(n6218) );
  AOI221_X1 U5781 ( .B1(n4688), .B2(n4687), .C1(n6224), .C2(n4687), .A(n6218), 
        .ZN(n4693) );
  NOR3_X1 U5782 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4689), .A3(n6224), 
        .ZN(n4692) );
  OAI21_X1 U5783 ( .B1(n6198), .B2(n5155), .A(n4690), .ZN(n4691) );
  NOR3_X1 U5784 ( .A1(n4693), .A2(n4692), .A3(n4691), .ZN(n4694) );
  OAI21_X1 U5785 ( .B1(n6184), .B2(n4695), .A(n4694), .ZN(U3013) );
  OAI21_X1 U5786 ( .B1(n4698), .B2(n4697), .A(n4696), .ZN(n6208) );
  NAND2_X1 U5787 ( .A1(n6240), .A2(REIP_REG_7__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U5788 ( .A1(n6161), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4699)
         );
  OAI211_X1 U5789 ( .C1(n6170), .C2(n4989), .A(n6205), .B(n4699), .ZN(n4700)
         );
  AOI21_X1 U5790 ( .B1(n4702), .B2(n5681), .A(n4700), .ZN(n4701) );
  OAI21_X1 U5791 ( .B1(n6208), .B2(n6144), .A(n4701), .ZN(U2979) );
  INV_X1 U5792 ( .A(DATAI_7_), .ZN(n4704) );
  INV_X1 U5793 ( .A(n4702), .ZN(n5011) );
  OAI222_X1 U5794 ( .A1(n4705), .A2(n4704), .B1(n5911), .B2(n5011), .C1(n4703), 
        .C2(n5581), .ZN(U2884) );
  INV_X1 U5795 ( .A(n4950), .ZN(n4953) );
  NOR2_X1 U5796 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4953), .ZN(n4736)
         );
  OAI21_X1 U5797 ( .B1(n6253), .B2(n5069), .A(n4872), .ZN(n6258) );
  NOR2_X1 U5798 ( .A1(n4712), .A2(n5069), .ZN(n6259) );
  NOR3_X1 U5799 ( .A1(n6258), .A2(n6263), .A3(n6259), .ZN(n4710) );
  NAND2_X1 U5800 ( .A1(n4418), .A2(n4806), .ZN(n6252) );
  AND2_X1 U5801 ( .A1(n2963), .A2(n4706), .ZN(n4707) );
  OAI21_X1 U5802 ( .B1(n4853), .B2(n4977), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4708) );
  NAND3_X1 U5803 ( .A1(n6252), .A2(n6310), .A3(n4708), .ZN(n4709) );
  OAI211_X1 U5804 ( .C1(n4736), .C2(n6508), .A(n4710), .B(n4709), .ZN(n4711)
         );
  INV_X1 U5805 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4716) );
  INV_X1 U5806 ( .A(n6253), .ZN(n4713) );
  AND2_X1 U5807 ( .A1(n4712), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6254) );
  INV_X1 U5808 ( .A(n6254), .ZN(n5103) );
  OAI33_X1 U5809 ( .A1(n4713), .A2(n6263), .A3(n5103), .B1(n6252), .B2(n6297), 
        .B3(n6052), .ZN(n4735) );
  AOI22_X1 U5810 ( .A1(n6256), .A2(n4735), .B1(n6312), .B2(n4853), .ZN(n4715)
         );
  INV_X1 U5811 ( .A(n6266), .ZN(n6303) );
  AOI22_X1 U5812 ( .A1(n6304), .A2(n4736), .B1(n6303), .B2(n4977), .ZN(n4714)
         );
  OAI211_X1 U5813 ( .C1(n4740), .C2(n4716), .A(n4715), .B(n4714), .ZN(U3132)
         );
  AOI22_X1 U5814 ( .A1(n6374), .A2(n4735), .B1(n6336), .B2(n4853), .ZN(n4718)
         );
  INV_X1 U5815 ( .A(n6283), .ZN(n6370) );
  AOI22_X1 U5816 ( .A1(n6372), .A2(n4736), .B1(n6370), .B2(n4977), .ZN(n4717)
         );
  OAI211_X1 U5817 ( .C1(n4740), .C2(n4719), .A(n4718), .B(n4717), .ZN(U3137)
         );
  INV_X1 U5818 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4722) );
  AOI22_X1 U5819 ( .A1(n6277), .A2(n4735), .B1(n6330), .B2(n4853), .ZN(n4721)
         );
  INV_X1 U5820 ( .A(n6280), .ZN(n6332) );
  AOI22_X1 U5821 ( .A1(n6331), .A2(n4736), .B1(n6332), .B2(n4977), .ZN(n4720)
         );
  OAI211_X1 U5822 ( .C1(n4740), .C2(n4722), .A(n4721), .B(n4720), .ZN(U3136)
         );
  INV_X1 U5823 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4725) );
  AOI22_X1 U5824 ( .A1(n6284), .A2(n4735), .B1(n6340), .B2(n4853), .ZN(n4724)
         );
  INV_X1 U5825 ( .A(n6287), .ZN(n6342) );
  AOI22_X1 U5826 ( .A1(n6341), .A2(n4736), .B1(n6342), .B2(n4977), .ZN(n4723)
         );
  OAI211_X1 U5827 ( .C1(n4740), .C2(n4725), .A(n4724), .B(n4723), .ZN(U3138)
         );
  AOI22_X1 U5828 ( .A1(n6365), .A2(n2988), .B1(n6326), .B2(n4853), .ZN(n4727)
         );
  INV_X1 U5829 ( .A(n6276), .ZN(n6363) );
  AOI22_X1 U5830 ( .A1(n6364), .A2(n4736), .B1(n6363), .B2(n4977), .ZN(n4726)
         );
  OAI211_X1 U5831 ( .C1(n4740), .C2(n4728), .A(n4727), .B(n4726), .ZN(U3135)
         );
  INV_X1 U5832 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4731) );
  AOI22_X1 U5833 ( .A1(n6290), .A2(n2988), .B1(n6347), .B2(n4853), .ZN(n4730)
         );
  INV_X1 U5834 ( .A(n6296), .ZN(n6351) );
  AOI22_X1 U5835 ( .A1(n6349), .A2(n4736), .B1(n6351), .B2(n4977), .ZN(n4729)
         );
  OAI211_X1 U5836 ( .C1(n4740), .C2(n4731), .A(n4730), .B(n4729), .ZN(U3139)
         );
  INV_X1 U5837 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4734) );
  AOI22_X1 U5838 ( .A1(n6359), .A2(n2988), .B1(n6316), .B2(n4853), .ZN(n4733)
         );
  INV_X1 U5839 ( .A(n6269), .ZN(n6357) );
  AOI22_X1 U5840 ( .A1(n6358), .A2(n4736), .B1(n6357), .B2(n4977), .ZN(n4732)
         );
  OAI211_X1 U5841 ( .C1(n4740), .C2(n4734), .A(n4733), .B(n4732), .ZN(U3133)
         );
  INV_X1 U5842 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4739) );
  AOI22_X1 U5843 ( .A1(n6270), .A2(n2988), .B1(n6320), .B2(n4853), .ZN(n4738)
         );
  INV_X1 U5844 ( .A(n6273), .ZN(n6322) );
  AOI22_X1 U5845 ( .A1(n6321), .A2(n4736), .B1(n6322), .B2(n4977), .ZN(n4737)
         );
  OAI211_X1 U5846 ( .C1(n4740), .C2(n4739), .A(n4738), .B(n4737), .ZN(U3134)
         );
  OAI21_X1 U5847 ( .B1(n4765), .B2(n5852), .A(n6310), .ZN(n4746) );
  NOR2_X1 U5848 ( .A1(n4742), .A2(n6263), .ZN(n6371) );
  AOI21_X1 U5849 ( .B1(n4768), .B2(n5361), .A(n6371), .ZN(n4743) );
  NAND3_X1 U5850 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n5030), .ZN(n4769) );
  OAI22_X1 U5851 ( .A1(n4746), .A2(n4743), .B1(n4769), .B2(n5069), .ZN(n6373)
         );
  INV_X1 U5852 ( .A(n6373), .ZN(n4764) );
  INV_X1 U5853 ( .A(n4743), .ZN(n4745) );
  AOI21_X1 U5854 ( .B1(n6297), .B2(n4769), .A(n5065), .ZN(n4744) );
  OAI21_X1 U5855 ( .B1(n4746), .B2(n4745), .A(n4744), .ZN(n6375) );
  NAND2_X1 U5856 ( .A1(n2963), .A2(n5098), .ZN(n4747) );
  NAND2_X1 U5857 ( .A1(n2963), .A2(n6250), .ZN(n4748) );
  AOI22_X1 U5858 ( .A1(n6321), .A2(n6371), .B1(n6322), .B2(n6369), .ZN(n4749)
         );
  OAI21_X1 U5859 ( .B1(n6378), .B2(n5126), .A(n4749), .ZN(n4750) );
  AOI21_X1 U5860 ( .B1(INSTQUEUE_REG_11__2__SCAN_IN), .B2(n6375), .A(n4750), 
        .ZN(n4751) );
  OAI21_X1 U5861 ( .B1(n4764), .B2(n6325), .A(n4751), .ZN(U3110) );
  AOI22_X1 U5862 ( .A1(n6304), .A2(n6371), .B1(n6303), .B2(n6369), .ZN(n4752)
         );
  OAI21_X1 U5863 ( .B1(n6378), .B2(n5118), .A(n4752), .ZN(n4753) );
  AOI21_X1 U5864 ( .B1(INSTQUEUE_REG_11__0__SCAN_IN), .B2(n6375), .A(n4753), 
        .ZN(n4754) );
  OAI21_X1 U5865 ( .B1(n4764), .B2(n6315), .A(n4754), .ZN(U3108) );
  AOI22_X1 U5866 ( .A1(n6341), .A2(n6371), .B1(n6342), .B2(n6369), .ZN(n4755)
         );
  OAI21_X1 U5867 ( .B1(n6378), .B2(n5108), .A(n4755), .ZN(n4756) );
  AOI21_X1 U5868 ( .B1(INSTQUEUE_REG_11__6__SCAN_IN), .B2(n6375), .A(n4756), 
        .ZN(n4757) );
  OAI21_X1 U5869 ( .B1(n4764), .B2(n6345), .A(n4757), .ZN(U3114) );
  AOI22_X1 U5870 ( .A1(n6331), .A2(n6371), .B1(n6332), .B2(n6369), .ZN(n4758)
         );
  OAI21_X1 U5871 ( .B1(n6378), .B2(n5130), .A(n4758), .ZN(n4759) );
  AOI21_X1 U5872 ( .B1(INSTQUEUE_REG_11__4__SCAN_IN), .B2(n6375), .A(n4759), 
        .ZN(n4760) );
  OAI21_X1 U5873 ( .B1(n4764), .B2(n6335), .A(n4760), .ZN(U3112) );
  AOI22_X1 U5874 ( .A1(n6349), .A2(n6371), .B1(n6351), .B2(n6369), .ZN(n4761)
         );
  OAI21_X1 U5875 ( .B1(n6378), .B2(n5122), .A(n4761), .ZN(n4762) );
  AOI21_X1 U5876 ( .B1(INSTQUEUE_REG_11__7__SCAN_IN), .B2(n6375), .A(n4762), 
        .ZN(n4763) );
  OAI21_X1 U5877 ( .B1(n4764), .B2(n6355), .A(n4763), .ZN(U3115) );
  NAND2_X1 U5878 ( .A1(n4803), .A2(n6250), .ZN(n4773) );
  NAND2_X1 U5879 ( .A1(n4773), .A2(n6378), .ZN(n4766) );
  AOI21_X1 U5880 ( .B1(n4766), .B2(STATEBS16_REG_SCAN_IN), .A(n6297), .ZN(
        n4771) );
  INV_X1 U5881 ( .A(n6259), .ZN(n4918) );
  NOR2_X1 U5882 ( .A1(n4918), .A2(n6263), .ZN(n4767) );
  AOI22_X1 U5883 ( .A1(n4771), .A2(n4768), .B1(n6253), .B2(n4767), .ZN(n4800)
         );
  NOR2_X1 U5884 ( .A1(n6254), .A2(n6258), .ZN(n5227) );
  INV_X1 U5885 ( .A(n4768), .ZN(n4770) );
  OR2_X1 U5886 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4769), .ZN(n4796)
         );
  AOI22_X1 U5887 ( .A1(n4771), .A2(n4770), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n4796), .ZN(n4772) );
  NAND2_X1 U5888 ( .A1(n4795), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4776)
         );
  OAI22_X1 U5889 ( .A1(n4796), .A2(n4857), .B1(n6378), .B2(n6273), .ZN(n4774)
         );
  AOI21_X1 U5890 ( .B1(n4867), .B2(n6320), .A(n4774), .ZN(n4775) );
  OAI211_X1 U5891 ( .C1(n4800), .C2(n6325), .A(n4776), .B(n4775), .ZN(U3102)
         );
  NAND2_X1 U5892 ( .A1(n4795), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4779)
         );
  OAI22_X1 U5893 ( .A1(n4796), .A2(n4835), .B1(n6378), .B2(n6287), .ZN(n4777)
         );
  AOI21_X1 U5894 ( .B1(n4867), .B2(n6340), .A(n4777), .ZN(n4778) );
  OAI211_X1 U5895 ( .C1(n4800), .C2(n6345), .A(n4779), .B(n4778), .ZN(U3106)
         );
  NAND2_X1 U5896 ( .A1(n4795), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4782)
         );
  OAI22_X1 U5897 ( .A1(n4796), .A2(n4841), .B1(n6378), .B2(n6280), .ZN(n4780)
         );
  AOI21_X1 U5898 ( .B1(n4867), .B2(n6330), .A(n4780), .ZN(n4781) );
  OAI211_X1 U5899 ( .C1(n4800), .C2(n6335), .A(n4782), .B(n4781), .ZN(U3104)
         );
  NAND2_X1 U5900 ( .A1(n4795), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4785)
         );
  OAI22_X1 U5901 ( .A1(n4796), .A2(n4844), .B1(n6378), .B2(n6283), .ZN(n4783)
         );
  AOI21_X1 U5902 ( .B1(n4867), .B2(n6336), .A(n4783), .ZN(n4784) );
  OAI211_X1 U5903 ( .C1(n4800), .C2(n6339), .A(n4785), .B(n4784), .ZN(U3105)
         );
  NAND2_X1 U5904 ( .A1(n4795), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4788)
         );
  OAI22_X1 U5905 ( .A1(n4796), .A2(n4828), .B1(n6378), .B2(n6276), .ZN(n4786)
         );
  AOI21_X1 U5906 ( .B1(n4867), .B2(n6326), .A(n4786), .ZN(n4787) );
  OAI211_X1 U5907 ( .C1(n4800), .C2(n6329), .A(n4788), .B(n4787), .ZN(U3103)
         );
  NAND2_X1 U5908 ( .A1(n4795), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4791)
         );
  OAI22_X1 U5909 ( .A1(n4796), .A2(n4850), .B1(n6378), .B2(n6269), .ZN(n4789)
         );
  AOI21_X1 U5910 ( .B1(n4867), .B2(n6316), .A(n4789), .ZN(n4790) );
  OAI211_X1 U5911 ( .C1(n4800), .C2(n6319), .A(n4791), .B(n4790), .ZN(U3101)
         );
  NAND2_X1 U5912 ( .A1(n4795), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4794)
         );
  OAI22_X1 U5913 ( .A1(n4796), .A2(n4838), .B1(n6378), .B2(n6296), .ZN(n4792)
         );
  AOI21_X1 U5914 ( .B1(n4867), .B2(n6347), .A(n4792), .ZN(n4793) );
  OAI211_X1 U5915 ( .C1(n4800), .C2(n6355), .A(n4794), .B(n4793), .ZN(U3107)
         );
  NAND2_X1 U5916 ( .A1(n4795), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4799)
         );
  OAI22_X1 U5917 ( .A1(n4847), .A2(n4796), .B1(n6378), .B2(n6266), .ZN(n4797)
         );
  AOI21_X1 U5918 ( .B1(n4867), .B2(n6312), .A(n4797), .ZN(n4798) );
  OAI211_X1 U5919 ( .C1(n4800), .C2(n6315), .A(n4799), .B(n4798), .ZN(U3100)
         );
  XNOR2_X1 U5920 ( .A(n4802), .B(n4801), .ZN(n6197) );
  OAI222_X1 U5921 ( .A1(n5579), .A2(n5197), .B1(n6076), .B2(n5191), .C1(n5578), 
        .C2(n6197), .ZN(U2851) );
  INV_X1 U5922 ( .A(n2963), .ZN(n5024) );
  NAND3_X1 U5923 ( .A1(n4804), .A2(n5024), .A3(STATEBS16_REG_SCAN_IN), .ZN(
        n4805) );
  NAND2_X1 U5924 ( .A1(n4805), .A2(n6310), .ZN(n4809) );
  AND2_X1 U5925 ( .A1(n5361), .A2(n2961), .ZN(n4949) );
  OR2_X1 U5926 ( .A1(n4418), .A2(n4806), .ZN(n5027) );
  INV_X1 U5927 ( .A(n5027), .ZN(n5094) );
  NAND3_X1 U5928 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5030), .A3(n6394), .ZN(n5093) );
  NOR2_X1 U5929 ( .A1(n6388), .A2(n5093), .ZN(n4866) );
  AOI21_X1 U5930 ( .B1(n4949), .B2(n5094), .A(n4866), .ZN(n4810) );
  INV_X1 U5931 ( .A(n4810), .ZN(n4808) );
  AOI21_X1 U5932 ( .B1(n6297), .B2(n5093), .A(n5065), .ZN(n4807) );
  OAI21_X1 U5933 ( .B1(n4809), .B2(n4808), .A(n4807), .ZN(n4865) );
  OAI22_X1 U5934 ( .A1(n4810), .A2(n4809), .B1(n5069), .B2(n5093), .ZN(n4864)
         );
  AOI22_X1 U5935 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4865), .B1(n6256), 
        .B2(n4864), .ZN(n4812) );
  AOI22_X1 U5936 ( .A1(n4867), .A2(n6303), .B1(n6304), .B2(n4866), .ZN(n4811)
         );
  OAI211_X1 U5937 ( .C1(n5118), .C2(n5137), .A(n4812), .B(n4811), .ZN(U3092)
         );
  AOI22_X1 U5938 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4865), .B1(n6365), 
        .B2(n4864), .ZN(n4814) );
  AOI22_X1 U5939 ( .A1(n4867), .A2(n6363), .B1(n6364), .B2(n4866), .ZN(n4813)
         );
  OAI211_X1 U5940 ( .C1(n6368), .C2(n5137), .A(n4814), .B(n4813), .ZN(U3095)
         );
  NAND2_X1 U5941 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4815), .ZN(n4907) );
  NOR2_X1 U5942 ( .A1(n6388), .A2(n4907), .ZN(n4816) );
  INV_X1 U5943 ( .A(n4816), .ZN(n4856) );
  INV_X1 U5944 ( .A(n4915), .ZN(n4817) );
  AOI21_X1 U5945 ( .B1(n4949), .B2(n4817), .A(n4816), .ZN(n4824) );
  INV_X1 U5946 ( .A(n4824), .ZN(n4820) );
  NAND2_X1 U5947 ( .A1(n6310), .A2(n4818), .ZN(n4823) );
  AOI21_X1 U5948 ( .B1(n6297), .B2(n4907), .A(n5065), .ZN(n4819) );
  OAI21_X1 U5949 ( .B1(n4820), .B2(n4823), .A(n4819), .ZN(n4852) );
  NAND2_X1 U5950 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4821) );
  OAI22_X1 U5951 ( .A1(n4824), .A2(n4823), .B1(n4822), .B2(n4821), .ZN(n4851)
         );
  AOI22_X1 U5952 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4852), .B1(n6365), 
        .B2(n4851), .ZN(n4827) );
  AOI22_X1 U5953 ( .A1(n6326), .A2(n4913), .B1(n4853), .B2(n6363), .ZN(n4826)
         );
  OAI211_X1 U5954 ( .C1(n4828), .C2(n4856), .A(n4827), .B(n4826), .ZN(U3127)
         );
  AOI22_X1 U5955 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4865), .B1(n6270), 
        .B2(n4864), .ZN(n4830) );
  AOI22_X1 U5956 ( .A1(n4867), .A2(n6322), .B1(n6321), .B2(n4866), .ZN(n4829)
         );
  OAI211_X1 U5957 ( .C1(n5126), .C2(n5137), .A(n4830), .B(n4829), .ZN(U3094)
         );
  AOI22_X1 U5958 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4865), .B1(n6359), 
        .B2(n4864), .ZN(n4832) );
  AOI22_X1 U5959 ( .A1(n4867), .A2(n6357), .B1(n6358), .B2(n4866), .ZN(n4831)
         );
  OAI211_X1 U5960 ( .C1(n6362), .C2(n5137), .A(n4832), .B(n4831), .ZN(U3093)
         );
  AOI22_X1 U5961 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4852), .B1(n6284), 
        .B2(n4851), .ZN(n4834) );
  AOI22_X1 U5962 ( .A1(n6340), .A2(n4913), .B1(n4853), .B2(n6342), .ZN(n4833)
         );
  OAI211_X1 U5963 ( .C1(n4835), .C2(n4856), .A(n4834), .B(n4833), .ZN(U3130)
         );
  AOI22_X1 U5964 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4852), .B1(n6290), 
        .B2(n4851), .ZN(n4837) );
  AOI22_X1 U5965 ( .A1(n6347), .A2(n4913), .B1(n4853), .B2(n6351), .ZN(n4836)
         );
  OAI211_X1 U5966 ( .C1(n4838), .C2(n4856), .A(n4837), .B(n4836), .ZN(U3131)
         );
  AOI22_X1 U5967 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4852), .B1(n6277), 
        .B2(n4851), .ZN(n4840) );
  AOI22_X1 U5968 ( .A1(n6330), .A2(n4913), .B1(n4853), .B2(n6332), .ZN(n4839)
         );
  OAI211_X1 U5969 ( .C1(n4841), .C2(n4856), .A(n4840), .B(n4839), .ZN(U3128)
         );
  AOI22_X1 U5970 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4852), .B1(n6374), 
        .B2(n4851), .ZN(n4843) );
  AOI22_X1 U5971 ( .A1(n6336), .A2(n4913), .B1(n4853), .B2(n6370), .ZN(n4842)
         );
  OAI211_X1 U5972 ( .C1(n4844), .C2(n4856), .A(n4843), .B(n4842), .ZN(U3129)
         );
  AOI22_X1 U5973 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4852), .B1(n6256), 
        .B2(n4851), .ZN(n4846) );
  AOI22_X1 U5974 ( .A1(n6312), .A2(n4913), .B1(n4853), .B2(n6303), .ZN(n4845)
         );
  OAI211_X1 U5975 ( .C1(n4847), .C2(n4856), .A(n4846), .B(n4845), .ZN(U3124)
         );
  AOI22_X1 U5976 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4852), .B1(n6359), 
        .B2(n4851), .ZN(n4849) );
  AOI22_X1 U5977 ( .A1(n6316), .A2(n4913), .B1(n4853), .B2(n6357), .ZN(n4848)
         );
  OAI211_X1 U5978 ( .C1(n4850), .C2(n4856), .A(n4849), .B(n4848), .ZN(U3125)
         );
  AOI22_X1 U5979 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4852), .B1(n6270), 
        .B2(n4851), .ZN(n4855) );
  AOI22_X1 U5980 ( .A1(n6320), .A2(n4913), .B1(n4853), .B2(n6322), .ZN(n4854)
         );
  OAI211_X1 U5981 ( .C1(n4857), .C2(n4856), .A(n4855), .B(n4854), .ZN(U3126)
         );
  AOI22_X1 U5982 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4865), .B1(n6277), 
        .B2(n4864), .ZN(n4859) );
  AOI22_X1 U5983 ( .A1(n4867), .A2(n6332), .B1(n6331), .B2(n4866), .ZN(n4858)
         );
  OAI211_X1 U5984 ( .C1(n5130), .C2(n5137), .A(n4859), .B(n4858), .ZN(U3096)
         );
  AOI22_X1 U5985 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4865), .B1(n6374), 
        .B2(n4864), .ZN(n4861) );
  AOI22_X1 U5986 ( .A1(n4867), .A2(n6370), .B1(n6372), .B2(n4866), .ZN(n4860)
         );
  OAI211_X1 U5987 ( .C1(n6379), .C2(n5137), .A(n4861), .B(n4860), .ZN(U3097)
         );
  AOI22_X1 U5988 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4865), .B1(n6290), 
        .B2(n4864), .ZN(n4863) );
  AOI22_X1 U5989 ( .A1(n4867), .A2(n6351), .B1(n6349), .B2(n4866), .ZN(n4862)
         );
  OAI211_X1 U5990 ( .C1(n5122), .C2(n5137), .A(n4863), .B(n4862), .ZN(U3099)
         );
  AOI22_X1 U5991 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4865), .B1(n6284), 
        .B2(n4864), .ZN(n4869) );
  AOI22_X1 U5992 ( .A1(n4867), .A2(n6342), .B1(n6341), .B2(n4866), .ZN(n4868)
         );
  OAI211_X1 U5993 ( .C1(n5108), .C2(n5137), .A(n4869), .B(n4868), .ZN(U3098)
         );
  NOR2_X1 U5994 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4870), .ZN(n4903)
         );
  INV_X1 U5995 ( .A(n4903), .ZN(n4873) );
  INV_X1 U5996 ( .A(n4908), .ZN(n4871) );
  OAI21_X1 U5997 ( .B1(n3075), .B2(n5069), .A(n4872), .ZN(n5031) );
  AOI211_X1 U5998 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4873), .A(n6259), .B(
        n5031), .ZN(n4877) );
  OAI211_X1 U5999 ( .C1(n4906), .C2(n5028), .A(n4875), .B(n4874), .ZN(n4876)
         );
  NAND2_X1 U6000 ( .A1(n4877), .A2(n4876), .ZN(n4899) );
  NAND2_X1 U6001 ( .A1(n4899), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4880) );
  NOR2_X1 U6002 ( .A1(n4915), .A2(n6297), .ZN(n4909) );
  AOI22_X1 U6003 ( .A1(n4909), .A2(n6052), .B1(n6254), .B2(n3075), .ZN(n4901)
         );
  OAI22_X1 U6004 ( .A1(n6335), .A2(n4901), .B1(n6280), .B2(n4900), .ZN(n4878)
         );
  AOI21_X1 U6005 ( .B1(n6331), .B2(n4903), .A(n4878), .ZN(n4879) );
  OAI211_X1 U6006 ( .C1(n4906), .C2(n5130), .A(n4880), .B(n4879), .ZN(U3056)
         );
  NAND2_X1 U6007 ( .A1(n4899), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4883) );
  OAI22_X1 U6008 ( .A1(n6339), .A2(n4901), .B1(n6283), .B2(n4900), .ZN(n4881)
         );
  AOI21_X1 U6009 ( .B1(n6372), .B2(n4903), .A(n4881), .ZN(n4882) );
  OAI211_X1 U6010 ( .C1(n4906), .C2(n6379), .A(n4883), .B(n4882), .ZN(U3057)
         );
  NAND2_X1 U6011 ( .A1(n4899), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4886) );
  OAI22_X1 U6012 ( .A1(n6315), .A2(n4901), .B1(n6266), .B2(n4900), .ZN(n4884)
         );
  AOI21_X1 U6013 ( .B1(n6304), .B2(n4903), .A(n4884), .ZN(n4885) );
  OAI211_X1 U6014 ( .C1(n4906), .C2(n5118), .A(n4886), .B(n4885), .ZN(U3052)
         );
  NAND2_X1 U6015 ( .A1(n4899), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4889) );
  OAI22_X1 U6016 ( .A1(n6329), .A2(n4901), .B1(n6276), .B2(n4900), .ZN(n4887)
         );
  AOI21_X1 U6017 ( .B1(n6364), .B2(n4903), .A(n4887), .ZN(n4888) );
  OAI211_X1 U6018 ( .C1(n4906), .C2(n6368), .A(n4889), .B(n4888), .ZN(U3055)
         );
  NAND2_X1 U6019 ( .A1(n4899), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4892) );
  OAI22_X1 U6020 ( .A1(n6325), .A2(n4901), .B1(n6273), .B2(n4900), .ZN(n4890)
         );
  AOI21_X1 U6021 ( .B1(n6321), .B2(n4903), .A(n4890), .ZN(n4891) );
  OAI211_X1 U6022 ( .C1(n4906), .C2(n5126), .A(n4892), .B(n4891), .ZN(U3054)
         );
  NAND2_X1 U6023 ( .A1(n4899), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4895) );
  OAI22_X1 U6024 ( .A1(n6319), .A2(n4901), .B1(n6269), .B2(n4900), .ZN(n4893)
         );
  AOI21_X1 U6025 ( .B1(n6358), .B2(n4903), .A(n4893), .ZN(n4894) );
  OAI211_X1 U6026 ( .C1(n4906), .C2(n6362), .A(n4895), .B(n4894), .ZN(U3053)
         );
  NAND2_X1 U6027 ( .A1(n4899), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4898) );
  OAI22_X1 U6028 ( .A1(n6345), .A2(n4901), .B1(n6287), .B2(n4900), .ZN(n4896)
         );
  AOI21_X1 U6029 ( .B1(n6341), .B2(n4903), .A(n4896), .ZN(n4897) );
  OAI211_X1 U6030 ( .C1(n4906), .C2(n5108), .A(n4898), .B(n4897), .ZN(U3058)
         );
  NAND2_X1 U6031 ( .A1(n4899), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4905) );
  OAI22_X1 U6032 ( .A1(n6355), .A2(n4901), .B1(n6296), .B2(n4900), .ZN(n4902)
         );
  AOI21_X1 U6033 ( .B1(n6349), .B2(n4903), .A(n4902), .ZN(n4904) );
  OAI211_X1 U6034 ( .C1(n4906), .C2(n5122), .A(n4905), .B(n4904), .ZN(U3059)
         );
  NOR2_X1 U6035 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4907), .ZN(n4942)
         );
  OR2_X1 U6036 ( .A1(n6253), .A2(n4908), .ZN(n4912) );
  INV_X1 U6037 ( .A(n4912), .ZN(n5095) );
  AOI22_X1 U6038 ( .A1(n4909), .A2(n2961), .B1(n6254), .B2(n5095), .ZN(n4940)
         );
  OAI22_X1 U6039 ( .A1(n6319), .A2(n4940), .B1(n6269), .B2(n4939), .ZN(n4910)
         );
  AOI21_X1 U6040 ( .B1(n6358), .B2(n4942), .A(n4910), .ZN(n4920) );
  AOI21_X1 U6041 ( .B1(n4912), .B2(STATE2_REG_2__SCAN_IN), .A(n4911), .ZN(
        n5102) );
  OAI21_X1 U6042 ( .B1(n6369), .B2(n4913), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4914) );
  OAI211_X1 U6043 ( .C1(n6052), .C2(n4915), .A(n4914), .B(n6310), .ZN(n4917)
         );
  OR2_X1 U6044 ( .A1(n4942), .A2(n6508), .ZN(n4916) );
  NAND4_X1 U6045 ( .A1(n5102), .A2(n4918), .A3(n4917), .A4(n4916), .ZN(n4943)
         );
  NAND2_X1 U6046 ( .A1(n4943), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4919)
         );
  OAI211_X1 U6047 ( .C1(n4946), .C2(n6362), .A(n4920), .B(n4919), .ZN(U3117)
         );
  OAI22_X1 U6048 ( .A1(n6315), .A2(n4940), .B1(n6266), .B2(n4939), .ZN(n4921)
         );
  AOI21_X1 U6049 ( .B1(n6304), .B2(n4942), .A(n4921), .ZN(n4923) );
  NAND2_X1 U6050 ( .A1(n4943), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4922)
         );
  OAI211_X1 U6051 ( .C1(n4946), .C2(n5118), .A(n4923), .B(n4922), .ZN(U3116)
         );
  OAI22_X1 U6052 ( .A1(n6325), .A2(n4940), .B1(n6273), .B2(n4939), .ZN(n4924)
         );
  AOI21_X1 U6053 ( .B1(n6321), .B2(n4942), .A(n4924), .ZN(n4926) );
  NAND2_X1 U6054 ( .A1(n4943), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4925)
         );
  OAI211_X1 U6055 ( .C1(n4946), .C2(n5126), .A(n4926), .B(n4925), .ZN(U3118)
         );
  OAI22_X1 U6056 ( .A1(n6355), .A2(n4940), .B1(n6296), .B2(n4939), .ZN(n4927)
         );
  AOI21_X1 U6057 ( .B1(n6349), .B2(n4942), .A(n4927), .ZN(n4929) );
  NAND2_X1 U6058 ( .A1(n4943), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4928)
         );
  OAI211_X1 U6059 ( .C1(n4946), .C2(n5122), .A(n4929), .B(n4928), .ZN(U3123)
         );
  OAI22_X1 U6060 ( .A1(n6345), .A2(n4940), .B1(n6287), .B2(n4939), .ZN(n4930)
         );
  AOI21_X1 U6061 ( .B1(n6341), .B2(n4942), .A(n4930), .ZN(n4932) );
  NAND2_X1 U6062 ( .A1(n4943), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4931)
         );
  OAI211_X1 U6063 ( .C1(n4946), .C2(n5108), .A(n4932), .B(n4931), .ZN(U3122)
         );
  OAI22_X1 U6064 ( .A1(n6335), .A2(n4940), .B1(n6280), .B2(n4939), .ZN(n4933)
         );
  AOI21_X1 U6065 ( .B1(n6331), .B2(n4942), .A(n4933), .ZN(n4935) );
  NAND2_X1 U6066 ( .A1(n4943), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4934)
         );
  OAI211_X1 U6067 ( .C1(n4946), .C2(n5130), .A(n4935), .B(n4934), .ZN(U3120)
         );
  OAI22_X1 U6068 ( .A1(n6339), .A2(n4940), .B1(n6283), .B2(n4939), .ZN(n4936)
         );
  AOI21_X1 U6069 ( .B1(n6372), .B2(n4942), .A(n4936), .ZN(n4938) );
  NAND2_X1 U6070 ( .A1(n4943), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4937)
         );
  OAI211_X1 U6071 ( .C1(n4946), .C2(n6379), .A(n4938), .B(n4937), .ZN(U3121)
         );
  OAI22_X1 U6072 ( .A1(n6329), .A2(n4940), .B1(n6276), .B2(n4939), .ZN(n4941)
         );
  AOI21_X1 U6073 ( .B1(n6364), .B2(n4942), .A(n4941), .ZN(n4945) );
  NAND2_X1 U6074 ( .A1(n4943), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4944)
         );
  OAI211_X1 U6075 ( .C1(n4946), .C2(n6368), .A(n4945), .B(n4944), .ZN(U3119)
         );
  INV_X1 U6076 ( .A(n6252), .ZN(n4948) );
  INV_X1 U6077 ( .A(n4947), .ZN(n4978) );
  AOI21_X1 U6078 ( .B1(n4949), .B2(n4948), .A(n4978), .ZN(n4954) );
  OAI21_X1 U6079 ( .B1(n4955), .B2(n6139), .A(n5225), .ZN(n4952) );
  NOR2_X1 U6080 ( .A1(n6310), .A2(n4950), .ZN(n4951) );
  AOI211_X2 U6081 ( .C1(n4954), .C2(n4952), .A(n4951), .B(n5065), .ZN(n4982)
         );
  INV_X1 U6082 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4958) );
  OAI22_X1 U6083 ( .A1(n4954), .A2(n6297), .B1(n4953), .B2(n5069), .ZN(n4976)
         );
  AOI22_X1 U6084 ( .A1(n6277), .A2(n4976), .B1(n6332), .B2(n5035), .ZN(n4957)
         );
  AOI22_X1 U6085 ( .A1(n6331), .A2(n4978), .B1(n6330), .B2(n4977), .ZN(n4956)
         );
  OAI211_X1 U6086 ( .C1(n4982), .C2(n4958), .A(n4957), .B(n4956), .ZN(U3144)
         );
  INV_X1 U6087 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4961) );
  AOI22_X1 U6088 ( .A1(n6374), .A2(n4976), .B1(n6370), .B2(n5035), .ZN(n4960)
         );
  AOI22_X1 U6089 ( .A1(n6372), .A2(n4978), .B1(n6336), .B2(n4977), .ZN(n4959)
         );
  OAI211_X1 U6090 ( .C1(n4982), .C2(n4961), .A(n4960), .B(n4959), .ZN(U3145)
         );
  INV_X1 U6091 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4964) );
  AOI22_X1 U6092 ( .A1(n6256), .A2(n4976), .B1(n6303), .B2(n5035), .ZN(n4963)
         );
  AOI22_X1 U6093 ( .A1(n6304), .A2(n4978), .B1(n6312), .B2(n4977), .ZN(n4962)
         );
  OAI211_X1 U6094 ( .C1(n4982), .C2(n4964), .A(n4963), .B(n4962), .ZN(U3140)
         );
  INV_X1 U6095 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4967) );
  AOI22_X1 U6096 ( .A1(n6359), .A2(n4976), .B1(n6357), .B2(n5035), .ZN(n4966)
         );
  AOI22_X1 U6097 ( .A1(n6358), .A2(n4978), .B1(n6316), .B2(n4977), .ZN(n4965)
         );
  OAI211_X1 U6098 ( .C1(n4982), .C2(n4967), .A(n4966), .B(n4965), .ZN(U3141)
         );
  INV_X1 U6099 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4970) );
  AOI22_X1 U6100 ( .A1(n6365), .A2(n4976), .B1(n6363), .B2(n5035), .ZN(n4969)
         );
  AOI22_X1 U6101 ( .A1(n6364), .A2(n4978), .B1(n6326), .B2(n4977), .ZN(n4968)
         );
  OAI211_X1 U6102 ( .C1(n4982), .C2(n4970), .A(n4969), .B(n4968), .ZN(U3143)
         );
  AOI22_X1 U6103 ( .A1(n6270), .A2(n4976), .B1(n6322), .B2(n5035), .ZN(n4972)
         );
  AOI22_X1 U6104 ( .A1(n6321), .A2(n4978), .B1(n6320), .B2(n4977), .ZN(n4971)
         );
  OAI211_X1 U6105 ( .C1(n4982), .C2(n6568), .A(n4972), .B(n4971), .ZN(U3142)
         );
  INV_X1 U6106 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4975) );
  AOI22_X1 U6107 ( .A1(n6290), .A2(n4976), .B1(n6351), .B2(n5035), .ZN(n4974)
         );
  AOI22_X1 U6108 ( .A1(n6349), .A2(n4978), .B1(n6347), .B2(n4977), .ZN(n4973)
         );
  OAI211_X1 U6109 ( .C1(n4982), .C2(n4975), .A(n4974), .B(n4973), .ZN(U3147)
         );
  INV_X1 U6110 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4981) );
  AOI22_X1 U6111 ( .A1(n6284), .A2(n4976), .B1(n6342), .B2(n5035), .ZN(n4980)
         );
  AOI22_X1 U6112 ( .A1(n6341), .A2(n4978), .B1(n6340), .B2(n4977), .ZN(n4979)
         );
  OAI211_X1 U6113 ( .C1(n4982), .C2(n4981), .A(n4980), .B(n4979), .ZN(U3146)
         );
  NOR3_X1 U6114 ( .A1(n6421), .A2(n6508), .A3(n6430), .ZN(n6413) );
  OR3_X1 U6115 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6425), .A3(n5362), .ZN(n4983) );
  NAND2_X1 U6116 ( .A1(n6196), .A2(n4983), .ZN(n4984) );
  OR2_X1 U6117 ( .A1(n6413), .A2(n4984), .ZN(n4985) );
  NAND2_X1 U6118 ( .A1(n5378), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4986) );
  INV_X1 U6119 ( .A(n4986), .ZN(n4987) );
  INV_X1 U6120 ( .A(n4989), .ZN(n5009) );
  NOR2_X1 U6121 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6407) );
  NAND2_X1 U6122 ( .A1(n6408), .A2(n6407), .ZN(n4990) );
  NAND2_X1 U6123 ( .A1(n3335), .A2(n4990), .ZN(n5374) );
  INV_X1 U6124 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5528) );
  INV_X1 U6125 ( .A(n6407), .ZN(n4997) );
  NAND3_X1 U6126 ( .A1(n4993), .A2(n5528), .A3(n4997), .ZN(n4991) );
  AND2_X1 U6127 ( .A1(n5374), .A2(n4991), .ZN(n4992) );
  INV_X1 U6128 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6456) );
  NAND3_X1 U6129 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5166) );
  NOR2_X1 U6130 ( .A1(n6456), .A2(n5166), .ZN(n5153) );
  NAND2_X1 U6131 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5153), .ZN(n5002) );
  INV_X1 U6132 ( .A(n5002), .ZN(n4996) );
  NAND3_X1 U6133 ( .A1(n4994), .A2(n6407), .A3(n4993), .ZN(n4995) );
  NAND2_X1 U6134 ( .A1(n6016), .A2(n5378), .ZN(n5499) );
  INV_X1 U6135 ( .A(n5499), .ZN(n5888) );
  AOI21_X1 U6136 ( .B1(n5378), .B2(n4996), .A(n5888), .ZN(n6032) );
  NOR3_X1 U6137 ( .A1(n6016), .A2(n5002), .A3(REIP_REG_6__SCAN_IN), .ZN(n6031)
         );
  OAI21_X1 U6138 ( .B1(n6032), .B2(n6031), .A(REIP_REG_7__SCAN_IN), .ZN(n5006)
         );
  NAND3_X1 U6139 ( .A1(n4998), .A2(EBX_REG_31__SCAN_IN), .A3(n4997), .ZN(n4999) );
  INV_X1 U6140 ( .A(n5000), .ZN(n6207) );
  NAND2_X1 U6141 ( .A1(n5378), .A2(n5001), .ZN(n6033) );
  INV_X1 U6142 ( .A(n6016), .ZN(n6002) );
  INV_X1 U6143 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6531) );
  INV_X1 U6144 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6459) );
  NOR2_X1 U6145 ( .A1(n6459), .A2(n5002), .ZN(n5187) );
  NAND3_X1 U6146 ( .A1(n6002), .A2(n6531), .A3(n5187), .ZN(n5003) );
  OAI211_X1 U6147 ( .C1(n6035), .C2(n6628), .A(n6033), .B(n5003), .ZN(n5004)
         );
  AOI21_X1 U6148 ( .B1(n6047), .B2(n6207), .A(n5004), .ZN(n5005) );
  OAI211_X1 U6149 ( .C1(n5007), .C2(n6029), .A(n5006), .B(n5005), .ZN(n5008)
         );
  AOI21_X1 U6150 ( .B1(n6057), .B2(n5009), .A(n5008), .ZN(n5010) );
  OAI21_X1 U6151 ( .B1(n5011), .B2(n6024), .A(n5010), .ZN(U2820) );
  NAND2_X1 U6152 ( .A1(n4642), .A2(n5013), .ZN(n5014) );
  NAND2_X1 U6153 ( .A1(n5012), .A2(n5014), .ZN(n6066) );
  AOI22_X1 U6154 ( .A1(n5357), .A2(DATAI_9_), .B1(n6084), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n5015) );
  OAI21_X1 U6155 ( .B1(n6066), .B2(n5911), .A(n5015), .ZN(U2882) );
  OAI21_X1 U6156 ( .B1(n5018), .B2(n5017), .A(n5016), .ZN(n6200) );
  INV_X1 U6157 ( .A(n5197), .ZN(n5021) );
  AOI22_X1 U6158 ( .A1(n6161), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6240), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5019) );
  OAI21_X1 U6159 ( .B1(n5192), .B2(n6170), .A(n5019), .ZN(n5020) );
  AOI21_X1 U6160 ( .B1(n5021), .B2(n5681), .A(n5020), .ZN(n5022) );
  OAI21_X1 U6161 ( .B1(n6200), .B2(n6144), .A(n5022), .ZN(U2978) );
  NAND3_X1 U6162 ( .A1(n5025), .A2(n5024), .A3(n5023), .ZN(n5072) );
  INV_X1 U6163 ( .A(n5072), .ZN(n5026) );
  NOR2_X1 U6164 ( .A1(n2961), .A2(n5027), .ZN(n5064) );
  NOR2_X1 U6165 ( .A1(n5035), .A2(n6297), .ZN(n5029) );
  AOI21_X1 U6166 ( .B1(n5092), .B2(n5029), .A(n5028), .ZN(n5034) );
  NAND3_X1 U6167 ( .A1(n6263), .A2(n5030), .A3(n6394), .ZN(n5068) );
  NOR2_X1 U6168 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5068), .ZN(n5061)
         );
  INV_X1 U6169 ( .A(n5061), .ZN(n5032) );
  AOI211_X1 U6170 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5032), .A(n6254), .B(
        n5031), .ZN(n5033) );
  NAND2_X1 U6171 ( .A1(n5057), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5038) );
  AOI22_X1 U6172 ( .A1(n5064), .A2(n6310), .B1(n6259), .B2(n3075), .ZN(n5059)
         );
  OAI22_X1 U6173 ( .A1(n6325), .A2(n5059), .B1(n5126), .B2(n5058), .ZN(n5036)
         );
  AOI21_X1 U6174 ( .B1(n6321), .B2(n5061), .A(n5036), .ZN(n5037) );
  OAI211_X1 U6175 ( .C1(n5092), .C2(n6273), .A(n5038), .B(n5037), .ZN(U3022)
         );
  NAND2_X1 U6176 ( .A1(n5057), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5041) );
  OAI22_X1 U6177 ( .A1(n6315), .A2(n5059), .B1(n5118), .B2(n5058), .ZN(n5039)
         );
  AOI21_X1 U6178 ( .B1(n6304), .B2(n5061), .A(n5039), .ZN(n5040) );
  OAI211_X1 U6179 ( .C1(n5092), .C2(n6266), .A(n5041), .B(n5040), .ZN(U3020)
         );
  NAND2_X1 U6180 ( .A1(n5057), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5044) );
  OAI22_X1 U6181 ( .A1(n6339), .A2(n5059), .B1(n6379), .B2(n5058), .ZN(n5042)
         );
  AOI21_X1 U6182 ( .B1(n6372), .B2(n5061), .A(n5042), .ZN(n5043) );
  OAI211_X1 U6183 ( .C1(n5092), .C2(n6283), .A(n5044), .B(n5043), .ZN(U3025)
         );
  NAND2_X1 U6184 ( .A1(n5057), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5047) );
  OAI22_X1 U6185 ( .A1(n6319), .A2(n5059), .B1(n6362), .B2(n5058), .ZN(n5045)
         );
  AOI21_X1 U6186 ( .B1(n6358), .B2(n5061), .A(n5045), .ZN(n5046) );
  OAI211_X1 U6187 ( .C1(n5092), .C2(n6269), .A(n5047), .B(n5046), .ZN(U3021)
         );
  NAND2_X1 U6188 ( .A1(n5057), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5050) );
  OAI22_X1 U6189 ( .A1(n6355), .A2(n5059), .B1(n5122), .B2(n5058), .ZN(n5048)
         );
  AOI21_X1 U6190 ( .B1(n6349), .B2(n5061), .A(n5048), .ZN(n5049) );
  OAI211_X1 U6191 ( .C1(n5092), .C2(n6296), .A(n5050), .B(n5049), .ZN(U3027)
         );
  NAND2_X1 U6192 ( .A1(n5057), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5053) );
  OAI22_X1 U6193 ( .A1(n6335), .A2(n5059), .B1(n5130), .B2(n5058), .ZN(n5051)
         );
  AOI21_X1 U6194 ( .B1(n6331), .B2(n5061), .A(n5051), .ZN(n5052) );
  OAI211_X1 U6195 ( .C1(n5092), .C2(n6280), .A(n5053), .B(n5052), .ZN(U3024)
         );
  NAND2_X1 U6196 ( .A1(n5057), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5056) );
  OAI22_X1 U6197 ( .A1(n6329), .A2(n5059), .B1(n6368), .B2(n5058), .ZN(n5054)
         );
  AOI21_X1 U6198 ( .B1(n6364), .B2(n5061), .A(n5054), .ZN(n5055) );
  OAI211_X1 U6199 ( .C1(n5092), .C2(n6276), .A(n5056), .B(n5055), .ZN(U3023)
         );
  NAND2_X1 U6200 ( .A1(n5057), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5063) );
  OAI22_X1 U6201 ( .A1(n6345), .A2(n5059), .B1(n5108), .B2(n5058), .ZN(n5060)
         );
  AOI21_X1 U6202 ( .B1(n6341), .B2(n5061), .A(n5060), .ZN(n5062) );
  OAI211_X1 U6203 ( .C1(n5092), .C2(n6287), .A(n5063), .B(n5062), .ZN(U3026)
         );
  OAI21_X1 U6204 ( .B1(n5072), .B2(n6424), .A(n6310), .ZN(n5071) );
  NOR2_X1 U6205 ( .A1(n6388), .A2(n5068), .ZN(n5089) );
  AOI21_X1 U6206 ( .B1(n5064), .B2(n5361), .A(n5089), .ZN(n5070) );
  INV_X1 U6207 ( .A(n5070), .ZN(n5067) );
  AOI21_X1 U6208 ( .B1(n6297), .B2(n5068), .A(n5065), .ZN(n5066) );
  OAI21_X1 U6209 ( .B1(n5071), .B2(n5067), .A(n5066), .ZN(n5088) );
  OAI22_X1 U6210 ( .A1(n5071), .A2(n5070), .B1(n5069), .B2(n5068), .ZN(n5087)
         );
  AOI22_X1 U6211 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5088), .B1(n6374), 
        .B2(n5087), .ZN(n5074) );
  NOR2_X2 U6212 ( .A1(n5072), .A2(n5098), .ZN(n5256) );
  AOI22_X1 U6213 ( .A1(n5256), .A2(n6370), .B1(n6372), .B2(n5089), .ZN(n5073)
         );
  OAI211_X1 U6214 ( .C1(n6379), .C2(n5092), .A(n5074), .B(n5073), .ZN(U3033)
         );
  AOI22_X1 U6215 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5088), .B1(n6277), 
        .B2(n5087), .ZN(n5076) );
  AOI22_X1 U6216 ( .A1(n5256), .A2(n6332), .B1(n6331), .B2(n5089), .ZN(n5075)
         );
  OAI211_X1 U6217 ( .C1(n5130), .C2(n5092), .A(n5076), .B(n5075), .ZN(U3032)
         );
  AOI22_X1 U6218 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5088), .B1(n6270), 
        .B2(n5087), .ZN(n5078) );
  AOI22_X1 U6219 ( .A1(n5256), .A2(n6322), .B1(n6321), .B2(n5089), .ZN(n5077)
         );
  OAI211_X1 U6220 ( .C1(n5126), .C2(n5092), .A(n5078), .B(n5077), .ZN(U3030)
         );
  AOI22_X1 U6221 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5088), .B1(n6290), 
        .B2(n5087), .ZN(n5080) );
  AOI22_X1 U6222 ( .A1(n5256), .A2(n6351), .B1(n6349), .B2(n5089), .ZN(n5079)
         );
  OAI211_X1 U6223 ( .C1(n5122), .C2(n5092), .A(n5080), .B(n5079), .ZN(U3035)
         );
  AOI22_X1 U6224 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5088), .B1(n6256), 
        .B2(n5087), .ZN(n5082) );
  AOI22_X1 U6225 ( .A1(n5256), .A2(n6303), .B1(n6304), .B2(n5089), .ZN(n5081)
         );
  OAI211_X1 U6226 ( .C1(n5118), .C2(n5092), .A(n5082), .B(n5081), .ZN(U3028)
         );
  AOI22_X1 U6227 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5088), .B1(n6365), 
        .B2(n5087), .ZN(n5084) );
  AOI22_X1 U6228 ( .A1(n5256), .A2(n6363), .B1(n6364), .B2(n5089), .ZN(n5083)
         );
  OAI211_X1 U6229 ( .C1(n6368), .C2(n5092), .A(n5084), .B(n5083), .ZN(U3031)
         );
  AOI22_X1 U6230 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5088), .B1(n6284), 
        .B2(n5087), .ZN(n5086) );
  AOI22_X1 U6231 ( .A1(n5256), .A2(n6342), .B1(n6341), .B2(n5089), .ZN(n5085)
         );
  OAI211_X1 U6232 ( .C1(n5108), .C2(n5092), .A(n5086), .B(n5085), .ZN(U3034)
         );
  AOI22_X1 U6233 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5088), .B1(n6359), 
        .B2(n5087), .ZN(n5091) );
  AOI22_X1 U6234 ( .A1(n5256), .A2(n6357), .B1(n6358), .B2(n5089), .ZN(n5090)
         );
  OAI211_X1 U6235 ( .C1(n6362), .C2(n5092), .A(n5091), .B(n5090), .ZN(U3029)
         );
  NOR2_X1 U6236 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5093), .ZN(n5133)
         );
  AND2_X1 U6237 ( .A1(n5094), .A2(n2961), .ZN(n5100) );
  AOI22_X1 U6238 ( .A1(n5100), .A2(n6310), .B1(n6259), .B2(n5095), .ZN(n5131)
         );
  AND2_X1 U6239 ( .A1(n2963), .A2(n5096), .ZN(n5097) );
  NAND2_X1 U6240 ( .A1(n5857), .A2(n5097), .ZN(n6251) );
  OAI22_X1 U6241 ( .A1(n6339), .A2(n5131), .B1(n6379), .B2(n6302), .ZN(n5099)
         );
  AOI21_X1 U6242 ( .B1(n6372), .B2(n5133), .A(n5099), .ZN(n5107) );
  NAND3_X1 U6243 ( .A1(n5137), .A2(n6310), .A3(n6302), .ZN(n5101) );
  AOI21_X1 U6244 ( .B1(n5101), .B2(n5225), .A(n5100), .ZN(n5105) );
  OAI211_X1 U6245 ( .C1(n6508), .C2(n5133), .A(n5103), .B(n5102), .ZN(n5104)
         );
  NAND2_X1 U6246 ( .A1(n5134), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5106) );
  OAI211_X1 U6247 ( .C1(n5137), .C2(n6283), .A(n5107), .B(n5106), .ZN(U3089)
         );
  OAI22_X1 U6248 ( .A1(n6345), .A2(n5131), .B1(n5108), .B2(n6302), .ZN(n5109)
         );
  AOI21_X1 U6249 ( .B1(n6341), .B2(n5133), .A(n5109), .ZN(n5111) );
  NAND2_X1 U6250 ( .A1(n5134), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5110) );
  OAI211_X1 U6251 ( .C1(n5137), .C2(n6287), .A(n5111), .B(n5110), .ZN(U3090)
         );
  OAI22_X1 U6252 ( .A1(n6329), .A2(n5131), .B1(n6368), .B2(n6302), .ZN(n5112)
         );
  AOI21_X1 U6253 ( .B1(n6364), .B2(n5133), .A(n5112), .ZN(n5114) );
  NAND2_X1 U6254 ( .A1(n5134), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5113) );
  OAI211_X1 U6255 ( .C1(n5137), .C2(n6276), .A(n5114), .B(n5113), .ZN(U3087)
         );
  OAI22_X1 U6256 ( .A1(n6319), .A2(n5131), .B1(n6362), .B2(n6302), .ZN(n5115)
         );
  AOI21_X1 U6257 ( .B1(n6358), .B2(n5133), .A(n5115), .ZN(n5117) );
  NAND2_X1 U6258 ( .A1(n5134), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5116) );
  OAI211_X1 U6259 ( .C1(n5137), .C2(n6269), .A(n5117), .B(n5116), .ZN(U3085)
         );
  OAI22_X1 U6260 ( .A1(n6315), .A2(n5131), .B1(n5118), .B2(n6302), .ZN(n5119)
         );
  AOI21_X1 U6261 ( .B1(n6304), .B2(n5133), .A(n5119), .ZN(n5121) );
  NAND2_X1 U6262 ( .A1(n5134), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5120) );
  OAI211_X1 U6263 ( .C1(n5137), .C2(n6266), .A(n5121), .B(n5120), .ZN(U3084)
         );
  OAI22_X1 U6264 ( .A1(n6355), .A2(n5131), .B1(n5122), .B2(n6302), .ZN(n5123)
         );
  AOI21_X1 U6265 ( .B1(n6349), .B2(n5133), .A(n5123), .ZN(n5125) );
  NAND2_X1 U6266 ( .A1(n5134), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5124) );
  OAI211_X1 U6267 ( .C1(n5137), .C2(n6296), .A(n5125), .B(n5124), .ZN(U3091)
         );
  OAI22_X1 U6268 ( .A1(n6325), .A2(n5131), .B1(n5126), .B2(n6302), .ZN(n5127)
         );
  AOI21_X1 U6269 ( .B1(n6321), .B2(n5133), .A(n5127), .ZN(n5129) );
  NAND2_X1 U6270 ( .A1(n5134), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5128) );
  OAI211_X1 U6271 ( .C1(n5137), .C2(n6273), .A(n5129), .B(n5128), .ZN(U3086)
         );
  OAI22_X1 U6272 ( .A1(n6335), .A2(n5131), .B1(n5130), .B2(n6302), .ZN(n5132)
         );
  AOI21_X1 U6273 ( .B1(n6331), .B2(n5133), .A(n5132), .ZN(n5136) );
  NAND2_X1 U6274 ( .A1(n5134), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5135) );
  OAI211_X1 U6275 ( .C1(n5137), .C2(n6280), .A(n5136), .B(n5135), .ZN(U3088)
         );
  INV_X1 U6276 ( .A(n5138), .ZN(n5139) );
  AOI21_X1 U6277 ( .B1(n5140), .B2(n5012), .A(n5139), .ZN(n5267) );
  INV_X1 U6278 ( .A(n5267), .ZN(n5217) );
  AOI22_X1 U6279 ( .A1(n5357), .A2(DATAI_10_), .B1(n6084), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5141) );
  OAI21_X1 U6280 ( .B1(n5217), .B2(n5911), .A(n5141), .ZN(U2881) );
  OR2_X1 U6281 ( .A1(n5142), .A2(n6011), .ZN(n5143) );
  AND2_X1 U6282 ( .A1(n5143), .A2(n2984), .ZN(n5278) );
  INV_X1 U6283 ( .A(n5278), .ZN(n5210) );
  OAI222_X1 U6284 ( .A1(n5217), .A2(n5579), .B1(n6076), .B2(n3642), .C1(n5210), 
        .C2(n5578), .ZN(U2849) );
  INV_X1 U6285 ( .A(n5375), .ZN(n5144) );
  OR2_X1 U6286 ( .A1(n5375), .A2(n5145), .ZN(n6051) );
  NOR2_X1 U6287 ( .A1(n6016), .A2(REIP_REG_1__SCAN_IN), .ZN(n5202) );
  INV_X1 U6288 ( .A(n5378), .ZN(n5201) );
  AOI22_X1 U6289 ( .A1(n6046), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n5201), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5146) );
  OAI21_X1 U6290 ( .B1(n5988), .B2(n5147), .A(n5146), .ZN(n5148) );
  AOI211_X1 U6291 ( .C1(n6048), .C2(EBX_REG_1__SCAN_IN), .A(n5202), .B(n5148), 
        .ZN(n5149) );
  OAI21_X1 U6292 ( .B1(n5854), .B2(n6051), .A(n5149), .ZN(n5150) );
  AOI21_X1 U6293 ( .B1(n6057), .B2(n6623), .A(n5150), .ZN(n5151) );
  OAI21_X1 U6294 ( .B1(n6053), .B2(n5152), .A(n5151), .ZN(U2826) );
  INV_X1 U6295 ( .A(n6032), .ZN(n5159) );
  AOI21_X1 U6296 ( .B1(n6002), .B2(n5153), .A(REIP_REG_5__SCAN_IN), .ZN(n5158)
         );
  AOI21_X1 U6297 ( .B1(n6046), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n6020), 
        .ZN(n5154) );
  OAI21_X1 U6298 ( .B1(n5155), .B2(n5988), .A(n5154), .ZN(n5156) );
  AOI21_X1 U6299 ( .B1(n6048), .B2(EBX_REG_5__SCAN_IN), .A(n5156), .ZN(n5157)
         );
  OAI21_X1 U6300 ( .B1(n5159), .B2(n5158), .A(n5157), .ZN(n5160) );
  AOI21_X1 U6301 ( .B1(n6057), .B2(n5161), .A(n5160), .ZN(n5162) );
  OAI21_X1 U6302 ( .B1(n6053), .B2(n5163), .A(n5162), .ZN(U2822) );
  INV_X1 U6303 ( .A(n5164), .ZN(n5172) );
  OAI21_X1 U6304 ( .B1(n5201), .B2(n5166), .A(n5499), .ZN(n6060) );
  OAI22_X1 U6305 ( .A1(n6060), .A2(n6456), .B1(n6536), .B2(n6035), .ZN(n5165)
         );
  AOI211_X1 U6306 ( .C1(n6047), .C2(n6223), .A(n5165), .B(n6020), .ZN(n5169)
         );
  NOR3_X1 U6307 ( .A1(n6016), .A2(REIP_REG_4__SCAN_IN), .A3(n5166), .ZN(n5167)
         );
  AOI21_X1 U6308 ( .B1(n6048), .B2(EBX_REG_4__SCAN_IN), .A(n5167), .ZN(n5168)
         );
  OAI211_X1 U6309 ( .C1(n5170), .C2(n6051), .A(n5169), .B(n5168), .ZN(n5171)
         );
  AOI21_X1 U6310 ( .B1(n6057), .B2(n5172), .A(n5171), .ZN(n5173) );
  OAI21_X1 U6311 ( .B1(n6053), .B2(n5174), .A(n5173), .ZN(U2823) );
  NOR2_X1 U6312 ( .A1(n6051), .A2(n6299), .ZN(n5177) );
  OAI22_X1 U6313 ( .A1(n6626), .A2(n6029), .B1(n5988), .B2(n5175), .ZN(n5176)
         );
  AOI211_X1 U6314 ( .C1(REIP_REG_0__SCAN_IN), .C2(n5499), .A(n5177), .B(n5176), 
        .ZN(n5179) );
  OAI21_X1 U6315 ( .B1(n6057), .B2(n6046), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5178) );
  OAI211_X1 U6316 ( .C1(n6053), .C2(n5180), .A(n5179), .B(n5178), .ZN(U2827)
         );
  NAND2_X1 U6317 ( .A1(n5182), .A2(n5181), .ZN(n5183) );
  NAND2_X1 U6318 ( .A1(n6190), .A2(n6165), .ZN(n5186) );
  NAND2_X1 U6319 ( .A1(n6240), .A2(REIP_REG_9__SCAN_IN), .ZN(n6186) );
  OAI21_X1 U6320 ( .B1(n5725), .B2(n6018), .A(n6186), .ZN(n5184) );
  AOI21_X1 U6321 ( .B1(n5728), .B2(n6022), .A(n5184), .ZN(n5185) );
  OAI211_X1 U6322 ( .C1(n6139), .C2(n6066), .A(n5186), .B(n5185), .ZN(U2977)
         );
  INV_X1 U6323 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U6324 ( .A1(REIP_REG_7__SCAN_IN), .A2(n5187), .ZN(n5188) );
  NOR2_X1 U6325 ( .A1(n6462), .A2(n5188), .ZN(n6014) );
  OAI21_X1 U6326 ( .B1(n6016), .B2(n6014), .A(n5378), .ZN(n6021) );
  OAI21_X1 U6327 ( .B1(n6016), .B2(n5188), .A(n6462), .ZN(n5195) );
  NOR2_X1 U6328 ( .A1(n5988), .A2(n6197), .ZN(n5189) );
  AOI211_X1 U6329 ( .C1(n6046), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6020), 
        .B(n5189), .ZN(n5190) );
  OAI21_X1 U6330 ( .B1(n6029), .B2(n5191), .A(n5190), .ZN(n5194) );
  NOR2_X1 U6331 ( .A1(n6041), .A2(n5192), .ZN(n5193) );
  AOI211_X1 U6332 ( .C1(n6021), .C2(n5195), .A(n5194), .B(n5193), .ZN(n5196)
         );
  OAI21_X1 U6333 ( .B1(n6024), .B2(n5197), .A(n5196), .ZN(U2819) );
  XOR2_X1 U6334 ( .A(n5199), .B(n5198), .Z(n6238) );
  INV_X1 U6335 ( .A(n4418), .ZN(n5859) );
  INV_X1 U6336 ( .A(REIP_REG_2__SCAN_IN), .ZN(n5203) );
  NAND3_X1 U6337 ( .A1(n6002), .A2(REIP_REG_1__SCAN_IN), .A3(n5203), .ZN(n5200) );
  OAI21_X1 U6338 ( .B1(n6035), .B2(n6591), .A(n5200), .ZN(n5205) );
  NOR2_X1 U6339 ( .A1(n5202), .A2(n5201), .ZN(n6042) );
  NOR2_X1 U6340 ( .A1(n6042), .A2(n5203), .ZN(n5204) );
  AOI211_X1 U6341 ( .C1(n6048), .C2(EBX_REG_2__SCAN_IN), .A(n5205), .B(n5204), 
        .ZN(n5206) );
  OAI21_X1 U6342 ( .B1(n5859), .B2(n6051), .A(n5206), .ZN(n5208) );
  NOR2_X1 U6343 ( .A1(n6041), .A2(n6169), .ZN(n5207) );
  AOI211_X1 U6344 ( .C1(n6047), .C2(n6238), .A(n5208), .B(n5207), .ZN(n5209)
         );
  OAI21_X1 U6345 ( .B1(n6053), .B2(n6072), .A(n5209), .ZN(U2825) );
  NAND2_X1 U6346 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6014), .ZN(n5283) );
  MUX2_X1 U6347 ( .A(n5283), .B(REIP_REG_9__SCAN_IN), .S(REIP_REG_10__SCAN_IN), 
        .Z(n5213) );
  OAI22_X1 U6348 ( .A1(n3642), .A2(n6029), .B1(n5988), .B2(n5210), .ZN(n5211)
         );
  AOI211_X1 U6349 ( .C1(n6046), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5211), 
        .B(n6020), .ZN(n5212) );
  OAI21_X1 U6350 ( .B1(n6016), .B2(n5213), .A(n5212), .ZN(n5215) );
  NOR2_X1 U6351 ( .A1(n6041), .A2(n5265), .ZN(n5214) );
  AOI211_X1 U6352 ( .C1(REIP_REG_10__SCAN_IN), .C2(n6021), .A(n5215), .B(n5214), .ZN(n5216) );
  OAI21_X1 U6353 ( .B1(n5217), .B2(n6024), .A(n5216), .ZN(U2817) );
  AND2_X1 U6354 ( .A1(n5138), .A2(n5218), .ZN(n5220) );
  OR2_X1 U6355 ( .A1(n5220), .A2(n5219), .ZN(n6140) );
  AOI22_X1 U6356 ( .A1(n5357), .A2(DATAI_11_), .B1(n6084), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5221) );
  OAI21_X1 U6357 ( .B1(n6140), .B2(n5911), .A(n5221), .ZN(U2880) );
  AOI21_X1 U6358 ( .B1(n5222), .B2(n2984), .A(n5286), .ZN(n6178) );
  AOI22_X1 U6359 ( .A1(n4255), .A2(n6178), .B1(EBX_REG_11__SCAN_IN), .B2(n5544), .ZN(n5223) );
  OAI21_X1 U6360 ( .B1(n6140), .B2(n5579), .A(n5223), .ZN(U2848) );
  NOR2_X1 U6361 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5224), .ZN(n5253)
         );
  OAI21_X1 U6362 ( .B1(n5256), .B2(n5255), .A(n5225), .ZN(n5226) );
  NAND2_X1 U6363 ( .A1(n5226), .A2(n5231), .ZN(n5228) );
  OAI221_X1 U6364 ( .B1(n5253), .B2(n6508), .C1(n5253), .C2(n5228), .A(n5227), 
        .ZN(n5229) );
  INV_X1 U6365 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5234) );
  NAND3_X1 U6366 ( .A1(n6259), .A2(n6253), .A3(n6263), .ZN(n5230) );
  OAI21_X1 U6367 ( .B1(n5231), .B2(n6297), .A(n5230), .ZN(n5254) );
  AOI22_X1 U6368 ( .A1(n6270), .A2(n5254), .B1(n6321), .B2(n5253), .ZN(n5233)
         );
  AOI22_X1 U6369 ( .A1(n6320), .A2(n5256), .B1(n5255), .B2(n6322), .ZN(n5232)
         );
  OAI211_X1 U6370 ( .C1(n5260), .C2(n5234), .A(n5233), .B(n5232), .ZN(U3038)
         );
  INV_X1 U6371 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5237) );
  AOI22_X1 U6372 ( .A1(n6290), .A2(n5254), .B1(n6349), .B2(n5253), .ZN(n5236)
         );
  AOI22_X1 U6373 ( .A1(n6347), .A2(n5256), .B1(n5255), .B2(n6351), .ZN(n5235)
         );
  OAI211_X1 U6374 ( .C1(n5260), .C2(n5237), .A(n5236), .B(n5235), .ZN(U3043)
         );
  INV_X1 U6375 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5240) );
  AOI22_X1 U6376 ( .A1(n6284), .A2(n5254), .B1(n6341), .B2(n5253), .ZN(n5239)
         );
  AOI22_X1 U6377 ( .A1(n6340), .A2(n5256), .B1(n5255), .B2(n6342), .ZN(n5238)
         );
  OAI211_X1 U6378 ( .C1(n5260), .C2(n5240), .A(n5239), .B(n5238), .ZN(U3042)
         );
  INV_X1 U6379 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5243) );
  AOI22_X1 U6380 ( .A1(n6359), .A2(n5254), .B1(n6358), .B2(n5253), .ZN(n5242)
         );
  AOI22_X1 U6381 ( .A1(n6316), .A2(n5256), .B1(n5255), .B2(n6357), .ZN(n5241)
         );
  OAI211_X1 U6382 ( .C1(n5260), .C2(n5243), .A(n5242), .B(n5241), .ZN(U3037)
         );
  INV_X1 U6383 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5246) );
  AOI22_X1 U6384 ( .A1(n6277), .A2(n5254), .B1(n6331), .B2(n5253), .ZN(n5245)
         );
  AOI22_X1 U6385 ( .A1(n6330), .A2(n5256), .B1(n5255), .B2(n6332), .ZN(n5244)
         );
  OAI211_X1 U6386 ( .C1(n5260), .C2(n5246), .A(n5245), .B(n5244), .ZN(U3040)
         );
  INV_X1 U6387 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5249) );
  AOI22_X1 U6388 ( .A1(n6365), .A2(n5254), .B1(n6364), .B2(n5253), .ZN(n5248)
         );
  AOI22_X1 U6389 ( .A1(n6326), .A2(n5256), .B1(n5255), .B2(n6363), .ZN(n5247)
         );
  OAI211_X1 U6390 ( .C1(n5260), .C2(n5249), .A(n5248), .B(n5247), .ZN(U3039)
         );
  INV_X1 U6391 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5252) );
  AOI22_X1 U6392 ( .A1(n6256), .A2(n5254), .B1(n6304), .B2(n5253), .ZN(n5251)
         );
  AOI22_X1 U6393 ( .A1(n6312), .A2(n5256), .B1(n5255), .B2(n6303), .ZN(n5250)
         );
  OAI211_X1 U6394 ( .C1(n5260), .C2(n5252), .A(n5251), .B(n5250), .ZN(U3036)
         );
  INV_X1 U6395 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5259) );
  AOI22_X1 U6396 ( .A1(n6374), .A2(n5254), .B1(n6372), .B2(n5253), .ZN(n5258)
         );
  AOI22_X1 U6397 ( .A1(n6336), .A2(n5256), .B1(n5255), .B2(n6370), .ZN(n5257)
         );
  OAI211_X1 U6398 ( .C1(n5260), .C2(n5259), .A(n5258), .B(n5257), .ZN(U3041)
         );
  NAND2_X1 U6399 ( .A1(n6134), .A2(n5261), .ZN(n5263) );
  XOR2_X1 U6400 ( .A(n5263), .B(n5262), .Z(n5281) );
  NAND2_X1 U6401 ( .A1(n6240), .A2(REIP_REG_10__SCAN_IN), .ZN(n5276) );
  NAND2_X1 U6402 ( .A1(n6161), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5264)
         );
  OAI211_X1 U6403 ( .C1(n6170), .C2(n5265), .A(n5276), .B(n5264), .ZN(n5266)
         );
  AOI21_X1 U6404 ( .B1(n5267), .B2(n5681), .A(n5266), .ZN(n5268) );
  OAI21_X1 U6405 ( .B1(n5281), .B2(n6144), .A(n5268), .ZN(U2976) );
  INV_X1 U6406 ( .A(n5269), .ZN(n5272) );
  AOI22_X1 U6407 ( .A1(n6234), .A2(n5272), .B1(n5831), .B2(n5270), .ZN(n6210)
         );
  AOI21_X1 U6408 ( .B1(n6195), .B2(n5271), .A(n6210), .ZN(n6194) );
  NAND2_X1 U6409 ( .A1(n5272), .A2(n6230), .ZN(n6213) );
  NOR2_X1 U6410 ( .A1(n6195), .A2(n6213), .ZN(n6189) );
  NAND2_X1 U6411 ( .A1(n6189), .A2(n5273), .ZN(n5274) );
  OAI21_X1 U6412 ( .B1(n6194), .B2(n3494), .A(n5274), .ZN(n5275) );
  OAI21_X1 U6413 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A(n5275), .ZN(n5280) );
  INV_X1 U6414 ( .A(n5276), .ZN(n5277) );
  AOI21_X1 U6415 ( .B1(n6237), .B2(n5278), .A(n5277), .ZN(n5279) );
  OAI211_X1 U6416 ( .C1(n5281), .C2(n6184), .A(n5280), .B(n5279), .ZN(U3008)
         );
  XOR2_X1 U6417 ( .A(n5282), .B(n5219), .Z(n5305) );
  INV_X1 U6418 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5285) );
  INV_X1 U6419 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6465) );
  NOR2_X1 U6420 ( .A1(n6465), .A2(n5283), .ZN(n6001) );
  NAND2_X1 U6421 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6001), .ZN(n5316) );
  INV_X1 U6422 ( .A(n5316), .ZN(n5289) );
  OAI21_X1 U6423 ( .B1(n6016), .B2(n5289), .A(n5378), .ZN(n6003) );
  AOI22_X1 U6424 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6048), .B1(
        REIP_REG_12__SCAN_IN), .B2(n6003), .ZN(n5284) );
  OAI211_X1 U6425 ( .C1(n6035), .C2(n5285), .A(n5284), .B(n6033), .ZN(n5292)
         );
  NOR2_X1 U6426 ( .A1(n6016), .A2(REIP_REG_12__SCAN_IN), .ZN(n5995) );
  OR2_X1 U6427 ( .A1(n5287), .A2(n5286), .ZN(n5288) );
  AND2_X1 U6428 ( .A1(n5288), .A2(n2971), .ZN(n6171) );
  AOI22_X1 U6429 ( .A1(n5995), .A2(n5289), .B1(n6047), .B2(n6171), .ZN(n5290)
         );
  OAI21_X1 U6430 ( .B1(n6041), .B2(n5303), .A(n5290), .ZN(n5291) );
  AOI211_X1 U6431 ( .C1(n5305), .C2(n6038), .A(n5292), .B(n5291), .ZN(n5293)
         );
  INV_X1 U6432 ( .A(n5293), .ZN(U2815) );
  INV_X1 U6433 ( .A(n5305), .ZN(n5295) );
  AOI22_X1 U6434 ( .A1(n5357), .A2(DATAI_12_), .B1(n6084), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5294) );
  OAI21_X1 U6435 ( .B1(n5295), .B2(n5911), .A(n5294), .ZN(U2879) );
  INV_X1 U6436 ( .A(n6171), .ZN(n5296) );
  OAI222_X1 U6437 ( .A1(n5578), .A2(n5296), .B1(n6076), .B2(n3648), .C1(n5579), 
        .C2(n5295), .ZN(U2847) );
  INV_X1 U6438 ( .A(n5297), .ZN(n5299) );
  NAND2_X1 U6439 ( .A1(n5299), .A2(n5298), .ZN(n5300) );
  XNOR2_X1 U6440 ( .A(n5301), .B(n5300), .ZN(n6172) );
  INV_X1 U6441 ( .A(n6172), .ZN(n5307) );
  AOI22_X1 U6442 ( .A1(n6161), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n6240), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n5302) );
  OAI21_X1 U6443 ( .B1(n5303), .B2(n6170), .A(n5302), .ZN(n5304) );
  AOI21_X1 U6444 ( .B1(n5305), .B2(n5681), .A(n5304), .ZN(n5306) );
  OAI21_X1 U6445 ( .B1(n5307), .B2(n6144), .A(n5306), .ZN(U2974) );
  NAND2_X1 U6446 ( .A1(n5310), .A2(n5309), .ZN(n5311) );
  AOI22_X1 U6447 ( .A1(n5357), .A2(DATAI_13_), .B1(n6084), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5312) );
  OAI21_X1 U6448 ( .B1(n5331), .B2(n5911), .A(n5312), .ZN(U2878) );
  NAND2_X1 U6449 ( .A1(n5308), .A2(n5313), .ZN(n5315) );
  NAND2_X1 U6450 ( .A1(n5315), .A2(n5314), .ZN(n5354) );
  OAI21_X1 U6451 ( .B1(n5315), .B2(n5314), .A(n5354), .ZN(n5731) );
  INV_X1 U6452 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6471) );
  INV_X1 U6453 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6468) );
  NOR2_X1 U6454 ( .A1(n6468), .A2(n5316), .ZN(n5990) );
  NAND2_X1 U6455 ( .A1(REIP_REG_13__SCAN_IN), .A2(n5990), .ZN(n5321) );
  NOR2_X1 U6456 ( .A1(n6471), .A2(n5321), .ZN(n5371) );
  INV_X1 U6457 ( .A(n5371), .ZN(n5520) );
  NAND2_X1 U6458 ( .A1(n6002), .A2(n5520), .ZN(n5322) );
  NAND2_X1 U6459 ( .A1(n5322), .A2(n5378), .ZN(n5976) );
  INV_X1 U6460 ( .A(n5976), .ZN(n5326) );
  OR2_X1 U6461 ( .A1(n5318), .A2(n5317), .ZN(n5319) );
  NAND2_X1 U6462 ( .A1(n5319), .A2(n5835), .ZN(n5844) );
  NAND2_X1 U6463 ( .A1(n6046), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5320)
         );
  OAI211_X1 U6464 ( .C1(n5988), .C2(n5844), .A(n6033), .B(n5320), .ZN(n5324)
         );
  NOR2_X1 U6465 ( .A1(n5322), .A2(n5321), .ZN(n5323) );
  AOI211_X1 U6466 ( .C1(EBX_REG_14__SCAN_IN), .C2(n6048), .A(n5324), .B(n5323), 
        .ZN(n5325) );
  OAI21_X1 U6467 ( .B1(n6471), .B2(n5326), .A(n5325), .ZN(n5327) );
  AOI21_X1 U6468 ( .B1(n6057), .B2(n5727), .A(n5327), .ZN(n5328) );
  OAI21_X1 U6469 ( .B1(n5731), .B2(n6024), .A(n5328), .ZN(U2813) );
  AOI22_X1 U6470 ( .A1(n5357), .A2(DATAI_14_), .B1(n6084), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5329) );
  OAI21_X1 U6471 ( .B1(n5731), .B2(n5911), .A(n5329), .ZN(U2877) );
  XNOR2_X1 U6472 ( .A(n5330), .B(n2971), .ZN(n5987) );
  OAI222_X1 U6473 ( .A1(n5579), .A2(n5331), .B1(n6076), .B2(n3652), .C1(n5578), 
        .C2(n5987), .ZN(U2846) );
  INV_X1 U6474 ( .A(n5332), .ZN(n5800) );
  AOI22_X1 U6475 ( .A1(n5800), .A2(n5345), .B1(n5334), .B2(n5333), .ZN(n6180)
         );
  NAND2_X1 U6476 ( .A1(n6173), .A2(n5335), .ZN(n5336) );
  OAI211_X1 U6477 ( .C1(n5843), .C2(n5346), .A(n6180), .B(n5336), .ZN(n5846)
         );
  INV_X1 U6478 ( .A(n5846), .ZN(n5352) );
  XNOR2_X1 U6479 ( .A(n5337), .B(n5338), .ZN(n5925) );
  NAND2_X1 U6480 ( .A1(n5925), .A2(n6242), .ZN(n5351) );
  AND2_X1 U6481 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5339), .ZN(n6235)
         );
  AOI21_X1 U6482 ( .B1(n5341), .B2(n6235), .A(n5340), .ZN(n5344) );
  INV_X1 U6483 ( .A(n5342), .ZN(n5343) );
  NOR4_X1 U6484 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5344), .A3(n5343), 
        .A4(n6173), .ZN(n5847) );
  NOR4_X1 U6485 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5346), .A3(n6173), 
        .A4(n5345), .ZN(n5349) );
  INV_X1 U6486 ( .A(REIP_REG_13__SCAN_IN), .ZN(n5347) );
  OAI22_X1 U6487 ( .A1(n6198), .A2(n5987), .B1(n6196), .B2(n5347), .ZN(n5348)
         );
  NOR3_X1 U6488 ( .A1(n5847), .A2(n5349), .A3(n5348), .ZN(n5350) );
  OAI211_X1 U6489 ( .C1(n5352), .C2(n3726), .A(n5351), .B(n5350), .ZN(U3005)
         );
  AND2_X1 U6490 ( .A1(n5354), .A2(n5353), .ZN(n5356) );
  OR2_X1 U6491 ( .A1(n5356), .A2(n5355), .ZN(n5980) );
  AOI22_X1 U6492 ( .A1(n5357), .A2(DATAI_15_), .B1(n6084), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5358) );
  OAI21_X1 U6493 ( .B1(n5980), .B2(n5911), .A(n5358), .ZN(U2876) );
  AOI22_X1 U6494 ( .A1(n5361), .A2(n5360), .B1(n5359), .B2(n5367), .ZN(n6391)
         );
  OAI21_X1 U6495 ( .B1(n6391), .B2(STATE2_REG_3__SCAN_IN), .A(n5362), .ZN(
        n5365) );
  AOI22_X1 U6496 ( .A1(n5365), .A2(n5364), .B1(n5363), .B2(n5367), .ZN(n5370)
         );
  AOI21_X1 U6497 ( .B1(n6389), .B2(n5366), .A(n5369), .ZN(n5368) );
  OAI22_X1 U6498 ( .A1(n5370), .A2(n5369), .B1(n5368), .B2(n5367), .ZN(U3461)
         );
  NAND3_X1 U6499 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .A3(
        n5371), .ZN(n5377) );
  NOR2_X1 U6500 ( .A1(n6016), .A2(n5377), .ZN(n5510) );
  NAND2_X1 U6501 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5510), .ZN(n5969) );
  NAND2_X1 U6502 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5497) );
  NOR2_X1 U6503 ( .A1(n5969), .A2(n5497), .ZN(n5906) );
  NAND2_X1 U6504 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5906), .ZN(n5889) );
  NAND3_X1 U6505 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5372) );
  NAND3_X1 U6506 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5445) );
  INV_X1 U6507 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6489) );
  NOR2_X1 U6508 ( .A1(n5445), .A2(n6489), .ZN(n5373) );
  NAND2_X1 U6509 ( .A1(n5878), .A2(n5373), .ZN(n5435) );
  INV_X1 U6510 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6491) );
  OR3_X1 U6511 ( .A1(n5435), .A2(n5418), .A3(n6491), .ZN(n5411) );
  NOR3_X1 U6512 ( .A1(n5411), .A2(REIP_REG_31__SCAN_IN), .A3(n6498), .ZN(n5387) );
  NOR3_X1 U6513 ( .A1(n5375), .A2(n5528), .A3(n5374), .ZN(n5376) );
  AOI21_X1 U6514 ( .B1(n6046), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5376), 
        .ZN(n5386) );
  INV_X1 U6515 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6479) );
  INV_X1 U6516 ( .A(n5377), .ZN(n5379) );
  NAND3_X1 U6517 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5379), .A3(n5378), .ZN(
        n5498) );
  NOR3_X1 U6518 ( .A1(n6479), .A2(n5497), .A3(n5498), .ZN(n5887) );
  INV_X1 U6519 ( .A(n5445), .ZN(n5380) );
  AND3_X1 U6520 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5467) );
  NAND3_X1 U6521 ( .A1(n5887), .A2(n5380), .A3(n5467), .ZN(n5381) );
  NAND2_X1 U6522 ( .A1(n5381), .A2(n5499), .ZN(n5439) );
  AND2_X1 U6523 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5439), .ZN(n5382) );
  NAND2_X1 U6524 ( .A1(REIP_REG_28__SCAN_IN), .A2(n5382), .ZN(n5383) );
  NAND2_X1 U6525 ( .A1(n5499), .A2(n5383), .ZN(n5429) );
  OAI21_X1 U6526 ( .B1(REIP_REG_29__SCAN_IN), .B2(n6016), .A(n5429), .ZN(n5407) );
  NOR2_X1 U6527 ( .A1(n6016), .A2(REIP_REG_30__SCAN_IN), .ZN(n5384) );
  OAI21_X1 U6528 ( .B1(n5407), .B2(n5384), .A(REIP_REG_31__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U6529 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(n5389), .ZN(n5391) );
  NAND3_X1 U6530 ( .A1(n5391), .A2(n5390), .A3(n5947), .ZN(U2788) );
  NAND2_X1 U6531 ( .A1(n5392), .A2(n5401), .ZN(n5400) );
  NAND3_X1 U6532 ( .A1(n5394), .A2(n5393), .A3(n4331), .ZN(n5398) );
  INV_X1 U6533 ( .A(n5401), .ZN(n5397) );
  AOI22_X1 U6534 ( .A1(n5398), .A2(n5397), .B1(n5396), .B2(n5395), .ZN(n5399)
         );
  AND2_X1 U6535 ( .A1(n5400), .A2(n5399), .ZN(n6381) );
  INV_X1 U6536 ( .A(n6381), .ZN(n5406) );
  OAI22_X1 U6537 ( .A1(n5404), .A2(n5403), .B1(n5402), .B2(n5401), .ZN(n5945)
         );
  AOI21_X1 U6538 ( .B1(n5405), .B2(n6440), .A(READY_N), .ZN(n6522) );
  OR2_X1 U6539 ( .A1(n5945), .A2(n6522), .ZN(n6382) );
  AND2_X1 U6540 ( .A1(n6382), .A2(n6422), .ZN(n5951) );
  MUX2_X1 U6541 ( .A(MORE_REG_SCAN_IN), .B(n5406), .S(n5951), .Z(U3471) );
  INV_X1 U6542 ( .A(n5608), .ZN(n5584) );
  INV_X1 U6543 ( .A(n5606), .ZN(n5414) );
  AOI22_X1 U6544 ( .A1(n6048), .A2(EBX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6046), .ZN(n5409) );
  NAND2_X1 U6545 ( .A1(n5407), .A2(REIP_REG_30__SCAN_IN), .ZN(n5408) );
  OAI211_X1 U6546 ( .C1(n5410), .C2(n5988), .A(n5409), .B(n5408), .ZN(n5413)
         );
  NOR2_X1 U6547 ( .A1(n5411), .A2(REIP_REG_30__SCAN_IN), .ZN(n5412) );
  AOI211_X1 U6548 ( .C1(n5414), .C2(n6057), .A(n5413), .B(n5412), .ZN(n5415)
         );
  OAI21_X1 U6549 ( .B1(n5584), .B2(n6024), .A(n5415), .ZN(U2797) );
  NAND2_X1 U6550 ( .A1(n5530), .A2(n6047), .ZN(n5417) );
  AOI22_X1 U6551 ( .A1(n6048), .A2(EBX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6046), .ZN(n5416) );
  OAI211_X1 U6552 ( .C1(n5429), .C2(n5418), .A(n5417), .B(n5416), .ZN(n5419)
         );
  AOI21_X1 U6553 ( .B1(n6057), .B2(n5420), .A(n5419), .ZN(n5422) );
  OR3_X1 U6554 ( .A1(n5435), .A2(REIP_REG_29__SCAN_IN), .A3(n6491), .ZN(n5421)
         );
  OAI211_X1 U6555 ( .C1(n5587), .C2(n6024), .A(n5422), .B(n5421), .ZN(U2798)
         );
  AOI21_X1 U6556 ( .B1(n5424), .B2(n5437), .A(n4307), .ZN(n5620) );
  NAND2_X1 U6557 ( .A1(n5620), .A2(n6038), .ZN(n5434) );
  INV_X1 U6558 ( .A(n5618), .ZN(n5432) );
  AND2_X1 U6559 ( .A1(n5442), .A2(n5425), .ZN(n5427) );
  NOR2_X1 U6560 ( .A1(n5732), .A2(n5988), .ZN(n5431) );
  AOI22_X1 U6561 ( .A1(n6048), .A2(EBX_REG_28__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6046), .ZN(n5428) );
  OAI21_X1 U6562 ( .B1(n5429), .B2(n6491), .A(n5428), .ZN(n5430) );
  AOI211_X1 U6563 ( .C1(n6057), .C2(n5432), .A(n5431), .B(n5430), .ZN(n5433)
         );
  OAI211_X1 U6564 ( .C1(REIP_REG_28__SCAN_IN), .C2(n5435), .A(n5434), .B(n5433), .ZN(U2799) );
  INV_X1 U6565 ( .A(n5439), .ZN(n5459) );
  NAND2_X1 U6566 ( .A1(n5455), .A2(n5440), .ZN(n5441) );
  NAND2_X1 U6567 ( .A1(n5442), .A2(n5441), .ZN(n5742) );
  NAND2_X1 U6568 ( .A1(n6057), .A2(n5629), .ZN(n5444) );
  AOI22_X1 U6569 ( .A1(n6048), .A2(EBX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6046), .ZN(n5443) );
  OAI211_X1 U6570 ( .C1(n5988), .C2(n5742), .A(n5444), .B(n5443), .ZN(n5447)
         );
  INV_X1 U6571 ( .A(n5878), .ZN(n5452) );
  NOR3_X1 U6572 ( .A1(n5452), .A2(REIP_REG_27__SCAN_IN), .A3(n5445), .ZN(n5446) );
  AOI211_X1 U6573 ( .C1(REIP_REG_27__SCAN_IN), .C2(n5459), .A(n5447), .B(n5446), .ZN(n5448) );
  OAI21_X1 U6574 ( .B1(n5626), .B2(n6024), .A(n5448), .ZN(U2800) );
  AOI21_X1 U6575 ( .B1(n5450), .B2(n5449), .A(n5436), .ZN(n5635) );
  INV_X1 U6576 ( .A(n5635), .ZN(n5595) );
  NAND2_X1 U6577 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5471) );
  INV_X1 U6578 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5451) );
  OAI21_X1 U6579 ( .B1(n5452), .B2(n5471), .A(n5451), .ZN(n5460) );
  NOR2_X1 U6580 ( .A1(n6041), .A2(n5633), .ZN(n5458) );
  NAND2_X1 U6581 ( .A1(n5464), .A2(n5453), .ZN(n5454) );
  NAND2_X1 U6582 ( .A1(n5455), .A2(n5454), .ZN(n5750) );
  AOI22_X1 U6583 ( .A1(n6048), .A2(EBX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6046), .ZN(n5456) );
  OAI21_X1 U6584 ( .B1(n5750), .B2(n5988), .A(n5456), .ZN(n5457) );
  AOI211_X1 U6585 ( .C1(n5460), .C2(n5459), .A(n5458), .B(n5457), .ZN(n5461)
         );
  OAI21_X1 U6586 ( .B1(n5595), .B2(n6024), .A(n5461), .ZN(U2801) );
  OAI21_X1 U6587 ( .B1(n5462), .B2(n5463), .A(n5449), .ZN(n5644) );
  OAI21_X1 U6588 ( .B1(n5540), .B2(n5465), .A(n5464), .ZN(n5761) );
  AOI22_X1 U6589 ( .A1(n6048), .A2(EBX_REG_25__SCAN_IN), .B1(n6046), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5466) );
  OAI21_X1 U6590 ( .B1(n5761), .B2(n5988), .A(n5466), .ZN(n5470) );
  NAND2_X1 U6591 ( .A1(n5887), .A2(n5467), .ZN(n5468) );
  NAND2_X1 U6592 ( .A1(n5468), .A2(n5499), .ZN(n5870) );
  INV_X1 U6593 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6571) );
  NOR2_X1 U6594 ( .A1(n5870), .A2(n6571), .ZN(n5469) );
  AOI211_X1 U6595 ( .C1(n6057), .C2(n5639), .A(n5470), .B(n5469), .ZN(n5473)
         );
  OAI211_X1 U6596 ( .C1(REIP_REG_24__SCAN_IN), .C2(REIP_REG_25__SCAN_IN), .A(
        n5878), .B(n5471), .ZN(n5472) );
  OAI211_X1 U6597 ( .C1(n5644), .C2(n6024), .A(n5473), .B(n5472), .ZN(U2802)
         );
  INV_X1 U6598 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6481) );
  NOR2_X1 U6599 ( .A1(n6481), .A2(n5889), .ZN(n5883) );
  AOI21_X1 U6600 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5883), .A(
        REIP_REG_23__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U6601 ( .A1(n5475), .A2(n5476), .ZN(n5477) );
  NAND2_X1 U6602 ( .A1(n5474), .A2(n5477), .ZN(n5659) );
  INV_X1 U6603 ( .A(n5659), .ZN(n5478) );
  NAND2_X1 U6604 ( .A1(n5478), .A2(n6038), .ZN(n5485) );
  INV_X1 U6605 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5479) );
  OAI22_X1 U6606 ( .A1(n5479), .A2(n6029), .B1(n5658), .B2(n6035), .ZN(n5483)
         );
  AOI21_X1 U6607 ( .B1(n5480), .B2(n5551), .A(n5539), .ZN(n5773) );
  INV_X1 U6608 ( .A(n5773), .ZN(n5481) );
  NOR2_X1 U6609 ( .A1(n5481), .A2(n5988), .ZN(n5482) );
  AOI211_X1 U6610 ( .C1(n6057), .C2(n5662), .A(n5483), .B(n5482), .ZN(n5484)
         );
  OAI211_X1 U6611 ( .C1(n5486), .C2(n5870), .A(n5485), .B(n5484), .ZN(U2804)
         );
  INV_X1 U6612 ( .A(n5488), .ZN(n5489) );
  INV_X1 U6613 ( .A(n5490), .ZN(n5562) );
  NOR2_X1 U6614 ( .A1(n3617), .A2(n5491), .ZN(n5492) );
  AOI21_X1 U6615 ( .B1(n5562), .B2(n3617), .A(n5492), .ZN(n5569) );
  OR2_X1 U6616 ( .A1(n5569), .A2(n5493), .ZN(n5571) );
  XNOR2_X1 U6617 ( .A(n5571), .B(n2985), .ZN(n5818) );
  OAI21_X1 U6618 ( .B1(n6035), .B2(n5685), .A(n6033), .ZN(n5494) );
  AOI21_X1 U6619 ( .B1(n6047), .B2(n5818), .A(n5494), .ZN(n5495) );
  OAI21_X1 U6620 ( .B1(n5496), .B2(n6029), .A(n5495), .ZN(n5502) );
  OAI21_X1 U6621 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n5497), .ZN(n5500) );
  INV_X1 U6622 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6574) );
  NAND2_X1 U6623 ( .A1(n5499), .A2(n5498), .ZN(n5968) );
  OAI22_X1 U6624 ( .A1(n5969), .A2(n5500), .B1(n6574), .B2(n5968), .ZN(n5501)
         );
  AOI211_X1 U6625 ( .C1(n6057), .C2(n5687), .A(n5502), .B(n5501), .ZN(n5503)
         );
  OAI21_X1 U6626 ( .B1(n5921), .B2(n6024), .A(n5503), .ZN(U2808) );
  INV_X1 U6627 ( .A(n5504), .ZN(n5506) );
  OAI21_X1 U6628 ( .B1(n5506), .B2(n3070), .A(n5567), .ZN(n5708) );
  OR2_X1 U6629 ( .A1(n5518), .A2(n5507), .ZN(n5508) );
  AND2_X1 U6630 ( .A1(n5493), .A2(n5508), .ZN(n5929) );
  INV_X1 U6631 ( .A(n5929), .ZN(n5574) );
  NAND2_X1 U6632 ( .A1(n6048), .A2(EBX_REG_17__SCAN_IN), .ZN(n5509) );
  OAI211_X1 U6633 ( .C1(n5574), .C2(n5988), .A(n5509), .B(n6033), .ZN(n5513)
         );
  NOR2_X1 U6634 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5510), .ZN(n5511) );
  OAI22_X1 U6635 ( .A1(n5511), .A2(n5968), .B1(n5703), .B2(n6035), .ZN(n5512)
         );
  AOI211_X1 U6636 ( .C1(n6057), .C2(n5705), .A(n5513), .B(n5512), .ZN(n5514)
         );
  OAI21_X1 U6637 ( .B1(n5708), .B2(n6024), .A(n5514), .ZN(U2810) );
  OAI21_X1 U6638 ( .B1(n5355), .B2(n5515), .A(n5504), .ZN(n6080) );
  NOR2_X1 U6639 ( .A1(n5516), .A2(n5834), .ZN(n5517) );
  OR2_X1 U6640 ( .A1(n5518), .A2(n5517), .ZN(n5936) );
  AOI21_X1 U6641 ( .B1(n6046), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6020), 
        .ZN(n5519) );
  OAI21_X1 U6642 ( .B1(n5988), .B2(n5936), .A(n5519), .ZN(n5526) );
  INV_X1 U6643 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5577) );
  NOR2_X1 U6644 ( .A1(n6016), .A2(n5520), .ZN(n5522) );
  INV_X1 U6645 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5521) );
  AND2_X1 U6646 ( .A1(n5522), .A2(n5521), .ZN(n5977) );
  OAI21_X1 U6647 ( .B1(n5976), .B2(n5977), .A(REIP_REG_16__SCAN_IN), .ZN(n5524) );
  INV_X1 U6648 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6474) );
  NAND3_X1 U6649 ( .A1(n5522), .A2(REIP_REG_15__SCAN_IN), .A3(n6474), .ZN(
        n5523) );
  OAI211_X1 U6650 ( .C1(n6029), .C2(n5577), .A(n5524), .B(n5523), .ZN(n5525)
         );
  AOI211_X1 U6651 ( .C1(n5715), .C2(n6057), .A(n5526), .B(n5525), .ZN(n5527)
         );
  OAI21_X1 U6652 ( .B1(n6080), .B2(n6024), .A(n5527), .ZN(U2811) );
  OAI22_X1 U6653 ( .A1(n5529), .A2(n5578), .B1(n6076), .B2(n5528), .ZN(U2828)
         );
  AOI22_X1 U6654 ( .A1(n5530), .A2(n4255), .B1(EBX_REG_29__SCAN_IN), .B2(n5544), .ZN(n5531) );
  OAI21_X1 U6655 ( .B1(n5587), .B2(n5579), .A(n5531), .ZN(U2830) );
  INV_X1 U6656 ( .A(n5620), .ZN(n5590) );
  OAI222_X1 U6657 ( .A1(n5579), .A2(n5590), .B1(n5532), .B2(n6076), .C1(n5732), 
        .C2(n5578), .ZN(U2831) );
  INV_X1 U6658 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5533) );
  OAI222_X1 U6659 ( .A1(n5579), .A2(n5626), .B1(n5533), .B2(n6076), .C1(n5742), 
        .C2(n5578), .ZN(U2832) );
  OAI222_X1 U6660 ( .A1(n5579), .A2(n5595), .B1(n5534), .B2(n6076), .C1(n5750), 
        .C2(n5578), .ZN(U2833) );
  INV_X1 U6661 ( .A(n5761), .ZN(n5535) );
  AOI22_X1 U6662 ( .A1(n5535), .A2(n4255), .B1(EBX_REG_25__SCAN_IN), .B2(n5544), .ZN(n5536) );
  OAI21_X1 U6663 ( .B1(n5644), .B2(n5579), .A(n5536), .ZN(U2834) );
  AOI21_X1 U6664 ( .B1(n5537), .B2(n5474), .A(n5462), .ZN(n5652) );
  INV_X1 U6665 ( .A(n5652), .ZN(n5875) );
  INV_X1 U6666 ( .A(n5538), .ZN(n5542) );
  INV_X1 U6667 ( .A(n5539), .ZN(n5541) );
  AOI21_X1 U6668 ( .B1(n5542), .B2(n5541), .A(n5540), .ZN(n5873) );
  AOI22_X1 U6669 ( .A1(n5873), .A2(n4255), .B1(EBX_REG_24__SCAN_IN), .B2(n5544), .ZN(n5543) );
  OAI21_X1 U6670 ( .B1(n5875), .B2(n5579), .A(n5543), .ZN(U2835) );
  AOI22_X1 U6671 ( .A1(n5773), .A2(n4255), .B1(EBX_REG_23__SCAN_IN), .B2(n5544), .ZN(n5545) );
  OAI21_X1 U6672 ( .B1(n5659), .B2(n5579), .A(n5545), .ZN(U2836) );
  INV_X1 U6673 ( .A(n5475), .ZN(n5546) );
  AOI21_X1 U6674 ( .B1(n5547), .B2(n2965), .A(n5546), .ZN(n5912) );
  INV_X1 U6675 ( .A(n5912), .ZN(n5553) );
  NAND2_X1 U6676 ( .A1(n5548), .A2(n5549), .ZN(n5550) );
  NAND2_X1 U6677 ( .A1(n5551), .A2(n5550), .ZN(n5885) );
  OAI222_X1 U6678 ( .A1(n5579), .A2(n5553), .B1(n5552), .B2(n6076), .C1(n5885), 
        .C2(n5578), .ZN(U2837) );
  OAI21_X1 U6679 ( .B1(n5554), .B2(n2972), .A(n2965), .ZN(n5895) );
  OR2_X1 U6680 ( .A1(n5556), .A2(n5555), .ZN(n5557) );
  NAND2_X1 U6681 ( .A1(n5548), .A2(n5557), .ZN(n5896) );
  OAI222_X1 U6682 ( .A1(n5579), .A2(n5895), .B1(n5558), .B2(n6076), .C1(n5896), 
        .C2(n5578), .ZN(U2838) );
  AOI21_X1 U6683 ( .B1(n5559), .B2(n2966), .A(n2972), .ZN(n5918) );
  INV_X1 U6684 ( .A(n5918), .ZN(n5904) );
  MUX2_X1 U6685 ( .A(n5562), .B(n5561), .S(n5560), .Z(n5564) );
  XNOR2_X1 U6686 ( .A(n5564), .B(n5563), .ZN(n5903) );
  OAI222_X1 U6687 ( .A1(n5579), .A2(n5904), .B1(n6076), .B2(n3671), .C1(n5903), 
        .C2(n5578), .ZN(U2839) );
  INV_X1 U6688 ( .A(n5818), .ZN(n5565) );
  OAI222_X1 U6689 ( .A1(n5921), .A2(n5579), .B1(n6076), .B2(n5496), .C1(n5578), 
        .C2(n5565), .ZN(U2840) );
  NAND2_X1 U6690 ( .A1(n5567), .A2(n5566), .ZN(n5568) );
  NAND2_X1 U6691 ( .A1(n5488), .A2(n5568), .ZN(n5971) );
  NAND2_X1 U6692 ( .A1(n5569), .A2(n5493), .ZN(n5570) );
  INV_X1 U6693 ( .A(n5972), .ZN(n5572) );
  OAI222_X1 U6694 ( .A1(n5579), .A2(n5971), .B1(n5573), .B2(n6076), .C1(n5572), 
        .C2(n5578), .ZN(U2841) );
  OAI22_X1 U6695 ( .A1(n5578), .A2(n5574), .B1(n6639), .B2(n6076), .ZN(n5575)
         );
  INV_X1 U6696 ( .A(n5575), .ZN(n5576) );
  OAI21_X1 U6697 ( .B1(n5708), .B2(n5579), .A(n5576), .ZN(U2842) );
  OAI222_X1 U6698 ( .A1(n6080), .A2(n5579), .B1(n6076), .B2(n5577), .C1(n5936), 
        .C2(n5578), .ZN(U2843) );
  OAI222_X1 U6699 ( .A1(n5731), .A2(n5579), .B1(n6076), .B2(n3655), .C1(n5844), 
        .C2(n5578), .ZN(U2845) );
  AOI22_X1 U6700 ( .A1(n6081), .A2(DATAI_30_), .B1(n6084), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U6701 ( .A1(n6085), .A2(DATAI_14_), .ZN(n5582) );
  OAI211_X1 U6702 ( .C1(n5584), .C2(n5911), .A(n5583), .B(n5582), .ZN(U2861)
         );
  AOI22_X1 U6703 ( .A1(n6081), .A2(DATAI_29_), .B1(n6084), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U6704 ( .A1(n6085), .A2(DATAI_13_), .ZN(n5585) );
  OAI211_X1 U6705 ( .C1(n5587), .C2(n5911), .A(n5586), .B(n5585), .ZN(U2862)
         );
  AOI22_X1 U6706 ( .A1(n6081), .A2(DATAI_28_), .B1(n6084), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U6707 ( .A1(n6085), .A2(DATAI_12_), .ZN(n5588) );
  OAI211_X1 U6708 ( .C1(n5590), .C2(n5911), .A(n5589), .B(n5588), .ZN(U2863)
         );
  AOI22_X1 U6709 ( .A1(n6081), .A2(DATAI_27_), .B1(n6084), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U6710 ( .A1(n6085), .A2(DATAI_11_), .ZN(n5591) );
  OAI211_X1 U6711 ( .C1(n5626), .C2(n5911), .A(n5592), .B(n5591), .ZN(U2864)
         );
  AOI22_X1 U6712 ( .A1(n6081), .A2(DATAI_26_), .B1(n6084), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U6713 ( .A1(n6085), .A2(DATAI_10_), .ZN(n5593) );
  OAI211_X1 U6714 ( .C1(n5595), .C2(n5911), .A(n5594), .B(n5593), .ZN(U2865)
         );
  AOI22_X1 U6715 ( .A1(n6081), .A2(DATAI_25_), .B1(n6084), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U6716 ( .A1(n6085), .A2(DATAI_9_), .ZN(n5596) );
  OAI211_X1 U6717 ( .C1(n5644), .C2(n5911), .A(n5597), .B(n5596), .ZN(U2866)
         );
  AOI22_X1 U6718 ( .A1(n6085), .A2(DATAI_8_), .B1(n6084), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U6719 ( .A1(n6081), .A2(DATAI_24_), .ZN(n5598) );
  OAI211_X1 U6720 ( .C1(n5875), .C2(n5911), .A(n5599), .B(n5598), .ZN(U2867)
         );
  AOI22_X1 U6721 ( .A1(n6081), .A2(DATAI_23_), .B1(n6084), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5601) );
  NAND2_X1 U6722 ( .A1(n6085), .A2(DATAI_7_), .ZN(n5600) );
  OAI211_X1 U6723 ( .C1(n5659), .C2(n5911), .A(n5601), .B(n5600), .ZN(U2868)
         );
  AOI22_X1 U6724 ( .A1(n6081), .A2(DATAI_17_), .B1(n6084), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U6725 ( .A1(n6085), .A2(DATAI_1_), .ZN(n5602) );
  OAI211_X1 U6726 ( .C1(n5708), .C2(n5911), .A(n5603), .B(n5602), .ZN(U2874)
         );
  AOI21_X1 U6727 ( .B1(n6161), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5604), 
        .ZN(n5605) );
  OAI21_X1 U6728 ( .B1(n5606), .B2(n6170), .A(n5605), .ZN(n5607) );
  OAI21_X1 U6729 ( .B1(n5610), .B2(n6144), .A(n5609), .ZN(U2956) );
  NAND3_X1 U6730 ( .A1(n5611), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5648), .ZN(n5615) );
  NAND2_X1 U6731 ( .A1(n5612), .A2(n5614), .ZN(n5753) );
  NOR2_X1 U6732 ( .A1(n5648), .A2(n5753), .ZN(n5613) );
  NAND2_X1 U6733 ( .A1(n5640), .A2(n5613), .ZN(n5622) );
  AOI22_X1 U6734 ( .A1(n5615), .A2(n5622), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5614), .ZN(n5616) );
  XNOR2_X1 U6735 ( .A(n5616), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5740)
         );
  NOR2_X1 U6736 ( .A1(n6196), .A2(n6491), .ZN(n5734) );
  AOI21_X1 U6737 ( .B1(n6161), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5734), 
        .ZN(n5617) );
  OAI21_X1 U6738 ( .B1(n5618), .B2(n6170), .A(n5617), .ZN(n5619) );
  AOI21_X1 U6739 ( .B1(n5620), .B2(n5681), .A(n5619), .ZN(n5621) );
  OAI21_X1 U6740 ( .B1(n6144), .B2(n5740), .A(n5621), .ZN(U2958) );
  NAND2_X1 U6741 ( .A1(n5623), .A2(n5622), .ZN(n5624) );
  XNOR2_X1 U6742 ( .A(n5624), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5748)
         );
  NAND2_X1 U6743 ( .A1(n6240), .A2(REIP_REG_27__SCAN_IN), .ZN(n5741) );
  OAI21_X1 U6744 ( .B1(n5725), .B2(n5625), .A(n5741), .ZN(n5628) );
  NOR2_X1 U6745 ( .A1(n5626), .A2(n6139), .ZN(n5627) );
  OAI21_X1 U6746 ( .B1(n5748), .B2(n6144), .A(n5630), .ZN(U2959) );
  XNOR2_X1 U6747 ( .A(n5648), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5631)
         );
  XNOR2_X1 U6748 ( .A(n5611), .B(n5631), .ZN(n5757) );
  NAND2_X1 U6749 ( .A1(n6240), .A2(REIP_REG_26__SCAN_IN), .ZN(n5749) );
  NAND2_X1 U6750 ( .A1(n6161), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5632)
         );
  OAI211_X1 U6751 ( .C1(n5633), .C2(n6170), .A(n5749), .B(n5632), .ZN(n5634)
         );
  AOI21_X1 U6752 ( .B1(n5635), .B2(n5681), .A(n5634), .ZN(n5636) );
  OAI21_X1 U6753 ( .B1(n6144), .B2(n5757), .A(n5636), .ZN(U2960) );
  NAND2_X1 U6754 ( .A1(n6240), .A2(REIP_REG_25__SCAN_IN), .ZN(n5760) );
  OAI21_X1 U6755 ( .B1(n5725), .B2(n5637), .A(n5760), .ZN(n5638) );
  AOI21_X1 U6756 ( .B1(n5639), .B2(n5728), .A(n5638), .ZN(n5643) );
  OAI21_X1 U6757 ( .B1(n5641), .B2(n5640), .A(n3513), .ZN(n5759) );
  NAND2_X1 U6758 ( .A1(n5759), .A2(n6165), .ZN(n5642) );
  OAI211_X1 U6759 ( .C1(n5644), .C2(n6139), .A(n5643), .B(n5642), .ZN(U2961)
         );
  XNOR2_X1 U6760 ( .A(n5648), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5683)
         );
  NAND2_X1 U6761 ( .A1(n3492), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U6762 ( .A1(n5654), .A2(n5645), .ZN(n5677) );
  INV_X1 U6763 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U6764 ( .A1(n5648), .A2(n6638), .ZN(n5646) );
  XNOR2_X1 U6765 ( .A(n5648), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5671)
         );
  NOR2_X1 U6766 ( .A1(n5648), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5664)
         );
  INV_X1 U6767 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6549) );
  XNOR2_X1 U6768 ( .A(n5649), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5772)
         );
  AND2_X1 U6769 ( .A1(n6240), .A2(REIP_REG_24__SCAN_IN), .ZN(n5770) );
  AOI21_X1 U6770 ( .B1(n6161), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5770), 
        .ZN(n5650) );
  OAI21_X1 U6771 ( .B1(n5868), .B2(n6170), .A(n5650), .ZN(n5651) );
  AOI21_X1 U6772 ( .B1(n5652), .B2(n5681), .A(n5651), .ZN(n5653) );
  OAI21_X1 U6773 ( .B1(n5772), .B2(n6144), .A(n5653), .ZN(U2962) );
  NAND2_X1 U6774 ( .A1(n5786), .A2(n5808), .ZN(n5656) );
  OAI21_X1 U6775 ( .B1(n5654), .B2(n5656), .A(n5655), .ZN(n5657) );
  XNOR2_X1 U6776 ( .A(n5657), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5781)
         );
  NAND2_X1 U6777 ( .A1(n6240), .A2(REIP_REG_23__SCAN_IN), .ZN(n5775) );
  OAI21_X1 U6778 ( .B1(n5725), .B2(n5658), .A(n5775), .ZN(n5661) );
  NOR2_X1 U6779 ( .A1(n5659), .A2(n6139), .ZN(n5660) );
  AOI211_X1 U6780 ( .C1(n5728), .C2(n5662), .A(n5661), .B(n5660), .ZN(n5663)
         );
  OAI21_X1 U6781 ( .B1(n5781), .B2(n6144), .A(n5663), .ZN(U2963) );
  AOI21_X1 U6782 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5648), .A(n5664), 
        .ZN(n5666) );
  XOR2_X1 U6783 ( .A(n5666), .B(n5665), .Z(n5790) );
  NAND2_X1 U6784 ( .A1(n6240), .A2(REIP_REG_22__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U6785 ( .A1(n6161), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5667)
         );
  OAI211_X1 U6786 ( .C1(n5882), .C2(n6170), .A(n5783), .B(n5667), .ZN(n5668)
         );
  AOI21_X1 U6787 ( .B1(n5912), .B2(n5681), .A(n5668), .ZN(n5669) );
  OAI21_X1 U6788 ( .B1(n5790), .B2(n6144), .A(n5669), .ZN(U2964) );
  OAI21_X1 U6789 ( .B1(n5671), .B2(n5670), .A(n2975), .ZN(n5791) );
  NAND2_X1 U6790 ( .A1(n5791), .A2(n6165), .ZN(n5675) );
  NAND2_X1 U6791 ( .A1(n6240), .A2(REIP_REG_21__SCAN_IN), .ZN(n5792) );
  OAI21_X1 U6792 ( .B1(n5725), .B2(n5672), .A(n5792), .ZN(n5673) );
  AOI21_X1 U6793 ( .B1(n5894), .B2(n5728), .A(n5673), .ZN(n5674) );
  OAI211_X1 U6794 ( .C1(n6139), .C2(n5895), .A(n5675), .B(n5674), .ZN(U2965)
         );
  XNOR2_X1 U6795 ( .A(n5648), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5676)
         );
  XNOR2_X1 U6796 ( .A(n5677), .B(n5676), .ZN(n5812) );
  NOR2_X1 U6797 ( .A1(n5910), .A2(n6170), .ZN(n5680) );
  NAND2_X1 U6798 ( .A1(n6240), .A2(REIP_REG_20__SCAN_IN), .ZN(n5804) );
  OAI21_X1 U6799 ( .B1(n5725), .B2(n5678), .A(n5804), .ZN(n5679) );
  AOI211_X1 U6800 ( .C1(n5918), .C2(n5681), .A(n5680), .B(n5679), .ZN(n5682)
         );
  OAI21_X1 U6801 ( .B1(n5812), .B2(n6144), .A(n5682), .ZN(U2966) );
  OR2_X1 U6802 ( .A1(n5684), .A2(n5683), .ZN(n5814) );
  NAND3_X1 U6803 ( .A1(n5814), .A2(n6165), .A3(n5654), .ZN(n5689) );
  NOR2_X1 U6804 ( .A1(n6196), .A2(n6574), .ZN(n5817) );
  NOR2_X1 U6805 ( .A1(n5725), .A2(n5685), .ZN(n5686) );
  AOI211_X1 U6806 ( .C1(n5687), .C2(n5728), .A(n5817), .B(n5686), .ZN(n5688)
         );
  OAI211_X1 U6807 ( .C1(n6139), .C2(n5921), .A(n5689), .B(n5688), .ZN(U2967)
         );
  NOR3_X1 U6808 ( .A1(n5696), .A2(n3492), .A3(n5824), .ZN(n5700) );
  NAND2_X1 U6809 ( .A1(n3492), .A2(n5934), .ZN(n5709) );
  NOR3_X1 U6810 ( .A1(n5690), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5709), 
        .ZN(n5698) );
  NOR2_X1 U6811 ( .A1(n5700), .A2(n5698), .ZN(n5691) );
  XNOR2_X1 U6812 ( .A(n5691), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5823)
         );
  NAND2_X1 U6813 ( .A1(n5823), .A2(n6165), .ZN(n5695) );
  INV_X1 U6814 ( .A(REIP_REG_18__SCAN_IN), .ZN(n5692) );
  NOR2_X1 U6815 ( .A1(n6196), .A2(n5692), .ZN(n5826) );
  NOR2_X1 U6816 ( .A1(n5975), .A2(n6170), .ZN(n5693) );
  AOI211_X1 U6817 ( .C1(n6161), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5826), 
        .B(n5693), .ZN(n5694) );
  OAI211_X1 U6818 ( .C1(n6139), .C2(n5971), .A(n5695), .B(n5694), .ZN(U2968)
         );
  AOI21_X1 U6819 ( .B1(n3492), .B2(n5824), .A(n5696), .ZN(n5697) );
  AOI21_X1 U6820 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5709), .A(n5697), 
        .ZN(n5701) );
  INV_X1 U6821 ( .A(n5698), .ZN(n5699) );
  OAI21_X1 U6822 ( .B1(n5701), .B2(n5700), .A(n5699), .ZN(n5930) );
  NAND2_X1 U6823 ( .A1(n5930), .A2(n6165), .ZN(n5707) );
  INV_X1 U6824 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5702) );
  OAI22_X1 U6825 ( .A1(n5725), .A2(n5703), .B1(n6196), .B2(n5702), .ZN(n5704)
         );
  AOI21_X1 U6826 ( .B1(n5728), .B2(n5705), .A(n5704), .ZN(n5706) );
  OAI211_X1 U6827 ( .C1(n6139), .C2(n5708), .A(n5707), .B(n5706), .ZN(U2969)
         );
  OAI21_X1 U6828 ( .B1(n3492), .B2(n5934), .A(n5709), .ZN(n5711) );
  XOR2_X1 U6829 ( .A(n5711), .B(n5710), .Z(n5937) );
  INV_X1 U6830 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5712) );
  OAI22_X1 U6831 ( .A1(n5725), .A2(n5712), .B1(n6196), .B2(n6474), .ZN(n5714)
         );
  NOR2_X1 U6832 ( .A1(n6080), .A2(n6139), .ZN(n5713) );
  AOI211_X1 U6833 ( .C1(n5728), .C2(n5715), .A(n5714), .B(n5713), .ZN(n5716)
         );
  OAI21_X1 U6834 ( .B1(n5937), .B2(n6144), .A(n5716), .ZN(U2970) );
  INV_X1 U6835 ( .A(n5690), .ZN(n5718) );
  AOI21_X1 U6836 ( .B1(n5719), .B2(n5717), .A(n5718), .ZN(n5841) );
  INV_X1 U6837 ( .A(n5980), .ZN(n6062) );
  NAND2_X1 U6838 ( .A1(n6161), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5720)
         );
  NAND2_X1 U6839 ( .A1(n6240), .A2(REIP_REG_15__SCAN_IN), .ZN(n5837) );
  OAI211_X1 U6840 ( .C1(n6170), .C2(n5982), .A(n5720), .B(n5837), .ZN(n5721)
         );
  AOI21_X1 U6841 ( .B1(n6062), .B2(n5681), .A(n5721), .ZN(n5722) );
  OAI21_X1 U6842 ( .B1(n5841), .B2(n6144), .A(n5722), .ZN(U2971) );
  XNOR2_X1 U6843 ( .A(n5648), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5724)
         );
  XNOR2_X1 U6844 ( .A(n5723), .B(n5724), .ZN(n5842) );
  NAND2_X1 U6845 ( .A1(n5842), .A2(n6165), .ZN(n5730) );
  OAI22_X1 U6846 ( .A1(n5725), .A2(n3928), .B1(n6196), .B2(n6471), .ZN(n5726)
         );
  AOI21_X1 U6847 ( .B1(n5728), .B2(n5727), .A(n5726), .ZN(n5729) );
  OAI211_X1 U6848 ( .C1(n6139), .C2(n5731), .A(n5730), .B(n5729), .ZN(U2972)
         );
  NOR2_X1 U6849 ( .A1(n5732), .A2(n6198), .ZN(n5733) );
  AOI211_X1 U6850 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5746), .A(n5734), .B(n5733), .ZN(n5739) );
  NAND3_X1 U6851 ( .A1(n5737), .A2(n5736), .A3(n5735), .ZN(n5738) );
  OAI211_X1 U6852 ( .C1(n5740), .C2(n6184), .A(n5739), .B(n5738), .ZN(U2990)
         );
  OAI21_X1 U6853 ( .B1(n5742), .B2(n6198), .A(n5741), .ZN(n5745) );
  NOR2_X1 U6854 ( .A1(n5743), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5744)
         );
  AOI211_X1 U6855 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5746), .A(n5745), .B(n5744), .ZN(n5747) );
  OAI21_X1 U6856 ( .B1(n5748), .B2(n6184), .A(n5747), .ZN(U2991) );
  INV_X1 U6857 ( .A(n5767), .ZN(n5763) );
  OAI21_X1 U6858 ( .B1(n5750), .B2(n6198), .A(n5749), .ZN(n5751) );
  AOI21_X1 U6859 ( .B1(n5763), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5751), 
        .ZN(n5756) );
  INV_X1 U6860 ( .A(n5752), .ZN(n5754) );
  NAND3_X1 U6861 ( .A1(n5758), .A2(n5754), .A3(n5753), .ZN(n5755) );
  OAI211_X1 U6862 ( .C1(n5757), .C2(n6184), .A(n5756), .B(n5755), .ZN(U2992)
         );
  INV_X1 U6863 ( .A(n5758), .ZN(n5766) );
  NAND2_X1 U6864 ( .A1(n5759), .A2(n6242), .ZN(n5765) );
  OAI21_X1 U6865 ( .B1(n5761), .B2(n6198), .A(n5760), .ZN(n5762) );
  AOI21_X1 U6866 ( .B1(n5763), .B2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5762), 
        .ZN(n5764) );
  OAI211_X1 U6867 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5766), .A(n5765), .B(n5764), .ZN(U2993) );
  AOI21_X1 U6868 ( .B1(n5779), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5768) );
  NOR2_X1 U6869 ( .A1(n5768), .A2(n5767), .ZN(n5769) );
  AOI211_X1 U6870 ( .C1(n6237), .C2(n5873), .A(n5770), .B(n5769), .ZN(n5771)
         );
  OAI21_X1 U6871 ( .B1(n5772), .B2(n6184), .A(n5771), .ZN(U2994) );
  NAND2_X1 U6872 ( .A1(n5773), .A2(n6237), .ZN(n5774) );
  OAI211_X1 U6873 ( .C1(n5776), .C2(n5778), .A(n5775), .B(n5774), .ZN(n5777)
         );
  AOI21_X1 U6874 ( .B1(n5779), .B2(n5778), .A(n5777), .ZN(n5780) );
  OAI21_X1 U6875 ( .B1(n5781), .B2(n6184), .A(n5780), .ZN(U2995) );
  INV_X1 U6876 ( .A(n5782), .ZN(n5794) );
  OAI21_X1 U6877 ( .B1(n6198), .B2(n5885), .A(n5783), .ZN(n5788) );
  INV_X1 U6878 ( .A(n5784), .ZN(n5797) );
  NOR3_X1 U6879 ( .A1(n5797), .A2(n5786), .A3(n5785), .ZN(n5787) );
  AOI211_X1 U6880 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5794), .A(n5788), .B(n5787), .ZN(n5789) );
  OAI21_X1 U6881 ( .B1(n5790), .B2(n6184), .A(n5789), .ZN(U2996) );
  NAND2_X1 U6882 ( .A1(n5791), .A2(n6242), .ZN(n5796) );
  OAI21_X1 U6883 ( .B1(n6198), .B2(n5896), .A(n5792), .ZN(n5793) );
  AOI21_X1 U6884 ( .B1(n5794), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5793), 
        .ZN(n5795) );
  OAI211_X1 U6885 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5797), .A(n5796), .B(n5795), .ZN(U2997) );
  AND2_X1 U6886 ( .A1(n5798), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5803)
         );
  NAND2_X1 U6887 ( .A1(n5800), .A2(n5799), .ZN(n5801) );
  OAI21_X1 U6888 ( .B1(n5803), .B2(n5802), .A(n5801), .ZN(n5928) );
  AOI21_X1 U6889 ( .B1(n6244), .B2(n5824), .A(n5928), .ZN(n5830) );
  OAI21_X1 U6890 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5831), .A(n5830), 
        .ZN(n5813) );
  OAI21_X1 U6891 ( .B1(n6198), .B2(n5903), .A(n5804), .ZN(n5810) );
  INV_X1 U6892 ( .A(n5933), .ZN(n5806) );
  NAND2_X1 U6893 ( .A1(n5806), .A2(n5805), .ZN(n5815) );
  NOR3_X1 U6894 ( .A1(n5815), .A2(n5808), .A3(n5807), .ZN(n5809) );
  AOI211_X1 U6895 ( .C1(n5813), .C2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5810), .B(n5809), .ZN(n5811) );
  OAI21_X1 U6896 ( .B1(n5812), .B2(n6184), .A(n5811), .ZN(U2998) );
  INV_X1 U6897 ( .A(n5813), .ZN(n5822) );
  INV_X1 U6898 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5821) );
  NAND3_X1 U6899 ( .A1(n5814), .A2(n6242), .A3(n5654), .ZN(n5820) );
  NOR2_X1 U6900 ( .A1(n5815), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5816)
         );
  AOI211_X1 U6901 ( .C1(n6237), .C2(n5818), .A(n5817), .B(n5816), .ZN(n5819)
         );
  OAI211_X1 U6902 ( .C1(n5822), .C2(n5821), .A(n5820), .B(n5819), .ZN(U2999)
         );
  NAND2_X1 U6903 ( .A1(n5823), .A2(n6242), .ZN(n5828) );
  NOR3_X1 U6904 ( .A1(n5933), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n5824), 
        .ZN(n5825) );
  AOI211_X1 U6905 ( .C1(n6237), .C2(n5972), .A(n5826), .B(n5825), .ZN(n5827)
         );
  OAI211_X1 U6906 ( .C1(n5830), .C2(n5829), .A(n5828), .B(n5827), .ZN(U3000)
         );
  INV_X1 U6907 ( .A(n5833), .ZN(n5832) );
  OAI21_X1 U6908 ( .B1(n5832), .B2(n5831), .A(n6180), .ZN(n5939) );
  NOR3_X1 U6909 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n6179), .A3(n5833), 
        .ZN(n5940) );
  AOI21_X1 U6910 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n5939), .A(n5940), 
        .ZN(n5840) );
  AOI21_X1 U6911 ( .B1(n5836), .B2(n5835), .A(n5834), .ZN(n6061) );
  INV_X1 U6912 ( .A(n5837), .ZN(n5838) );
  AOI21_X1 U6913 ( .B1(n6237), .B2(n6061), .A(n5838), .ZN(n5839) );
  OAI211_X1 U6914 ( .C1(n5841), .C2(n6184), .A(n5840), .B(n5839), .ZN(U3003)
         );
  NAND2_X1 U6915 ( .A1(n5842), .A2(n6242), .ZN(n5851) );
  INV_X1 U6916 ( .A(n6179), .ZN(n6174) );
  NAND3_X1 U6917 ( .A1(n6174), .A2(n5843), .A3(n3502), .ZN(n5850) );
  OAI22_X1 U6918 ( .A1(n6198), .A2(n5844), .B1(n6471), .B2(n6196), .ZN(n5845)
         );
  INV_X1 U6919 ( .A(n5845), .ZN(n5849) );
  OAI21_X1 U6920 ( .B1(n5847), .B2(n5846), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5848) );
  NAND4_X1 U6921 ( .A1(n5851), .A2(n5850), .A3(n5849), .A4(n5848), .ZN(U3004)
         );
  OAI211_X1 U6922 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n2963), .A(n5852), .B(
        n6310), .ZN(n5853) );
  OAI21_X1 U6923 ( .B1(n5858), .B2(n5854), .A(n5853), .ZN(n5855) );
  MUX2_X1 U6924 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5855), .S(n6249), 
        .Z(U3464) );
  XNOR2_X1 U6925 ( .A(n5857), .B(n5856), .ZN(n5860) );
  OAI22_X1 U6926 ( .A1(n5860), .A2(n6297), .B1(n5859), .B2(n5858), .ZN(n5861)
         );
  MUX2_X1 U6927 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5861), .S(n6249), 
        .Z(U3463) );
  INV_X1 U6928 ( .A(n5862), .ZN(n5864) );
  OAI22_X1 U6929 ( .A1(n5864), .A2(n6420), .B1(n5863), .B2(n6415), .ZN(n5866)
         );
  MUX2_X1 U6930 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5866), .S(n5865), 
        .Z(U3456) );
  AND2_X1 U6931 ( .A1(n5867), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U6932 ( .A(n5868), .ZN(n5872) );
  INV_X1 U6933 ( .A(REIP_REG_24__SCAN_IN), .ZN(n5877) );
  OAI22_X1 U6934 ( .A1(n5877), .A2(n5870), .B1(n5869), .B2(n6035), .ZN(n5871)
         );
  AOI21_X1 U6935 ( .B1(n5872), .B2(n6057), .A(n5871), .ZN(n5880) );
  INV_X1 U6936 ( .A(n5873), .ZN(n5874) );
  OAI22_X1 U6937 ( .A1(n5875), .A2(n6024), .B1(n5874), .B2(n5988), .ZN(n5876)
         );
  AOI21_X1 U6938 ( .B1(n5878), .B2(n5877), .A(n5876), .ZN(n5879) );
  OAI211_X1 U6939 ( .C1(n5881), .C2(n6029), .A(n5880), .B(n5879), .ZN(U2803)
         );
  AOI22_X1 U6940 ( .A1(EBX_REG_22__SCAN_IN), .A2(n6048), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6046), .ZN(n5893) );
  INV_X1 U6941 ( .A(n5882), .ZN(n5884) );
  INV_X1 U6942 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6483) );
  AOI22_X1 U6943 ( .A1(n5884), .A2(n6057), .B1(n5883), .B2(n6483), .ZN(n5892)
         );
  INV_X1 U6944 ( .A(n5885), .ZN(n5886) );
  AOI22_X1 U6945 ( .A1(n5912), .A2(n6038), .B1(n5886), .B2(n6047), .ZN(n5891)
         );
  NOR2_X1 U6946 ( .A1(n5888), .A2(n5887), .ZN(n5907) );
  NOR2_X1 U6947 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5889), .ZN(n5898) );
  OAI21_X1 U6948 ( .B1(n5907), .B2(n5898), .A(REIP_REG_22__SCAN_IN), .ZN(n5890) );
  NAND4_X1 U6949 ( .A1(n5893), .A2(n5892), .A3(n5891), .A4(n5890), .ZN(U2805)
         );
  AOI22_X1 U6950 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6048), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6046), .ZN(n5902) );
  AOI22_X1 U6951 ( .A1(n5894), .A2(n6057), .B1(REIP_REG_21__SCAN_IN), .B2(
        n5907), .ZN(n5901) );
  INV_X1 U6952 ( .A(n5895), .ZN(n5915) );
  INV_X1 U6953 ( .A(n5896), .ZN(n5897) );
  AOI22_X1 U6954 ( .A1(n5915), .A2(n6038), .B1(n6047), .B2(n5897), .ZN(n5900)
         );
  INV_X1 U6955 ( .A(n5898), .ZN(n5899) );
  NAND4_X1 U6956 ( .A1(n5902), .A2(n5901), .A3(n5900), .A4(n5899), .ZN(U2806)
         );
  AOI22_X1 U6957 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6048), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6046), .ZN(n5909) );
  OAI22_X1 U6958 ( .A1(n5904), .A2(n6024), .B1(n5988), .B2(n5903), .ZN(n5905)
         );
  AOI221_X1 U6959 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5907), .C1(n5906), .C2(
        n5907), .A(n5905), .ZN(n5908) );
  OAI211_X1 U6960 ( .C1(n5910), .C2(n6041), .A(n5909), .B(n5908), .ZN(U2807)
         );
  INV_X1 U6961 ( .A(n5911), .ZN(n6082) );
  AOI22_X1 U6962 ( .A1(n5912), .A2(n6082), .B1(n6081), .B2(DATAI_22_), .ZN(
        n5914) );
  AOI22_X1 U6963 ( .A1(n6085), .A2(DATAI_6_), .B1(n6084), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U6964 ( .A1(n5914), .A2(n5913), .ZN(U2869) );
  AOI22_X1 U6965 ( .A1(n5915), .A2(n6082), .B1(n6081), .B2(DATAI_21_), .ZN(
        n5917) );
  AOI22_X1 U6966 ( .A1(n6085), .A2(DATAI_5_), .B1(n6084), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U6967 ( .A1(n5917), .A2(n5916), .ZN(U2870) );
  AOI22_X1 U6968 ( .A1(n5918), .A2(n6082), .B1(n6081), .B2(DATAI_20_), .ZN(
        n5920) );
  AOI22_X1 U6969 ( .A1(n6085), .A2(DATAI_4_), .B1(n6084), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U6970 ( .A1(n5920), .A2(n5919), .ZN(U2871) );
  INV_X1 U6971 ( .A(n5921), .ZN(n5922) );
  AOI22_X1 U6972 ( .A1(n5922), .A2(n6082), .B1(n6081), .B2(DATAI_19_), .ZN(
        n5924) );
  AOI22_X1 U6973 ( .A1(n6085), .A2(DATAI_3_), .B1(n6084), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U6974 ( .A1(n5924), .A2(n5923), .ZN(U2872) );
  AOI22_X1 U6975 ( .A1(n6240), .A2(REIP_REG_13__SCAN_IN), .B1(n6161), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5927) );
  AOI22_X1 U6976 ( .A1(n5925), .A2(n6165), .B1(n5681), .B2(n5994), .ZN(n5926)
         );
  OAI211_X1 U6977 ( .C1(n6170), .C2(n5998), .A(n5927), .B(n5926), .ZN(U2973)
         );
  AOI22_X1 U6978 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5928), .B1(n6240), .B2(REIP_REG_17__SCAN_IN), .ZN(n5932) );
  AOI22_X1 U6979 ( .A1(n5930), .A2(n6242), .B1(n6237), .B2(n5929), .ZN(n5931)
         );
  OAI211_X1 U6980 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5933), .A(n5932), .B(n5931), .ZN(U3001) );
  NAND2_X1 U6981 ( .A1(n5935), .A2(n5934), .ZN(n5943) );
  OAI22_X1 U6982 ( .A1(n5937), .A2(n6184), .B1(n6198), .B2(n5936), .ZN(n5938)
         );
  AOI221_X1 U6983 ( .B1(n5940), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .C1(
        n5939), .C2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5938), .ZN(n5942) );
  NAND2_X1 U6984 ( .A1(n6240), .A2(REIP_REG_16__SCAN_IN), .ZN(n5941) );
  OAI211_X1 U6985 ( .C1(n6179), .C2(n5943), .A(n5942), .B(n5941), .ZN(U3002)
         );
  INV_X1 U6986 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6441) );
  NOR2_X1 U6987 ( .A1(n6441), .A2(STATE_REG_0__SCAN_IN), .ZN(n6500) );
  OAI21_X1 U6988 ( .B1(STATE_REG_2__SCAN_IN), .B2(n6441), .A(
        STATE_REG_0__SCAN_IN), .ZN(n5949) );
  NOR2_X1 U6989 ( .A1(ADS_N_REG_SCAN_IN), .A2(n5949), .ZN(n5944) );
  NOR2_X1 U6990 ( .A1(n6500), .A2(n5944), .ZN(U2789) );
  OAI21_X1 U6991 ( .B1(n5945), .B2(n6418), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5946) );
  OAI21_X1 U6992 ( .B1(n5947), .B2(n6421), .A(n5946), .ZN(U2790) );
  INV_X2 U6993 ( .A(n6500), .ZN(n6529) );
  NOR2_X1 U6994 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5950) );
  OAI21_X1 U6995 ( .B1(n5950), .B2(D_C_N_REG_SCAN_IN), .A(n6529), .ZN(n5948)
         );
  OAI21_X1 U6996 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6529), .A(n5948), .ZN(
        U2791) );
  NAND2_X1 U6997 ( .A1(n6529), .A2(n5949), .ZN(n6688) );
  INV_X1 U6998 ( .A(n6688), .ZN(n6505) );
  OAI21_X1 U6999 ( .B1(n5950), .B2(BS16_N), .A(n6505), .ZN(n6503) );
  OAI21_X1 U7000 ( .B1(n6505), .B2(n6424), .A(n6503), .ZN(U2792) );
  OAI21_X1 U7001 ( .B1(n5951), .B2(n6577), .A(n6144), .ZN(U2793) );
  NOR4_X1 U7002 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n5955) );
  NOR4_X1 U7003 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n5954) );
  NOR4_X1 U7004 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5953) );
  NOR4_X1 U7005 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5952) );
  NAND4_X1 U7006 ( .A1(n5955), .A2(n5954), .A3(n5953), .A4(n5952), .ZN(n5961)
         );
  NOR4_X1 U7007 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_24__SCAN_IN), .ZN(n5959) );
  AOI211_X1 U7008 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_2__SCAN_IN), .B(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n5958) );
  NOR4_X1 U7009 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(
        n5957) );
  NOR4_X1 U7010 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n5956) );
  NAND4_X1 U7011 ( .A1(n5959), .A2(n5958), .A3(n5957), .A4(n5956), .ZN(n5960)
         );
  NOR2_X1 U7012 ( .A1(n5961), .A2(n5960), .ZN(n6516) );
  INV_X1 U7013 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5963) );
  NOR3_X1 U7014 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5964) );
  OAI21_X1 U7015 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5964), .A(n6516), .ZN(n5962)
         );
  OAI21_X1 U7016 ( .B1(n6516), .B2(n5963), .A(n5962), .ZN(U2794) );
  INV_X1 U7017 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6504) );
  AOI21_X1 U7018 ( .B1(n6509), .B2(n6504), .A(n5964), .ZN(n5966) );
  INV_X1 U7019 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5965) );
  INV_X1 U7020 ( .A(n6516), .ZN(n6511) );
  AOI22_X1 U7021 ( .A1(n6516), .A2(n5966), .B1(n5965), .B2(n6511), .ZN(U2795)
         );
  AOI21_X1 U7022 ( .B1(n6046), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6020), 
        .ZN(n5967) );
  OAI221_X1 U7023 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5969), .C1(n5692), .C2(
        n5968), .A(n5967), .ZN(n5970) );
  AOI21_X1 U7024 ( .B1(EBX_REG_18__SCAN_IN), .B2(n6048), .A(n5970), .ZN(n5974)
         );
  INV_X1 U7025 ( .A(n5971), .ZN(n6077) );
  AOI22_X1 U7026 ( .A1(n6077), .A2(n6038), .B1(n6047), .B2(n5972), .ZN(n5973)
         );
  OAI211_X1 U7027 ( .C1(n5975), .C2(n6041), .A(n5974), .B(n5973), .ZN(U2809)
         );
  AOI22_X1 U7028 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6048), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5976), .ZN(n5979) );
  AOI211_X1 U7029 ( .C1(n6046), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6020), 
        .B(n5977), .ZN(n5978) );
  OAI211_X1 U7030 ( .C1(n5980), .C2(n6024), .A(n5979), .B(n5978), .ZN(n5981)
         );
  INV_X1 U7031 ( .A(n5981), .ZN(n5985) );
  INV_X1 U7032 ( .A(n5982), .ZN(n5983) );
  AOI22_X1 U7033 ( .A1(n6057), .A2(n5983), .B1(n6061), .B2(n6047), .ZN(n5984)
         );
  NAND2_X1 U7034 ( .A1(n5985), .A2(n5984), .ZN(U2812) );
  NAND2_X1 U7035 ( .A1(n6046), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5986)
         );
  OAI211_X1 U7036 ( .C1(n5988), .C2(n5987), .A(n6033), .B(n5986), .ZN(n5989)
         );
  INV_X1 U7037 ( .A(n5989), .ZN(n5992) );
  NAND3_X1 U7038 ( .A1(n6002), .A2(n5347), .A3(n5990), .ZN(n5991) );
  OAI211_X1 U7039 ( .C1(n3652), .C2(n6029), .A(n5992), .B(n5991), .ZN(n5993)
         );
  AOI21_X1 U7040 ( .B1(n5994), .B2(n6038), .A(n5993), .ZN(n5997) );
  OAI21_X1 U7041 ( .B1(n5995), .B2(n6003), .A(REIP_REG_13__SCAN_IN), .ZN(n5996) );
  OAI211_X1 U7042 ( .C1(n6041), .C2(n5998), .A(n5997), .B(n5996), .ZN(U2814)
         );
  AOI22_X1 U7043 ( .A1(EBX_REG_11__SCAN_IN), .A2(n6048), .B1(
        PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n6046), .ZN(n6008) );
  AOI21_X1 U7044 ( .B1(n6047), .B2(n6178), .A(n6020), .ZN(n6007) );
  INV_X1 U7045 ( .A(n5999), .ZN(n6138) );
  OAI22_X1 U7046 ( .A1(n6140), .A2(n6024), .B1(n6041), .B2(n6138), .ZN(n6000)
         );
  INV_X1 U7047 ( .A(n6000), .ZN(n6006) );
  AND2_X1 U7048 ( .A1(n6002), .A2(n6001), .ZN(n6004) );
  OAI21_X1 U7049 ( .B1(n6004), .B2(REIP_REG_11__SCAN_IN), .A(n6003), .ZN(n6005) );
  NAND4_X1 U7050 ( .A1(n6008), .A2(n6007), .A3(n6006), .A4(n6005), .ZN(U2816)
         );
  NAND2_X1 U7051 ( .A1(n6010), .A2(n6009), .ZN(n6013) );
  INV_X1 U7052 ( .A(n6011), .ZN(n6012) );
  NAND2_X1 U7053 ( .A1(n6013), .A2(n6012), .ZN(n6065) );
  INV_X1 U7054 ( .A(n6065), .ZN(n6188) );
  INV_X1 U7055 ( .A(n6014), .ZN(n6015) );
  NOR3_X1 U7056 ( .A1(n6016), .A2(REIP_REG_9__SCAN_IN), .A3(n6015), .ZN(n6017)
         );
  AOI21_X1 U7057 ( .B1(n6188), .B2(n6047), .A(n6017), .ZN(n6028) );
  OAI22_X1 U7058 ( .A1(n6576), .A2(n6029), .B1(n6018), .B2(n6035), .ZN(n6019)
         );
  AOI211_X1 U7059 ( .C1(REIP_REG_9__SCAN_IN), .C2(n6021), .A(n6020), .B(n6019), 
        .ZN(n6027) );
  INV_X1 U7060 ( .A(n6022), .ZN(n6023) );
  OAI22_X1 U7061 ( .A1(n6066), .A2(n6024), .B1(n6041), .B2(n6023), .ZN(n6025)
         );
  INV_X1 U7062 ( .A(n6025), .ZN(n6026) );
  NAND3_X1 U7063 ( .A1(n6028), .A2(n6027), .A3(n6026), .ZN(U2818) );
  NOR2_X1 U7064 ( .A1(n6537), .A2(n6029), .ZN(n6030) );
  AOI211_X1 U7065 ( .C1(n6032), .C2(REIP_REG_6__SCAN_IN), .A(n6031), .B(n6030), 
        .ZN(n6040) );
  INV_X1 U7066 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7067 ( .A1(n6047), .A2(n6216), .ZN(n6034) );
  OAI211_X1 U7068 ( .C1(n6036), .C2(n6035), .A(n6034), .B(n6033), .ZN(n6037)
         );
  AOI21_X1 U7069 ( .B1(n6149), .B2(n6038), .A(n6037), .ZN(n6039) );
  OAI211_X1 U7070 ( .C1(n6152), .C2(n6041), .A(n6040), .B(n6039), .ZN(U2821)
         );
  INV_X1 U7071 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6453) );
  NAND2_X1 U7072 ( .A1(n6042), .A2(REIP_REG_2__SCAN_IN), .ZN(n6059) );
  INV_X1 U7073 ( .A(n6160), .ZN(n6056) );
  AOI21_X1 U7074 ( .B1(n6045), .B2(n6044), .A(n6043), .ZN(n6228) );
  AOI22_X1 U7075 ( .A1(n6047), .A2(n6228), .B1(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .B2(n6046), .ZN(n6050) );
  NAND2_X1 U7076 ( .A1(n6048), .A2(EBX_REG_3__SCAN_IN), .ZN(n6049) );
  OAI211_X1 U7077 ( .C1(n6052), .C2(n6051), .A(n6050), .B(n6049), .ZN(n6055)
         );
  NOR2_X1 U7078 ( .A1(n6053), .A2(n6069), .ZN(n6054) );
  AOI211_X1 U7079 ( .C1(n6057), .C2(n6056), .A(n6055), .B(n6054), .ZN(n6058)
         );
  OAI221_X1 U7080 ( .B1(n6060), .B2(n6453), .C1(n6060), .C2(n6059), .A(n6058), 
        .ZN(U2824) );
  AOI22_X1 U7081 ( .A1(n6062), .A2(n6073), .B1(n4255), .B2(n6061), .ZN(n6063)
         );
  OAI21_X1 U7082 ( .B1(n6076), .B2(n6064), .A(n6063), .ZN(U2844) );
  OAI22_X1 U7083 ( .A1(n6066), .A2(n5579), .B1(n5578), .B2(n6065), .ZN(n6067)
         );
  INV_X1 U7084 ( .A(n6067), .ZN(n6068) );
  OAI21_X1 U7085 ( .B1(n6076), .B2(n6576), .A(n6068), .ZN(U2850) );
  INV_X1 U7086 ( .A(n6069), .ZN(n6157) );
  AOI22_X1 U7087 ( .A1(n6157), .A2(n6073), .B1(n4255), .B2(n6228), .ZN(n6070)
         );
  OAI21_X1 U7088 ( .B1(n6076), .B2(n6071), .A(n6070), .ZN(U2856) );
  INV_X1 U7089 ( .A(n6072), .ZN(n6166) );
  AOI22_X1 U7090 ( .A1(n6166), .A2(n6073), .B1(n4255), .B2(n6238), .ZN(n6074)
         );
  OAI21_X1 U7091 ( .B1(n6076), .B2(n6075), .A(n6074), .ZN(U2857) );
  AOI22_X1 U7092 ( .A1(n6077), .A2(n6082), .B1(n6081), .B2(DATAI_18_), .ZN(
        n6079) );
  AOI22_X1 U7093 ( .A1(n6085), .A2(DATAI_2_), .B1(n6084), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7094 ( .A1(n6079), .A2(n6078), .ZN(U2873) );
  INV_X1 U7095 ( .A(n6080), .ZN(n6083) );
  AOI22_X1 U7096 ( .A1(n6083), .A2(n6082), .B1(n6081), .B2(DATAI_16_), .ZN(
        n6087) );
  AOI22_X1 U7097 ( .A1(n6085), .A2(DATAI_0_), .B1(n6084), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7098 ( .A1(n6087), .A2(n6086), .ZN(U2875) );
  AOI22_X1 U7099 ( .A1(n6521), .A2(LWORD_REG_15__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6089) );
  OAI21_X1 U7100 ( .B1(n6090), .B2(n6115), .A(n6089), .ZN(U2908) );
  INV_X1 U7101 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6092) );
  AOI22_X1 U7102 ( .A1(n6521), .A2(LWORD_REG_14__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6091) );
  OAI21_X1 U7103 ( .B1(n6092), .B2(n6115), .A(n6091), .ZN(U2909) );
  INV_X1 U7104 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6094) );
  AOI22_X1 U7105 ( .A1(n6521), .A2(LWORD_REG_13__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6093) );
  OAI21_X1 U7106 ( .B1(n6094), .B2(n6115), .A(n6093), .ZN(U2910) );
  AOI22_X1 U7107 ( .A1(n6521), .A2(LWORD_REG_12__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6095) );
  OAI21_X1 U7108 ( .B1(n6598), .B2(n6115), .A(n6095), .ZN(U2911) );
  INV_X1 U7109 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6097) );
  AOI22_X1 U7110 ( .A1(n6521), .A2(LWORD_REG_11__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6096) );
  OAI21_X1 U7111 ( .B1(n6097), .B2(n6115), .A(n6096), .ZN(U2912) );
  AOI22_X1 U7112 ( .A1(n6521), .A2(LWORD_REG_10__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6098) );
  OAI21_X1 U7113 ( .B1(n6641), .B2(n6115), .A(n6098), .ZN(U2913) );
  INV_X1 U7114 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6100) );
  AOI22_X1 U7115 ( .A1(n6521), .A2(LWORD_REG_9__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6099) );
  OAI21_X1 U7116 ( .B1(n6100), .B2(n6115), .A(n6099), .ZN(U2914) );
  INV_X1 U7117 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6102) );
  AOI22_X1 U7118 ( .A1(n6521), .A2(LWORD_REG_8__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6101) );
  OAI21_X1 U7119 ( .B1(n6102), .B2(n6115), .A(n6101), .ZN(U2915) );
  AOI22_X1 U7120 ( .A1(n6521), .A2(LWORD_REG_7__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6103) );
  OAI21_X1 U7121 ( .B1(n4703), .B2(n6115), .A(n6103), .ZN(U2916) );
  AOI22_X1 U7122 ( .A1(n6521), .A2(LWORD_REG_6__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6104) );
  OAI21_X1 U7123 ( .B1(n4579), .B2(n6115), .A(n6104), .ZN(U2917) );
  AOI22_X1 U7124 ( .A1(n6521), .A2(LWORD_REG_5__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6105) );
  OAI21_X1 U7125 ( .B1(n6106), .B2(n6115), .A(n6105), .ZN(U2918) );
  AOI22_X1 U7126 ( .A1(n6521), .A2(LWORD_REG_4__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6107) );
  OAI21_X1 U7127 ( .B1(n6108), .B2(n6115), .A(n6107), .ZN(U2919) );
  AOI22_X1 U7128 ( .A1(n6521), .A2(LWORD_REG_3__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6109) );
  OAI21_X1 U7129 ( .B1(n6608), .B2(n6115), .A(n6109), .ZN(U2920) );
  AOI22_X1 U7130 ( .A1(n6521), .A2(LWORD_REG_2__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6110) );
  OAI21_X1 U7131 ( .B1(n6111), .B2(n6115), .A(n6110), .ZN(U2921) );
  AOI22_X1 U7132 ( .A1(n6521), .A2(LWORD_REG_1__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6112) );
  OAI21_X1 U7133 ( .B1(n6113), .B2(n6115), .A(n6112), .ZN(U2922) );
  AOI22_X1 U7134 ( .A1(n6521), .A2(LWORD_REG_0__SCAN_IN), .B1(n5867), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6114) );
  OAI21_X1 U7135 ( .B1(n6116), .B2(n6115), .A(n6114), .ZN(U2923) );
  AOI22_X1 U7136 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6130), .B1(n6129), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n6117) );
  OAI21_X1 U7137 ( .B1(n6119), .B2(n4578), .A(n6117), .ZN(U2945) );
  AOI22_X1 U7138 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6130), .B1(n6129), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n6118) );
  OAI21_X1 U7139 ( .B1(n6119), .B2(n4704), .A(n6118), .ZN(U2946) );
  AOI22_X1 U7140 ( .A1(LWORD_REG_8__SCAN_IN), .A2(n6126), .B1(n6129), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7141 ( .A1(n6131), .A2(DATAI_8_), .ZN(n6120) );
  NAND2_X1 U7142 ( .A1(n6121), .A2(n6120), .ZN(U2947) );
  AOI22_X1 U7143 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n6126), .B1(n6129), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7144 ( .A1(n6131), .A2(DATAI_9_), .ZN(n6122) );
  NAND2_X1 U7145 ( .A1(n6123), .A2(n6122), .ZN(U2948) );
  AOI22_X1 U7146 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6126), .B1(n6129), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n6125) );
  NAND2_X1 U7147 ( .A1(n6131), .A2(DATAI_11_), .ZN(n6124) );
  NAND2_X1 U7148 ( .A1(n6125), .A2(n6124), .ZN(U2950) );
  AOI22_X1 U7149 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n6126), .B1(n6129), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7150 ( .A1(n6131), .A2(DATAI_13_), .ZN(n6127) );
  NAND2_X1 U7151 ( .A1(n6128), .A2(n6127), .ZN(U2952) );
  AOI22_X1 U7152 ( .A1(LWORD_REG_14__SCAN_IN), .A2(n6130), .B1(n6129), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n6133) );
  NAND2_X1 U7153 ( .A1(n6131), .A2(DATAI_14_), .ZN(n6132) );
  NAND2_X1 U7154 ( .A1(n6133), .A2(n6132), .ZN(U2953) );
  NAND2_X1 U7155 ( .A1(n6135), .A2(n6134), .ZN(n6137) );
  XNOR2_X1 U7156 ( .A(n5648), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6136)
         );
  XNOR2_X1 U7157 ( .A(n6137), .B(n6136), .ZN(n6185) );
  AOI22_X1 U7158 ( .A1(n6240), .A2(REIP_REG_11__SCAN_IN), .B1(n6161), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6143) );
  OAI22_X1 U7159 ( .A1(n6140), .A2(n6139), .B1(n6170), .B2(n6138), .ZN(n6141)
         );
  INV_X1 U7160 ( .A(n6141), .ZN(n6142) );
  OAI211_X1 U7161 ( .C1(n6185), .C2(n6144), .A(n6143), .B(n6142), .ZN(U2975)
         );
  AOI22_X1 U7162 ( .A1(n6240), .A2(REIP_REG_6__SCAN_IN), .B1(n6161), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6151) );
  OAI21_X1 U7163 ( .B1(n6147), .B2(n6146), .A(n6145), .ZN(n6148) );
  INV_X1 U7164 ( .A(n6148), .ZN(n6215) );
  AOI22_X1 U7165 ( .A1(n6215), .A2(n6165), .B1(n5681), .B2(n6149), .ZN(n6150)
         );
  OAI211_X1 U7166 ( .C1(n6170), .C2(n6152), .A(n6151), .B(n6150), .ZN(U2980)
         );
  AOI22_X1 U7167 ( .A1(n6240), .A2(REIP_REG_3__SCAN_IN), .B1(n6161), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6159) );
  OR2_X1 U7168 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  AND2_X1 U7169 ( .A1(n6156), .A2(n6155), .ZN(n6229) );
  AOI22_X1 U7170 ( .A1(n6165), .A2(n6229), .B1(n6157), .B2(n5681), .ZN(n6158)
         );
  OAI211_X1 U7171 ( .C1(n6170), .C2(n6160), .A(n6159), .B(n6158), .ZN(U2983)
         );
  AOI22_X1 U7172 ( .A1(n6240), .A2(REIP_REG_2__SCAN_IN), .B1(n6161), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6168) );
  XOR2_X1 U7173 ( .A(n6162), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n6164) );
  XNOR2_X1 U7174 ( .A(n6164), .B(n6163), .ZN(n6241) );
  AOI22_X1 U7175 ( .A1(n6166), .A2(n5681), .B1(n6241), .B2(n6165), .ZN(n6167)
         );
  OAI211_X1 U7176 ( .C1(n6170), .C2(n6169), .A(n6168), .B(n6167), .ZN(U2984)
         );
  AOI222_X1 U7177 ( .A1(n6172), .A2(n6242), .B1(n6237), .B2(n6171), .C1(
        REIP_REG_12__SCAN_IN), .C2(n6240), .ZN(n6176) );
  OAI211_X1 U7178 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A(n6174), .B(n6173), .ZN(n6175) );
  OAI211_X1 U7179 ( .C1(n6180), .C2(n6177), .A(n6176), .B(n6175), .ZN(U3006)
         );
  AOI22_X1 U7180 ( .A1(n6237), .A2(n6178), .B1(n6240), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n6183) );
  OAI22_X1 U7181 ( .A1(n3495), .A2(n6180), .B1(n6179), .B2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6181) );
  INV_X1 U7182 ( .A(n6181), .ZN(n6182) );
  OAI211_X1 U7183 ( .C1(n6185), .C2(n6184), .A(n6183), .B(n6182), .ZN(U3007)
         );
  INV_X1 U7184 ( .A(n6186), .ZN(n6187) );
  AOI21_X1 U7185 ( .B1(n6237), .B2(n6188), .A(n6187), .ZN(n6192) );
  AOI22_X1 U7186 ( .A1(n6190), .A2(n6242), .B1(n6189), .B2(n6193), .ZN(n6191)
         );
  OAI211_X1 U7187 ( .C1(n6194), .C2(n6193), .A(n6192), .B(n6191), .ZN(U3009)
         );
  OAI21_X1 U7188 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6195), .ZN(n6204) );
  OAI22_X1 U7189 ( .A1(n6198), .A2(n6197), .B1(n6462), .B2(n6196), .ZN(n6199)
         );
  INV_X1 U7190 ( .A(n6199), .ZN(n6203) );
  INV_X1 U7191 ( .A(n6200), .ZN(n6201) );
  AOI22_X1 U7192 ( .A1(n6201), .A2(n6242), .B1(INSTADDRPOINTER_REG_8__SCAN_IN), 
        .B2(n6210), .ZN(n6202) );
  OAI211_X1 U7193 ( .C1(n6213), .C2(n6204), .A(n6203), .B(n6202), .ZN(U3010)
         );
  INV_X1 U7194 ( .A(n6205), .ZN(n6206) );
  AOI21_X1 U7195 ( .B1(n6237), .B2(n6207), .A(n6206), .ZN(n6212) );
  INV_X1 U7196 ( .A(n6208), .ZN(n6209) );
  AOI22_X1 U7197 ( .A1(n6210), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .B1(n6209), 
        .B2(n6242), .ZN(n6211) );
  OAI211_X1 U7198 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6213), .A(n6212), 
        .B(n6211), .ZN(U3011) );
  NAND2_X1 U7199 ( .A1(n6214), .A2(n6230), .ZN(n6220) );
  AOI222_X1 U7200 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6240), .B1(n6237), .B2(
        n6216), .C1(n6242), .C2(n6215), .ZN(n6217) );
  OAI221_X1 U7201 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6220), .C1(n6219), .C2(n6218), .A(n6217), .ZN(U3012) );
  INV_X1 U7202 ( .A(n6221), .ZN(n6222) );
  AOI222_X1 U7203 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6240), .B1(n6237), .B2(
        n6223), .C1(n6242), .C2(n6222), .ZN(n6226) );
  OAI211_X1 U7204 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6224), .B(n6230), .ZN(n6225) );
  OAI211_X1 U7205 ( .C1(n6234), .C2(n6227), .A(n6226), .B(n6225), .ZN(U3014)
         );
  AOI22_X1 U7206 ( .A1(n6237), .A2(n6228), .B1(n6240), .B2(REIP_REG_3__SCAN_IN), .ZN(n6232) );
  AOI22_X1 U7207 ( .A1(n6230), .A2(n6233), .B1(n6229), .B2(n6242), .ZN(n6231)
         );
  OAI211_X1 U7208 ( .C1(n6234), .C2(n6233), .A(n6232), .B(n6231), .ZN(U3015)
         );
  AOI22_X1 U7209 ( .A1(n6238), .A2(n6237), .B1(n6236), .B2(n6235), .ZN(n6248)
         );
  AOI21_X1 U7210 ( .B1(REIP_REG_2__SCAN_IN), .B2(n6240), .A(n6239), .ZN(n6247)
         );
  AOI22_X1 U7211 ( .A1(n6243), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6242), 
        .B2(n6241), .ZN(n6246) );
  NAND3_X1 U7212 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6244), .A3(n6643), 
        .ZN(n6245) );
  NAND4_X1 U7213 ( .A1(n6248), .A2(n6247), .A3(n6246), .A4(n6245), .ZN(U3016)
         );
  NOR2_X1 U7214 ( .A1(n6614), .A2(n6249), .ZN(U3019) );
  OR2_X1 U7215 ( .A1(n2961), .A2(n6252), .ZN(n6300) );
  NAND3_X1 U7216 ( .A1(n6254), .A2(n6253), .A3(n6263), .ZN(n6255) );
  OAI21_X1 U7217 ( .B1(n6300), .B2(n6297), .A(n6255), .ZN(n6289) );
  NAND2_X1 U7218 ( .A1(n6388), .A2(n6311), .ZN(n6260) );
  INV_X1 U7219 ( .A(n6260), .ZN(n6288) );
  AOI22_X1 U7220 ( .A1(n6256), .A2(n6289), .B1(n6304), .B2(n6288), .ZN(n6265)
         );
  OAI21_X1 U7221 ( .B1(n6346), .B2(n6291), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6257) );
  NAND3_X1 U7222 ( .A1(n6257), .A2(n6310), .A3(n6300), .ZN(n6262) );
  AOI211_X1 U7223 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6260), .A(n6259), .B(
        n6258), .ZN(n6261) );
  NAND3_X1 U7224 ( .A1(n6263), .A2(n6262), .A3(n6261), .ZN(n6292) );
  AOI22_X1 U7225 ( .A1(n6292), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6312), 
        .B2(n6291), .ZN(n6264) );
  OAI211_X1 U7226 ( .C1(n6266), .C2(n6295), .A(n6265), .B(n6264), .ZN(U3068)
         );
  AOI22_X1 U7227 ( .A1(n6359), .A2(n6289), .B1(n6358), .B2(n6288), .ZN(n6268)
         );
  AOI22_X1 U7228 ( .A1(n6292), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6316), 
        .B2(n6291), .ZN(n6267) );
  OAI211_X1 U7229 ( .C1(n6269), .C2(n6295), .A(n6268), .B(n6267), .ZN(U3069)
         );
  AOI22_X1 U7230 ( .A1(n6270), .A2(n6289), .B1(n6321), .B2(n6288), .ZN(n6272)
         );
  AOI22_X1 U7231 ( .A1(n6292), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6320), 
        .B2(n6291), .ZN(n6271) );
  OAI211_X1 U7232 ( .C1(n6273), .C2(n6295), .A(n6272), .B(n6271), .ZN(U3070)
         );
  AOI22_X1 U7233 ( .A1(n6365), .A2(n6289), .B1(n6364), .B2(n6288), .ZN(n6275)
         );
  AOI22_X1 U7234 ( .A1(n6292), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6326), 
        .B2(n6291), .ZN(n6274) );
  OAI211_X1 U7235 ( .C1(n6276), .C2(n6295), .A(n6275), .B(n6274), .ZN(U3071)
         );
  AOI22_X1 U7236 ( .A1(n6277), .A2(n6289), .B1(n6331), .B2(n6288), .ZN(n6279)
         );
  AOI22_X1 U7237 ( .A1(n6292), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6330), 
        .B2(n6291), .ZN(n6278) );
  OAI211_X1 U7238 ( .C1(n6280), .C2(n6295), .A(n6279), .B(n6278), .ZN(U3072)
         );
  AOI22_X1 U7239 ( .A1(n6374), .A2(n6289), .B1(n6372), .B2(n6288), .ZN(n6282)
         );
  AOI22_X1 U7240 ( .A1(n6292), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6336), 
        .B2(n6291), .ZN(n6281) );
  OAI211_X1 U7241 ( .C1(n6283), .C2(n6295), .A(n6282), .B(n6281), .ZN(U3073)
         );
  AOI22_X1 U7242 ( .A1(n6284), .A2(n6289), .B1(n6341), .B2(n6288), .ZN(n6286)
         );
  AOI22_X1 U7243 ( .A1(n6292), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6340), 
        .B2(n6291), .ZN(n6285) );
  OAI211_X1 U7244 ( .C1(n6287), .C2(n6295), .A(n6286), .B(n6285), .ZN(U3074)
         );
  AOI22_X1 U7245 ( .A1(n6290), .A2(n6289), .B1(n6349), .B2(n6288), .ZN(n6294)
         );
  AOI22_X1 U7246 ( .A1(n6292), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6347), 
        .B2(n6291), .ZN(n6293) );
  OAI211_X1 U7247 ( .C1(n6296), .C2(n6295), .A(n6294), .B(n6293), .ZN(U3075)
         );
  NOR2_X1 U7248 ( .A1(n6298), .A2(n6297), .ZN(n6307) );
  OAI21_X1 U7249 ( .B1(n6300), .B2(n6299), .A(n6301), .ZN(n6305) );
  AOI22_X1 U7250 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6311), .B1(n6307), .B2(
        n6305), .ZN(n6356) );
  INV_X1 U7251 ( .A(n6301), .ZN(n6348) );
  AOI22_X1 U7252 ( .A1(n6304), .A2(n6348), .B1(n6303), .B2(n6350), .ZN(n6314)
         );
  INV_X1 U7253 ( .A(n6305), .ZN(n6306) );
  NAND2_X1 U7254 ( .A1(n6307), .A2(n6306), .ZN(n6308) );
  OAI211_X1 U7255 ( .C1(n6311), .C2(n6310), .A(n6309), .B(n6308), .ZN(n6352)
         );
  AOI22_X1 U7256 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6352), .B1(n6312), 
        .B2(n6346), .ZN(n6313) );
  OAI211_X1 U7257 ( .C1(n6356), .C2(n6315), .A(n6314), .B(n6313), .ZN(U3076)
         );
  AOI22_X1 U7258 ( .A1(n6358), .A2(n6348), .B1(n6316), .B2(n6346), .ZN(n6318)
         );
  AOI22_X1 U7259 ( .A1(n6352), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n6357), 
        .B2(n6350), .ZN(n6317) );
  OAI211_X1 U7260 ( .C1(n6356), .C2(n6319), .A(n6318), .B(n6317), .ZN(U3077)
         );
  AOI22_X1 U7261 ( .A1(n6321), .A2(n6348), .B1(n6320), .B2(n6346), .ZN(n6324)
         );
  AOI22_X1 U7262 ( .A1(n6352), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n6322), 
        .B2(n6350), .ZN(n6323) );
  OAI211_X1 U7263 ( .C1(n6356), .C2(n6325), .A(n6324), .B(n6323), .ZN(U3078)
         );
  AOI22_X1 U7264 ( .A1(n6364), .A2(n6348), .B1(n6363), .B2(n6350), .ZN(n6328)
         );
  AOI22_X1 U7265 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6352), .B1(n6326), 
        .B2(n6346), .ZN(n6327) );
  OAI211_X1 U7266 ( .C1(n6356), .C2(n6329), .A(n6328), .B(n6327), .ZN(U3079)
         );
  AOI22_X1 U7267 ( .A1(n6331), .A2(n6348), .B1(n6330), .B2(n6346), .ZN(n6334)
         );
  AOI22_X1 U7268 ( .A1(n6352), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n6332), 
        .B2(n6350), .ZN(n6333) );
  OAI211_X1 U7269 ( .C1(n6356), .C2(n6335), .A(n6334), .B(n6333), .ZN(U3080)
         );
  AOI22_X1 U7270 ( .A1(n6372), .A2(n6348), .B1(n6336), .B2(n6346), .ZN(n6338)
         );
  AOI22_X1 U7271 ( .A1(n6352), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n6370), 
        .B2(n6350), .ZN(n6337) );
  OAI211_X1 U7272 ( .C1(n6356), .C2(n6339), .A(n6338), .B(n6337), .ZN(U3081)
         );
  AOI22_X1 U7273 ( .A1(n6341), .A2(n6348), .B1(n6340), .B2(n6346), .ZN(n6344)
         );
  AOI22_X1 U7274 ( .A1(n6352), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n6342), 
        .B2(n6350), .ZN(n6343) );
  OAI211_X1 U7275 ( .C1(n6356), .C2(n6345), .A(n6344), .B(n6343), .ZN(U3082)
         );
  AOI22_X1 U7276 ( .A1(n6349), .A2(n6348), .B1(n6347), .B2(n6346), .ZN(n6354)
         );
  AOI22_X1 U7277 ( .A1(n6352), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n6351), 
        .B2(n6350), .ZN(n6353) );
  OAI211_X1 U7278 ( .C1(n6356), .C2(n6355), .A(n6354), .B(n6353), .ZN(U3083)
         );
  AOI22_X1 U7279 ( .A1(n6358), .A2(n6371), .B1(n6357), .B2(n6369), .ZN(n6361)
         );
  AOI22_X1 U7280 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6375), .B1(n6359), 
        .B2(n6373), .ZN(n6360) );
  OAI211_X1 U7281 ( .C1(n6362), .C2(n6378), .A(n6361), .B(n6360), .ZN(U3109)
         );
  AOI22_X1 U7282 ( .A1(n6364), .A2(n6371), .B1(n6363), .B2(n6369), .ZN(n6367)
         );
  AOI22_X1 U7283 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6375), .B1(n6365), 
        .B2(n6373), .ZN(n6366) );
  OAI211_X1 U7284 ( .C1(n6368), .C2(n6378), .A(n6367), .B(n6366), .ZN(U3111)
         );
  AOI22_X1 U7285 ( .A1(n6372), .A2(n6371), .B1(n6370), .B2(n6369), .ZN(n6377)
         );
  AOI22_X1 U7286 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6375), .B1(n6374), 
        .B2(n6373), .ZN(n6376) );
  OAI211_X1 U7287 ( .C1(n6379), .C2(n6378), .A(n6377), .B(n6376), .ZN(U3113)
         );
  NOR2_X1 U7288 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6383) );
  OAI211_X1 U7289 ( .C1(n6383), .C2(n6382), .A(n6381), .B(n6380), .ZN(n6384)
         );
  NOR2_X1 U7290 ( .A1(n6385), .A2(n6384), .ZN(n6404) );
  NAND2_X1 U7291 ( .A1(n6387), .A2(n6386), .ZN(n6392) );
  INV_X1 U7292 ( .A(n6392), .ZN(n6395) );
  AOI21_X1 U7293 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6389), .A(n6388), 
        .ZN(n6390) );
  OAI211_X1 U7294 ( .C1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n6392), .A(n6391), .B(n6390), .ZN(n6393) );
  OAI21_X1 U7295 ( .B1(n6395), .B2(n6394), .A(n6393), .ZN(n6396) );
  AOI222_X1 U7296 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6397), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6396), .C1(n6397), .C2(n6396), 
        .ZN(n6398) );
  INV_X1 U7297 ( .A(n6398), .ZN(n6399) );
  AND2_X1 U7298 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6399), .ZN(n6400)
         );
  OAI22_X1 U7299 ( .A1(n6401), .A2(n6400), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6399), .ZN(n6402) );
  NAND2_X1 U7300 ( .A1(n6402), .A2(n6614), .ZN(n6403) );
  NAND2_X1 U7301 ( .A1(n6419), .A2(n6422), .ZN(n6406) );
  NAND2_X1 U7302 ( .A1(READY_N), .A2(n6521), .ZN(n6405) );
  NAND2_X1 U7303 ( .A1(n6406), .A2(n6405), .ZN(n6412) );
  AND2_X1 U7304 ( .A1(n6408), .A2(n6407), .ZN(n6409) );
  NAND2_X1 U7305 ( .A1(n6410), .A2(n6409), .ZN(n6411) );
  OAI21_X1 U7306 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6520), .A(n6507), .ZN(
        n6426) );
  AOI221_X1 U7307 ( .B1(n6414), .B2(STATE2_REG_0__SCAN_IN), .C1(n6426), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6413), .ZN(n6417) );
  OAI211_X1 U7308 ( .C1(n6430), .C2(n6415), .A(n6421), .B(n6507), .ZN(n6416)
         );
  OAI211_X1 U7309 ( .C1(n6419), .C2(n6418), .A(n6417), .B(n6416), .ZN(U3148)
         );
  NOR2_X1 U7310 ( .A1(n6421), .A2(n6420), .ZN(n6423) );
  AOI21_X1 U7311 ( .B1(n6423), .B2(n6520), .A(n6422), .ZN(n6428) );
  INV_X1 U7312 ( .A(n6425), .ZN(n6433) );
  OAI221_X1 U7313 ( .B1(n6433), .B2(n6426), .C1(n6425), .C2(n6424), .A(
        STATE2_REG_1__SCAN_IN), .ZN(n6427) );
  OAI21_X1 U7314 ( .B1(n6429), .B2(n6428), .A(n6427), .ZN(U3149) );
  OAI211_X1 U7315 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6520), .A(n6506), .B(
        n6430), .ZN(n6432) );
  OAI21_X1 U7316 ( .B1(n6433), .B2(n6432), .A(n6431), .ZN(U3150) );
  AND2_X1 U7317 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6688), .ZN(U3151) );
  AND2_X1 U7318 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6688), .ZN(U3152) );
  AND2_X1 U7319 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6688), .ZN(U3153) );
  AND2_X1 U7320 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6688), .ZN(U3154) );
  AND2_X1 U7321 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6688), .ZN(U3155) );
  AND2_X1 U7322 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6688), .ZN(U3156) );
  AND2_X1 U7323 ( .A1(n6688), .A2(DATAWIDTH_REG_25__SCAN_IN), .ZN(U3157) );
  AND2_X1 U7324 ( .A1(n6688), .A2(DATAWIDTH_REG_24__SCAN_IN), .ZN(U3158) );
  AND2_X1 U7325 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6688), .ZN(U3159) );
  AND2_X1 U7326 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6688), .ZN(U3160) );
  AND2_X1 U7327 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6688), .ZN(U3161) );
  AND2_X1 U7328 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6688), .ZN(U3162) );
  AND2_X1 U7329 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6688), .ZN(U3163) );
  AND2_X1 U7330 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6688), .ZN(U3164) );
  AND2_X1 U7331 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6688), .ZN(U3165) );
  AND2_X1 U7332 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6688), .ZN(U3166) );
  AND2_X1 U7333 ( .A1(n6688), .A2(DATAWIDTH_REG_15__SCAN_IN), .ZN(U3167) );
  AND2_X1 U7334 ( .A1(n6688), .A2(DATAWIDTH_REG_14__SCAN_IN), .ZN(U3168) );
  AND2_X1 U7335 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6688), .ZN(U3169) );
  AND2_X1 U7336 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6688), .ZN(U3170) );
  INV_X1 U7337 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6584) );
  NOR2_X1 U7338 ( .A1(n6505), .A2(n6584), .ZN(U3171) );
  AND2_X1 U7339 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6688), .ZN(U3172) );
  AND2_X1 U7340 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6688), .ZN(U3173) );
  AND2_X1 U7341 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6688), .ZN(U3174) );
  AND2_X1 U7342 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6688), .ZN(U3175) );
  AND2_X1 U7343 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6688), .ZN(U3176) );
  AND2_X1 U7344 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6688), .ZN(U3177) );
  AND2_X1 U7345 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6688), .ZN(U3178) );
  AND2_X1 U7346 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6688), .ZN(U3179) );
  INV_X1 U7347 ( .A(n6434), .ZN(n6442) );
  AOI22_X1 U7348 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6450) );
  AND2_X1 U7349 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6438) );
  INV_X1 U7350 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6436) );
  INV_X1 U7351 ( .A(NA_N), .ZN(n6443) );
  AOI221_X1 U7352 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6443), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6447) );
  AOI221_X1 U7353 ( .B1(n6438), .B2(n6529), .C1(n6436), .C2(n6529), .A(n6447), 
        .ZN(n6435) );
  OAI21_X1 U7354 ( .B1(n6442), .B2(n6450), .A(n6435), .ZN(U3181) );
  INV_X1 U7355 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6445) );
  NOR2_X1 U7356 ( .A1(n6445), .A2(n6436), .ZN(n6444) );
  NAND2_X1 U7357 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6437) );
  OAI21_X1 U7358 ( .B1(n6444), .B2(n6438), .A(n6437), .ZN(n6439) );
  OAI211_X1 U7359 ( .C1(n6441), .C2(n6520), .A(n6440), .B(n6439), .ZN(U3182)
         );
  AOI21_X1 U7360 ( .B1(n6444), .B2(n6443), .A(n6442), .ZN(n6449) );
  AOI221_X1 U7361 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6520), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6446) );
  AOI221_X1 U7362 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6446), .C2(HOLD), .A(n6445), .ZN(n6448) );
  OAI22_X1 U7363 ( .A1(n6450), .A2(n6449), .B1(n6448), .B2(n6447), .ZN(U3183)
         );
  NAND2_X1 U7364 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6500), .ZN(n6497) );
  NOR2_X2 U7365 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6529), .ZN(n6495) );
  AOI22_X1 U7366 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6495), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6529), .ZN(n6451) );
  OAI21_X1 U7367 ( .B1(n6509), .B2(n6497), .A(n6451), .ZN(U3184) );
  INV_X1 U7368 ( .A(n6497), .ZN(n6492) );
  AOI22_X1 U7369 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6529), .ZN(n6452) );
  OAI21_X1 U7370 ( .B1(n6453), .B2(n6494), .A(n6452), .ZN(U3185) );
  AOI22_X1 U7371 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6529), .ZN(n6454) );
  OAI21_X1 U7372 ( .B1(n6456), .B2(n6494), .A(n6454), .ZN(U3186) );
  AOI22_X1 U7373 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6495), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6529), .ZN(n6455) );
  OAI21_X1 U7374 ( .B1(n6456), .B2(n6497), .A(n6455), .ZN(U3187) );
  AOI22_X1 U7375 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6529), .ZN(n6457) );
  OAI21_X1 U7376 ( .B1(n6459), .B2(n6494), .A(n6457), .ZN(U3188) );
  AOI22_X1 U7377 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6495), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6529), .ZN(n6458) );
  OAI21_X1 U7378 ( .B1(n6459), .B2(n6497), .A(n6458), .ZN(U3189) );
  AOI22_X1 U7379 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6529), .ZN(n6460) );
  OAI21_X1 U7380 ( .B1(n6462), .B2(n6494), .A(n6460), .ZN(U3190) );
  AOI22_X1 U7381 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6495), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6529), .ZN(n6461) );
  OAI21_X1 U7382 ( .B1(n6462), .B2(n6497), .A(n6461), .ZN(U3191) );
  AOI22_X1 U7383 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6529), .ZN(n6463) );
  OAI21_X1 U7384 ( .B1(n6465), .B2(n6494), .A(n6463), .ZN(U3192) );
  AOI22_X1 U7385 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6495), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6529), .ZN(n6464) );
  OAI21_X1 U7386 ( .B1(n6465), .B2(n6497), .A(n6464), .ZN(U3193) );
  AOI22_X1 U7387 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6529), .ZN(n6466) );
  OAI21_X1 U7388 ( .B1(n6468), .B2(n6494), .A(n6466), .ZN(U3194) );
  AOI22_X1 U7389 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6495), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6529), .ZN(n6467) );
  OAI21_X1 U7390 ( .B1(n6468), .B2(n6497), .A(n6467), .ZN(U3195) );
  AOI22_X1 U7391 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6529), .ZN(n6469) );
  OAI21_X1 U7392 ( .B1(n6471), .B2(n6494), .A(n6469), .ZN(U3196) );
  AOI22_X1 U7393 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6495), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6529), .ZN(n6470) );
  OAI21_X1 U7394 ( .B1(n6471), .B2(n6497), .A(n6470), .ZN(U3197) );
  AOI22_X1 U7395 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6529), .ZN(n6472) );
  OAI21_X1 U7396 ( .B1(n6474), .B2(n6494), .A(n6472), .ZN(U3198) );
  AOI22_X1 U7397 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6495), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6529), .ZN(n6473) );
  OAI21_X1 U7398 ( .B1(n6474), .B2(n6497), .A(n6473), .ZN(U3199) );
  AOI22_X1 U7399 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6529), .ZN(n6475) );
  OAI21_X1 U7400 ( .B1(n5692), .B2(n6494), .A(n6475), .ZN(U3200) );
  AOI22_X1 U7401 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6529), .ZN(n6476) );
  OAI21_X1 U7402 ( .B1(n6574), .B2(n6494), .A(n6476), .ZN(U3201) );
  AOI22_X1 U7403 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6529), .ZN(n6477) );
  OAI21_X1 U7404 ( .B1(n6479), .B2(n6494), .A(n6477), .ZN(U3202) );
  AOI22_X1 U7405 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6495), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6529), .ZN(n6478) );
  OAI21_X1 U7406 ( .B1(n6479), .B2(n6497), .A(n6478), .ZN(U3203) );
  AOI22_X1 U7407 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6495), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6529), .ZN(n6480) );
  OAI21_X1 U7408 ( .B1(n6481), .B2(n6497), .A(n6480), .ZN(U3204) );
  AOI22_X1 U7409 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6495), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6529), .ZN(n6482) );
  OAI21_X1 U7410 ( .B1(n6483), .B2(n6497), .A(n6482), .ZN(U3205) );
  AOI222_X1 U7411 ( .A1(n6492), .A2(REIP_REG_23__SCAN_IN), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6529), .C1(REIP_REG_24__SCAN_IN), .C2(
        n6495), .ZN(n6484) );
  INV_X1 U7412 ( .A(n6484), .ZN(U3206) );
  AOI22_X1 U7413 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6529), .ZN(n6485) );
  OAI21_X1 U7414 ( .B1(n6571), .B2(n6494), .A(n6485), .ZN(U3207) );
  AOI22_X1 U7415 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6495), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6529), .ZN(n6486) );
  OAI21_X1 U7416 ( .B1(n6571), .B2(n6497), .A(n6486), .ZN(U3208) );
  AOI22_X1 U7417 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6529), .ZN(n6487) );
  OAI21_X1 U7418 ( .B1(n6489), .B2(n6494), .A(n6487), .ZN(U3209) );
  AOI22_X1 U7419 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6495), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6529), .ZN(n6488) );
  OAI21_X1 U7420 ( .B1(n6489), .B2(n6497), .A(n6488), .ZN(U3210) );
  AOI22_X1 U7421 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6495), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6529), .ZN(n6490) );
  OAI21_X1 U7422 ( .B1(n6491), .B2(n6497), .A(n6490), .ZN(U3211) );
  AOI22_X1 U7423 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6492), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6529), .ZN(n6493) );
  OAI21_X1 U7424 ( .B1(n6498), .B2(n6494), .A(n6493), .ZN(U3212) );
  AOI22_X1 U7425 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6495), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6529), .ZN(n6496) );
  OAI21_X1 U7426 ( .B1(n6498), .B2(n6497), .A(n6496), .ZN(U3213) );
  OAI22_X1 U7427 ( .A1(n6529), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6500), .ZN(n6499) );
  INV_X1 U7428 ( .A(n6499), .ZN(U3445) );
  MUX2_X1 U7429 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6529), .Z(U3446) );
  MUX2_X1 U7430 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6529), .Z(U3447) );
  OAI22_X1 U7431 ( .A1(n6529), .A2(BYTEENABLE_REG_0__SCAN_IN), .B1(
        BE_N_REG_0__SCAN_IN), .B2(n6500), .ZN(n6501) );
  INV_X1 U7432 ( .A(n6501), .ZN(U3448) );
  OAI21_X1 U7433 ( .B1(n6505), .B2(DATAWIDTH_REG_0__SCAN_IN), .A(n6503), .ZN(
        n6502) );
  INV_X1 U7434 ( .A(n6502), .ZN(U3451) );
  OAI21_X1 U7435 ( .B1(n6505), .B2(n6504), .A(n6503), .ZN(U3452) );
  OAI221_X1 U7436 ( .B1(n6508), .B2(STATE2_REG_0__SCAN_IN), .C1(n6508), .C2(
        n6507), .A(n6506), .ZN(U3453) );
  AOI21_X1 U7437 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6510) );
  AOI22_X1 U7438 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6510), .B2(n6509), .ZN(n6513) );
  INV_X1 U7439 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6512) );
  AOI22_X1 U7440 ( .A1(n6516), .A2(n6513), .B1(n6512), .B2(n6511), .ZN(U3468)
         );
  INV_X1 U7441 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6515) );
  OAI21_X1 U7442 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6516), .ZN(n6514) );
  OAI21_X1 U7443 ( .B1(n6516), .B2(n6515), .A(n6514), .ZN(U3469) );
  NAND2_X1 U7444 ( .A1(n6529), .A2(W_R_N_REG_SCAN_IN), .ZN(n6517) );
  OAI21_X1 U7445 ( .B1(n6529), .B2(READREQUEST_REG_SCAN_IN), .A(n6517), .ZN(
        U3470) );
  AOI211_X1 U7446 ( .C1(n6521), .C2(n6520), .A(n6519), .B(n6518), .ZN(n6528)
         );
  OAI211_X1 U7447 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6523), .A(n6522), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6525) );
  AOI21_X1 U7448 ( .B1(n6525), .B2(STATE2_REG_0__SCAN_IN), .A(n6524), .ZN(
        n6527) );
  NAND2_X1 U7449 ( .A1(n6528), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6526) );
  OAI21_X1 U7450 ( .B1(n6528), .B2(n6527), .A(n6526), .ZN(U3472) );
  MUX2_X1 U7451 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6529), .Z(U3473) );
  AOI22_X1 U7452 ( .A1(n6531), .A2(keyinput12), .B1(n4703), .B2(keyinput25), 
        .ZN(n6530) );
  OAI221_X1 U7453 ( .B1(n6531), .B2(keyinput12), .C1(n4703), .C2(keyinput25), 
        .A(n6530), .ZN(n6544) );
  INV_X1 U7454 ( .A(keyinput4), .ZN(n6534) );
  INV_X1 U7455 ( .A(keyinput41), .ZN(n6533) );
  AOI22_X1 U7456 ( .A1(n6534), .A2(ADDRESS_REG_16__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6533), .ZN(n6532) );
  OAI221_X1 U7457 ( .B1(n6534), .B2(ADDRESS_REG_16__SCAN_IN), .C1(n6533), .C2(
        BE_N_REG_3__SCAN_IN), .A(n6532), .ZN(n6543) );
  AOI22_X1 U7458 ( .A1(n6537), .A2(keyinput15), .B1(keyinput50), .B2(n6536), 
        .ZN(n6535) );
  OAI221_X1 U7459 ( .B1(n6537), .B2(keyinput15), .C1(n6536), .C2(keyinput50), 
        .A(n6535), .ZN(n6542) );
  INV_X1 U7460 ( .A(keyinput35), .ZN(n6540) );
  INV_X1 U7461 ( .A(keyinput20), .ZN(n6539) );
  AOI22_X1 U7462 ( .A1(n6540), .A2(M_IO_N_REG_SCAN_IN), .B1(
        BE_N_REG_0__SCAN_IN), .B2(n6539), .ZN(n6538) );
  OAI221_X1 U7463 ( .B1(n6540), .B2(M_IO_N_REG_SCAN_IN), .C1(n6539), .C2(
        BE_N_REG_0__SCAN_IN), .A(n6538), .ZN(n6541) );
  NOR4_X1 U7464 ( .A1(n6544), .A2(n6543), .A3(n6542), .A4(n6541), .ZN(n6687)
         );
  INV_X1 U7465 ( .A(DATAI_18_), .ZN(n6547) );
  INV_X1 U7466 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n6546) );
  AOI22_X1 U7467 ( .A1(n6547), .A2(keyinput52), .B1(keyinput6), .B2(n6546), 
        .ZN(n6545) );
  OAI221_X1 U7468 ( .B1(n6547), .B2(keyinput52), .C1(n6546), .C2(keyinput6), 
        .A(n6545), .ZN(n6559) );
  AOI22_X1 U7469 ( .A1(n6549), .A2(keyinput3), .B1(keyinput9), .B2(n3652), 
        .ZN(n6548) );
  OAI221_X1 U7470 ( .B1(n6549), .B2(keyinput3), .C1(n3652), .C2(keyinput9), 
        .A(n6548), .ZN(n6558) );
  INV_X1 U7471 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n6552) );
  INV_X1 U7472 ( .A(keyinput61), .ZN(n6551) );
  AOI22_X1 U7473 ( .A1(n6552), .A2(keyinput33), .B1(DATAO_REG_31__SCAN_IN), 
        .B2(n6551), .ZN(n6550) );
  OAI221_X1 U7474 ( .B1(n6552), .B2(keyinput33), .C1(n6551), .C2(
        DATAO_REG_31__SCAN_IN), .A(n6550), .ZN(n6557) );
  INV_X1 U7475 ( .A(keyinput40), .ZN(n6553) );
  XOR2_X1 U7476 ( .A(DATAWIDTH_REG_24__SCAN_IN), .B(n6553), .Z(n6555) );
  XNOR2_X1 U7477 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .B(keyinput19), .ZN(n6554)
         );
  NAND2_X1 U7478 ( .A1(n6555), .A2(n6554), .ZN(n6556) );
  NOR4_X1 U7479 ( .A1(n6559), .A2(n6558), .A3(n6557), .A4(n6556), .ZN(n6686)
         );
  INV_X1 U7480 ( .A(keyinput31), .ZN(n6561) );
  AOI22_X1 U7481 ( .A1(n6562), .A2(keyinput62), .B1(DATAWIDTH_REG_15__SCAN_IN), 
        .B2(n6561), .ZN(n6560) );
  OAI221_X1 U7482 ( .B1(n6562), .B2(keyinput62), .C1(n6561), .C2(
        DATAWIDTH_REG_15__SCAN_IN), .A(n6560), .ZN(n6656) );
  INV_X1 U7483 ( .A(keyinput51), .ZN(n6564) );
  AOI22_X1 U7484 ( .A1(n6565), .A2(keyinput58), .B1(DATAO_REG_22__SCAN_IN), 
        .B2(n6564), .ZN(n6563) );
  OAI221_X1 U7485 ( .B1(n6565), .B2(keyinput58), .C1(n6564), .C2(
        DATAO_REG_22__SCAN_IN), .A(n6563), .ZN(n6655) );
  INV_X1 U7486 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n6568) );
  INV_X1 U7487 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6567) );
  AOI22_X1 U7488 ( .A1(n6568), .A2(keyinput39), .B1(n6567), .B2(keyinput14), 
        .ZN(n6566) );
  OAI221_X1 U7489 ( .B1(n6568), .B2(keyinput39), .C1(n6567), .C2(keyinput14), 
        .A(n6566), .ZN(n6581) );
  AOI22_X1 U7490 ( .A1(n6571), .A2(keyinput55), .B1(n6570), .B2(keyinput54), 
        .ZN(n6569) );
  OAI221_X1 U7491 ( .B1(n6571), .B2(keyinput55), .C1(n6570), .C2(keyinput54), 
        .A(n6569), .ZN(n6580) );
  INV_X1 U7492 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n6573) );
  AOI22_X1 U7493 ( .A1(n6574), .A2(keyinput23), .B1(n6573), .B2(keyinput21), 
        .ZN(n6572) );
  OAI221_X1 U7494 ( .B1(n6574), .B2(keyinput23), .C1(n6573), .C2(keyinput21), 
        .A(n6572), .ZN(n6579) );
  AOI22_X1 U7495 ( .A1(n6577), .A2(keyinput1), .B1(n6576), .B2(keyinput45), 
        .ZN(n6575) );
  OAI221_X1 U7496 ( .B1(n6577), .B2(keyinput1), .C1(n6576), .C2(keyinput45), 
        .A(n6575), .ZN(n6578) );
  NOR4_X1 U7497 ( .A1(n6581), .A2(n6580), .A3(n6579), .A4(n6578), .ZN(n6588)
         );
  INV_X1 U7498 ( .A(keyinput43), .ZN(n6583) );
  OAI22_X1 U7499 ( .A1(keyinput5), .A2(n6584), .B1(n6583), .B2(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n6582) );
  AOI221_X1 U7500 ( .B1(n6584), .B2(keyinput5), .C1(n6583), .C2(
        DATAWIDTH_REG_25__SCAN_IN), .A(n6582), .ZN(n6587) );
  XNOR2_X1 U7501 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .B(keyinput0), .ZN(n6586)
         );
  XNOR2_X1 U7502 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .B(keyinput47), .ZN(n6585) );
  NAND4_X1 U7503 ( .A1(n6588), .A2(n6587), .A3(n6586), .A4(n6585), .ZN(n6654)
         );
  INV_X1 U7504 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n6590) );
  AOI22_X1 U7505 ( .A1(n6591), .A2(keyinput7), .B1(keyinput60), .B2(n6590), 
        .ZN(n6589) );
  OAI221_X1 U7506 ( .B1(n6591), .B2(keyinput7), .C1(n6590), .C2(keyinput60), 
        .A(n6589), .ZN(n6603) );
  INV_X1 U7507 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n6593) );
  AOI22_X1 U7508 ( .A1(n4579), .A2(keyinput36), .B1(n6593), .B2(keyinput26), 
        .ZN(n6592) );
  OAI221_X1 U7509 ( .B1(n4579), .B2(keyinput36), .C1(n6593), .C2(keyinput26), 
        .A(n6592), .ZN(n6602) );
  INV_X1 U7510 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6596) );
  INV_X1 U7511 ( .A(keyinput8), .ZN(n6595) );
  AOI22_X1 U7512 ( .A1(n6596), .A2(keyinput63), .B1(ADDRESS_REG_22__SCAN_IN), 
        .B2(n6595), .ZN(n6594) );
  OAI221_X1 U7513 ( .B1(n6596), .B2(keyinput63), .C1(n6595), .C2(
        ADDRESS_REG_22__SCAN_IN), .A(n6594), .ZN(n6601) );
  AOI22_X1 U7514 ( .A1(n6599), .A2(keyinput38), .B1(keyinput30), .B2(n6598), 
        .ZN(n6597) );
  OAI221_X1 U7515 ( .B1(n6599), .B2(keyinput38), .C1(n6598), .C2(keyinput30), 
        .A(n6597), .ZN(n6600) );
  NOR4_X1 U7516 ( .A1(n6603), .A2(n6602), .A3(n6601), .A4(n6600), .ZN(n6652)
         );
  INV_X1 U7517 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n6605) );
  AOI22_X1 U7518 ( .A1(n5558), .A2(keyinput59), .B1(n6605), .B2(keyinput42), 
        .ZN(n6604) );
  OAI221_X1 U7519 ( .B1(n5558), .B2(keyinput59), .C1(n6605), .C2(keyinput42), 
        .A(n6604), .ZN(n6618) );
  INV_X1 U7520 ( .A(keyinput16), .ZN(n6607) );
  AOI22_X1 U7521 ( .A1(n6608), .A2(keyinput29), .B1(DATAWIDTH_REG_14__SCAN_IN), 
        .B2(n6607), .ZN(n6606) );
  OAI221_X1 U7522 ( .B1(n6608), .B2(keyinput29), .C1(n6607), .C2(
        DATAWIDTH_REG_14__SCAN_IN), .A(n6606), .ZN(n6617) );
  INV_X1 U7523 ( .A(DATAI_23_), .ZN(n6611) );
  INV_X1 U7524 ( .A(DATAI_31_), .ZN(n6610) );
  AOI22_X1 U7525 ( .A1(n6611), .A2(keyinput2), .B1(n6610), .B2(keyinput37), 
        .ZN(n6609) );
  OAI221_X1 U7526 ( .B1(n6611), .B2(keyinput2), .C1(n6610), .C2(keyinput37), 
        .A(n6609), .ZN(n6616) );
  INV_X1 U7527 ( .A(keyinput18), .ZN(n6613) );
  AOI22_X1 U7528 ( .A1(n6614), .A2(keyinput17), .B1(ADDRESS_REG_4__SCAN_IN), 
        .B2(n6613), .ZN(n6612) );
  OAI221_X1 U7529 ( .B1(n6614), .B2(keyinput17), .C1(n6613), .C2(
        ADDRESS_REG_4__SCAN_IN), .A(n6612), .ZN(n6615) );
  NOR4_X1 U7530 ( .A1(n6618), .A2(n6617), .A3(n6616), .A4(n6615), .ZN(n6651)
         );
  INV_X1 U7531 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n6621) );
  INV_X1 U7532 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6620) );
  AOI22_X1 U7533 ( .A1(n6621), .A2(keyinput53), .B1(n6620), .B2(keyinput57), 
        .ZN(n6619) );
  OAI221_X1 U7534 ( .B1(n6621), .B2(keyinput53), .C1(n6620), .C2(keyinput57), 
        .A(n6619), .ZN(n6633) );
  AOI22_X1 U7535 ( .A1(n3620), .A2(keyinput28), .B1(keyinput10), .B2(n6623), 
        .ZN(n6622) );
  OAI221_X1 U7536 ( .B1(n3620), .B2(keyinput28), .C1(n6623), .C2(keyinput10), 
        .A(n6622), .ZN(n6632) );
  INV_X1 U7537 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n6625) );
  AOI22_X1 U7538 ( .A1(n6626), .A2(keyinput11), .B1(n6625), .B2(keyinput56), 
        .ZN(n6624) );
  OAI221_X1 U7539 ( .B1(n6626), .B2(keyinput11), .C1(n6625), .C2(keyinput56), 
        .A(n6624), .ZN(n6631) );
  INV_X1 U7540 ( .A(DATAI_9_), .ZN(n6629) );
  AOI22_X1 U7541 ( .A1(n6629), .A2(keyinput22), .B1(n6628), .B2(keyinput34), 
        .ZN(n6627) );
  OAI221_X1 U7542 ( .B1(n6629), .B2(keyinput22), .C1(n6628), .C2(keyinput34), 
        .A(n6627), .ZN(n6630) );
  NOR4_X1 U7543 ( .A1(n6633), .A2(n6632), .A3(n6631), .A4(n6630), .ZN(n6650)
         );
  INV_X1 U7544 ( .A(EAX_REG_31__SCAN_IN), .ZN(n6636) );
  INV_X1 U7545 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n6635) );
  AOI22_X1 U7546 ( .A1(n6636), .A2(keyinput44), .B1(n6635), .B2(keyinput49), 
        .ZN(n6634) );
  OAI221_X1 U7547 ( .B1(n6636), .B2(keyinput44), .C1(n6635), .C2(keyinput49), 
        .A(n6634), .ZN(n6648) );
  AOI22_X1 U7548 ( .A1(n6639), .A2(keyinput13), .B1(keyinput32), .B2(n6638), 
        .ZN(n6637) );
  OAI221_X1 U7549 ( .B1(n6639), .B2(keyinput13), .C1(n6638), .C2(keyinput32), 
        .A(n6637), .ZN(n6647) );
  AOI22_X1 U7550 ( .A1(n6641), .A2(keyinput46), .B1(n4734), .B2(keyinput48), 
        .ZN(n6640) );
  OAI221_X1 U7551 ( .B1(n6641), .B2(keyinput46), .C1(n4734), .C2(keyinput48), 
        .A(n6640), .ZN(n6646) );
  INV_X1 U7552 ( .A(LWORD_REG_8__SCAN_IN), .ZN(n6644) );
  AOI22_X1 U7553 ( .A1(n6644), .A2(keyinput27), .B1(n6643), .B2(keyinput24), 
        .ZN(n6642) );
  OAI221_X1 U7554 ( .B1(n6644), .B2(keyinput27), .C1(n6643), .C2(keyinput24), 
        .A(n6642), .ZN(n6645) );
  NOR4_X1 U7555 ( .A1(n6648), .A2(n6647), .A3(n6646), .A4(n6645), .ZN(n6649)
         );
  NAND4_X1 U7556 ( .A1(n6652), .A2(n6651), .A3(n6650), .A4(n6649), .ZN(n6653)
         );
  NOR4_X1 U7557 ( .A1(n6656), .A2(n6655), .A3(n6654), .A4(n6653), .ZN(n6685)
         );
  NAND4_X1 U7558 ( .A1(keyinput63), .A2(keyinput8), .A3(keyinput38), .A4(
        keyinput30), .ZN(n6661) );
  NAND3_X1 U7559 ( .A1(keyinput59), .A2(keyinput16), .A3(keyinput29), .ZN(
        n6660) );
  NOR3_X1 U7560 ( .A1(keyinput7), .A2(keyinput60), .A3(keyinput26), .ZN(n6658)
         );
  NOR3_X1 U7561 ( .A1(keyinput2), .A2(keyinput37), .A3(keyinput17), .ZN(n6657)
         );
  NAND4_X1 U7562 ( .A1(keyinput36), .A2(n6658), .A3(keyinput18), .A4(n6657), 
        .ZN(n6659) );
  NOR4_X1 U7563 ( .A1(keyinput42), .A2(n6661), .A3(n6660), .A4(n6659), .ZN(
        n6683) );
  NAND2_X1 U7564 ( .A1(keyinput44), .A2(keyinput49), .ZN(n6664) );
  INV_X1 U7565 ( .A(keyinput48), .ZN(n6662) );
  NAND4_X1 U7566 ( .A1(keyinput46), .A2(keyinput27), .A3(keyinput24), .A4(
        n6662), .ZN(n6663) );
  NOR4_X1 U7567 ( .A1(keyinput13), .A2(keyinput32), .A3(n6664), .A4(n6663), 
        .ZN(n6682) );
  NAND3_X1 U7568 ( .A1(keyinput53), .A2(keyinput57), .A3(keyinput28), .ZN(
        n6666) );
  NAND3_X1 U7569 ( .A1(keyinput11), .A2(keyinput56), .A3(keyinput22), .ZN(
        n6665) );
  NOR4_X1 U7570 ( .A1(keyinput10), .A2(keyinput34), .A3(n6666), .A4(n6665), 
        .ZN(n6681) );
  NOR2_X1 U7571 ( .A1(keyinput51), .A2(keyinput62), .ZN(n6672) );
  NAND2_X1 U7572 ( .A1(keyinput55), .A2(keyinput54), .ZN(n6670) );
  NOR3_X1 U7573 ( .A1(keyinput5), .A2(keyinput43), .A3(keyinput0), .ZN(n6668)
         );
  NOR3_X1 U7574 ( .A1(keyinput1), .A2(keyinput23), .A3(keyinput21), .ZN(n6667)
         );
  NAND4_X1 U7575 ( .A1(keyinput47), .A2(n6668), .A3(keyinput45), .A4(n6667), 
        .ZN(n6669) );
  NOR4_X1 U7576 ( .A1(keyinput39), .A2(keyinput14), .A3(n6670), .A4(n6669), 
        .ZN(n6671) );
  NAND4_X1 U7577 ( .A1(keyinput58), .A2(keyinput31), .A3(n6672), .A4(n6671), 
        .ZN(n6679) );
  NAND3_X1 U7578 ( .A1(keyinput20), .A2(keyinput15), .A3(keyinput50), .ZN(
        n6678) );
  NOR3_X1 U7579 ( .A1(keyinput52), .A2(keyinput6), .A3(keyinput9), .ZN(n6676)
         );
  INV_X1 U7580 ( .A(keyinput19), .ZN(n6673) );
  NOR4_X1 U7581 ( .A1(keyinput61), .A2(keyinput33), .A3(keyinput40), .A4(n6673), .ZN(n6675) );
  NOR4_X1 U7582 ( .A1(keyinput4), .A2(keyinput41), .A3(keyinput12), .A4(
        keyinput25), .ZN(n6674) );
  NAND4_X1 U7583 ( .A1(keyinput3), .A2(n6676), .A3(n6675), .A4(n6674), .ZN(
        n6677) );
  NOR4_X1 U7584 ( .A1(keyinput35), .A2(n6679), .A3(n6678), .A4(n6677), .ZN(
        n6680) );
  NAND4_X1 U7585 ( .A1(n6683), .A2(n6682), .A3(n6681), .A4(n6680), .ZN(n6684)
         );
  NAND4_X1 U7586 ( .A1(n6687), .A2(n6686), .A3(n6685), .A4(n6684), .ZN(n6690)
         );
  NAND2_X1 U7587 ( .A1(n6688), .A2(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6689) );
  XOR2_X1 U7588 ( .A(n6690), .B(n6689), .Z(U3180) );
  CLKBUF_X1 U3420 ( .A(n3333), .Z(n2957) );
  CLKBUF_X1 U3421 ( .A(n4527), .Z(n2961) );
  CLKBUF_X1 U3427 ( .A(n3198), .Z(n5402) );
  CLKBUF_X1 U3431 ( .A(n5423), .Z(n5437) );
  CLKBUF_X1 U3432 ( .A(n3218), .Z(n4607) );
endmodule

