

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940,
         n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
         n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
         n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964,
         n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972,
         n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
         n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
         n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
         n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
         n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
         n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036,
         n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044,
         n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
         n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
         n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068,
         n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076,
         n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
         n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
         n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
         n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108,
         n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
         n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
         n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132,
         n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
         n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
         n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156,
         n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164,
         n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
         n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180,
         n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
         n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196,
         n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204,
         n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212,
         n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220,
         n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228,
         n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236,
         n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
         n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252,
         n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260,
         n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268,
         n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276,
         n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284,
         n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292,
         n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300,
         n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308,
         n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
         n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324,
         n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332,
         n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340,
         n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348,
         n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356,
         n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364,
         n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372,
         n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380,
         n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388,
         n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396,
         n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404,
         n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412,
         n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420,
         n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428,
         n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436,
         n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444,
         n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452,
         n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460,
         n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468,
         n21469, n21470;

  CLKBUF_X1 U11024 ( .A(n16329), .Z(n9583) );
  INV_X1 U11025 ( .A(n17768), .ZN(n17785) );
  INV_X1 U11026 ( .A(n20781), .ZN(n20757) );
  NAND2_X1 U11027 ( .A1(n11209), .A2(n11208), .ZN(n16130) );
  CLKBUF_X2 U11028 ( .A(n17438), .Z(n17653) );
  NAND2_X1 U11029 ( .A1(n11351), .A2(n11350), .ZN(n13677) );
  CLKBUF_X2 U11030 ( .A(n13230), .Z(n17946) );
  CLKBUF_X1 U11031 ( .A(n11302), .Z(n11303) );
  INV_X2 U11032 ( .A(n11093), .ZN(n19989) );
  CLKBUF_X1 U11033 ( .A(n13082), .Z(n17824) );
  CLKBUF_X2 U11035 ( .A(n13202), .Z(n17945) );
  AND2_X1 U11036 ( .A1(n9872), .A2(n13839), .ZN(n15613) );
  CLKBUF_X2 U11037 ( .A(n13232), .Z(n18010) );
  CLKBUF_X1 U11038 ( .A(n13230), .Z(n18063) );
  CLKBUF_X3 U11039 ( .A(n13082), .Z(n9588) );
  INV_X1 U11040 ( .A(n13197), .ZN(n17961) );
  NAND2_X1 U11041 ( .A1(n10615), .A2(n10614), .ZN(n10782) );
  CLKBUF_X2 U11042 ( .A(n10895), .Z(n14541) );
  CLKBUF_X1 U11044 ( .A(n20758), .Z(n9580) );
  NOR2_X1 U11045 ( .A1(n15026), .A2(n12911), .ZN(n20758) );
  INV_X1 U11046 ( .A(n12351), .ZN(n12485) );
  NAND2_X1 U11047 ( .A1(n11268), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n9792) );
  INV_X1 U11048 ( .A(n11744), .ZN(n12199) );
  NAND2_X1 U11049 ( .A1(n13839), .A2(n12719), .ZN(n12977) );
  INV_X1 U11050 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15614) );
  NOR2_X1 U11051 ( .A1(n11570), .A2(n11569), .ZN(n11603) );
  INV_X1 U11052 ( .A(n12672), .ZN(n10793) );
  INV_X1 U11053 ( .A(n13622), .ZN(n13519) );
  AND2_X1 U11054 ( .A1(n13563), .A2(n12719), .ZN(n9699) );
  INV_X2 U11055 ( .A(n12943), .ZN(n12944) );
  INV_X2 U11056 ( .A(n21470), .ZN(n13741) );
  NAND2_X1 U11057 ( .A1(n13625), .A2(n15614), .ZN(n11767) );
  NOR2_X1 U11058 ( .A1(n11287), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11286) );
  AND2_X1 U11059 ( .A1(n11278), .A2(n10786), .ZN(n13574) );
  INV_X2 U11060 ( .A(n11542), .ZN(n11096) );
  NAND2_X2 U11061 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19508) );
  NOR2_X1 U11062 ( .A1(n9906), .A2(n9703), .ZN(n13008) );
  CLKBUF_X2 U11064 ( .A(n11304), .Z(n11475) );
  AND2_X1 U11065 ( .A1(n16391), .A2(n16389), .ZN(n14389) );
  INV_X1 U11066 ( .A(n18578), .ZN(n18566) );
  INV_X1 U11067 ( .A(n17743), .ZN(n19056) );
  NOR2_X1 U11068 ( .A1(n20735), .A2(n12927), .ZN(n17160) );
  INV_X1 U11069 ( .A(n19866), .ZN(n10245) );
  AND2_X1 U11070 ( .A1(n13927), .A2(n13874), .ZN(n20637) );
  INV_X1 U11071 ( .A(n13529), .ZN(n20685) );
  AOI211_X2 U11072 ( .C1(n13290), .C2(n13289), .A(n13293), .B(n13292), .ZN(
        n19529) );
  NOR2_X1 U11073 ( .A1(n18189), .A2(n21358), .ZN(n18188) );
  INV_X1 U11074 ( .A(n19084), .ZN(n18213) );
  INV_X1 U11075 ( .A(n10142), .ZN(n18634) );
  INV_X1 U11076 ( .A(n21303), .ZN(n21309) );
  INV_X1 U11078 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20276) );
  INV_X2 U11079 ( .A(n20700), .ZN(n20699) );
  NAND2_X1 U11080 ( .A1(n19059), .A2(n13326), .ZN(n18725) );
  INV_X2 U11081 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13162) );
  INV_X1 U11082 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13161) );
  CLKBUF_X3 U11083 ( .A(n11311), .Z(n9599) );
  NAND2_X1 U11084 ( .A1(n11680), .A2(n11679), .ZN(n9581) );
  INV_X2 U11085 ( .A(n13777), .ZN(n13818) );
  AND2_X2 U11086 ( .A1(n18596), .A2(n13337), .ZN(n18962) );
  INV_X1 U11087 ( .A(n19074), .ZN(n18113) );
  NAND2_X2 U11088 ( .A1(n10102), .A2(n11879), .ZN(n11880) );
  NOR2_X2 U11089 ( .A1(n14860), .A2(n12933), .ZN(n14824) );
  NOR2_X2 U11090 ( .A1(n17618), .A2(n17983), .ZN(n17996) );
  NOR2_X2 U11091 ( .A1(n18626), .A2(n13328), .ZN(n17434) );
  NAND2_X2 U11093 ( .A1(n17165), .A2(n12771), .ZN(n15385) );
  OAI21_X2 U11094 ( .B1(n14708), .B2(n10297), .A(n10294), .ZN(n9833) );
  NAND2_X2 U11095 ( .A1(n11826), .A2(n11825), .ZN(n11881) );
  NAND2_X2 U11096 ( .A1(n11287), .A2(n10784), .ZN(n12672) );
  XNOR2_X1 U11097 ( .A(n12725), .B(n13672), .ZN(n13792) );
  AOI211_X2 U11098 ( .C1(n9580), .C2(n15405), .A(n14768), .B(n14767), .ZN(
        n14769) );
  AOI211_X2 U11099 ( .C1(n15415), .C2(n9580), .A(n14782), .B(n14781), .ZN(
        n14783) );
  NAND2_X2 U11100 ( .A1(n10468), .A2(n10466), .ZN(n13766) );
  AND2_X4 U11101 ( .A1(n13624), .A2(n11565), .ZN(n11733) );
  AND2_X2 U11102 ( .A1(n9981), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11565) );
  AOI21_X2 U11103 ( .B1(n13863), .B2(n13862), .A(n13861), .ZN(n14056) );
  NOR2_X4 U11104 ( .A1(n17287), .A2(n18724), .ZN(n18636) );
  NAND2_X1 U11105 ( .A1(n13326), .A2(n19691), .ZN(n18724) );
  INV_X1 U11106 ( .A(n18062), .ZN(n9584) );
  INV_X4 U11107 ( .A(n17889), .ZN(n18062) );
  OAI211_X2 U11108 ( .C1(n10833), .C2(n10838), .A(n10837), .B(n9792), .ZN(
        n11182) );
  OAI21_X1 U11110 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19699), .A(n17401), 
        .ZN(n18721) );
  NAND2_X1 U11112 ( .A1(n14389), .A2(n14388), .ZN(n16378) );
  NAND2_X1 U11113 ( .A1(n14360), .A2(n14722), .ZN(n16410) );
  NAND2_X1 U11114 ( .A1(n10131), .A2(n9654), .ZN(n16329) );
  OAI21_X1 U11115 ( .B1(n10281), .B2(n10123), .A(n10077), .ZN(n12781) );
  OR2_X1 U11116 ( .A1(n10292), .A2(n9968), .ZN(n9817) );
  NOR2_X2 U11117 ( .A1(n15779), .A2(n15778), .ZN(n15781) );
  NAND2_X1 U11118 ( .A1(n13151), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n18382) );
  OR2_X1 U11119 ( .A1(n13151), .A2(n10139), .ZN(n13155) );
  INV_X1 U11120 ( .A(n20248), .ZN(n20292) );
  NAND2_X1 U11121 ( .A1(n9969), .A2(n11543), .ZN(n16517) );
  OAI211_X1 U11122 ( .C1(n18408), .C2(n18409), .A(n10536), .B(n18407), .ZN(
        n18393) );
  OR2_X1 U11123 ( .A1(n11039), .A2(n11038), .ZN(n15891) );
  NAND2_X2 U11124 ( .A1(n18514), .A2(n10142), .ZN(n18427) );
  CLKBUF_X2 U11125 ( .A(n12777), .Z(n15353) );
  AND2_X1 U11126 ( .A1(n14865), .A2(n14866), .ZN(n14868) );
  NOR2_X2 U11127 ( .A1(n10882), .A2(n16831), .ZN(n20035) );
  AND2_X1 U11128 ( .A1(n10874), .A2(n10875), .ZN(n20243) );
  AOI22_X1 U11129 ( .A1(n19529), .A2(n18893), .B1(n18954), .B2(n13356), .ZN(
        n19533) );
  INV_X1 U11130 ( .A(n16831), .ZN(n9927) );
  AND2_X1 U11131 ( .A1(n13650), .A2(n9668), .ZN(n15965) );
  NAND2_X1 U11132 ( .A1(n17415), .A2(n13268), .ZN(n13288) );
  OR3_X1 U11133 ( .A1(n12195), .A2(n15300), .A3(n14907), .ZN(n12178) );
  XNOR2_X1 U11134 ( .A(n13331), .B(n13330), .ZN(n17438) );
  NAND2_X1 U11135 ( .A1(n12515), .A2(n12514), .ZN(n12522) );
  OAI211_X2 U11136 ( .C1(n11523), .C2(n11443), .A(n11300), .B(n11289), .ZN(
        n13610) );
  NAND2_X1 U11137 ( .A1(n10196), .A2(n13262), .ZN(n13355) );
  NAND3_X1 U11138 ( .A1(n10544), .A2(n13048), .A3(n10538), .ZN(n13298) );
  NOR2_X1 U11139 ( .A1(n13218), .A2(n13217), .ZN(n19066) );
  INV_X1 U11140 ( .A(n10782), .ZN(n11278) );
  NOR2_X1 U11141 ( .A1(n10794), .A2(n10782), .ZN(n10797) );
  AND2_X1 U11142 ( .A1(n11287), .A2(n20276), .ZN(n11311) );
  NAND2_X1 U11143 ( .A1(n11603), .A2(n11602), .ZN(n12575) );
  NAND2_X1 U11144 ( .A1(n10598), .A2(n10597), .ZN(n11287) );
  BUF_X2 U11145 ( .A(n13061), .Z(n18066) );
  CLKBUF_X2 U11146 ( .A(n17816), .Z(n17043) );
  CLKBUF_X2 U11147 ( .A(n11733), .Z(n12430) );
  CLKBUF_X2 U11148 ( .A(n13252), .Z(n18001) );
  INV_X2 U11149 ( .A(n19024), .ZN(n9586) );
  CLKBUF_X2 U11150 ( .A(n13076), .Z(n18059) );
  BUF_X4 U11151 ( .A(n13253), .Z(n9587) );
  BUF_X4 U11152 ( .A(n13049), .Z(n9594) );
  CLKBUF_X2 U11153 ( .A(n10887), .Z(n9595) );
  INV_X1 U11154 ( .A(n13223), .ZN(n17830) );
  INV_X4 U11155 ( .A(n13197), .ZN(n9589) );
  NOR2_X1 U11156 ( .A1(n13041), .A2(n13040), .ZN(n13049) );
  INV_X4 U11157 ( .A(n11926), .ZN(n11732) );
  CLKBUF_X2 U11158 ( .A(n13232), .Z(n18046) );
  BUF_X4 U11159 ( .A(n13184), .Z(n9590) );
  AND2_X1 U11160 ( .A1(n14514), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10887) );
  AND2_X2 U11161 ( .A1(n14509), .A2(n10750), .ZN(n10620) );
  NAND2_X2 U11162 ( .A1(n15666), .A2(n11563), .ZN(n11926) );
  OR2_X1 U11163 ( .A1(n13044), .A2(n19508), .ZN(n13223) );
  NAND2_X2 U11164 ( .A1(n13625), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11667) );
  INV_X2 U11165 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n11830) );
  INV_X4 U11166 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19654) );
  INV_X4 U11167 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10750) );
  AND2_X1 U11168 ( .A1(n15370), .A2(n15369), .ZN(n15582) );
  AOI21_X1 U11169 ( .B1(n14730), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n14729), .ZN(n14731) );
  OAI21_X1 U11170 ( .B1(n16690), .B2(n16550), .A(n9965), .ZN(n9964) );
  AOI21_X1 U11171 ( .B1(n9884), .B2(n16351), .A(n9801), .ZN(n9800) );
  NAND2_X1 U11172 ( .A1(n12782), .A2(n15197), .ZN(n10174) );
  OR2_X1 U11173 ( .A1(n16292), .A2(n10357), .ZN(n10351) );
  OAI21_X1 U11174 ( .B1(n16711), .B2(n16550), .A(n9857), .ZN(n9856) );
  OAI21_X1 U11175 ( .B1(n9808), .B2(n10046), .A(n10044), .ZN(n9811) );
  OAI21_X1 U11176 ( .B1(n16643), .B2(n16550), .A(n9854), .ZN(n9853) );
  AND2_X1 U11177 ( .A1(n9851), .A2(n9850), .ZN(n16309) );
  NOR2_X1 U11178 ( .A1(n16431), .A2(n9683), .ZN(n9766) );
  AOI21_X1 U11179 ( .B1(n14749), .B2(n19945), .A(n14748), .ZN(n14750) );
  NAND2_X1 U11180 ( .A1(n10021), .A2(n10020), .ZN(n16292) );
  OAI21_X1 U11181 ( .B1(n16316), .B2(n9687), .A(n14318), .ZN(n14321) );
  AND2_X1 U11182 ( .A1(n9967), .A2(n14716), .ZN(n16664) );
  OAI21_X1 U11183 ( .B1(n15205), .B2(n15178), .A(n15374), .ZN(n15197) );
  AND2_X1 U11184 ( .A1(n9773), .A2(n9828), .ZN(n9772) );
  AOI21_X1 U11185 ( .B1(n16061), .B2(n10460), .A(n16056), .ZN(n16050) );
  NOR2_X1 U11186 ( .A1(n9916), .A2(n16450), .ZN(n16724) );
  AOI21_X1 U11187 ( .B1(n16378), .B2(n16377), .A(n16376), .ZN(n16382) );
  AND2_X1 U11188 ( .A1(n14398), .A2(n14364), .ZN(n14385) );
  NOR2_X1 U11189 ( .A1(n16353), .A2(n16354), .ZN(n16630) );
  OAI21_X1 U11190 ( .B1(n16410), .B2(n19970), .A(n14723), .ZN(n16662) );
  OR2_X1 U11191 ( .A1(n15207), .A2(n15448), .ZN(n15219) );
  AOI211_X1 U11192 ( .C1(BUF1_REG_30__SCAN_IN), .C2(n16259), .A(n14699), .B(
        n14698), .ZN(n14700) );
  AND2_X1 U11193 ( .A1(n9914), .A2(n16451), .ZN(n9916) );
  INV_X1 U11194 ( .A(n10067), .ZN(n16450) );
  AOI21_X1 U11195 ( .B1(n9847), .B2(n9844), .A(n9692), .ZN(n9970) );
  XNOR2_X1 U11196 ( .A(n11550), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14749) );
  NOR2_X1 U11197 ( .A1(n12674), .A2(n10242), .ZN(n10241) );
  OAI21_X1 U11198 ( .B1(n14389), .B2(n10217), .A(n10216), .ZN(n10214) );
  OAI21_X1 U11199 ( .B1(n16369), .B2(n16365), .A(n16366), .ZN(n16362) );
  NAND2_X1 U11200 ( .A1(n14360), .A2(n14396), .ZN(n10008) );
  AND2_X1 U11201 ( .A1(n14360), .A2(n9631), .ZN(n16351) );
  AND2_X1 U11202 ( .A1(n9933), .A2(n9697), .ZN(n9932) );
  NAND2_X1 U11203 ( .A1(n14360), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16476) );
  NAND2_X1 U11204 ( .A1(n9925), .A2(n10363), .ZN(n10009) );
  NAND2_X1 U11205 ( .A1(n10417), .A2(n9600), .ZN(n14708) );
  NAND2_X1 U11206 ( .A1(n14360), .A2(n10110), .ZN(n16394) );
  XNOR2_X1 U11207 ( .A(n11101), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11102) );
  NOR2_X1 U11208 ( .A1(n14629), .A2(n14628), .ZN(n16055) );
  OR2_X1 U11209 ( .A1(n16312), .A2(n10525), .ZN(n11550) );
  XNOR2_X1 U11210 ( .A(n15774), .B(n12680), .ZN(n14701) );
  NAND2_X1 U11211 ( .A1(n12683), .A2(n12682), .ZN(n14697) );
  AND2_X1 U11212 ( .A1(n10011), .A2(n16318), .ZN(n9934) );
  AND2_X1 U11213 ( .A1(n9860), .A2(n10136), .ZN(n10371) );
  AND2_X1 U11214 ( .A1(n10231), .A2(n10230), .ZN(n13159) );
  NOR2_X1 U11215 ( .A1(n18365), .A2(n18364), .ZN(n18363) );
  AND2_X1 U11216 ( .A1(n16328), .A2(n16333), .ZN(n10011) );
  NAND2_X1 U11217 ( .A1(n15781), .A2(n12681), .ZN(n12683) );
  AND3_X1 U11218 ( .A1(n10136), .A2(n10130), .A3(n11546), .ZN(n9795) );
  NAND2_X1 U11219 ( .A1(n9793), .A2(n11538), .ZN(n9860) );
  XNOR2_X1 U11220 ( .A(n11098), .B(n11094), .ZN(n12688) );
  AND2_X1 U11221 ( .A1(n9821), .A2(n9820), .ZN(n18365) );
  OR2_X1 U11222 ( .A1(n15812), .A2(n15811), .ZN(n16583) );
  INV_X1 U11223 ( .A(n11540), .ZN(n11538) );
  NAND2_X1 U11224 ( .A1(n10372), .A2(n10104), .ZN(n10370) );
  OR2_X1 U11225 ( .A1(n16457), .A2(n16456), .ZN(n16505) );
  NAND2_X1 U11226 ( .A1(n10287), .A2(n10290), .ZN(n10007) );
  NAND2_X1 U11227 ( .A1(n11006), .A2(n10530), .ZN(n10292) );
  NOR2_X1 U11228 ( .A1(n13155), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17134) );
  OR2_X1 U11229 ( .A1(n11068), .A2(n16354), .ZN(n16366) );
  NOR3_X1 U11230 ( .A1(n14793), .A2(n14765), .A3(n21272), .ZN(n12951) );
  NAND2_X1 U11231 ( .A1(n16514), .A2(n11008), .ZN(n10290) );
  NAND2_X1 U11232 ( .A1(n10108), .A2(n9794), .ZN(n11539) );
  AND3_X1 U11233 ( .A1(n11536), .A2(n16534), .A3(n16805), .ZN(n10104) );
  NAND2_X1 U11234 ( .A1(n9879), .A2(n9878), .ZN(n16805) );
  AND2_X1 U11235 ( .A1(n9954), .A2(n9953), .ZN(n11546) );
  NAND2_X1 U11236 ( .A1(n9961), .A2(n16791), .ZN(n16534) );
  OAI22_X1 U11237 ( .A1(n9651), .A2(n16807), .B1(n16792), .B2(n10972), .ZN(
        n16529) );
  AOI21_X1 U11238 ( .B1(n9771), .B2(n15976), .A(n16791), .ZN(n10293) );
  NAND2_X1 U11239 ( .A1(n16120), .A2(n9736), .ZN(n16078) );
  NAND2_X1 U11240 ( .A1(n20857), .A2(n12746), .ZN(n17180) );
  NAND2_X1 U11241 ( .A1(n10066), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11541) );
  OR2_X1 U11242 ( .A1(n20309), .A2(n20247), .ZN(n20248) );
  OR2_X1 U11243 ( .A1(n15891), .A2(n11542), .ZN(n11049) );
  NAND2_X2 U11244 ( .A1(n12913), .A2(n12912), .ZN(n12914) );
  NOR2_X2 U11245 ( .A1(n20309), .A2(n20629), .ZN(n10554) );
  NOR2_X2 U11246 ( .A1(n20405), .A2(n20630), .ZN(n20340) );
  NOR2_X2 U11247 ( .A1(n20405), .A2(n20247), .ZN(n10547) );
  NAND2_X2 U11248 ( .A1(n10983), .A2(n9802), .ZN(n11543) );
  NAND2_X1 U11249 ( .A1(n10039), .A2(n10142), .ZN(n18407) );
  AND2_X1 U11250 ( .A1(n9661), .A2(n11010), .ZN(n19752) );
  NAND2_X1 U11251 ( .A1(n20637), .A2(n20664), .ZN(n20309) );
  OR2_X1 U11252 ( .A1(n19763), .A2(n11542), .ZN(n11064) );
  OR2_X1 U11253 ( .A1(n20637), .A2(n20664), .ZN(n20146) );
  AND2_X1 U11254 ( .A1(n10212), .A2(n10954), .ZN(n9802) );
  AND3_X2 U11255 ( .A1(n10904), .A2(n9738), .A3(n9835), .ZN(n10983) );
  AND2_X1 U11256 ( .A1(n9770), .A2(n10937), .ZN(n10212) );
  NAND2_X1 U11257 ( .A1(n13148), .A2(n10226), .ZN(n10225) );
  OAI21_X1 U11258 ( .B1(n18518), .B2(n9745), .A(n10533), .ZN(n13148) );
  AND4_X1 U11259 ( .A1(n10914), .A2(n10913), .A3(n10912), .A4(n10911), .ZN(
        n10917) );
  NOR2_X1 U11260 ( .A1(n16810), .A2(n11505), .ZN(n16740) );
  XNOR2_X1 U11261 ( .A(n13859), .B(n13863), .ZN(n20647) );
  INV_X1 U11262 ( .A(n11917), .ZN(n10445) );
  NAND2_X1 U11263 ( .A1(n12696), .A2(n12695), .ZN(n12777) );
  NOR2_X2 U11264 ( .A1(n10882), .A2(n9927), .ZN(n16877) );
  AOI21_X1 U11265 ( .B1(n20243), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A(
        n20688), .ZN(n10878) );
  NAND2_X1 U11266 ( .A1(n11958), .A2(n11957), .ZN(n12696) );
  INV_X2 U11267 ( .A(n13600), .ZN(n13702) );
  OR2_X1 U11268 ( .A1(n10881), .A2(n10873), .ZN(n20143) );
  INV_X1 U11269 ( .A(n13976), .ZN(n11198) );
  OAI21_X1 U11270 ( .B1(n11826), .B2(n11825), .A(n11881), .ZN(n14006) );
  NAND2_X1 U11271 ( .A1(n10869), .A2(n10868), .ZN(n10882) );
  NAND2_X1 U11272 ( .A1(n10869), .A2(n10552), .ZN(n16890) );
  OAI21_X1 U11273 ( .B1(n18596), .B2(n10232), .A(n10142), .ZN(n13146) );
  INV_X1 U11274 ( .A(n11881), .ZN(n10083) );
  NOR2_X1 U11275 ( .A1(n13846), .A2(n13813), .ZN(n21184) );
  NAND2_X1 U11276 ( .A1(n13143), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13337) );
  NOR2_X2 U11277 ( .A1(n13846), .A2(n13818), .ZN(n21138) );
  AOI211_X1 U11278 ( .C1(n14712), .C2(n13659), .A(n13654), .B(n19961), .ZN(
        n17224) );
  AND2_X1 U11279 ( .A1(n16007), .A2(n14344), .ZN(n10861) );
  AND2_X1 U11280 ( .A1(n14994), .A2(n9712), .ZN(n14946) );
  NOR2_X2 U11281 ( .A1(n19533), .A2(n19547), .ZN(n13326) );
  INV_X1 U11282 ( .A(n10881), .ZN(n10869) );
  NOR2_X1 U11283 ( .A1(n13846), .A2(n13834), .ZN(n21193) );
  INV_X1 U11284 ( .A(n13766), .ZN(n10868) );
  NOR2_X1 U11285 ( .A1(n13846), .A2(n13823), .ZN(n21166) );
  NOR2_X1 U11286 ( .A1(n13846), .A2(n13829), .ZN(n21154) );
  NAND2_X1 U11287 ( .A1(n13867), .A2(n13866), .ZN(n14054) );
  AND2_X2 U11288 ( .A1(n20712), .A2(n12794), .ZN(n20882) );
  NOR2_X2 U11289 ( .A1(n14282), .A2(n14281), .ZN(n14994) );
  NOR2_X2 U11290 ( .A1(n17599), .A2(n17981), .ZN(n17954) );
  NAND2_X1 U11291 ( .A1(n13584), .A2(n13583), .ZN(n16826) );
  NAND2_X1 U11292 ( .A1(n10052), .A2(n10051), .ZN(n14754) );
  CLKBUF_X1 U11293 ( .A(n13938), .Z(n15657) );
  INV_X1 U11294 ( .A(n13775), .ZN(n10052) );
  NAND2_X1 U11295 ( .A1(n18639), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10223) );
  NAND2_X1 U11296 ( .A1(n10423), .A2(n10421), .ZN(n14282) );
  XNOR2_X1 U11297 ( .A(n13140), .B(n13139), .ZN(n18639) );
  NAND3_X1 U11298 ( .A1(n10846), .A2(n9829), .A3(n10033), .ZN(n10129) );
  CLKBUF_X1 U11299 ( .A(n14113), .Z(n21060) );
  NAND2_X1 U11300 ( .A1(n11076), .A2(n10716), .ZN(n10984) );
  INV_X4 U11301 ( .A(n19499), .ZN(n19494) );
  OR2_X1 U11302 ( .A1(n14175), .A2(n14176), .ZN(n14259) );
  NAND2_X1 U11303 ( .A1(n10843), .A2(n10107), .ZN(n9829) );
  AND2_X1 U11304 ( .A1(n9834), .A2(n10033), .ZN(n10843) );
  NAND2_X1 U11305 ( .A1(n11758), .A2(n10069), .ZN(n13797) );
  OR2_X2 U11306 ( .A1(n10986), .A2(n11093), .ZN(n11076) );
  OR2_X1 U11307 ( .A1(n10986), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10716) );
  NAND2_X1 U11308 ( .A1(n10851), .A2(n10850), .ZN(n10855) );
  NAND2_X1 U11309 ( .A1(n19491), .A2(n19486), .ZN(n17416) );
  NAND2_X1 U11310 ( .A1(n10990), .A2(n10991), .ZN(n10986) );
  OR2_X1 U11311 ( .A1(n10064), .A2(n10062), .ZN(n10061) );
  CLKBUF_X1 U11312 ( .A(n11722), .Z(n11723) );
  AND2_X1 U11313 ( .A1(n9789), .A2(n9788), .ZN(n10828) );
  INV_X4 U11314 ( .A(n11273), .ZN(n11268) );
  INV_X2 U11315 ( .A(n11247), .ZN(n11267) );
  CLKBUF_X1 U11316 ( .A(n16818), .Z(n16855) );
  NAND2_X1 U11317 ( .A1(n10259), .A2(n10257), .ZN(n17145) );
  NAND2_X1 U11318 ( .A1(n9841), .A2(n9838), .ZN(n10836) );
  NAND2_X1 U11319 ( .A1(n9791), .A2(n10798), .ZN(n10830) );
  AND3_X1 U11320 ( .A1(n11317), .A2(n11316), .A3(n11315), .ZN(n15996) );
  NAND2_X1 U11321 ( .A1(n13266), .A2(n19486), .ZN(n17400) );
  NOR2_X1 U11322 ( .A1(n10673), .A2(n10016), .ZN(n10015) );
  AND3_X1 U11323 ( .A1(n11323), .A2(n11322), .A3(n11321), .ZN(n15982) );
  CLKBUF_X1 U11324 ( .A(n12566), .Z(n17210) );
  OR2_X1 U11325 ( .A1(n11134), .A2(n11093), .ZN(n10650) );
  INV_X1 U11326 ( .A(n12543), .ZN(n12542) );
  NOR2_X1 U11327 ( .A1(n13125), .A2(n18229), .ZN(n13138) );
  INV_X1 U11328 ( .A(n10971), .ZN(n10673) );
  NOR2_X1 U11329 ( .A1(n10804), .A2(n20690), .ZN(n9838) );
  NOR2_X1 U11330 ( .A1(n13267), .A2(n19482), .ZN(n16966) );
  NAND2_X1 U11331 ( .A1(n10648), .A2(n10647), .ZN(n11134) );
  AND2_X1 U11332 ( .A1(n10792), .A2(n10793), .ZN(n9841) );
  AND2_X1 U11333 ( .A1(n10791), .A2(n20689), .ZN(n10138) );
  CLKBUF_X1 U11334 ( .A(n11166), .Z(n16960) );
  AND2_X1 U11335 ( .A1(n11708), .A2(n11707), .ZN(n12959) );
  NOR2_X1 U11336 ( .A1(n13278), .A2(n9681), .ZN(n9938) );
  NAND2_X1 U11337 ( .A1(n11180), .A2(n10801), .ZN(n11481) );
  NAND2_X1 U11338 ( .A1(n10795), .A2(n9832), .ZN(n10804) );
  INV_X1 U11339 ( .A(n13355), .ZN(n19078) );
  NAND3_X1 U11340 ( .A1(n13196), .A2(n13195), .A3(n13194), .ZN(n17743) );
  NAND2_X1 U11341 ( .A1(n11706), .A2(n11697), .ZN(n12120) );
  CLKBUF_X1 U11342 ( .A(n11935), .Z(n12511) );
  NAND2_X1 U11343 ( .A1(n10103), .A2(n10797), .ZN(n11166) );
  INV_X2 U11344 ( .A(n11280), .ZN(n20688) );
  NOR2_X1 U11345 ( .A1(n18236), .A2(n13102), .ZN(n13114) );
  AND2_X2 U11346 ( .A1(n9807), .A2(n10788), .ZN(n10792) );
  OR2_X1 U11347 ( .A1(n10666), .A2(n10665), .ZN(n11535) );
  NAND2_X1 U11348 ( .A1(n13298), .A2(n18247), .ZN(n13102) );
  INV_X1 U11349 ( .A(n12719), .ZN(n13823) );
  INV_X2 U11350 ( .A(n19059), .ZN(n19691) );
  INV_X1 U11351 ( .A(n11706), .ZN(n12958) );
  AOI21_X2 U11352 ( .B1(n12575), .B2(n13808), .A(n11627), .ZN(n11707) );
  NAND2_X1 U11353 ( .A1(n13829), .A2(n13777), .ZN(n13622) );
  CLKBUF_X1 U11354 ( .A(n11701), .Z(n13760) );
  NOR2_X1 U11355 ( .A1(n19084), .A2(n19066), .ZN(n13285) );
  NOR2_X1 U11356 ( .A1(n17432), .A2(n18472), .ZN(n18446) );
  CLKBUF_X1 U11357 ( .A(n11827), .Z(n13813) );
  BUF_X1 U11358 ( .A(n10789), .Z(n19984) );
  INV_X2 U11359 ( .A(U212), .ZN(n17351) );
  INV_X2 U11360 ( .A(n17304), .ZN(n17354) );
  OR2_X2 U11361 ( .A1(n13059), .A2(n13060), .ZN(n18247) );
  NOR2_X2 U11362 ( .A1(n13182), .A2(n13181), .ZN(n19059) );
  OR2_X1 U11363 ( .A1(n10629), .A2(n10628), .ZN(n11524) );
  INV_X1 U11364 ( .A(n10783), .ZN(n10788) );
  OR2_X1 U11365 ( .A1(n10641), .A2(n10640), .ZN(n10919) );
  CLKBUF_X1 U11366 ( .A(n11829), .Z(n13758) );
  INV_X2 U11368 ( .A(n13563), .ZN(n13829) );
  AND2_X1 U11369 ( .A1(n11602), .A2(n11603), .ZN(n11827) );
  NAND4_X2 U11370 ( .A1(n11626), .A2(n11625), .A3(n11624), .A4(n11623), .ZN(
        n11829) );
  INV_X1 U11371 ( .A(n10789), .ZN(n9591) );
  AND3_X1 U11372 ( .A1(n10555), .A2(n11674), .A3(n11673), .ZN(n11680) );
  AND2_X2 U11373 ( .A1(n11644), .A2(n11643), .ZN(n13839) );
  OAI21_X1 U11374 ( .B1(n10591), .B2(n10590), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10598) );
  NOR2_X2 U11375 ( .A1(n15085), .A2(n15382), .ZN(n13804) );
  AOI21_X1 U11376 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n19514), .A(
        n13164), .ZN(n13165) );
  NOR2_X1 U11377 ( .A1(n11596), .A2(n11595), .ZN(n11601) );
  AND4_X1 U11378 ( .A1(n11574), .A2(n11573), .A3(n11572), .A4(n11571), .ZN(
        n11607) );
  AND4_X1 U11379 ( .A1(n11578), .A2(n11577), .A3(n11576), .A4(n11575), .ZN(
        n11606) );
  AND4_X1 U11380 ( .A1(n11557), .A2(n11556), .A3(n11555), .A4(n11554), .ZN(
        n11602) );
  AND3_X1 U11381 ( .A1(n11691), .A2(n11690), .A3(n11689), .ZN(n11692) );
  AND4_X1 U11382 ( .A1(n11672), .A2(n11671), .A3(n11670), .A4(n11669), .ZN(
        n11673) );
  AND4_X1 U11383 ( .A1(n11619), .A2(n11618), .A3(n11617), .A4(n11616), .ZN(
        n11624) );
  CLKBUF_X2 U11384 ( .A(n10893), .Z(n14539) );
  INV_X1 U11385 ( .A(n9587), .ZN(n9592) );
  BUF_X2 U11386 ( .A(n10893), .Z(n14478) );
  CLKBUF_X3 U11387 ( .A(n17816), .Z(n16999) );
  NAND2_X2 U11388 ( .A1(n19708), .A2(n19696), .ZN(n19024) );
  NAND2_X1 U11389 ( .A1(n10154), .A2(n10255), .ZN(n17889) );
  BUF_X2 U11390 ( .A(n13061), .Z(n18044) );
  BUF_X2 U11391 ( .A(n13081), .Z(n17960) );
  INV_X2 U11392 ( .A(n13183), .ZN(n18045) );
  CLKBUF_X3 U11393 ( .A(n13252), .Z(n18058) );
  INV_X2 U11394 ( .A(n12246), .ZN(n9593) );
  NAND2_X2 U11395 ( .A1(n20699), .A2(n20565), .ZN(n20614) );
  NAND2_X2 U11396 ( .A1(n19707), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19630) );
  AND2_X1 U11397 ( .A1(n14512), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10686) );
  AOI21_X1 U11398 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n21428), .A(
        n13163), .ZN(n13168) );
  INV_X2 U11399 ( .A(n17388), .ZN(n17390) );
  AND2_X2 U11400 ( .A1(n11564), .A2(n11563), .ZN(n11772) );
  AND2_X2 U11401 ( .A1(n11565), .A2(n15666), .ZN(n11868) );
  AND2_X2 U11402 ( .A1(n11565), .A2(n11564), .ZN(n11787) );
  AND2_X2 U11403 ( .A1(n14556), .A2(n10750), .ZN(n14533) );
  INV_X2 U11404 ( .A(n19705), .ZN(n19707) );
  AND2_X2 U11405 ( .A1(n14515), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14531) );
  INV_X1 U11406 ( .A(n18026), .ZN(n13183) );
  CLKBUF_X1 U11407 ( .A(n14509), .Z(n16854) );
  NAND2_X1 U11408 ( .A1(n14516), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10678) );
  CLKBUF_X3 U11409 ( .A(n10775), .Z(n14668) );
  NOR2_X1 U11410 ( .A1(n13033), .A2(n13042), .ZN(n13076) );
  INV_X1 U11411 ( .A(n13033), .ZN(n10154) );
  NOR2_X1 U11412 ( .A1(n13040), .A2(n13043), .ZN(n13230) );
  NAND2_X1 U11413 ( .A1(n10255), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n19493) );
  NOR2_X1 U11414 ( .A1(n13040), .A2(n13042), .ZN(n13082) );
  NOR2_X1 U11415 ( .A1(n13041), .A2(n17789), .ZN(n13252) );
  INV_X2 U11416 ( .A(n11767), .ZN(n12487) );
  AND2_X1 U11417 ( .A1(n10099), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10086) );
  AND2_X1 U11418 ( .A1(n13664), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11564) );
  AND3_X2 U11419 ( .A1(n10556), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14556) );
  AND2_X2 U11420 ( .A1(n13624), .A2(n11563), .ZN(n11739) );
  AND2_X2 U11421 ( .A1(n9836), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n16832) );
  AND2_X2 U11422 ( .A1(n15615), .A2(n11558), .ZN(n11738) );
  CLKBUF_X1 U11423 ( .A(n21029), .Z(n21149) );
  NAND2_X1 U11424 ( .A1(n13161), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13033) );
  NAND2_X1 U11425 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19654), .ZN(
        n13043) );
  NAND2_X1 U11426 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n13162), .ZN(
        n13040) );
  NAND2_X1 U11427 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19663), .ZN(
        n13041) );
  INV_X1 U11428 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16920) );
  INV_X1 U11429 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10556) );
  INV_X1 U11430 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9836) );
  NOR2_X2 U11431 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10560) );
  INV_X1 U11432 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16821) );
  AND2_X1 U11433 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15615) );
  AND2_X1 U11434 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11553) );
  NOR2_X2 U11435 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11563) );
  AND2_X1 U11436 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13624) );
  OR2_X2 U11437 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17789) );
  INV_X2 U11438 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19663) );
  INV_X4 U11439 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21428) );
  NOR3_X2 U11440 ( .A1(n17806), .A2(n17805), .A3(n17855), .ZN(n17848) );
  AOI21_X1 U11441 ( .B1(n12548), .B2(n12547), .A(n12546), .ZN(n12557) );
  NOR2_X2 U11442 ( .A1(n15871), .A2(n10516), .ZN(n15798) );
  NOR2_X2 U11443 ( .A1(n15026), .A2(n12923), .ZN(n20783) );
  INV_X2 U11444 ( .A(n10784), .ZN(n12597) );
  AND2_X2 U11445 ( .A1(n14712), .A2(n14714), .ZN(n19961) );
  AND2_X1 U11446 ( .A1(n13875), .A2(n10858), .ZN(n20069) );
  AND2_X1 U11447 ( .A1(n13875), .A2(n10859), .ZN(n20176) );
  NOR2_X2 U11448 ( .A1(n13934), .A2(n10508), .ZN(n14726) );
  NAND2_X2 U11449 ( .A1(n11417), .A2(n11416), .ZN(n13934) );
  NAND2_X2 U11450 ( .A1(n12811), .A2(n12912), .ZN(n20749) );
  NOR2_X2 U11451 ( .A1(n14369), .A2(n14370), .ZN(n14368) );
  NOR2_X2 U11452 ( .A1(n13677), .A2(n10502), .ZN(n13854) );
  CLKBUF_X2 U11453 ( .A(n10887), .Z(n9596) );
  INV_X4 U11454 ( .A(n17157), .ZN(n15023) );
  INV_X1 U11455 ( .A(n10678), .ZN(n9597) );
  INV_X1 U11456 ( .A(n10678), .ZN(n9598) );
  NOR2_X4 U11457 ( .A1(n19493), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13253) );
  NOR2_X2 U11458 ( .A1(n19656), .A2(n18716), .ZN(n18578) );
  NAND2_X1 U11459 ( .A1(n10289), .A2(n10288), .ZN(n10287) );
  AOI21_X1 U11460 ( .B1(n10293), .B2(n10530), .A(n10291), .ZN(n10288) );
  INV_X1 U11461 ( .A(n10797), .ZN(n10524) );
  NAND2_X1 U11462 ( .A1(n13845), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11862) );
  NOR2_X1 U11463 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11558) );
  NAND2_X1 U11464 ( .A1(n10820), .A2(n9730), .ZN(n10065) );
  NAND4_X1 U11465 ( .A1(n10808), .A2(n10529), .A3(n9591), .A4(n10788), .ZN(
        n10812) );
  NAND2_X2 U11466 ( .A1(n11862), .A2(n11861), .ZN(n12559) );
  INV_X1 U11467 ( .A(n13523), .ZN(n11861) );
  OR2_X1 U11468 ( .A1(n11794), .A2(n11793), .ZN(n12765) );
  AND2_X1 U11469 ( .A1(n16380), .A2(n11066), .ZN(n16346) );
  NAND2_X1 U11470 ( .A1(n10066), .A2(n11542), .ZN(n9771) );
  OAI211_X1 U11471 ( .C1(n10468), .C2(n16963), .A(n10464), .B(n10465), .ZN(
        n9787) );
  AND2_X1 U11472 ( .A1(n9948), .A2(n9947), .ZN(n19516) );
  NAND2_X1 U11473 ( .A1(n19660), .A2(n19534), .ZN(n9948) );
  NAND2_X1 U11474 ( .A1(n14861), .A2(n10097), .ZN(n14784) );
  AND2_X1 U11475 ( .A1(n9653), .A2(n14796), .ZN(n10097) );
  NOR2_X1 U11476 ( .A1(n17168), .A2(n10163), .ZN(n10162) );
  INV_X1 U11477 ( .A(n12763), .ZN(n10163) );
  NAND4_X2 U11478 ( .A1(n9795), .A2(n10370), .A3(n11539), .A4(n9860), .ZN(
        n10131) );
  AND2_X1 U11479 ( .A1(n9631), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10522) );
  NAND2_X1 U11480 ( .A1(n14360), .A2(n16409), .ZN(n16422) );
  NAND2_X1 U11481 ( .A1(n17073), .A2(n9763), .ZN(n13157) );
  NOR2_X1 U11482 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n9981), .ZN(
        n11552) );
  INV_X1 U11483 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10099) );
  NAND2_X1 U11484 ( .A1(n9764), .A2(n10524), .ZN(n11165) );
  NAND2_X1 U11485 ( .A1(n10803), .A2(n19984), .ZN(n11155) );
  CLKBUF_X1 U11486 ( .A(n12403), .Z(n12455) );
  NAND2_X1 U11487 ( .A1(n11934), .A2(n11933), .ZN(n11942) );
  AND3_X1 U11488 ( .A1(n11752), .A2(n13777), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12543) );
  NAND2_X1 U11489 ( .A1(n10830), .A2(n10799), .ZN(n9790) );
  INV_X1 U11490 ( .A(n11543), .ZN(n9955) );
  OAI21_X1 U11491 ( .B1(n10809), .B2(n10808), .A(n10807), .ZN(n10811) );
  NAND2_X1 U11492 ( .A1(n10803), .A2(n16914), .ZN(n10810) );
  NAND2_X1 U11493 ( .A1(n9779), .A2(n9778), .ZN(n10783) );
  OAI21_X1 U11494 ( .B1(n10729), .B2(n10730), .A(n10750), .ZN(n9779) );
  NAND2_X1 U11495 ( .A1(n14772), .A2(n10453), .ZN(n10452) );
  INV_X1 U11496 ( .A(n14785), .ZN(n10453) );
  INV_X1 U11497 ( .A(n14827), .ZN(n10446) );
  INV_X1 U11498 ( .A(n11935), .ZN(n12505) );
  NOR2_X1 U11499 ( .A1(n15374), .A2(n10006), .ZN(n10005) );
  INV_X1 U11500 ( .A(n12779), .ZN(n10006) );
  NAND2_X1 U11501 ( .A1(n12781), .A2(n15430), .ZN(n12780) );
  OR2_X1 U11502 ( .A1(n12784), .A2(n15207), .ZN(n12782) );
  NAND2_X1 U11503 ( .A1(n12776), .A2(n10285), .ZN(n10284) );
  OR2_X1 U11504 ( .A1(n12709), .A2(n12704), .ZN(n10283) );
  OAI21_X1 U11505 ( .B1(n12755), .B2(n12754), .A(n12761), .ZN(n12762) );
  OAI211_X1 U11506 ( .C1(n10445), .C2(n9991), .A(n12750), .B(n9989), .ZN(
        n12752) );
  NAND2_X1 U11507 ( .A1(n9995), .A2(n12960), .ZN(n9991) );
  NAND2_X1 U11508 ( .A1(n10159), .A2(n12744), .ZN(n12745) );
  INV_X1 U11509 ( .A(n13760), .ZN(n11828) );
  AND2_X1 U11510 ( .A1(n11717), .A2(n9985), .ZN(n9984) );
  NAND2_X1 U11511 ( .A1(n11714), .A2(n13519), .ZN(n9985) );
  OAI211_X1 U11512 ( .C1(n13845), .C2(n13622), .A(n15020), .B(n10160), .ZN(
        n10161) );
  OR2_X1 U11513 ( .A1(n12804), .A2(n13839), .ZN(n10160) );
  NAND2_X1 U11514 ( .A1(n11818), .A2(n11817), .ZN(n11823) );
  NAND2_X1 U11515 ( .A1(n12120), .A2(n11699), .ZN(n11704) );
  INV_X1 U11516 ( .A(n11011), .ZN(n10473) );
  NOR2_X1 U11517 ( .A1(n11012), .A2(n11009), .ZN(n10472) );
  NAND2_X1 U11518 ( .A1(n10017), .A2(n10015), .ZN(n10955) );
  INV_X1 U11519 ( .A(n10959), .ZN(n10017) );
  MUX2_X1 U11520 ( .A(n13773), .B(n11130), .S(n10787), .Z(n10963) );
  NAND2_X1 U11521 ( .A1(n13868), .A2(n13869), .ZN(n14062) );
  INV_X1 U11522 ( .A(n10834), .ZN(n10833) );
  NOR2_X1 U11523 ( .A1(n15873), .A2(n10521), .ZN(n10520) );
  INV_X1 U11524 ( .A(n15862), .ZN(n10521) );
  NAND2_X1 U11525 ( .A1(n10507), .A2(n10506), .ZN(n10505) );
  INV_X1 U11526 ( .A(n13783), .ZN(n10506) );
  INV_X1 U11527 ( .A(n13756), .ZN(n10507) );
  INV_X1 U11528 ( .A(n10499), .ZN(n10498) );
  OAI21_X1 U11529 ( .B1(n13567), .B2(n11333), .A(n13595), .ZN(n10499) );
  AND2_X1 U11530 ( .A1(n13602), .A2(n13585), .ZN(n14625) );
  AND2_X1 U11531 ( .A1(n19972), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13602) );
  NAND4_X1 U11532 ( .A1(n10032), .A2(n10860), .A3(n10061), .A4(n9834), .ZN(
        n10846) );
  AND2_X1 U11533 ( .A1(n10842), .A2(n10033), .ZN(n10032) );
  AND3_X1 U11534 ( .A1(n15821), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n11096), .ZN(n14315) );
  AND2_X1 U11535 ( .A1(n10953), .A2(n10952), .ZN(n10954) );
  OAI21_X1 U11536 ( .B1(n9769), .B2(n10983), .A(n10982), .ZN(n9831) );
  AOI22_X1 U11537 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n16877), .B1(
        n10921), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10916) );
  NAND2_X1 U11538 ( .A1(n10650), .A2(n10649), .ZN(n10961) );
  INV_X1 U11539 ( .A(n10809), .ZN(n10791) );
  AND2_X1 U11540 ( .A1(n14062), .A2(n13925), .ZN(n13872) );
  NAND2_X1 U11541 ( .A1(n9927), .A2(n13766), .ZN(n10873) );
  NOR2_X1 U11542 ( .A1(n11485), .A2(n11484), .ZN(n16926) );
  OAI21_X1 U11543 ( .B1(n13276), .B2(n19066), .A(n10204), .ZN(n13286) );
  NOR2_X1 U11544 ( .A1(n10205), .A2(n9678), .ZN(n10204) );
  INV_X1 U11545 ( .A(n19529), .ZN(n17061) );
  AND2_X2 U11546 ( .A1(n14757), .A2(n12810), .ZN(n20784) );
  AND2_X1 U11547 ( .A1(n12832), .A2(n12943), .ZN(n13750) );
  AND2_X1 U11548 ( .A1(n11830), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12510) );
  AND4_X1 U11549 ( .A1(n11678), .A2(n11677), .A3(n11676), .A4(n11675), .ZN(
        n11679) );
  NAND2_X1 U11550 ( .A1(n12276), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12342) );
  AND2_X1 U11551 ( .A1(n14873), .A2(n12216), .ZN(n14861) );
  NOR2_X1 U11552 ( .A1(n12215), .A2(n12214), .ZN(n12216) );
  OR2_X1 U11553 ( .A1(n14875), .A2(n14902), .ZN(n12214) );
  INV_X1 U11554 ( .A(n14159), .ZN(n10095) );
  INV_X1 U11555 ( .A(n14098), .ZN(n10096) );
  INV_X1 U11556 ( .A(n10174), .ZN(n10112) );
  AND2_X2 U11557 ( .A1(n14853), .A2(n10434), .ZN(n14786) );
  AND2_X1 U11558 ( .A1(n9627), .A2(n14807), .ZN(n10434) );
  NAND2_X1 U11559 ( .A1(n10318), .A2(n9987), .ZN(n10317) );
  INV_X1 U11560 ( .A(n17179), .ZN(n9987) );
  NAND2_X1 U11561 ( .A1(n10165), .A2(n10318), .ZN(n10164) );
  NAND2_X1 U11562 ( .A1(n12973), .A2(n9907), .ZN(n13030) );
  OR2_X1 U11563 ( .A1(n17107), .A2(n9904), .ZN(n9907) );
  NAND2_X1 U11564 ( .A1(n9615), .A2(n9905), .ZN(n9904) );
  NAND2_X1 U11565 ( .A1(n13797), .A2(n11756), .ZN(n14113) );
  NAND3_X1 U11566 ( .A1(n11700), .A2(n17109), .A3(n11704), .ZN(n12566) );
  AND2_X1 U11567 ( .A1(n12804), .A2(n11703), .ZN(n11700) );
  AND2_X1 U11568 ( .A1(n10493), .A2(n10492), .ZN(n10491) );
  INV_X1 U11569 ( .A(n15825), .ZN(n10492) );
  INV_X1 U11570 ( .A(n10026), .ZN(n10020) );
  AND2_X1 U11571 ( .A1(n16347), .A2(n16346), .ZN(n16369) );
  NAND2_X1 U11572 ( .A1(n14360), .A2(n11547), .ZN(n16353) );
  NAND2_X1 U11573 ( .A1(n11061), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16418) );
  INV_X1 U11574 ( .A(n10221), .ZN(n10013) );
  AND2_X1 U11575 ( .A1(n10292), .A2(n14350), .ZN(n10014) );
  NAND2_X1 U11576 ( .A1(n14360), .A2(n9762), .ZN(n16443) );
  AND4_X1 U11577 ( .A1(n10708), .A2(n10707), .A3(n10706), .A4(n10705), .ZN(
        n10714) );
  AND4_X1 U11578 ( .A1(n10712), .A2(n10711), .A3(n10710), .A4(n10709), .ZN(
        n10713) );
  NOR2_X1 U11579 ( .A1(n10704), .A2(n10703), .ZN(n10715) );
  NAND2_X1 U11580 ( .A1(n11479), .A2(n9804), .ZN(n16818) );
  INV_X1 U11581 ( .A(n9861), .ZN(n13475) );
  AND2_X1 U11582 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20313) );
  NAND2_X1 U11583 ( .A1(n19529), .A2(n10258), .ZN(n10257) );
  INV_X1 U11584 ( .A(n17060), .ZN(n10258) );
  OAI21_X1 U11585 ( .B1(n17133), .B2(n10142), .A(n13159), .ZN(n13160) );
  INV_X1 U11586 ( .A(n13158), .ZN(n10230) );
  NAND2_X1 U11587 ( .A1(n10229), .A2(n10227), .ZN(n10231) );
  INV_X1 U11588 ( .A(n13157), .ZN(n17133) );
  NOR2_X2 U11589 ( .A1(n18392), .A2(n10303), .ZN(n13151) );
  NAND2_X1 U11590 ( .A1(n10534), .A2(n10535), .ZN(n10303) );
  NAND2_X1 U11591 ( .A1(n19066), .A2(n19062), .ZN(n19482) );
  INV_X1 U11592 ( .A(n12952), .ZN(n10048) );
  AND2_X1 U11593 ( .A1(n12599), .A2(n19716), .ZN(n20682) );
  NAND2_X1 U11594 ( .A1(n9810), .A2(n9809), .ZN(n16690) );
  AOI21_X1 U11595 ( .B1(n9583), .B2(n9883), .A(n9690), .ZN(n9882) );
  NOR2_X1 U11596 ( .A1(n19970), .A2(n9891), .ZN(n9883) );
  NOR2_X1 U11597 ( .A1(n9958), .A2(n9957), .ZN(n9956) );
  INV_X1 U11598 ( .A(n14728), .ZN(n9958) );
  NOR2_X1 U11599 ( .A1(n16123), .A2(n16782), .ZN(n9957) );
  AOI21_X1 U11600 ( .B1(n12541), .B2(n12540), .A(n12539), .ZN(n12549) );
  INV_X1 U11601 ( .A(n11731), .ZN(n12452) );
  NAND2_X1 U11602 ( .A1(n20651), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10645) );
  NOR2_X1 U11603 ( .A1(n11166), .A2(n20567), .ZN(n9859) );
  AND2_X1 U11604 ( .A1(n10783), .A2(n10786), .ZN(n11160) );
  NAND2_X1 U11605 ( .A1(n13475), .A2(n12597), .ZN(n9862) );
  NOR2_X1 U11606 ( .A1(n13168), .A2(n13167), .ZN(n13164) );
  OAI21_X1 U11607 ( .B1(n9902), .B2(n9607), .A(n9895), .ZN(n9894) );
  AND2_X1 U11608 ( .A1(n9893), .A2(n12532), .ZN(n9892) );
  INV_X1 U11609 ( .A(n12538), .ZN(n9893) );
  INV_X1 U11610 ( .A(n13829), .ZN(n9903) );
  AND2_X1 U11611 ( .A1(n9655), .A2(n10120), .ZN(n10119) );
  NAND2_X1 U11612 ( .A1(n15374), .A2(n12778), .ZN(n10120) );
  AND2_X1 U11613 ( .A1(n15383), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12776) );
  INV_X1 U11614 ( .A(n11960), .ZN(n11958) );
  OR2_X1 U11615 ( .A1(n11956), .A2(n11955), .ZN(n12758) );
  INV_X1 U11616 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9981) );
  XNOR2_X1 U11617 ( .A(n10750), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10667) );
  NOR2_X1 U11618 ( .A1(n12672), .A2(n20690), .ZN(n10799) );
  AOI21_X1 U11619 ( .B1(n10834), .B2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n10796), .ZN(n10816) );
  NAND2_X1 U11620 ( .A1(n9842), .A2(n9837), .ZN(n10796) );
  NAND2_X1 U11621 ( .A1(n9841), .A2(n9839), .ZN(n9842) );
  AOI21_X1 U11622 ( .B1(n9613), .B2(n11169), .A(n9739), .ZN(n9837) );
  NOR2_X1 U11623 ( .A1(n14355), .A2(n14353), .ZN(n14354) );
  XNOR2_X1 U11624 ( .A(n10644), .B(n10642), .ZN(n11144) );
  NAND2_X1 U11625 ( .A1(n10524), .A2(n10523), .ZN(n11157) );
  NAND2_X1 U11626 ( .A1(n10059), .A2(n10058), .ZN(n11172) );
  NAND2_X1 U11627 ( .A1(n20690), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10058) );
  NAND2_X1 U11628 ( .A1(n11123), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10059) );
  OAI21_X1 U11629 ( .B1(n13183), .B2(n18061), .A(n13185), .ZN(n13186) );
  NOR2_X1 U11630 ( .A1(n17400), .A2(n13270), .ZN(n17065) );
  INV_X1 U11631 ( .A(n19500), .ZN(n9939) );
  INV_X1 U11632 ( .A(n19070), .ZN(n13278) );
  NAND2_X1 U11633 ( .A1(n11701), .A2(n11696), .ZN(n11698) );
  NAND2_X1 U11634 ( .A1(n12575), .A2(n11829), .ZN(n11701) );
  INV_X1 U11635 ( .A(n14805), .ZN(n10098) );
  NOR2_X1 U11636 ( .A1(n14851), .A2(n10448), .ZN(n10447) );
  INV_X1 U11637 ( .A(n14862), .ZN(n10448) );
  INV_X1 U11638 ( .A(n12471), .ZN(n12507) );
  AND2_X1 U11639 ( .A1(n12092), .A2(n10440), .ZN(n10439) );
  NAND2_X1 U11640 ( .A1(n10441), .A2(n12054), .ZN(n10440) );
  INV_X1 U11641 ( .A(n10442), .ZN(n10441) );
  AND2_X1 U11642 ( .A1(n10443), .A2(n14280), .ZN(n10442) );
  INV_X1 U11643 ( .A(n14271), .ZN(n10443) );
  NOR2_X1 U11644 ( .A1(n14258), .A2(n14263), .ZN(n11993) );
  NOR2_X1 U11645 ( .A1(n14260), .A2(n10425), .ZN(n10424) );
  INV_X1 U11646 ( .A(n14266), .ZN(n10425) );
  INV_X1 U11647 ( .A(n14259), .ZN(n10423) );
  NAND2_X1 U11648 ( .A1(n21470), .A2(n12943), .ZN(n12897) );
  NAND2_X1 U11649 ( .A1(n9875), .A2(n12712), .ZN(n12736) );
  INV_X1 U11650 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11594) );
  OR2_X1 U11651 ( .A1(n11810), .A2(n11809), .ZN(n12720) );
  NOR2_X1 U11652 ( .A1(n13818), .A2(n12915), .ZN(n10117) );
  INV_X1 U11653 ( .A(n15646), .ZN(n14121) );
  NAND2_X1 U11654 ( .A1(n13938), .A2(n11759), .ZN(n10102) );
  AND2_X2 U11655 ( .A1(n10794), .A2(n10782), .ZN(n10808) );
  OR2_X1 U11656 ( .A1(n10573), .A2(n10572), .ZN(n10902) );
  INV_X1 U11657 ( .A(n10248), .ZN(n10247) );
  OAI21_X1 U11658 ( .B1(n10245), .B2(n9718), .A(n10249), .ZN(n10248) );
  INV_X1 U11659 ( .A(n16341), .ZN(n10249) );
  NOR2_X1 U11660 ( .A1(n12602), .A2(n10399), .ZN(n10398) );
  OR2_X1 U11661 ( .A1(n11022), .A2(n11023), .ZN(n11025) );
  AND2_X1 U11662 ( .A1(n9626), .A2(n16102), .ZN(n10462) );
  NAND2_X1 U11663 ( .A1(n10513), .A2(n16257), .ZN(n10512) );
  INV_X1 U11664 ( .A(n10514), .ZN(n10513) );
  NAND2_X1 U11665 ( .A1(n16925), .A2(n19972), .ZN(n11173) );
  INV_X1 U11666 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10389) );
  NOR2_X1 U11667 ( .A1(n11088), .A2(n10025), .ZN(n10024) );
  INV_X1 U11668 ( .A(n16344), .ZN(n10025) );
  AND2_X1 U11669 ( .A1(n15851), .A2(n11096), .ZN(n11072) );
  INV_X1 U11670 ( .A(n15839), .ZN(n10518) );
  OR2_X1 U11671 ( .A1(n13677), .A2(n13756), .ZN(n13754) );
  NAND2_X1 U11672 ( .A1(n9815), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9814) );
  INV_X1 U11673 ( .A(n16498), .ZN(n9815) );
  NAND2_X1 U11674 ( .A1(n9819), .A2(n19861), .ZN(n9818) );
  NAND2_X1 U11675 ( .A1(n9969), .A2(n11542), .ZN(n9819) );
  NAND3_X1 U11676 ( .A1(n9969), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n11543), .ZN(n11522) );
  NAND2_X1 U11677 ( .A1(n16804), .A2(n16792), .ZN(n11536) );
  NOR2_X1 U11678 ( .A1(n10684), .A2(n10683), .ZN(n11327) );
  INV_X1 U11679 ( .A(n10212), .ZN(n9962) );
  NOR2_X1 U11680 ( .A1(n9728), .A2(n11096), .ZN(n9920) );
  INV_X1 U11681 ( .A(n16003), .ZN(n10286) );
  INV_X1 U11682 ( .A(n13768), .ZN(n13767) );
  NAND2_X1 U11683 ( .A1(n20688), .A2(n10803), .ZN(n11486) );
  AOI21_X1 U11684 ( .B1(n16819), .B2(n11489), .A(n10788), .ZN(n11496) );
  NAND2_X1 U11685 ( .A1(n10813), .A2(n9863), .ZN(n11492) );
  NAND2_X1 U11686 ( .A1(n10804), .A2(n10788), .ZN(n10798) );
  NAND2_X1 U11687 ( .A1(n11488), .A2(n16914), .ZN(n9791) );
  AND2_X1 U11688 ( .A1(n13766), .A2(n16831), .ZN(n10552) );
  AOI22_X1 U11689 ( .A1(n14516), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10776) );
  NAND2_X1 U11690 ( .A1(n18018), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10261) );
  NOR2_X1 U11691 ( .A1(n17458), .A2(n18362), .ZN(n10326) );
  NOR2_X1 U11692 ( .A1(n13043), .A2(n17789), .ZN(n13061) );
  NOR2_X1 U11693 ( .A1(n18524), .A2(n10345), .ZN(n10344) );
  INV_X1 U11694 ( .A(n18522), .ZN(n10343) );
  NAND2_X1 U11695 ( .A1(n10140), .A2(n18734), .ZN(n10139) );
  NOR2_X1 U11696 ( .A1(n18634), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10140) );
  NAND2_X1 U11697 ( .A1(n18634), .A2(n18856), .ZN(n13145) );
  AND2_X1 U11698 ( .A1(n18596), .A2(n9603), .ZN(n10042) );
  NOR2_X1 U11699 ( .A1(n17062), .A2(n17065), .ZN(n17415) );
  NAND2_X1 U11700 ( .A1(n13138), .A2(n13300), .ZN(n17288) );
  INV_X1 U11701 ( .A(n13322), .ZN(n10082) );
  NAND2_X1 U11702 ( .A1(n18649), .A2(n13127), .ZN(n13140) );
  NAND2_X1 U11703 ( .A1(n18665), .A2(n13314), .ZN(n13316) );
  NAND2_X1 U11704 ( .A1(n18687), .A2(n13090), .ZN(n13103) );
  XNOR2_X1 U11705 ( .A(n13306), .B(n10072), .ZN(n13307) );
  INV_X1 U11706 ( .A(n18236), .ZN(n10072) );
  XNOR2_X1 U11707 ( .A(n13101), .B(n13102), .ZN(n13089) );
  NAND2_X1 U11708 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10200) );
  NOR2_X1 U11709 ( .A1(n13183), .A2(n17829), .ZN(n10198) );
  NAND2_X1 U11710 ( .A1(n20783), .A2(n9758), .ZN(n20773) );
  AND2_X1 U11711 ( .A1(n12823), .A2(n12822), .ZN(n13787) );
  NAND2_X1 U11712 ( .A1(n12559), .A2(n12558), .ZN(n12560) );
  AND4_X1 U11713 ( .A1(n11688), .A2(n11687), .A3(n11686), .A4(n11685), .ZN(
        n11693) );
  AND4_X1 U11714 ( .A1(n11684), .A2(n11683), .A3(n11682), .A4(n11681), .ZN(
        n11694) );
  INV_X1 U11715 ( .A(n10451), .ZN(n10449) );
  OR2_X1 U11716 ( .A1(n14784), .A2(n10452), .ZN(n14771) );
  NAND2_X1 U11717 ( .A1(n12391), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12441) );
  OAI21_X1 U11718 ( .B1(n15230), .B2(n12503), .A(n12315), .ZN(n14827) );
  NAND2_X1 U11719 ( .A1(n12116), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12234) );
  NAND2_X1 U11720 ( .A1(n12115), .A2(n12114), .ZN(n12195) );
  AND2_X1 U11721 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12114) );
  INV_X1 U11722 ( .A(n12156), .ZN(n12115) );
  INV_X1 U11723 ( .A(n12073), .ZN(n12094) );
  INV_X1 U11724 ( .A(n14097), .ZN(n10094) );
  AOI21_X1 U11725 ( .B1(n12747), .B2(n12107), .A(n11941), .ZN(n14159) );
  OAI211_X1 U11726 ( .C1(n10445), .C2(n9998), .A(n9997), .B(n9992), .ZN(n12747) );
  AOI21_X1 U11727 ( .B1(n12738), .B2(n12107), .A(n11916), .ZN(n14098) );
  NAND2_X1 U11728 ( .A1(n11856), .A2(n11855), .ZN(n13974) );
  NAND2_X1 U11729 ( .A1(n10002), .A2(n10000), .ZN(n10070) );
  NAND2_X1 U11730 ( .A1(n10001), .A2(n13020), .ZN(n10000) );
  NAND2_X1 U11731 ( .A1(n9912), .A2(n15422), .ZN(n15404) );
  OR2_X1 U11732 ( .A1(n13005), .A2(n15400), .ZN(n9912) );
  OR2_X1 U11733 ( .A1(n14773), .A2(n14776), .ZN(n14774) );
  NAND2_X1 U11734 ( .A1(n15237), .A2(n10005), .ZN(n9999) );
  NAND2_X1 U11735 ( .A1(n10118), .A2(n15353), .ZN(n10004) );
  NOR2_X1 U11736 ( .A1(n15447), .A2(n13003), .ZN(n15428) );
  AND2_X2 U11737 ( .A1(n14868), .A2(n14855), .ZN(n14853) );
  INV_X1 U11738 ( .A(n14890), .ZN(n10430) );
  INV_X1 U11739 ( .A(n12777), .ZN(n15286) );
  INV_X1 U11740 ( .A(n14947), .ZN(n10432) );
  INV_X1 U11741 ( .A(n17171), .ZN(n9988) );
  XNOR2_X1 U11742 ( .A(n12762), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17171) );
  NAND2_X1 U11743 ( .A1(n17180), .A2(n17179), .ZN(n17178) );
  NOR3_X1 U11744 ( .A1(n17204), .A2(n10429), .A3(n14045), .ZN(n10426) );
  OR2_X1 U11745 ( .A1(n14046), .A2(n10428), .ZN(n17203) );
  XNOR2_X1 U11746 ( .A(n12745), .B(n20900), .ZN(n20858) );
  INV_X1 U11747 ( .A(n13030), .ZN(n9906) );
  AND2_X1 U11748 ( .A1(n13030), .A2(n17101), .ZN(n20891) );
  NOR2_X1 U11749 ( .A1(n10170), .A2(n9665), .ZN(n10169) );
  NAND2_X1 U11750 ( .A1(n14755), .A2(n11715), .ZN(n9983) );
  INV_X1 U11751 ( .A(n10124), .ZN(n12713) );
  OAI21_X1 U11752 ( .B1(n14113), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11779), 
        .ZN(n10124) );
  XNOR2_X1 U11753 ( .A(n11823), .B(n11821), .ZN(n11836) );
  INV_X1 U11754 ( .A(n14077), .ZN(n14066) );
  OAI21_X1 U11755 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n21064), .A(
        n14121), .ZN(n14071) );
  AND2_X1 U11756 ( .A1(n15658), .A2(n14006), .ZN(n14077) );
  OR2_X1 U11757 ( .A1(n14006), .A2(n11880), .ZN(n15659) );
  AND2_X1 U11758 ( .A1(n14014), .A2(n15640), .ZN(n15679) );
  INV_X1 U11759 ( .A(n14220), .ZN(n20993) );
  NOR2_X1 U11760 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21029) );
  OR2_X1 U11761 ( .A1(n15658), .A2(n15653), .ZN(n21031) );
  INV_X1 U11762 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n14084) );
  OR2_X1 U11763 ( .A1(n14014), .A2(n15640), .ZN(n14089) );
  OR2_X1 U11764 ( .A1(n14014), .A2(n14013), .ZN(n14088) );
  NOR2_X1 U11765 ( .A1(n15683), .A2(n15646), .ZN(n21098) );
  INV_X1 U11766 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21136) );
  NAND2_X1 U11767 ( .A1(n11759), .A2(n13807), .ZN(n15646) );
  OR2_X1 U11768 ( .A1(n14006), .A2(n14005), .ZN(n21140) );
  INV_X1 U11769 ( .A(n14071), .ZN(n21147) );
  NAND2_X1 U11770 ( .A1(n10785), .A2(n12597), .ZN(n10790) );
  NAND2_X1 U11771 ( .A1(n16825), .A2(n20690), .ZN(n20681) );
  INV_X1 U11772 ( .A(n11081), .ZN(n11099) );
  NOR2_X1 U11773 ( .A1(n11042), .A2(n10477), .ZN(n10476) );
  NOR2_X1 U11774 ( .A1(n15879), .A2(n10384), .ZN(n10380) );
  NOR2_X1 U11775 ( .A1(n10471), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10470) );
  OR2_X1 U11776 ( .A1(n10019), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10018) );
  NAND2_X1 U11777 ( .A1(n19787), .A2(n12637), .ZN(n19773) );
  NOR2_X1 U11778 ( .A1(n19989), .A2(n10718), .ZN(n11027) );
  AND2_X1 U11779 ( .A1(n19829), .A2(n9628), .ZN(n15930) );
  NAND2_X1 U11780 ( .A1(n10401), .A2(n10403), .ZN(n12617) );
  INV_X1 U11781 ( .A(n12618), .ZN(n10401) );
  AND2_X1 U11782 ( .A1(n19837), .A2(n19817), .ZN(n10480) );
  NAND2_X1 U11783 ( .A1(n19845), .A2(n19848), .ZN(n15952) );
  NAND2_X1 U11784 ( .A1(n10652), .A2(n10651), .ZN(n10959) );
  INV_X1 U11785 ( .A(n10961), .ZN(n10651) );
  CLKBUF_X1 U11786 ( .A(n10955), .Z(n10976) );
  AND2_X1 U11787 ( .A1(n11147), .A2(n11146), .ZN(n16931) );
  OR2_X1 U11788 ( .A1(n11145), .A2(n11148), .ZN(n11146) );
  NAND2_X1 U11789 ( .A1(n15800), .A2(n9724), .ZN(n15775) );
  NAND2_X1 U11790 ( .A1(n14062), .A2(n14061), .ZN(n10459) );
  INV_X1 U11791 ( .A(n14429), .ZN(n10461) );
  INV_X1 U11792 ( .A(n14181), .ZN(n14184) );
  OR2_X1 U11793 ( .A1(n13677), .A2(n10505), .ZN(n13879) );
  NAND2_X1 U11794 ( .A1(n10504), .A2(n10503), .ZN(n10502) );
  INV_X1 U11795 ( .A(n13878), .ZN(n10503) );
  INV_X1 U11796 ( .A(n10505), .ZN(n10504) );
  AND3_X1 U11797 ( .A1(n11349), .A2(n11348), .A3(n11347), .ZN(n13679) );
  CLKBUF_X1 U11798 ( .A(n13593), .Z(n13594) );
  INV_X1 U11799 ( .A(n10786), .ZN(n9832) );
  AND2_X1 U11800 ( .A1(n13927), .A2(n13926), .ZN(n14104) );
  NAND2_X1 U11801 ( .A1(n9695), .A2(n11288), .ZN(n11289) );
  OR2_X1 U11802 ( .A1(n12651), .A2(n12603), .ZN(n12653) );
  OR2_X1 U11803 ( .A1(n12649), .A2(n16338), .ZN(n12651) );
  CLKBUF_X1 U11804 ( .A(n15867), .Z(n15868) );
  OR2_X1 U11805 ( .A1(n12632), .A2(n15921), .ZN(n12636) );
  NOR2_X1 U11806 ( .A1(n12636), .A2(n19793), .ZN(n12635) );
  INV_X1 U11807 ( .A(n10843), .ZN(n10844) );
  AND2_X1 U11808 ( .A1(n10847), .A2(n10842), .ZN(n10845) );
  AND2_X1 U11809 ( .A1(n9724), .A2(n10489), .ZN(n10488) );
  INV_X1 U11810 ( .A(n15776), .ZN(n10489) );
  NOR2_X1 U11811 ( .A1(n16568), .A2(n16570), .ZN(n16554) );
  NAND2_X1 U11812 ( .A1(n9852), .A2(n9849), .ZN(n9850) );
  NOR2_X1 U11813 ( .A1(n10528), .A2(n11548), .ZN(n9849) );
  NAND2_X1 U11814 ( .A1(n9852), .A2(n9761), .ZN(n16313) );
  AND2_X1 U11815 ( .A1(n16738), .A2(n11547), .ZN(n16623) );
  NAND2_X1 U11816 ( .A1(n10218), .A2(n16388), .ZN(n10217) );
  NAND2_X1 U11817 ( .A1(n14359), .A2(n14358), .ZN(n10216) );
  OR2_X1 U11818 ( .A1(n11064), .A2(n16650), .ZN(n16389) );
  NAND2_X1 U11819 ( .A1(n9816), .A2(n14357), .ZN(n16391) );
  OAI211_X1 U11820 ( .C1(n10007), .C2(n9968), .A(n9817), .B(n9616), .ZN(n9816)
         );
  NAND2_X1 U11821 ( .A1(n10482), .A2(n9676), .ZN(n10481) );
  INV_X1 U11822 ( .A(n10483), .ZN(n10482) );
  NAND2_X1 U11823 ( .A1(n16476), .A2(n10376), .ZN(n9809) );
  NAND2_X1 U11824 ( .A1(n14360), .A2(n9915), .ZN(n9914) );
  NOR2_X1 U11825 ( .A1(n16465), .A2(n16739), .ZN(n9915) );
  AND2_X1 U11826 ( .A1(n11198), .A2(n9610), .ZN(n16148) );
  INV_X1 U11827 ( .A(n15982), .ZN(n10501) );
  NAND2_X1 U11828 ( .A1(n10983), .A2(n10147), .ZN(n10146) );
  INV_X1 U11829 ( .A(n9831), .ZN(n9830) );
  NAND2_X1 U11830 ( .A1(n10957), .A2(n10958), .ZN(n9949) );
  NAND2_X1 U11831 ( .A1(n11501), .A2(n13654), .ZN(n10057) );
  NAND2_X1 U11832 ( .A1(n13582), .A2(n20276), .ZN(n13865) );
  CLKBUF_X1 U11833 ( .A(n11137), .Z(n11138) );
  OR3_X1 U11834 ( .A1(n20008), .A2(n20028), .A3(n20463), .ZN(n20011) );
  NAND2_X1 U11835 ( .A1(n10861), .A2(n10868), .ZN(n9798) );
  NAND2_X1 U11836 ( .A1(n10868), .A2(n9927), .ZN(n9796) );
  NOR2_X1 U11837 ( .A1(n20315), .A2(n20314), .ZN(n20319) );
  NAND2_X2 U11838 ( .A1(n10861), .A2(n10552), .ZN(n9866) );
  NAND2_X1 U11839 ( .A1(n20647), .A2(n20655), .ZN(n20114) );
  AND2_X1 U11840 ( .A1(n20637), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20472) );
  NAND2_X1 U11841 ( .A1(n13546), .A2(n13545), .ZN(n20476) );
  OR2_X1 U11842 ( .A1(n20695), .A2(n13544), .ZN(n13545) );
  NAND2_X1 U11843 ( .A1(n17251), .A2(n20690), .ZN(n13546) );
  INV_X1 U11844 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20463) );
  NOR2_X1 U11845 ( .A1(n17456), .A2(n17653), .ZN(n17451) );
  NAND2_X1 U11846 ( .A1(n17468), .A2(n17847), .ZN(n17450) );
  NOR2_X1 U11847 ( .A1(n18464), .A2(n18451), .ZN(n10332) );
  OR2_X1 U11848 ( .A1(n18375), .A2(n10346), .ZN(n13331) );
  OR2_X1 U11849 ( .A1(n10348), .A2(n10347), .ZN(n10346) );
  NAND2_X1 U11850 ( .A1(n19710), .A2(n17743), .ZN(n17421) );
  NOR2_X1 U11851 ( .A1(n17924), .A2(n10267), .ZN(n10265) );
  INV_X1 U11852 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n10267) );
  NOR2_X1 U11853 ( .A1(n18109), .A2(n10211), .ZN(n10210) );
  AND2_X1 U11854 ( .A1(n18389), .A2(n18369), .ZN(n18370) );
  NAND2_X1 U11855 ( .A1(n13327), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13328) );
  NOR2_X1 U11856 ( .A1(n18652), .A2(n10337), .ZN(n10340) );
  INV_X1 U11857 ( .A(n18859), .ZN(n18786) );
  NAND2_X1 U11858 ( .A1(n18513), .A2(n18839), .ZN(n18514) );
  OAI22_X1 U11859 ( .A1(n18786), .A2(n19527), .B1(n18860), .B2(n18910), .ZN(
        n18801) );
  NAND2_X1 U11860 ( .A1(n18655), .A2(n13317), .ZN(n18642) );
  XNOR2_X1 U11861 ( .A(n13316), .B(n10153), .ZN(n18656) );
  INV_X1 U11862 ( .A(n13315), .ZN(n10153) );
  NAND2_X1 U11863 ( .A1(n18656), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18655) );
  XNOR2_X1 U11864 ( .A(n13103), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18680) );
  OR2_X1 U11865 ( .A1(n21354), .A2(n13074), .ZN(n13075) );
  INV_X1 U11866 ( .A(n13288), .ZN(n13287) );
  NAND2_X1 U11867 ( .A1(n19501), .A2(n9940), .ZN(n19502) );
  NAND2_X1 U11868 ( .A1(n19499), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9940) );
  NOR2_X2 U11869 ( .A1(n19711), .A2(n17060), .ZN(n19512) );
  OAI211_X1 U11870 ( .C1(n9666), .C2(n19516), .A(n9946), .B(n9944), .ZN(n9943)
         );
  AOI21_X1 U11871 ( .B1(n19519), .B2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n9946) );
  NAND2_X1 U11872 ( .A1(n9945), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n9944) );
  OR2_X1 U11873 ( .A1(n12953), .A2(n21276), .ZN(n10049) );
  AND2_X1 U11874 ( .A1(n14835), .A2(n12936), .ZN(n14800) );
  INV_X1 U11875 ( .A(n12913), .ZN(n12811) );
  XNOR2_X1 U11876 ( .A(n9639), .B(n12513), .ZN(n12955) );
  INV_X1 U11877 ( .A(n15170), .ZN(n15077) );
  OR2_X1 U11878 ( .A1(n13638), .A2(n12577), .ZN(n12578) );
  NAND2_X1 U11879 ( .A1(n10112), .A2(n10176), .ZN(n10175) );
  AND2_X1 U11880 ( .A1(n12783), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10176) );
  NAND2_X1 U11881 ( .A1(n10181), .A2(n10178), .ZN(n10177) );
  OR2_X1 U11882 ( .A1(n12787), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10181) );
  NAND2_X1 U11883 ( .A1(n12787), .A2(n10179), .ZN(n10178) );
  NAND2_X1 U11884 ( .A1(n10180), .A2(n13019), .ZN(n10179) );
  XNOR2_X1 U11885 ( .A(n12950), .B(n12949), .ZN(n15043) );
  NAND2_X1 U11886 ( .A1(n12947), .A2(n12946), .ZN(n12950) );
  OR2_X1 U11887 ( .A1(n15404), .A2(n9910), .ZN(n9909) );
  INV_X1 U11888 ( .A(n9911), .ZN(n9910) );
  AOI21_X1 U11889 ( .B1(n15521), .B2(n21452), .A(n13006), .ZN(n9911) );
  XNOR2_X1 U11890 ( .A(n10420), .B(n12945), .ZN(n15397) );
  NAND2_X1 U11891 ( .A1(n9650), .A2(n10418), .ZN(n10420) );
  OAI21_X1 U11892 ( .B1(n14773), .B2(n10419), .A(n12944), .ZN(n10418) );
  OAI21_X1 U11893 ( .B1(n15189), .B2(n10541), .A(n10319), .ZN(n15165) );
  NAND2_X1 U11894 ( .A1(n10174), .A2(n10320), .ZN(n10319) );
  XNOR2_X1 U11895 ( .A(n9722), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10276) );
  INV_X1 U11896 ( .A(n15409), .ZN(n10277) );
  NAND2_X1 U11897 ( .A1(n12998), .A2(n15474), .ZN(n15459) );
  AND2_X1 U11898 ( .A1(n10314), .A2(n12566), .ZN(n13028) );
  NAND2_X1 U11899 ( .A1(n14007), .A2(n21057), .ZN(n21145) );
  OR2_X1 U11900 ( .A1(n14014), .A2(n21141), .ZN(n14007) );
  NAND2_X1 U11901 ( .A1(n12668), .A2(n12669), .ZN(n10242) );
  NAND2_X1 U11902 ( .A1(n10245), .A2(n19875), .ZN(n19806) );
  NAND2_X1 U11903 ( .A1(n12690), .A2(n12689), .ZN(n12691) );
  AOI21_X1 U11904 ( .B1(n12688), .B2(n19832), .A(n12687), .ZN(n12689) );
  AOI21_X1 U11905 ( .B1(n16559), .B2(n19803), .A(n10414), .ZN(n10413) );
  NAND2_X1 U11906 ( .A1(n15784), .A2(n15785), .ZN(n10414) );
  AND2_X1 U11907 ( .A1(n19866), .A2(n19875), .ZN(n19810) );
  INV_X1 U11908 ( .A(n19870), .ZN(n19803) );
  INV_X1 U11909 ( .A(n19810), .ZN(n16046) );
  INV_X1 U11910 ( .A(n19860), .ZN(n19832) );
  NAND2_X1 U11911 ( .A1(n9602), .A2(n10456), .ZN(n14181) );
  NOR2_X1 U11912 ( .A1(n11400), .A2(n11399), .ZN(n14063) );
  XNOR2_X1 U11913 ( .A(n10840), .B(n11182), .ZN(n10841) );
  AND2_X1 U11914 ( .A1(n16287), .A2(n13574), .ZN(n16260) );
  XNOR2_X1 U11915 ( .A(n10030), .B(n16328), .ZN(n16586) );
  NAND2_X1 U11916 ( .A1(n10031), .A2(n16334), .ZN(n10030) );
  AND2_X1 U11917 ( .A1(n16312), .A2(n9848), .ZN(n9843) );
  AND2_X1 U11918 ( .A1(n9583), .A2(n19945), .ZN(n9774) );
  AOI21_X1 U11919 ( .B1(n16633), .B2(n16547), .A(n16375), .ZN(n10134) );
  INV_X1 U11920 ( .A(n16501), .ZN(n10105) );
  AND2_X1 U11921 ( .A1(n19955), .A2(n14341), .ZN(n19943) );
  INV_X1 U11922 ( .A(n19943), .ZN(n16544) );
  INV_X1 U11923 ( .A(n19955), .ZN(n16510) );
  NAND3_X1 U11924 ( .A1(n20634), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20476), 
        .ZN(n19950) );
  NAND2_X1 U11925 ( .A1(n10354), .A2(n10353), .ZN(n10352) );
  NAND2_X1 U11926 ( .A1(n11102), .A2(n10361), .ZN(n10353) );
  OAI21_X1 U11927 ( .B1(n10358), .B2(n10362), .A(n10355), .ZN(n10354) );
  NAND2_X1 U11928 ( .A1(n16292), .A2(n9667), .ZN(n10356) );
  NAND2_X1 U11929 ( .A1(n11074), .A2(n16344), .ZN(n9926) );
  NOR2_X1 U11930 ( .A1(n19970), .A2(n9846), .ZN(n9845) );
  INV_X1 U11931 ( .A(n9848), .ZN(n9846) );
  INV_X1 U11932 ( .A(n16586), .ZN(n10035) );
  NAND2_X1 U11933 ( .A1(n9583), .A2(n16579), .ZN(n9847) );
  OAI21_X1 U11934 ( .B1(n9636), .B2(n9887), .A(n9886), .ZN(n9885) );
  NAND2_X1 U11935 ( .A1(n16362), .A2(n9663), .ZN(n9775) );
  NOR2_X1 U11936 ( .A1(n16374), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16631) );
  NAND2_X1 U11937 ( .A1(n9855), .A2(n16353), .ZN(n16643) );
  NAND2_X1 U11938 ( .A1(n10008), .A2(n16637), .ZN(n9855) );
  NAND2_X1 U11939 ( .A1(n16662), .A2(n9960), .ZN(n9959) );
  AND2_X1 U11940 ( .A1(n14724), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9960) );
  NAND2_X1 U11941 ( .A1(n9966), .A2(n9729), .ZN(n9967) );
  AND2_X1 U11942 ( .A1(n16714), .A2(n16692), .ZN(n10045) );
  NAND2_X1 U11943 ( .A1(n9809), .A2(n16799), .ZN(n9808) );
  NAND2_X1 U11944 ( .A1(n10374), .A2(n10376), .ZN(n10373) );
  XNOR2_X1 U11945 ( .A(n10125), .B(n16419), .ZN(n16693) );
  NAND2_X1 U11946 ( .A1(n10417), .A2(n14352), .ZN(n10125) );
  NOR2_X1 U11947 ( .A1(n16476), .A2(n10374), .ZN(n16431) );
  INV_X1 U11948 ( .A(n10417), .ZN(n16424) );
  NAND2_X1 U11949 ( .A1(n9858), .A2(n16443), .ZN(n16711) );
  NAND2_X1 U11950 ( .A1(n10067), .A2(n16713), .ZN(n9858) );
  AND2_X1 U11951 ( .A1(n16714), .A2(n16713), .ZN(n10252) );
  AOI22_X1 U11952 ( .A1(n16437), .A2(n16451), .B1(n10012), .B2(n16447), .ZN(
        n16438) );
  INV_X1 U11953 ( .A(n16449), .ZN(n16437) );
  AND2_X1 U11954 ( .A1(n16762), .A2(n11545), .ZN(n16738) );
  NOR2_X1 U11955 ( .A1(n16499), .A2(n16500), .ZN(n16758) );
  AND2_X1 U11956 ( .A1(n16762), .A2(n16760), .ZN(n10128) );
  AND2_X1 U11957 ( .A1(n16499), .A2(n16500), .ZN(n16757) );
  NOR2_X1 U11958 ( .A1(n16789), .A2(n11512), .ZN(n16762) );
  NAND2_X1 U11959 ( .A1(n11551), .A2(n11483), .ZN(n17237) );
  NAND2_X1 U11960 ( .A1(n10822), .A2(n10137), .ZN(n10365) );
  NAND2_X1 U11961 ( .A1(n16818), .A2(n20688), .ZN(n10137) );
  INV_X1 U11962 ( .A(n19958), .ZN(n16802) );
  INV_X1 U11963 ( .A(n16782), .ZN(n19967) );
  INV_X1 U11964 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20667) );
  INV_X1 U11965 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20660) );
  INV_X1 U11966 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20651) );
  INV_X1 U11967 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20643) );
  INV_X1 U11968 ( .A(n20219), .ZN(n20216) );
  NOR2_X1 U11969 ( .A1(n20309), .A2(n20630), .ZN(n20350) );
  NOR4_X1 U11970 ( .A1(n16957), .A2(n16956), .A3(n20671), .A4(n16955), .ZN(
        n17255) );
  NAND4_X1 U11971 ( .A1(n19024), .A2(n19698), .A3(n19555), .A4(n19545), .ZN(
        n17801) );
  NOR2_X2 U11972 ( .A1(n13208), .A2(n13207), .ZN(n19084) );
  AND2_X1 U11973 ( .A1(n18140), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n18141) );
  NOR2_X2 U11974 ( .A1(n18113), .A2(n18177), .ZN(n18183) );
  NOR2_X1 U11975 ( .A1(n9629), .A2(n10209), .ZN(n10208) );
  NOR2_X1 U11976 ( .A1(n13137), .A2(n13136), .ZN(n18222) );
  NOR2_X1 U11977 ( .A1(n13113), .A2(n13112), .ZN(n18229) );
  INV_X1 U11978 ( .A(n18242), .ZN(n18248) );
  INV_X1 U11979 ( .A(n18248), .ZN(n18237) );
  NOR2_X2 U11980 ( .A1(n18222), .A2(n18724), .ZN(n18635) );
  OAI211_X1 U11981 ( .C1(n13156), .C2(n10036), .A(n13160), .B(n10037), .ZN(
        n13359) );
  NAND2_X1 U11982 ( .A1(n13158), .A2(n10038), .ZN(n10037) );
  NAND2_X1 U11983 ( .A1(n9664), .A2(n13158), .ZN(n10036) );
  NAND2_X2 U11984 ( .A1(n18929), .A2(n19494), .ZN(n18851) );
  INV_X1 U11985 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19517) );
  NAND2_X1 U11986 ( .A1(n12536), .A2(n12535), .ZN(n12541) );
  OAI21_X1 U11987 ( .B1(n12522), .B2(n9901), .A(n12523), .ZN(n9900) );
  NAND2_X1 U11988 ( .A1(n9903), .A2(n12567), .ZN(n9901) );
  INV_X1 U11989 ( .A(n11738), .ZN(n12317) );
  NAND2_X1 U11990 ( .A1(P2_EBX_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n9840) );
  NAND2_X1 U11991 ( .A1(n10645), .A2(n10602), .ZN(n10642) );
  NAND2_X1 U11992 ( .A1(n10601), .A2(n10600), .ZN(n10644) );
  OR2_X1 U11993 ( .A1(n11127), .A2(n11103), .ZN(n10601) );
  INV_X1 U11994 ( .A(n10808), .ZN(n10523) );
  BUF_X1 U11995 ( .A(n12460), .Z(n12493) );
  AND2_X1 U11996 ( .A1(n11918), .A2(n9998), .ZN(n9996) );
  NAND2_X1 U11997 ( .A1(n12696), .A2(n11961), .ZN(n12755) );
  OR2_X1 U11998 ( .A1(n11932), .A2(n11931), .ZN(n12756) );
  NOR2_X1 U11999 ( .A1(n9993), .A2(n12754), .ZN(n9990) );
  NOR2_X1 U12000 ( .A1(n9994), .A2(n9996), .ZN(n9993) );
  INV_X1 U12001 ( .A(n9997), .ZN(n9994) );
  NAND2_X1 U12002 ( .A1(n9997), .A2(n9998), .ZN(n9995) );
  INV_X1 U12003 ( .A(n9982), .ZN(n11757) );
  OAI211_X1 U12004 ( .C1(n11722), .C2(n9986), .A(n10167), .B(n11845), .ZN(
        n9982) );
  NAND2_X1 U12005 ( .A1(n11811), .A2(n10168), .ZN(n10167) );
  INV_X1 U12006 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10168) );
  OR2_X1 U12007 ( .A1(n11878), .A2(n11877), .ZN(n12739) );
  NAND2_X1 U12008 ( .A1(n20660), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10600) );
  NOR2_X1 U12009 ( .A1(n11333), .A2(n10496), .ZN(n10495) );
  INV_X1 U12010 ( .A(n11329), .ZN(n10496) );
  OAI211_X1 U12011 ( .C1(n10836), .C2(n10819), .A(n10817), .B(n10818), .ZN(
        n10063) );
  NAND2_X1 U12012 ( .A1(n9859), .A2(n10799), .ZN(n10817) );
  INV_X1 U12013 ( .A(n10816), .ZN(n9950) );
  NOR2_X1 U12014 ( .A1(n10696), .A2(n10695), .ZN(n11328) );
  NOR2_X2 U12015 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10565) );
  AND2_X1 U12016 ( .A1(n14668), .A2(n10750), .ZN(n10893) );
  NAND2_X1 U12017 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20667), .ZN(
        n11103) );
  AND2_X1 U12018 ( .A1(n10812), .A2(n12597), .ZN(n9863) );
  NAND2_X1 U12019 ( .A1(n11156), .A2(n9862), .ZN(n11164) );
  AND2_X1 U12020 ( .A1(n13290), .A2(n13291), .ZN(n13163) );
  NAND2_X1 U12021 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n13329), .ZN(
        n10349) );
  NOR2_X1 U12022 ( .A1(n13317), .A2(n13318), .ZN(n10074) );
  INV_X1 U12023 ( .A(n19066), .ZN(n13271) );
  OAI21_X1 U12024 ( .B1(n13277), .B2(n19084), .A(n13278), .ZN(n10206) );
  NAND2_X1 U12025 ( .A1(n9898), .A2(n9896), .ZN(n12548) );
  INV_X1 U12026 ( .A(n9897), .ZN(n9896) );
  OAI21_X1 U12027 ( .B1(n12538), .B2(n9614), .A(n9693), .ZN(n9897) );
  NAND2_X1 U12028 ( .A1(n9899), .A2(n9903), .ZN(n12545) );
  INV_X1 U12029 ( .A(n12522), .ZN(n9899) );
  NAND2_X1 U12030 ( .A1(n12543), .A2(n12960), .ZN(n12555) );
  OR2_X1 U12031 ( .A1(n12551), .A2(n12550), .ZN(n12554) );
  AND4_X1 U12032 ( .A1(n11611), .A2(n11610), .A3(n11609), .A4(n11608), .ZN(
        n11626) );
  AND4_X1 U12033 ( .A1(n11615), .A2(n11614), .A3(n11613), .A4(n11612), .ZN(
        n11625) );
  AND4_X1 U12034 ( .A1(n11663), .A2(n11662), .A3(n11661), .A4(n11660), .ZN(
        n10555) );
  INV_X1 U12035 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11666) );
  AOI22_X1 U12036 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11689) );
  NOR2_X1 U12037 ( .A1(n10452), .A2(n14761), .ZN(n10451) );
  OR4_X1 U12038 ( .A1(n12335), .A2(n12334), .A3(n12333), .A4(n12332), .ZN(
        n12362) );
  XNOR2_X1 U12039 ( .A(n12696), .B(n11970), .ZN(n12764) );
  NAND2_X1 U12040 ( .A1(n10445), .A2(n9996), .ZN(n9992) );
  OR2_X1 U12041 ( .A1(n11918), .A2(n9998), .ZN(n9997) );
  INV_X1 U12042 ( .A(n11942), .ZN(n9998) );
  AND2_X1 U12043 ( .A1(n11910), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11936) );
  AND2_X1 U12044 ( .A1(n10005), .A2(n13020), .ZN(n10003) );
  INV_X1 U12045 ( .A(n10004), .ZN(n10001) );
  NAND2_X1 U12046 ( .A1(n10121), .A2(n9680), .ZN(n15205) );
  NAND2_X1 U12047 ( .A1(n15237), .A2(n10122), .ZN(n10121) );
  INV_X1 U12048 ( .A(n14817), .ZN(n10435) );
  AND2_X1 U12049 ( .A1(n10437), .A2(n14843), .ZN(n10436) );
  INV_X1 U12050 ( .A(n14829), .ZN(n10437) );
  AOI21_X1 U12051 ( .B1(n15237), .B2(n12779), .A(n9876), .ZN(n15207) );
  NAND2_X1 U12052 ( .A1(n9655), .A2(n15353), .ZN(n9876) );
  INV_X1 U12053 ( .A(n10078), .ZN(n10077) );
  OAI21_X1 U12054 ( .B1(n10279), .B2(n10123), .A(n10119), .ZN(n10078) );
  INV_X1 U12055 ( .A(n14920), .ZN(n10431) );
  AND2_X1 U12056 ( .A1(n15309), .A2(n15312), .ZN(n15283) );
  INV_X1 U12057 ( .A(n14962), .ZN(n10433) );
  OR2_X1 U12058 ( .A1(n15353), .A2(n21418), .ZN(n15281) );
  INV_X1 U12059 ( .A(n14168), .ZN(n10429) );
  INV_X1 U12060 ( .A(n12984), .ZN(n10170) );
  OAI211_X1 U12061 ( .C1(n12542), .C2(n11815), .A(n11814), .B(n11813), .ZN(
        n11843) );
  OAI22_X1 U12062 ( .A1(n11812), .A2(n11862), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n9986), .ZN(n11844) );
  OR2_X1 U12063 ( .A1(n11778), .A2(n11777), .ZN(n12714) );
  AND2_X1 U12064 ( .A1(n15613), .A2(n13808), .ZN(n10315) );
  NAND2_X1 U12065 ( .A1(n10313), .A2(n11721), .ZN(n11728) );
  AND2_X1 U12066 ( .A1(n21203), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11724) );
  OR2_X2 U12067 ( .A1(n11658), .A2(n11657), .ZN(n12719) );
  INV_X1 U12068 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n17091) );
  AOI21_X1 U12069 ( .B1(n10670), .B2(n10669), .A(n10668), .ZN(n11117) );
  INV_X1 U12070 ( .A(n10667), .ZN(n10669) );
  AND2_X1 U12071 ( .A1(n10478), .A2(n11075), .ZN(n10475) );
  NOR2_X1 U12072 ( .A1(n11042), .A2(n10479), .ZN(n10478) );
  NAND2_X1 U12073 ( .A1(n10722), .A2(n11044), .ZN(n10479) );
  OR2_X1 U12074 ( .A1(n10385), .A2(n12604), .ZN(n10379) );
  NAND2_X1 U12075 ( .A1(n12642), .A2(n10378), .ZN(n10383) );
  INV_X1 U12076 ( .A(n12605), .ZN(n10378) );
  NAND2_X1 U12077 ( .A1(n10472), .A2(n10721), .ZN(n10471) );
  NOR2_X1 U12078 ( .A1(n10405), .A2(n10404), .ZN(n10403) );
  CLKBUF_X1 U12079 ( .A(n10984), .Z(n10985) );
  NAND2_X1 U12080 ( .A1(n10815), .A2(n10816), .ZN(n10033) );
  CLKBUF_X1 U12081 ( .A(n14512), .Z(n14682) );
  CLKBUF_X1 U12082 ( .A(n14556), .Z(n14683) );
  CLKBUF_X1 U12083 ( .A(n14514), .Z(n14681) );
  CLKBUF_X1 U12084 ( .A(n14515), .Z(n14679) );
  INV_X1 U12085 ( .A(n14625), .ZN(n14605) );
  INV_X1 U12086 ( .A(n16108), .ZN(n10463) );
  AND2_X1 U12087 ( .A1(n15856), .A2(n15842), .ZN(n10493) );
  NAND2_X1 U12088 ( .A1(n12641), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12643) );
  NAND2_X1 U12089 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10410) );
  OR2_X1 U12090 ( .A1(n10410), .A2(n10409), .ZN(n10408) );
  INV_X1 U12091 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10409) );
  NAND2_X1 U12092 ( .A1(n10486), .A2(n14052), .ZN(n10485) );
  INV_X1 U12093 ( .A(n16131), .ZN(n10486) );
  NAND2_X1 U12094 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10405) );
  NAND2_X1 U12095 ( .A1(n10061), .A2(n10842), .ZN(n9918) );
  NAND2_X1 U12096 ( .A1(n10824), .A2(n10823), .ZN(n10849) );
  NAND2_X1 U12097 ( .A1(n10821), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10824) );
  INV_X1 U12098 ( .A(n14328), .ZN(n10490) );
  NAND2_X1 U12099 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10528) );
  NOR2_X1 U12100 ( .A1(n15804), .A2(n11542), .ZN(n16317) );
  INV_X1 U12101 ( .A(n16318), .ZN(n9936) );
  INV_X1 U12102 ( .A(n15871), .ZN(n10519) );
  NAND2_X1 U12103 ( .A1(n9955), .A2(n9952), .ZN(n9954) );
  NAND2_X1 U12104 ( .A1(n16495), .A2(n11545), .ZN(n9953) );
  AND2_X1 U12105 ( .A1(n11096), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9952) );
  NAND2_X1 U12106 ( .A1(n11072), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16345) );
  NAND2_X1 U12107 ( .A1(n11069), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10010) );
  INV_X1 U12108 ( .A(n10010), .ZN(n9889) );
  NAND2_X1 U12109 ( .A1(n10220), .A2(n14346), .ZN(n10219) );
  NAND2_X1 U12110 ( .A1(n9600), .A2(n16425), .ZN(n10416) );
  INV_X1 U12111 ( .A(n10220), .ZN(n9968) );
  NAND2_X1 U12112 ( .A1(n10484), .A2(n14152), .ZN(n10483) );
  INV_X1 U12113 ( .A(n10485), .ZN(n10484) );
  NAND2_X1 U12114 ( .A1(n16268), .A2(n10515), .ZN(n10514) );
  INV_X1 U12115 ( .A(n14162), .ZN(n10515) );
  OR2_X1 U12116 ( .A1(n15922), .A2(n11542), .ZN(n11060) );
  NAND2_X1 U12117 ( .A1(n14348), .A2(n14349), .ZN(n10221) );
  NOR2_X1 U12118 ( .A1(n16716), .A2(n16713), .ZN(n10375) );
  OR2_X1 U12119 ( .A1(n15948), .A2(n11542), .ZN(n14349) );
  AND3_X1 U12120 ( .A1(n11377), .A2(n11376), .A3(n11375), .ZN(n13783) );
  INV_X1 U12121 ( .A(n14207), .ZN(n10487) );
  NAND2_X1 U12122 ( .A1(n9765), .A2(n10372), .ZN(n10130) );
  NAND2_X1 U12123 ( .A1(n9955), .A2(n11096), .ZN(n16498) );
  NAND2_X1 U12124 ( .A1(n11543), .A2(n11542), .ZN(n16495) );
  INV_X1 U12125 ( .A(n11522), .ZN(n11537) );
  AND2_X1 U12126 ( .A1(n9777), .A2(n16534), .ZN(n9793) );
  AND2_X1 U12127 ( .A1(n16517), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9777) );
  NAND2_X1 U12129 ( .A1(n11536), .A2(n16805), .ZN(n11540) );
  AND4_X1 U12130 ( .A1(n10925), .A2(n10924), .A3(n10923), .A4(n10922), .ZN(
        n10934) );
  XNOR2_X1 U12131 ( .A(n11534), .B(n11535), .ZN(n9880) );
  NAND2_X1 U12132 ( .A1(n9827), .A2(n11533), .ZN(n9881) );
  INV_X1 U12133 ( .A(n16538), .ZN(n10182) );
  NAND2_X1 U12134 ( .A1(n9806), .A2(n9805), .ZN(n11479) );
  AND2_X1 U12135 ( .A1(n10785), .A2(n10788), .ZN(n10366) );
  AND2_X1 U12136 ( .A1(n10556), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10566) );
  NOR2_X1 U12137 ( .A1(n14605), .A2(n13603), .ZN(n13769) );
  NAND2_X1 U12138 ( .A1(n13871), .A2(n13872), .ZN(n13927) );
  NAND2_X1 U12139 ( .A1(n10770), .A2(n10769), .ZN(n10789) );
  NAND2_X1 U12140 ( .A1(n11172), .A2(n11126), .ZN(n16925) );
  NAND2_X1 U12141 ( .A1(n11125), .A2(n11124), .ZN(n11126) );
  OAI211_X1 U12142 ( .C1(n13197), .C2(n13192), .A(n13191), .B(n9646), .ZN(
        n13193) );
  NOR2_X1 U12143 ( .A1(n13042), .A2(n19508), .ZN(n13232) );
  NOR2_X1 U12144 ( .A1(n13033), .A2(n13043), .ZN(n13184) );
  OR2_X1 U12145 ( .A1(n10349), .A2(n17459), .ZN(n10348) );
  NAND2_X1 U12146 ( .A1(n13155), .A2(n10142), .ZN(n10229) );
  AND2_X1 U12147 ( .A1(n10228), .A2(n21367), .ZN(n10227) );
  OR2_X1 U12148 ( .A1(n18634), .A2(n17269), .ZN(n10228) );
  AND2_X1 U12149 ( .A1(n18213), .A2(n17146), .ZN(n13274) );
  NAND2_X1 U12150 ( .A1(n10223), .A2(n13142), .ZN(n13143) );
  AND2_X1 U12151 ( .A1(n10142), .A2(n10141), .ZN(n13141) );
  NAND2_X1 U12152 ( .A1(n17288), .A2(n18222), .ZN(n10141) );
  XNOR2_X1 U12153 ( .A(n13298), .B(n18247), .ZN(n13074) );
  NAND2_X1 U12154 ( .A1(n13263), .A2(n9937), .ZN(n13264) );
  AOI22_X1 U12155 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n21428), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n13161), .ZN(n13290) );
  OAI21_X1 U12156 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n21439), .A(
        n13172), .ZN(n13292) );
  INV_X1 U12157 ( .A(n13044), .ZN(n10255) );
  OAI21_X1 U12158 ( .B1(n13332), .B2(n19537), .A(n19658), .ZN(n19054) );
  INV_X1 U12159 ( .A(n19515), .ZN(n9945) );
  NOR2_X2 U12160 ( .A1(n13777), .A2(n13563), .ZN(n17109) );
  NOR2_X1 U12161 ( .A1(n17097), .A2(n17103), .ZN(n17108) );
  NAND2_X2 U12162 ( .A1(n13818), .A2(n13563), .ZN(n15020) );
  NOR2_X1 U12163 ( .A1(n20784), .A2(n17222), .ZN(n12912) );
  NAND2_X1 U12164 ( .A1(n10451), .A2(n12802), .ZN(n10450) );
  NAND2_X1 U12165 ( .A1(n12574), .A2(n12573), .ZN(n13638) );
  OR2_X1 U12166 ( .A1(n17107), .A2(n12565), .ZN(n12574) );
  OR2_X1 U12167 ( .A1(n15154), .A2(n13760), .ZN(n13763) );
  AOI21_X1 U12168 ( .B1(n20856), .B2(n13776), .A(n17142), .ZN(n20801) );
  OR2_X1 U12169 ( .A1(n13775), .A2(n15669), .ZN(n13776) );
  INV_X1 U12170 ( .A(n20842), .ZN(n13729) );
  INV_X1 U12171 ( .A(n15085), .ZN(n13803) );
  AND2_X1 U12172 ( .A1(n12442), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12443) );
  AOI21_X1 U12173 ( .B1(n15187), .B2(n12273), .A(n12440), .ZN(n14772) );
  OAI21_X1 U12174 ( .B1(n15192), .B2(n12503), .A(n12418), .ZN(n14785) );
  OR2_X1 U12175 ( .A1(n12342), .A2(n15221), .ZN(n12344) );
  OAI21_X1 U12176 ( .B1(n15214), .B2(n12503), .A(n12367), .ZN(n14805) );
  AND2_X1 U12177 ( .A1(n12275), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12276) );
  AND2_X1 U12178 ( .A1(n12235), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12236) );
  INV_X1 U12179 ( .A(n12234), .ZN(n12235) );
  OAI21_X1 U12180 ( .B1(n15249), .B2(n12503), .A(n12257), .ZN(n14851) );
  NOR2_X1 U12181 ( .A1(n12178), .A2(n15271), .ZN(n12116) );
  AND2_X1 U12182 ( .A1(n12140), .A2(n12139), .ZN(n14876) );
  AOI21_X1 U12183 ( .B1(n15291), .B2(n11907), .A(n12213), .ZN(n14902) );
  NOR2_X1 U12184 ( .A1(n14915), .A2(n14902), .ZN(n14901) );
  NOR2_X1 U12185 ( .A1(n14942), .A2(n14874), .ZN(n14928) );
  AND2_X1 U12186 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12093) );
  INV_X1 U12187 ( .A(n10088), .ZN(n10087) );
  OAI21_X1 U12188 ( .B1(n11993), .B2(n10089), .A(n10439), .ZN(n10088) );
  INV_X1 U12189 ( .A(n12054), .ZN(n10089) );
  NAND2_X1 U12190 ( .A1(n12037), .A2(n12036), .ZN(n12073) );
  NOR2_X1 U12191 ( .A1(n14990), .A2(n14989), .ZN(n14988) );
  NOR2_X1 U12192 ( .A1(n12014), .A2(n12013), .ZN(n12037) );
  INV_X1 U12193 ( .A(n14264), .ZN(n10444) );
  OR2_X1 U12194 ( .A1(n12008), .A2(n15010), .ZN(n12014) );
  AND3_X1 U12195 ( .A1(n12012), .A2(n12011), .A3(n12010), .ZN(n14271) );
  AND3_X1 U12196 ( .A1(n11992), .A2(n11991), .A3(n11990), .ZN(n14263) );
  INV_X1 U12197 ( .A(n11971), .ZN(n11972) );
  NAND2_X1 U12198 ( .A1(n11972), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12008) );
  NAND2_X1 U12199 ( .A1(n11963), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11971) );
  AND2_X1 U12200 ( .A1(n11936), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11963) );
  AND2_X1 U12201 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11909), .ZN(
        n11910) );
  NAND2_X1 U12202 ( .A1(n11888), .A2(n11887), .ZN(n13975) );
  NAND2_X1 U12203 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11883) );
  OAI21_X1 U12204 ( .B1(n14006), .B2(n12172), .A(n11834), .ZN(n11835) );
  INV_X1 U12205 ( .A(n12783), .ZN(n10180) );
  OR2_X1 U12206 ( .A1(n14762), .A2(n12944), .ZN(n12947) );
  NAND2_X1 U12207 ( .A1(n14762), .A2(n12945), .ZN(n12946) );
  OR2_X1 U12208 ( .A1(n14763), .A2(n14776), .ZN(n10419) );
  NOR2_X1 U12209 ( .A1(n15374), .A2(n15391), .ZN(n10320) );
  NAND2_X1 U12210 ( .A1(n14853), .A2(n10436), .ZN(n14831) );
  INV_X1 U12211 ( .A(n12781), .ZN(n15228) );
  AND2_X1 U12212 ( .A1(n12876), .A2(n12875), .ZN(n14890) );
  NAND2_X1 U12213 ( .A1(n14919), .A2(n9721), .ZN(n14906) );
  AND2_X1 U12214 ( .A1(n12868), .A2(n12867), .ZN(n14932) );
  OR2_X1 U12215 ( .A1(n15353), .A2(n15534), .ZN(n15312) );
  AND2_X1 U12216 ( .A1(n12866), .A2(n12865), .ZN(n14947) );
  NAND2_X1 U12217 ( .A1(n14994), .A2(n9649), .ZN(n14960) );
  AND2_X1 U12218 ( .A1(n12857), .A2(n12856), .ZN(n14993) );
  AND2_X1 U12219 ( .A1(n10424), .A2(n10422), .ZN(n10421) );
  INV_X1 U12220 ( .A(n14273), .ZN(n10422) );
  NAND2_X1 U12221 ( .A1(n10423), .A2(n10424), .ZN(n14274) );
  NAND2_X1 U12222 ( .A1(n15366), .A2(n12708), .ZN(n15383) );
  NOR2_X1 U12223 ( .A1(n14259), .A2(n14260), .ZN(n14267) );
  AND2_X1 U12224 ( .A1(n12840), .A2(n12839), .ZN(n14176) );
  INV_X1 U12225 ( .A(n20867), .ZN(n10071) );
  INV_X1 U12226 ( .A(n13787), .ZN(n12824) );
  INV_X1 U12227 ( .A(n13786), .ZN(n12825) );
  NOR2_X1 U12228 ( .A1(n14046), .A2(n14045), .ZN(n14169) );
  NAND2_X1 U12229 ( .A1(n20867), .A2(n20866), .ZN(n20865) );
  NAND2_X1 U12230 ( .A1(n13748), .A2(n21470), .ZN(n13746) );
  NAND2_X1 U12231 ( .A1(n9871), .A2(n11828), .ZN(n13025) );
  AND2_X1 U12232 ( .A1(n10315), .A2(n17109), .ZN(n9871) );
  OAI211_X1 U12233 ( .C1(n11667), .C2(n11594), .A(n11593), .B(n11592), .ZN(
        n11595) );
  INV_X1 U12234 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13664) );
  NOR2_X1 U12235 ( .A1(n17097), .A2(n13829), .ZN(n17084) );
  AND4_X1 U12236 ( .A1(n11632), .A2(n11631), .A3(n11630), .A4(n11629), .ZN(
        n11644) );
  NOR2_X1 U12237 ( .A1(n11642), .A2(n11641), .ZN(n11643) );
  INV_X1 U12238 ( .A(n15679), .ZN(n21030) );
  INV_X1 U12239 ( .A(n14076), .ZN(n21091) );
  NAND3_X1 U12240 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n11759), .A3(n13807), 
        .ZN(n13846) );
  OR2_X1 U12241 ( .A1(n17107), .A2(n21064), .ZN(n13798) );
  NAND2_X1 U12242 ( .A1(n10919), .A2(n10793), .ZN(n10648) );
  NAND2_X1 U12243 ( .A1(n10603), .A2(n11112), .ZN(n11130) );
  NAND2_X1 U12244 ( .A1(n9698), .A2(n19866), .ZN(n10244) );
  OR2_X1 U12246 ( .A1(n15857), .A2(n10245), .ZN(n10246) );
  NAND2_X1 U12247 ( .A1(n11099), .A2(n11083), .ZN(n11085) );
  AND2_X1 U12248 ( .A1(n15857), .A2(n16356), .ZN(n15844) );
  NAND2_X1 U12249 ( .A1(n10383), .A2(n10381), .ZN(n15874) );
  NOR2_X1 U12250 ( .A1(n10382), .A2(n10384), .ZN(n10381) );
  INV_X1 U12251 ( .A(n10379), .ZN(n10382) );
  NAND2_X1 U12252 ( .A1(n12640), .A2(n10235), .ZN(n15897) );
  NOR2_X1 U12253 ( .A1(n19747), .A2(n10236), .ZN(n10235) );
  INV_X1 U12254 ( .A(n19760), .ZN(n10236) );
  NAND2_X1 U12255 ( .A1(n19866), .A2(n12642), .ZN(n15886) );
  NAND2_X1 U12256 ( .A1(n10473), .A2(n10474), .ZN(n11014) );
  NOR2_X1 U12257 ( .A1(n10029), .A2(n10028), .ZN(n10027) );
  INV_X1 U12258 ( .A(n11015), .ZN(n10028) );
  INV_X1 U12259 ( .A(n10472), .ZN(n10029) );
  NAND2_X1 U12260 ( .A1(n10720), .A2(n9733), .ZN(n10019) );
  INV_X1 U12261 ( .A(n11027), .ZN(n10719) );
  NAND2_X1 U12262 ( .A1(n11029), .A2(n11032), .ZN(n11026) );
  NOR2_X1 U12263 ( .A1(n12618), .A2(n10402), .ZN(n12614) );
  NAND2_X1 U12264 ( .A1(n10403), .A2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10402) );
  CLKBUF_X1 U12265 ( .A(n10986), .Z(n10995) );
  NOR2_X1 U12266 ( .A1(n19865), .A2(n19868), .ZN(n19845) );
  NAND2_X1 U12267 ( .A1(n15968), .A2(n16530), .ZN(n19865) );
  NOR2_X1 U12268 ( .A1(n15983), .A2(n19942), .ZN(n15968) );
  NAND2_X1 U12269 ( .A1(n10238), .A2(n10237), .ZN(n15999) );
  INV_X1 U12270 ( .A(n16027), .ZN(n10238) );
  NAND2_X1 U12271 ( .A1(n16028), .A2(n16823), .ZN(n16027) );
  INV_X1 U12272 ( .A(n19806), .ZN(n16043) );
  INV_X1 U12273 ( .A(n14063), .ZN(n10455) );
  INV_X1 U12274 ( .A(n14608), .ZN(n14629) );
  NAND2_X1 U12275 ( .A1(n9623), .A2(n10517), .ZN(n10516) );
  INV_X1 U12276 ( .A(n15835), .ZN(n10517) );
  XNOR2_X1 U12277 ( .A(n14604), .B(n14603), .ZN(n16075) );
  NAND2_X1 U12278 ( .A1(n10519), .A2(n10520), .ZN(n15838) );
  AND2_X1 U12279 ( .A1(n11459), .A2(n11458), .ZN(n15873) );
  NOR2_X1 U12280 ( .A1(n15871), .A2(n15873), .ZN(n15861) );
  AND2_X1 U12281 ( .A1(n16120), .A2(n10462), .ZN(n16093) );
  AND2_X1 U12282 ( .A1(n11449), .A2(n11448), .ZN(n16239) );
  NAND2_X1 U12283 ( .A1(n16120), .A2(n14463), .ZN(n16113) );
  NAND2_X1 U12284 ( .A1(n10510), .A2(n10509), .ZN(n10508) );
  INV_X1 U12285 ( .A(n14727), .ZN(n10509) );
  INV_X1 U12286 ( .A(n10512), .ZN(n10510) );
  AND3_X1 U12287 ( .A1(n11415), .A2(n11414), .A3(n11413), .ZN(n13935) );
  CLKBUF_X1 U12288 ( .A(n13855), .Z(n13856) );
  AND3_X1 U12289 ( .A1(n11390), .A2(n11389), .A3(n11388), .ZN(n13878) );
  INV_X1 U12290 ( .A(n13679), .ZN(n11350) );
  NOR2_X1 U12291 ( .A1(n19887), .A2(n13576), .ZN(n14694) );
  NAND2_X1 U12292 ( .A1(n10784), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13493) );
  INV_X1 U12293 ( .A(n11173), .ZN(n13489) );
  NOR2_X1 U12294 ( .A1(n12598), .A2(n9861), .ZN(n13488) );
  NAND2_X1 U12295 ( .A1(n10391), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10386) );
  OR2_X1 U12296 ( .A1(n12656), .A2(n10389), .ZN(n10388) );
  NAND2_X1 U12297 ( .A1(n12656), .A2(n9751), .ZN(n10387) );
  NOR2_X1 U12298 ( .A1(n12653), .A2(n16319), .ZN(n12656) );
  AND2_X1 U12299 ( .A1(n9622), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10397) );
  NAND2_X1 U12300 ( .A1(n12641), .A2(n9622), .ZN(n12646) );
  AND2_X1 U12301 ( .A1(n12607), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12641) );
  NOR2_X1 U12302 ( .A1(n12636), .A2(n10406), .ZN(n12607) );
  NAND2_X1 U12303 ( .A1(n10407), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10406) );
  INV_X1 U12304 ( .A(n10408), .ZN(n10407) );
  NOR2_X1 U12305 ( .A1(n12636), .A2(n10410), .ZN(n12639) );
  AND2_X1 U12306 ( .A1(n14722), .A2(n10111), .ZN(n10110) );
  INV_X1 U12307 ( .A(n14362), .ZN(n10111) );
  NAND2_X1 U12308 ( .A1(n12601), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12632) );
  INV_X1 U12309 ( .A(n12630), .ZN(n12601) );
  AND2_X1 U12310 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10392) );
  NAND2_X1 U12311 ( .A1(n10395), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12626) );
  NOR2_X1 U12312 ( .A1(n10396), .A2(n12624), .ZN(n10395) );
  NOR2_X1 U12313 ( .A1(n10396), .A2(n16013), .ZN(n10394) );
  NOR2_X1 U12314 ( .A1(n12624), .A2(n19954), .ZN(n10393) );
  NAND2_X1 U12315 ( .A1(n10849), .A2(n10848), .ZN(n10860) );
  INV_X1 U12316 ( .A(n11102), .ZN(n10355) );
  OR2_X1 U12317 ( .A1(n10528), .A2(n16557), .ZN(n10527) );
  NOR2_X1 U12318 ( .A1(n14302), .A2(n10359), .ZN(n10358) );
  INV_X1 U12319 ( .A(n16294), .ZN(n10359) );
  INV_X1 U12320 ( .A(n10023), .ZN(n10022) );
  OAI21_X1 U12321 ( .B1(n10024), .B2(n10026), .A(n16294), .ZN(n10023) );
  NAND2_X1 U12322 ( .A1(n16327), .A2(n10011), .ZN(n16316) );
  NAND2_X1 U12323 ( .A1(n16625), .A2(n10060), .ZN(n16570) );
  AND2_X1 U12324 ( .A1(n9609), .A2(n9701), .ZN(n10060) );
  NAND2_X1 U12325 ( .A1(n16315), .A2(n9936), .ZN(n9935) );
  NAND2_X1 U12326 ( .A1(n10152), .A2(n10292), .ZN(n10150) );
  INV_X1 U12327 ( .A(n10290), .ZN(n10152) );
  NAND2_X1 U12328 ( .A1(n10149), .A2(n10292), .ZN(n10151) );
  NAND2_X1 U12329 ( .A1(n16348), .A2(n16616), .ZN(n10364) );
  NAND2_X1 U12330 ( .A1(n16578), .A2(n16579), .ZN(n9848) );
  NAND2_X1 U12331 ( .A1(n16625), .A2(n9609), .ZN(n16588) );
  NAND2_X1 U12332 ( .A1(n16625), .A2(n11508), .ZN(n16601) );
  OR2_X1 U12333 ( .A1(n9636), .A2(n9889), .ZN(n9888) );
  NAND2_X1 U12334 ( .A1(n9636), .A2(n10010), .ZN(n9886) );
  NOR2_X1 U12335 ( .A1(n16361), .A2(n9889), .ZN(n9887) );
  CLKBUF_X1 U12336 ( .A(n14366), .Z(n14401) );
  NAND2_X1 U12337 ( .A1(n14360), .A2(n10109), .ZN(n14398) );
  AND2_X1 U12338 ( .A1(n10110), .A2(n16638), .ZN(n10109) );
  INV_X1 U12339 ( .A(n16110), .ZN(n11233) );
  CLKBUF_X1 U12340 ( .A(n14718), .Z(n14719) );
  AOI21_X1 U12341 ( .B1(n10296), .B2(n10300), .A(n10295), .ZN(n10294) );
  INV_X1 U12342 ( .A(n14710), .ZN(n10295) );
  OR2_X1 U12343 ( .A1(n15914), .A2(n11054), .ZN(n14706) );
  NAND2_X1 U12344 ( .A1(n14360), .A2(n9634), .ZN(n9966) );
  OR2_X1 U12345 ( .A1(n14349), .A2(n16713), .ZN(n16435) );
  NAND2_X1 U12346 ( .A1(n14360), .A2(n10068), .ZN(n10067) );
  NOR2_X1 U12347 ( .A1(n16716), .A2(n16739), .ZN(n10068) );
  INV_X1 U12348 ( .A(n16142), .ZN(n11209) );
  NAND2_X1 U12349 ( .A1(n11198), .A2(n11197), .ZN(n14208) );
  INV_X1 U12350 ( .A(n10997), .ZN(n16456) );
  OAI21_X1 U12351 ( .B1(n16534), .B2(n11522), .A(n11541), .ZN(n10108) );
  NAND2_X1 U12352 ( .A1(n9765), .A2(n9686), .ZN(n9794) );
  CLKBUF_X1 U12353 ( .A(n11479), .Z(n16934) );
  NAND2_X1 U12354 ( .A1(n9880), .A2(n9881), .ZN(n16804) );
  AOI21_X1 U12355 ( .B1(n16540), .B2(n9734), .A(n9922), .ZN(n9921) );
  NOR2_X1 U12356 ( .A1(n16003), .A2(n10838), .ZN(n9922) );
  NAND2_X1 U12357 ( .A1(n11502), .A2(n17233), .ZN(n16810) );
  NAND2_X1 U12358 ( .A1(n13650), .A2(n11310), .ZN(n15997) );
  NAND2_X1 U12359 ( .A1(n16024), .A2(n16023), .ZN(n16025) );
  NAND2_X1 U12360 ( .A1(n9786), .A2(n13768), .ZN(n9785) );
  AND2_X1 U12361 ( .A1(n11306), .A2(n11305), .ZN(n13647) );
  AND2_X1 U12362 ( .A1(n11498), .A2(n11497), .ZN(n16830) );
  XNOR2_X1 U12363 ( .A(n16826), .B(n13769), .ZN(n13771) );
  INV_X1 U12364 ( .A(n20247), .ZN(n20249) );
  NOR2_X1 U12365 ( .A1(n20637), .A2(n16907), .ZN(n20007) );
  INV_X1 U12366 ( .A(n20007), .ZN(n20174) );
  NOR2_X1 U12367 ( .A1(n20629), .A2(n20174), .ZN(n20213) );
  OR2_X1 U12368 ( .A1(n16903), .A2(n16902), .ZN(n16909) );
  NAND2_X1 U12369 ( .A1(n10780), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9783) );
  NAND2_X1 U12370 ( .A1(n20637), .A2(n16907), .ZN(n20405) );
  NAND2_X1 U12371 ( .A1(n10740), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9780) );
  NAND2_X1 U12372 ( .A1(n10745), .A2(n10750), .ZN(n9781) );
  AND2_X1 U12373 ( .A1(n20476), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19998) );
  NOR2_X2 U12374 ( .A1(n16873), .A2(n19950), .ZN(n20001) );
  NOR2_X2 U12375 ( .A1(n16872), .A2(n19950), .ZN(n20002) );
  AND2_X1 U12376 ( .A1(n16925), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17251) );
  OR3_X1 U12377 ( .A1(n10260), .A2(n13237), .A3(n13238), .ZN(n13266) );
  NAND2_X1 U12378 ( .A1(n10325), .A2(n10323), .ZN(n17456) );
  NAND2_X1 U12379 ( .A1(n17653), .A2(n10324), .ZN(n10323) );
  INV_X1 U12380 ( .A(n17458), .ZN(n10324) );
  NOR2_X1 U12381 ( .A1(n17489), .A2(n18399), .ZN(n17488) );
  NAND2_X1 U12382 ( .A1(n17612), .A2(n17603), .ZN(n17601) );
  NOR2_X1 U12383 ( .A1(n17634), .A2(P3_EBX_REG_14__SCAN_IN), .ZN(n17612) );
  NOR2_X1 U12384 ( .A1(n17764), .A2(P3_EBX_REG_4__SCAN_IN), .ZN(n17745) );
  NAND2_X1 U12385 ( .A1(n19522), .A2(n17417), .ZN(n19698) );
  NAND2_X1 U12386 ( .A1(n17954), .A2(n10263), .ZN(n17887) );
  NOR2_X1 U12387 ( .A1(n21333), .A2(n17953), .ZN(n10266) );
  NOR2_X1 U12388 ( .A1(n17667), .A2(n17686), .ZN(n10269) );
  NOR2_X1 U12389 ( .A1(n19059), .A2(n19056), .ZN(n16967) );
  NOR2_X1 U12390 ( .A1(n18324), .A2(n10202), .ZN(n10201) );
  NOR2_X1 U12391 ( .A1(n10195), .A2(n10193), .ZN(n10192) );
  NAND2_X1 U12392 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .ZN(n10195) );
  NAND2_X1 U12393 ( .A1(n9757), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n10193) );
  NAND2_X1 U12394 ( .A1(n10549), .A2(n10542), .ZN(n18109) );
  OR2_X1 U12395 ( .A1(n13088), .A2(n13087), .ZN(n13101) );
  AOI21_X1 U12396 ( .B1(n17416), .B2(n17064), .A(n17067), .ZN(n17147) );
  NOR2_X1 U12397 ( .A1(n19691), .A2(n17743), .ZN(n17146) );
  INV_X1 U12398 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21312) );
  NOR2_X1 U12399 ( .A1(n18304), .A2(n18255), .ZN(n18257) );
  NOR2_X1 U12400 ( .A1(n18375), .A2(n10348), .ZN(n17270) );
  NOR2_X1 U12401 ( .A1(n18375), .A2(n18714), .ZN(n17439) );
  NOR2_X1 U12402 ( .A1(n18412), .A2(n18413), .ZN(n18394) );
  NAND2_X1 U12403 ( .A1(n18433), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18412) );
  INV_X1 U12404 ( .A(n18446), .ZN(n18444) );
  INV_X1 U12405 ( .A(n18486), .ZN(n10342) );
  NAND2_X1 U12406 ( .A1(n10343), .A2(n10344), .ZN(n18485) );
  NOR2_X1 U12407 ( .A1(n18522), .A2(n18524), .ZN(n18508) );
  NAND3_X1 U12408 ( .A1(n17434), .A2(n18562), .A3(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18522) );
  OAI21_X1 U12409 ( .B1(n18714), .B2(n18441), .A(n19335), .ZN(n18561) );
  AND3_X1 U12410 ( .A1(n10340), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        n10341), .ZN(n18627) );
  NOR2_X1 U12411 ( .A1(n19655), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10038) );
  OR2_X1 U12412 ( .A1(n18731), .A2(n17136), .ZN(n10158) );
  NAND2_X1 U12413 ( .A1(n13154), .A2(n13155), .ZN(n17073) );
  INV_X1 U12414 ( .A(n18382), .ZN(n13153) );
  NAND2_X1 U12415 ( .A1(n18406), .A2(n13324), .ZN(n18731) );
  NOR2_X1 U12416 ( .A1(n18859), .A2(n18748), .ZN(n18406) );
  NAND2_X1 U12417 ( .A1(n9823), .A2(n10225), .ZN(n9822) );
  INV_X1 U12418 ( .A(n18465), .ZN(n9823) );
  INV_X1 U12419 ( .A(n18518), .ZN(n18453) );
  NAND2_X1 U12420 ( .A1(n9657), .A2(n18856), .ZN(n10041) );
  NAND2_X1 U12421 ( .A1(n18633), .A2(n18596), .ZN(n18539) );
  INV_X1 U12422 ( .A(n18532), .ZN(n18860) );
  NAND2_X1 U12423 ( .A1(n18909), .A2(n13336), .ZN(n18554) );
  NOR2_X1 U12424 ( .A1(n18847), .A2(n13337), .ZN(n18550) );
  INV_X1 U12425 ( .A(n18596), .ZN(n18538) );
  INV_X1 U12426 ( .A(n13337), .ZN(n18911) );
  NAND2_X1 U12427 ( .A1(n18622), .A2(n13323), .ZN(n18909) );
  NAND3_X1 U12428 ( .A1(n10081), .A2(n13320), .A3(n9715), .ZN(n18623) );
  NAND2_X1 U12429 ( .A1(n18623), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18622) );
  NAND2_X1 U12430 ( .A1(n18663), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10306) );
  NAND2_X1 U12431 ( .A1(n18690), .A2(n13312), .ZN(n18676) );
  XNOR2_X1 U12432 ( .A(n13307), .B(n19011), .ZN(n18692) );
  NAND2_X1 U12433 ( .A1(n18691), .A2(n18692), .ZN(n18690) );
  XNOR2_X1 U12434 ( .A(n13074), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18702) );
  NAND2_X1 U12435 ( .A1(n10302), .A2(n13073), .ZN(n9826) );
  NOR2_X1 U12436 ( .A1(n18851), .A2(n13358), .ZN(n19525) );
  NOR3_X1 U12437 ( .A1(n10199), .A2(n10198), .A3(n10197), .ZN(n10196) );
  NOR2_X1 U12438 ( .A1(n13358), .A2(n19524), .ZN(n13356) );
  INV_X1 U12439 ( .A(n17063), .ZN(n19523) );
  INV_X1 U12440 ( .A(n19502), .ZN(n19509) );
  NOR2_X1 U12441 ( .A1(n13288), .A2(n13286), .ZN(n19491) );
  INV_X1 U12442 ( .A(n19334), .ZN(n19394) );
  NOR2_X2 U12443 ( .A1(n13250), .A2(n13249), .ZN(n19070) );
  NOR2_X2 U12444 ( .A1(n13229), .A2(n13228), .ZN(n19074) );
  NAND2_X1 U12445 ( .A1(n19696), .A2(n19054), .ZN(n19334) );
  AND2_X1 U12446 ( .A1(n15027), .A2(n12943), .ZN(n14755) );
  NOR2_X1 U12447 ( .A1(n9581), .A2(n11759), .ZN(n13523) );
  NAND2_X1 U12448 ( .A1(n15001), .A2(n10053), .ZN(n14860) );
  AND2_X1 U12449 ( .A1(n9756), .A2(n10054), .ZN(n10053) );
  INV_X1 U12450 ( .A(n12931), .ZN(n10054) );
  NAND2_X1 U12451 ( .A1(n15001), .A2(n9756), .ZN(n14896) );
  AND2_X1 U12452 ( .A1(n15001), .A2(n12925), .ZN(n14925) );
  AND2_X1 U12453 ( .A1(n17160), .A2(n12928), .ZN(n15001) );
  INV_X1 U12454 ( .A(n20729), .ZN(n20755) );
  NAND2_X1 U12455 ( .A1(n20764), .A2(n9759), .ZN(n20735) );
  OR2_X1 U12456 ( .A1(n20784), .A2(n20706), .ZN(n20759) );
  OR2_X1 U12457 ( .A1(n20784), .A2(n21064), .ZN(n20762) );
  NOR2_X1 U12458 ( .A1(n20773), .A2(n21226), .ZN(n20764) );
  OR2_X1 U12459 ( .A1(n15026), .A2(n12918), .ZN(n20781) );
  INV_X1 U12460 ( .A(n20762), .ZN(n20785) );
  OR2_X1 U12461 ( .A1(n20783), .A2(n20784), .ZN(n20729) );
  INV_X1 U12462 ( .A(n20800), .ZN(n15065) );
  AND2_X1 U12463 ( .A1(n20800), .A2(n13834), .ZN(n20795) );
  AND2_X1 U12464 ( .A1(n13745), .A2(n9905), .ZN(n20800) );
  INV_X1 U12465 ( .A(n20796), .ZN(n15067) );
  INV_X1 U12466 ( .A(n20795), .ZN(n15068) );
  NAND2_X1 U12467 ( .A1(n15150), .A2(n13762), .ZN(n15144) );
  INV_X1 U12468 ( .A(n15138), .ZN(n15146) );
  NAND2_X2 U12469 ( .A1(n15150), .A2(n13761), .ZN(n15163) );
  OR2_X1 U12471 ( .A1(n14754), .A2(n13563), .ZN(n20856) );
  XNOR2_X1 U12472 ( .A(n14760), .B(n12803), .ZN(n15170) );
  NAND2_X1 U12473 ( .A1(n10093), .A2(n14771), .ZN(n15185) );
  OR2_X1 U12474 ( .A1(n14770), .A2(n14772), .ZN(n10093) );
  NAND2_X1 U12475 ( .A1(n14861), .A2(n9647), .ZN(n14826) );
  INV_X1 U12476 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15300) );
  INV_X1 U12477 ( .A(n20881), .ZN(n15304) );
  AND3_X1 U12478 ( .A1(n10094), .A2(n10096), .A3(n10095), .ZN(n14173) );
  NAND2_X1 U12479 ( .A1(n21149), .A2(n12800), .ZN(n15382) );
  INV_X1 U12480 ( .A(n20882), .ZN(n15301) );
  NAND2_X1 U12481 ( .A1(n9909), .A2(n9672), .ZN(n9908) );
  NAND2_X1 U12482 ( .A1(n13004), .A2(n13007), .ZN(n15422) );
  AOI21_X1 U12483 ( .B1(n14790), .B2(n14789), .A(n14788), .ZN(n15424) );
  NAND2_X1 U12484 ( .A1(n12786), .A2(n12785), .ZN(n15188) );
  NAND2_X1 U12485 ( .A1(n9999), .A2(n10004), .ZN(n12785) );
  NAND2_X1 U12486 ( .A1(n9913), .A2(n9684), .ZN(n15447) );
  INV_X1 U12487 ( .A(n15459), .ZN(n9913) );
  OAI21_X1 U12488 ( .B1(n15237), .B2(n12778), .A(n15374), .ZN(n15238) );
  NAND2_X1 U12489 ( .A1(n12996), .A2(n15585), .ZN(n15474) );
  OR2_X1 U12490 ( .A1(n17200), .A2(n21388), .ZN(n17196) );
  NAND2_X1 U12491 ( .A1(n10164), .A2(n9688), .ZN(n17167) );
  OR2_X1 U12492 ( .A1(n20903), .A2(n15541), .ZN(n17200) );
  NAND2_X1 U12493 ( .A1(n17178), .A2(n12753), .ZN(n17172) );
  OR2_X1 U12494 ( .A1(n20936), .A2(n13008), .ZN(n20912) );
  AND2_X1 U12495 ( .A1(n20931), .A2(n12986), .ZN(n15583) );
  AND2_X1 U12496 ( .A1(n13030), .A2(n17084), .ZN(n20936) );
  NAND2_X1 U12497 ( .A1(n10166), .A2(n11811), .ZN(n11847) );
  INV_X1 U12498 ( .A(n12713), .ZN(n11838) );
  NAND2_X1 U12499 ( .A1(n10270), .A2(n13883), .ZN(n15634) );
  INV_X1 U12500 ( .A(n20951), .ZN(n14244) );
  NOR2_X1 U12501 ( .A1(n14066), .A2(n14088), .ZN(n14247) );
  OAI21_X1 U12502 ( .B1(n14075), .B2(n14073), .A(n14072), .ZN(n20954) );
  AND2_X1 U12503 ( .A1(n14077), .A2(n14076), .ZN(n20951) );
  OAI21_X1 U12504 ( .B1(n14192), .B2(n20966), .A(n21098), .ZN(n20969) );
  AOI22_X1 U12505 ( .A1(n15735), .A2(n15732), .B1(n15730), .B2(n15729), .ZN(
        n15773) );
  OAI21_X1 U12506 ( .B1(n14012), .B2(n14015), .A(n21147), .ZN(n14038) );
  INV_X1 U12507 ( .A(n14112), .ZN(n14147) );
  OAI211_X1 U12508 ( .C1(n21029), .C2(n14087), .A(n21147), .B(n14086), .ZN(
        n20988) );
  INV_X1 U12509 ( .A(n20995), .ZN(n21017) );
  OR2_X1 U12510 ( .A1(n21031), .A2(n21091), .ZN(n21044) );
  OAI211_X1 U12511 ( .C1(n21029), .C2(n21028), .A(n21147), .B(n21027), .ZN(
        n21050) );
  INV_X1 U12512 ( .A(n21044), .ZN(n21049) );
  OAI211_X1 U12513 ( .C1(n10548), .C2(n21064), .A(n21098), .B(n21063), .ZN(
        n21087) );
  INV_X1 U12514 ( .A(n21054), .ZN(n21085) );
  OAI211_X1 U12515 ( .C1(n21099), .C2(n21124), .A(n21098), .B(n21097), .ZN(
        n21128) );
  NOR2_X1 U12516 ( .A1(n15646), .A2(n15143), .ZN(n21139) );
  NOR2_X1 U12517 ( .A1(n15646), .A2(n13828), .ZN(n21155) );
  NOR2_X1 U12518 ( .A1(n15646), .A2(n15126), .ZN(n21167) );
  NOR2_X1 U12519 ( .A1(n15646), .A2(n15122), .ZN(n21173) );
  NOR2_X1 U12520 ( .A1(n15646), .A2(n15112), .ZN(n21185) );
  OR2_X1 U12521 ( .A1(n21140), .A2(n21091), .ZN(n21201) );
  INV_X1 U12522 ( .A(n21190), .ZN(n21197) );
  NOR2_X1 U12523 ( .A1(n15646), .A2(n15107), .ZN(n21195) );
  NAND2_X1 U12524 ( .A1(n17222), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21203) );
  INV_X1 U12525 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21064) );
  NOR2_X1 U12526 ( .A1(n16960), .A2(n12596), .ZN(n19715) );
  XNOR2_X1 U12527 ( .A(n11089), .B(n11090), .ZN(n15795) );
  INV_X1 U12528 ( .A(n11085), .ZN(n15821) );
  AOI21_X1 U12529 ( .B1(n15857), .B2(n9718), .A(n10245), .ZN(n15828) );
  AND2_X1 U12530 ( .A1(n11048), .A2(n11082), .ZN(n15851) );
  NAND2_X1 U12531 ( .A1(n11039), .A2(n10476), .ZN(n11047) );
  NOR2_X1 U12532 ( .A1(n19773), .A2(n12638), .ZN(n15911) );
  NAND2_X1 U12533 ( .A1(n15911), .A2(n15910), .ZN(n19745) );
  NOR2_X1 U12534 ( .A1(n15917), .A2(n12634), .ZN(n19787) );
  NAND2_X1 U12535 ( .A1(n19829), .A2(n9604), .ZN(n19809) );
  INV_X1 U12536 ( .A(n19864), .ZN(n19838) );
  NAND2_X1 U12537 ( .A1(n19829), .A2(n12628), .ZN(n19820) );
  NAND2_X1 U12538 ( .A1(n10984), .A2(n19837), .ZN(n11000) );
  INV_X1 U12539 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19879) );
  OR2_X1 U12540 ( .A1(n10959), .A2(n10673), .ZN(n10974) );
  NAND2_X1 U12541 ( .A1(n14184), .A2(n14183), .ZN(n14430) );
  NOR2_X1 U12542 ( .A1(n10454), .A2(n10458), .ZN(n14156) );
  OR2_X1 U12543 ( .A1(n10459), .A2(n14063), .ZN(n10454) );
  NAND2_X1 U12544 ( .A1(n10456), .A2(n10457), .ZN(n16136) );
  INV_X1 U12545 ( .A(n10459), .ZN(n10457) );
  OR2_X1 U12546 ( .A1(n11361), .A2(n11360), .ZN(n16152) );
  OR2_X1 U12547 ( .A1(n11345), .A2(n11344), .ZN(n14212) );
  INV_X1 U12548 ( .A(n9716), .ZN(n16150) );
  INV_X1 U12549 ( .A(n20664), .ZN(n16907) );
  AND2_X1 U12550 ( .A1(n14694), .A2(n16873), .ZN(n16259) );
  AND2_X1 U12551 ( .A1(n14184), .A2(n9725), .ZN(n16127) );
  NAND2_X1 U12552 ( .A1(n13566), .A2(n13567), .ZN(n10497) );
  AND2_X1 U12553 ( .A1(n16227), .A2(n16282), .ZN(n16275) );
  INV_X1 U12554 ( .A(n19896), .ZN(n16279) );
  OR2_X1 U12555 ( .A1(n13572), .A2(n13571), .ZN(n13573) );
  INV_X2 U12556 ( .A(n16287), .ZN(n19887) );
  INV_X1 U12557 ( .A(n16282), .ZN(n19888) );
  INV_X1 U12558 ( .A(n13528), .ZN(n19899) );
  NAND2_X1 U12559 ( .A1(n19933), .A2(n13529), .ZN(n19902) );
  INV_X1 U12560 ( .A(n19902), .ZN(n19931) );
  INV_X1 U12561 ( .A(n13402), .ZN(n19937) );
  INV_X1 U12562 ( .A(n13490), .ZN(n19938) );
  OAI211_X1 U12563 ( .C1(n16327), .C2(n9935), .A(n9928), .B(n9932), .ZN(n16566) );
  NAND2_X1 U12564 ( .A1(n16327), .A2(n9934), .ZN(n9928) );
  INV_X1 U12565 ( .A(n9966), .ZN(n14736) );
  NAND2_X1 U12566 ( .A1(n16502), .A2(n16547), .ZN(n10106) );
  NAND2_X1 U12567 ( .A1(n19725), .A2(n13551), .ZN(n19955) );
  CLKBUF_X1 U12568 ( .A(n16007), .Z(n16008) );
  INV_X1 U12569 ( .A(n10467), .ZN(n10466) );
  AND2_X1 U12570 ( .A1(n10532), .A2(n11517), .ZN(n11518) );
  INV_X1 U12571 ( .A(n9850), .ZN(n16296) );
  NAND2_X1 U12572 ( .A1(n16313), .A2(n16551), .ZN(n9851) );
  NAND2_X1 U12573 ( .A1(n9932), .A2(n9935), .ZN(n9931) );
  INV_X1 U12574 ( .A(n9934), .ZN(n9930) );
  INV_X1 U12575 ( .A(n16312), .ZN(n16314) );
  INV_X1 U12576 ( .A(n16327), .ZN(n16336) );
  NAND2_X1 U12577 ( .A1(n16362), .A2(n16361), .ZN(n16609) );
  AND2_X1 U12578 ( .A1(n10187), .A2(n10186), .ZN(n10185) );
  NAND2_X1 U12579 ( .A1(n16633), .A2(n19967), .ZN(n10187) );
  INV_X1 U12580 ( .A(n16632), .ZN(n10186) );
  CLKBUF_X1 U12581 ( .A(n14402), .Z(n14403) );
  NAND2_X1 U12582 ( .A1(n10215), .A2(n10213), .ZN(n14387) );
  NAND2_X1 U12583 ( .A1(n14389), .A2(n14359), .ZN(n10215) );
  NAND2_X1 U12584 ( .A1(n9868), .A2(n9867), .ZN(n16399) );
  NAND2_X1 U12585 ( .A1(n10298), .A2(n10296), .ZN(n16397) );
  NAND2_X1 U12586 ( .A1(n10301), .A2(n10300), .ZN(n9867) );
  INV_X1 U12587 ( .A(n9914), .ZN(n16464) );
  INV_X1 U12588 ( .A(n14360), .ZN(n16478) );
  AND2_X1 U12589 ( .A1(n10057), .A2(n10056), .ZN(n17233) );
  NOR2_X1 U12590 ( .A1(n13651), .A2(n17241), .ZN(n10056) );
  NAND2_X1 U12591 ( .A1(n9923), .A2(n16003), .ZN(n16542) );
  INV_X1 U12592 ( .A(n10057), .ZN(n13656) );
  INV_X1 U12593 ( .A(n17237), .ZN(n19956) );
  INV_X1 U12594 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19964) );
  INV_X1 U12595 ( .A(n20655), .ZN(n20656) );
  NAND2_X1 U12596 ( .A1(n20647), .A2(n20656), .ZN(n20629) );
  INV_X1 U12597 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17144) );
  CLKBUF_X1 U12598 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n21340) );
  NAND2_X1 U12599 ( .A1(n9754), .A2(n13475), .ZN(n16951) );
  AND2_X1 U12600 ( .A1(n20011), .A2(n20010), .ZN(n20029) );
  OAI211_X1 U12601 ( .C1(n20057), .C2(n20042), .A(n20041), .B(n20476), .ZN(
        n20059) );
  NAND2_X1 U12602 ( .A1(n20034), .A2(n20039), .ZN(n20058) );
  OAI21_X1 U12603 ( .B1(n20072), .B2(n20071), .A(n20070), .ZN(n20090) );
  NOR2_X1 U12604 ( .A1(n20174), .A2(n20630), .ZN(n20089) );
  OAI21_X1 U12605 ( .B1(n16893), .B2(n20628), .A(n16892), .ZN(n20108) );
  NOR2_X2 U12606 ( .A1(n20146), .A2(n20114), .ZN(n20134) );
  OAI21_X1 U12607 ( .B1(n20121), .B2(n20118), .A(n20117), .ZN(n20139) );
  NOR2_X1 U12608 ( .A1(n20174), .A2(n20114), .ZN(n20147) );
  AOI21_X1 U12609 ( .B1(n20463), .B2(n20145), .A(n20150), .ZN(n20169) );
  OR2_X1 U12610 ( .A1(n20181), .A2(n20178), .ZN(n20206) );
  OAI21_X1 U12611 ( .B1(n20237), .B2(n20218), .A(n20476), .ZN(n20239) );
  INV_X1 U12612 ( .A(n20293), .ZN(n20306) );
  OAI221_X1 U12613 ( .B1(n20322), .B2(n20321), .C1(n20322), .C2(n20472), .A(
        n20320), .ZN(n20341) );
  AOI21_X1 U12614 ( .B1(n20463), .B2(n20316), .A(n20319), .ZN(n20339) );
  NOR2_X1 U12615 ( .A1(n20369), .A2(n20634), .ZN(n9865) );
  AND2_X1 U12616 ( .A1(n19998), .A2(n10784), .ZN(n20407) );
  AND2_X1 U12617 ( .A1(n20476), .A2(n16881), .ZN(n20418) );
  INV_X1 U12618 ( .A(n20482), .ZN(n20408) );
  INV_X1 U12619 ( .A(n20489), .ZN(n20423) );
  AND2_X1 U12620 ( .A1(n19998), .A2(n19972), .ZN(n20422) );
  AND2_X1 U12621 ( .A1(n19998), .A2(n19989), .ZN(n20444) );
  OAI21_X1 U12622 ( .B1(n20417), .B2(n20416), .A(n20415), .ZN(n20457) );
  INV_X1 U12623 ( .A(n20421), .ZN(n20479) );
  INV_X1 U12624 ( .A(n20427), .ZN(n20486) );
  INV_X1 U12625 ( .A(n20433), .ZN(n20493) );
  INV_X1 U12626 ( .A(n20386), .ZN(n20507) );
  INV_X1 U12627 ( .A(n20449), .ZN(n20514) );
  INV_X1 U12628 ( .A(n20395), .ZN(n20521) );
  OR2_X1 U12629 ( .A1(n20473), .A2(n20467), .ZN(n20528) );
  INV_X1 U12630 ( .A(n20344), .ZN(n20530) );
  AOI211_X1 U12631 ( .C1(n16964), .C2(n16963), .A(n16962), .B(n16961), .ZN(
        n20537) );
  INV_X1 U12632 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n20690) );
  NAND2_X1 U12633 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20562), .ZN(n20700) );
  INV_X1 U12634 ( .A(n17062), .ZN(n18305) );
  INV_X1 U12635 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19696) );
  NOR2_X1 U12636 ( .A1(n10336), .A2(n19555), .ZN(n9976) );
  XNOR2_X1 U12637 ( .A(n17451), .B(n17452), .ZN(n10336) );
  OR2_X1 U12638 ( .A1(n17454), .A2(n17453), .ZN(n9975) );
  NOR2_X1 U12639 ( .A1(n17463), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n10335) );
  NOR2_X1 U12640 ( .A1(n17482), .A2(P3_EBX_REG_28__SCAN_IN), .ZN(n17468) );
  NOR2_X1 U12641 ( .A1(n17501), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n17487) );
  NAND2_X1 U12642 ( .A1(n17487), .A2(n17805), .ZN(n17482) );
  NOR2_X1 U12643 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17523), .ZN(n17506) );
  NOR2_X1 U12644 ( .A1(n17544), .A2(P3_EBX_REG_22__SCAN_IN), .ZN(n17532) );
  NAND2_X1 U12645 ( .A1(n17532), .A2(n17524), .ZN(n17523) );
  NAND2_X1 U12646 ( .A1(n17653), .A2(n10330), .ZN(n10329) );
  INV_X1 U12647 ( .A(n18451), .ZN(n10330) );
  OR2_X1 U12648 ( .A1(n17550), .A2(n17653), .ZN(n10334) );
  NOR2_X1 U12649 ( .A1(n17564), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n17548) );
  NAND2_X1 U12650 ( .A1(n17548), .A2(n17901), .ZN(n17544) );
  OAI21_X1 U12651 ( .B1(n17437), .B2(n17653), .A(n17594), .ZN(n17551) );
  NOR2_X1 U12652 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17584), .ZN(n17568) );
  NOR2_X1 U12653 ( .A1(n17601), .A2(P3_EBX_REG_16__SCAN_IN), .ZN(n17588) );
  NAND2_X1 U12654 ( .A1(n17588), .A2(n17953), .ZN(n17584) );
  OAI21_X1 U12655 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17600), .A(
        n17436), .ZN(n17594) );
  NOR2_X1 U12656 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17685), .ZN(n17666) );
  NAND2_X1 U12657 ( .A1(n17690), .A2(n17686), .ZN(n17685) );
  NOR2_X1 U12658 ( .A1(n17710), .A2(P3_EBX_REG_8__SCAN_IN), .ZN(n17690) );
  NOR2_X1 U12659 ( .A1(n17731), .A2(P3_EBX_REG_6__SCAN_IN), .ZN(n17716) );
  NAND2_X1 U12660 ( .A1(n17716), .A2(n17711), .ZN(n17710) );
  AND3_X1 U12661 ( .A1(n9973), .A2(n9972), .A3(n9971), .ZN(n17769) );
  INV_X1 U12662 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n9971) );
  NAND2_X1 U12663 ( .A1(n17769), .A2(n17765), .ZN(n17764) );
  NOR2_X2 U12664 ( .A1(n19540), .A2(n17421), .ZN(n17782) );
  INV_X1 U12665 ( .A(n17800), .ZN(n17787) );
  INV_X1 U12666 ( .A(n17782), .ZN(n17788) );
  NOR2_X1 U12667 ( .A1(n17814), .A2(n17813), .ZN(n17843) );
  NAND2_X1 U12668 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17863), .ZN(n17855) );
  AND2_X1 U12669 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17867), .ZN(n17863) );
  NOR2_X1 U12670 ( .A1(n17873), .A2(n17807), .ZN(n17867) );
  AND2_X1 U12671 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17886), .ZN(n17872) );
  NAND2_X1 U12672 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17899), .ZN(n17873) );
  NOR2_X1 U12673 ( .A1(n17864), .A2(n17873), .ZN(n17886) );
  AND2_X1 U12674 ( .A1(n17954), .A2(n10262), .ZN(n17899) );
  NOR2_X1 U12675 ( .A1(n18213), .A2(n10264), .ZN(n10262) );
  NAND2_X1 U12676 ( .A1(n17954), .A2(P3_EBX_REG_17__SCAN_IN), .ZN(n17937) );
  NAND2_X1 U12677 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17996), .ZN(n17981) );
  AND2_X1 U12678 ( .A1(n18055), .A2(n10268), .ZN(n17053) );
  AND2_X1 U12679 ( .A1(n9630), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n10268) );
  NAND2_X1 U12680 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17053), .ZN(n17983) );
  NAND2_X1 U12681 ( .A1(n18055), .A2(n9630), .ZN(n18022) );
  NAND2_X1 U12682 ( .A1(n18055), .A2(P3_EBX_REG_9__SCAN_IN), .ZN(n18053) );
  NAND3_X1 U12683 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(n18080), .ZN(n18056) );
  NOR2_X1 U12684 ( .A1(n18057), .A2(n18056), .ZN(n18055) );
  AND2_X1 U12685 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n18084), .ZN(n18080) );
  NOR2_X1 U12686 ( .A1(n18105), .A2(n18090), .ZN(n18084) );
  OR3_X1 U12687 ( .A1(n18088), .A2(n17765), .A3(n18087), .ZN(n18090) );
  INV_X1 U12688 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18100) );
  NAND2_X1 U12689 ( .A1(n17145), .A2(n10256), .ZN(n18105) );
  AND2_X1 U12690 ( .A1(n16967), .A2(n19700), .ZN(n10256) );
  NOR2_X2 U12691 ( .A1(n19084), .A2(n18105), .ZN(n18106) );
  NAND2_X1 U12692 ( .A1(n18118), .A2(n18177), .ZN(n18117) );
  NAND2_X1 U12693 ( .A1(n18123), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n18118) );
  AND2_X1 U12694 ( .A1(n18125), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n18123) );
  INV_X1 U12695 ( .A(n18128), .ZN(n18125) );
  NAND2_X1 U12696 ( .A1(n18141), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n18136) );
  NOR2_X1 U12697 ( .A1(n18213), .A2(n10191), .ZN(n10189) );
  NOR2_X1 U12698 ( .A1(n18310), .A2(n18176), .ZN(n18171) );
  OR3_X1 U12699 ( .A1(n18213), .A2(n18184), .A3(n18308), .ZN(n18176) );
  NOR2_X1 U12700 ( .A1(n18250), .A2(n9629), .ZN(n18193) );
  NAND2_X1 U12701 ( .A1(n10207), .A2(n10210), .ZN(n18219) );
  NOR2_X1 U12702 ( .A1(n18250), .A2(n18109), .ZN(n18224) );
  NOR2_X1 U12703 ( .A1(n18294), .A2(n18232), .ZN(n18235) );
  INV_X1 U12704 ( .A(n13101), .ZN(n18236) );
  INV_X1 U12705 ( .A(n13298), .ZN(n18241) );
  AND2_X1 U12706 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18240), .ZN(n18244) );
  INV_X1 U12707 ( .A(n18245), .ZN(n18249) );
  INV_X1 U12708 ( .A(n21311), .ZN(n18272) );
  CLKBUF_X1 U12709 ( .A(n18355), .Z(n18341) );
  INV_X1 U12710 ( .A(n18352), .ZN(n18358) );
  INV_X1 U12711 ( .A(n10158), .ZN(n17281) );
  AOI21_X1 U12712 ( .B1(n18374), .B2(n18373), .A(n18372), .ZN(n18379) );
  OR2_X1 U12713 ( .A1(n18371), .A2(n18370), .ZN(n18372) );
  AND2_X1 U12714 ( .A1(n18446), .A2(n10322), .ZN(n18433) );
  INV_X1 U12715 ( .A(n18447), .ZN(n10322) );
  INV_X1 U12716 ( .A(n18531), .ZN(n18459) );
  NAND2_X1 U12717 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18524) );
  INV_X1 U12718 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18581) );
  NOR2_X1 U12719 ( .A1(n17738), .A2(n10338), .ZN(n10339) );
  INV_X1 U12720 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18652) );
  INV_X1 U12721 ( .A(n19335), .ZN(n19427) );
  INV_X1 U12722 ( .A(n18715), .ZN(n18707) );
  INV_X1 U12723 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19656) );
  OR2_X1 U12724 ( .A1(n13360), .A2(n19006), .ZN(n13375) );
  AOI21_X1 U12725 ( .B1(n10158), .B2(n19040), .A(n10155), .ZN(n17137) );
  INV_X1 U12726 ( .A(n10156), .ZN(n10155) );
  AOI21_X1 U12727 ( .B1(n17260), .B2(n18961), .A(n10157), .ZN(n10156) );
  INV_X1 U12728 ( .A(n18851), .ZN(n18954) );
  NAND2_X1 U12729 ( .A1(n18427), .A2(n13148), .ZN(n18418) );
  INV_X1 U12730 ( .A(n10039), .ZN(n18417) );
  NAND2_X1 U12731 ( .A1(n18504), .A2(n13150), .ZN(n18428) );
  INV_X1 U12732 ( .A(n18852), .ZN(n18831) );
  NOR2_X1 U12733 ( .A1(n18852), .A2(n10084), .ZN(n18840) );
  OR2_X1 U12734 ( .A1(n18832), .A2(n18833), .ZN(n10084) );
  OR2_X1 U12735 ( .A1(n18801), .A2(n19026), .ZN(n18852) );
  INV_X1 U12736 ( .A(n13146), .ZN(n18519) );
  OAI21_X1 U12737 ( .B1(n18623), .B2(n10080), .A(n10079), .ZN(n18859) );
  AOI21_X1 U12738 ( .B1(n13323), .B2(n18957), .A(n18780), .ZN(n10079) );
  INV_X1 U12739 ( .A(n13323), .ZN(n10080) );
  OR2_X1 U12740 ( .A1(n13288), .A2(n19482), .ZN(n9941) );
  NOR2_X2 U12741 ( .A1(n19512), .A2(n19032), .ZN(n18929) );
  NOR2_X1 U12742 ( .A1(n17287), .A2(n19035), .ZN(n18961) );
  INV_X1 U12743 ( .A(n18643), .ZN(n10076) );
  NAND2_X1 U12744 ( .A1(n10307), .A2(n9748), .ZN(n18661) );
  AND2_X1 U12745 ( .A1(n10307), .A2(n10305), .ZN(n18662) );
  INV_X1 U12746 ( .A(n19032), .ZN(n19501) );
  INV_X1 U12747 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19195) );
  NOR2_X1 U12748 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19650), .ZN(
        n19671) );
  AOI211_X1 U12749 ( .C1(n19700), .C2(n19534), .A(n19055), .B(n17070), .ZN(
        n19677) );
  INV_X1 U12750 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n21439) );
  INV_X1 U12751 ( .A(n19677), .ZN(n19675) );
  NOR2_X1 U12752 ( .A1(n9942), .A2(n19536), .ZN(n19548) );
  NAND2_X1 U12753 ( .A1(n9943), .A2(n9675), .ZN(n9942) );
  AND2_X2 U12754 ( .A1(n12589), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n15085)
         );
  CLKBUF_X1 U12755 ( .A(n17383), .Z(n17385) );
  NAND2_X1 U12756 ( .A1(n10050), .A2(n9670), .ZN(P1_U2809) );
  NAND2_X1 U12757 ( .A1(n9877), .A2(n9685), .ZN(P1_U2968) );
  NAND2_X1 U12758 ( .A1(n10275), .A2(n10274), .ZN(n15408) );
  OAI21_X1 U12759 ( .B1(n15417), .B2(n20712), .A(n10090), .ZN(P1_U2971) );
  INV_X1 U12760 ( .A(n10091), .ZN(n10090) );
  OAI21_X1 U12761 ( .B1(n15185), .B2(n15382), .A(n10092), .ZN(n10091) );
  AOI21_X1 U12762 ( .B1(n15304), .B2(n15187), .A(n15186), .ZN(n10092) );
  INV_X1 U12763 ( .A(n9909), .ZN(n15395) );
  AND2_X1 U12764 ( .A1(n15407), .A2(n15406), .ZN(n10278) );
  OAI21_X1 U12765 ( .B1(n12676), .B2(n16046), .A(n10239), .ZN(P2_U2824) );
  INV_X1 U12766 ( .A(n10240), .ZN(n10239) );
  OAI211_X1 U12767 ( .C1(n14747), .C2(n19871), .A(n9691), .B(n10241), .ZN(
        n10240) );
  INV_X1 U12768 ( .A(n12679), .ZN(n12694) );
  AOI21_X1 U12769 ( .B1(n15777), .B2(n19768), .A(n10412), .ZN(n10411) );
  NAND2_X1 U12770 ( .A1(n9656), .A2(n10413), .ZN(n10412) );
  OAI21_X1 U12771 ( .B1(n10144), .B2(n10143), .A(n14750), .ZN(P2_U2983) );
  INV_X1 U12772 ( .A(n10356), .ZN(n10143) );
  AOI21_X1 U12773 ( .B1(n16585), .B2(n16547), .A(n16332), .ZN(n9980) );
  NAND2_X1 U12774 ( .A1(n9696), .A2(n19945), .ZN(n9979) );
  AOI21_X1 U12775 ( .B1(n16607), .B2(n16547), .A(n16352), .ZN(n9828) );
  OAI21_X1 U12776 ( .B1(n16351), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n9774), .ZN(n9773) );
  OAI21_X1 U12777 ( .B1(n16631), .B2(n10135), .A(n10132), .ZN(P2_U2992) );
  OR2_X1 U12778 ( .A1(n16630), .A2(n16550), .ZN(n10135) );
  INV_X1 U12779 ( .A(n10133), .ZN(n10132) );
  INV_X1 U12780 ( .A(n9853), .ZN(n16387) );
  AOI21_X1 U12781 ( .B1(n16645), .B2(n16547), .A(n16386), .ZN(n9854) );
  INV_X1 U12782 ( .A(n9964), .ZN(n9963) );
  AOI21_X1 U12783 ( .B1(n16682), .B2(n16547), .A(n16423), .ZN(n9965) );
  INV_X1 U12784 ( .A(n9856), .ZN(n16446) );
  AOI21_X1 U12785 ( .B1(n16445), .B2(n16547), .A(n16444), .ZN(n9857) );
  NAND2_X1 U12786 ( .A1(n10034), .A2(n9970), .ZN(P2_U3020) );
  NAND2_X1 U12787 ( .A1(n10035), .A2(n19958), .ZN(n10034) );
  AND2_X1 U12788 ( .A1(n16312), .A2(n9845), .ZN(n9844) );
  OAI21_X1 U12789 ( .B1(n16608), .B2(n16802), .A(n9800), .ZN(P2_U3022) );
  AND2_X1 U12790 ( .A1(n9583), .A2(n16799), .ZN(n9884) );
  INV_X1 U12791 ( .A(n9882), .ZN(n9801) );
  OAI21_X1 U12792 ( .B1(n16631), .B2(n10188), .A(n10183), .ZN(P2_U3024) );
  INV_X1 U12793 ( .A(n10184), .ZN(n10183) );
  OR2_X1 U12794 ( .A1(n16630), .A2(n19970), .ZN(n10188) );
  OAI21_X1 U12795 ( .B1(n16634), .B2(n16802), .A(n10185), .ZN(n10184) );
  INV_X1 U12796 ( .A(n9864), .ZN(n16646) );
  NAND2_X1 U12797 ( .A1(n9959), .A2(n9956), .ZN(n14729) );
  OAI21_X1 U12798 ( .B1(n16693), .B2(n16802), .A(n10043), .ZN(P2_U3032) );
  NOR2_X1 U12799 ( .A1(n16691), .A2(n10045), .ZN(n10044) );
  NAND2_X1 U12800 ( .A1(n9766), .A2(n16799), .ZN(n16702) );
  NOR2_X1 U12801 ( .A1(n16712), .A2(n10252), .ZN(n10251) );
  OAI211_X1 U12802 ( .C1(n9652), .C2(n16757), .A(n10127), .B(n10126), .ZN(
        P2_U3038) );
  NOR2_X1 U12803 ( .A1(n16759), .A2(n10128), .ZN(n10127) );
  OR2_X1 U12804 ( .A1(n16761), .A2(n16802), .ZN(n10126) );
  AOI211_X1 U12805 ( .C1(n17455), .C2(n17814), .A(n17447), .B(n17446), .ZN(
        n17448) );
  NAND2_X1 U12806 ( .A1(n9977), .A2(n9974), .ZN(P3_U2641) );
  NAND2_X1 U12807 ( .A1(n9978), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9977) );
  NOR3_X1 U12808 ( .A1(n10335), .A2(n9976), .A3(n9975), .ZN(n9974) );
  OR2_X1 U12809 ( .A1(n17455), .A2(n17800), .ZN(n9978) );
  NAND2_X1 U12810 ( .A1(n18188), .A2(n10190), .ZN(n18146) );
  AND2_X1 U12811 ( .A1(n13345), .A2(n13344), .ZN(n13346) );
  INV_X2 U12812 ( .A(n12287), .ZN(n11795) );
  NAND2_X1 U12813 ( .A1(n12605), .A2(n12604), .ZN(n19866) );
  AND2_X1 U12814 ( .A1(n14352), .A2(n16417), .ZN(n9600) );
  CLKBUF_X3 U12815 ( .A(n13202), .Z(n17041) );
  AND2_X1 U12816 ( .A1(n10100), .A2(n12983), .ZN(n9601) );
  AND2_X1 U12817 ( .A1(n9600), .A2(n10221), .ZN(n10220) );
  AND2_X1 U12818 ( .A1(n14062), .A2(n9612), .ZN(n9602) );
  INV_X1 U12819 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19954) );
  AND3_X2 U12820 ( .A1(n10715), .A2(n10714), .A3(n10713), .ZN(n11542) );
  AND2_X1 U12821 ( .A1(n13336), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9603) );
  AND2_X1 U12822 ( .A1(n9624), .A2(n19811), .ZN(n9604) );
  NAND2_X2 U12823 ( .A1(n13823), .A2(n13777), .ZN(n12832) );
  CLKBUF_X3 U12824 ( .A(n10631), .Z(n14532) );
  NAND2_X1 U12825 ( .A1(n10444), .A2(n10442), .ZN(n14279) );
  NAND2_X1 U12826 ( .A1(n9799), .A2(n9841), .ZN(n9605) );
  AND2_X1 U12827 ( .A1(n14861), .A2(n9653), .ZN(n9606) );
  NAND2_X1 U12828 ( .A1(n14861), .A2(n14862), .ZN(n14850) );
  AND2_X1 U12829 ( .A1(n15854), .A2(n15856), .ZN(n15841) );
  OAI21_X1 U12830 ( .B1(n11994), .B2(n10089), .A(n10087), .ZN(n14939) );
  NOR2_X1 U12831 ( .A1(n16013), .A2(n12624), .ZN(n12623) );
  AND2_X1 U12832 ( .A1(n12520), .A2(n12555), .ZN(n9607) );
  OR2_X1 U12833 ( .A1(n13934), .A2(n10512), .ZN(n14725) );
  INV_X1 U12834 ( .A(n9655), .ZN(n10118) );
  NOR2_X1 U12835 ( .A1(n13934), .A2(n14162), .ZN(n9608) );
  INV_X1 U12836 ( .A(n10316), .ZN(n12561) );
  AND2_X1 U12837 ( .A1(n11508), .A2(n9671), .ZN(n9609) );
  AND2_X1 U12838 ( .A1(n11197), .A2(n10487), .ZN(n9610) );
  AND3_X1 U12839 ( .A1(n16377), .A2(n16379), .A3(n11040), .ZN(n9611) );
  INV_X1 U12840 ( .A(n11541), .ZN(n9765) );
  AND2_X1 U12841 ( .A1(n12753), .A2(n9988), .ZN(n10318) );
  AND2_X1 U12842 ( .A1(n14061), .A2(n9735), .ZN(n9612) );
  AND2_X1 U12843 ( .A1(n10799), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n9613) );
  INV_X1 U12844 ( .A(n15777), .ZN(n16562) );
  OR2_X1 U12845 ( .A1(n12531), .A2(n12530), .ZN(n9614) );
  AND2_X1 U12846 ( .A1(n12972), .A2(n13839), .ZN(n9615) );
  AND2_X1 U12847 ( .A1(n9694), .A2(n10219), .ZN(n9616) );
  AND2_X1 U12848 ( .A1(n9662), .A2(n14816), .ZN(n9617) );
  INV_X1 U12849 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12624) );
  INV_X1 U12850 ( .A(n16405), .ZN(n10301) );
  OR2_X1 U12851 ( .A1(n15897), .A2(n10234), .ZN(n12642) );
  INV_X1 U12852 ( .A(n12642), .ZN(n10385) );
  INV_X1 U12853 ( .A(n10511), .ZN(n16256) );
  AND2_X1 U12854 ( .A1(n10344), .A2(n10342), .ZN(n9618) );
  AND2_X1 U12855 ( .A1(n9610), .A2(n16147), .ZN(n9619) );
  AND2_X1 U12856 ( .A1(n9767), .A2(n9732), .ZN(n9620) );
  NAND2_X1 U12857 ( .A1(n13650), .A2(n9726), .ZN(n15981) );
  NAND4_X1 U12858 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A4(n10392), .ZN(n12620) );
  NAND2_X1 U12859 ( .A1(n10427), .A2(n10426), .ZN(n14175) );
  INV_X1 U12860 ( .A(n10456), .ZN(n10458) );
  NAND2_X1 U12861 ( .A1(n12641), .A2(n10398), .ZN(n9621) );
  AND2_X1 U12862 ( .A1(n10398), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9622) );
  AND2_X1 U12863 ( .A1(n10520), .A2(n10518), .ZN(n9623) );
  AND2_X1 U12864 ( .A1(n12628), .A2(n16466), .ZN(n9624) );
  AND3_X1 U12865 ( .A1(n13317), .A2(n10076), .A3(n18655), .ZN(n9625) );
  AND2_X1 U12866 ( .A1(n12656), .A2(n9747), .ZN(n12658) );
  NAND2_X1 U12867 ( .A1(n11917), .A2(n11882), .ZN(n15658) );
  AND2_X1 U12868 ( .A1(n14463), .A2(n10463), .ZN(n9626) );
  AND2_X1 U12869 ( .A1(n10436), .A2(n10435), .ZN(n9627) );
  AND2_X1 U12870 ( .A1(n9604), .A2(n16442), .ZN(n9628) );
  NAND2_X1 U12871 ( .A1(n10210), .A2(n9752), .ZN(n9629) );
  AND2_X1 U12872 ( .A1(n10269), .A2(P3_EBX_REG_11__SCAN_IN), .ZN(n9630) );
  AND2_X1 U12873 ( .A1(n11547), .A2(n16602), .ZN(n9631) );
  NAND2_X1 U12874 ( .A1(n13150), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9632) );
  AND4_X1 U12875 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .A4(P3_EAX_REG_10__SCAN_IN), .ZN(n9633)
         );
  NOR2_X2 U12876 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20634) );
  AND2_X1 U12877 ( .A1(n14722), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9634) );
  AND2_X2 U12878 ( .A1(n16832), .A2(n14507), .ZN(n10621) );
  AND2_X2 U12879 ( .A1(n14507), .A2(n10567), .ZN(n10623) );
  AND2_X1 U12880 ( .A1(n13875), .A2(n10876), .ZN(n9635) );
  AND2_X1 U12881 ( .A1(n16345), .A2(n16344), .ZN(n9636) );
  NAND2_X1 U12882 ( .A1(n16315), .A2(n11087), .ZN(n10026) );
  AND2_X1 U12883 ( .A1(n14861), .A2(n10447), .ZN(n14840) );
  NAND2_X1 U12884 ( .A1(n10519), .A2(n9623), .ZN(n9637) );
  OR2_X1 U12885 ( .A1(n16130), .A2(n10483), .ZN(n9638) );
  OR2_X1 U12886 ( .A1(n14784), .A2(n10450), .ZN(n9639) );
  NOR2_X1 U12887 ( .A1(n14939), .A2(n14940), .ZN(n14873) );
  NAND2_X1 U12888 ( .A1(n14861), .A2(n9617), .ZN(n14804) );
  AND2_X1 U12889 ( .A1(n14853), .A2(n9627), .ZN(n9640) );
  NOR2_X1 U12890 ( .A1(n14264), .A2(n14271), .ZN(n14270) );
  AND2_X1 U12891 ( .A1(n10246), .A2(n10247), .ZN(n9641) );
  AND2_X1 U12892 ( .A1(n10138), .A2(n10367), .ZN(n11480) );
  NOR2_X1 U12893 ( .A1(n12618), .A2(n16493), .ZN(n12619) );
  NAND2_X1 U12894 ( .A1(n15854), .A2(n10493), .ZN(n15824) );
  AND2_X1 U12895 ( .A1(n16120), .A2(n9626), .ZN(n9642) );
  NOR2_X1 U12896 ( .A1(n20756), .A2(n20755), .ZN(n9643) );
  AND2_X1 U12897 ( .A1(n10394), .A2(n10393), .ZN(n12622) );
  AND4_X1 U12898 ( .A1(n11600), .A2(n11599), .A3(n11598), .A4(n11597), .ZN(
        n9644) );
  INV_X1 U12899 ( .A(n12352), .ZN(n12495) );
  INV_X2 U12900 ( .A(n12495), .ZN(n12302) );
  AND2_X2 U12901 ( .A1(n11552), .A2(n15666), .ZN(n12352) );
  INV_X2 U12902 ( .A(n12321), .ZN(n11804) );
  NAND2_X1 U12903 ( .A1(n9785), .A2(n13860), .ZN(n13859) );
  INV_X1 U12904 ( .A(n10085), .ZN(n13297) );
  OR2_X1 U12905 ( .A1(n13071), .A2(n13070), .ZN(n10085) );
  INV_X1 U12906 ( .A(n11332), .ZN(n11333) );
  OR2_X1 U12907 ( .A1(n9583), .A2(n16578), .ZN(n9645) );
  NAND2_X1 U12908 ( .A1(n14706), .A2(n14710), .ZN(n14355) );
  AND4_X1 U12909 ( .A1(n13190), .A2(n13189), .A3(n13188), .A4(n13187), .ZN(
        n9646) );
  INV_X1 U12910 ( .A(n10123), .ZN(n10122) );
  NOR2_X1 U12911 ( .A1(n15374), .A2(n12779), .ZN(n10123) );
  AND2_X1 U12912 ( .A1(n10447), .A2(n14841), .ZN(n9647) );
  AND2_X1 U12913 ( .A1(n14993), .A2(n14977), .ZN(n9648) );
  AND2_X1 U12914 ( .A1(n9648), .A2(n10433), .ZN(n9649) );
  INV_X1 U12915 ( .A(n14359), .ZN(n10218) );
  OR3_X1 U12916 ( .A1(n14773), .A2(n12910), .A3(n14776), .ZN(n9650) );
  AND2_X1 U12917 ( .A1(n9919), .A2(n9921), .ZN(n9651) );
  OR2_X1 U12918 ( .A1(n16758), .A2(n19970), .ZN(n9652) );
  AND2_X1 U12919 ( .A1(n9617), .A2(n10098), .ZN(n9653) );
  INV_X1 U12920 ( .A(n18381), .ZN(n9821) );
  AND2_X1 U12921 ( .A1(n10369), .A2(n10522), .ZN(n9654) );
  OR2_X1 U12922 ( .A1(n15366), .A2(n15467), .ZN(n9655) );
  INV_X1 U12923 ( .A(n10362), .ZN(n10361) );
  OR2_X1 U12924 ( .A1(n15782), .A2(n19860), .ZN(n9656) );
  AND2_X1 U12925 ( .A1(n13146), .A2(n13145), .ZN(n9657) );
  OR2_X1 U12926 ( .A1(n18663), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9658) );
  AND2_X1 U12927 ( .A1(n16585), .A2(n19967), .ZN(n9659) );
  AND2_X1 U12928 ( .A1(n18247), .A2(n10085), .ZN(n9660) );
  INV_X1 U12929 ( .A(n20688), .ZN(n19972) );
  INV_X1 U12930 ( .A(n10785), .ZN(n11280) );
  NAND2_X1 U12931 ( .A1(n11016), .A2(n10027), .ZN(n9661) );
  AND2_X1 U12932 ( .A1(n9647), .A2(n10446), .ZN(n9662) );
  NOR2_X1 U12933 ( .A1(n12618), .A2(n10405), .ZN(n12616) );
  INV_X1 U12934 ( .A(n18464), .ZN(n10333) );
  AND2_X1 U12935 ( .A1(n9636), .A2(n16361), .ZN(n9663) );
  OR2_X1 U12936 ( .A1(n17134), .A2(n18634), .ZN(n9664) );
  OR2_X1 U12937 ( .A1(n17211), .A2(n11759), .ZN(n9665) );
  INV_X1 U12938 ( .A(n10114), .ZN(n12788) );
  AND2_X1 U12939 ( .A1(n19515), .A2(n19514), .ZN(n9666) );
  AND2_X1 U12940 ( .A1(n11102), .A2(n10358), .ZN(n9667) );
  NAND2_X1 U12941 ( .A1(n17073), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17072) );
  AND2_X1 U12942 ( .A1(n11310), .A2(n10500), .ZN(n9668) );
  AND2_X1 U12943 ( .A1(n15321), .A2(n15343), .ZN(n9669) );
  AND3_X1 U12944 ( .A1(n10049), .A2(n12956), .A3(n10047), .ZN(n9670) );
  NAND2_X1 U12945 ( .A1(n18443), .A2(n18721), .ZN(n18441) );
  OR2_X1 U12946 ( .A1(n19961), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9671) );
  AND2_X1 U12947 ( .A1(n13007), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9672) );
  AND2_X1 U12948 ( .A1(n16645), .A2(n19967), .ZN(n9673) );
  AND2_X1 U12949 ( .A1(n11719), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9674) );
  NOR2_X1 U12950 ( .A1(n19689), .A2(n19535), .ZN(n9675) );
  NOR2_X1 U12951 ( .A1(n14252), .A2(n14179), .ZN(n9676) );
  INV_X1 U12952 ( .A(n10835), .ZN(n11247) );
  AND2_X1 U12953 ( .A1(n11169), .A2(n10799), .ZN(n10835) );
  NAND2_X1 U12954 ( .A1(n10855), .A2(n10860), .ZN(n14344) );
  OR2_X1 U12955 ( .A1(n11022), .A2(n10019), .ZN(n9677) );
  INV_X1 U12956 ( .A(n11008), .ZN(n10291) );
  NOR2_X1 U12957 ( .A1(n13274), .A2(n13273), .ZN(n9678) );
  AND2_X1 U12958 ( .A1(n20688), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9679) );
  AND2_X1 U12959 ( .A1(n10119), .A2(n15448), .ZN(n9680) );
  AND2_X1 U12960 ( .A1(n13355), .A2(n19074), .ZN(n9681) );
  AND2_X1 U12961 ( .A1(n18643), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9682) );
  NAND2_X1 U12962 ( .A1(n11016), .A2(n11015), .ZN(n11011) );
  AND2_X1 U12963 ( .A1(n16443), .A2(n16694), .ZN(n9683) );
  NAND2_X1 U12964 ( .A1(n20891), .A2(n15448), .ZN(n9684) );
  AND2_X1 U12965 ( .A1(n12801), .A2(n12799), .ZN(n9685) );
  NAND2_X1 U12966 ( .A1(n16519), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9686) );
  NOR2_X1 U12967 ( .A1(n16317), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9687) );
  AND2_X1 U12968 ( .A1(n10317), .A2(n12763), .ZN(n9688) );
  NAND2_X1 U12969 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13044) );
  NAND2_X1 U12970 ( .A1(n10758), .A2(n10757), .ZN(n10800) );
  AND2_X1 U12971 ( .A1(n10352), .A2(n19958), .ZN(n9689) );
  INV_X1 U12972 ( .A(n10788), .ZN(n16914) );
  INV_X1 U12973 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12613) );
  OR2_X1 U12974 ( .A1(n16606), .A2(n9890), .ZN(n9690) );
  NAND2_X1 U12975 ( .A1(n12673), .A2(n19832), .ZN(n9691) );
  OR2_X1 U12976 ( .A1(n16584), .A2(n9659), .ZN(n9692) );
  NAND2_X1 U12977 ( .A1(n11994), .A2(n11993), .ZN(n14264) );
  INV_X1 U12978 ( .A(n10101), .ZN(n15180) );
  INV_X1 U12979 ( .A(n10297), .ZN(n10296) );
  NAND2_X1 U12980 ( .A1(n16398), .A2(n10301), .ZN(n10297) );
  OR2_X1 U12981 ( .A1(n12555), .A2(n12537), .ZN(n9693) );
  INV_X1 U12982 ( .A(n10046), .ZN(n9810) );
  NAND2_X1 U12983 ( .A1(n16422), .A2(n10373), .ZN(n10046) );
  AND2_X1 U12984 ( .A1(n14354), .A2(n10416), .ZN(n9694) );
  NAND2_X1 U12985 ( .A1(n10786), .A2(n20276), .ZN(n9695) );
  AND2_X1 U12986 ( .A1(n9847), .A2(n9843), .ZN(n9696) );
  NAND2_X1 U12987 ( .A1(n14853), .A2(n14843), .ZN(n14828) );
  INV_X1 U12988 ( .A(n11074), .ZN(n10363) );
  INV_X1 U12989 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16493) );
  OR2_X1 U12990 ( .A1(n16315), .A2(n9936), .ZN(n9697) );
  INV_X1 U12991 ( .A(n11811), .ZN(n9986) );
  INV_X1 U12992 ( .A(n16517), .ZN(n10372) );
  NAND2_X1 U12993 ( .A1(n10247), .A2(n16331), .ZN(n9698) );
  AND2_X1 U12994 ( .A1(n16344), .A2(n16333), .ZN(n9700) );
  OR2_X1 U12995 ( .A1(n19961), .A2(n11549), .ZN(n9701) );
  AND2_X1 U12996 ( .A1(n11918), .A2(n11942), .ZN(n9702) );
  NOR2_X1 U12997 ( .A1(n13620), .A2(n12985), .ZN(n9703) );
  INV_X1 U12998 ( .A(n10804), .ZN(n9799) );
  AND2_X1 U12999 ( .A1(n10148), .A2(n16344), .ZN(n9704) );
  NOR2_X1 U13000 ( .A1(n16644), .A2(n9673), .ZN(n9705) );
  OR2_X1 U13001 ( .A1(n11011), .A2(n10471), .ZN(n9706) );
  AND2_X1 U13002 ( .A1(n15283), .A2(n12775), .ZN(n9707) );
  OR2_X1 U13003 ( .A1(n12727), .A2(n11862), .ZN(n9708) );
  AND2_X1 U13004 ( .A1(n11712), .A2(n13621), .ZN(n9709) );
  NAND2_X1 U13005 ( .A1(n15353), .A2(n15430), .ZN(n9710) );
  AND2_X1 U13006 ( .A1(n10301), .A2(n9600), .ZN(n9711) );
  AND2_X1 U13007 ( .A1(n9649), .A2(n10432), .ZN(n9712) );
  AND2_X1 U13008 ( .A1(n10328), .A2(n10327), .ZN(n9713) );
  AND2_X1 U13009 ( .A1(n16367), .A2(n10364), .ZN(n9714) );
  INV_X1 U13010 ( .A(n13839), .ZN(n13636) );
  INV_X1 U13011 ( .A(n12704), .ZN(n10285) );
  NAND2_X1 U13012 ( .A1(n10075), .A2(n10073), .ZN(n13319) );
  NAND2_X1 U13013 ( .A1(n18643), .A2(n18642), .ZN(n9715) );
  INV_X2 U13014 ( .A(n18106), .ZN(n18101) );
  OR2_X1 U13015 ( .A1(n16154), .A2(n9832), .ZN(n9716) );
  INV_X1 U13016 ( .A(n19027), .ZN(n10157) );
  NOR2_X1 U13017 ( .A1(n14097), .A2(n14098), .ZN(n9717) );
  NAND2_X1 U13018 ( .A1(n14919), .A2(n14920), .ZN(n14903) );
  AND2_X1 U13019 ( .A1(n16350), .A2(n16356), .ZN(n9718) );
  OR2_X1 U13020 ( .A1(n12636), .A2(n10408), .ZN(n9719) );
  AND2_X1 U13021 ( .A1(n18141), .A2(n10201), .ZN(n9720) );
  NOR2_X1 U13022 ( .A1(n10431), .A2(n14904), .ZN(n9721) );
  NOR2_X1 U13023 ( .A1(n16130), .A2(n16131), .ZN(n14051) );
  AND2_X1 U13024 ( .A1(n15374), .A2(n10277), .ZN(n9722) );
  AND2_X1 U13025 ( .A1(n10903), .A2(n10920), .ZN(n9723) );
  NAND2_X1 U13026 ( .A1(n14994), .A2(n9648), .ZN(n14959) );
  AND2_X1 U13027 ( .A1(n12641), .A2(n10397), .ZN(n12647) );
  AND2_X1 U13028 ( .A1(n10490), .A2(n15801), .ZN(n9724) );
  NAND2_X1 U13029 ( .A1(n15963), .A2(n11329), .ZN(n13566) );
  AND2_X1 U13030 ( .A1(n14183), .A2(n10461), .ZN(n9725) );
  NOR2_X1 U13031 ( .A1(n16130), .A2(n10485), .ZN(n14050) );
  AND2_X1 U13032 ( .A1(n14994), .A2(n14993), .ZN(n14976) );
  INV_X1 U13033 ( .A(n17099), .ZN(n10051) );
  AOI21_X1 U13034 ( .B1(n12764), .B2(n12107), .A(n11975), .ZN(n14258) );
  AND2_X1 U13035 ( .A1(n14099), .A2(n14100), .ZN(n13928) );
  NOR2_X1 U13036 ( .A1(n12620), .A2(n19879), .ZN(n12621) );
  AND2_X1 U13037 ( .A1(n18188), .A2(n10189), .ZN(n18140) );
  INV_X1 U13038 ( .A(n10973), .ZN(n10016) );
  NAND2_X1 U13039 ( .A1(n10497), .A2(n11332), .ZN(n13592) );
  INV_X1 U13040 ( .A(n19861), .ZN(n10222) );
  OR2_X1 U13041 ( .A1(n21203), .A2(n11759), .ZN(n20710) );
  INV_X1 U13042 ( .A(n20710), .ZN(n9905) );
  INV_X1 U13043 ( .A(n11012), .ZN(n10474) );
  AND2_X1 U13044 ( .A1(n11310), .A2(n11318), .ZN(n9726) );
  AND2_X1 U13045 ( .A1(n17954), .A2(n10266), .ZN(n9727) );
  NOR2_X1 U13046 ( .A1(n16540), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9728) );
  OR2_X1 U13047 ( .A1(n13934), .A2(n10514), .ZN(n10511) );
  NAND2_X1 U13048 ( .A1(n19970), .A2(n14712), .ZN(n9729) );
  AND2_X1 U13049 ( .A1(n12656), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12655) );
  INV_X1 U13050 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16013) );
  OR2_X1 U13051 ( .A1(n20681), .A2(n20660), .ZN(n9730) );
  AND2_X1 U13052 ( .A1(n18188), .A2(n10192), .ZN(n9731) );
  AND2_X1 U13053 ( .A1(n10106), .A2(n10105), .ZN(n9732) );
  NAND2_X1 U13054 ( .A1(n11860), .A2(n11859), .ZN(n13883) );
  OR2_X1 U13055 ( .A1(n19989), .A2(n11219), .ZN(n9733) );
  OR2_X1 U13056 ( .A1(n10286), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9734) );
  AND2_X1 U13057 ( .A1(n10455), .A2(n14155), .ZN(n9735) );
  AND2_X1 U13058 ( .A1(n10462), .A2(n14506), .ZN(n9736) );
  INV_X1 U13059 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13621) );
  INV_X1 U13060 ( .A(n10300), .ZN(n10299) );
  NAND2_X1 U13061 ( .A1(n16418), .A2(n16406), .ZN(n10300) );
  NAND2_X1 U13062 ( .A1(n10315), .A2(n17109), .ZN(n9737) );
  NAND2_X1 U13063 ( .A1(n11628), .A2(n11707), .ZN(n10114) );
  INV_X1 U13064 ( .A(n10794), .ZN(n13585) );
  AND2_X1 U13065 ( .A1(n9723), .A2(n11535), .ZN(n9738) );
  NOR2_X1 U13066 ( .A1(n14892), .A2(n14878), .ZN(n14865) );
  AND2_X1 U13067 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n9739) );
  OAI221_X1 U13068 ( .B1(n17147), .B2(n17146), .C1(n17147), .C2(n17145), .A(
        n19700), .ZN(n18250) );
  NOR2_X1 U13069 ( .A1(n19989), .A2(n11223), .ZN(n11023) );
  XOR2_X1 U13070 ( .A(n15172), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n9740) );
  AND2_X1 U13071 ( .A1(n10719), .A2(n11032), .ZN(n9741) );
  AND2_X1 U13072 ( .A1(n9721), .A2(n10430), .ZN(n9742) );
  AND2_X1 U13073 ( .A1(n9725), .A2(n16126), .ZN(n9743) );
  AND2_X1 U13074 ( .A1(n10334), .A2(n10333), .ZN(n9744) );
  INV_X2 U13075 ( .A(n11667), .ZN(n11744) );
  OR2_X1 U13076 ( .A1(n18726), .A2(n18767), .ZN(n9745) );
  INV_X1 U13077 ( .A(n16331), .ZN(n10250) );
  INV_X1 U13078 ( .A(n15896), .ZN(n10234) );
  AND2_X1 U13079 ( .A1(n18055), .A2(n10269), .ZN(n9746) );
  OR2_X1 U13080 ( .A1(n19725), .A2(n19972), .ZN(n16550) );
  INV_X1 U13081 ( .A(n16550), .ZN(n19945) );
  AND2_X1 U13082 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9747) );
  OR2_X1 U13083 ( .A1(n13103), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10305) );
  INV_X1 U13084 ( .A(n10722), .ZN(n10477) );
  AND2_X1 U13085 ( .A1(n10305), .A2(n18663), .ZN(n9748) );
  OR2_X1 U13086 ( .A1(n18375), .A2(n10349), .ZN(n9749) );
  AND2_X1 U13087 ( .A1(n19829), .A2(n9624), .ZN(n9750) );
  INV_X1 U13088 ( .A(n16384), .ZN(n10384) );
  OR2_X1 U13089 ( .A1(n13775), .A2(n17112), .ZN(n20712) );
  INV_X1 U13090 ( .A(n20712), .ZN(n20887) );
  NAND2_X1 U13091 ( .A1(n12825), .A2(n12824), .ZN(n14046) );
  INV_X1 U13092 ( .A(n14046), .ZN(n10427) );
  AND2_X1 U13093 ( .A1(n10390), .A2(n10389), .ZN(n9751) );
  OR2_X1 U13094 ( .A1(n14045), .A2(n10429), .ZN(n10428) );
  AND2_X1 U13095 ( .A1(n9633), .A2(P3_EAX_REG_9__SCAN_IN), .ZN(n9752) );
  AND3_X2 U13096 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13625) );
  NAND2_X1 U13097 ( .A1(n11456), .A2(n11455), .ZN(n9753) );
  AND2_X1 U13098 ( .A1(n13485), .A2(n13484), .ZN(n9754) );
  INV_X1 U13099 ( .A(n10391), .ZN(n10390) );
  NAND2_X1 U13100 ( .A1(n9747), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10391) );
  AND2_X1 U13101 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n9755) );
  INV_X1 U13102 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n11759) );
  INV_X1 U13103 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10338) );
  INV_X1 U13104 ( .A(n17753), .ZN(n19555) );
  INV_X1 U13105 ( .A(n16016), .ZN(n10237) );
  NOR2_X1 U13106 ( .A1(n18686), .A2(n17738), .ZN(n17727) );
  INV_X1 U13107 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10345) );
  INV_X1 U13108 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10400) );
  AND2_X1 U13109 ( .A1(n12925), .A2(n12930), .ZN(n9756) );
  AND4_X1 U13110 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_22__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .A4(P3_EAX_REG_18__SCAN_IN), .ZN(n9757)
         );
  AND3_X1 U13111 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .ZN(n9758) );
  INV_X1 U13112 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19514) );
  AND2_X1 U13113 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .ZN(n9759) );
  INV_X1 U13114 ( .A(n10191), .ZN(n10190) );
  NAND2_X1 U13115 ( .A1(n10192), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n10191) );
  INV_X1 U13116 ( .A(n10264), .ZN(n10263) );
  NAND2_X1 U13117 ( .A1(n10266), .A2(n10265), .ZN(n10264) );
  AND2_X1 U13118 ( .A1(n10201), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n9760) );
  NAND2_X1 U13119 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12604) );
  NAND2_X1 U13120 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17738) );
  INV_X1 U13121 ( .A(n17738), .ZN(n10341) );
  INV_X1 U13122 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10233) );
  INV_X1 U13123 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n10209) );
  INV_X1 U13124 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n10194) );
  INV_X1 U13125 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n10202) );
  INV_X1 U13126 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n10203) );
  INV_X1 U13127 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10347) );
  INV_X1 U13128 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n9973) );
  INV_X1 U13129 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10337) );
  INV_X1 U13130 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10396) );
  AND2_X1 U13131 ( .A1(n11549), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9761) );
  AND2_X1 U13132 ( .A1(n10375), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9762) );
  INV_X1 U13133 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10399) );
  INV_X1 U13134 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n10211) );
  INV_X1 U13135 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10226) );
  AND2_X1 U13136 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n9763) );
  INV_X1 U13137 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n9972) );
  INV_X1 U13138 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10404) );
  INV_X1 U13139 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10376) );
  INV_X1 U13140 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n9891) );
  NAND2_X1 U13141 ( .A1(n10375), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10374) );
  OAI21_X1 U13142 ( .B1(n16693), .B2(n16483), .A(n9963), .ZN(P2_U3000) );
  OAI211_X1 U13143 ( .C1(n16586), .C2(n16483), .A(n9980), .B(n9979), .ZN(
        P2_U2988) );
  INV_X1 U13144 ( .A(n16483), .ZN(n10145) );
  OAI21_X1 U13145 ( .B1(n16634), .B2(n16483), .A(n10134), .ZN(n10133) );
  OR2_X1 U13146 ( .A1(n16761), .A2(n16483), .ZN(n9767) );
  AOI21_X1 U13147 ( .B1(n15043), .B2(n20758), .A(n10048), .ZN(n10047) );
  INV_X1 U13148 ( .A(n20758), .ZN(n20780) );
  OR2_X1 U13149 ( .A1(n20784), .A2(n11830), .ZN(n15026) );
  NAND2_X1 U13150 ( .A1(n19024), .A2(n19026), .ZN(n19027) );
  AOI22_X2 U13151 ( .A1(DATAI_22_), .A2(n13804), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n13844), .ZN(n21191) );
  NAND3_X1 U13152 ( .A1(n11165), .A2(n11155), .A3(n10786), .ZN(n11488) );
  NAND2_X2 U13153 ( .A1(n10787), .A2(n13585), .ZN(n10803) );
  NOR2_X1 U13154 ( .A1(n10808), .A2(n19984), .ZN(n9764) );
  NAND3_X1 U13155 ( .A1(n11540), .A2(n11541), .A3(n11537), .ZN(n10136) );
  NAND2_X1 U13156 ( .A1(n9766), .A2(n19945), .ZN(n16432) );
  OAI21_X1 U13157 ( .B1(n9768), .B2(n16757), .A(n9620), .ZN(P2_U3006) );
  OR2_X1 U13158 ( .A1(n16758), .A2(n16550), .ZN(n9768) );
  MUX2_X1 U13159 ( .A(n10977), .B(n10978), .S(n10212), .Z(n9769) );
  NAND4_X1 U13160 ( .A1(n10935), .A2(n10934), .A3(n10933), .A4(n10936), .ZN(
        n9770) );
  OAI21_X1 U13161 ( .B1(n16608), .B2(n16483), .A(n9772), .ZN(P2_U2990) );
  NAND3_X1 U13162 ( .A1(n9776), .A2(n9775), .A3(n9885), .ZN(n16608) );
  OR2_X1 U13163 ( .A1(n16362), .A2(n9888), .ZN(n9776) );
  NAND2_X2 U13164 ( .A1(n9784), .A2(n9783), .ZN(n10794) );
  AND4_X2 U13165 ( .A1(n9591), .A2(n9782), .A3(n10786), .A4(n10783), .ZN(
        n10103) );
  NAND2_X1 U13166 ( .A1(n10735), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9778) );
  NAND2_X4 U13167 ( .A1(n9781), .A2(n9780), .ZN(n10786) );
  INV_X1 U13168 ( .A(n10800), .ZN(n9782) );
  NAND2_X2 U13169 ( .A1(n10103), .A2(n10808), .ZN(n11180) );
  NAND2_X1 U13170 ( .A1(n10781), .A2(n10750), .ZN(n9784) );
  NAND2_X1 U13171 ( .A1(n16060), .A2(n16062), .ZN(n16061) );
  XNOR2_X1 U13172 ( .A(n14608), .B(n14628), .ZN(n16060) );
  INV_X1 U13173 ( .A(n13859), .ZN(n13862) );
  NAND2_X1 U13174 ( .A1(n9787), .A2(n13767), .ZN(n13860) );
  INV_X1 U13175 ( .A(n9787), .ZN(n9786) );
  NAND3_X1 U13176 ( .A1(n10813), .A2(n9863), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n9788) );
  NAND3_X1 U13177 ( .A1(n10806), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10805), 
        .ZN(n9789) );
  NAND2_X2 U13178 ( .A1(n10828), .A2(n9790), .ZN(n10821) );
  NAND3_X1 U13179 ( .A1(n9602), .A2(n10456), .A3(n9743), .ZN(n16119) );
  INV_X1 U13180 ( .A(n16119), .ZN(n14452) );
  NAND3_X1 U13181 ( .A1(n10061), .A2(n10842), .A3(n10860), .ZN(n10847) );
  OAI211_X2 U13182 ( .C1(n10833), .C2(n19964), .A(n10831), .B(n10832), .ZN(
        n10848) );
  NOR2_X2 U13183 ( .A1(n9797), .A2(n9796), .ZN(n20283) );
  INV_X1 U13184 ( .A(n10861), .ZN(n9797) );
  NOR2_X2 U13185 ( .A1(n9798), .A2(n9927), .ZN(n10921) );
  NAND2_X2 U13186 ( .A1(n9803), .A2(n16519), .ZN(n9969) );
  NAND2_X1 U13187 ( .A1(n10983), .A2(n10212), .ZN(n9803) );
  NAND2_X1 U13188 ( .A1(n11166), .A2(n10784), .ZN(n9805) );
  NAND4_X1 U13189 ( .A1(n10792), .A2(n13485), .A3(n13575), .A4(n11093), .ZN(
        n9804) );
  NAND2_X1 U13190 ( .A1(n12597), .A2(n10812), .ZN(n9806) );
  INV_X1 U13191 ( .A(n19976), .ZN(n9807) );
  INV_X1 U13192 ( .A(n9811), .ZN(n10043) );
  NAND2_X2 U13193 ( .A1(n9813), .A2(n9812), .ZN(n10834) );
  NAND4_X1 U13194 ( .A1(n10138), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10367), 
        .A4(n10792), .ZN(n9812) );
  NAND2_X1 U13195 ( .A1(n9679), .A2(n16818), .ZN(n9813) );
  AND2_X1 U13196 ( .A1(n10792), .A2(n10367), .ZN(n9917) );
  NAND3_X1 U13197 ( .A1(n11546), .A2(n11544), .A3(n9814), .ZN(n10369) );
  OAI211_X1 U13198 ( .C1(n11543), .C2(n10222), .A(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n9818), .ZN(n10997) );
  INV_X1 U13199 ( .A(n9582), .ZN(n9852) );
  NAND3_X1 U13200 ( .A1(n9654), .A2(n10131), .A3(n11549), .ZN(n16312) );
  NAND2_X1 U13201 ( .A1(n18382), .A2(n18634), .ZN(n9820) );
  NOR2_X1 U13202 ( .A1(n13151), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n18381) );
  AOI21_X2 U13203 ( .B1(n9822), .B2(n18427), .A(n9632), .ZN(n18408) );
  NAND3_X1 U13204 ( .A1(n9824), .A2(n10306), .A3(n10304), .ZN(n18650) );
  NAND3_X1 U13205 ( .A1(n9658), .A2(n10305), .A3(n18680), .ZN(n9824) );
  NAND2_X1 U13206 ( .A1(n18650), .A2(n18651), .ZN(n18649) );
  NAND2_X1 U13207 ( .A1(n9825), .A2(n18701), .ZN(n19023) );
  NAND2_X1 U13208 ( .A1(n18702), .A2(n9826), .ZN(n18701) );
  OR2_X1 U13209 ( .A1(n9826), .A2(n18702), .ZN(n9825) );
  OR2_X2 U13210 ( .A1(n13143), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18596) );
  NAND3_X1 U13211 ( .A1(n9949), .A2(n11534), .A3(n10182), .ZN(n9827) );
  NAND2_X1 U13212 ( .A1(n9829), .A2(n10846), .ZN(n10467) );
  NAND3_X1 U13213 ( .A1(n16529), .A2(n10530), .A3(n16528), .ZN(n10289) );
  NAND2_X2 U13214 ( .A1(n10146), .A2(n9830), .ZN(n16528) );
  NOR2_X1 U13215 ( .A1(n11292), .A2(n9832), .ZN(n11293) );
  NAND2_X1 U13216 ( .A1(n16287), .A2(n9832), .ZN(n16282) );
  XNOR2_X1 U13217 ( .A(n9833), .B(n14711), .ZN(n14739) );
  OR2_X2 U13218 ( .A1(n16426), .A2(n16425), .ZN(n10417) );
  NAND2_X1 U13219 ( .A1(n9950), .A2(n9951), .ZN(n9834) );
  NAND2_X1 U13220 ( .A1(n9835), .A2(n10920), .ZN(n10958) );
  NAND3_X2 U13221 ( .A1(n10904), .A2(n9723), .A3(n9835), .ZN(n11534) );
  NAND4_X2 U13222 ( .A1(n10916), .A2(n10917), .A3(n10915), .A4(n10918), .ZN(
        n9835) );
  INV_X1 U13223 ( .A(n11166), .ZN(n11169) );
  NOR2_X1 U13224 ( .A1(n10804), .A2(n9840), .ZN(n9839) );
  CLKBUF_X1 U13225 ( .A(n10812), .Z(n9861) );
  OAI21_X1 U13226 ( .B1(n16643), .B2(n19970), .A(n9705), .ZN(n9864) );
  INV_X1 U13227 ( .A(n9866), .ZN(n20347) );
  OAI21_X1 U13228 ( .B1(n9866), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n9865), .ZN(
        n20353) );
  OAI22_X1 U13229 ( .A1(n16890), .A2(n10870), .B1(n9866), .B2(n10871), .ZN(
        n10872) );
  OAI22_X1 U13230 ( .A1(n16890), .A2(n10930), .B1(n9866), .B2(n10929), .ZN(
        n10931) );
  OAI22_X1 U13231 ( .A1(n20143), .A2(n10906), .B1(n9866), .B2(n10905), .ZN(
        n10910) );
  OAI22_X1 U13232 ( .A1(n20143), .A2(n10945), .B1(n9866), .B2(n10944), .ZN(
        n10946) );
  NAND2_X1 U13233 ( .A1(n10417), .A2(n9711), .ZN(n9868) );
  NAND2_X1 U13234 ( .A1(n14708), .A2(n10299), .ZN(n10298) );
  NAND2_X1 U13235 ( .A1(n9869), .A2(n19861), .ZN(n9870) );
  NAND3_X1 U13236 ( .A1(n9969), .A2(n11543), .A3(n11542), .ZN(n9869) );
  XNOR2_X2 U13237 ( .A(n9870), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16514) );
  INV_X1 U13238 ( .A(n12719), .ZN(n9872) );
  INV_X1 U13239 ( .A(n17180), .ZN(n10165) );
  NAND3_X1 U13240 ( .A1(n9874), .A2(n9873), .A3(n20858), .ZN(n20857) );
  NAND2_X1 U13241 ( .A1(n10071), .A2(n12737), .ZN(n9873) );
  NAND2_X1 U13242 ( .A1(n10308), .A2(n12737), .ZN(n9874) );
  XNOR2_X1 U13243 ( .A(n12736), .B(n20908), .ZN(n20867) );
  NAND3_X1 U13244 ( .A1(n11917), .A2(n12960), .A3(n11882), .ZN(n9875) );
  NAND2_X2 U13245 ( .A1(n10281), .A2(n10279), .ZN(n15237) );
  NAND4_X1 U13246 ( .A1(n10175), .A2(n10173), .A3(n20887), .A4(n10177), .ZN(
        n9877) );
  INV_X1 U13247 ( .A(n9880), .ZN(n9878) );
  INV_X1 U13248 ( .A(n9881), .ZN(n9879) );
  AND2_X1 U13249 ( .A1(n16607), .A2(n19967), .ZN(n9890) );
  NAND2_X1 U13250 ( .A1(n9894), .A2(n9892), .ZN(n9898) );
  INV_X1 U13251 ( .A(n9900), .ZN(n9895) );
  OAI21_X1 U13252 ( .B1(n12522), .B2(n12524), .A(n12521), .ZN(n9902) );
  OR2_X2 U13253 ( .A1(n17107), .A2(n20710), .ZN(n13775) );
  NAND3_X1 U13254 ( .A1(n9908), .A2(n13023), .A3(n13022), .ZN(n13024) );
  MUX2_X1 U13255 ( .A(n16516), .B(n16517), .S(n10104), .Z(n16518) );
  NAND2_X1 U13256 ( .A1(n9917), .A2(n10138), .ZN(n10822) );
  XNOR2_X1 U13257 ( .A(n10860), .B(n9918), .ZN(n13606) );
  NAND2_X1 U13258 ( .A1(n13581), .A2(n9918), .ZN(n10856) );
  NAND3_X1 U13259 ( .A1(n9949), .A2(n9920), .A3(n11534), .ZN(n9919) );
  NAND3_X1 U13260 ( .A1(n9949), .A2(n11534), .A3(n11542), .ZN(n9923) );
  NAND2_X2 U13261 ( .A1(n9924), .A2(n9926), .ZN(n16327) );
  NAND3_X1 U13262 ( .A1(n10150), .A2(n9704), .A3(n10151), .ZN(n9924) );
  NAND3_X1 U13263 ( .A1(n10150), .A2(n10151), .A3(n10148), .ZN(n9925) );
  OAI211_X1 U13264 ( .C1(n9931), .C2(n16327), .A(n19958), .B(n9929), .ZN(
        n16576) );
  NAND3_X1 U13265 ( .A1(n16327), .A2(n9932), .A3(n9930), .ZN(n9929) );
  OR2_X1 U13266 ( .A1(n10011), .A2(n9935), .ZN(n9933) );
  NAND3_X1 U13267 ( .A1(n9939), .A2(n17743), .A3(n9938), .ZN(n9937) );
  NOR2_X2 U13268 ( .A1(n13355), .A2(n19074), .ZN(n19500) );
  NAND2_X2 U13269 ( .A1(n19485), .A2(n9941), .ZN(n19499) );
  NAND2_X1 U13270 ( .A1(n19513), .A2(n19663), .ZN(n9947) );
  NAND2_X1 U13271 ( .A1(n9949), .A2(n11534), .ZN(n16539) );
  INV_X1 U13272 ( .A(n10815), .ZN(n9951) );
  INV_X1 U13273 ( .A(n10066), .ZN(n9961) );
  XNOR2_X2 U13274 ( .A(n10983), .B(n9962), .ZN(n10066) );
  AOI21_X1 U13275 ( .B1(n10821), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10839), .ZN(n11181) );
  AOI21_X1 U13276 ( .B1(n14749), .B2(n16799), .A(n11521), .ZN(n10360) );
  MUX2_X1 U13277 ( .A(n10980), .B(n10981), .S(n10212), .Z(n10147) );
  NAND2_X1 U13278 ( .A1(n10007), .A2(n10292), .ZN(n16449) );
  NAND4_X1 U13279 ( .A1(n10171), .A2(n10169), .A3(n9984), .A4(n9983), .ZN(
        n11845) );
  NAND2_X2 U13280 ( .A1(n11710), .A2(n11719), .ZN(n11722) );
  NAND3_X1 U13281 ( .A1(n10164), .A2(n10162), .A3(n10317), .ZN(n17165) );
  NAND2_X1 U13282 ( .A1(n10445), .A2(n9990), .ZN(n9989) );
  NAND2_X1 U13283 ( .A1(n15237), .A2(n10003), .ZN(n10002) );
  AOI21_X1 U13284 ( .B1(n10014), .B2(n10007), .A(n10013), .ZN(n16426) );
  INV_X1 U13285 ( .A(n10008), .ZN(n16385) );
  AND2_X4 U13286 ( .A1(n10131), .A2(n10369), .ZN(n14360) );
  NAND2_X1 U13287 ( .A1(n10009), .A2(n10024), .ZN(n10021) );
  NAND2_X1 U13288 ( .A1(n10009), .A2(n9700), .ZN(n10031) );
  OAI21_X1 U13289 ( .B1(n10009), .B2(n10026), .A(n10022), .ZN(n14299) );
  NAND2_X1 U13290 ( .A1(n16449), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10012) );
  NAND2_X2 U13291 ( .A1(n10584), .A2(n10585), .ZN(n10784) );
  NAND2_X1 U13292 ( .A1(n10902), .A2(n10793), .ZN(n10603) );
  NOR2_X2 U13293 ( .A1(n10955), .A2(n10956), .ZN(n10990) );
  OR2_X2 U13294 ( .A1(n11022), .A2(n10018), .ZN(n11021) );
  NAND2_X1 U13295 ( .A1(n18719), .A2(n18711), .ZN(n10302) );
  XNOR2_X1 U13296 ( .A(n18247), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18711) );
  NAND2_X1 U13297 ( .A1(n18688), .A2(n18689), .ZN(n18687) );
  NAND2_X1 U13298 ( .A1(n13359), .A2(n18960), .ZN(n13377) );
  NAND2_X1 U13299 ( .A1(n10224), .A2(n18427), .ZN(n10039) );
  NOR2_X2 U13300 ( .A1(n18393), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n18392) );
  NAND2_X1 U13301 ( .A1(n18633), .A2(n10042), .ZN(n18518) );
  NAND2_X1 U13302 ( .A1(n10040), .A2(n10041), .ZN(n18513) );
  NAND3_X1 U13303 ( .A1(n9657), .A2(n18633), .A3(n10042), .ZN(n10040) );
  NAND3_X1 U13304 ( .A1(n12951), .A2(n21276), .A3(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n10050) );
  OAI21_X2 U13305 ( .B1(n12557), .B2(n12556), .A(n12560), .ZN(n17107) );
  NAND3_X1 U13306 ( .A1(n11106), .A2(n11107), .A3(n10055), .ZN(n11115) );
  OAI211_X1 U13307 ( .C1(n11105), .C2(n11280), .A(n12597), .B(n11104), .ZN(
        n10055) );
  NAND2_X1 U13308 ( .A1(n10064), .A2(n10062), .ZN(n10842) );
  AOI21_X1 U13309 ( .B1(n10834), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n10063), .ZN(n10062) );
  AOI21_X2 U13310 ( .B1(n10821), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n10065), .ZN(n10064) );
  INV_X1 U13311 ( .A(n11757), .ZN(n10069) );
  NAND2_X1 U13312 ( .A1(n12786), .A2(n10070), .ZN(n12787) );
  NAND2_X1 U13313 ( .A1(n18656), .A2(n9755), .ZN(n10075) );
  NOR2_X1 U13314 ( .A1(n10074), .A2(n9682), .ZN(n10073) );
  NAND2_X1 U13315 ( .A1(n13319), .A2(n10082), .ZN(n10081) );
  INV_X1 U13316 ( .A(n11880), .ZN(n14005) );
  NAND2_X2 U13317 ( .A1(n10083), .A2(n11880), .ZN(n11917) );
  AOI21_X2 U13318 ( .B1(n12713), .B2(n11836), .A(n11824), .ZN(n11825) );
  XNOR2_X2 U13319 ( .A(n11755), .B(n11754), .ZN(n11826) );
  NOR2_X1 U13320 ( .A1(n17789), .A2(n13044), .ZN(n13054) );
  AND2_X2 U13321 ( .A1(n10086), .A2(n11553), .ZN(n11761) );
  AND2_X2 U13322 ( .A1(n10086), .A2(n11563), .ZN(n12218) );
  AND2_X2 U13323 ( .A1(n10086), .A2(n11565), .ZN(n11745) );
  AND2_X2 U13324 ( .A1(n10086), .A2(n11552), .ZN(n11731) );
  NAND4_X1 U13325 ( .A1(n10094), .A2(n14172), .A3(n10095), .A4(n10096), .ZN(
        n14171) );
  AND2_X1 U13326 ( .A1(n14861), .A2(n9662), .ZN(n14815) );
  INV_X1 U13327 ( .A(n12804), .ZN(n12976) );
  NAND2_X1 U13328 ( .A1(n9699), .A2(n12804), .ZN(n10100) );
  AND2_X2 U13329 ( .A1(n11695), .A2(n13845), .ZN(n12804) );
  INV_X4 U13330 ( .A(n11752), .ZN(n13845) );
  NAND2_X1 U13331 ( .A1(n12781), .A2(n9710), .ZN(n10101) );
  NAND4_X1 U13332 ( .A1(n11880), .A2(n11825), .A3(n11826), .A4(n9702), .ZN(
        n11960) );
  NAND4_X1 U13333 ( .A1(n10371), .A2(n10130), .A3(n11539), .A4(n10370), .ZN(
        n16494) );
  INV_X1 U13334 ( .A(n10842), .ZN(n10107) );
  NAND2_X1 U13335 ( .A1(n10473), .A2(n10470), .ZN(n10723) );
  AOI21_X2 U13336 ( .B1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n10921), .A(
        n10880), .ZN(n10884) );
  NAND4_X2 U13337 ( .A1(n10884), .A2(n10885), .A3(n10886), .A4(n10883), .ZN(
        n10904) );
  NAND2_X1 U13338 ( .A1(n12738), .A2(n12960), .ZN(n10159) );
  NAND2_X1 U13339 ( .A1(n10282), .A2(n15385), .ZN(n10281) );
  INV_X1 U13340 ( .A(n15658), .ZN(n10321) );
  NAND3_X1 U13341 ( .A1(n12782), .A2(n15197), .A3(n15374), .ZN(n15189) );
  NAND2_X1 U13342 ( .A1(n10112), .A2(n10276), .ZN(n10275) );
  NAND2_X1 U13343 ( .A1(n10174), .A2(n9740), .ZN(n10274) );
  NAND3_X1 U13344 ( .A1(n13025), .A2(n12566), .A3(n10113), .ZN(n11702) );
  OAI21_X1 U13345 ( .B1(n10117), .B2(n21470), .A(n10316), .ZN(n10113) );
  AND4_X2 U13346 ( .A1(n10115), .A2(n10116), .A3(n11707), .A4(n11628), .ZN(
        n10316) );
  NAND2_X1 U13347 ( .A1(n10316), .A2(n21470), .ZN(n10314) );
  NOR2_X1 U13348 ( .A1(n11698), .A2(n12977), .ZN(n11659) );
  INV_X1 U13349 ( .A(n12977), .ZN(n10115) );
  INV_X1 U13350 ( .A(n11698), .ZN(n10116) );
  AOI21_X1 U13351 ( .B1(n11184), .B2(n10129), .A(n11183), .ZN(n14099) );
  XNOR2_X2 U13352 ( .A(n10129), .B(n10841), .ZN(n13875) );
  OR2_X1 U13353 ( .A1(n18247), .A2(n13072), .ZN(n13073) );
  OR2_X2 U13354 ( .A1(n17288), .A2(n18222), .ZN(n10142) );
  NAND3_X1 U13355 ( .A1(n10352), .A2(n10351), .A3(n10145), .ZN(n10144) );
  INV_X1 U13356 ( .A(n10287), .ZN(n10149) );
  AND2_X1 U13357 ( .A1(n9611), .A2(n9714), .ZN(n10148) );
  NAND3_X1 U13358 ( .A1(n10151), .A2(n10150), .A3(n9611), .ZN(n16347) );
  XNOR2_X2 U13359 ( .A(n11917), .B(n11918), .ZN(n12738) );
  INV_X1 U13360 ( .A(n10161), .ZN(n11705) );
  NAND2_X1 U13361 ( .A1(n11722), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10166) );
  INV_X1 U13362 ( .A(n11718), .ZN(n10171) );
  NAND3_X1 U13363 ( .A1(n10173), .A2(n10172), .A3(n10177), .ZN(n13031) );
  AND2_X1 U13364 ( .A1(n10175), .A2(n20922), .ZN(n10172) );
  NAND3_X1 U13365 ( .A1(n10174), .A2(n12787), .A3(n13019), .ZN(n10173) );
  NAND2_X1 U13366 ( .A1(n18188), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n18184) );
  NAND3_X1 U13367 ( .A1(n13256), .A2(n13251), .A3(n13257), .ZN(n10197) );
  NAND3_X1 U13368 ( .A1(n13255), .A2(n10200), .A3(n13254), .ZN(n10199) );
  NAND2_X1 U13369 ( .A1(n18141), .A2(n9760), .ZN(n18128) );
  NAND3_X1 U13370 ( .A1(n13284), .A2(n13275), .A3(n10206), .ZN(n10205) );
  INV_X1 U13371 ( .A(n18250), .ZN(n10207) );
  NAND2_X1 U13372 ( .A1(n10207), .A2(n10208), .ZN(n18189) );
  OR2_X2 U13373 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13042) );
  INV_X1 U13374 ( .A(n10214), .ZN(n10213) );
  OAI21_X1 U13375 ( .B1(n16483), .B2(n14387), .A(n14386), .ZN(P2_U2995) );
  OAI21_X1 U13376 ( .B1(n18639), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n10223), .ZN(n18974) );
  INV_X1 U13377 ( .A(n10225), .ZN(n10224) );
  NAND2_X1 U13378 ( .A1(n18427), .A2(n18465), .ZN(n18504) );
  NAND3_X1 U13379 ( .A1(n13144), .A2(n21454), .A3(n10233), .ZN(n10232) );
  MUX2_X1 U13380 ( .A(n19964), .B(n12625), .S(n20690), .Z(n16823) );
  OR2_X1 U13381 ( .A1(n15857), .A2(n10245), .ZN(n10243) );
  NAND2_X1 U13382 ( .A1(n10243), .A2(n10244), .ZN(n15802) );
  INV_X1 U13383 ( .A(n13875), .ZN(n10875) );
  NAND3_X1 U13384 ( .A1(n10254), .A2(n10253), .A3(n10251), .ZN(P2_U3034) );
  OR2_X1 U13385 ( .A1(n16711), .A2(n19970), .ZN(n10253) );
  OR2_X1 U13386 ( .A1(n16715), .A2(n16802), .ZN(n10254) );
  NAND3_X1 U13387 ( .A1(n16966), .A2(n19084), .A3(n19070), .ZN(n10259) );
  INV_X2 U13388 ( .A(n13266), .ZN(n19062) );
  NAND3_X1 U13389 ( .A1(n13239), .A2(n13240), .A3(n10261), .ZN(n10260) );
  NAND3_X1 U13390 ( .A1(n10271), .A2(n11730), .A3(n11759), .ZN(n10438) );
  INV_X1 U13391 ( .A(n10271), .ZN(n10270) );
  NAND2_X1 U13392 ( .A1(n10271), .A2(n11730), .ZN(n13618) );
  XNOR2_X1 U13393 ( .A(n10271), .B(n13883), .ZN(n13938) );
  NAND2_X2 U13394 ( .A1(n11726), .A2(n11725), .ZN(n10271) );
  NAND4_X1 U13395 ( .A1(n15330), .A2(n12698), .A3(n9669), .A4(n12699), .ZN(
        n15296) );
  NOR2_X1 U13396 ( .A1(n10272), .A2(n15331), .ZN(n15320) );
  NAND2_X1 U13397 ( .A1(n12698), .A2(n9669), .ZN(n10272) );
  NAND2_X1 U13398 ( .A1(n15296), .A2(n15283), .ZN(n12702) );
  NAND2_X1 U13399 ( .A1(n12698), .A2(n15321), .ZN(n15334) );
  NAND2_X1 U13400 ( .A1(n10273), .A2(n10278), .ZN(P1_U3002) );
  NAND3_X1 U13401 ( .A1(n10275), .A2(n10274), .A3(n20922), .ZN(n10273) );
  INV_X1 U13402 ( .A(n10280), .ZN(n10279) );
  OAI21_X1 U13403 ( .B1(n15284), .B2(n10284), .A(n9707), .ZN(n10280) );
  NOR2_X1 U13404 ( .A1(n15284), .A2(n10283), .ZN(n10282) );
  AOI21_X1 U13405 ( .B1(n16529), .B2(n16528), .A(n10293), .ZN(n16515) );
  NOR2_X1 U13406 ( .A1(n16514), .A2(n16515), .ZN(n16457) );
  AND2_X1 U13407 ( .A1(n14708), .A2(n16418), .ZN(n16408) );
  OAI21_X1 U13408 ( .B1(n18711), .B2(n18719), .A(n10302), .ZN(n19036) );
  OR2_X1 U13409 ( .A1(n18680), .A2(n18681), .ZN(n10307) );
  NAND3_X1 U13410 ( .A1(n9658), .A2(n10305), .A3(n18681), .ZN(n10304) );
  INV_X1 U13411 ( .A(n10307), .ZN(n18679) );
  NAND2_X2 U13412 ( .A1(n18962), .A2(n18634), .ZN(n18633) );
  INV_X1 U13413 ( .A(n20866), .ZN(n10308) );
  NAND2_X1 U13414 ( .A1(n20873), .A2(n12735), .ZN(n20866) );
  NAND2_X1 U13415 ( .A1(n20865), .A2(n12737), .ZN(n20859) );
  NOR2_X4 U13416 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15666) );
  OAI211_X2 U13417 ( .C1(n11722), .C2(n10312), .A(n10310), .B(n10309), .ZN(
        n14010) );
  NAND2_X1 U13418 ( .A1(n11722), .A2(n9674), .ZN(n10309) );
  OAI21_X1 U13419 ( .B1(n11719), .B2(n9709), .A(n10311), .ZN(n10310) );
  NAND2_X1 U13420 ( .A1(n11719), .A2(n11712), .ZN(n10311) );
  NAND2_X1 U13421 ( .A1(n10313), .A2(n11712), .ZN(n10312) );
  INV_X1 U13422 ( .A(n11719), .ZN(n10313) );
  NAND3_X1 U13423 ( .A1(n12788), .A2(n11659), .A3(n9581), .ZN(n17099) );
  NAND2_X1 U13424 ( .A1(n17178), .A2(n10318), .ZN(n17174) );
  NAND2_X1 U13425 ( .A1(n10321), .A2(n12107), .ZN(n11888) );
  OR2_X1 U13426 ( .A1(n17477), .A2(n17653), .ZN(n10328) );
  AOI21_X1 U13427 ( .B1(n17477), .B2(n10327), .A(n17653), .ZN(n17457) );
  NAND2_X1 U13428 ( .A1(n17477), .A2(n10326), .ZN(n10325) );
  INV_X1 U13429 ( .A(n10328), .ZN(n17469) );
  INV_X1 U13430 ( .A(n18362), .ZN(n10327) );
  AOI21_X1 U13431 ( .B1(n17550), .B2(n10333), .A(n17653), .ZN(n17531) );
  NAND2_X1 U13432 ( .A1(n10331), .A2(n10329), .ZN(n17530) );
  NAND2_X1 U13433 ( .A1(n17550), .A2(n10332), .ZN(n10331) );
  INV_X1 U13434 ( .A(n10334), .ZN(n17541) );
  NAND3_X1 U13435 ( .A1(n10339), .A2(n10340), .A3(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18626) );
  NAND3_X1 U13436 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n10341), .A3(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17714) );
  NAND2_X1 U13437 ( .A1(n10343), .A2(n9618), .ZN(n17432) );
  NAND2_X1 U13438 ( .A1(n10350), .A2(n10360), .ZN(P2_U3015) );
  NAND3_X1 U13439 ( .A1(n10351), .A2(n10356), .A3(n9689), .ZN(n10350) );
  OR2_X1 U13440 ( .A1(n11102), .A2(n10362), .ZN(n10357) );
  NAND2_X1 U13441 ( .A1(n14300), .A2(n16293), .ZN(n10362) );
  NAND2_X1 U13442 ( .A1(n11551), .A2(n10365), .ZN(n16782) );
  NAND2_X1 U13443 ( .A1(n10797), .A2(n10366), .ZN(n10368) );
  NAND2_X2 U13444 ( .A1(n10790), .A2(n12672), .ZN(n20689) );
  OAI21_X1 U13445 ( .B1(n10803), .B2(n10788), .A(n10368), .ZN(n10367) );
  NAND2_X1 U13446 ( .A1(n10371), .A2(n11539), .ZN(n16521) );
  NAND2_X1 U13447 ( .A1(n10377), .A2(n19866), .ZN(n15857) );
  NAND3_X1 U13448 ( .A1(n10383), .A2(n10380), .A3(n10379), .ZN(n10377) );
  NAND3_X1 U13449 ( .A1(n10388), .A2(n10387), .A3(n10386), .ZN(n14742) );
  OAI21_X1 U13450 ( .B1(n10415), .B2(n20545), .A(n10411), .ZN(P2_U2826) );
  XNOR2_X1 U13451 ( .A(n15783), .B(n10537), .ZN(n10415) );
  NOR2_X1 U13452 ( .A1(n14773), .A2(n10419), .ZN(n14762) );
  NAND2_X1 U13453 ( .A1(n14919), .A2(n9742), .ZN(n14892) );
  NAND2_X1 U13454 ( .A1(n10438), .A2(n9708), .ZN(n11755) );
  NOR2_X1 U13455 ( .A1(n14784), .A2(n10449), .ZN(n14760) );
  NOR2_X1 U13456 ( .A1(n14784), .A2(n14785), .ZN(n14770) );
  NAND2_X1 U13457 ( .A1(n14056), .A2(n14055), .ZN(n10456) );
  AND2_X4 U13458 ( .A1(n11137), .A2(n16821), .ZN(n14516) );
  AND2_X2 U13459 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11137) );
  INV_X1 U13460 ( .A(n16055), .ZN(n10460) );
  NAND2_X1 U13461 ( .A1(n10467), .A2(n13580), .ZN(n10464) );
  NAND2_X1 U13462 ( .A1(n10845), .A2(n10844), .ZN(n10468) );
  INV_X1 U13463 ( .A(n13765), .ZN(n10465) );
  NAND3_X1 U13464 ( .A1(n10804), .A2(n10803), .A3(n13485), .ZN(n10805) );
  OR2_X2 U13465 ( .A1(n10469), .A2(n11092), .ZN(n11098) );
  XNOR2_X1 U13466 ( .A(n10469), .B(n11092), .ZN(n15782) );
  NAND2_X1 U13467 ( .A1(n11091), .A2(n11090), .ZN(n10469) );
  NAND2_X1 U13468 ( .A1(n11029), .A2(n9741), .ZN(n11022) );
  AND2_X1 U13469 ( .A1(n11039), .A2(n10478), .ZN(n15827) );
  NAND2_X1 U13470 ( .A1(n11039), .A2(n10475), .ZN(n11079) );
  NAND2_X1 U13471 ( .A1(n11039), .A2(n10722), .ZN(n11043) );
  NAND2_X1 U13472 ( .A1(n10984), .A2(n10480), .ZN(n10998) );
  INV_X1 U13473 ( .A(n10998), .ZN(n10717) );
  NAND2_X1 U13474 ( .A1(n14366), .A2(n14400), .ZN(n14399) );
  NOR2_X2 U13475 ( .A1(n16112), .A2(n14365), .ZN(n14366) );
  NAND2_X1 U13476 ( .A1(n14718), .A2(n11233), .ZN(n16112) );
  NOR2_X2 U13477 ( .A1(n14717), .A2(n14721), .ZN(n14718) );
  NOR2_X2 U13478 ( .A1(n16130), .A2(n10481), .ZN(n14254) );
  NAND2_X1 U13479 ( .A1(n11198), .A2(n9619), .ZN(n16142) );
  NAND2_X1 U13480 ( .A1(n15800), .A2(n15801), .ZN(n14326) );
  AND2_X2 U13481 ( .A1(n15800), .A2(n10488), .ZN(n15774) );
  AND2_X4 U13482 ( .A1(n10560), .A2(n16821), .ZN(n14513) );
  NOR2_X1 U13483 ( .A1(n11138), .A2(n10560), .ZN(n16841) );
  INV_X1 U13484 ( .A(n10803), .ZN(n11292) );
  NAND2_X1 U13485 ( .A1(n15854), .A2(n10491), .ZN(n15813) );
  NAND2_X2 U13486 ( .A1(n10787), .A2(n11286), .ZN(n11443) );
  MUX2_X1 U13487 ( .A(n10630), .B(n11524), .S(n10787), .Z(n10966) );
  NAND2_X1 U13488 ( .A1(n15963), .A2(n10495), .ZN(n10494) );
  NAND2_X1 U13489 ( .A1(n10494), .A2(n10498), .ZN(n13593) );
  AND2_X1 U13490 ( .A1(n11318), .A2(n10501), .ZN(n10500) );
  NAND2_X1 U13491 ( .A1(n10904), .A2(n10903), .ZN(n10957) );
  NOR2_X1 U13492 ( .A1(n16312), .A2(n10527), .ZN(n16298) );
  NAND2_X1 U13493 ( .A1(n10526), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10525) );
  INV_X1 U13494 ( .A(n10527), .ZN(n10526) );
  INV_X1 U13495 ( .A(n14402), .ZN(n11457) );
  OAI211_X1 U13496 ( .C1(n14697), .C2(n17237), .A(n14308), .B(n10531), .ZN(
        n14309) );
  NAND2_X1 U13497 ( .A1(n11457), .A2(n9753), .ZN(n15871) );
  CLKBUF_X1 U13498 ( .A(n14513), .Z(n14680) );
  INV_X1 U13499 ( .A(n12777), .ZN(n15374) );
  OR2_X1 U13500 ( .A1(n12777), .A2(n15511), .ZN(n15321) );
  AND2_X2 U13501 ( .A1(n14516), .A2(n10750), .ZN(n10888) );
  INV_X1 U13502 ( .A(n13860), .ZN(n13861) );
  NAND2_X1 U13503 ( .A1(n12955), .A2(n12579), .ZN(n12595) );
  AND2_X1 U13504 ( .A1(n16378), .A2(n14391), .ZN(n14395) );
  INV_X1 U13505 ( .A(n14056), .ZN(n13871) );
  AOI21_X1 U13506 ( .B1(n14426), .B2(n16799), .A(n14311), .ZN(n14312) );
  AND2_X1 U13507 ( .A1(n10875), .A2(n10876), .ZN(n16903) );
  AND2_X1 U13508 ( .A1(n10875), .A2(n10859), .ZN(n20465) );
  AND2_X1 U13509 ( .A1(n10875), .A2(n10858), .ZN(n20315) );
  OR2_X1 U13510 ( .A1(n13875), .A2(n16963), .ZN(n13867) );
  AND2_X1 U13511 ( .A1(n13875), .A2(n10874), .ZN(n20008) );
  CLKBUF_X3 U13512 ( .A(n10686), .Z(n14529) );
  AND2_X1 U13513 ( .A1(n10800), .A2(n10786), .ZN(n10529) );
  AND2_X1 U13514 ( .A1(n11005), .A2(n11004), .ZN(n10530) );
  NAND2_X1 U13515 ( .A1(n12578), .A2(n9905), .ZN(n15154) );
  INV_X2 U13516 ( .A(n15154), .ZN(n15150) );
  OR2_X1 U13517 ( .A1(n14307), .A2(n14306), .ZN(n10531) );
  OR3_X1 U13518 ( .A1(n14306), .A2(n11511), .A3(n11510), .ZN(n10532) );
  OR3_X1 U13519 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n18452), .ZN(n10533) );
  OR2_X1 U13520 ( .A1(n18408), .A2(n10142), .ZN(n10534) );
  NAND2_X1 U13521 ( .A1(n18634), .A2(n18730), .ZN(n10535) );
  INV_X1 U13522 ( .A(n11907), .ZN(n12503) );
  INV_X1 U13523 ( .A(n12503), .ZN(n12273) );
  OR2_X1 U13524 ( .A1(n10142), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10536) );
  NOR2_X1 U13525 ( .A1(n12658), .A2(n12659), .ZN(n10537) );
  AND3_X1 U13526 ( .A1(n13047), .A2(n13046), .A3(n13045), .ZN(n10538) );
  OR2_X1 U13527 ( .A1(n16074), .A2(n16066), .ZN(n10539) );
  AND4_X1 U13528 ( .A1(n11737), .A2(n11736), .A3(n11735), .A4(n11734), .ZN(
        n10540) );
  OR2_X1 U13529 ( .A1(n15409), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10541) );
  AND4_X1 U13530 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(P3_EAX_REG_1__SCAN_IN), .A4(P3_EAX_REG_0__SCAN_IN), .ZN(n10542) );
  INV_X1 U13531 ( .A(n16104), .ZN(n16154) );
  OR2_X1 U13532 ( .A1(n13281), .A2(n13266), .ZN(n10543) );
  AND4_X1 U13533 ( .A1(n13037), .A2(n13036), .A3(n13035), .A4(n13034), .ZN(
        n10544) );
  AND3_X1 U13534 ( .A1(n19819), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n11096), .ZN(n10545) );
  NOR2_X1 U13535 ( .A1(n16298), .A2(n16297), .ZN(n10546) );
  NAND2_X1 U13536 ( .A1(n13813), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12172) );
  INV_X1 U13537 ( .A(n12172), .ZN(n12107) );
  NOR2_X1 U13538 ( .A1(n21053), .A2(n21135), .ZN(n10548) );
  INV_X1 U13539 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12013) );
  INV_X1 U13540 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12602) );
  AND4_X1 U13541 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_5__SCAN_IN), .A4(P3_EAX_REG_4__SCAN_IN), .ZN(n10549) );
  INV_X1 U13542 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13330) );
  INV_X1 U13543 ( .A(n18177), .ZN(n18194) );
  NAND2_X2 U13544 ( .A1(n10207), .A2(n18213), .ZN(n18177) );
  NOR2_X1 U13545 ( .A1(n13041), .A2(n13033), .ZN(n17816) );
  INV_X1 U13546 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16921) );
  AND2_X1 U13547 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10550) );
  NAND2_X1 U13548 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATEBS16_REG_SCAN_IN), .ZN(n10551) );
  INV_X1 U13549 ( .A(n15868), .ZN(n15884) );
  NOR2_X1 U13550 ( .A1(n20309), .A2(n20114), .ZN(n10553) );
  INV_X1 U13551 ( .A(n14726), .ZN(n16240) );
  INV_X1 U13552 ( .A(n11733), .ZN(n12490) );
  INV_X1 U13553 ( .A(n11803), .ZN(n12447) );
  NAND2_X1 U13554 ( .A1(n9635), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10877) );
  INV_X1 U13555 ( .A(n12403), .ZN(n12479) );
  OR2_X1 U13556 ( .A1(n10926), .A2(n10863), .ZN(n10864) );
  AOI22_X1 U13557 ( .A1(n14514), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14513), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10612) );
  OR2_X1 U13558 ( .A1(n12383), .A2(n12382), .ZN(n12413) );
  INV_X1 U13559 ( .A(n11760), .ZN(n12460) );
  OR2_X1 U13560 ( .A1(n11901), .A2(n11900), .ZN(n12741) );
  INV_X1 U13561 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10721) );
  AND4_X1 U13562 ( .A1(n10941), .A2(n10940), .A3(n10939), .A4(n10938), .ZN(
        n10949) );
  NAND2_X1 U13563 ( .A1(n19984), .A2(n10786), .ZN(n10809) );
  INV_X1 U13564 ( .A(n12517), .ZN(n12525) );
  INV_X1 U13565 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12491) );
  NAND2_X1 U13566 ( .A1(n11745), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11664) );
  AND2_X1 U13567 ( .A1(n13563), .A2(n11695), .ZN(n12960) );
  OR2_X1 U13568 ( .A1(n11767), .A2(n11633), .ZN(n11636) );
  NAND2_X1 U13569 ( .A1(n11076), .A2(n11021), .ZN(n11016) );
  NAND2_X1 U13570 ( .A1(n11093), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10649) );
  NAND2_X1 U13571 ( .A1(n10646), .A2(n10645), .ZN(n10670) );
  NOR2_X1 U13572 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14507) );
  INV_X1 U13573 ( .A(n20661), .ZN(n11288) );
  INV_X1 U13574 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15010) );
  INV_X1 U13575 ( .A(n12274), .ZN(n12275) );
  NOR2_X1 U13576 ( .A1(n13758), .A2(n11830), .ZN(n11935) );
  OR2_X1 U13577 ( .A1(n12120), .A2(n11759), .ZN(n12471) );
  AND2_X1 U13578 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12036) );
  NAND2_X1 U13579 ( .A1(n12672), .A2(n11108), .ZN(n10647) );
  INV_X1 U13580 ( .A(n11023), .ZN(n10720) );
  AND2_X1 U13581 ( .A1(n11109), .A2(n11108), .ZN(n11143) );
  INV_X1 U13582 ( .A(n16143), .ZN(n11208) );
  INV_X1 U13583 ( .A(n11181), .ZN(n10840) );
  NOR2_X1 U13584 ( .A1(n16081), .A2(n16080), .ZN(n14570) );
  INV_X1 U13585 ( .A(n13935), .ZN(n11416) );
  INV_X1 U13586 ( .A(n14719), .ZN(n14720) );
  NAND2_X1 U13587 ( .A1(n10997), .A2(n10996), .ZN(n11006) );
  AOI22_X1 U13588 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n19514), .B2(n19663), .ZN(
        n13167) );
  INV_X1 U13589 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17829) );
  NAND2_X1 U13590 ( .A1(n17961), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n13045) );
  NAND2_X1 U13591 ( .A1(n16966), .A2(n13274), .ZN(n13268) );
  NAND2_X1 U13592 ( .A1(n12554), .A2(n12553), .ZN(n12572) );
  OR2_X1 U13593 ( .A1(n12790), .A2(n15168), .ZN(n12792) );
  AND2_X1 U13594 ( .A1(n12855), .A2(n12854), .ZN(n14281) );
  INV_X1 U13595 ( .A(n11966), .ZN(n11967) );
  NAND2_X1 U13596 ( .A1(n12443), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12790) );
  INV_X1 U13597 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14907) );
  NAND2_X1 U13598 ( .A1(n12094), .A2(n12093), .ZN(n12156) );
  AND2_X1 U13599 ( .A1(n12107), .A2(n12053), .ZN(n14953) );
  AND2_X1 U13600 ( .A1(n12894), .A2(n12893), .ZN(n14817) );
  OAI211_X1 U13601 ( .C1(n15766), .C2(n21064), .A(n21098), .B(n15736), .ZN(
        n15765) );
  INV_X1 U13602 ( .A(n11836), .ZN(n11837) );
  AND4_X1 U13603 ( .A1(n11582), .A2(n11581), .A3(n11580), .A4(n11579), .ZN(
        n11605) );
  INV_X1 U13604 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n17089) );
  NAND2_X1 U13605 ( .A1(n10583), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10584) );
  INV_X1 U13606 ( .A(n15869), .ZN(n11246) );
  INV_X1 U13607 ( .A(n14107), .ZN(n11197) );
  OR2_X1 U13608 ( .A1(n15781), .A2(n12681), .ZN(n12682) );
  OAI211_X1 U13609 ( .C1(n14627), .C2(n14626), .A(n14625), .B(n14660), .ZN(
        n14628) );
  OAI21_X1 U13610 ( .B1(n14316), .B2(n15804), .A(n16334), .ZN(n14317) );
  INV_X1 U13611 ( .A(n11548), .ZN(n11549) );
  NOR2_X1 U13612 ( .A1(n10545), .A2(n11007), .ZN(n11008) );
  NAND2_X1 U13613 ( .A1(n14742), .A2(n20690), .ZN(n12605) );
  INV_X1 U13614 ( .A(n13473), .ZN(n16924) );
  NOR2_X1 U13615 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13162), .ZN(
        n13291) );
  INV_X1 U13616 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18061) );
  NOR2_X1 U13617 ( .A1(n13261), .A2(n13260), .ZN(n13262) );
  OR2_X1 U13618 ( .A1(n18305), .A2(n19059), .ZN(n17064) );
  INV_X1 U13619 ( .A(n17286), .ZN(n13152) );
  NAND2_X1 U13620 ( .A1(n13114), .A2(n13299), .ZN(n13125) );
  NAND2_X1 U13621 ( .A1(n13285), .A2(n13264), .ZN(n13350) );
  INV_X1 U13622 ( .A(n19695), .ZN(n19537) );
  OR2_X1 U13623 ( .A1(n12806), .A2(n12805), .ZN(n17097) );
  OR2_X1 U13624 ( .A1(n12344), .A2(n12343), .ZN(n12390) );
  AND2_X1 U13625 ( .A1(n15009), .A2(n12928), .ZN(n14991) );
  XNOR2_X1 U13626 ( .A(n12792), .B(n12791), .ZN(n12913) );
  OR2_X1 U13627 ( .A1(n9699), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12815) );
  NAND2_X1 U13628 ( .A1(n11968), .A2(n11967), .ZN(n14172) );
  NOR2_X1 U13629 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11907) );
  INV_X1 U13630 ( .A(n12802), .ZN(n12803) );
  AOI21_X1 U13631 ( .B1(n15199), .B2(n12273), .A(n12389), .ZN(n14796) );
  NAND2_X1 U13632 ( .A1(n12236), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12274) );
  INV_X1 U13633 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15271) );
  INV_X1 U13634 ( .A(n14873), .ZN(n14942) );
  OR2_X1 U13635 ( .A1(n15504), .A2(n15502), .ZN(n15493) );
  OR2_X1 U13636 ( .A1(n12796), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20893) );
  OAI21_X1 U13637 ( .B1(n17128), .B2(n13799), .A(n13798), .ZN(n13807) );
  OR3_X1 U13638 ( .A1(n13639), .A2(n13638), .A3(n13637), .ZN(n15635) );
  INV_X1 U13639 ( .A(n13940), .ZN(n13968) );
  OR2_X1 U13640 ( .A1(n15659), .A2(n14089), .ZN(n14193) );
  OR2_X1 U13641 ( .A1(n15659), .A2(n21091), .ZN(n15768) );
  OR2_X1 U13642 ( .A1(n21140), .A2(n14089), .ZN(n21054) );
  AND2_X1 U13643 ( .A1(n14014), .A2(n14013), .ZN(n14076) );
  INV_X1 U13644 ( .A(n12639), .ZN(n12611) );
  INV_X1 U13645 ( .A(n16930), .ZN(n13474) );
  NAND2_X1 U13646 ( .A1(n11119), .A2(n11118), .ZN(n11147) );
  NOR2_X1 U13647 ( .A1(n14604), .A2(n14603), .ZN(n16065) );
  AND2_X1 U13648 ( .A1(n11452), .A2(n11451), .ZN(n14370) );
  AND2_X1 U13649 ( .A1(n11447), .A2(n11446), .ZN(n14727) );
  AND3_X1 U13650 ( .A1(n11430), .A2(n11429), .A3(n11428), .ZN(n14162) );
  AND3_X1 U13651 ( .A1(n11364), .A2(n11363), .A3(n11362), .ZN(n13756) );
  OAI21_X1 U13652 ( .B1(n13390), .B2(n13389), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n14164) );
  OR2_X1 U13653 ( .A1(n20637), .A2(n20687), .ZN(n20640) );
  OR2_X1 U13654 ( .A1(n20647), .A2(n20656), .ZN(n20247) );
  NOR3_X1 U13655 ( .A1(n20144), .A2(n20168), .A3(n20463), .ZN(n20150) );
  AND2_X1 U13656 ( .A1(n20313), .A2(n20148), .ZN(n20219) );
  INV_X1 U13657 ( .A(n20634), .ZN(n20628) );
  OR2_X1 U13658 ( .A1(n20647), .A2(n20655), .ZN(n20630) );
  BUF_X1 U13659 ( .A(n10800), .Z(n19976) );
  INV_X1 U13660 ( .A(n20681), .ZN(n16962) );
  NOR2_X1 U13661 ( .A1(n13169), .A2(n13296), .ZN(n13293) );
  INV_X1 U13662 ( .A(n17438), .ZN(n17436) );
  INV_X1 U13663 ( .A(n17799), .ZN(n17791) );
  NOR2_X1 U13664 ( .A1(n19547), .A2(n19523), .ZN(n17417) );
  INV_X1 U13665 ( .A(n18561), .ZN(n18523) );
  INV_X1 U13666 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18567) );
  INV_X1 U13667 ( .A(n13371), .ZN(n13372) );
  NOR2_X1 U13668 ( .A1(n18730), .A2(n18405), .ZN(n18733) );
  INV_X1 U13669 ( .A(n13141), .ZN(n13139) );
  INV_X1 U13670 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13072) );
  NAND2_X1 U13671 ( .A1(n19394), .A2(n19108), .ZN(n19335) );
  INV_X1 U13672 ( .A(n20749), .ZN(n12954) );
  INV_X1 U13673 ( .A(n20759), .ZN(n20772) );
  INV_X1 U13674 ( .A(n12591), .ZN(n12592) );
  INV_X1 U13675 ( .A(n20856), .ZN(n13735) );
  OR2_X1 U13676 ( .A1(n12957), .A2(n12976), .ZN(n17112) );
  INV_X1 U13677 ( .A(n11883), .ZN(n11909) );
  INV_X1 U13678 ( .A(n20933), .ZN(n20922) );
  INV_X1 U13679 ( .A(n20893), .ZN(n20916) );
  NOR2_X1 U13680 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n21291) );
  OAI211_X1 U13681 ( .C1(n15690), .C2(n15689), .A(n15688), .B(n20993), .ZN(
        n15719) );
  OAI211_X1 U13682 ( .C1(n21149), .C2(n13946), .A(n21147), .B(n13945), .ZN(
        n13970) );
  NOR2_X2 U13683 ( .A1(n14066), .A2(n14089), .ZN(n15723) );
  OAI21_X1 U13684 ( .B1(n14223), .B2(n14222), .A(n14221), .ZN(n14248) );
  OAI22_X1 U13685 ( .A1(n14075), .A2(n14074), .B1(n11830), .B2(n14218), .ZN(
        n20953) );
  INV_X1 U13686 ( .A(n14193), .ZN(n20968) );
  NOR2_X2 U13687 ( .A1(n15659), .A2(n14088), .ZN(n15770) );
  INV_X1 U13688 ( .A(n15768), .ZN(n14042) );
  OAI211_X1 U13689 ( .C1(n14123), .C2(n21064), .A(n14122), .B(n20993), .ZN(
        n14148) );
  NOR2_X1 U13690 ( .A1(n21031), .A2(n14089), .ZN(n20987) );
  OAI22_X1 U13691 ( .A1(n20999), .A2(n20998), .B1(n20997), .B2(n21093), .ZN(
        n21016) );
  INV_X1 U13692 ( .A(n21090), .ZN(n21056) );
  OAI22_X1 U13693 ( .A1(n21067), .A2(n21066), .B1(n21094), .B2(n21065), .ZN(
        n21086) );
  NOR2_X2 U13694 ( .A1(n21140), .A2(n14088), .ZN(n21127) );
  NOR2_X1 U13695 ( .A1(n15646), .A2(n15131), .ZN(n21161) );
  NOR2_X1 U13696 ( .A1(n15646), .A2(n15117), .ZN(n21179) );
  OAI211_X1 U13697 ( .C1(n21149), .C2(n21148), .A(n21147), .B(n21146), .ZN(
        n21198) );
  AND2_X1 U13698 ( .A1(n10784), .A2(n20542), .ZN(n13549) );
  AND2_X1 U13699 ( .A1(n11031), .A2(n11030), .ZN(n19805) );
  INV_X1 U13700 ( .A(n19878), .ZN(n19856) );
  AND2_X1 U13701 ( .A1(n12667), .A2(n16958), .ZN(n19864) );
  INV_X1 U13702 ( .A(n19871), .ZN(n19768) );
  OR2_X1 U13703 ( .A1(n11374), .A2(n11373), .ZN(n16140) );
  NOR2_X1 U13704 ( .A1(n14104), .A2(n14103), .ZN(n14102) );
  INV_X1 U13705 ( .A(n13770), .ZN(n13607) );
  INV_X1 U13706 ( .A(n16227), .ZN(n19892) );
  INV_X1 U13707 ( .A(n13399), .ZN(n19935) );
  INV_X1 U13708 ( .A(n14164), .ZN(n16873) );
  AND2_X1 U13709 ( .A1(n14253), .A2(n14180), .ZN(n16682) );
  NOR2_X1 U13710 ( .A1(n14314), .A2(n14315), .ZN(n16328) );
  INV_X1 U13711 ( .A(n19970), .ZN(n16799) );
  AND2_X1 U13712 ( .A1(n11551), .A2(n20674), .ZN(n19958) );
  AND2_X1 U13713 ( .A1(n20634), .A2(n16962), .ZN(n19941) );
  NOR2_X1 U13714 ( .A1(n16826), .A2(n13587), .ZN(n20664) );
  OAI21_X1 U13715 ( .B1(n16880), .B2(n16879), .A(n16878), .ZN(n20003) );
  NOR2_X2 U13716 ( .A1(n20247), .A2(n20146), .ZN(n20030) );
  INV_X1 U13717 ( .A(n20094), .ZN(n20085) );
  OAI21_X1 U13718 ( .B1(n16889), .B2(n20107), .A(n16888), .ZN(n20109) );
  OAI21_X1 U13719 ( .B1(n20121), .B2(n20120), .A(n20119), .ZN(n20138) );
  OAI21_X1 U13720 ( .B1(n20168), .B2(n20276), .A(n20153), .ZN(n20170) );
  NOR2_X2 U13721 ( .A1(n20629), .A2(n20146), .ZN(n20208) );
  OAI21_X1 U13722 ( .B1(n20222), .B2(n20221), .A(n20220), .ZN(n20238) );
  OAI21_X1 U13723 ( .B1(n20311), .B2(n20285), .A(n20284), .ZN(n20305) );
  OAI21_X1 U13724 ( .B1(n20349), .B2(n20352), .A(n20348), .ZN(n20370) );
  NOR2_X2 U13725 ( .A1(n20405), .A2(n20114), .ZN(n20400) );
  NAND2_X1 U13726 ( .A1(n16906), .A2(n16905), .ZN(n20392) );
  AND2_X1 U13727 ( .A1(n20476), .A2(n16913), .ZN(n20436) );
  INV_X1 U13728 ( .A(n20439), .ZN(n20500) );
  NOR2_X1 U13729 ( .A1(n20405), .A2(n20629), .ZN(n20456) );
  INV_X1 U13730 ( .A(n19723), .ZN(n20542) );
  AND3_X1 U13731 ( .A1(n20562), .A2(n20615), .A3(n20547), .ZN(n20692) );
  NOR3_X1 U13732 ( .A1(n21372), .A2(n17498), .A3(n19624), .ZN(n17476) );
  NOR2_X1 U13733 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17660), .ZN(n17638) );
  INV_X1 U13734 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17765) );
  NOR2_X1 U13735 ( .A1(n19056), .A2(n18302), .ZN(n21311) );
  INV_X1 U13736 ( .A(n17417), .ZN(n18304) );
  INV_X1 U13737 ( .A(n18318), .ZN(n18355) );
  OR2_X1 U13738 ( .A1(n13360), .A2(n18725), .ZN(n13345) );
  NAND2_X1 U13739 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18550), .ZN(
        n18532) );
  NOR2_X1 U13740 ( .A1(n18581), .A2(n18567), .ZN(n18562) );
  INV_X1 U13741 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21454) );
  NOR2_X2 U13742 ( .A1(n18222), .A2(n19035), .ZN(n18960) );
  INV_X1 U13743 ( .A(n19193), .ZN(n19186) );
  INV_X1 U13744 ( .A(n19213), .ZN(n19215) );
  INV_X1 U13745 ( .A(n19258), .ZN(n19260) );
  INV_X1 U13746 ( .A(n19317), .ZN(n19329) );
  INV_X1 U13747 ( .A(n19547), .ZN(n19700) );
  AND3_X1 U13748 ( .A1(n19572), .A2(n19630), .A3(n19560), .ZN(n19690) );
  INV_X1 U13749 ( .A(n16873), .ZN(n16872) );
  NAND2_X1 U13750 ( .A1(n15170), .A2(n12954), .ZN(n12942) );
  NAND2_X1 U13751 ( .A1(n20800), .A2(n13758), .ZN(n15070) );
  INV_X1 U13752 ( .A(n15328), .ZN(n15153) );
  INV_X1 U13753 ( .A(n15389), .ZN(n15018) );
  INV_X1 U13754 ( .A(n15155), .ZN(n15161) );
  INV_X1 U13755 ( .A(n20801), .ZN(n20826) );
  NOR2_X1 U13756 ( .A1(n14754), .A2(n13562), .ZN(n13600) );
  OAI21_X1 U13757 ( .B1(n14873), .B2(n14930), .A(n14929), .ZN(n15319) );
  OR2_X1 U13758 ( .A1(n20882), .A2(n13671), .ZN(n20881) );
  INV_X1 U13759 ( .A(n17191), .ZN(n20895) );
  NAND2_X1 U13760 ( .A1(n13030), .A2(n13029), .ZN(n20933) );
  AND2_X1 U13761 ( .A1(n15596), .A2(n15540), .ZN(n20903) );
  INV_X1 U13762 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20942) );
  INV_X1 U13763 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17214) );
  AOI22_X1 U13764 ( .A1(n15684), .A2(n15689), .B1(n15683), .B2(n15682), .ZN(
        n15726) );
  INV_X1 U13765 ( .A(n14247), .ZN(n13973) );
  AOI22_X1 U13766 ( .A1(n14217), .A2(n14222), .B1(n15683), .B2(n15730), .ZN(
        n14251) );
  NAND2_X1 U13767 ( .A1(n14077), .A2(n15679), .ZN(n20972) );
  INV_X1 U13768 ( .A(n13802), .ZN(n13853) );
  INV_X1 U13769 ( .A(n21173), .ZN(n15756) );
  NAND2_X1 U13770 ( .A1(n14004), .A2(n15679), .ZN(n14112) );
  INV_X1 U13771 ( .A(n20987), .ZN(n14151) );
  OR2_X1 U13772 ( .A1(n21031), .A2(n14088), .ZN(n21020) );
  OR2_X1 U13773 ( .A1(n21031), .A2(n21030), .ZN(n21090) );
  INV_X1 U13774 ( .A(n13885), .ZN(n13923) );
  OR2_X1 U13775 ( .A1(n21140), .A2(n21030), .ZN(n21190) );
  INV_X1 U13776 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n17222) );
  INV_X1 U13777 ( .A(n21288), .ZN(n21284) );
  INV_X1 U13778 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20702) );
  INV_X1 U13779 ( .A(n21269), .ZN(n21275) );
  OR2_X1 U13780 ( .A1(n13490), .A2(n16958), .ZN(n19870) );
  OR2_X1 U13781 ( .A1(n19834), .A2(n20276), .ZN(n19878) );
  AND2_X1 U13782 ( .A1(n13589), .A2(n20542), .ZN(n16104) );
  XNOR2_X1 U13783 ( .A(n13771), .B(n13607), .ZN(n20655) );
  AND2_X1 U13784 ( .A1(n13573), .A2(n20542), .ZN(n16287) );
  AND2_X1 U13785 ( .A1(n13578), .A2(n13577), .ZN(n19896) );
  OR2_X1 U13786 ( .A1(n19933), .A2(n13493), .ZN(n13528) );
  NAND2_X1 U13787 ( .A1(n13492), .A2(n20692), .ZN(n19933) );
  NAND2_X1 U13788 ( .A1(n19715), .A2(n20688), .ZN(n13490) );
  OR2_X1 U13789 ( .A1(n16664), .A2(n16663), .ZN(n16665) );
  NAND2_X1 U13790 ( .A1(n11551), .A2(n20670), .ZN(n19970) );
  AOI211_X2 U13791 ( .C1(n16871), .C2(n16879), .A(n20182), .B(n16870), .ZN(
        n20006) );
  NAND2_X1 U13792 ( .A1(n20249), .A2(n20007), .ZN(n20062) );
  NAND2_X1 U13793 ( .A1(n20037), .A2(n20321), .ZN(n20094) );
  INV_X1 U13794 ( .A(n20089), .ZN(n20112) );
  INV_X1 U13795 ( .A(n20134), .ZN(n20142) );
  INV_X1 U13796 ( .A(n20147), .ZN(n20173) );
  INV_X1 U13797 ( .A(n20213), .ZN(n20242) );
  AND2_X1 U13798 ( .A1(n20281), .A2(n20476), .ZN(n20293) );
  INV_X1 U13799 ( .A(n20340), .ZN(n20337) );
  INV_X1 U13800 ( .A(n20350), .ZN(n20374) );
  INV_X1 U13801 ( .A(n20392), .ZN(n20404) );
  INV_X1 U13802 ( .A(n10553), .ZN(n20462) );
  INV_X1 U13803 ( .A(n20456), .ZN(n20534) );
  OR2_X1 U13804 ( .A1(n13552), .A2(n12660), .ZN(n20545) );
  INV_X1 U13805 ( .A(n20627), .ZN(n20546) );
  INV_X1 U13806 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20562) );
  INV_X1 U13807 ( .A(n19698), .ZN(n19710) );
  INV_X1 U13808 ( .A(n13326), .ZN(n17401) );
  NAND2_X1 U13809 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17801), .ZN(n17768) );
  INV_X1 U13810 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18092) );
  OR2_X1 U13811 ( .A1(n18118), .A2(n18259), .ZN(n18112) );
  NAND2_X1 U13812 ( .A1(n19500), .A2(n10207), .ZN(n18242) );
  OR2_X1 U13813 ( .A1(n18300), .A2(n18257), .ZN(n18292) );
  INV_X1 U13814 ( .A(n18257), .ZN(n18302) );
  AOI211_X1 U13815 ( .C1(n19693), .C2(n19691), .A(n18305), .B(n18304), .ZN(
        n18318) );
  INV_X1 U13816 ( .A(n18356), .ZN(n18354) );
  INV_X1 U13817 ( .A(n18635), .ZN(n18609) );
  INV_X1 U13818 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18686) );
  AND2_X1 U13819 ( .A1(n13375), .A2(n13374), .ZN(n13376) );
  INV_X1 U13820 ( .A(n19037), .ZN(n19026) );
  INV_X1 U13821 ( .A(n18960), .ZN(n18935) );
  NAND2_X1 U13822 ( .A1(n18893), .A2(n19037), .ZN(n19006) );
  NAND2_X1 U13823 ( .A1(n19037), .A2(n19525), .ZN(n19035) );
  INV_X1 U13824 ( .A(n19434), .ZN(n19343) );
  INV_X1 U13825 ( .A(n19428), .ZN(n19397) );
  NAND2_X1 U13826 ( .A1(n19552), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19547) );
  INV_X1 U13827 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19650) );
  INV_X1 U13828 ( .A(n19647), .ZN(n19559) );
  INV_X1 U13829 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19572) );
  NAND2_X1 U13830 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19572), .ZN(n19705) );
  NOR2_X1 U13831 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13391), .ZN(n17383)
         );
  NAND2_X1 U13832 ( .A1(n12595), .A2(n12594), .ZN(P1_U2873) );
  NAND2_X1 U13833 ( .A1(n12694), .A2(n12693), .ZN(P2_U2825) );
  INV_X1 U13834 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16616) );
  INV_X1 U13835 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13773) );
  INV_X1 U13836 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10558) );
  AND2_X4 U13837 ( .A1(n16832), .A2(n16920), .ZN(n14512) );
  INV_X1 U13838 ( .A(n10686), .ZN(n10654) );
  NAND2_X1 U13839 ( .A1(n14556), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11139) );
  INV_X1 U13840 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10557) );
  OAI22_X1 U13841 ( .A1(n10558), .A2(n10654), .B1(n11139), .B2(n10557), .ZN(
        n10559) );
  INV_X1 U13842 ( .A(n10559), .ZN(n10564) );
  AND2_X1 U13843 ( .A1(n14513), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10631) );
  AND2_X2 U13844 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10567) );
  AND2_X4 U13845 ( .A1(n10567), .A2(n16920), .ZN(n14515) );
  AOI22_X1 U13846 ( .A1(n14532), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10563) );
  AND2_X4 U13847 ( .A1(n10560), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14514) );
  AOI22_X1 U13848 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n14533), .B1(
        n9596), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10562) );
  AND2_X4 U13849 ( .A1(n11137), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14509) );
  AOI22_X1 U13850 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10888), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10561) );
  NAND4_X1 U13851 ( .A1(n10564), .A2(n10563), .A3(n10562), .A4(n10561), .ZN(
        n10573) );
  AND2_X4 U13852 ( .A1(n10565), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10775) );
  AND2_X4 U13853 ( .A1(n14668), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14538) );
  AOI22_X1 U13854 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n14478), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10571) );
  AND2_X2 U13855 ( .A1(n14509), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10894) );
  AOI22_X1 U13856 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10894), .B1(
        n9597), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10570) );
  AND2_X1 U13857 ( .A1(n10565), .A2(n14507), .ZN(n10895) );
  AOI22_X1 U13858 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U13860 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10568) );
  NAND4_X1 U13861 ( .A1(n10571), .A2(n10570), .A3(n10569), .A4(n10568), .ZN(
        n10572) );
  AOI22_X1 U13862 ( .A1(n14556), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14513), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10577) );
  AOI22_X1 U13863 ( .A1(n14514), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10775), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10576) );
  AOI22_X1 U13864 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14515), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10575) );
  AOI22_X1 U13865 ( .A1(n14516), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10574) );
  NAND4_X1 U13866 ( .A1(n10577), .A2(n10576), .A3(n10575), .A4(n10574), .ZN(
        n10578) );
  NAND2_X1 U13867 ( .A1(n10578), .A2(n10750), .ZN(n10585) );
  AOI22_X1 U13868 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14514), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10582) );
  AOI22_X1 U13869 ( .A1(n14556), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14513), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10581) );
  AOI22_X1 U13870 ( .A1(n14516), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10580) );
  BUF_X4 U13871 ( .A(n10775), .Z(n14678) );
  AOI22_X1 U13872 ( .A1(n14678), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14515), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10579) );
  NAND4_X1 U13873 ( .A1(n10582), .A2(n10581), .A3(n10580), .A4(n10579), .ZN(
        n10583) );
  AOI22_X1 U13874 ( .A1(n14514), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14513), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10587) );
  AOI22_X1 U13875 ( .A1(n14516), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10586) );
  NAND2_X1 U13876 ( .A1(n10587), .A2(n10586), .ZN(n10591) );
  AOI22_X1 U13877 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14556), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U13878 ( .A1(n14678), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14515), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10588) );
  NAND2_X1 U13879 ( .A1(n10589), .A2(n10588), .ZN(n10590) );
  AOI22_X1 U13880 ( .A1(n14514), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14513), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10595) );
  AOI22_X1 U13881 ( .A1(n14516), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10594) );
  AOI22_X1 U13882 ( .A1(n14678), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14515), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U13883 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14556), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10592) );
  NAND4_X1 U13884 ( .A1(n10595), .A2(n10594), .A3(n10593), .A4(n10592), .ZN(
        n10596) );
  NAND2_X1 U13885 ( .A1(n10596), .A2(n10750), .ZN(n10597) );
  NAND2_X1 U13886 ( .A1(n21312), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10599) );
  NAND2_X1 U13887 ( .A1(n10600), .A2(n10599), .ZN(n11127) );
  NAND2_X1 U13888 ( .A1(n16920), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10602) );
  NAND2_X1 U13889 ( .A1(n12672), .A2(n11144), .ZN(n11112) );
  AOI22_X1 U13890 ( .A1(n14513), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14514), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U13891 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14515), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U13892 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14556), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10605) );
  AOI22_X1 U13893 ( .A1(n14516), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10604) );
  NAND4_X1 U13894 ( .A1(n10607), .A2(n10606), .A3(n10605), .A4(n10604), .ZN(
        n10608) );
  NAND2_X1 U13895 ( .A1(n10608), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10615) );
  AOI22_X1 U13896 ( .A1(n14516), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10611) );
  AOI22_X1 U13897 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14515), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10610) );
  AOI22_X1 U13898 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14556), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10609) );
  NAND4_X1 U13899 ( .A1(n10612), .A2(n10611), .A3(n10610), .A4(n10609), .ZN(
        n10613) );
  NAND2_X1 U13900 ( .A1(n10613), .A2(n10750), .ZN(n10614) );
  NOR2_X1 U13901 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10630) );
  AOI22_X1 U13902 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10686), .B1(
        n14533), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10619) );
  INV_X4 U13903 ( .A(n11139), .ZN(n14530) );
  AOI22_X1 U13904 ( .A1(n14530), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9595), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10618) );
  AOI22_X1 U13905 ( .A1(n14532), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10617) );
  AOI22_X1 U13906 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10888), .B1(
        n9598), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10616) );
  NAND4_X1 U13907 ( .A1(n10619), .A2(n10618), .A3(n10617), .A4(n10616), .ZN(
        n10629) );
  AOI22_X1 U13908 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n14539), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10627) );
  AOI22_X1 U13909 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10894), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10626) );
  AOI22_X1 U13910 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10625) );
  AOI22_X1 U13911 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10624) );
  NAND4_X1 U13912 ( .A1(n10627), .A2(n10626), .A3(n10625), .A4(n10624), .ZN(
        n10628) );
  NAND2_X1 U13913 ( .A1(n10963), .A2(n10966), .ZN(n10960) );
  INV_X1 U13914 ( .A(n10960), .ZN(n10652) );
  AOI22_X1 U13915 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n14530), .B1(
        n10686), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10635) );
  AOI22_X1 U13916 ( .A1(n14533), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10634) );
  AOI22_X1 U13917 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n9596), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10633) );
  AOI22_X1 U13918 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10888), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10632) );
  NAND4_X1 U13919 ( .A1(n10635), .A2(n10634), .A3(n10633), .A4(n10632), .ZN(
        n10641) );
  AOI22_X1 U13920 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n14539), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10639) );
  AOI22_X1 U13921 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10894), .B1(
        n9598), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10638) );
  AOI22_X1 U13922 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10637) );
  AOI22_X1 U13923 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10636) );
  NAND4_X1 U13924 ( .A1(n10639), .A2(n10638), .A3(n10637), .A4(n10636), .ZN(
        n10640) );
  INV_X1 U13925 ( .A(n10642), .ZN(n10643) );
  NAND2_X1 U13926 ( .A1(n10644), .A2(n10643), .ZN(n10646) );
  XNOR2_X1 U13927 ( .A(n10670), .B(n10667), .ZN(n11108) );
  INV_X1 U13928 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10655) );
  INV_X1 U13929 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10653) );
  OAI22_X1 U13930 ( .A1(n10655), .A2(n10654), .B1(n11139), .B2(n10653), .ZN(
        n10656) );
  INV_X1 U13931 ( .A(n10656), .ZN(n10660) );
  AOI22_X1 U13932 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10659) );
  AOI22_X1 U13933 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n14533), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U13934 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10888), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10657) );
  NAND4_X1 U13935 ( .A1(n10660), .A2(n10659), .A3(n10658), .A4(n10657), .ZN(
        n10666) );
  AOI22_X1 U13936 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n14539), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10664) );
  AOI22_X1 U13937 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10894), .B1(
        n9598), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10663) );
  AOI22_X1 U13938 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10662) );
  AOI22_X1 U13939 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10661) );
  NAND4_X1 U13940 ( .A1(n10664), .A2(n10663), .A3(n10662), .A4(n10661), .ZN(
        n10665) );
  NOR2_X1 U13941 ( .A1(n10750), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10668) );
  NOR2_X1 U13942 ( .A1(n17144), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10671) );
  NAND2_X1 U13943 ( .A1(n11117), .A2(n10671), .ZN(n11109) );
  MUX2_X1 U13944 ( .A(n11535), .B(n11109), .S(n12672), .Z(n11133) );
  INV_X1 U13945 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n10672) );
  MUX2_X1 U13946 ( .A(n11133), .B(n10672), .S(n11093), .Z(n10971) );
  INV_X1 U13947 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13931) );
  AOI22_X1 U13948 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n14530), .B1(
        n14529), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10677) );
  AOI22_X1 U13949 ( .A1(n9595), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10676) );
  AOI22_X1 U13950 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n14533), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10675) );
  AOI22_X1 U13951 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n10888), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10674) );
  NAND4_X1 U13952 ( .A1(n10677), .A2(n10676), .A3(n10675), .A4(n10674), .ZN(
        n10684) );
  AOI22_X1 U13953 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n14478), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U13954 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n10894), .B1(
        n9597), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U13955 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U13956 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10679) );
  NAND4_X1 U13957 ( .A1(n10682), .A2(n10681), .A3(n10680), .A4(n10679), .ZN(
        n10683) );
  INV_X1 U13958 ( .A(n11327), .ZN(n10685) );
  MUX2_X1 U13959 ( .A(n13931), .B(n10685), .S(n19989), .Z(n10973) );
  AOI22_X1 U13960 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n14530), .B1(
        n14529), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U13961 ( .A1(n9595), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10689) );
  AOI22_X1 U13962 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n14533), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U13963 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10888), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10687) );
  NAND4_X1 U13964 ( .A1(n10690), .A2(n10689), .A3(n10688), .A4(n10687), .ZN(
        n10696) );
  AOI22_X1 U13965 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n14539), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10694) );
  AOI22_X1 U13966 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10894), .B1(
        n9598), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U13967 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U13968 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10691) );
  NAND4_X1 U13969 ( .A1(n10694), .A2(n10693), .A3(n10692), .A4(n10691), .ZN(
        n10695) );
  MUX2_X1 U13970 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n11328), .S(n19989), .Z(
        n10956) );
  INV_X1 U13971 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n14109) );
  AOI22_X1 U13972 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10621), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10700) );
  AOI22_X1 U13973 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10623), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10699) );
  NAND2_X1 U13974 ( .A1(n14478), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10698) );
  NAND2_X1 U13975 ( .A1(n14538), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10697) );
  NAND4_X1 U13976 ( .A1(n10700), .A2(n10699), .A3(n10698), .A4(n10697), .ZN(
        n10704) );
  NAND2_X1 U13977 ( .A1(n10894), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10702) );
  NAND2_X1 U13978 ( .A1(n9598), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10701) );
  NAND2_X1 U13979 ( .A1(n10702), .A2(n10701), .ZN(n10703) );
  NAND2_X1 U13980 ( .A1(n14530), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10708) );
  NAND2_X1 U13981 ( .A1(n14531), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10707) );
  NAND2_X1 U13982 ( .A1(n14532), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10706) );
  NAND2_X1 U13983 ( .A1(n9595), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10705) );
  NAND2_X1 U13984 ( .A1(n14529), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10712) );
  NAND2_X1 U13985 ( .A1(n14533), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10711) );
  NAND2_X1 U13986 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10710) );
  NAND2_X1 U13987 ( .A1(n10888), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10709) );
  MUX2_X1 U13988 ( .A(n14109), .B(n11096), .S(n19989), .Z(n10991) );
  INV_X1 U13989 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n19837) );
  INV_X1 U13990 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n19817) );
  INV_X1 U13991 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n19801) );
  NAND2_X1 U13992 ( .A1(n10717), .A2(n19801), .ZN(n11034) );
  NAND2_X2 U13993 ( .A1(n11034), .A2(n11076), .ZN(n11029) );
  NAND2_X1 U13994 ( .A1(n11093), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11032) );
  INV_X1 U13995 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10718) );
  INV_X1 U13996 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11223) );
  INV_X1 U13997 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11219) );
  INV_X1 U13998 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11018) );
  NAND2_X1 U13999 ( .A1(n11093), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11015) );
  INV_X1 U14000 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n19762) );
  NOR2_X1 U14001 ( .A1(n19989), .A2(n19762), .ZN(n11012) );
  INV_X1 U14002 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n19750) );
  NOR2_X1 U14003 ( .A1(n19989), .A2(n19750), .ZN(n11009) );
  INV_X1 U14004 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n15890) );
  NAND2_X2 U14005 ( .A1(n10723), .A2(n11076), .ZN(n11039) );
  NAND2_X1 U14006 ( .A1(n11093), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10722) );
  NAND2_X1 U14007 ( .A1(n11093), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11041) );
  XNOR2_X1 U14008 ( .A(n11043), .B(n11041), .ZN(n15865) );
  NAND2_X1 U14009 ( .A1(n15865), .A2(n11096), .ZN(n16348) );
  NAND2_X1 U14010 ( .A1(n10723), .A2(n10477), .ZN(n10724) );
  NAND2_X1 U14011 ( .A1(n11043), .A2(n10724), .ZN(n15881) );
  NOR2_X1 U14012 ( .A1(n15881), .A2(n11542), .ZN(n11067) );
  NOR2_X1 U14013 ( .A1(n11067), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16365) );
  AOI22_X1 U14014 ( .A1(n14514), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14513), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U14015 ( .A1(n14516), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10725) );
  NAND2_X1 U14016 ( .A1(n10726), .A2(n10725), .ZN(n10730) );
  AOI22_X1 U14017 ( .A1(n14678), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14515), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10728) );
  AOI22_X1 U14018 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14556), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10727) );
  NAND2_X1 U14019 ( .A1(n10728), .A2(n10727), .ZN(n10729) );
  AOI22_X1 U14020 ( .A1(n14556), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14514), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U14021 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14513), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10733) );
  AOI22_X1 U14022 ( .A1(n14516), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10732) );
  AOI22_X1 U14023 ( .A1(n14678), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14515), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10731) );
  NAND4_X1 U14024 ( .A1(n10734), .A2(n10733), .A3(n10732), .A4(n10731), .ZN(
        n10735) );
  AOI22_X1 U14025 ( .A1(n14514), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14513), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10739) );
  AOI22_X1 U14026 ( .A1(n14516), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10738) );
  AOI22_X1 U14027 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14515), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10737) );
  AOI22_X1 U14028 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14556), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10736) );
  NAND4_X1 U14029 ( .A1(n10739), .A2(n10738), .A3(n10737), .A4(n10736), .ZN(
        n10740) );
  AOI22_X1 U14030 ( .A1(n14514), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14513), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U14031 ( .A1(n14678), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14515), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10743) );
  AOI22_X1 U14032 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n14556), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10742) );
  AOI22_X1 U14033 ( .A1(n14516), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10741) );
  NAND4_X1 U14034 ( .A1(n10744), .A2(n10743), .A3(n10742), .A4(n10741), .ZN(
        n10745) );
  AOI22_X1 U14035 ( .A1(n14514), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14513), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U14036 ( .A1(n14678), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14515), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10748) );
  AOI22_X1 U14037 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14556), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U14038 ( .A1(n14516), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10746) );
  NAND4_X1 U14039 ( .A1(n10749), .A2(n10748), .A3(n10747), .A4(n10746), .ZN(
        n10751) );
  NAND2_X1 U14040 ( .A1(n10751), .A2(n10750), .ZN(n10758) );
  AOI22_X1 U14041 ( .A1(n14678), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14515), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10755) );
  AOI22_X1 U14042 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14556), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10754) );
  AOI22_X1 U14043 ( .A1(n14516), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10753) );
  AOI22_X1 U14044 ( .A1(n14513), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__2__SCAN_IN), .B2(n14514), .ZN(n10752) );
  NAND4_X1 U14045 ( .A1(n10755), .A2(n10754), .A3(n10753), .A4(n10752), .ZN(
        n10756) );
  NAND2_X1 U14046 ( .A1(n10756), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10757) );
  AOI22_X1 U14047 ( .A1(n14514), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14513), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10762) );
  AOI22_X1 U14048 ( .A1(n14678), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14515), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10761) );
  AOI22_X1 U14049 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14556), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10760) );
  AOI22_X1 U14050 ( .A1(n14516), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10759) );
  NAND4_X1 U14051 ( .A1(n10762), .A2(n10761), .A3(n10760), .A4(n10759), .ZN(
        n10763) );
  NAND2_X1 U14052 ( .A1(n10763), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10770) );
  AOI22_X1 U14053 ( .A1(n14514), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14513), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10767) );
  AOI22_X1 U14054 ( .A1(n14678), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14515), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10766) );
  AOI22_X1 U14055 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14556), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10765) );
  AOI22_X1 U14056 ( .A1(n14516), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10764) );
  NAND4_X1 U14057 ( .A1(n10767), .A2(n10766), .A3(n10765), .A4(n10764), .ZN(
        n10768) );
  NAND2_X1 U14058 ( .A1(n10768), .A2(n10750), .ZN(n10769) );
  AOI22_X1 U14059 ( .A1(n14513), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n14514), .ZN(n10774) );
  AOI22_X1 U14060 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n14556), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U14061 ( .A1(n14678), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14515), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U14062 ( .A1(n14516), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14509), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10771) );
  NAND4_X1 U14063 ( .A1(n10774), .A2(n10773), .A3(n10772), .A4(n10771), .ZN(
        n10781) );
  AOI22_X1 U14064 ( .A1(n14513), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__6__SCAN_IN), .B2(n14514), .ZN(n10779) );
  AOI22_X1 U14065 ( .A1(n14512), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14556), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10778) );
  AOI22_X1 U14066 ( .A1(n10775), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14515), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10777) );
  NAND4_X1 U14067 ( .A1(n10779), .A2(n10778), .A3(n10777), .A4(n10776), .ZN(
        n10780) );
  INV_X1 U14068 ( .A(n11287), .ZN(n10785) );
  INV_X2 U14069 ( .A(n10790), .ZN(n13485) );
  AND2_X1 U14070 ( .A1(n10794), .A2(n10786), .ZN(n13575) );
  NAND3_X1 U14071 ( .A1(n11278), .A2(n9591), .A3(n10794), .ZN(n10807) );
  INV_X1 U14072 ( .A(n10807), .ZN(n10795) );
  AND2_X1 U14073 ( .A1(n9782), .A2(n11287), .ZN(n10801) );
  NAND2_X1 U14074 ( .A1(n11481), .A2(n11166), .ZN(n10802) );
  NAND2_X1 U14075 ( .A1(n10802), .A2(n10784), .ZN(n10806) );
  NAND3_X1 U14076 ( .A1(n10811), .A2(n10810), .A3(n9807), .ZN(n10813) );
  INV_X1 U14077 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16825) );
  OAI21_X1 U14078 ( .B1(n20651), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16825), 
        .ZN(n10814) );
  AOI21_X2 U14079 ( .B1(n10821), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10814), .ZN(n10815) );
  INV_X1 U14080 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n10819) );
  NAND2_X1 U14081 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10818) );
  NAND2_X1 U14082 ( .A1(n16818), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10820) );
  NAND2_X1 U14083 ( .A1(n10822), .A2(n9605), .ZN(n16850) );
  AOI22_X1 U14084 ( .A1(n16850), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16962), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10823) );
  INV_X1 U14085 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n16040) );
  NAND2_X1 U14086 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10825) );
  NAND2_X1 U14087 ( .A1(n20681), .A2(n10825), .ZN(n10826) );
  AOI21_X1 U14088 ( .B1(n10835), .B2(P2_REIP_REG_0__SCAN_IN), .A(n10826), .ZN(
        n10827) );
  OAI211_X1 U14089 ( .C1(n16040), .C2(n10836), .A(n10828), .B(n10827), .ZN(
        n10829) );
  INV_X1 U14090 ( .A(n10829), .ZN(n10832) );
  NAND3_X1 U14091 ( .A1(n10830), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n11486), 
        .ZN(n10831) );
  INV_X1 U14092 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U14093 ( .A1(n10835), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10837) );
  BUF_X4 U14094 ( .A(n10836), .Z(n11273) );
  NOR2_X1 U14095 ( .A1(n20681), .A2(n20643), .ZN(n10839) );
  INV_X1 U14096 ( .A(n10847), .ZN(n10852) );
  INV_X1 U14097 ( .A(n10848), .ZN(n10851) );
  INV_X1 U14098 ( .A(n10849), .ZN(n10850) );
  NAND2_X1 U14099 ( .A1(n10852), .A2(n10855), .ZN(n10853) );
  NOR2_X1 U14100 ( .A1(n13766), .A2(n10853), .ZN(n10858) );
  INV_X1 U14101 ( .A(n10853), .ZN(n10854) );
  AND2_X1 U14102 ( .A1(n13766), .A2(n10854), .ZN(n10859) );
  AOI22_X1 U14103 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20315), .B1(
        n20465), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10867) );
  NOR2_X1 U14104 ( .A1(n13766), .A2(n10856), .ZN(n10874) );
  INV_X1 U14105 ( .A(n10856), .ZN(n10857) );
  AND2_X1 U14106 ( .A1(n13766), .A2(n10857), .ZN(n10876) );
  AOI22_X1 U14107 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20008), .B1(
        n16903), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10866) );
  AOI22_X1 U14108 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20069), .B1(
        n20176), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10865) );
  INV_X1 U14109 ( .A(n10873), .ZN(n10862) );
  INV_X1 U14110 ( .A(n13875), .ZN(n16007) );
  NAND2_X2 U14111 ( .A1(n10862), .A2(n10861), .ZN(n10926) );
  INV_X1 U14112 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10863) );
  AND4_X2 U14113 ( .A1(n10867), .A2(n10866), .A3(n10865), .A4(n10864), .ZN(
        n10886) );
  INV_X1 U14114 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10871) );
  NAND2_X1 U14115 ( .A1(n13875), .A2(n14344), .ZN(n10881) );
  INV_X1 U14116 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10870) );
  AOI21_X1 U14117 ( .B1(n20283), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n10872), .ZN(n10885) );
  INV_X1 U14118 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10879) );
  OAI211_X1 U14119 ( .C1(n20143), .C2(n10879), .A(n10878), .B(n10877), .ZN(
        n10880) );
  AOI22_X1 U14120 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16877), .B1(
        n20035), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10883) );
  AOI22_X1 U14121 ( .A1(n14530), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14533), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10892) );
  AOI22_X1 U14122 ( .A1(n14529), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10891) );
  AOI22_X1 U14123 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n10887), .B1(
        n10631), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10890) );
  AOI22_X1 U14124 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n9597), .B1(
        n10888), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10889) );
  NAND4_X1 U14125 ( .A1(n10892), .A2(n10891), .A3(n10890), .A4(n10889), .ZN(
        n10901) );
  AOI22_X1 U14126 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n10893), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10899) );
  AOI22_X1 U14127 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n10620), .B1(
        n10894), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10898) );
  AOI22_X1 U14128 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n10621), .B1(
        n10895), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10897) );
  AOI22_X1 U14129 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10896) );
  NAND4_X1 U14130 ( .A1(n10899), .A2(n10898), .A3(n10897), .A4(n10896), .ZN(
        n10900) );
  OR2_X2 U14131 ( .A1(n10901), .A2(n10900), .ZN(n14338) );
  NAND3_X1 U14132 ( .A1(n20688), .A2(n14338), .A3(n11524), .ZN(n11528) );
  INV_X1 U14133 ( .A(n10902), .ZN(n11527) );
  NAND2_X1 U14134 ( .A1(n11528), .A2(n11527), .ZN(n10903) );
  INV_X1 U14135 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10906) );
  INV_X1 U14136 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10905) );
  INV_X1 U14137 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10908) );
  INV_X1 U14138 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10907) );
  OAI22_X1 U14139 ( .A1(n10908), .A2(n16890), .B1(n10926), .B2(n10907), .ZN(
        n10909) );
  NOR2_X1 U14140 ( .A1(n10910), .A2(n10909), .ZN(n10918) );
  AOI22_X1 U14141 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n9635), .B1(
        n20176), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10914) );
  AOI22_X1 U14142 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20069), .B1(
        n20465), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10913) );
  AOI22_X1 U14143 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20008), .B1(
        n20243), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U14144 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20315), .B1(
        n16903), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U14145 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20035), .B1(
        n20283), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10915) );
  INV_X1 U14146 ( .A(n10919), .ZN(n11314) );
  NAND2_X1 U14147 ( .A1(n11314), .A2(n20688), .ZN(n10920) );
  INV_X1 U14148 ( .A(n11535), .ZN(n11320) );
  AOI22_X1 U14149 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20035), .B1(
        n20283), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10936) );
  AOI22_X1 U14150 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n16877), .B1(
        n10921), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10935) );
  AOI22_X1 U14151 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20008), .B1(
        n16903), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10925) );
  AOI22_X1 U14152 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20315), .B1(
        n20243), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U14153 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n9635), .B1(
        n20465), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U14154 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20069), .B1(
        n20176), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10922) );
  INV_X1 U14155 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10928) );
  INV_X1 U14156 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10927) );
  OAI22_X1 U14157 ( .A1(n10928), .A2(n20143), .B1(n10926), .B2(n10927), .ZN(
        n10932) );
  INV_X1 U14158 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10930) );
  INV_X1 U14159 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10929) );
  NOR2_X1 U14160 ( .A1(n10932), .A2(n10931), .ZN(n10933) );
  NAND2_X1 U14161 ( .A1(n11327), .A2(n20688), .ZN(n10937) );
  AOI22_X1 U14162 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n16877), .B1(
        n20283), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10951) );
  AOI22_X1 U14163 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20035), .B1(
        n10921), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10950) );
  AOI22_X1 U14164 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20176), .B1(
        n16903), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U14165 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20069), .B1(
        n9635), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U14166 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20008), .B1(
        n20243), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U14167 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20315), .B1(
        n20465), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10938) );
  INV_X1 U14168 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10943) );
  INV_X1 U14169 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10942) );
  OAI22_X1 U14170 ( .A1(n10943), .A2(n16890), .B1(n10926), .B2(n10942), .ZN(
        n10947) );
  INV_X1 U14171 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10945) );
  INV_X1 U14172 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10944) );
  NOR2_X1 U14173 ( .A1(n10947), .A2(n10946), .ZN(n10948) );
  NAND4_X1 U14174 ( .A1(n10951), .A2(n10950), .A3(n10949), .A4(n10948), .ZN(
        n10953) );
  NAND2_X1 U14175 ( .A1(n11328), .A2(n20688), .ZN(n10952) );
  INV_X1 U14176 ( .A(n10954), .ZN(n16519) );
  XNOR2_X1 U14177 ( .A(n10976), .B(n10956), .ZN(n19861) );
  NAND2_X1 U14178 ( .A1(n10961), .A2(n10960), .ZN(n10962) );
  NAND2_X1 U14179 ( .A1(n10959), .A2(n10962), .ZN(n16003) );
  INV_X1 U14180 ( .A(n10963), .ZN(n10964) );
  XNOR2_X1 U14181 ( .A(n10964), .B(n10966), .ZN(n16017) );
  INV_X1 U14182 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10965) );
  XNOR2_X1 U14183 ( .A(n16017), .B(n10965), .ZN(n13556) );
  INV_X1 U14184 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19963) );
  OAI21_X1 U14185 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20667), .A(
        n11103), .ZN(n11149) );
  INV_X1 U14186 ( .A(n11149), .ZN(n11105) );
  MUX2_X1 U14187 ( .A(n14338), .B(n11105), .S(n12672), .Z(n11129) );
  MUX2_X1 U14188 ( .A(n11129), .B(P2_EBX_REG_0__SCAN_IN), .S(n11093), .Z(
        n16042) );
  NAND2_X1 U14189 ( .A1(n16042), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14337) );
  AND2_X1 U14190 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19962) );
  NAND2_X1 U14191 ( .A1(n16042), .A2(n19962), .ZN(n10969) );
  INV_X1 U14192 ( .A(n10966), .ZN(n10968) );
  NAND3_X1 U14193 ( .A1(n11093), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n10967) );
  NAND2_X1 U14194 ( .A1(n10968), .A2(n10967), .ZN(n16031) );
  AOI22_X1 U14195 ( .A1(n19963), .A2(n14337), .B1(n10969), .B2(n16031), .ZN(
        n13555) );
  NAND2_X1 U14196 ( .A1(n13556), .A2(n13555), .ZN(n13645) );
  NAND2_X1 U14197 ( .A1(n16017), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10970) );
  NAND2_X1 U14198 ( .A1(n13645), .A2(n10970), .ZN(n16540) );
  XNOR2_X1 U14199 ( .A(n10959), .B(n10971), .ZN(n15991) );
  XNOR2_X1 U14200 ( .A(n15991), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n16807) );
  INV_X1 U14201 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16792) );
  INV_X1 U14202 ( .A(n15991), .ZN(n10972) );
  NOR2_X1 U14203 ( .A1(n11096), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10980) );
  INV_X1 U14204 ( .A(n10980), .ZN(n10978) );
  NAND2_X1 U14205 ( .A1(n10974), .A2(n10016), .ZN(n10975) );
  NAND2_X1 U14206 ( .A1(n10976), .A2(n10975), .ZN(n15976) );
  AND2_X1 U14207 ( .A1(n15976), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10981) );
  INV_X1 U14208 ( .A(n10981), .ZN(n10977) );
  NAND2_X1 U14209 ( .A1(n11096), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10979) );
  MUX2_X1 U14210 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n10979), .S(
        n15976), .Z(n10982) );
  INV_X1 U14211 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16775) );
  INV_X1 U14212 ( .A(n10985), .ZN(n10988) );
  NAND3_X1 U14213 ( .A1(n10995), .A2(n11093), .A3(P2_EBX_REG_8__SCAN_IN), .ZN(
        n10987) );
  AND2_X1 U14214 ( .A1(n10988), .A2(n10987), .ZN(n11003) );
  AND2_X1 U14215 ( .A1(n11096), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10989) );
  NAND2_X1 U14216 ( .A1(n11003), .A2(n10989), .ZN(n16485) );
  INV_X1 U14217 ( .A(n10990), .ZN(n10993) );
  INV_X1 U14218 ( .A(n10991), .ZN(n10992) );
  NAND2_X1 U14219 ( .A1(n10993), .A2(n10992), .ZN(n10994) );
  NAND2_X1 U14220 ( .A1(n10995), .A2(n10994), .ZN(n19851) );
  INV_X1 U14221 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16763) );
  OR2_X1 U14222 ( .A1(n19851), .A2(n16763), .ZN(n16504) );
  NAND2_X1 U14223 ( .A1(n16485), .A2(n16504), .ZN(n16460) );
  INV_X1 U14224 ( .A(n16460), .ZN(n10996) );
  NOR2_X1 U14225 ( .A1(n19989), .A2(n19817), .ZN(n10999) );
  INV_X1 U14226 ( .A(n11076), .ZN(n11045) );
  AOI21_X1 U14227 ( .B1(n11000), .B2(n10999), .A(n11045), .ZN(n11001) );
  AND2_X1 U14228 ( .A1(n10998), .A2(n11001), .ZN(n19819) );
  AOI21_X1 U14229 ( .B1(n19819), .B2(n11096), .A(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16461) );
  INV_X1 U14230 ( .A(n16461), .ZN(n11005) );
  NOR2_X1 U14231 ( .A1(n19989), .A2(n19837), .ZN(n11002) );
  XNOR2_X1 U14232 ( .A(n10985), .B(n11002), .ZN(n19833) );
  AOI21_X1 U14233 ( .B1(n19833), .B2(n11096), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16471) );
  INV_X1 U14234 ( .A(n11003), .ZN(n15960) );
  INV_X1 U14235 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16752) );
  OAI21_X1 U14236 ( .B1(n15960), .B2(n11542), .A(n16752), .ZN(n16486) );
  NAND2_X1 U14237 ( .A1(n19851), .A2(n16763), .ZN(n16503) );
  NAND2_X1 U14238 ( .A1(n16486), .A2(n16503), .ZN(n16458) );
  NOR2_X1 U14239 ( .A1(n16471), .A2(n16458), .ZN(n11004) );
  NAND3_X1 U14240 ( .A1(n19833), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n11096), .ZN(n16472) );
  INV_X1 U14241 ( .A(n16472), .ZN(n11007) );
  NAND2_X1 U14242 ( .A1(n11014), .A2(n11009), .ZN(n11010) );
  NAND2_X1 U14243 ( .A1(n19752), .A2(n11096), .ZN(n11051) );
  INV_X1 U14244 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14363) );
  NAND2_X1 U14245 ( .A1(n11051), .A2(n14363), .ZN(n14345) );
  NAND2_X1 U14246 ( .A1(n11011), .A2(n11012), .ZN(n11013) );
  NAND2_X1 U14247 ( .A1(n11014), .A2(n11013), .ZN(n19763) );
  INV_X1 U14248 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16650) );
  NAND2_X1 U14249 ( .A1(n11064), .A2(n16650), .ZN(n16388) );
  NAND2_X1 U14250 ( .A1(n14345), .A2(n16388), .ZN(n14390) );
  AND2_X1 U14251 ( .A1(n11076), .A2(n11096), .ZN(n11086) );
  NOR2_X1 U14252 ( .A1(n11086), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14393) );
  NOR2_X1 U14253 ( .A1(n14390), .A2(n14393), .ZN(n16377) );
  OR2_X1 U14254 ( .A1(n11016), .A2(n11015), .ZN(n11017) );
  AND2_X1 U14255 ( .A1(n11011), .A2(n11017), .ZN(n11053) );
  AOI21_X1 U14256 ( .B1(n11053), .B2(n11096), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14705) );
  NOR2_X1 U14257 ( .A1(n19989), .A2(n11018), .ZN(n11019) );
  AOI21_X1 U14258 ( .B1(n9677), .B2(n11019), .A(n11045), .ZN(n11020) );
  AND2_X1 U14259 ( .A1(n11021), .A2(n11020), .ZN(n19780) );
  NAND2_X1 U14260 ( .A1(n19780), .A2(n11096), .ZN(n11055) );
  INV_X1 U14261 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16663) );
  XNOR2_X1 U14262 ( .A(n11055), .B(n16663), .ZN(n14709) );
  XNOR2_X1 U14263 ( .A(n11025), .B(n9733), .ZN(n19790) );
  AOI21_X1 U14264 ( .B1(n19790), .B2(n11096), .A(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16405) );
  NAND2_X1 U14265 ( .A1(n11022), .A2(n11023), .ZN(n11024) );
  NAND2_X1 U14266 ( .A1(n11025), .A2(n11024), .ZN(n15922) );
  NAND2_X1 U14267 ( .A1(n11060), .A2(n10376), .ZN(n16417) );
  NAND2_X1 U14268 ( .A1(n11026), .A2(n11027), .ZN(n11028) );
  NAND2_X1 U14269 ( .A1(n11022), .A2(n11028), .ZN(n15928) );
  INV_X1 U14270 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16694) );
  OAI21_X1 U14271 ( .B1(n15928), .B2(n11542), .A(n16694), .ZN(n14352) );
  INV_X1 U14272 ( .A(n11029), .ZN(n11031) );
  NAND3_X1 U14273 ( .A1(n10998), .A2(n11093), .A3(P2_EBX_REG_11__SCAN_IN), 
        .ZN(n11030) );
  NAND2_X1 U14274 ( .A1(n19805), .A2(n11096), .ZN(n16447) );
  INV_X1 U14275 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16451) );
  NAND2_X1 U14276 ( .A1(n16447), .A2(n16451), .ZN(n14347) );
  INV_X1 U14277 ( .A(n11032), .ZN(n11033) );
  NAND2_X1 U14278 ( .A1(n11034), .A2(n11033), .ZN(n11035) );
  NAND2_X1 U14279 ( .A1(n11026), .A2(n11035), .ZN(n15948) );
  INV_X1 U14280 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16713) );
  NAND2_X1 U14281 ( .A1(n14349), .A2(n16713), .ZN(n16434) );
  NAND4_X1 U14282 ( .A1(n16417), .A2(n14352), .A3(n14347), .A4(n16434), .ZN(
        n11036) );
  NOR4_X1 U14283 ( .A1(n14705), .A2(n14709), .A3(n16405), .A4(n11036), .ZN(
        n11040) );
  NOR2_X1 U14284 ( .A1(n19989), .A2(n15890), .ZN(n11037) );
  AND2_X1 U14285 ( .A1(n9706), .A2(n11037), .ZN(n11038) );
  INV_X1 U14286 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16637) );
  NAND2_X1 U14287 ( .A1(n11049), .A2(n16637), .ZN(n16379) );
  INV_X1 U14288 ( .A(n11041), .ZN(n11042) );
  INV_X1 U14289 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n11044) );
  NOR2_X1 U14290 ( .A1(n19989), .A2(n11044), .ZN(n11046) );
  AOI21_X1 U14291 ( .B1(n11047), .B2(n11046), .A(n11045), .ZN(n11048) );
  INV_X1 U14292 ( .A(n15827), .ZN(n11082) );
  INV_X1 U14293 ( .A(n11049), .ZN(n11050) );
  NAND2_X1 U14294 ( .A1(n11050), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16380) );
  INV_X1 U14295 ( .A(n11051), .ZN(n11052) );
  NAND2_X1 U14296 ( .A1(n11052), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14388) );
  INV_X1 U14297 ( .A(n11053), .ZN(n15914) );
  NAND2_X1 U14298 ( .A1(n11096), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11054) );
  INV_X1 U14299 ( .A(n11055), .ZN(n11056) );
  NAND2_X1 U14300 ( .A1(n11056), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14710) );
  INV_X1 U14301 ( .A(n11086), .ZN(n11084) );
  INV_X1 U14302 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14397) );
  OR2_X1 U14303 ( .A1(n11084), .A2(n14397), .ZN(n14392) );
  INV_X1 U14304 ( .A(n16447), .ZN(n16436) );
  NAND2_X1 U14305 ( .A1(n16436), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11057) );
  NAND2_X1 U14306 ( .A1(n16435), .A2(n11057), .ZN(n14346) );
  OR3_X1 U14307 ( .A1(n15928), .A2(n11542), .A3(n16694), .ZN(n14351) );
  INV_X1 U14308 ( .A(n14351), .ZN(n11058) );
  NOR2_X1 U14309 ( .A1(n14346), .A2(n11058), .ZN(n11062) );
  AND2_X1 U14310 ( .A1(n11096), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11059) );
  NAND2_X1 U14311 ( .A1(n19790), .A2(n11059), .ZN(n16406) );
  INV_X1 U14312 ( .A(n11060), .ZN(n11061) );
  NAND4_X1 U14313 ( .A1(n14392), .A2(n11062), .A3(n16406), .A4(n16418), .ZN(
        n11063) );
  NOR2_X1 U14314 ( .A1(n14355), .A2(n11063), .ZN(n11065) );
  AND3_X1 U14315 ( .A1(n14388), .A2(n11065), .A3(n16389), .ZN(n11066) );
  INV_X1 U14316 ( .A(n11067), .ZN(n11068) );
  INV_X1 U14317 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16354) );
  NAND2_X1 U14318 ( .A1(n16366), .A2(n16616), .ZN(n11070) );
  INV_X1 U14319 ( .A(n16348), .ZN(n11069) );
  NAND2_X1 U14320 ( .A1(n11070), .A2(n11069), .ZN(n11071) );
  NAND3_X1 U14321 ( .A1(n16345), .A2(n16346), .A3(n11071), .ZN(n11074) );
  INV_X1 U14322 ( .A(n11072), .ZN(n11073) );
  NAND2_X1 U14323 ( .A1(n11073), .A2(n9891), .ZN(n16344) );
  NOR2_X1 U14324 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(P2_EBX_REG_25__SCAN_IN), 
        .ZN(n11075) );
  NAND2_X1 U14325 ( .A1(n11079), .A2(n11076), .ZN(n11081) );
  NAND2_X1 U14326 ( .A1(n11093), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11077) );
  NAND2_X1 U14327 ( .A1(n11081), .A2(n11077), .ZN(n11089) );
  INV_X1 U14328 ( .A(n11077), .ZN(n11078) );
  NAND2_X1 U14329 ( .A1(n11079), .A2(n11078), .ZN(n11080) );
  NAND2_X1 U14330 ( .A1(n11089), .A2(n11080), .ZN(n15804) );
  INV_X1 U14331 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16551) );
  INV_X1 U14332 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14329) );
  NOR2_X1 U14333 ( .A1(n16551), .A2(n14329), .ZN(n11514) );
  OAI211_X1 U14334 ( .C1(n11082), .C2(P2_EBX_REG_25__SCAN_IN), .A(
        P2_EBX_REG_26__SCAN_IN), .B(n11093), .ZN(n11083) );
  INV_X1 U14335 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16579) );
  OAI21_X1 U14336 ( .B1(n11085), .B2(n11542), .A(n16579), .ZN(n14313) );
  INV_X1 U14337 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16578) );
  NAND2_X1 U14338 ( .A1(n11084), .A2(n16578), .ZN(n16333) );
  OAI211_X1 U14339 ( .C1(n16317), .C2(n11514), .A(n14313), .B(n16333), .ZN(
        n11088) );
  AND2_X1 U14340 ( .A1(n11086), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16326) );
  NOR2_X1 U14341 ( .A1(n14315), .A2(n16326), .ZN(n16315) );
  NAND2_X1 U14342 ( .A1(n11093), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11090) );
  OAI211_X1 U14343 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n15795), .B(n11096), .ZN(
        n11087) );
  INV_X1 U14344 ( .A(n11089), .ZN(n11091) );
  INV_X1 U14345 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n11265) );
  NOR2_X1 U14346 ( .A1(n19989), .A2(n11265), .ZN(n11092) );
  INV_X1 U14347 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16557) );
  OAI21_X1 U14348 ( .B1(n15782), .B2(n11542), .A(n16557), .ZN(n16294) );
  NAND2_X1 U14349 ( .A1(n11093), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11094) );
  AOI21_X1 U14350 ( .B1(n12688), .B2(n11096), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14302) );
  AND2_X1 U14351 ( .A1(n11096), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11095) );
  NAND2_X1 U14352 ( .A1(n12688), .A2(n11095), .ZN(n14300) );
  INV_X1 U14353 ( .A(n15782), .ZN(n11097) );
  NAND3_X1 U14354 ( .A1(n11097), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11096), .ZN(n16293) );
  NOR2_X2 U14355 ( .A1(n11098), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11100) );
  MUX2_X2 U14356 ( .A(n11100), .B(n11099), .S(n19989), .Z(n12673) );
  NAND2_X1 U14357 ( .A1(n12673), .A2(n11096), .ZN(n11101) );
  NAND2_X1 U14358 ( .A1(n13485), .A2(n11144), .ZN(n11107) );
  OAI21_X1 U14359 ( .B1(n11149), .B2(n11127), .A(n10793), .ZN(n11106) );
  XNOR2_X1 U14360 ( .A(n11127), .B(n11103), .ZN(n11145) );
  INV_X1 U14361 ( .A(n11145), .ZN(n11104) );
  NAND2_X1 U14362 ( .A1(n13493), .A2(n11280), .ZN(n11111) );
  INV_X1 U14363 ( .A(n11144), .ZN(n11110) );
  NAND2_X1 U14364 ( .A1(n11111), .A2(n11110), .ZN(n11113) );
  NAND2_X1 U14365 ( .A1(n11113), .A2(n11112), .ZN(n11114) );
  NAND3_X1 U14366 ( .A1(n11115), .A2(n11143), .A3(n11114), .ZN(n11122) );
  NAND2_X1 U14367 ( .A1(n17144), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11116) );
  NAND2_X1 U14368 ( .A1(n11117), .A2(n11116), .ZN(n11119) );
  NAND2_X1 U14369 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16921), .ZN(
        n11118) );
  OAI21_X1 U14370 ( .B1(n11143), .B2(n12672), .A(n11147), .ZN(n11120) );
  INV_X1 U14371 ( .A(n11120), .ZN(n11121) );
  NAND2_X1 U14372 ( .A1(n11122), .A2(n11121), .ZN(n11123) );
  INV_X1 U14373 ( .A(n11147), .ZN(n11125) );
  INV_X1 U14374 ( .A(n13493), .ZN(n11124) );
  NAND2_X2 U14375 ( .A1(n20699), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n20615) );
  NOR2_X1 U14376 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20559) );
  INV_X1 U14377 ( .A(n20559), .ZN(n20547) );
  NAND2_X1 U14378 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20686) );
  NAND2_X1 U14379 ( .A1(n20692), .A2(n20686), .ZN(n16930) );
  NAND3_X1 U14380 ( .A1(n13489), .A2(n13474), .A3(n19976), .ZN(n11178) );
  INV_X1 U14381 ( .A(n11127), .ZN(n11128) );
  NAND2_X1 U14382 ( .A1(n11129), .A2(n11128), .ZN(n11132) );
  INV_X1 U14383 ( .A(n11130), .ZN(n11131) );
  NAND2_X1 U14384 ( .A1(n11132), .A2(n11131), .ZN(n11135) );
  NAND3_X1 U14385 ( .A1(n11135), .A2(n11134), .A3(n11133), .ZN(n11136) );
  AND2_X1 U14386 ( .A1(n11136), .A2(n11147), .ZN(n20678) );
  NAND2_X1 U14387 ( .A1(n20688), .A2(n10784), .ZN(n16959) );
  NOR2_X1 U14388 ( .A1(n11180), .A2(n16959), .ZN(n20670) );
  NAND2_X1 U14389 ( .A1(n20678), .A2(n20670), .ZN(n11154) );
  INV_X1 U14390 ( .A(n11180), .ZN(n16935) );
  AOI21_X1 U14391 ( .B1(n11138), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13483) );
  NAND2_X1 U14392 ( .A1(n11139), .A2(n13483), .ZN(n11141) );
  INV_X1 U14393 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n11140) );
  NAND2_X1 U14394 ( .A1(n11141), .A2(n11140), .ZN(n11142) );
  NAND2_X1 U14395 ( .A1(n11142), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n17247) );
  NAND2_X1 U14396 ( .A1(n11144), .A2(n11143), .ZN(n11148) );
  OAI21_X1 U14397 ( .B1(n11149), .B2(n11148), .A(n16931), .ZN(n11150) );
  INV_X1 U14398 ( .A(n11150), .ZN(n11151) );
  NAND2_X1 U14399 ( .A1(n16825), .A2(n11151), .ZN(n11152) );
  NAND2_X1 U14400 ( .A1(n17247), .A2(n11152), .ZN(n20672) );
  NAND3_X1 U14401 ( .A1(n16935), .A2(n19972), .A3(n20672), .ZN(n11153) );
  NAND2_X1 U14402 ( .A1(n11154), .A2(n11153), .ZN(n13550) );
  INV_X1 U14403 ( .A(n13550), .ZN(n11177) );
  NAND2_X1 U14404 ( .A1(n11155), .A2(n9807), .ZN(n11156) );
  NAND2_X1 U14405 ( .A1(n11157), .A2(n10786), .ZN(n11159) );
  INV_X1 U14406 ( .A(n16959), .ZN(n11158) );
  NAND2_X1 U14407 ( .A1(n11159), .A2(n11158), .ZN(n11489) );
  NAND2_X1 U14408 ( .A1(n20688), .A2(n19984), .ZN(n11484) );
  NAND2_X1 U14409 ( .A1(n11484), .A2(n12597), .ZN(n11161) );
  NAND2_X1 U14410 ( .A1(n11161), .A2(n11160), .ZN(n11162) );
  NAND2_X1 U14411 ( .A1(n11162), .A2(n9807), .ZN(n11163) );
  NAND4_X1 U14412 ( .A1(n11165), .A2(n11164), .A3(n11489), .A4(n11163), .ZN(
        n11485) );
  NAND2_X1 U14413 ( .A1(n16931), .A2(n13474), .ZN(n11167) );
  NOR2_X1 U14414 ( .A1(n16960), .A2(n11167), .ZN(n11168) );
  NOR2_X1 U14415 ( .A1(n11485), .A2(n11168), .ZN(n13477) );
  MUX2_X1 U14416 ( .A(n11169), .B(n19976), .S(n20688), .Z(n11170) );
  NAND3_X1 U14417 ( .A1(n11170), .A2(n16931), .A3(n20686), .ZN(n11171) );
  AND2_X1 U14418 ( .A1(n13477), .A2(n11171), .ZN(n11176) );
  INV_X1 U14419 ( .A(n11172), .ZN(n11174) );
  OAI211_X1 U14420 ( .C1(n11174), .C2(n10784), .A(n11173), .B(n19984), .ZN(
        n11175) );
  NAND4_X1 U14421 ( .A1(n11178), .A2(n11177), .A3(n11176), .A4(n11175), .ZN(
        n11179) );
  AND2_X1 U14422 ( .A1(n16825), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12661) );
  NAND2_X1 U14423 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n12661), .ZN(n19723) );
  AND2_X2 U14424 ( .A1(n11179), .A2(n20542), .ZN(n11551) );
  NOR2_X1 U14425 ( .A1(n11180), .A2(n12672), .ZN(n20674) );
  XNOR2_X1 U14426 ( .A(n11182), .B(n11181), .ZN(n11184) );
  NOR2_X1 U14427 ( .A1(n11182), .A2(n10840), .ZN(n11183) );
  AOI22_X1 U14428 ( .A1(n11267), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11186) );
  NAND2_X1 U14429 ( .A1(n11268), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11185) );
  OAI211_X1 U14430 ( .C1(n11271), .C2(n16792), .A(n11186), .B(n11185), .ZN(
        n14100) );
  INV_X1 U14431 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13980) );
  NAND2_X1 U14432 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11188) );
  NAND2_X1 U14433 ( .A1(n11267), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11187) );
  OAI211_X1 U14434 ( .C1(n11273), .C2(n13980), .A(n11188), .B(n11187), .ZN(
        n11189) );
  AOI21_X1 U14435 ( .B1(n11275), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n11189), .ZN(n13977) );
  INV_X1 U14436 ( .A(n13977), .ZN(n11192) );
  INV_X1 U14437 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16791) );
  AOI22_X1 U14438 ( .A1(n11267), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11191) );
  NAND2_X1 U14439 ( .A1(n11268), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11190) );
  OAI211_X1 U14440 ( .C1(n11271), .C2(n16791), .A(n11191), .B(n11190), .ZN(
        n13929) );
  AND2_X1 U14441 ( .A1(n11192), .A2(n13929), .ZN(n11193) );
  NAND2_X1 U14442 ( .A1(n13928), .A2(n11193), .ZN(n13976) );
  NAND2_X1 U14443 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11195) );
  NAND2_X1 U14444 ( .A1(n11267), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11194) );
  OAI211_X1 U14445 ( .C1(n11273), .C2(n14109), .A(n11195), .B(n11194), .ZN(
        n11196) );
  AOI21_X1 U14446 ( .B1(n11275), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n11196), .ZN(n14107) );
  INV_X1 U14447 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n11201) );
  NAND2_X1 U14448 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11200) );
  NAND2_X1 U14449 ( .A1(n11267), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n11199) );
  OAI211_X1 U14450 ( .C1(n11273), .C2(n11201), .A(n11200), .B(n11199), .ZN(
        n11202) );
  AOI21_X1 U14451 ( .B1(n11275), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n11202), .ZN(n14207) );
  INV_X1 U14452 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16739) );
  AOI22_X1 U14453 ( .A1(n11267), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11204) );
  NAND2_X1 U14454 ( .A1(n11268), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11203) );
  OAI211_X1 U14455 ( .C1(n11271), .C2(n16739), .A(n11204), .B(n11203), .ZN(
        n16147) );
  NAND2_X1 U14456 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11206) );
  NAND2_X1 U14457 ( .A1(n11267), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n11205) );
  OAI211_X1 U14458 ( .C1(n11273), .C2(n19817), .A(n11206), .B(n11205), .ZN(
        n11207) );
  AOI21_X1 U14459 ( .B1(n11275), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n11207), .ZN(n16143) );
  NAND2_X1 U14460 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11211) );
  NAND2_X1 U14461 ( .A1(n11267), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n11210) );
  OAI211_X1 U14462 ( .C1(n11273), .C2(n19801), .A(n11211), .B(n11210), .ZN(
        n11212) );
  AOI21_X1 U14463 ( .B1(n11275), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11212), .ZN(n16131) );
  AOI22_X1 U14464 ( .A1(n11267), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11214) );
  NAND2_X1 U14465 ( .A1(n11268), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11213) );
  OAI211_X1 U14466 ( .C1(n11271), .C2(n16713), .A(n11214), .B(n11213), .ZN(
        n14052) );
  AOI22_X1 U14467 ( .A1(n11267), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11216) );
  NAND2_X1 U14468 ( .A1(n11268), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11215) );
  OAI211_X1 U14469 ( .C1(n11271), .C2(n16694), .A(n11216), .B(n11215), .ZN(
        n14152) );
  NAND2_X1 U14470 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11218) );
  NAND2_X1 U14471 ( .A1(n11267), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11217) );
  OAI211_X1 U14472 ( .C1(n11273), .C2(n11219), .A(n11218), .B(n11217), .ZN(
        n11220) );
  AOI21_X1 U14473 ( .B1(n11275), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n11220), .ZN(n14252) );
  NAND2_X1 U14474 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11222) );
  NAND2_X1 U14475 ( .A1(n11267), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n11221) );
  OAI211_X1 U14476 ( .C1(n11273), .C2(n11223), .A(n11222), .B(n11221), .ZN(
        n11224) );
  AOI21_X1 U14477 ( .B1(n11275), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11224), .ZN(n14179) );
  AOI22_X1 U14478 ( .A1(n11267), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11226) );
  NAND2_X1 U14479 ( .A1(n11268), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11225) );
  OAI211_X1 U14480 ( .C1(n11271), .C2(n16663), .A(n11226), .B(n11225), .ZN(
        n16124) );
  NAND2_X1 U14481 ( .A1(n14254), .A2(n16124), .ZN(n14717) );
  INV_X1 U14482 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n15907) );
  NAND2_X1 U14483 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11228) );
  NAND2_X1 U14484 ( .A1(n11267), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11227) );
  OAI211_X1 U14485 ( .C1(n11273), .C2(n15907), .A(n11228), .B(n11227), .ZN(
        n11229) );
  AOI21_X1 U14486 ( .B1(n11275), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11229), .ZN(n14721) );
  NAND2_X1 U14487 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11231) );
  NAND2_X1 U14488 ( .A1(n11267), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11230) );
  OAI211_X1 U14489 ( .C1(n11273), .C2(n19762), .A(n11231), .B(n11230), .ZN(
        n11232) );
  AOI21_X1 U14490 ( .B1(n11275), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n11232), .ZN(n16110) );
  NAND2_X1 U14491 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11235) );
  NAND2_X1 U14492 ( .A1(n11267), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11234) );
  OAI211_X1 U14493 ( .C1(n11273), .C2(n19750), .A(n11235), .B(n11234), .ZN(
        n11236) );
  AOI21_X1 U14494 ( .B1(n11275), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11236), .ZN(n14365) );
  AOI22_X1 U14495 ( .A1(n11267), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11238) );
  NAND2_X1 U14496 ( .A1(n11268), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11237) );
  OAI211_X1 U14497 ( .C1(n11271), .C2(n14397), .A(n11238), .B(n11237), .ZN(
        n14400) );
  NAND2_X1 U14498 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11240) );
  NAND2_X1 U14499 ( .A1(n11267), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11239) );
  OAI211_X1 U14500 ( .C1(n11273), .C2(n15890), .A(n11240), .B(n11239), .ZN(
        n11241) );
  AOI21_X1 U14501 ( .B1(n11275), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n11241), .ZN(n15885) );
  NOR2_X2 U14502 ( .A1(n14399), .A2(n15885), .ZN(n15867) );
  INV_X1 U14503 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n11244) );
  NAND2_X1 U14504 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11243) );
  NAND2_X1 U14505 ( .A1(n11267), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11242) );
  OAI211_X1 U14506 ( .C1(n11273), .C2(n11244), .A(n11243), .B(n11242), .ZN(
        n11245) );
  AOI21_X1 U14507 ( .B1(n11275), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n11245), .ZN(n15869) );
  AND2_X2 U14508 ( .A1(n15867), .A2(n11246), .ZN(n15854) );
  INV_X1 U14509 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20601) );
  INV_X1 U14510 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16357) );
  OAI22_X1 U14511 ( .A1(n11247), .A2(n20601), .B1(n16825), .B2(n16357), .ZN(
        n11248) );
  AOI21_X1 U14512 ( .B1(n11268), .B2(P2_EBX_REG_23__SCAN_IN), .A(n11248), .ZN(
        n11249) );
  OAI21_X1 U14513 ( .B1(n11271), .B2(n16616), .A(n11249), .ZN(n15856) );
  AOI22_X1 U14514 ( .A1(n11267), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11251) );
  NAND2_X1 U14515 ( .A1(n11268), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11250) );
  OAI211_X1 U14516 ( .C1(n11271), .C2(n9891), .A(n11251), .B(n11250), .ZN(
        n15842) );
  INV_X1 U14517 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15829) );
  NAND2_X1 U14518 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11253) );
  NAND2_X1 U14519 ( .A1(n11267), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11252) );
  OAI211_X1 U14520 ( .C1(n11273), .C2(n15829), .A(n11253), .B(n11252), .ZN(
        n11254) );
  AOI21_X1 U14521 ( .B1(n11275), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n11254), .ZN(n15825) );
  INV_X1 U14522 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n15815) );
  NAND2_X1 U14523 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11256) );
  NAND2_X1 U14524 ( .A1(n11267), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11255) );
  OAI211_X1 U14525 ( .C1(n11273), .C2(n15815), .A(n11256), .B(n11255), .ZN(
        n11257) );
  AOI21_X1 U14526 ( .B1(n11275), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11257), .ZN(n15814) );
  NOR2_X2 U14527 ( .A1(n15813), .A2(n15814), .ZN(n15800) );
  AOI22_X1 U14528 ( .A1(n11267), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11259) );
  NAND2_X1 U14529 ( .A1(n11268), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11258) );
  OAI211_X1 U14530 ( .C1(n11271), .C2(n14329), .A(n11259), .B(n11258), .ZN(
        n15801) );
  INV_X1 U14531 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n15786) );
  NAND2_X1 U14532 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11261) );
  NAND2_X1 U14533 ( .A1(n11267), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11260) );
  OAI211_X1 U14534 ( .C1(n11273), .C2(n15786), .A(n11261), .B(n11260), .ZN(
        n11262) );
  AOI21_X1 U14535 ( .B1(n11275), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n11262), .ZN(n14328) );
  NAND2_X1 U14536 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11264) );
  NAND2_X1 U14537 ( .A1(n11267), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11263) );
  OAI211_X1 U14538 ( .C1(n11273), .C2(n11265), .A(n11264), .B(n11263), .ZN(
        n11266) );
  AOI21_X1 U14539 ( .B1(n11275), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11266), .ZN(n15776) );
  INV_X1 U14540 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11515) );
  AOI22_X1 U14541 ( .A1(n11267), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11270) );
  NAND2_X1 U14542 ( .A1(n11268), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11269) );
  OAI211_X1 U14543 ( .C1(n11271), .C2(n11515), .A(n11270), .B(n11269), .ZN(
        n12680) );
  NAND2_X1 U14544 ( .A1(n15774), .A2(n12680), .ZN(n11277) );
  INV_X1 U14545 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U14546 ( .A1(n11267), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11272) );
  OAI21_X1 U14547 ( .B1(n11273), .B2(n12663), .A(n11272), .ZN(n11274) );
  AOI21_X1 U14548 ( .B1(n11275), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n11274), .ZN(n11276) );
  XNOR2_X2 U14549 ( .A(n11277), .B(n11276), .ZN(n14747) );
  NAND2_X1 U14550 ( .A1(n13574), .A2(n11286), .ZN(n11302) );
  INV_X1 U14551 ( .A(n11302), .ZN(n11279) );
  NAND2_X1 U14552 ( .A1(n11279), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11285) );
  INV_X1 U14553 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n11282) );
  NAND2_X1 U14554 ( .A1(n11280), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11281) );
  OAI211_X1 U14555 ( .C1(n10786), .C2(n11282), .A(n11281), .B(n20276), .ZN(
        n11283) );
  INV_X1 U14556 ( .A(n11283), .ZN(n11284) );
  NAND2_X1 U14557 ( .A1(n11285), .A2(n11284), .ZN(n13609) );
  INV_X1 U14558 ( .A(n14338), .ZN(n11523) );
  NAND2_X1 U14559 ( .A1(n11292), .A2(n11311), .ZN(n11300) );
  AND2_X1 U14560 ( .A1(n20667), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20661) );
  NAND2_X1 U14561 ( .A1(n13609), .A2(n13610), .ZN(n13613) );
  INV_X1 U14562 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20567) );
  OR2_X1 U14563 ( .A1(n11302), .A2(n20567), .ZN(n11291) );
  NOR2_X1 U14564 ( .A1(n10786), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11304) );
  AOI22_X1 U14565 ( .A1(n11304), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11311), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11290) );
  NAND2_X1 U14566 ( .A1(n11291), .A2(n11290), .ZN(n11297) );
  XNOR2_X1 U14567 ( .A(n13613), .B(n11297), .ZN(n16024) );
  MUX2_X1 U14568 ( .A(n11293), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_STATE2_REG_3__SCAN_IN), .Z(n11296) );
  INV_X1 U14569 ( .A(n11524), .ZN(n11294) );
  NOR2_X1 U14570 ( .A1(n11443), .A2(n11294), .ZN(n11295) );
  NOR2_X1 U14571 ( .A1(n11296), .A2(n11295), .ZN(n16023) );
  INV_X1 U14572 ( .A(n11297), .ZN(n11298) );
  NAND2_X1 U14573 ( .A1(n13613), .A2(n11298), .ZN(n11299) );
  NAND2_X1 U14574 ( .A1(n16025), .A2(n11299), .ZN(n11309) );
  OR2_X1 U14575 ( .A1(n11443), .A2(n11527), .ZN(n11301) );
  OAI211_X1 U14576 ( .C1(n20276), .C2(n20651), .A(n11301), .B(n11300), .ZN(
        n11307) );
  XNOR2_X1 U14577 ( .A(n11309), .B(n11307), .ZN(n13648) );
  INV_X1 U14578 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20569) );
  OR2_X1 U14579 ( .A1(n11303), .A2(n20569), .ZN(n11306) );
  AOI22_X1 U14580 ( .A1(n11475), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11305) );
  NAND2_X2 U14581 ( .A1(n13648), .A2(n13647), .ZN(n13650) );
  INV_X1 U14582 ( .A(n11307), .ZN(n11308) );
  NAND2_X1 U14583 ( .A1(n11309), .A2(n11308), .ZN(n11310) );
  AOI22_X1 U14584 ( .A1(n9599), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11313) );
  NAND2_X1 U14585 ( .A1(n11475), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11312) );
  AND2_X1 U14586 ( .A1(n11313), .A2(n11312), .ZN(n11317) );
  OR2_X1 U14587 ( .A1(n11303), .A2(n20571), .ZN(n11316) );
  OR2_X1 U14588 ( .A1(n11443), .A2(n11314), .ZN(n11315) );
  INV_X1 U14589 ( .A(n15996), .ZN(n11318) );
  INV_X1 U14590 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11319) );
  OR2_X1 U14591 ( .A1(n11303), .A2(n11319), .ZN(n11323) );
  AOI22_X1 U14592 ( .A1(n11475), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11322) );
  OR2_X1 U14593 ( .A1(n11443), .A2(n11320), .ZN(n11321) );
  INV_X1 U14594 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n11324) );
  OR2_X1 U14595 ( .A1(n11303), .A2(n11324), .ZN(n11326) );
  AOI22_X1 U14596 ( .A1(n11475), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11325) );
  OAI211_X1 U14597 ( .C1(n11327), .C2(n11443), .A(n11326), .B(n11325), .ZN(
        n15964) );
  NAND2_X1 U14598 ( .A1(n15965), .A2(n15964), .ZN(n15963) );
  OR2_X1 U14599 ( .A1(n11443), .A2(n11328), .ZN(n11329) );
  INV_X1 U14600 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20574) );
  OR2_X1 U14601 ( .A1(n11303), .A2(n20574), .ZN(n11331) );
  AOI22_X1 U14602 ( .A1(n11475), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11330) );
  NAND2_X1 U14603 ( .A1(n11331), .A2(n11330), .ZN(n13567) );
  OR2_X1 U14604 ( .A1(n11443), .A2(n11542), .ZN(n11332) );
  INV_X1 U14605 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20576) );
  OR2_X1 U14606 ( .A1(n11303), .A2(n20576), .ZN(n11335) );
  AOI22_X1 U14607 ( .A1(n11475), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11334) );
  NAND2_X1 U14608 ( .A1(n11335), .A2(n11334), .ZN(n13595) );
  INV_X1 U14609 ( .A(n13593), .ZN(n11351) );
  INV_X1 U14610 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n16490) );
  OR2_X1 U14611 ( .A1(n11303), .A2(n16490), .ZN(n11349) );
  AOI22_X1 U14612 ( .A1(n11475), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11348) );
  AOI22_X1 U14613 ( .A1(n14530), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14529), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11339) );
  AOI22_X1 U14614 ( .A1(n14532), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11338) );
  AOI22_X1 U14615 ( .A1(n14533), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9596), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11337) );
  AOI22_X1 U14616 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n10888), .B1(
        n10894), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11336) );
  NAND4_X1 U14617 ( .A1(n11339), .A2(n11338), .A3(n11337), .A4(n11336), .ZN(
        n11345) );
  AOI22_X1 U14618 ( .A1(n14478), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14619 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9597), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14620 ( .A1(n10621), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U14621 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11340) );
  NAND4_X1 U14622 ( .A1(n11343), .A2(n11342), .A3(n11341), .A4(n11340), .ZN(
        n11344) );
  INV_X1 U14623 ( .A(n14212), .ZN(n11346) );
  OR2_X1 U14624 ( .A1(n11443), .A2(n11346), .ZN(n11347) );
  INV_X1 U14625 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n20579) );
  OR2_X1 U14626 ( .A1(n11303), .A2(n20579), .ZN(n11364) );
  AOI22_X1 U14627 ( .A1(n11475), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14628 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n14530), .B1(
        n14529), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U14629 ( .A1(n9595), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U14630 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n14533), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14631 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n10620), .B1(
        n10888), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11352) );
  NAND4_X1 U14632 ( .A1(n11355), .A2(n11354), .A3(n11353), .A4(n11352), .ZN(
        n11361) );
  AOI22_X1 U14633 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n14478), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U14634 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n10894), .B1(
        n9597), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14635 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14636 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11356) );
  NAND4_X1 U14637 ( .A1(n11359), .A2(n11358), .A3(n11357), .A4(n11356), .ZN(
        n11360) );
  INV_X1 U14638 ( .A(n16152), .ZN(n16133) );
  OR2_X1 U14639 ( .A1(n11443), .A2(n16133), .ZN(n11362) );
  INV_X1 U14640 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20581) );
  OR2_X1 U14641 ( .A1(n11303), .A2(n20581), .ZN(n11377) );
  AOI22_X1 U14642 ( .A1(n11475), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11376) );
  AOI22_X1 U14643 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n14530), .B1(
        n14529), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11368) );
  AOI22_X1 U14644 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11367) );
  AOI22_X1 U14645 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n14533), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11366) );
  AOI22_X1 U14646 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n10620), .B1(
        n10888), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11365) );
  NAND4_X1 U14647 ( .A1(n11368), .A2(n11367), .A3(n11366), .A4(n11365), .ZN(
        n11374) );
  AOI22_X1 U14648 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n14478), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11372) );
  AOI22_X1 U14649 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n9598), .B1(
        n10894), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11371) );
  AOI22_X1 U14650 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11370) );
  AOI22_X1 U14651 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11369) );
  NAND4_X1 U14652 ( .A1(n11372), .A2(n11371), .A3(n11370), .A4(n11369), .ZN(
        n11373) );
  INV_X1 U14653 ( .A(n16140), .ZN(n16135) );
  OR2_X1 U14654 ( .A1(n11443), .A2(n16135), .ZN(n11375) );
  INV_X1 U14655 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n20583) );
  OR2_X1 U14656 ( .A1(n11303), .A2(n20583), .ZN(n11390) );
  AOI22_X1 U14657 ( .A1(n11475), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11389) );
  AOI22_X1 U14658 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n14530), .B1(
        n14529), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11381) );
  AOI22_X1 U14659 ( .A1(n9595), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11380) );
  AOI22_X1 U14660 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n14533), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11379) );
  AOI22_X1 U14661 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10888), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11378) );
  NAND4_X1 U14662 ( .A1(n11381), .A2(n11380), .A3(n11379), .A4(n11378), .ZN(
        n11387) );
  AOI22_X1 U14663 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n14539), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11385) );
  AOI22_X1 U14664 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10894), .B1(
        n9598), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11384) );
  AOI22_X1 U14665 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14666 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11382) );
  NAND4_X1 U14667 ( .A1(n11385), .A2(n11384), .A3(n11383), .A4(n11382), .ZN(
        n11386) );
  NOR2_X1 U14668 ( .A1(n11387), .A2(n11386), .ZN(n16134) );
  OR2_X1 U14669 ( .A1(n11443), .A2(n16134), .ZN(n11388) );
  AOI22_X1 U14670 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n14530), .B1(
        n14529), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11394) );
  AOI22_X1 U14671 ( .A1(n14533), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14672 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n9595), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11392) );
  AOI22_X1 U14673 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n9597), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11391) );
  NAND4_X1 U14674 ( .A1(n11394), .A2(n11393), .A3(n11392), .A4(n11391), .ZN(
        n11400) );
  AOI22_X1 U14675 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n14478), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U14676 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10894), .B1(
        n10888), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14677 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U14678 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11395) );
  NAND4_X1 U14679 ( .A1(n11398), .A2(n11397), .A3(n11396), .A4(n11395), .ZN(
        n11399) );
  INV_X1 U14680 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n16440) );
  OR2_X1 U14681 ( .A1(n11303), .A2(n16440), .ZN(n11402) );
  AOI22_X1 U14682 ( .A1(n11475), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11401) );
  OAI211_X1 U14683 ( .C1(n14063), .C2(n11443), .A(n11402), .B(n11401), .ZN(
        n13857) );
  NAND2_X1 U14684 ( .A1(n13854), .A2(n13857), .ZN(n13855) );
  INV_X1 U14685 ( .A(n13855), .ZN(n11417) );
  INV_X1 U14686 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n16427) );
  OR2_X1 U14687 ( .A1(n11303), .A2(n16427), .ZN(n11415) );
  AOI22_X1 U14688 ( .A1(n11475), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14689 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n14530), .B1(
        n14529), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11406) );
  AOI22_X1 U14690 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11405) );
  AOI22_X1 U14691 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n14533), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11404) );
  AOI22_X1 U14692 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n10620), .B1(
        n10888), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11403) );
  NAND4_X1 U14693 ( .A1(n11406), .A2(n11405), .A3(n11404), .A4(n11403), .ZN(
        n11412) );
  AOI22_X1 U14694 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n14478), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14695 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n10894), .B1(
        n9598), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11409) );
  AOI22_X1 U14696 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11408) );
  AOI22_X1 U14697 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11407) );
  NAND4_X1 U14698 ( .A1(n11410), .A2(n11409), .A3(n11408), .A4(n11407), .ZN(
        n11411) );
  NOR2_X1 U14699 ( .A1(n11412), .A2(n11411), .ZN(n14154) );
  OR2_X1 U14700 ( .A1(n11443), .A2(n14154), .ZN(n11413) );
  INV_X1 U14701 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20587) );
  OR2_X1 U14702 ( .A1(n11303), .A2(n20587), .ZN(n11430) );
  AOI22_X1 U14703 ( .A1(n11475), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11429) );
  AOI22_X1 U14704 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n14530), .B1(
        n14529), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11421) );
  AOI22_X1 U14705 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11420) );
  AOI22_X1 U14706 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n14533), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14707 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10620), .B1(
        n10888), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11418) );
  NAND4_X1 U14708 ( .A1(n11421), .A2(n11420), .A3(n11419), .A4(n11418), .ZN(
        n11427) );
  AOI22_X1 U14709 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n14539), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U14710 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10894), .B1(
        n9598), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U14711 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14712 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11422) );
  NAND4_X1 U14713 ( .A1(n11425), .A2(n11424), .A3(n11423), .A4(n11422), .ZN(
        n11426) );
  NOR2_X1 U14714 ( .A1(n11427), .A2(n11426), .ZN(n14182) );
  OR2_X1 U14715 ( .A1(n11443), .A2(n14182), .ZN(n11428) );
  AOI22_X1 U14716 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n14530), .B1(
        n14529), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U14717 ( .A1(n9595), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11433) );
  AOI22_X1 U14718 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n14533), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11432) );
  AOI22_X1 U14719 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n10620), .B1(
        n10888), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11431) );
  NAND4_X1 U14720 ( .A1(n11434), .A2(n11433), .A3(n11432), .A4(n11431), .ZN(
        n11440) );
  AOI22_X1 U14721 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n14478), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11438) );
  AOI22_X1 U14722 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10894), .B1(
        n9597), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11437) );
  AOI22_X1 U14723 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11436) );
  AOI22_X1 U14724 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11435) );
  NAND4_X1 U14725 ( .A1(n11438), .A2(n11437), .A3(n11436), .A4(n11435), .ZN(
        n11439) );
  NOR2_X1 U14726 ( .A1(n11440), .A2(n11439), .ZN(n14429) );
  INV_X1 U14727 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20589) );
  OR2_X1 U14728 ( .A1(n11303), .A2(n20589), .ZN(n11442) );
  AOI22_X1 U14729 ( .A1(n11475), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11441) );
  OAI211_X1 U14730 ( .C1(n14429), .C2(n11443), .A(n11442), .B(n11441), .ZN(
        n16268) );
  INV_X1 U14731 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20591) );
  OR2_X1 U14732 ( .A1(n11303), .A2(n20591), .ZN(n11445) );
  AOI22_X1 U14733 ( .A1(n11475), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11444) );
  NAND2_X1 U14734 ( .A1(n11445), .A2(n11444), .ZN(n16257) );
  INV_X1 U14735 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20593) );
  OR2_X1 U14736 ( .A1(n11303), .A2(n20593), .ZN(n11447) );
  AOI22_X1 U14737 ( .A1(n11475), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11446) );
  NAND2_X1 U14738 ( .A1(n11279), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U14739 ( .A1(n11475), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11448) );
  INV_X1 U14740 ( .A(n16239), .ZN(n11450) );
  NAND2_X1 U14741 ( .A1(n14726), .A2(n11450), .ZN(n14369) );
  INV_X1 U14742 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20596) );
  OR2_X1 U14743 ( .A1(n11303), .A2(n20596), .ZN(n11452) );
  AOI22_X1 U14744 ( .A1(n11475), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11451) );
  INV_X1 U14745 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n14405) );
  OR2_X1 U14746 ( .A1(n11303), .A2(n14405), .ZN(n11454) );
  AOI22_X1 U14747 ( .A1(n11475), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11311), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11453) );
  NAND2_X1 U14748 ( .A1(n11454), .A2(n11453), .ZN(n14404) );
  NAND2_X1 U14749 ( .A1(n14368), .A2(n14404), .ZN(n14402) );
  INV_X1 U14750 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20599) );
  OR2_X1 U14751 ( .A1(n11303), .A2(n20599), .ZN(n11456) );
  AOI22_X1 U14752 ( .A1(n11475), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11455) );
  NAND2_X1 U14753 ( .A1(n11279), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11459) );
  AOI22_X1 U14754 ( .A1(n11475), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11311), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11458) );
  OR2_X1 U14755 ( .A1(n11303), .A2(n20601), .ZN(n11461) );
  AOI22_X1 U14756 ( .A1(n11475), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11460) );
  NAND2_X1 U14757 ( .A1(n11461), .A2(n11460), .ZN(n15862) );
  NAND2_X1 U14758 ( .A1(n11279), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U14759 ( .A1(n11475), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11462) );
  AND2_X1 U14760 ( .A1(n11463), .A2(n11462), .ZN(n15839) );
  INV_X1 U14761 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20605) );
  OR2_X1 U14762 ( .A1(n11303), .A2(n20605), .ZN(n11465) );
  AOI22_X1 U14763 ( .A1(n11475), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11311), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11464) );
  AND2_X1 U14764 ( .A1(n11465), .A2(n11464), .ZN(n15835) );
  INV_X1 U14765 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20610) );
  OR2_X1 U14766 ( .A1(n11303), .A2(n20610), .ZN(n11467) );
  AOI22_X1 U14767 ( .A1(n11475), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11466) );
  NAND2_X1 U14768 ( .A1(n11467), .A2(n11466), .ZN(n15799) );
  INV_X1 U14769 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20607) );
  OR2_X1 U14770 ( .A1(n11303), .A2(n20607), .ZN(n11469) );
  AOI22_X1 U14771 ( .A1(n11475), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11311), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11468) );
  NAND2_X1 U14772 ( .A1(n11469), .A2(n11468), .ZN(n15810) );
  AND2_X1 U14773 ( .A1(n15799), .A2(n15810), .ZN(n11470) );
  NAND2_X1 U14774 ( .A1(n15798), .A2(n11470), .ZN(n14322) );
  NAND2_X1 U14775 ( .A1(n11279), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11472) );
  AOI22_X1 U14776 ( .A1(n11475), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11311), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11471) );
  AND2_X1 U14777 ( .A1(n11472), .A2(n11471), .ZN(n14323) );
  OR2_X2 U14778 ( .A1(n14322), .A2(n14323), .ZN(n15779) );
  INV_X1 U14779 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20612) );
  OR2_X1 U14780 ( .A1(n11303), .A2(n20612), .ZN(n11474) );
  AOI22_X1 U14781 ( .A1(n11475), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11473) );
  AND2_X1 U14782 ( .A1(n11474), .A2(n11473), .ZN(n15778) );
  INV_X1 U14783 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20616) );
  OR2_X1 U14784 ( .A1(n11303), .A2(n20616), .ZN(n11477) );
  AOI22_X1 U14785 ( .A1(n11475), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n9599), .B2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11476) );
  NAND2_X1 U14786 ( .A1(n11477), .A2(n11476), .ZN(n12681) );
  AOI222_X1 U14787 ( .A1(n11279), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n11475), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11311), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11478) );
  XNOR2_X2 U14788 ( .A(n12683), .B(n11478), .ZN(n12600) );
  INV_X1 U14789 ( .A(n11481), .ZN(n11482) );
  NAND2_X1 U14790 ( .A1(n11480), .A2(n11482), .ZN(n13473) );
  OAI21_X1 U14791 ( .B1(n20688), .B2(n16934), .A(n13473), .ZN(n11483) );
  NAND2_X1 U14792 ( .A1(n11551), .A2(n16926), .ZN(n14712) );
  AND2_X1 U14793 ( .A1(n10792), .A2(n11486), .ZN(n11487) );
  NAND2_X1 U14794 ( .A1(n10830), .A2(n11487), .ZN(n11498) );
  NAND2_X1 U14795 ( .A1(n11488), .A2(n19972), .ZN(n16819) );
  NAND2_X1 U14796 ( .A1(n9799), .A2(n13485), .ZN(n13570) );
  NAND2_X1 U14797 ( .A1(n13570), .A2(n20689), .ZN(n11490) );
  NAND2_X1 U14798 ( .A1(n11490), .A2(n10792), .ZN(n11494) );
  OAI22_X1 U14799 ( .A1(n20689), .A2(n9591), .B1(n9807), .B2(n12597), .ZN(
        n11491) );
  INV_X1 U14800 ( .A(n11491), .ZN(n11493) );
  NAND3_X1 U14801 ( .A1(n11494), .A2(n11493), .A3(n11492), .ZN(n11495) );
  NOR2_X1 U14802 ( .A1(n11496), .A2(n11495), .ZN(n11497) );
  NAND2_X1 U14803 ( .A1(n16830), .A2(n9605), .ZN(n11499) );
  NAND2_X1 U14804 ( .A1(n11551), .A2(n11499), .ZN(n14714) );
  OR2_X1 U14805 ( .A1(n19961), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11502) );
  NOR2_X1 U14806 ( .A1(n11551), .A2(n19941), .ZN(n17241) );
  NAND2_X1 U14807 ( .A1(n19962), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13659) );
  INV_X1 U14808 ( .A(n13659), .ZN(n11500) );
  NOR2_X1 U14809 ( .A1(n14714), .A2(n11500), .ZN(n13651) );
  INV_X1 U14810 ( .A(n14712), .ZN(n11501) );
  NOR2_X1 U14811 ( .A1(n19962), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13654) );
  AND2_X1 U14812 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11545) );
  NOR2_X1 U14813 ( .A1(n16792), .A2(n16791), .ZN(n16790) );
  NAND2_X1 U14814 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16790), .ZN(
        n11512) );
  INV_X1 U14815 ( .A(n11512), .ZN(n11503) );
  AND2_X1 U14816 ( .A1(n11545), .A2(n11503), .ZN(n11504) );
  NOR2_X1 U14817 ( .A1(n19961), .A2(n11504), .ZN(n11505) );
  NAND2_X1 U14818 ( .A1(n16740), .A2(n19961), .ZN(n16685) );
  NAND2_X1 U14819 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16716) );
  NOR2_X1 U14820 ( .A1(n16716), .A2(n16739), .ZN(n16683) );
  NAND2_X1 U14821 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16679) );
  NOR2_X1 U14822 ( .A1(n16679), .A2(n10376), .ZN(n16681) );
  NAND2_X1 U14823 ( .A1(n16683), .A2(n16681), .ZN(n16668) );
  INV_X1 U14824 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16412) );
  OR2_X1 U14825 ( .A1(n16668), .A2(n16412), .ZN(n14361) );
  NAND2_X1 U14826 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14362) );
  OR2_X1 U14827 ( .A1(n14361), .A2(n14362), .ZN(n14373) );
  AND2_X1 U14828 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16638) );
  NAND2_X1 U14829 ( .A1(n16638), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11506) );
  NOR2_X1 U14830 ( .A1(n14373), .A2(n11506), .ZN(n14396) );
  AND2_X1 U14831 ( .A1(n14396), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11547) );
  NAND2_X1 U14832 ( .A1(n16740), .A2(n11547), .ZN(n11507) );
  NAND2_X1 U14833 ( .A1(n16685), .A2(n11507), .ZN(n16625) );
  NAND2_X1 U14834 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16613) );
  INV_X1 U14835 ( .A(n16613), .ZN(n16602) );
  OR2_X1 U14836 ( .A1(n19961), .A2(n16602), .ZN(n11508) );
  NAND2_X1 U14837 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11548) );
  AOI21_X1 U14838 ( .B1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n11514), .A(
        n19961), .ZN(n11509) );
  NOR3_X1 U14839 ( .A1(n16570), .A2(n11509), .A3(n11515), .ZN(n14306) );
  INV_X1 U14840 ( .A(n16685), .ZN(n11511) );
  INV_X1 U14841 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11510) );
  NAND2_X1 U14842 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17224), .ZN(
        n16789) );
  NOR2_X1 U14843 ( .A1(n16613), .A2(n9891), .ZN(n11513) );
  NAND2_X1 U14844 ( .A1(n16623), .A2(n11513), .ZN(n16590) );
  NOR2_X1 U14845 ( .A1(n16590), .A2(n11548), .ZN(n16552) );
  NAND2_X1 U14846 ( .A1(n16552), .A2(n11514), .ZN(n14305) );
  NOR4_X1 U14847 ( .A1(n14305), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16557), .A4(n11515), .ZN(n11516) );
  INV_X2 U14848 ( .A(n19941), .ZN(n16491) );
  INV_X1 U14849 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20618) );
  NOR2_X1 U14850 ( .A1(n16491), .A2(n20618), .ZN(n14743) );
  NOR2_X1 U14851 ( .A1(n11516), .A2(n14743), .ZN(n11517) );
  OAI21_X1 U14852 ( .B1(n12600), .B2(n17237), .A(n11518), .ZN(n11519) );
  INV_X1 U14853 ( .A(n11519), .ZN(n11520) );
  OAI21_X1 U14854 ( .B1(n14747), .B2(n16782), .A(n11520), .ZN(n11521) );
  NAND3_X1 U14855 ( .A1(n11523), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n11524), .ZN(n11526) );
  NOR2_X1 U14856 ( .A1(n14338), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11525) );
  XNOR2_X1 U14857 ( .A(n11525), .B(n11524), .ZN(n14294) );
  NAND2_X1 U14858 ( .A1(n14294), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14293) );
  NAND2_X1 U14859 ( .A1(n11526), .A2(n14293), .ZN(n11529) );
  XOR2_X1 U14860 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11529), .Z(
        n13548) );
  XNOR2_X1 U14861 ( .A(n11528), .B(n11527), .ZN(n13547) );
  NAND2_X1 U14862 ( .A1(n13548), .A2(n13547), .ZN(n11531) );
  NAND2_X1 U14863 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11529), .ZN(
        n11530) );
  NAND2_X1 U14864 ( .A1(n11531), .A2(n11530), .ZN(n11532) );
  XNOR2_X1 U14865 ( .A(n11532), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16538) );
  NAND2_X1 U14866 ( .A1(n11532), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11533) );
  OAI21_X1 U14867 ( .B1(n16495), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11544) );
  AOI22_X1 U14868 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U14869 ( .A1(n11761), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12352), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U14870 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11555) );
  AND2_X4 U14871 ( .A1(n15666), .A2(n11553), .ZN(n12403) );
  AOI22_X1 U14872 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11554) );
  INV_X1 U14873 ( .A(n11767), .ZN(n11587) );
  NAND2_X1 U14874 ( .A1(n11587), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11562) );
  AND3_X2 U14875 ( .A1(n15615), .A2(n13664), .A3(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12295) );
  AOI22_X1 U14876 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11561) );
  NAND2_X1 U14877 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11560) );
  NAND2_X1 U14878 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11559) );
  NAND4_X1 U14879 ( .A1(n11562), .A2(n11561), .A3(n11560), .A4(n11559), .ZN(
        n11570) );
  INV_X1 U14880 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11568) );
  NAND2_X1 U14881 ( .A1(n11772), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11567) );
  NAND2_X1 U14882 ( .A1(n11745), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11566) );
  OAI211_X1 U14883 ( .C1(n11667), .C2(n11568), .A(n11567), .B(n11566), .ZN(
        n11569) );
  NAND2_X1 U14884 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11574) );
  AOI22_X1 U14885 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11573) );
  NAND2_X1 U14886 ( .A1(n12218), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11572) );
  NAND2_X1 U14887 ( .A1(n11732), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11571) );
  NAND2_X1 U14888 ( .A1(n11745), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11578) );
  NAND2_X1 U14889 ( .A1(n11761), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11577) );
  NAND2_X1 U14890 ( .A1(n12352), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11576) );
  NAND2_X1 U14891 ( .A1(n12403), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11575) );
  NAND2_X1 U14892 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11582) );
  NAND2_X1 U14893 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11581) );
  NAND2_X1 U14894 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11580) );
  NAND2_X1 U14895 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11579) );
  INV_X1 U14896 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11585) );
  NAND2_X1 U14897 ( .A1(n11772), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11584) );
  NAND2_X1 U14898 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11583) );
  OAI211_X1 U14899 ( .C1(n11767), .C2(n11585), .A(n11584), .B(n11583), .ZN(
        n11586) );
  INV_X1 U14900 ( .A(n11586), .ZN(n11604) );
  NAND4_X2 U14901 ( .A1(n11607), .A2(n11606), .A3(n11605), .A4(n11604), .ZN(
        n11695) );
  AND2_X2 U14902 ( .A1(n11827), .A2(n11695), .ZN(n11706) );
  NAND2_X1 U14903 ( .A1(n11587), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11591) );
  AOI22_X1 U14904 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11590) );
  NAND2_X1 U14905 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11589) );
  NAND2_X1 U14906 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11588) );
  NAND4_X1 U14907 ( .A1(n11591), .A2(n11590), .A3(n11589), .A4(n11588), .ZN(
        n11596) );
  NAND2_X1 U14908 ( .A1(n11772), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11593) );
  NAND2_X1 U14909 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11592) );
  AOI22_X1 U14910 ( .A1(n12352), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U14911 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U14912 ( .A1(n11745), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U14913 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11597) );
  NAND2_X2 U14914 ( .A1(n11601), .A2(n9644), .ZN(n11752) );
  NAND2_X1 U14915 ( .A1(n11706), .A2(n13845), .ZN(n11628) );
  AND4_X2 U14916 ( .A1(n11607), .A2(n11606), .A3(n11605), .A4(n11604), .ZN(
        n13808) );
  NAND2_X1 U14917 ( .A1(n11587), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11611) );
  AOI22_X1 U14918 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11610) );
  NAND2_X1 U14919 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11609) );
  NAND2_X1 U14920 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11608) );
  NAND2_X1 U14921 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11615) );
  NAND2_X1 U14922 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11614) );
  NAND2_X1 U14923 ( .A1(n12218), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11613) );
  NAND2_X1 U14924 ( .A1(n11732), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11612) );
  NAND2_X1 U14925 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11619) );
  NAND2_X1 U14926 ( .A1(n11761), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11618) );
  NAND2_X1 U14927 ( .A1(n12352), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11617) );
  NAND2_X1 U14928 ( .A1(n12403), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11616) );
  NAND2_X1 U14929 ( .A1(n11772), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11621) );
  NAND2_X1 U14930 ( .A1(n11745), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11620) );
  OAI211_X1 U14931 ( .C1(n11667), .C2(n12491), .A(n11621), .B(n11620), .ZN(
        n11622) );
  INV_X1 U14932 ( .A(n11622), .ZN(n11623) );
  INV_X1 U14933 ( .A(n11829), .ZN(n11627) );
  NAND2_X1 U14934 ( .A1(n11752), .A2(n11829), .ZN(n11696) );
  AOI22_X1 U14935 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11632) );
  AOI22_X1 U14936 ( .A1(n11761), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12352), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11631) );
  AOI22_X1 U14937 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U14938 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U14939 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11637) );
  INV_X1 U14940 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11633) );
  NAND2_X1 U14941 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11635) );
  NAND2_X1 U14942 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11634) );
  NAND4_X1 U14943 ( .A1(n11637), .A2(n11636), .A3(n11635), .A4(n11634), .ZN(
        n11642) );
  INV_X1 U14944 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11640) );
  NAND2_X1 U14945 ( .A1(n11772), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11639) );
  NAND2_X1 U14946 ( .A1(n11745), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11638) );
  OAI211_X1 U14947 ( .C1(n11667), .C2(n11640), .A(n11639), .B(n11638), .ZN(
        n11641) );
  INV_X1 U14948 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11647) );
  NAND2_X1 U14949 ( .A1(n11772), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11646) );
  NAND2_X1 U14950 ( .A1(n11745), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11645) );
  OAI211_X1 U14951 ( .C1(n11667), .C2(n11647), .A(n11646), .B(n11645), .ZN(
        n11648) );
  INV_X1 U14952 ( .A(n11648), .ZN(n11652) );
  AOI22_X1 U14953 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14954 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11650) );
  NAND2_X1 U14955 ( .A1(n11587), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11649) );
  NAND4_X1 U14956 ( .A1(n11652), .A2(n11651), .A3(n11650), .A4(n11649), .ZN(
        n11658) );
  AOI22_X1 U14957 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11732), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U14958 ( .A1(n11761), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12352), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11655) );
  AOI22_X1 U14959 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12218), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11654) );
  AOI22_X1 U14960 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11653) );
  NAND4_X1 U14961 ( .A1(n11656), .A2(n11655), .A3(n11654), .A4(n11653), .ZN(
        n11657) );
  NAND2_X1 U14962 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11663) );
  NAND2_X1 U14963 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11662) );
  NAND2_X1 U14964 ( .A1(n12218), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11661) );
  NAND2_X1 U14965 ( .A1(n11732), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11660) );
  NAND2_X1 U14966 ( .A1(n11772), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11665) );
  OAI211_X1 U14967 ( .C1(n11667), .C2(n11666), .A(n11665), .B(n11664), .ZN(
        n11668) );
  INV_X1 U14968 ( .A(n11668), .ZN(n11674) );
  NAND2_X1 U14969 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11672) );
  NAND2_X1 U14970 ( .A1(n11761), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11671) );
  NAND2_X1 U14971 ( .A1(n12352), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11670) );
  NAND2_X1 U14972 ( .A1(n12403), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11669) );
  AOI22_X1 U14973 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11678) );
  NAND2_X1 U14974 ( .A1(n11587), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11677) );
  NAND2_X1 U14975 ( .A1(n11868), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11676) );
  NAND2_X1 U14976 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11675) );
  NAND2_X4 U14977 ( .A1(n11680), .A2(n11679), .ZN(n13777) );
  NAND2_X1 U14978 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n21220) );
  OAI21_X1 U14979 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(n21220), .ZN(n12915) );
  AOI22_X1 U14980 ( .A1(n11787), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11868), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11684) );
  AOI22_X1 U14981 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12352), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14982 ( .A1(n11772), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U14983 ( .A1(n11745), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11681) );
  NAND2_X1 U14984 ( .A1(n12218), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11688) );
  NAND2_X1 U14985 ( .A1(n11732), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11687) );
  NAND2_X1 U14986 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11686) );
  NAND2_X1 U14987 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11685) );
  NAND2_X1 U14988 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11691) );
  NAND2_X1 U14989 ( .A1(n11587), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11690) );
  NAND3_X4 U14990 ( .A1(n11694), .A2(n11693), .A3(n11692), .ZN(n13563) );
  NAND3_X1 U14992 ( .A1(n13839), .A2(n11695), .A3(n12575), .ZN(n11703) );
  INV_X1 U14993 ( .A(n11696), .ZN(n11697) );
  NAND2_X1 U14994 ( .A1(n11698), .A2(n13823), .ZN(n11699) );
  NAND2_X2 U14995 ( .A1(n11702), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11719) );
  NAND2_X1 U14996 ( .A1(n11704), .A2(n11703), .ZN(n12806) );
  NAND2_X1 U14997 ( .A1(n12806), .A2(n13818), .ZN(n12980) );
  NAND2_X1 U14998 ( .A1(n13777), .A2(n13636), .ZN(n12983) );
  NAND3_X1 U14999 ( .A1(n11705), .A2(n12980), .A3(n9601), .ZN(n11718) );
  XNOR2_X1 U15000 ( .A(n12958), .B(n13845), .ZN(n11708) );
  INV_X1 U15001 ( .A(n15613), .ZN(n11716) );
  NAND2_X1 U15002 ( .A1(n12959), .A2(n11716), .ZN(n11709) );
  OAI21_X2 U15003 ( .B1(n11718), .B2(n11709), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11710) );
  NAND2_X1 U15004 ( .A1(n21291), .A2(n11759), .ZN(n12796) );
  NAND2_X1 U15005 ( .A1(n21136), .A2(n14084), .ZN(n21053) );
  NAND2_X1 U15006 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21132) );
  NAND2_X1 U15007 ( .A1(n21053), .A2(n21132), .ZN(n20992) );
  NAND2_X1 U15008 ( .A1(n21203), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11720) );
  OAI21_X1 U15009 ( .B1(n12796), .B2(n20992), .A(n11720), .ZN(n11711) );
  INV_X1 U15010 ( .A(n11711), .ZN(n11712) );
  INV_X1 U15011 ( .A(n21203), .ZN(n17124) );
  MUX2_X1 U15012 ( .A(n17124), .B(n12796), .S(n14084), .Z(n11811) );
  INV_X1 U15013 ( .A(n12959), .ZN(n11713) );
  NAND2_X1 U15014 ( .A1(n11713), .A2(n13563), .ZN(n11717) );
  INV_X1 U15015 ( .A(n17109), .ZN(n15027) );
  INV_X4 U15016 ( .A(n9699), .ZN(n12943) );
  NAND2_X1 U15017 ( .A1(n12958), .A2(n12719), .ZN(n11715) );
  INV_X1 U15018 ( .A(n11707), .ZN(n11714) );
  INV_X1 U15019 ( .A(n21291), .ZN(n17211) );
  OR2_X1 U15020 ( .A1(n11716), .A2(n12575), .ZN(n12984) );
  NAND2_X2 U15021 ( .A1(n14010), .A2(n11757), .ZN(n11756) );
  NAND2_X1 U15022 ( .A1(n11720), .A2(n13621), .ZN(n11721) );
  NAND2_X1 U15023 ( .A1(n11756), .A2(n11728), .ZN(n11726) );
  AOI21_X2 U15024 ( .B1(n11723), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11724), .ZN(n11729) );
  INV_X1 U15025 ( .A(n12796), .ZN(n13515) );
  XNOR2_X1 U15026 ( .A(n21132), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14120) );
  NAND2_X1 U15027 ( .A1(n13515), .A2(n14120), .ZN(n11727) );
  NAND2_X1 U15028 ( .A1(n11729), .A2(n11727), .ZN(n11725) );
  NAND4_X1 U15029 ( .A1(n11756), .A2(n11729), .A3(n11728), .A4(n11727), .ZN(
        n11730) );
  INV_X1 U15030 ( .A(n12218), .ZN(n12246) );
  AOI22_X1 U15031 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U15032 ( .A1(n11795), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U15033 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11735) );
  AOI22_X1 U15034 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11734) );
  INV_X1 U15035 ( .A(n12295), .ZN(n12351) );
  INV_X2 U15036 ( .A(n12317), .ZN(n11867) );
  AOI22_X1 U15037 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11743) );
  NAND2_X1 U15038 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n11742) );
  NAND2_X1 U15039 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11741) );
  INV_X1 U15040 ( .A(n11739), .ZN(n11766) );
  NAND2_X1 U15041 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11740) );
  NAND4_X1 U15042 ( .A1(n11743), .A2(n11742), .A3(n11741), .A4(n11740), .ZN(
        n11750) );
  INV_X1 U15043 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11748) );
  INV_X2 U15044 ( .A(n12407), .ZN(n12459) );
  NAND2_X1 U15045 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11747) );
  INV_X1 U15046 ( .A(n11745), .ZN(n11760) );
  NAND2_X1 U15047 ( .A1(n12460), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11746) );
  OAI211_X1 U15048 ( .C1(n12199), .C2(n11748), .A(n11747), .B(n11746), .ZN(
        n11749) );
  NOR2_X1 U15049 ( .A1(n11750), .A2(n11749), .ZN(n11751) );
  AND2_X1 U15050 ( .A1(n10540), .A2(n11751), .ZN(n12727) );
  INV_X1 U15051 ( .A(n12727), .ZN(n11753) );
  AOI22_X1 U15052 ( .A1(n13523), .A2(n11753), .B1(n12543), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11754) );
  INV_X1 U15053 ( .A(n14010), .ZN(n11758) );
  INV_X1 U15054 ( .A(n11862), .ZN(n11816) );
  INV_X1 U15055 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11764) );
  NAND2_X1 U15056 ( .A1(n12460), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11763) );
  INV_X1 U15057 ( .A(n11761), .ZN(n12287) );
  NAND2_X1 U15058 ( .A1(n11795), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11762) );
  OAI211_X1 U15059 ( .C1(n12199), .C2(n11764), .A(n11763), .B(n11762), .ZN(
        n11765) );
  INV_X1 U15060 ( .A(n11765), .ZN(n11771) );
  AOI22_X1 U15061 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11770) );
  AOI22_X1 U15062 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11769) );
  NAND2_X1 U15063 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11768) );
  NAND4_X1 U15064 ( .A1(n11771), .A2(n11770), .A3(n11769), .A4(n11768), .ZN(
        n11778) );
  INV_X1 U15065 ( .A(n11772), .ZN(n12407) );
  AOI22_X1 U15066 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U15067 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U15068 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U15069 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11773) );
  NAND4_X1 U15070 ( .A1(n11776), .A2(n11775), .A3(n11774), .A4(n11773), .ZN(
        n11777) );
  NAND2_X1 U15071 ( .A1(n11816), .A2(n12714), .ZN(n11779) );
  INV_X1 U15072 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12478) );
  NAND2_X1 U15073 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11781) );
  NAND2_X1 U15074 ( .A1(n12460), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11780) );
  OAI211_X1 U15075 ( .C1(n12199), .C2(n12478), .A(n11781), .B(n11780), .ZN(
        n11782) );
  INV_X1 U15076 ( .A(n11782), .ZN(n11786) );
  AOI22_X1 U15077 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11785) );
  AOI22_X1 U15078 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11784) );
  NAND2_X1 U15079 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11783) );
  NAND4_X1 U15080 ( .A1(n11786), .A2(n11785), .A3(n11784), .A4(n11783), .ZN(
        n11794) );
  INV_X1 U15081 ( .A(n11787), .ZN(n11803) );
  INV_X1 U15082 ( .A(n11803), .ZN(n11788) );
  AOI22_X1 U15083 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U15084 ( .A1(n11795), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U15085 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11790) );
  AOI22_X1 U15086 ( .A1(n11733), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11789) );
  NAND4_X1 U15087 ( .A1(n11792), .A2(n11791), .A3(n11790), .A4(n11789), .ZN(
        n11793) );
  INV_X1 U15088 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11815) );
  NAND2_X1 U15089 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11797) );
  NAND2_X1 U15090 ( .A1(n11795), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11796) );
  OAI211_X1 U15091 ( .C1(n12199), .C2(n11815), .A(n11797), .B(n11796), .ZN(
        n11798) );
  INV_X1 U15092 ( .A(n11798), .ZN(n11802) );
  AOI22_X1 U15093 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U15094 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11800) );
  NAND2_X1 U15095 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11799) );
  NAND4_X1 U15096 ( .A1(n11802), .A2(n11801), .A3(n11800), .A4(n11799), .ZN(
        n11810) );
  AOI22_X1 U15097 ( .A1(n12460), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11733), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11808) );
  AOI22_X1 U15098 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11804), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11807) );
  AOI22_X1 U15099 ( .A1(n11731), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11806) );
  AOI22_X1 U15100 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11805) );
  NAND4_X1 U15101 ( .A1(n11808), .A2(n11807), .A3(n11806), .A4(n11805), .ZN(
        n11809) );
  XNOR2_X1 U15102 ( .A(n12765), .B(n12720), .ZN(n11812) );
  AOI21_X1 U15103 ( .B1(n13845), .B2(n12765), .A(n11759), .ZN(n11814) );
  NAND2_X1 U15104 ( .A1(n13818), .A2(n12720), .ZN(n11813) );
  NAND2_X1 U15105 ( .A1(n11844), .A2(n11843), .ZN(n11818) );
  NAND2_X1 U15106 ( .A1(n11816), .A2(n12765), .ZN(n11817) );
  NAND2_X1 U15107 ( .A1(n13523), .A2(n12714), .ZN(n11820) );
  NAND2_X1 U15108 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11819) );
  OAI211_X1 U15109 ( .C1(n11862), .C2(n12765), .A(n11820), .B(n11819), .ZN(
        n11822) );
  INV_X1 U15110 ( .A(n11822), .ZN(n11821) );
  NOR2_X1 U15111 ( .A1(n11823), .A2(n11822), .ZN(n11824) );
  NAND2_X1 U15112 ( .A1(n11828), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11906) );
  NAND2_X1 U15113 ( .A1(n12511), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11832) );
  OAI21_X1 U15114 ( .B1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n11883), .ZN(n20880) );
  OAI21_X1 U15115 ( .B1(n20880), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n11830), 
        .ZN(n11831) );
  OAI211_X1 U15116 ( .C1(n11906), .C2(n9981), .A(n11832), .B(n11831), .ZN(
        n11833) );
  INV_X1 U15117 ( .A(n11833), .ZN(n11834) );
  NAND2_X1 U15118 ( .A1(n12510), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11855) );
  NAND2_X1 U15119 ( .A1(n11835), .A2(n11855), .ZN(n13785) );
  INV_X1 U15120 ( .A(n13785), .ZN(n11854) );
  XNOR2_X2 U15121 ( .A(n11838), .B(n11837), .ZN(n14014) );
  NAND2_X1 U15122 ( .A1(n14014), .A2(n12107), .ZN(n11842) );
  AOI22_X1 U15123 ( .A1(n12511), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n11830), .ZN(n11840) );
  INV_X1 U15124 ( .A(n11906), .ZN(n11848) );
  NAND2_X1 U15125 ( .A1(n11848), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11839) );
  AND2_X1 U15126 ( .A1(n11840), .A2(n11839), .ZN(n11841) );
  NAND2_X1 U15127 ( .A1(n11842), .A2(n11841), .ZN(n13740) );
  XNOR2_X1 U15128 ( .A(n11844), .B(n11843), .ZN(n14013) );
  AOI21_X1 U15129 ( .B1(n14013), .B2(n13813), .A(n11830), .ZN(n13669) );
  INV_X1 U15130 ( .A(n11845), .ZN(n11846) );
  XNOR2_X1 U15131 ( .A(n11847), .B(n11846), .ZN(n15641) );
  NAND2_X1 U15132 ( .A1(n15641), .A2(n12107), .ZN(n11852) );
  AOI22_X1 U15133 ( .A1(n11935), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n11830), .ZN(n11850) );
  NAND2_X1 U15134 ( .A1(n11848), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11849) );
  AND2_X1 U15135 ( .A1(n11850), .A2(n11849), .ZN(n11851) );
  NAND2_X1 U15136 ( .A1(n11852), .A2(n11851), .ZN(n13670) );
  MUX2_X1 U15137 ( .A(n11907), .B(n13669), .S(n13670), .Z(n13739) );
  NAND2_X1 U15138 ( .A1(n13740), .A2(n13739), .ZN(n13738) );
  INV_X1 U15139 ( .A(n13738), .ZN(n11853) );
  NAND2_X1 U15140 ( .A1(n11854), .A2(n11853), .ZN(n11856) );
  NAND2_X1 U15141 ( .A1(n11723), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11860) );
  OAI21_X1 U15142 ( .B1(n21132), .B2(n17091), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11858) );
  INV_X1 U15143 ( .A(n21132), .ZN(n11857) );
  NOR2_X1 U15144 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n17091), .ZN(
        n14190) );
  NAND2_X1 U15145 ( .A1(n11857), .A2(n14190), .ZN(n14039) );
  NAND2_X1 U15146 ( .A1(n11858), .A2(n14039), .ZN(n14195) );
  AOI22_X1 U15147 ( .A1(n14195), .A2(n13515), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n21203), .ZN(n11859) );
  INV_X1 U15148 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11865) );
  NAND2_X1 U15149 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11864) );
  NAND2_X1 U15150 ( .A1(n12460), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11863) );
  OAI211_X1 U15151 ( .C1(n12199), .C2(n11865), .A(n11864), .B(n11863), .ZN(
        n11866) );
  INV_X1 U15152 ( .A(n11866), .ZN(n11872) );
  AOI22_X1 U15153 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11871) );
  INV_X1 U15154 ( .A(n11868), .ZN(n12321) );
  INV_X2 U15155 ( .A(n11766), .ZN(n12476) );
  AOI22_X1 U15156 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11870) );
  NAND2_X1 U15157 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11869) );
  NAND4_X1 U15158 ( .A1(n11872), .A2(n11871), .A3(n11870), .A4(n11869), .ZN(
        n11878) );
  AOI22_X1 U15159 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U15160 ( .A1(n11795), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U15161 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U15162 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11873) );
  NAND4_X1 U15163 ( .A1(n11876), .A2(n11875), .A3(n11874), .A4(n11873), .ZN(
        n11877) );
  AOI22_X1 U15164 ( .A1(n12559), .A2(n12739), .B1(n12543), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11879) );
  NAND2_X1 U15165 ( .A1(n11881), .A2(n14005), .ZN(n11882) );
  XNOR2_X1 U15166 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B(n11909), .ZN(
        n20872) );
  AOI22_X1 U15167 ( .A1(n11907), .A2(n20872), .B1(n12510), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11885) );
  NAND2_X1 U15168 ( .A1(n12511), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11884) );
  OAI211_X1 U15169 ( .C1(n11906), .C2(n15614), .A(n11885), .B(n11884), .ZN(
        n11886) );
  INV_X1 U15170 ( .A(n11886), .ZN(n11887) );
  NAND2_X1 U15171 ( .A1(n13974), .A2(n13975), .ZN(n14097) );
  INV_X1 U15172 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12404) );
  NAND2_X1 U15173 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11890) );
  NAND2_X1 U15174 ( .A1(n12455), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11889) );
  OAI211_X1 U15175 ( .C1(n12199), .C2(n12404), .A(n11890), .B(n11889), .ZN(
        n11891) );
  INV_X1 U15176 ( .A(n11891), .ZN(n11895) );
  AOI22_X1 U15177 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U15178 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11804), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11893) );
  NAND2_X1 U15179 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11892) );
  NAND4_X1 U15180 ( .A1(n11895), .A2(n11894), .A3(n11893), .A4(n11892), .ZN(
        n11901) );
  AOI22_X1 U15181 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12493), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U15182 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11898) );
  AOI22_X1 U15183 ( .A1(n11795), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11897) );
  AOI22_X1 U15184 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11896) );
  NAND4_X1 U15185 ( .A1(n11899), .A2(n11898), .A3(n11897), .A4(n11896), .ZN(
        n11900) );
  NAND2_X1 U15186 ( .A1(n12559), .A2(n12741), .ZN(n11903) );
  NAND2_X1 U15187 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11902) );
  NAND2_X1 U15188 ( .A1(n11903), .A2(n11902), .ZN(n11918) );
  NAND2_X1 U15189 ( .A1(n11830), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11905) );
  NAND2_X1 U15190 ( .A1(n12511), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11904) );
  OAI211_X1 U15191 ( .C1(n11906), .C2(n17214), .A(n11905), .B(n11904), .ZN(
        n11908) );
  NAND2_X1 U15192 ( .A1(n11908), .A2(n12503), .ZN(n11915) );
  INV_X1 U15193 ( .A(n11936), .ZN(n11937) );
  INV_X1 U15194 ( .A(n11910), .ZN(n11912) );
  INV_X1 U15195 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11911) );
  NAND2_X1 U15196 ( .A1(n11912), .A2(n11911), .ZN(n11913) );
  NAND2_X1 U15197 ( .A1(n11937), .A2(n11913), .ZN(n20864) );
  NAND2_X1 U15198 ( .A1(n20864), .A2(n12273), .ZN(n11914) );
  NAND2_X1 U15199 ( .A1(n11915), .A2(n11914), .ZN(n11916) );
  INV_X1 U15200 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12429) );
  NAND2_X1 U15201 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11920) );
  NAND2_X1 U15202 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11919) );
  OAI211_X1 U15203 ( .C1(n12199), .C2(n12429), .A(n11920), .B(n11919), .ZN(
        n11921) );
  INV_X1 U15204 ( .A(n11921), .ZN(n11925) );
  AOI22_X1 U15205 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U15206 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11923) );
  NAND2_X1 U15207 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11922) );
  NAND4_X1 U15208 ( .A1(n11925), .A2(n11924), .A3(n11923), .A4(n11922), .ZN(
        n11932) );
  AOI22_X1 U15209 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U15210 ( .A1(n11795), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11929) );
  INV_X2 U15211 ( .A(n11926), .ZN(n12486) );
  AOI22_X1 U15212 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11928) );
  AOI22_X1 U15213 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11927) );
  NAND4_X1 U15214 ( .A1(n11930), .A2(n11929), .A3(n11928), .A4(n11927), .ZN(
        n11931) );
  NAND2_X1 U15215 ( .A1(n12559), .A2(n12756), .ZN(n11934) );
  NAND2_X1 U15216 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11933) );
  INV_X1 U15217 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n14160) );
  INV_X1 U15218 ( .A(n11963), .ZN(n11939) );
  INV_X1 U15219 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20761) );
  NAND2_X1 U15220 ( .A1(n11937), .A2(n20761), .ZN(n11938) );
  NAND2_X1 U15221 ( .A1(n11939), .A2(n11938), .ZN(n20767) );
  AOI22_X1 U15222 ( .A1(n20767), .A2(n12273), .B1(n12510), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11940) );
  OAI21_X1 U15223 ( .B1(n12505), .B2(n14160), .A(n11940), .ZN(n11941) );
  INV_X1 U15224 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11945) );
  NAND2_X1 U15225 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11944) );
  NAND2_X1 U15226 ( .A1(n11795), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11943) );
  OAI211_X1 U15227 ( .C1(n12199), .C2(n11945), .A(n11944), .B(n11943), .ZN(
        n11946) );
  INV_X1 U15228 ( .A(n11946), .ZN(n11950) );
  AOI22_X1 U15229 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U15230 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11948) );
  NAND2_X1 U15231 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11947) );
  NAND4_X1 U15232 ( .A1(n11950), .A2(n11949), .A3(n11948), .A4(n11947), .ZN(
        n11956) );
  AOI22_X1 U15233 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11954) );
  AOI22_X1 U15234 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U15235 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U15236 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11951) );
  NAND4_X1 U15237 ( .A1(n11954), .A2(n11953), .A3(n11952), .A4(n11951), .ZN(
        n11955) );
  AOI22_X1 U15238 ( .A1(n12559), .A2(n12758), .B1(n12543), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11959) );
  INV_X1 U15239 ( .A(n11959), .ZN(n11957) );
  NAND2_X1 U15240 ( .A1(n11960), .A2(n11959), .ZN(n11961) );
  INV_X1 U15241 ( .A(n12755), .ZN(n11962) );
  NAND2_X1 U15242 ( .A1(n11962), .A2(n12107), .ZN(n11968) );
  INV_X1 U15243 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11965) );
  OAI21_X1 U15244 ( .B1(n11963), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n11971), .ZN(n20754) );
  AOI22_X1 U15245 ( .A1(n20754), .A2(n12273), .B1(n12510), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11964) );
  OAI21_X1 U15246 ( .B1(n12505), .B2(n11965), .A(n11964), .ZN(n11966) );
  INV_X1 U15247 ( .A(n14171), .ZN(n11994) );
  NAND2_X1 U15248 ( .A1(n12559), .A2(n12765), .ZN(n11969) );
  OAI21_X1 U15249 ( .B1(n12478), .B2(n12542), .A(n11969), .ZN(n11970) );
  INV_X1 U15250 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11974) );
  OAI21_X1 U15251 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n11972), .A(
        n12008), .ZN(n20739) );
  AOI22_X1 U15252 ( .A1(n12273), .A2(n20739), .B1(n12510), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11973) );
  OAI21_X1 U15253 ( .B1(n12505), .B2(n11974), .A(n11973), .ZN(n11975) );
  NAND2_X1 U15254 ( .A1(n12511), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11992) );
  XOR2_X1 U15255 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n12008), .Z(n15387) );
  AOI22_X1 U15256 ( .A1(n12510), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n12273), .B2(n15387), .ZN(n11991) );
  AOI22_X1 U15257 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11979) );
  AOI22_X1 U15258 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11978) );
  INV_X2 U15259 ( .A(n12452), .ZN(n12481) );
  AOI22_X1 U15260 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U15261 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11976) );
  NAND4_X1 U15262 ( .A1(n11979), .A2(n11978), .A3(n11977), .A4(n11976), .ZN(
        n11988) );
  AOI22_X1 U15263 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11982) );
  NAND2_X1 U15264 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11981) );
  AOI22_X1 U15265 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11980) );
  NAND3_X1 U15266 ( .A1(n11982), .A2(n11981), .A3(n11980), .ZN(n11987) );
  INV_X1 U15267 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11985) );
  NAND2_X1 U15268 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11984) );
  NAND2_X1 U15269 ( .A1(n11795), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11983) );
  OAI211_X1 U15270 ( .C1(n12479), .C2(n11985), .A(n11984), .B(n11983), .ZN(
        n11986) );
  NOR3_X1 U15271 ( .A1(n11988), .A2(n11987), .A3(n11986), .ZN(n11989) );
  OR2_X1 U15272 ( .A1(n12172), .A2(n11989), .ZN(n11990) );
  AOI22_X1 U15273 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U15274 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11997) );
  AOI22_X1 U15275 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11996) );
  AOI22_X1 U15276 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11995) );
  NAND4_X1 U15277 ( .A1(n11998), .A2(n11997), .A3(n11996), .A4(n11995), .ZN(
        n12007) );
  INV_X1 U15278 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12330) );
  NAND2_X1 U15279 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12000) );
  NAND2_X1 U15280 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11999) );
  OAI211_X1 U15281 ( .C1(n12199), .C2(n12330), .A(n12000), .B(n11999), .ZN(
        n12001) );
  INV_X1 U15282 ( .A(n12001), .ZN(n12005) );
  AOI22_X1 U15283 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U15284 ( .A1(n11795), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12003) );
  NAND2_X1 U15285 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12002) );
  NAND4_X1 U15286 ( .A1(n12005), .A2(n12004), .A3(n12003), .A4(n12002), .ZN(
        n12006) );
  OAI21_X1 U15287 ( .B1(n12007), .B2(n12006), .A(n12107), .ZN(n12012) );
  INV_X1 U15288 ( .A(n12014), .ZN(n12009) );
  XNOR2_X1 U15289 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n12009), .ZN(
        n15377) );
  AOI22_X1 U15290 ( .A1(n11907), .A2(n15377), .B1(n12510), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12011) );
  NAND2_X1 U15291 ( .A1(n12511), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12010) );
  XNOR2_X1 U15292 ( .A(n12037), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17156) );
  NAND2_X1 U15293 ( .A1(n17156), .A2(n12273), .ZN(n12033) );
  AOI22_X1 U15294 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11804), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U15295 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U15296 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U15297 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12015) );
  NAND4_X1 U15298 ( .A1(n12018), .A2(n12017), .A3(n12016), .A4(n12015), .ZN(
        n12028) );
  INV_X1 U15299 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12021) );
  NAND2_X1 U15300 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12020) );
  NAND2_X1 U15301 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n12019) );
  OAI211_X1 U15302 ( .C1(n12199), .C2(n12021), .A(n12020), .B(n12019), .ZN(
        n12022) );
  INV_X1 U15303 ( .A(n12022), .ZN(n12026) );
  AOI22_X1 U15304 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12025) );
  AOI22_X1 U15305 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12024) );
  NAND2_X1 U15306 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12023) );
  NAND4_X1 U15307 ( .A1(n12026), .A2(n12025), .A3(n12024), .A4(n12023), .ZN(
        n12027) );
  OAI21_X1 U15308 ( .B1(n12028), .B2(n12027), .A(n12107), .ZN(n12031) );
  NAND2_X1 U15309 ( .A1(n12511), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12030) );
  NAND2_X1 U15310 ( .A1(n12510), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12029) );
  AND3_X1 U15311 ( .A1(n12031), .A2(n12030), .A3(n12029), .ZN(n12032) );
  NAND2_X1 U15312 ( .A1(n12033), .A2(n12032), .ZN(n14280) );
  NAND2_X1 U15313 ( .A1(n12037), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12035) );
  INV_X1 U15314 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12034) );
  NAND2_X1 U15315 ( .A1(n12035), .A2(n12034), .ZN(n12038) );
  NAND2_X1 U15316 ( .A1(n12038), .A2(n12073), .ZN(n15359) );
  NAND2_X1 U15317 ( .A1(n15359), .A2(n12273), .ZN(n12040) );
  AOI22_X1 U15318 ( .A1(n12511), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12510), .ZN(n12039) );
  NAND2_X1 U15319 ( .A1(n12040), .A2(n12039), .ZN(n14954) );
  AOI22_X1 U15320 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12044) );
  AOI22_X1 U15321 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12043) );
  AOI22_X1 U15322 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U15323 ( .A1(n11795), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12041) );
  AND4_X1 U15324 ( .A1(n12044), .A2(n12043), .A3(n12042), .A4(n12041), .ZN(
        n12052) );
  AOI22_X1 U15325 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12051) );
  NAND2_X1 U15326 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12048) );
  AOI22_X1 U15327 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12047) );
  NAND2_X1 U15328 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12046) );
  NAND2_X1 U15329 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12045) );
  AND4_X1 U15330 ( .A1(n12048), .A2(n12047), .A3(n12046), .A4(n12045), .ZN(
        n12050) );
  NAND2_X1 U15331 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12049) );
  NAND4_X1 U15332 ( .A1(n12052), .A2(n12051), .A3(n12050), .A4(n12049), .ZN(
        n12053) );
  NAND2_X1 U15333 ( .A1(n14954), .A2(n14953), .ZN(n12054) );
  NAND2_X1 U15334 ( .A1(n12094), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12055) );
  INV_X1 U15335 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14964) );
  XNOR2_X1 U15336 ( .A(n12055), .B(n14964), .ZN(n15336) );
  AOI22_X1 U15337 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12059) );
  AOI22_X1 U15338 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U15339 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U15340 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12056) );
  NAND4_X1 U15341 ( .A1(n12059), .A2(n12058), .A3(n12057), .A4(n12056), .ZN(
        n12068) );
  INV_X1 U15342 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12244) );
  NAND2_X1 U15343 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12061) );
  NAND2_X1 U15344 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12060) );
  OAI211_X1 U15345 ( .C1(n12199), .C2(n12244), .A(n12061), .B(n12060), .ZN(
        n12062) );
  INV_X1 U15346 ( .A(n12062), .ZN(n12066) );
  AOI22_X1 U15347 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U15348 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12064) );
  NAND2_X1 U15349 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12063) );
  NAND4_X1 U15350 ( .A1(n12066), .A2(n12065), .A3(n12064), .A4(n12063), .ZN(
        n12067) );
  OAI21_X1 U15351 ( .B1(n12068), .B2(n12067), .A(n12107), .ZN(n12071) );
  NAND2_X1 U15352 ( .A1(n12511), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12070) );
  NAND2_X1 U15353 ( .A1(n12510), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12069) );
  NAND3_X1 U15354 ( .A1(n12071), .A2(n12070), .A3(n12069), .ZN(n12072) );
  AOI21_X1 U15355 ( .B1(n15336), .B2(n11907), .A(n12072), .ZN(n14957) );
  INV_X1 U15356 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n14980) );
  XNOR2_X1 U15357 ( .A(n12073), .B(n14980), .ZN(n15349) );
  NAND2_X1 U15358 ( .A1(n15349), .A2(n12273), .ZN(n12090) );
  INV_X1 U15359 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n15158) );
  AOI22_X1 U15360 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12430), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12077) );
  AOI22_X1 U15361 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12076) );
  AOI22_X1 U15362 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12075) );
  AOI22_X1 U15363 ( .A1(n11795), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12074) );
  AND4_X1 U15364 ( .A1(n12077), .A2(n12076), .A3(n12075), .A4(n12074), .ZN(
        n12084) );
  AOI22_X1 U15365 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U15366 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11804), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U15367 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12079) );
  NAND2_X1 U15368 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12078) );
  AND3_X1 U15369 ( .A1(n12080), .A2(n12079), .A3(n12078), .ZN(n12082) );
  NAND2_X1 U15370 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12081) );
  NAND4_X1 U15371 ( .A1(n12084), .A2(n12083), .A3(n12082), .A4(n12081), .ZN(
        n12085) );
  NAND2_X1 U15372 ( .A1(n12107), .A2(n12085), .ZN(n12087) );
  NAND2_X1 U15373 ( .A1(n12510), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12086) );
  OAI211_X1 U15374 ( .C1(n12505), .C2(n15158), .A(n12087), .B(n12086), .ZN(
        n12088) );
  INV_X1 U15375 ( .A(n12088), .ZN(n12089) );
  NAND2_X1 U15376 ( .A1(n12090), .A2(n12089), .ZN(n14972) );
  OAI21_X1 U15377 ( .B1(n14953), .B2(n14954), .A(n14972), .ZN(n12091) );
  NOR2_X1 U15378 ( .A1(n14957), .A2(n12091), .ZN(n12092) );
  INV_X1 U15379 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12155) );
  XNOR2_X1 U15380 ( .A(n12156), .B(n12155), .ZN(n15326) );
  AOI22_X1 U15381 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U15382 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U15383 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15384 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12095) );
  NAND4_X1 U15385 ( .A1(n12098), .A2(n12097), .A3(n12096), .A4(n12095), .ZN(
        n12109) );
  INV_X1 U15386 ( .A(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12101) );
  NAND2_X1 U15387 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12100) );
  NAND2_X1 U15388 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12099) );
  OAI211_X1 U15389 ( .C1(n12199), .C2(n12101), .A(n12100), .B(n12099), .ZN(
        n12102) );
  INV_X1 U15390 ( .A(n12102), .ZN(n12106) );
  AOI22_X1 U15391 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U15392 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12104) );
  NAND2_X1 U15393 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12103) );
  NAND4_X1 U15394 ( .A1(n12106), .A2(n12105), .A3(n12104), .A4(n12103), .ZN(
        n12108) );
  OAI21_X1 U15395 ( .B1(n12109), .B2(n12108), .A(n12107), .ZN(n12112) );
  NAND2_X1 U15396 ( .A1(n12511), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12111) );
  NAND2_X1 U15397 ( .A1(n12510), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12110) );
  NAND3_X1 U15398 ( .A1(n12112), .A2(n12111), .A3(n12110), .ZN(n12113) );
  AOI21_X1 U15399 ( .B1(n15326), .B2(n12273), .A(n12113), .ZN(n14940) );
  INV_X1 U15400 ( .A(n12116), .ZN(n12118) );
  INV_X1 U15401 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12117) );
  NAND2_X1 U15402 ( .A1(n12118), .A2(n12117), .ZN(n12119) );
  NAND2_X1 U15403 ( .A1(n12234), .A2(n12119), .ZN(n15267) );
  OR2_X1 U15404 ( .A1(n15267), .A2(n12503), .ZN(n12140) );
  INV_X1 U15405 ( .A(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12123) );
  NAND2_X1 U15406 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12122) );
  NAND2_X1 U15407 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12121) );
  OAI211_X1 U15408 ( .C1(n12199), .C2(n12123), .A(n12122), .B(n12121), .ZN(
        n12124) );
  INV_X1 U15409 ( .A(n12124), .ZN(n12128) );
  AOI22_X1 U15410 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U15411 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12126) );
  NAND2_X1 U15412 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12125) );
  NAND4_X1 U15413 ( .A1(n12128), .A2(n12127), .A3(n12126), .A4(n12125), .ZN(
        n12134) );
  AOI22_X1 U15414 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12481), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12132) );
  AOI22_X1 U15415 ( .A1(n11761), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12352), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U15416 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12130) );
  AOI22_X1 U15417 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12129) );
  NAND4_X1 U15418 ( .A1(n12132), .A2(n12131), .A3(n12130), .A4(n12129), .ZN(
        n12133) );
  NOR2_X1 U15419 ( .A1(n12134), .A2(n12133), .ZN(n12138) );
  NAND2_X1 U15420 ( .A1(n11830), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12135) );
  NAND2_X1 U15421 ( .A1(n12503), .A2(n12135), .ZN(n12136) );
  AOI21_X1 U15422 ( .B1(n12511), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12136), .ZN(
        n12137) );
  OAI21_X1 U15423 ( .B1(n12471), .B2(n12138), .A(n12137), .ZN(n12139) );
  XNOR2_X1 U15424 ( .A(n12195), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15303) );
  NAND2_X1 U15425 ( .A1(n12471), .A2(n12503), .ZN(n12268) );
  AOI22_X1 U15426 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11804), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12144) );
  AOI22_X1 U15427 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12143) );
  AOI22_X1 U15428 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12142) );
  AOI22_X1 U15429 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12141) );
  AND4_X1 U15430 ( .A1(n12144), .A2(n12143), .A3(n12142), .A4(n12141), .ZN(
        n12151) );
  AOI22_X1 U15431 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12148) );
  AOI21_X1 U15432 ( .B1(n12485), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n11907), .ZN(n12147) );
  AOI22_X1 U15433 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12146) );
  NAND2_X1 U15434 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12145) );
  AND4_X1 U15435 ( .A1(n12148), .A2(n12147), .A3(n12146), .A4(n12145), .ZN(
        n12150) );
  AOI22_X1 U15436 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12149) );
  NAND3_X1 U15437 ( .A1(n12151), .A2(n12150), .A3(n12149), .ZN(n12153) );
  INV_X1 U15438 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n15142) );
  OAI22_X1 U15439 ( .A1(n12505), .A2(n15142), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15300), .ZN(n12152) );
  AOI21_X1 U15440 ( .B1(n12268), .B2(n12153), .A(n12152), .ZN(n12154) );
  AOI21_X1 U15441 ( .B1(n15303), .B2(n11907), .A(n12154), .ZN(n14916) );
  INV_X1 U15442 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n21369) );
  OAI21_X1 U15443 ( .B1(n12156), .B2(n12155), .A(n21369), .ZN(n12157) );
  NAND2_X1 U15444 ( .A1(n12157), .A2(n12195), .ZN(n15315) );
  NAND2_X1 U15445 ( .A1(n15315), .A2(n12273), .ZN(n12177) );
  INV_X1 U15446 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20803) );
  INV_X1 U15447 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12492) );
  NAND2_X1 U15448 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12159) );
  NAND2_X1 U15449 ( .A1(n12455), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12158) );
  OAI211_X1 U15450 ( .C1(n12199), .C2(n12492), .A(n12159), .B(n12158), .ZN(
        n12160) );
  INV_X1 U15451 ( .A(n12160), .ZN(n12164) );
  AOI22_X1 U15452 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12163) );
  AOI22_X1 U15453 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12162) );
  NAND2_X1 U15454 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12161) );
  NAND4_X1 U15455 ( .A1(n12164), .A2(n12163), .A3(n12162), .A4(n12161), .ZN(
        n12170) );
  AOI22_X1 U15456 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15457 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U15458 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12166) );
  AOI22_X1 U15459 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12165) );
  NAND4_X1 U15460 ( .A1(n12168), .A2(n12167), .A3(n12166), .A4(n12165), .ZN(
        n12169) );
  NOR2_X1 U15461 ( .A1(n12170), .A2(n12169), .ZN(n12171) );
  OR2_X1 U15462 ( .A1(n12172), .A2(n12171), .ZN(n12174) );
  NAND2_X1 U15463 ( .A1(n12510), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12173) );
  OAI211_X1 U15464 ( .C1(n12505), .C2(n20803), .A(n12174), .B(n12173), .ZN(
        n12175) );
  INV_X1 U15465 ( .A(n12175), .ZN(n12176) );
  NAND2_X1 U15466 ( .A1(n12177), .A2(n12176), .ZN(n14930) );
  NAND3_X1 U15467 ( .A1(n14876), .A2(n14916), .A3(n14930), .ZN(n12215) );
  XNOR2_X1 U15468 ( .A(n12178), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15276) );
  NAND2_X1 U15469 ( .A1(n15276), .A2(n12273), .ZN(n12194) );
  AOI22_X1 U15470 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11804), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12182) );
  AOI22_X1 U15471 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12481), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15472 ( .A1(n11761), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12352), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15473 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12179) );
  NAND4_X1 U15474 ( .A1(n12182), .A2(n12181), .A3(n12180), .A4(n12179), .ZN(
        n12190) );
  AOI22_X1 U15475 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12188) );
  NAND2_X1 U15476 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12184) );
  AOI21_X1 U15477 ( .B1(n11867), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n11907), .ZN(n12183) );
  AND2_X1 U15478 ( .A1(n12184), .A2(n12183), .ZN(n12187) );
  AOI22_X1 U15479 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12485), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U15480 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12185) );
  NAND4_X1 U15481 ( .A1(n12188), .A2(n12187), .A3(n12186), .A4(n12185), .ZN(
        n12189) );
  OAI21_X1 U15482 ( .B1(n12190), .B2(n12189), .A(n12268), .ZN(n12192) );
  AOI22_X1 U15483 ( .A1(n12511), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n11830), .ZN(n12191) );
  NAND2_X1 U15484 ( .A1(n12192), .A2(n12191), .ZN(n12193) );
  NAND2_X1 U15485 ( .A1(n12194), .A2(n12193), .ZN(n14875) );
  OR2_X1 U15486 ( .A1(n12195), .A2(n15300), .ZN(n12196) );
  XNOR2_X1 U15487 ( .A(n12196), .B(n14907), .ZN(n15291) );
  INV_X1 U15488 ( .A(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12318) );
  NAND2_X1 U15489 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12198) );
  NAND2_X1 U15490 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12197) );
  OAI211_X1 U15491 ( .C1(n12199), .C2(n12318), .A(n12198), .B(n12197), .ZN(
        n12200) );
  INV_X1 U15492 ( .A(n12200), .ZN(n12204) );
  AOI22_X1 U15493 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15494 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12202) );
  NAND2_X1 U15495 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12201) );
  NAND4_X1 U15496 ( .A1(n12204), .A2(n12203), .A3(n12202), .A4(n12201), .ZN(
        n12210) );
  AOI22_X1 U15497 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15498 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15499 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15500 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12205) );
  NAND4_X1 U15501 ( .A1(n12208), .A2(n12207), .A3(n12206), .A4(n12205), .ZN(
        n12209) );
  NOR2_X1 U15502 ( .A1(n12210), .A2(n12209), .ZN(n12212) );
  AOI22_X1 U15503 ( .A1(n12511), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n12510), .ZN(n12211) );
  OAI21_X1 U15504 ( .B1(n12471), .B2(n12212), .A(n12211), .ZN(n12213) );
  XNOR2_X1 U15505 ( .A(n12234), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15259) );
  INV_X1 U15506 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15257) );
  AOI21_X1 U15507 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15257), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12217) );
  AOI21_X1 U15508 ( .B1(n12511), .B2(P1_EAX_REG_20__SCAN_IN), .A(n12217), .ZN(
        n12233) );
  AOI22_X1 U15509 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U15510 ( .A1(n11795), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U15511 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15512 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12219) );
  NAND4_X1 U15513 ( .A1(n12222), .A2(n12221), .A3(n12220), .A4(n12219), .ZN(
        n12231) );
  INV_X1 U15514 ( .A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12229) );
  INV_X1 U15515 ( .A(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12396) );
  INV_X1 U15516 ( .A(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12223) );
  OAI22_X1 U15517 ( .A1(n12351), .A2(n12396), .B1(n12317), .B2(n12223), .ZN(
        n12226) );
  INV_X1 U15518 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12224) );
  INV_X1 U15519 ( .A(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12406) );
  OAI22_X1 U15520 ( .A1(n12321), .A2(n12224), .B1(n11766), .B2(n12406), .ZN(
        n12225) );
  AOI211_X1 U15521 ( .C1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .C2(n12487), .A(
        n12226), .B(n12225), .ZN(n12228) );
  AOI22_X1 U15522 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12227) );
  OAI211_X1 U15523 ( .C1(n12199), .C2(n12229), .A(n12228), .B(n12227), .ZN(
        n12230) );
  OAI21_X1 U15524 ( .B1(n12231), .B2(n12230), .A(n12507), .ZN(n12232) );
  AOI22_X1 U15525 ( .A1(n15259), .A2(n12273), .B1(n12233), .B2(n12232), .ZN(
        n14862) );
  INV_X1 U15526 ( .A(n12236), .ZN(n12238) );
  INV_X1 U15527 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12237) );
  NAND2_X1 U15528 ( .A1(n12238), .A2(n12237), .ZN(n12239) );
  NAND2_X1 U15529 ( .A1(n12274), .A2(n12239), .ZN(n15249) );
  INV_X1 U15530 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n15116) );
  AOI22_X1 U15531 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12243) );
  AOI22_X1 U15532 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12242) );
  AOI22_X1 U15533 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U15534 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12240) );
  NAND4_X1 U15535 ( .A1(n12243), .A2(n12242), .A3(n12241), .A4(n12240), .ZN(
        n12254) );
  INV_X1 U15536 ( .A(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12252) );
  INV_X1 U15537 ( .A(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14095) );
  OAI22_X1 U15538 ( .A1(n12351), .A2(n12244), .B1(n12317), .B2(n14095), .ZN(
        n12249) );
  INV_X1 U15539 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12247) );
  INV_X1 U15540 ( .A(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12245) );
  OAI22_X1 U15541 ( .A1(n12321), .A2(n12247), .B1(n12246), .B2(n12245), .ZN(
        n12248) );
  AOI211_X1 U15542 ( .C1(n12487), .C2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n12249), .B(n12248), .ZN(n12251) );
  AOI22_X1 U15543 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12250) );
  OAI211_X1 U15544 ( .C1(n12199), .C2(n12252), .A(n12251), .B(n12250), .ZN(
        n12253) );
  OAI21_X1 U15545 ( .B1(n12254), .B2(n12253), .A(n12507), .ZN(n12256) );
  AOI21_X1 U15546 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n11830), .A(
        n12273), .ZN(n12255) );
  OAI211_X1 U15547 ( .C1(n12505), .C2(n15116), .A(n12256), .B(n12255), .ZN(
        n12257) );
  XNOR2_X1 U15548 ( .A(n12274), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15236) );
  AOI22_X1 U15549 ( .A1(n12511), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n11830), .ZN(n12272) );
  AOI22_X1 U15550 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11804), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12261) );
  AOI22_X1 U15551 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12260) );
  AOI22_X1 U15552 ( .A1(n12302), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12259) );
  AOI22_X1 U15553 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12258) );
  NAND4_X1 U15554 ( .A1(n12261), .A2(n12260), .A3(n12259), .A4(n12258), .ZN(
        n12270) );
  AOI22_X1 U15555 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12267) );
  AOI21_X1 U15556 ( .B1(n12485), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n11907), .ZN(n12263) );
  NAND2_X1 U15557 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12262) );
  AND2_X1 U15558 ( .A1(n12263), .A2(n12262), .ZN(n12266) );
  AOI22_X1 U15559 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15560 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12264) );
  NAND4_X1 U15561 ( .A1(n12267), .A2(n12266), .A3(n12265), .A4(n12264), .ZN(
        n12269) );
  OAI21_X1 U15562 ( .B1(n12270), .B2(n12269), .A(n12268), .ZN(n12271) );
  AOI22_X1 U15563 ( .A1(n15236), .A2(n12273), .B1(n12272), .B2(n12271), .ZN(
        n14841) );
  INV_X1 U15564 ( .A(n12276), .ZN(n12278) );
  INV_X1 U15565 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12277) );
  NAND2_X1 U15566 ( .A1(n12278), .A2(n12277), .ZN(n12279) );
  NAND2_X1 U15567 ( .A1(n12342), .A2(n12279), .ZN(n15230) );
  INV_X1 U15568 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12282) );
  AOI22_X1 U15569 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12281) );
  NAND2_X1 U15570 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12280) );
  OAI211_X1 U15571 ( .C1(n12282), .C2(n12199), .A(n12281), .B(n12280), .ZN(
        n12283) );
  INV_X1 U15572 ( .A(n12283), .ZN(n12286) );
  AOI22_X1 U15573 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12285) );
  AOI22_X1 U15574 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12284) );
  NAND3_X1 U15575 ( .A1(n12286), .A2(n12285), .A3(n12284), .ZN(n12294) );
  INV_X1 U15576 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12494) );
  OAI22_X1 U15577 ( .A1(n12452), .A2(n12494), .B1(n12287), .B2(n12478), .ZN(
        n12288) );
  AOI21_X1 U15578 ( .B1(n12493), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n12288), .ZN(n12292) );
  AOI22_X1 U15579 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U15580 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12290) );
  NAND2_X1 U15581 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12289) );
  NAND4_X1 U15582 ( .A1(n12292), .A2(n12291), .A3(n12290), .A4(n12289), .ZN(
        n12293) );
  NOR2_X1 U15583 ( .A1(n12294), .A2(n12293), .ZN(n12336) );
  AOI22_X1 U15584 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12299) );
  AOI22_X1 U15585 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15586 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U15587 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12296) );
  NAND4_X1 U15588 ( .A1(n12299), .A2(n12298), .A3(n12297), .A4(n12296), .ZN(
        n12311) );
  INV_X1 U15589 ( .A(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12309) );
  INV_X1 U15590 ( .A(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12301) );
  INV_X1 U15591 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12300) );
  OAI22_X1 U15592 ( .A1(n12321), .A2(n12301), .B1(n11766), .B2(n12300), .ZN(
        n12306) );
  INV_X1 U15593 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12304) );
  INV_X1 U15594 ( .A(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12303) );
  OAI22_X1 U15595 ( .A1(n12495), .A2(n12304), .B1(n11926), .B2(n12303), .ZN(
        n12305) );
  AOI211_X1 U15596 ( .C1(n12487), .C2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n12306), .B(n12305), .ZN(n12308) );
  AOI22_X1 U15597 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11795), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12307) );
  OAI211_X1 U15598 ( .C1(n12199), .C2(n12309), .A(n12308), .B(n12307), .ZN(
        n12310) );
  NOR2_X1 U15599 ( .A1(n12311), .A2(n12310), .ZN(n12337) );
  XNOR2_X1 U15600 ( .A(n12336), .B(n12337), .ZN(n12314) );
  AOI21_X1 U15601 ( .B1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n11830), .A(
        n12273), .ZN(n12313) );
  NAND2_X1 U15602 ( .A1(n12511), .A2(P1_EAX_REG_23__SCAN_IN), .ZN(n12312) );
  OAI211_X1 U15603 ( .C1(n12314), .C2(n12471), .A(n12313), .B(n12312), .ZN(
        n12315) );
  XNOR2_X1 U15604 ( .A(n12342), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15225) );
  INV_X1 U15605 ( .A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12326) );
  INV_X1 U15606 ( .A(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12316) );
  OAI22_X1 U15607 ( .A1(n12351), .A2(n12318), .B1(n12317), .B2(n12316), .ZN(
        n12323) );
  INV_X1 U15608 ( .A(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12320) );
  INV_X1 U15609 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12319) );
  OAI22_X1 U15610 ( .A1(n12321), .A2(n12320), .B1(n11766), .B2(n12319), .ZN(
        n12322) );
  AOI211_X1 U15611 ( .C1(n12487), .C2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n12323), .B(n12322), .ZN(n12325) );
  AOI22_X1 U15612 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12324) );
  OAI211_X1 U15613 ( .C1(n12199), .C2(n12326), .A(n12325), .B(n12324), .ZN(
        n12335) );
  AOI22_X1 U15614 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12328) );
  AOI22_X1 U15615 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12327) );
  NAND2_X1 U15616 ( .A1(n12328), .A2(n12327), .ZN(n12334) );
  INV_X1 U15617 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12329) );
  OAI22_X1 U15618 ( .A1(n12287), .A2(n12330), .B1(n12495), .B2(n12329), .ZN(
        n12333) );
  INV_X1 U15619 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12331) );
  OAI22_X1 U15620 ( .A1(n12490), .A2(n12331), .B1(n12479), .B2(n11764), .ZN(
        n12332) );
  NOR2_X1 U15621 ( .A1(n12337), .A2(n12336), .ZN(n12363) );
  XOR2_X1 U15622 ( .A(n12362), .B(n12363), .Z(n12340) );
  INV_X1 U15623 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n15102) );
  INV_X1 U15624 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20709) );
  NOR2_X1 U15625 ( .A1(n20709), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12338) );
  OAI22_X1 U15626 ( .A1(n12505), .A2(n15102), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12338), .ZN(n12339) );
  AOI21_X1 U15627 ( .B1(n12340), .B2(n12507), .A(n12339), .ZN(n12341) );
  AOI21_X1 U15628 ( .B1(n15225), .B2(n12273), .A(n12341), .ZN(n14816) );
  INV_X1 U15629 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15221) );
  INV_X1 U15630 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12343) );
  NAND2_X1 U15631 ( .A1(n12344), .A2(n12343), .ZN(n12345) );
  NAND2_X1 U15632 ( .A1(n12390), .A2(n12345), .ZN(n15214) );
  AOI22_X1 U15633 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11804), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12349) );
  AOI22_X1 U15634 ( .A1(n11795), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12348) );
  AOI22_X1 U15635 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U15636 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12346) );
  NAND4_X1 U15637 ( .A1(n12349), .A2(n12348), .A3(n12347), .A4(n12346), .ZN(
        n12361) );
  INV_X1 U15638 ( .A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12359) );
  INV_X1 U15639 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13843) );
  INV_X1 U15640 ( .A(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12350) );
  OAI22_X1 U15641 ( .A1(n12246), .A2(n13843), .B1(n12351), .B2(n12350), .ZN(
        n12356) );
  INV_X1 U15642 ( .A(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12354) );
  INV_X1 U15643 ( .A(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12353) );
  OAI22_X1 U15644 ( .A1(n12452), .A2(n12354), .B1(n12495), .B2(n12353), .ZN(
        n12355) );
  AOI211_X1 U15645 ( .C1(n12487), .C2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n12356), .B(n12355), .ZN(n12358) );
  AOI22_X1 U15646 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12430), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12357) );
  OAI211_X1 U15647 ( .C1(n12199), .C2(n12359), .A(n12358), .B(n12357), .ZN(
        n12360) );
  NOR2_X1 U15648 ( .A1(n12361), .A2(n12360), .ZN(n12369) );
  NAND2_X1 U15649 ( .A1(n12363), .A2(n12362), .ZN(n12368) );
  XNOR2_X1 U15650 ( .A(n12369), .B(n12368), .ZN(n12366) );
  AOI21_X1 U15651 ( .B1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n11830), .A(
        n12273), .ZN(n12365) );
  NAND2_X1 U15652 ( .A1(n12511), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n12364) );
  OAI211_X1 U15653 ( .C1(n12366), .C2(n12471), .A(n12365), .B(n12364), .ZN(
        n12367) );
  XNOR2_X1 U15654 ( .A(n12390), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15199) );
  NOR2_X1 U15655 ( .A1(n12369), .A2(n12368), .ZN(n12414) );
  INV_X1 U15656 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12372) );
  NAND2_X1 U15657 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12371) );
  NAND2_X1 U15658 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12370) );
  OAI211_X1 U15659 ( .C1(n12199), .C2(n12372), .A(n12371), .B(n12370), .ZN(
        n12373) );
  INV_X1 U15660 ( .A(n12373), .ZN(n12377) );
  AOI22_X1 U15661 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15662 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12375) );
  NAND2_X1 U15663 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12374) );
  NAND4_X1 U15664 ( .A1(n12377), .A2(n12376), .A3(n12375), .A4(n12374), .ZN(
        n12383) );
  AOI22_X1 U15665 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U15666 ( .A1(n11795), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12380) );
  AOI22_X1 U15667 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12379) );
  AOI22_X1 U15668 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12378) );
  NAND4_X1 U15669 ( .A1(n12381), .A2(n12380), .A3(n12379), .A4(n12378), .ZN(
        n12382) );
  INV_X1 U15670 ( .A(n12413), .ZN(n12384) );
  XNOR2_X1 U15671 ( .A(n12414), .B(n12384), .ZN(n12388) );
  INV_X1 U15672 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n12386) );
  NAND2_X1 U15673 ( .A1(n11830), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12385) );
  OAI211_X1 U15674 ( .C1(n12505), .C2(n12386), .A(n12503), .B(n12385), .ZN(
        n12387) );
  AOI21_X1 U15675 ( .B1(n12388), .B2(n12507), .A(n12387), .ZN(n12389) );
  INV_X1 U15676 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15201) );
  NOR2_X2 U15677 ( .A1(n12390), .A2(n15201), .ZN(n12391) );
  INV_X1 U15678 ( .A(n12391), .ZN(n12393) );
  INV_X1 U15679 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12392) );
  NAND2_X1 U15680 ( .A1(n12393), .A2(n12392), .ZN(n12394) );
  NAND2_X1 U15681 ( .A1(n12441), .A2(n12394), .ZN(n15192) );
  AOI22_X1 U15682 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12485), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12395) );
  OAI21_X1 U15683 ( .B1(n12396), .B2(n12287), .A(n12395), .ZN(n12397) );
  AOI21_X1 U15684 ( .B1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B2(n12487), .A(
        n12397), .ZN(n12400) );
  AOI22_X1 U15685 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15686 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12430), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12398) );
  NAND3_X1 U15687 ( .A1(n12400), .A2(n12399), .A3(n12398), .ZN(n12412) );
  INV_X1 U15688 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13892) );
  AOI22_X1 U15689 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12402) );
  NAND2_X1 U15690 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12401) );
  OAI211_X1 U15691 ( .C1(n11760), .C2(n13892), .A(n12402), .B(n12401), .ZN(
        n12410) );
  INV_X1 U15692 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13852) );
  OAI22_X1 U15693 ( .A1(n12246), .A2(n13852), .B1(n12479), .B2(n12404), .ZN(
        n12409) );
  INV_X1 U15694 ( .A(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12405) );
  OAI22_X1 U15695 ( .A1(n12407), .A2(n12406), .B1(n12495), .B2(n12405), .ZN(
        n12408) );
  OR3_X1 U15696 ( .A1(n12410), .A2(n12409), .A3(n12408), .ZN(n12411) );
  NOR2_X1 U15697 ( .A1(n12412), .A2(n12411), .ZN(n12420) );
  NAND2_X1 U15698 ( .A1(n12414), .A2(n12413), .ZN(n12419) );
  XNOR2_X1 U15699 ( .A(n12420), .B(n12419), .ZN(n12417) );
  AOI21_X1 U15700 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n11830), .A(
        n12273), .ZN(n12416) );
  NAND2_X1 U15701 ( .A1(n11935), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n12415) );
  OAI211_X1 U15702 ( .C1(n12417), .C2(n12471), .A(n12416), .B(n12415), .ZN(
        n12418) );
  XNOR2_X1 U15703 ( .A(n12441), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15187) );
  INV_X1 U15704 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15184) );
  OAI21_X1 U15705 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15184), .A(n12503), 
        .ZN(n12439) );
  NOR2_X1 U15706 ( .A1(n12420), .A2(n12419), .ZN(n12468) );
  INV_X1 U15707 ( .A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12423) );
  NAND2_X1 U15708 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12422) );
  NAND2_X1 U15709 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12421) );
  OAI211_X1 U15710 ( .C1(n12199), .C2(n12423), .A(n12422), .B(n12421), .ZN(
        n12424) );
  INV_X1 U15711 ( .A(n12424), .ZN(n12428) );
  AOI22_X1 U15712 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12427) );
  AOI22_X1 U15713 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12426) );
  NAND2_X1 U15714 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12425) );
  NAND4_X1 U15715 ( .A1(n12428), .A2(n12427), .A3(n12426), .A4(n12425), .ZN(
        n12436) );
  AOI22_X1 U15716 ( .A1(n12447), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12434) );
  AOI22_X1 U15717 ( .A1(n11795), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12302), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12433) );
  AOI22_X1 U15718 ( .A1(n12481), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U15719 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12403), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12431) );
  NAND4_X1 U15720 ( .A1(n12434), .A2(n12433), .A3(n12432), .A4(n12431), .ZN(
        n12435) );
  OR2_X1 U15721 ( .A1(n12436), .A2(n12435), .ZN(n12467) );
  XNOR2_X1 U15722 ( .A(n12468), .B(n12467), .ZN(n12437) );
  NOR2_X1 U15723 ( .A1(n12437), .A2(n12471), .ZN(n12438) );
  AOI211_X1 U15724 ( .C1(n12511), .C2(P1_EAX_REG_28__SCAN_IN), .A(n12439), .B(
        n12438), .ZN(n12440) );
  INV_X1 U15725 ( .A(n12441), .ZN(n12442) );
  INV_X1 U15726 ( .A(n12443), .ZN(n12445) );
  INV_X1 U15727 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12444) );
  NAND2_X1 U15728 ( .A1(n12445), .A2(n12444), .ZN(n12446) );
  NAND2_X1 U15729 ( .A1(n12790), .A2(n12446), .ZN(n15174) );
  INV_X1 U15730 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12458) );
  INV_X1 U15731 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12449) );
  INV_X1 U15732 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12448) );
  OAI22_X1 U15733 ( .A1(n11803), .A2(n12449), .B1(n11766), .B2(n12448), .ZN(
        n12454) );
  INV_X1 U15734 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12451) );
  INV_X1 U15735 ( .A(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12450) );
  OAI22_X1 U15736 ( .A1(n12452), .A2(n12451), .B1(n12495), .B2(n12450), .ZN(
        n12453) );
  AOI211_X1 U15737 ( .C1(n12487), .C2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n12454), .B(n12453), .ZN(n12457) );
  AOI22_X1 U15738 ( .A1(n12430), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12455), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12456) );
  OAI211_X1 U15739 ( .C1(n12199), .C2(n12458), .A(n12457), .B(n12456), .ZN(
        n12466) );
  AOI22_X1 U15740 ( .A1(n12460), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U15741 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11761), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12463) );
  AOI22_X1 U15742 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12462) );
  AOI22_X1 U15743 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12461) );
  NAND4_X1 U15744 ( .A1(n12464), .A2(n12463), .A3(n12462), .A4(n12461), .ZN(
        n12465) );
  NOR2_X1 U15745 ( .A1(n12466), .A2(n12465), .ZN(n12475) );
  NAND2_X1 U15746 ( .A1(n12468), .A2(n12467), .ZN(n12474) );
  XNOR2_X1 U15747 ( .A(n12475), .B(n12474), .ZN(n12472) );
  AOI21_X1 U15748 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n11830), .A(
        n12273), .ZN(n12470) );
  NAND2_X1 U15749 ( .A1(n12511), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12469) );
  OAI211_X1 U15750 ( .C1(n12472), .C2(n12471), .A(n12470), .B(n12469), .ZN(
        n12473) );
  OAI21_X1 U15751 ( .B1(n15174), .B2(n12503), .A(n12473), .ZN(n14761) );
  XNOR2_X1 U15752 ( .A(n12790), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15166) );
  NOR2_X1 U15753 ( .A1(n12475), .A2(n12474), .ZN(n12502) );
  AOI22_X1 U15754 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11867), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12477) );
  OAI21_X1 U15755 ( .B1(n12479), .B2(n12478), .A(n12477), .ZN(n12480) );
  AOI21_X1 U15756 ( .B1(n11744), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n12480), .ZN(n12484) );
  AOI22_X1 U15757 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12481), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U15758 ( .A1(n11788), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12482) );
  NAND3_X1 U15759 ( .A1(n12484), .A2(n12483), .A3(n12482), .ZN(n12500) );
  AOI22_X1 U15760 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12485), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12489) );
  NAND2_X1 U15761 ( .A1(n12487), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12488) );
  OAI211_X1 U15762 ( .C1(n12491), .C2(n12490), .A(n12489), .B(n12488), .ZN(
        n12498) );
  INV_X1 U15763 ( .A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13838) );
  OAI22_X1 U15764 ( .A1(n12246), .A2(n13838), .B1(n12287), .B2(n12492), .ZN(
        n12497) );
  INV_X1 U15765 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13908) );
  OAI22_X1 U15766 ( .A1(n11760), .A2(n13908), .B1(n12495), .B2(n12494), .ZN(
        n12496) );
  OR3_X1 U15767 ( .A1(n12498), .A2(n12497), .A3(n12496), .ZN(n12499) );
  NOR2_X1 U15768 ( .A1(n12500), .A2(n12499), .ZN(n12501) );
  XNOR2_X1 U15769 ( .A(n12502), .B(n12501), .ZN(n12508) );
  INV_X1 U15770 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n15073) );
  NAND2_X1 U15771 ( .A1(n11830), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12504) );
  OAI211_X1 U15772 ( .C1(n12505), .C2(n15073), .A(n12504), .B(n12503), .ZN(
        n12506) );
  AOI21_X1 U15773 ( .B1(n12508), .B2(n12507), .A(n12506), .ZN(n12509) );
  AOI21_X1 U15774 ( .B1(n15166), .B2(n12273), .A(n12509), .ZN(n12802) );
  AOI22_X1 U15775 ( .A1(n12511), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12510), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12512) );
  INV_X1 U15776 ( .A(n12512), .ZN(n12513) );
  NAND2_X1 U15777 ( .A1(n12559), .A2(n13563), .ZN(n12515) );
  NAND2_X1 U15778 ( .A1(n13808), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12514) );
  XNOR2_X1 U15779 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12526) );
  NAND2_X1 U15780 ( .A1(n14084), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12517) );
  XNOR2_X1 U15781 ( .A(n12526), .B(n12525), .ZN(n12567) );
  INV_X1 U15782 ( .A(n12567), .ZN(n12524) );
  NAND2_X1 U15783 ( .A1(n13808), .A2(n13777), .ZN(n12516) );
  NAND2_X1 U15784 ( .A1(n12516), .A2(n13829), .ZN(n12530) );
  OAI21_X1 U15785 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14084), .A(
        n12517), .ZN(n12518) );
  INV_X1 U15786 ( .A(n12518), .ZN(n12519) );
  OAI211_X1 U15787 ( .C1(n12976), .C2(n13818), .A(n12530), .B(n12519), .ZN(
        n12521) );
  NAND2_X1 U15788 ( .A1(n12559), .A2(n12519), .ZN(n12520) );
  NAND2_X1 U15789 ( .A1(n12522), .A2(n12524), .ZN(n12523) );
  NAND2_X1 U15790 ( .A1(n12526), .A2(n12525), .ZN(n12528) );
  NAND2_X1 U15791 ( .A1(n21136), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12527) );
  NAND2_X1 U15792 ( .A1(n12528), .A2(n12527), .ZN(n12534) );
  XNOR2_X1 U15793 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12533) );
  XNOR2_X1 U15794 ( .A(n12534), .B(n12533), .ZN(n12568) );
  INV_X1 U15795 ( .A(n12568), .ZN(n12529) );
  NAND2_X1 U15796 ( .A1(n12559), .A2(n12529), .ZN(n12531) );
  OAI211_X1 U15797 ( .C1(n12529), .C2(n12542), .A(n12531), .B(n12530), .ZN(
        n12532) );
  NAND2_X1 U15798 ( .A1(n12534), .A2(n12533), .ZN(n12536) );
  NAND2_X1 U15799 ( .A1(n17091), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12535) );
  MUX2_X1 U15800 ( .A(n17089), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n12540) );
  XNOR2_X1 U15801 ( .A(n12541), .B(n12540), .ZN(n12569) );
  AND2_X1 U15802 ( .A1(n12542), .A2(n12569), .ZN(n12538) );
  INV_X1 U15803 ( .A(n12569), .ZN(n12537) );
  NOR2_X1 U15804 ( .A1(n15614), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12539) );
  NOR2_X1 U15805 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20942), .ZN(
        n12552) );
  AND2_X1 U15806 ( .A1(n12549), .A2(n12552), .ZN(n12570) );
  NAND2_X1 U15807 ( .A1(n12542), .A2(n12570), .ZN(n12547) );
  NAND2_X1 U15808 ( .A1(n12543), .A2(n12570), .ZN(n12544) );
  OAI22_X1 U15809 ( .A1(n12545), .A2(n12544), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n17214), .ZN(n12546) );
  INV_X1 U15810 ( .A(n12549), .ZN(n12551) );
  NOR2_X1 U15811 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n17214), .ZN(
        n12550) );
  INV_X1 U15812 ( .A(n12552), .ZN(n12553) );
  NOR2_X1 U15813 ( .A1(n12555), .A2(n12572), .ZN(n12556) );
  INV_X1 U15814 ( .A(n12572), .ZN(n12558) );
  NAND2_X1 U15816 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n17215) );
  NAND2_X1 U15817 ( .A1(n21470), .A2(n17215), .ZN(n12563) );
  NOR2_X1 U15818 ( .A1(n12120), .A2(n12977), .ZN(n13623) );
  NAND2_X1 U15819 ( .A1(n13623), .A2(n17109), .ZN(n17098) );
  OAI21_X1 U15820 ( .B1(n12561), .B2(n12563), .A(n17098), .ZN(n12564) );
  INV_X1 U15821 ( .A(n12564), .ZN(n12565) );
  OR4_X1 U15822 ( .A1(n12570), .A2(n12569), .A3(n12568), .A4(n12567), .ZN(
        n12571) );
  AND2_X1 U15823 ( .A1(n12572), .A2(n12571), .ZN(n12807) );
  NAND2_X1 U15824 ( .A1(n12807), .A2(n17215), .ZN(n12965) );
  OR2_X1 U15825 ( .A1(n17210), .A2(n12965), .ZN(n12573) );
  INV_X1 U15826 ( .A(n13758), .ZN(n13834) );
  AND4_X1 U15827 ( .A1(n13808), .A2(n13845), .A3(n13834), .A4(n12575), .ZN(
        n12576) );
  NAND2_X1 U15828 ( .A1(n12576), .A2(n15613), .ZN(n13742) );
  NOR2_X1 U15829 ( .A1(n13742), .A2(n15027), .ZN(n12577) );
  NOR2_X1 U15830 ( .A1(n15154), .A2(n13758), .ZN(n12579) );
  INV_X1 U15831 ( .A(n13763), .ZN(n12590) );
  NOR4_X1 U15832 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12583) );
  NOR4_X1 U15833 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12582) );
  NOR4_X1 U15834 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12581) );
  NOR4_X1 U15835 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12580) );
  AND4_X1 U15836 ( .A1(n12583), .A2(n12582), .A3(n12581), .A4(n12580), .ZN(
        n12588) );
  NOR4_X1 U15837 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12586) );
  NOR4_X1 U15838 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12585) );
  NOR4_X1 U15839 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12584) );
  INV_X1 U15840 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21224) );
  AND4_X1 U15841 ( .A1(n12586), .A2(n12585), .A3(n12584), .A4(n21224), .ZN(
        n12587) );
  NAND2_X1 U15842 ( .A1(n12588), .A2(n12587), .ZN(n12589) );
  NAND2_X1 U15843 ( .A1(n12590), .A2(n15085), .ZN(n15138) );
  INV_X1 U15844 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n17303) );
  NOR2_X1 U15845 ( .A1(n15138), .A2(n17303), .ZN(n12593) );
  NOR2_X2 U15846 ( .A1(n13763), .A2(n15085), .ZN(n15147) );
  AOI22_X1 U15847 ( .A1(n15147), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15154), .ZN(n12591) );
  NOR2_X1 U15848 ( .A1(n12593), .A2(n12592), .ZN(n12594) );
  NAND2_X1 U15849 ( .A1(n16931), .A2(n13549), .ZN(n12596) );
  INV_X1 U15850 ( .A(n19715), .ZN(n12599) );
  NAND2_X1 U15851 ( .A1(n12597), .A2(n20542), .ZN(n12598) );
  NAND2_X1 U15852 ( .A1(n13488), .A2(n16931), .ZN(n19716) );
  INV_X1 U15853 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20687) );
  NAND2_X1 U15854 ( .A1(n20686), .A2(n20687), .ZN(n12670) );
  OR3_X1 U15855 ( .A1(n20682), .A2(n12672), .A3(n12670), .ZN(n19871) );
  NAND2_X1 U15856 ( .A1(n20687), .A2(n13474), .ZN(n16958) );
  NOR2_X1 U15857 ( .A1(n12600), .A2(n19870), .ZN(n12674) );
  NAND2_X1 U15858 ( .A1(n12621), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12618) );
  NAND2_X1 U15859 ( .A1(n12614), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12630) );
  INV_X1 U15860 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12629) );
  INV_X1 U15861 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15921) );
  INV_X1 U15862 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19793) );
  NAND2_X1 U15863 ( .A1(n12647), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12649) );
  INV_X1 U15864 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16338) );
  INV_X1 U15865 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12603) );
  INV_X1 U15866 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16319) );
  NOR2_X1 U15867 ( .A1(n12607), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12606) );
  NOR2_X1 U15868 ( .A1(n12641), .A2(n12606), .ZN(n19747) );
  INV_X1 U15869 ( .A(n12607), .ZN(n12610) );
  INV_X1 U15870 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12608) );
  NAND2_X1 U15871 ( .A1(n9719), .A2(n12608), .ZN(n12609) );
  NAND2_X1 U15872 ( .A1(n12610), .A2(n12609), .ZN(n19760) );
  OAI21_X1 U15873 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12635), .A(
        n12611), .ZN(n19775) );
  INV_X1 U15874 ( .A(n19775), .ZN(n12638) );
  OR2_X1 U15875 ( .A1(n12614), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12612) );
  NAND2_X1 U15876 ( .A1(n12630), .A2(n12612), .ZN(n16442) );
  INV_X1 U15877 ( .A(n16442), .ZN(n15946) );
  AND2_X1 U15878 ( .A1(n12617), .A2(n12613), .ZN(n12615) );
  OR2_X1 U15879 ( .A1(n12615), .A2(n12614), .ZN(n19811) );
  OAI21_X1 U15880 ( .B1(n12616), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n12617), .ZN(n16466) );
  INV_X1 U15881 ( .A(n16466), .ZN(n19822) );
  AOI21_X1 U15882 ( .B1(n16493), .B2(n12618), .A(n12619), .ZN(n16489) );
  AOI21_X1 U15883 ( .B1(n12620), .B2(n19879), .A(n12621), .ZN(n19868) );
  AOI21_X1 U15884 ( .B1(n19954), .B2(n12626), .A(n12622), .ZN(n19942) );
  AOI21_X1 U15885 ( .B1(n16013), .B2(n12624), .A(n12623), .ZN(n16016) );
  INV_X1 U15886 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12625) );
  MUX2_X1 U15887 ( .A(n19963), .B(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .S(n20690), .Z(n16028) );
  INV_X1 U15888 ( .A(n15999), .ZN(n16002) );
  OAI21_X1 U15889 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12623), .A(
        n12626), .ZN(n16543) );
  NAND2_X1 U15890 ( .A1(n16002), .A2(n16543), .ZN(n15983) );
  OAI21_X1 U15891 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n12622), .A(
        n12620), .ZN(n16530) );
  OAI21_X1 U15892 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n12621), .A(
        n12618), .ZN(n19848) );
  NOR2_X1 U15893 ( .A1(n16489), .A2(n15952), .ZN(n19829) );
  NOR2_X1 U15894 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n12619), .ZN(
        n12627) );
  NOR2_X1 U15895 ( .A1(n12616), .A2(n12627), .ZN(n19830) );
  INV_X1 U15896 ( .A(n19830), .ZN(n12628) );
  NAND2_X1 U15897 ( .A1(n12630), .A2(n12629), .ZN(n12631) );
  NAND2_X1 U15898 ( .A1(n12632), .A2(n12631), .ZN(n16429) );
  NAND2_X1 U15899 ( .A1(n15930), .A2(n16429), .ZN(n15917) );
  NAND2_X1 U15900 ( .A1(n12632), .A2(n15921), .ZN(n12633) );
  NAND2_X1 U15901 ( .A1(n12636), .A2(n12633), .ZN(n16421) );
  INV_X1 U15902 ( .A(n16421), .ZN(n12634) );
  AOI21_X1 U15903 ( .B1(n12636), .B2(n19793), .A(n12635), .ZN(n19789) );
  INV_X1 U15904 ( .A(n19789), .ZN(n12637) );
  OAI21_X1 U15905 ( .B1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n12639), .A(
        n9719), .ZN(n15910) );
  INV_X1 U15906 ( .A(n19745), .ZN(n12640) );
  OAI21_X1 U15907 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12641), .A(
        n12643), .ZN(n15896) );
  NAND2_X1 U15908 ( .A1(n12602), .A2(n12643), .ZN(n12644) );
  NAND2_X1 U15909 ( .A1(n9621), .A2(n12644), .ZN(n16384) );
  NAND2_X1 U15910 ( .A1(n9621), .A2(n10400), .ZN(n12645) );
  AND2_X1 U15911 ( .A1(n12645), .A2(n12646), .ZN(n15879) );
  AND2_X1 U15912 ( .A1(n12646), .A2(n16357), .ZN(n12648) );
  OR2_X1 U15913 ( .A1(n12648), .A2(n12647), .ZN(n16356) );
  OAI21_X1 U15914 ( .B1(n12647), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n12649), .ZN(n16350) );
  NAND2_X1 U15915 ( .A1(n12649), .A2(n16338), .ZN(n12650) );
  AND2_X1 U15916 ( .A1(n12651), .A2(n12650), .ZN(n16341) );
  INV_X1 U15917 ( .A(n12651), .ZN(n12652) );
  OAI21_X1 U15918 ( .B1(n12652), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n12653), .ZN(n16331) );
  AND2_X1 U15919 ( .A1(n12653), .A2(n16319), .ZN(n12654) );
  NOR2_X1 U15920 ( .A1(n12656), .A2(n12654), .ZN(n16323) );
  NOR2_X1 U15921 ( .A1(n15802), .A2(n16323), .ZN(n15789) );
  NOR2_X1 U15922 ( .A1(n12656), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12657) );
  OR2_X1 U15923 ( .A1(n12655), .A2(n12657), .ZN(n16307) );
  AOI21_X1 U15924 ( .B1(n15789), .B2(n16307), .A(n10245), .ZN(n15783) );
  NOR2_X1 U15925 ( .A1(n12655), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12659) );
  NOR2_X1 U15926 ( .A1(n15783), .A2(n10537), .ZN(n12675) );
  XNOR2_X1 U15927 ( .A(n12658), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14421) );
  OAI21_X1 U15928 ( .B1(n12675), .B2(n10245), .A(n14421), .ZN(n12676) );
  NAND2_X1 U15929 ( .A1(n20687), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13552) );
  NAND2_X1 U15930 ( .A1(n20463), .A2(n20690), .ZN(n12660) );
  INV_X1 U15931 ( .A(n20545), .ZN(n19875) );
  NAND3_X1 U15932 ( .A1(n20463), .A2(P2_STATE2_REG_3__SCAN_IN), .A3(n12661), 
        .ZN(n17249) );
  AND3_X1 U15933 ( .A1(n20545), .A2(n16491), .A3(n17249), .ZN(n12662) );
  AND2_X2 U15934 ( .A1(n20682), .A2(n12662), .ZN(n19834) );
  INV_X1 U15935 ( .A(n20686), .ZN(n20539) );
  OAI21_X1 U15936 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n20539), .A(n12663), 
        .ZN(n12664) );
  INV_X1 U15937 ( .A(n12664), .ZN(n12665) );
  NAND2_X1 U15938 ( .A1(n19715), .A2(n12665), .ZN(n12666) );
  NAND2_X1 U15939 ( .A1(n13490), .A2(n12666), .ZN(n12667) );
  AOI22_X1 U15940 ( .A1(n19834), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_EBX_REG_31__SCAN_IN), .B2(n19864), .ZN(n12669) );
  NAND2_X1 U15941 ( .A1(n19856), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12668) );
  NAND2_X1 U15942 ( .A1(n12670), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n12671) );
  OR3_X1 U15943 ( .A1(n20682), .A2(n12672), .A3(n12671), .ZN(n19860) );
  OAI21_X1 U15944 ( .B1(n12675), .B2(n14421), .A(n19875), .ZN(n12678) );
  INV_X1 U15945 ( .A(n12676), .ZN(n12677) );
  AOI21_X1 U15946 ( .B1(n19806), .B2(n12678), .A(n12677), .ZN(n12679) );
  INV_X1 U15947 ( .A(n14701), .ZN(n12692) );
  INV_X1 U15948 ( .A(n14697), .ZN(n12684) );
  NAND2_X1 U15949 ( .A1(n12684), .A2(n19803), .ZN(n12690) );
  INV_X1 U15950 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12686) );
  AOI22_X1 U15951 ( .A1(n19834), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_EBX_REG_30__SCAN_IN), .B2(n19864), .ZN(n12685) );
  OAI21_X1 U15952 ( .B1(n19878), .B2(n12686), .A(n12685), .ZN(n12687) );
  AOI21_X1 U15953 ( .B1(n12692), .B2(n19768), .A(n12691), .ZN(n12693) );
  AND2_X1 U15954 ( .A1(n12960), .A2(n12765), .ZN(n12695) );
  INV_X1 U15955 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15565) );
  NAND2_X1 U15956 ( .A1(n12777), .A2(n15565), .ZN(n15343) );
  INV_X4 U15957 ( .A(n15286), .ZN(n15366) );
  NAND2_X1 U15958 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12697) );
  NAND2_X1 U15959 ( .A1(n15366), .A2(n12697), .ZN(n15330) );
  INV_X1 U15960 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15511) );
  NAND2_X1 U15961 ( .A1(n15366), .A2(n15511), .ZN(n12698) );
  INV_X1 U15962 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15522) );
  NAND2_X1 U15963 ( .A1(n15366), .A2(n15522), .ZN(n12699) );
  OR2_X1 U15964 ( .A1(n12777), .A2(n15522), .ZN(n12700) );
  AND2_X1 U15965 ( .A1(n15321), .A2(n12700), .ZN(n15309) );
  INV_X1 U15966 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15534) );
  XNOR2_X1 U15967 ( .A(n15366), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15298) );
  NAND2_X1 U15968 ( .A1(n15366), .A2(n15534), .ZN(n15311) );
  AND2_X1 U15969 ( .A1(n15298), .A2(n15311), .ZN(n12701) );
  NAND2_X1 U15970 ( .A1(n12702), .A2(n12701), .ZN(n15284) );
  NAND2_X1 U15971 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12703) );
  AND2_X1 U15972 ( .A1(n15353), .A2(n12703), .ZN(n12704) );
  NAND2_X1 U15973 ( .A1(n12720), .A2(n12714), .ZN(n12728) );
  NAND2_X1 U15974 ( .A1(n12728), .A2(n12727), .ZN(n12740) );
  AND2_X1 U15975 ( .A1(n12739), .A2(n12741), .ZN(n12705) );
  NAND2_X1 U15976 ( .A1(n12740), .A2(n12705), .ZN(n12748) );
  INV_X1 U15977 ( .A(n12748), .ZN(n12757) );
  AND2_X1 U15978 ( .A1(n12756), .A2(n12758), .ZN(n12706) );
  NAND2_X1 U15979 ( .A1(n12757), .A2(n12706), .ZN(n12766) );
  INV_X1 U15980 ( .A(n12766), .ZN(n12707) );
  NAND3_X1 U15981 ( .A1(n12707), .A2(n13519), .A3(n12765), .ZN(n12708) );
  NOR2_X1 U15982 ( .A1(n15383), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12709) );
  INV_X1 U15983 ( .A(n12960), .ZN(n12754) );
  INV_X1 U15984 ( .A(n12739), .ZN(n12710) );
  XNOR2_X1 U15985 ( .A(n12740), .B(n12710), .ZN(n12711) );
  NAND2_X1 U15986 ( .A1(n12711), .A2(n13519), .ZN(n12712) );
  INV_X1 U15987 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20908) );
  NAND2_X1 U15988 ( .A1(n12713), .A2(n13563), .ZN(n12718) );
  OAI21_X1 U15989 ( .B1(n12714), .B2(n12720), .A(n12728), .ZN(n12715) );
  OAI211_X1 U15990 ( .C1(n12715), .C2(n13622), .A(n10115), .B(n11695), .ZN(
        n12716) );
  INV_X1 U15991 ( .A(n12716), .ZN(n12717) );
  NAND2_X1 U15992 ( .A1(n12718), .A2(n12717), .ZN(n12725) );
  OR2_X1 U15993 ( .A1(n14013), .A2(n12754), .ZN(n12723) );
  NAND2_X1 U15994 ( .A1(n13818), .A2(n12719), .ZN(n12729) );
  OAI21_X1 U15995 ( .B1(n13622), .B2(n12720), .A(n12729), .ZN(n12721) );
  INV_X1 U15996 ( .A(n12721), .ZN(n12722) );
  NAND2_X1 U15997 ( .A1(n12723), .A2(n12722), .ZN(n13673) );
  NAND2_X1 U15998 ( .A1(n13673), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13672) );
  NAND2_X1 U15999 ( .A1(n13792), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13791) );
  INV_X1 U16000 ( .A(n13672), .ZN(n12724) );
  NAND2_X1 U16001 ( .A1(n12725), .A2(n12724), .ZN(n12726) );
  NAND2_X1 U16002 ( .A1(n13791), .A2(n12726), .ZN(n12734) );
  INV_X1 U16003 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20926) );
  XNOR2_X1 U16004 ( .A(n12734), .B(n20926), .ZN(n20875) );
  OR2_X1 U16005 ( .A1(n14006), .A2(n12754), .ZN(n12733) );
  XNOR2_X1 U16006 ( .A(n12728), .B(n12727), .ZN(n12731) );
  INV_X1 U16007 ( .A(n12729), .ZN(n12730) );
  AOI21_X1 U16008 ( .B1(n13519), .B2(n12731), .A(n12730), .ZN(n12732) );
  NAND2_X1 U16009 ( .A1(n12733), .A2(n12732), .ZN(n20874) );
  NAND2_X1 U16010 ( .A1(n20875), .A2(n20874), .ZN(n20873) );
  NAND2_X1 U16011 ( .A1(n12734), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12735) );
  NAND2_X1 U16012 ( .A1(n12736), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12737) );
  NAND2_X1 U16013 ( .A1(n12740), .A2(n12739), .ZN(n12742) );
  XNOR2_X1 U16014 ( .A(n12742), .B(n12741), .ZN(n12743) );
  NAND2_X1 U16015 ( .A1(n12743), .A2(n13519), .ZN(n12744) );
  INV_X1 U16016 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20900) );
  NAND2_X1 U16017 ( .A1(n12745), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12746) );
  XNOR2_X1 U16018 ( .A(n12748), .B(n12756), .ZN(n12749) );
  NAND2_X1 U16019 ( .A1(n12749), .A2(n13519), .ZN(n12750) );
  INV_X1 U16020 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12751) );
  XNOR2_X1 U16021 ( .A(n12752), .B(n12751), .ZN(n17179) );
  NAND2_X1 U16022 ( .A1(n12752), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12753) );
  NAND2_X1 U16023 ( .A1(n12757), .A2(n12756), .ZN(n12759) );
  XNOR2_X1 U16024 ( .A(n12759), .B(n12758), .ZN(n12760) );
  NAND2_X1 U16025 ( .A1(n12760), .A2(n13519), .ZN(n12761) );
  OR2_X1 U16026 ( .A1(n12762), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12763) );
  NAND2_X1 U16027 ( .A1(n12764), .A2(n12960), .ZN(n12769) );
  XNOR2_X1 U16028 ( .A(n12766), .B(n12765), .ZN(n12767) );
  NAND2_X1 U16029 ( .A1(n12767), .A2(n13519), .ZN(n12768) );
  NAND2_X1 U16030 ( .A1(n12769), .A2(n12768), .ZN(n12770) );
  XNOR2_X1 U16031 ( .A(n12770), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17168) );
  NAND2_X1 U16032 ( .A1(n12770), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12771) );
  OR2_X1 U16033 ( .A1(n15353), .A2(n15565), .ZN(n15344) );
  NOR2_X1 U16034 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12772) );
  OR2_X1 U16035 ( .A1(n15353), .A2(n12772), .ZN(n15340) );
  NAND2_X1 U16036 ( .A1(n15344), .A2(n15340), .ZN(n15332) );
  NOR2_X1 U16037 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12773) );
  INV_X1 U16038 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21418) );
  OAI21_X1 U16039 ( .B1(n12773), .B2(n15366), .A(n15281), .ZN(n12774) );
  NOR2_X1 U16040 ( .A1(n15332), .A2(n12774), .ZN(n12775) );
  INV_X1 U16041 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15246) );
  INV_X1 U16042 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21379) );
  INV_X1 U16043 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15253) );
  INV_X1 U16044 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15502) );
  NAND4_X1 U16045 ( .A1(n15246), .A2(n21379), .A3(n15253), .A4(n15502), .ZN(
        n12778) );
  AND2_X1 U16046 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12995) );
  AND2_X1 U16047 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13018) );
  AND3_X1 U16048 ( .A1(n12995), .A2(n13018), .A3(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12779) );
  INV_X1 U16049 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15467) );
  AND2_X1 U16050 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12999) );
  NAND2_X1 U16051 ( .A1(n12999), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15430) );
  NAND2_X1 U16052 ( .A1(n12780), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12784) );
  INV_X1 U16053 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15448) );
  INV_X1 U16054 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15452) );
  INV_X1 U16055 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15210) );
  NAND2_X1 U16056 ( .A1(n15452), .A2(n15210), .ZN(n15178) );
  INV_X1 U16057 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15421) );
  INV_X1 U16058 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15413) );
  NAND2_X1 U16059 ( .A1(n15421), .A2(n15413), .ZN(n15409) );
  NOR4_X1 U16060 ( .A1(n15366), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n15409), .ZN(n12783) );
  INV_X1 U16061 ( .A(n12784), .ZN(n12786) );
  AND2_X1 U16062 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15400) );
  NAND2_X1 U16063 ( .A1(n15400), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15391) );
  INV_X1 U16064 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13006) );
  NOR2_X1 U16065 ( .A1(n15391), .A2(n13006), .ZN(n13020) );
  NAND2_X1 U16066 ( .A1(n12120), .A2(n13818), .ZN(n12789) );
  NAND3_X1 U16067 ( .A1(n12788), .A2(n10115), .A3(n12789), .ZN(n12957) );
  INV_X1 U16068 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15168) );
  INV_X1 U16069 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12791) );
  INV_X1 U16070 ( .A(n21029), .ZN(n21141) );
  NAND2_X1 U16071 ( .A1(n21141), .A2(n12796), .ZN(n12793) );
  NAND2_X1 U16072 ( .A1(n12793), .A2(n11759), .ZN(n12794) );
  NAND2_X1 U16073 ( .A1(n11759), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17119) );
  NAND2_X1 U16074 ( .A1(n20709), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12795) );
  AND2_X1 U16075 ( .A1(n17119), .A2(n12795), .ZN(n13671) );
  INV_X1 U16076 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21276) );
  NOR2_X1 U16077 ( .A1(n20893), .A2(n21276), .ZN(n13021) );
  AOI21_X1 U16078 ( .B1(n20882), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13021), .ZN(n12797) );
  OAI21_X1 U16079 ( .B1(n12913), .B2(n20881), .A(n12797), .ZN(n12798) );
  INV_X1 U16080 ( .A(n12798), .ZN(n12799) );
  NOR2_X1 U16081 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17222), .ZN(n13516) );
  NAND2_X1 U16082 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n13516), .ZN(n17217) );
  INV_X1 U16083 ( .A(n17217), .ZN(n12800) );
  INV_X1 U16084 ( .A(n15382), .ZN(n20884) );
  NAND2_X1 U16085 ( .A1(n12955), .A2(n20884), .ZN(n12801) );
  NAND2_X1 U16086 ( .A1(n12804), .A2(n13818), .ZN(n12805) );
  INV_X1 U16087 ( .A(n12807), .ZN(n17103) );
  NAND2_X1 U16088 ( .A1(n17108), .A2(n9905), .ZN(n14752) );
  AND2_X2 U16089 ( .A1(n14754), .A2(n14752), .ZN(n14757) );
  NOR2_X1 U16090 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n17128) );
  NAND2_X1 U16091 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n17128), .ZN(n17126) );
  NAND2_X1 U16092 ( .A1(n11907), .A2(n13516), .ZN(n12808) );
  OAI211_X1 U16093 ( .C1(n17126), .C2(n11759), .A(n20893), .B(n12808), .ZN(
        n12809) );
  INV_X1 U16094 ( .A(n12809), .ZN(n12810) );
  INV_X1 U16095 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20913) );
  NAND2_X1 U16096 ( .A1(n12832), .A2(n20913), .ZN(n12812) );
  OAI211_X1 U16097 ( .C1(n13741), .C2(P1_EBX_REG_1__SCAN_IN), .A(n12812), .B(
        n12943), .ZN(n12814) );
  INV_X1 U16098 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n20782) );
  NAND2_X1 U16099 ( .A1(n12944), .A2(n20782), .ZN(n12813) );
  NAND2_X1 U16100 ( .A1(n12814), .A2(n12813), .ZN(n12817) );
  NAND2_X1 U16101 ( .A1(n12832), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12816) );
  NAND2_X1 U16102 ( .A1(n12816), .A2(n12815), .ZN(n13751) );
  XNOR2_X1 U16103 ( .A(n12817), .B(n13751), .ZN(n13748) );
  INV_X1 U16104 ( .A(n12817), .ZN(n12818) );
  NAND2_X1 U16105 ( .A1(n12818), .A2(n13751), .ZN(n12819) );
  NAND2_X1 U16106 ( .A1(n13746), .A2(n12819), .ZN(n13786) );
  NAND2_X1 U16107 ( .A1(n12832), .A2(n20926), .ZN(n12820) );
  OAI211_X1 U16108 ( .C1(n13741), .C2(P1_EBX_REG_2__SCAN_IN), .A(n12820), .B(
        n12943), .ZN(n12823) );
  INV_X1 U16109 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n12821) );
  NAND2_X1 U16110 ( .A1(n12944), .A2(n12821), .ZN(n12822) );
  MUX2_X1 U16111 ( .A(n12897), .B(n12943), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12827) );
  NAND2_X1 U16112 ( .A1(n13750), .A2(n20908), .ZN(n12826) );
  NAND2_X1 U16113 ( .A1(n12827), .A2(n12826), .ZN(n14045) );
  NAND2_X1 U16114 ( .A1(n12943), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12828) );
  NAND2_X1 U16115 ( .A1(n12828), .A2(n12832), .ZN(n12829) );
  OAI21_X1 U16116 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(n13741), .A(n12829), .ZN(
        n12831) );
  INV_X1 U16117 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n20768) );
  NAND2_X1 U16118 ( .A1(n12944), .A2(n20768), .ZN(n12830) );
  NAND2_X1 U16119 ( .A1(n12831), .A2(n12830), .ZN(n14168) );
  OR2_X1 U16120 ( .A1(n12897), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n12835) );
  NAND2_X1 U16121 ( .A1(n12943), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12833) );
  OAI211_X1 U16122 ( .C1(n13741), .C2(P1_EBX_REG_5__SCAN_IN), .A(n12833), .B(
        n12832), .ZN(n12834) );
  NAND2_X1 U16123 ( .A1(n12835), .A2(n12834), .ZN(n17204) );
  NAND2_X1 U16124 ( .A1(n12943), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12836) );
  NAND2_X1 U16125 ( .A1(n12836), .A2(n12832), .ZN(n12837) );
  OAI21_X1 U16126 ( .B1(P1_EBX_REG_6__SCAN_IN), .B2(n13741), .A(n12837), .ZN(
        n12840) );
  INV_X1 U16127 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n12838) );
  NAND2_X1 U16128 ( .A1(n12944), .A2(n12838), .ZN(n12839) );
  OR2_X1 U16129 ( .A1(n12897), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n12843) );
  NAND2_X1 U16130 ( .A1(n12943), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12841) );
  OAI211_X1 U16131 ( .C1(n13741), .C2(P1_EBX_REG_7__SCAN_IN), .A(n12841), .B(
        n12832), .ZN(n12842) );
  NAND2_X1 U16132 ( .A1(n12843), .A2(n12842), .ZN(n14260) );
  NAND2_X1 U16133 ( .A1(n12943), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12844) );
  NAND2_X1 U16134 ( .A1(n12844), .A2(n12832), .ZN(n12845) );
  OAI21_X1 U16135 ( .B1(P1_EBX_REG_8__SCAN_IN), .B2(n13741), .A(n12845), .ZN(
        n12848) );
  INV_X1 U16136 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n12846) );
  NAND2_X1 U16137 ( .A1(n12944), .A2(n12846), .ZN(n12847) );
  NAND2_X1 U16138 ( .A1(n12848), .A2(n12847), .ZN(n14266) );
  OR2_X1 U16139 ( .A1(n12897), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n12851) );
  NAND2_X1 U16140 ( .A1(n12943), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12849) );
  OAI211_X1 U16141 ( .C1(n13741), .C2(P1_EBX_REG_9__SCAN_IN), .A(n12849), .B(
        n12832), .ZN(n12850) );
  NAND2_X1 U16142 ( .A1(n12851), .A2(n12850), .ZN(n14273) );
  INV_X1 U16143 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15364) );
  NAND2_X1 U16144 ( .A1(n12832), .A2(n15364), .ZN(n12852) );
  OAI211_X1 U16145 ( .C1(n13741), .C2(P1_EBX_REG_10__SCAN_IN), .A(n12852), .B(
        n12943), .ZN(n12855) );
  INV_X1 U16146 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n12853) );
  NAND2_X1 U16147 ( .A1(n12944), .A2(n12853), .ZN(n12854) );
  MUX2_X1 U16148 ( .A(n12897), .B(n12943), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12857) );
  INV_X1 U16149 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15576) );
  NAND2_X1 U16150 ( .A1(n13750), .A2(n15576), .ZN(n12856) );
  NAND2_X1 U16151 ( .A1(n12832), .A2(n15565), .ZN(n12858) );
  OAI211_X1 U16152 ( .C1(P1_EBX_REG_12__SCAN_IN), .C2(n13741), .A(n12858), .B(
        n12943), .ZN(n12861) );
  INV_X1 U16153 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n12859) );
  NAND2_X1 U16154 ( .A1(n12944), .A2(n12859), .ZN(n12860) );
  NAND2_X1 U16155 ( .A1(n12861), .A2(n12860), .ZN(n14977) );
  MUX2_X1 U16156 ( .A(n12897), .B(n12943), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12863) );
  NAND2_X1 U16157 ( .A1(n13750), .A2(n15511), .ZN(n12862) );
  NAND2_X1 U16158 ( .A1(n12863), .A2(n12862), .ZN(n14962) );
  NAND2_X1 U16159 ( .A1(n12832), .A2(n15522), .ZN(n12864) );
  OAI211_X1 U16160 ( .C1(P1_EBX_REG_14__SCAN_IN), .C2(n13741), .A(n12864), .B(
        n12943), .ZN(n12866) );
  INV_X1 U16161 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n21352) );
  NAND2_X1 U16162 ( .A1(n12944), .A2(n21352), .ZN(n12865) );
  MUX2_X1 U16163 ( .A(n12897), .B(n12943), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12868) );
  NAND2_X1 U16164 ( .A1(n13750), .A2(n15534), .ZN(n12867) );
  AND2_X2 U16165 ( .A1(n14946), .A2(n14932), .ZN(n14919) );
  INV_X1 U16166 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15523) );
  NAND2_X1 U16167 ( .A1(n12832), .A2(n15523), .ZN(n12869) );
  OAI211_X1 U16168 ( .C1(P1_EBX_REG_16__SCAN_IN), .C2(n13741), .A(n12869), .B(
        n12943), .ZN(n12871) );
  INV_X1 U16169 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15061) );
  NAND2_X1 U16170 ( .A1(n12944), .A2(n15061), .ZN(n12870) );
  NAND2_X1 U16171 ( .A1(n12871), .A2(n12870), .ZN(n14920) );
  MUX2_X1 U16172 ( .A(n12897), .B(n12943), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12873) );
  INV_X1 U16173 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15514) );
  NAND2_X1 U16174 ( .A1(n13750), .A2(n15514), .ZN(n12872) );
  NAND2_X1 U16175 ( .A1(n12873), .A2(n12872), .ZN(n14904) );
  NAND2_X1 U16176 ( .A1(n12832), .A2(n15502), .ZN(n12874) );
  OAI211_X1 U16177 ( .C1(P1_EBX_REG_18__SCAN_IN), .C2(n13741), .A(n12874), .B(
        n12943), .ZN(n12876) );
  INV_X1 U16178 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15059) );
  NAND2_X1 U16179 ( .A1(n12944), .A2(n15059), .ZN(n12875) );
  MUX2_X1 U16180 ( .A(n12897), .B(n12943), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12878) );
  NAND2_X1 U16181 ( .A1(n13750), .A2(n15253), .ZN(n12877) );
  NAND2_X1 U16182 ( .A1(n12878), .A2(n12877), .ZN(n14878) );
  NAND2_X1 U16183 ( .A1(n12943), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12879) );
  NAND2_X1 U16184 ( .A1(n12879), .A2(n12832), .ZN(n12880) );
  OAI21_X1 U16185 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(n13741), .A(n12880), .ZN(
        n12882) );
  INV_X1 U16186 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15057) );
  NAND2_X1 U16187 ( .A1(n12944), .A2(n15057), .ZN(n12881) );
  NAND2_X1 U16188 ( .A1(n12882), .A2(n12881), .ZN(n14866) );
  MUX2_X1 U16189 ( .A(n12897), .B(n12943), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12884) );
  NAND2_X1 U16190 ( .A1(n13750), .A2(n21379), .ZN(n12883) );
  AND2_X1 U16191 ( .A1(n12884), .A2(n12883), .ZN(n14855) );
  NAND2_X1 U16192 ( .A1(n12832), .A2(n15467), .ZN(n12885) );
  OAI211_X1 U16193 ( .C1(P1_EBX_REG_22__SCAN_IN), .C2(n13741), .A(n12885), .B(
        n12943), .ZN(n12887) );
  INV_X1 U16194 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15055) );
  NAND2_X1 U16195 ( .A1(n12944), .A2(n15055), .ZN(n12886) );
  NAND2_X1 U16196 ( .A1(n12887), .A2(n12886), .ZN(n14843) );
  OR2_X1 U16197 ( .A1(n12897), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n12890) );
  NAND2_X1 U16198 ( .A1(n12943), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12888) );
  OAI211_X1 U16199 ( .C1(n13741), .C2(P1_EBX_REG_23__SCAN_IN), .A(n12888), .B(
        n12832), .ZN(n12889) );
  NAND2_X1 U16200 ( .A1(n12890), .A2(n12889), .ZN(n14829) );
  NAND2_X1 U16201 ( .A1(n12832), .A2(n15452), .ZN(n12891) );
  OAI211_X1 U16202 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n13741), .A(n12891), .B(
        n12943), .ZN(n12894) );
  INV_X1 U16203 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n12892) );
  NAND2_X1 U16204 ( .A1(n12944), .A2(n12892), .ZN(n12893) );
  MUX2_X1 U16205 ( .A(n12897), .B(n12943), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12896) );
  NAND2_X1 U16206 ( .A1(n13750), .A2(n15210), .ZN(n12895) );
  AND2_X1 U16207 ( .A1(n12896), .A2(n12895), .ZN(n14807) );
  MUX2_X1 U16208 ( .A(n12897), .B(n12943), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12899) );
  NAND2_X1 U16209 ( .A1(n13750), .A2(n15421), .ZN(n12898) );
  NAND2_X1 U16210 ( .A1(n12899), .A2(n12898), .ZN(n14790) );
  INV_X1 U16211 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15431) );
  NAND2_X1 U16212 ( .A1(n12832), .A2(n15431), .ZN(n12900) );
  OAI211_X1 U16213 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n13741), .A(n12900), .B(
        n12943), .ZN(n12902) );
  INV_X1 U16214 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15050) );
  NAND2_X1 U16215 ( .A1(n12944), .A2(n15050), .ZN(n12901) );
  AND2_X1 U16216 ( .A1(n12902), .A2(n12901), .ZN(n14787) );
  NOR2_X1 U16217 ( .A1(n14790), .A2(n14787), .ZN(n12903) );
  NAND2_X1 U16218 ( .A1(n14786), .A2(n12903), .ZN(n14773) );
  NAND2_X1 U16219 ( .A1(n12832), .A2(n15413), .ZN(n12904) );
  OAI211_X1 U16220 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n13741), .A(n12904), .B(
        n12943), .ZN(n12907) );
  INV_X1 U16221 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n12905) );
  NAND2_X1 U16222 ( .A1(n12944), .A2(n12905), .ZN(n12906) );
  AND2_X1 U16223 ( .A1(n12907), .A2(n12906), .ZN(n14776) );
  INV_X1 U16224 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n12908) );
  NAND2_X1 U16225 ( .A1(n21470), .A2(n12908), .ZN(n12909) );
  INV_X1 U16226 ( .A(n13750), .ZN(n12978) );
  OAI21_X1 U16227 ( .B1(n12978), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12909), .ZN(n12910) );
  MUX2_X1 U16228 ( .A(n12909), .B(n12910), .S(n12943), .Z(n14763) );
  AOI22_X1 U16229 ( .A1(n12978), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n13741), .ZN(n12945) );
  NAND2_X1 U16230 ( .A1(n17215), .A2(n20709), .ZN(n17120) );
  NAND3_X1 U16231 ( .A1(n21470), .A2(P1_EBX_REG_31__SCAN_IN), .A3(n17120), 
        .ZN(n12911) );
  INV_X2 U16232 ( .A(n12914), .ZN(n17157) );
  INV_X1 U16233 ( .A(n15166), .ZN(n12920) );
  INV_X1 U16234 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15044) );
  OR2_X1 U16235 ( .A1(n12915), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n17142) );
  INV_X1 U16236 ( .A(n17142), .ZN(n17105) );
  OR2_X1 U16237 ( .A1(n13563), .A2(n17105), .ZN(n12970) );
  INV_X1 U16238 ( .A(n17120), .ZN(n12916) );
  AND2_X1 U16239 ( .A1(n12970), .A2(n12916), .ZN(n12922) );
  INV_X1 U16240 ( .A(n12922), .ZN(n12917) );
  OAI211_X1 U16241 ( .C1(n13829), .C2(n15044), .A(n12917), .B(n13777), .ZN(
        n12918) );
  AOI22_X1 U16242 ( .A1(n20757), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20785), .ZN(n12919) );
  OAI21_X1 U16243 ( .B1(n15023), .B2(n12920), .A(n12919), .ZN(n12921) );
  AOI21_X1 U16244 ( .B1(n15397), .B2(n9580), .A(n12921), .ZN(n12941) );
  INV_X1 U16245 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21226) );
  NAND2_X1 U16246 ( .A1(n12922), .A2(n13777), .ZN(n12923) );
  NAND2_X1 U16247 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .ZN(n12927) );
  AND2_X1 U16248 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n12928) );
  INV_X1 U16249 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21247) );
  NAND3_X1 U16250 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(P1_REIP_REG_11__SCAN_IN), .ZN(n14943) );
  INV_X1 U16251 ( .A(n14943), .ZN(n12924) );
  NAND2_X1 U16252 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n12924), .ZN(n14917) );
  NOR2_X1 U16253 ( .A1(n21247), .A2(n14917), .ZN(n12925) );
  AND2_X1 U16254 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n12930) );
  NAND3_X1 U16255 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(P1_REIP_REG_18__SCAN_IN), .ZN(n12931) );
  NAND3_X1 U16256 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(P1_REIP_REG_21__SCAN_IN), .ZN(n12933) );
  NAND4_X1 U16257 ( .A1(n14824), .A2(P1_REIP_REG_25__SCAN_IN), .A3(
        P1_REIP_REG_24__SCAN_IN), .A4(P1_REIP_REG_26__SCAN_IN), .ZN(n14793) );
  NAND2_X1 U16258 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n14765) );
  INV_X1 U16259 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21272) );
  NAND2_X1 U16260 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n12938) );
  INV_X1 U16261 ( .A(n14765), .ZN(n12937) );
  NAND3_X1 U16262 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n12926) );
  NOR3_X1 U16263 ( .A1(n20784), .A2(n21226), .A3(n12926), .ZN(n20756) );
  NAND3_X1 U16264 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n20756), .ZN(n20728) );
  NOR2_X1 U16265 ( .A1(n12927), .A2(n20728), .ZN(n15009) );
  INV_X1 U16266 ( .A(n14917), .ZN(n12929) );
  NAND2_X1 U16267 ( .A1(n14991), .A2(n12929), .ZN(n14918) );
  NOR2_X1 U16268 ( .A1(n14918), .A2(n21247), .ZN(n14881) );
  INV_X1 U16269 ( .A(n12930), .ZN(n14882) );
  NOR2_X1 U16270 ( .A1(n14882), .A2(n12931), .ZN(n12932) );
  NAND2_X1 U16271 ( .A1(n14881), .A2(n12932), .ZN(n14842) );
  OR2_X1 U16272 ( .A1(n14842), .A2(n12933), .ZN(n12934) );
  NAND2_X1 U16273 ( .A1(n12934), .A2(n20729), .ZN(n14835) );
  NAND3_X1 U16274 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .A3(P1_REIP_REG_24__SCAN_IN), .ZN(n12935) );
  NAND2_X1 U16275 ( .A1(n20729), .A2(n12935), .ZN(n12936) );
  OAI21_X1 U16276 ( .B1(n20755), .B2(n12937), .A(n14800), .ZN(n14779) );
  AOI21_X1 U16277 ( .B1(n20729), .B2(n12938), .A(n14779), .ZN(n12953) );
  INV_X1 U16278 ( .A(n12953), .ZN(n12939) );
  OAI21_X1 U16279 ( .B1(n12951), .B2(P1_REIP_REG_30__SCAN_IN), .A(n12939), 
        .ZN(n12940) );
  NAND3_X1 U16280 ( .A1(n12942), .A2(n12941), .A3(n12940), .ZN(P1_U2810) );
  AOI22_X1 U16281 ( .A1(n12978), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13741), .ZN(n12948) );
  INV_X1 U16282 ( .A(n12948), .ZN(n12949) );
  AOI22_X1 U16283 ( .A1(n20757), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20785), .ZN(n12952) );
  NAND2_X1 U16284 ( .A1(n12955), .A2(n12954), .ZN(n12956) );
  INV_X1 U16285 ( .A(n12120), .ZN(n13663) );
  NAND3_X1 U16286 ( .A1(n17107), .A2(n13663), .A3(n13563), .ZN(n12968) );
  INV_X1 U16287 ( .A(n12957), .ZN(n12963) );
  NAND2_X1 U16288 ( .A1(n12959), .A2(n12958), .ZN(n12962) );
  AOI21_X1 U16289 ( .B1(n12960), .B2(n13813), .A(n13818), .ZN(n12961) );
  NAND2_X1 U16290 ( .A1(n12962), .A2(n12961), .ZN(n12982) );
  NAND2_X1 U16291 ( .A1(n12963), .A2(n12982), .ZN(n12964) );
  NAND2_X1 U16292 ( .A1(n12964), .A2(n17097), .ZN(n13635) );
  NAND2_X1 U16293 ( .A1(n13563), .A2(n17142), .ZN(n13518) );
  INV_X1 U16294 ( .A(n12965), .ZN(n12966) );
  NAND3_X1 U16295 ( .A1(n13636), .A2(n13518), .A3(n12966), .ZN(n12967) );
  NAND3_X1 U16296 ( .A1(n12968), .A2(n13635), .A3(n12967), .ZN(n12969) );
  NAND2_X1 U16297 ( .A1(n12969), .A2(n9905), .ZN(n12973) );
  NAND2_X1 U16298 ( .A1(n12970), .A2(n17215), .ZN(n12971) );
  OAI211_X1 U16299 ( .C1(n12561), .C2(n12971), .A(n13777), .B(n13760), .ZN(
        n12972) );
  NAND2_X1 U16300 ( .A1(n10051), .A2(n13829), .ZN(n17121) );
  OAI21_X1 U16301 ( .B1(n13025), .B2(n11752), .A(n17121), .ZN(n12974) );
  AND2_X2 U16302 ( .A1(n13030), .A2(n12974), .ZN(n17191) );
  INV_X1 U16303 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21452) );
  NAND2_X1 U16304 ( .A1(n15020), .A2(n13839), .ZN(n12975) );
  AOI22_X1 U16305 ( .A1(n12978), .A2(n12977), .B1(n12976), .B2(n12975), .ZN(
        n12981) );
  NAND2_X1 U16306 ( .A1(n10114), .A2(n12944), .ZN(n12979) );
  NAND4_X1 U16307 ( .A1(n12982), .A2(n12981), .A3(n12980), .A4(n12979), .ZN(
        n13620) );
  NAND2_X1 U16308 ( .A1(n12984), .A2(n12983), .ZN(n12985) );
  AND2_X1 U16309 ( .A1(n13623), .A2(n21470), .ZN(n17101) );
  NOR2_X1 U16310 ( .A1(n20912), .A2(n20891), .ZN(n15602) );
  INV_X1 U16311 ( .A(n15602), .ZN(n15521) );
  NAND2_X1 U16312 ( .A1(n13008), .A2(n13790), .ZN(n20931) );
  NOR2_X1 U16313 ( .A1(n20916), .A2(n13030), .ZN(n20935) );
  INV_X1 U16314 ( .A(n20935), .ZN(n12986) );
  NOR2_X1 U16315 ( .A1(n20900), .A2(n20908), .ZN(n20892) );
  NAND2_X1 U16316 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20892), .ZN(
        n15541) );
  AOI21_X1 U16317 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20914) );
  NOR2_X1 U16318 ( .A1(n15541), .A2(n20914), .ZN(n15587) );
  NAND3_X1 U16319 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15584) );
  INV_X1 U16320 ( .A(n15584), .ZN(n12987) );
  AND3_X1 U16321 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n12987), .ZN(n15577) );
  AND2_X1 U16322 ( .A1(n15577), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15563) );
  AND2_X1 U16323 ( .A1(n15563), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13011) );
  NAND2_X1 U16324 ( .A1(n15587), .A2(n13011), .ZN(n13013) );
  OR2_X1 U16325 ( .A1(n15511), .A2(n13013), .ZN(n12988) );
  NAND2_X1 U16326 ( .A1(n20891), .A2(n12988), .ZN(n12989) );
  AND2_X1 U16327 ( .A1(n15583), .A2(n12989), .ZN(n15499) );
  AND2_X1 U16328 ( .A1(n13011), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15542) );
  NOR2_X1 U16329 ( .A1(n20926), .A2(n20913), .ZN(n20915) );
  INV_X1 U16330 ( .A(n20915), .ZN(n12990) );
  NOR2_X1 U16331 ( .A1(n15541), .A2(n12990), .ZN(n15559) );
  NAND4_X1 U16332 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15501) );
  NOR2_X1 U16333 ( .A1(n15501), .A2(n15502), .ZN(n12991) );
  NAND3_X1 U16334 ( .A1(n15542), .A2(n15559), .A3(n12991), .ZN(n12993) );
  INV_X1 U16335 ( .A(n12991), .ZN(n12992) );
  AOI22_X1 U16336 ( .A1(n20912), .A2(n12993), .B1(n20891), .B2(n12992), .ZN(
        n12994) );
  NAND2_X1 U16337 ( .A1(n15499), .A2(n12994), .ZN(n15491) );
  INV_X1 U16338 ( .A(n12995), .ZN(n15244) );
  OR2_X1 U16339 ( .A1(n15491), .A2(n15244), .ZN(n12996) );
  NAND2_X1 U16340 ( .A1(n15602), .A2(n15583), .ZN(n15585) );
  INV_X1 U16341 ( .A(n13018), .ZN(n12997) );
  NAND2_X1 U16342 ( .A1(n15521), .A2(n12997), .ZN(n12998) );
  NAND2_X1 U16343 ( .A1(n20891), .A2(n15452), .ZN(n13002) );
  NAND2_X1 U16344 ( .A1(n20936), .A2(n15430), .ZN(n13001) );
  INV_X1 U16345 ( .A(n12999), .ZN(n15429) );
  NAND2_X1 U16346 ( .A1(n13008), .A2(n15429), .ZN(n13000) );
  NAND3_X1 U16347 ( .A1(n13002), .A2(n13001), .A3(n13000), .ZN(n13003) );
  NAND2_X1 U16348 ( .A1(n15428), .A2(n15602), .ZN(n13007) );
  INV_X1 U16349 ( .A(n13007), .ZN(n13005) );
  NAND3_X1 U16350 ( .A1(n15428), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13004) );
  INV_X1 U16351 ( .A(n20936), .ZN(n13010) );
  NAND2_X1 U16352 ( .A1(n13008), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13009) );
  NAND2_X1 U16353 ( .A1(n13010), .A2(n13009), .ZN(n20910) );
  AND2_X1 U16354 ( .A1(n13011), .A2(n15559), .ZN(n13012) );
  NAND2_X1 U16355 ( .A1(n20910), .A2(n13012), .ZN(n13016) );
  INV_X1 U16356 ( .A(n13013), .ZN(n13014) );
  NAND2_X1 U16357 ( .A1(n20891), .A2(n13014), .ZN(n13015) );
  NAND2_X1 U16358 ( .A1(n13016), .A2(n13015), .ZN(n15510) );
  NOR2_X1 U16359 ( .A1(n15501), .A2(n15511), .ZN(n13017) );
  NAND2_X1 U16360 ( .A1(n15510), .A2(n13017), .ZN(n15504) );
  NOR2_X1 U16361 ( .A1(n15493), .A2(n15244), .ZN(n15477) );
  NAND2_X1 U16362 ( .A1(n15477), .A2(n13018), .ZN(n15461) );
  NOR3_X1 U16363 ( .A1(n15461), .A2(n15430), .A3(n15431), .ZN(n15419) );
  INV_X1 U16364 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13019) );
  NAND3_X1 U16365 ( .A1(n15419), .A2(n13020), .A3(n13019), .ZN(n13023) );
  INV_X1 U16366 ( .A(n13021), .ZN(n13022) );
  AOI21_X1 U16367 ( .B1(n15043), .B2(n17191), .A(n13024), .ZN(n13032) );
  OAI21_X1 U16368 ( .B1(n13845), .B2(n13025), .A(n17098), .ZN(n13026) );
  INV_X1 U16369 ( .A(n13026), .ZN(n13027) );
  NAND3_X1 U16370 ( .A1(n13028), .A2(n13027), .A3(n17112), .ZN(n13029) );
  NAND2_X1 U16371 ( .A1(n13032), .A2(n13031), .ZN(P1_U3000) );
  INV_X1 U16372 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21367) );
  NOR2_X4 U16373 ( .A1(n17789), .A2(n13042), .ZN(n18026) );
  AOI22_X1 U16374 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13037) );
  AOI22_X1 U16375 ( .A1(n18063), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18059), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13036) );
  NOR2_X2 U16376 ( .A1(n13043), .A2(n19508), .ZN(n13081) );
  AOI22_X1 U16377 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18038), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13035) );
  AOI22_X1 U16378 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13253), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13034) );
  AOI22_X1 U16379 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18001), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13038) );
  OAI21_X1 U16380 ( .B1(n13223), .B2(n18100), .A(n13038), .ZN(n13039) );
  INV_X1 U16381 ( .A(n13039), .ZN(n13048) );
  NOR2_X2 U16382 ( .A1(n13041), .A2(n19508), .ZN(n13202) );
  AOI22_X1 U16383 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13047) );
  AOI22_X1 U16384 ( .A1(n13232), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13046) );
  INV_X2 U16385 ( .A(n13054), .ZN(n13197) );
  AOI22_X1 U16386 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n9594), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13053) );
  AOI22_X1 U16387 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18066), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n9588), .ZN(n13052) );
  AOI22_X1 U16388 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n17945), .ZN(n13051) );
  AOI22_X1 U16389 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9590), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n13253), .ZN(n13050) );
  NAND4_X1 U16390 ( .A1(n13053), .A2(n13052), .A3(n13051), .A4(n13050), .ZN(
        n13060) );
  AOI22_X1 U16391 ( .A1(n18063), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17830), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13058) );
  AOI22_X1 U16392 ( .A1(n13054), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18062), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13057) );
  AOI22_X1 U16393 ( .A1(n17960), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n18026), .ZN(n13056) );
  AOI22_X1 U16394 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18001), .B1(
        n18059), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13055) );
  NAND4_X1 U16395 ( .A1(n13058), .A2(n13057), .A3(n13056), .A4(n13055), .ZN(
        n13059) );
  AOI22_X1 U16396 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13065) );
  AOI22_X1 U16397 ( .A1(n17960), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18044), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13064) );
  AOI22_X1 U16398 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13063) );
  AOI22_X1 U16399 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13253), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13062) );
  NAND4_X1 U16400 ( .A1(n13065), .A2(n13064), .A3(n13063), .A4(n13062), .ZN(
        n13071) );
  AOI22_X1 U16401 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13069) );
  AOI22_X1 U16402 ( .A1(n18063), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17961), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13068) );
  AOI22_X1 U16403 ( .A1(n18059), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17830), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13067) );
  AOI22_X1 U16404 ( .A1(n18001), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13066) );
  NAND4_X1 U16405 ( .A1(n13069), .A2(n13068), .A3(n13067), .A4(n13066), .ZN(
        n13070) );
  INV_X1 U16406 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19674) );
  NOR2_X2 U16407 ( .A1(n13297), .A2(n19674), .ZN(n18719) );
  INV_X1 U16408 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21354) );
  NAND2_X1 U16409 ( .A1(n18701), .A2(n13075), .ZN(n18688) );
  INV_X1 U16410 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n19011) );
  AOI22_X1 U16411 ( .A1(n18063), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17945), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13080) );
  AOI22_X1 U16412 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18062), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13079) );
  CLKBUF_X3 U16413 ( .A(n13076), .Z(n18043) );
  AOI22_X1 U16414 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17830), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13078) );
  AOI22_X1 U16415 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13077) );
  NAND4_X1 U16416 ( .A1(n13080), .A2(n13079), .A3(n13078), .A4(n13077), .ZN(
        n13088) );
  BUF_X4 U16417 ( .A(n13081), .Z(n18038) );
  AOI22_X1 U16418 ( .A1(n18038), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13086) );
  INV_X2 U16419 ( .A(n13183), .ZN(n18064) );
  AOI22_X1 U16420 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18064), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13085) );
  AOI22_X1 U16421 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13084) );
  AOI22_X1 U16422 ( .A1(n18044), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13083) );
  NAND4_X1 U16423 ( .A1(n13086), .A2(n13085), .A3(n13084), .A4(n13083), .ZN(
        n13087) );
  XNOR2_X1 U16424 ( .A(n19011), .B(n13089), .ZN(n18689) );
  NAND2_X1 U16425 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13089), .ZN(
        n13090) );
  AOI22_X1 U16426 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18064), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13100) );
  AOI22_X1 U16427 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13099) );
  AOI22_X1 U16428 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n9587), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13091) );
  OAI21_X1 U16429 ( .B1(n13223), .B2(n18092), .A(n13091), .ZN(n13097) );
  AOI22_X1 U16430 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13095) );
  AOI22_X1 U16431 ( .A1(n18063), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18001), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13094) );
  AOI22_X1 U16432 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18044), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13093) );
  AOI22_X1 U16433 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17945), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13092) );
  NAND4_X1 U16434 ( .A1(n13095), .A2(n13094), .A3(n13093), .A4(n13092), .ZN(
        n13096) );
  AOI211_X1 U16435 ( .C1(n17960), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n13097), .B(n13096), .ZN(n13098) );
  NAND3_X1 U16436 ( .A1(n13100), .A2(n13099), .A3(n13098), .ZN(n13299) );
  INV_X1 U16437 ( .A(n13299), .ZN(n18233) );
  XNOR2_X1 U16438 ( .A(n18233), .B(n13114), .ZN(n18681) );
  AOI22_X1 U16439 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17830), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13107) );
  AOI22_X1 U16440 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13106) );
  AOI22_X1 U16441 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13105) );
  AOI22_X1 U16442 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13104) );
  NAND4_X1 U16443 ( .A1(n13107), .A2(n13106), .A3(n13105), .A4(n13104), .ZN(
        n13113) );
  AOI22_X1 U16444 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13111) );
  AOI22_X1 U16445 ( .A1(n18063), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18044), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13110) );
  AOI22_X1 U16446 ( .A1(n17960), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13109) );
  AOI22_X1 U16447 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18064), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13108) );
  NAND4_X1 U16448 ( .A1(n13111), .A2(n13110), .A3(n13109), .A4(n13108), .ZN(
        n13112) );
  XOR2_X1 U16449 ( .A(n18229), .B(n13125), .Z(n18663) );
  INV_X1 U16450 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18985) );
  AOI22_X1 U16451 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13124) );
  AOI22_X1 U16452 ( .A1(n18063), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17961), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13123) );
  AOI22_X1 U16453 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13115) );
  OAI21_X1 U16454 ( .B1(n13223), .B2(n17829), .A(n13115), .ZN(n13121) );
  AOI22_X1 U16455 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13119) );
  AOI22_X1 U16456 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18038), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13118) );
  AOI22_X1 U16457 ( .A1(n18064), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18001), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13117) );
  AOI22_X1 U16458 ( .A1(n9587), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13116) );
  NAND4_X1 U16459 ( .A1(n13119), .A2(n13118), .A3(n13117), .A4(n13116), .ZN(
        n13120) );
  AOI211_X1 U16460 ( .C1(n17041), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n13121), .B(n13120), .ZN(n13122) );
  NAND3_X1 U16461 ( .A1(n13124), .A2(n13123), .A3(n13122), .ZN(n13300) );
  INV_X1 U16462 ( .A(n13300), .ZN(n18226) );
  XNOR2_X1 U16463 ( .A(n18226), .B(n13138), .ZN(n13126) );
  XOR2_X1 U16464 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n13126), .Z(
        n18651) );
  NAND2_X1 U16465 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13126), .ZN(
        n13127) );
  AOI22_X1 U16466 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13131) );
  AOI22_X1 U16467 ( .A1(n18038), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18044), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13130) );
  AOI22_X1 U16468 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13129) );
  AOI22_X1 U16469 ( .A1(n18063), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13128) );
  NAND4_X1 U16470 ( .A1(n13131), .A2(n13130), .A3(n13129), .A4(n13128), .ZN(
        n13137) );
  AOI22_X1 U16471 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18064), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13135) );
  AOI22_X1 U16472 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13134) );
  AOI22_X1 U16473 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17830), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13133) );
  AOI22_X1 U16474 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13132) );
  NAND4_X1 U16475 ( .A1(n13135), .A2(n13134), .A3(n13133), .A4(n13132), .ZN(
        n13136) );
  NAND2_X1 U16476 ( .A1(n13141), .A2(n13140), .ZN(n13142) );
  INV_X1 U16477 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18940) );
  INV_X1 U16478 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18917) );
  NOR2_X1 U16479 ( .A1(n18940), .A2(n18917), .ZN(n18916) );
  NAND2_X1 U16480 ( .A1(n18916), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18903) );
  NOR2_X1 U16481 ( .A1(n21454), .A2(n18903), .ZN(n18873) );
  NAND2_X1 U16482 ( .A1(n18873), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18862) );
  INV_X1 U16483 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18876) );
  NOR2_X1 U16484 ( .A1(n18862), .A2(n18876), .ZN(n13336) );
  NAND2_X1 U16485 ( .A1(n13336), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18780) );
  NAND2_X1 U16486 ( .A1(n18940), .A2(n18917), .ZN(n18605) );
  NOR4_X1 U16487 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A4(n18605), .ZN(n13144) );
  INV_X1 U16488 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18856) );
  INV_X1 U16489 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18839) );
  NOR2_X1 U16490 ( .A1(n18856), .A2(n18839), .ZN(n18830) );
  NAND2_X1 U16491 ( .A1(n18830), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18782) );
  INV_X1 U16492 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18480) );
  INV_X1 U16493 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18471) );
  NOR2_X1 U16494 ( .A1(n18480), .A2(n18471), .ZN(n18803) );
  NAND2_X1 U16495 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18803), .ZN(
        n13149) );
  NOR2_X1 U16496 ( .A1(n18782), .A2(n13149), .ZN(n18792) );
  NAND2_X1 U16497 ( .A1(n18792), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18726) );
  INV_X1 U16498 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18767) );
  NOR2_X1 U16499 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18634), .ZN(
        n18503) );
  NAND2_X1 U16500 ( .A1(n18503), .A2(n18480), .ZN(n13147) );
  NOR2_X1 U16501 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n13147), .ZN(
        n18466) );
  INV_X1 U16502 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18800) );
  NAND2_X1 U16503 ( .A1(n18466), .A2(n18800), .ZN(n18452) );
  NAND2_X1 U16504 ( .A1(n18830), .A2(n18453), .ZN(n18465) );
  INV_X1 U16505 ( .A(n13149), .ZN(n18789) );
  AND2_X1 U16506 ( .A1(n18789), .A2(n10550), .ZN(n13150) );
  INV_X1 U16507 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18409) );
  NAND2_X1 U16508 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18730) );
  INV_X1 U16509 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n18367) );
  NAND2_X1 U16510 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18634), .ZN(
        n17286) );
  NAND2_X1 U16511 ( .A1(n13153), .A2(n13152), .ZN(n13154) );
  OAI21_X1 U16512 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n21367), .A(
        n13157), .ZN(n13156) );
  INV_X1 U16513 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19655) );
  AOI22_X1 U16514 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n10142), .B1(
        n18634), .B2(n19655), .ZN(n13158) );
  AOI22_X1 U16515 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n21439), .B1(
        n13165), .B2(n19654), .ZN(n13170) );
  NOR2_X1 U16516 ( .A1(n13165), .A2(n19654), .ZN(n13171) );
  NAND2_X1 U16517 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n21439), .ZN(
        n13166) );
  OAI22_X1 U16518 ( .A1(n13170), .A2(n19517), .B1(n13171), .B2(n13166), .ZN(
        n13169) );
  AOI211_X1 U16519 ( .C1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .C2(n13162), .A(
        n13291), .B(n13169), .ZN(n13289) );
  XNOR2_X1 U16520 ( .A(n13168), .B(n13167), .ZN(n13296) );
  OAI21_X1 U16521 ( .B1(n13171), .B2(n19517), .A(n13170), .ZN(n13172) );
  INV_X2 U16522 ( .A(n13223), .ZN(n18065) );
  AOI22_X1 U16523 ( .A1(n18065), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13176) );
  AOI22_X1 U16524 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13175) );
  AOI22_X1 U16525 ( .A1(n18058), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13174) );
  AOI22_X1 U16526 ( .A1(n9587), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13173) );
  NAND4_X1 U16527 ( .A1(n13176), .A2(n13175), .A3(n13174), .A4(n13173), .ZN(
        n13182) );
  AOI22_X1 U16528 ( .A1(n17961), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13180) );
  AOI22_X1 U16529 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17946), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13179) );
  AOI22_X1 U16530 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13178) );
  AOI22_X1 U16531 ( .A1(n18038), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18059), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13177) );
  NAND4_X1 U16532 ( .A1(n13180), .A2(n13179), .A3(n13178), .A4(n13177), .ZN(
        n13181) );
  AOI22_X1 U16533 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13196) );
  AOI22_X1 U16534 ( .A1(n17946), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13195) );
  INV_X1 U16535 ( .A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13192) );
  AOI22_X1 U16536 ( .A1(n18059), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13185) );
  INV_X1 U16537 ( .A(n13186), .ZN(n13191) );
  AOI22_X1 U16538 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13190) );
  AOI22_X1 U16539 ( .A1(n18065), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13252), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13189) );
  AOI22_X1 U16540 ( .A1(n17945), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18038), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13188) );
  AOI22_X1 U16541 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13253), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13187) );
  INV_X1 U16542 ( .A(n13193), .ZN(n13194) );
  NOR2_X1 U16543 ( .A1(n17146), .A2(n16967), .ZN(n19711) );
  AOI22_X1 U16544 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13201) );
  AOI22_X1 U16545 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18062), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13200) );
  AOI22_X1 U16546 ( .A1(n18044), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13253), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13199) );
  AOI22_X1 U16547 ( .A1(n18018), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13198) );
  NAND4_X1 U16548 ( .A1(n13201), .A2(n13200), .A3(n13199), .A4(n13198), .ZN(
        n13208) );
  AOI22_X1 U16549 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13206) );
  AOI22_X1 U16550 ( .A1(n18038), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13205) );
  AOI22_X1 U16551 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17830), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13204) );
  AOI22_X1 U16552 ( .A1(n18045), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13203) );
  NAND4_X1 U16553 ( .A1(n13206), .A2(n13205), .A3(n13204), .A4(n13203), .ZN(
        n13207) );
  AOI22_X1 U16554 ( .A1(n18059), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13212) );
  AOI22_X1 U16555 ( .A1(n18038), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13211) );
  AOI22_X1 U16556 ( .A1(n18065), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13210) );
  AOI22_X1 U16557 ( .A1(n9587), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18064), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13209) );
  NAND4_X1 U16558 ( .A1(n13212), .A2(n13211), .A3(n13210), .A4(n13209), .ZN(
        n13218) );
  AOI22_X1 U16559 ( .A1(n17946), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18062), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13216) );
  AOI22_X1 U16560 ( .A1(n17945), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13215) );
  AOI22_X1 U16561 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17961), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13214) );
  AOI22_X1 U16562 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13213) );
  NAND4_X1 U16563 ( .A1(n13216), .A2(n13215), .A3(n13214), .A4(n13213), .ZN(
        n13217) );
  AOI22_X1 U16564 ( .A1(n18038), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13222) );
  AOI22_X1 U16565 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13221) );
  AOI22_X1 U16566 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18062), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13220) );
  AOI22_X1 U16567 ( .A1(n13253), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13219) );
  NAND4_X1 U16568 ( .A1(n13222), .A2(n13221), .A3(n13220), .A4(n13219), .ZN(
        n13229) );
  AOI22_X1 U16569 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18065), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13227) );
  AOI22_X1 U16570 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17041), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13226) );
  AOI22_X1 U16571 ( .A1(n17946), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13225) );
  AOI22_X1 U16572 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9594), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13224) );
  NAND4_X1 U16573 ( .A1(n13227), .A2(n13226), .A3(n13225), .A4(n13224), .ZN(
        n13228) );
  AOI22_X1 U16574 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18065), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13240) );
  AOI22_X1 U16575 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13239) );
  BUF_X1 U16576 ( .A(n13230), .Z(n18018) );
  AOI22_X1 U16577 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13231) );
  OAI21_X1 U16578 ( .B1(n13183), .B2(n18100), .A(n13231), .ZN(n13238) );
  AOI22_X1 U16579 ( .A1(n17961), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13236) );
  AOI22_X1 U16580 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13235) );
  AOI22_X1 U16581 ( .A1(n17960), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18010), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13234) );
  AOI22_X1 U16582 ( .A1(n18044), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13253), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13233) );
  NAND4_X1 U16583 ( .A1(n13236), .A2(n13235), .A3(n13234), .A4(n13233), .ZN(
        n13237) );
  NOR2_X1 U16584 ( .A1(n19074), .A2(n13266), .ZN(n13269) );
  AOI22_X1 U16585 ( .A1(n18059), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18065), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13244) );
  AOI22_X1 U16586 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13243) );
  AOI22_X1 U16587 ( .A1(n17946), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13242) );
  AOI22_X1 U16588 ( .A1(n17945), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13241) );
  NAND4_X1 U16589 ( .A1(n13244), .A2(n13243), .A3(n13242), .A4(n13241), .ZN(
        n13250) );
  AOI22_X1 U16590 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13248) );
  AOI22_X1 U16591 ( .A1(n17961), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13247) );
  AOI22_X1 U16592 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13246) );
  AOI22_X1 U16593 ( .A1(n17960), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13245) );
  NAND4_X1 U16594 ( .A1(n13248), .A2(n13247), .A3(n13246), .A4(n13245), .ZN(
        n13249) );
  AOI22_X1 U16595 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13251) );
  AOI22_X1 U16596 ( .A1(n17945), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13257) );
  AOI22_X1 U16597 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18059), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13256) );
  AOI22_X1 U16598 ( .A1(n17946), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17830), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13255) );
  AOI22_X1 U16599 ( .A1(n13253), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13252), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13254) );
  AOI22_X1 U16600 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n9594), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13258) );
  INV_X1 U16601 ( .A(n13258), .ZN(n13261) );
  AOI22_X1 U16602 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18038), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13259) );
  INV_X1 U16603 ( .A(n13259), .ZN(n13260) );
  NOR2_X1 U16604 ( .A1(n19070), .A2(n13355), .ZN(n19483) );
  NAND3_X1 U16605 ( .A1(n13285), .A2(n13269), .A3(n19483), .ZN(n17060) );
  NAND2_X1 U16606 ( .A1(n19500), .A2(n13278), .ZN(n13263) );
  NAND2_X1 U16607 ( .A1(n19078), .A2(n19070), .ZN(n13281) );
  NOR2_X1 U16608 ( .A1(n13350), .A2(n10543), .ZN(n17062) );
  NAND2_X1 U16609 ( .A1(n18113), .A2(n13355), .ZN(n13280) );
  NOR2_X1 U16610 ( .A1(n19084), .A2(n13280), .ZN(n13265) );
  AND4_X2 U16611 ( .A1(n19056), .A2(n19066), .A3(n19070), .A4(n13265), .ZN(
        n19486) );
  NOR2_X1 U16612 ( .A1(n19059), .A2(n17743), .ZN(n13272) );
  INV_X1 U16613 ( .A(n13272), .ZN(n13270) );
  NAND2_X1 U16614 ( .A1(n19074), .A2(n13355), .ZN(n13267) );
  INV_X1 U16615 ( .A(n13280), .ZN(n13277) );
  INV_X1 U16616 ( .A(n13269), .ZN(n13352) );
  NOR2_X1 U16617 ( .A1(n19084), .A2(n19500), .ZN(n17148) );
  NOR3_X1 U16618 ( .A1(n19056), .A2(n17148), .A3(n19691), .ZN(n13348) );
  AOI21_X1 U16619 ( .B1(n13352), .B2(n10543), .A(n13348), .ZN(n13276) );
  NAND2_X1 U16620 ( .A1(n19062), .A2(n13270), .ZN(n13349) );
  NAND2_X1 U16621 ( .A1(n13280), .A2(n13349), .ZN(n13275) );
  OR2_X1 U16622 ( .A1(n13272), .A2(n13271), .ZN(n13273) );
  AOI21_X1 U16623 ( .B1(n19062), .B2(n19056), .A(n19500), .ZN(n13279) );
  INV_X1 U16624 ( .A(n13279), .ZN(n13283) );
  NAND2_X1 U16625 ( .A1(n13281), .A2(n13280), .ZN(n13282) );
  NAND2_X1 U16626 ( .A1(n13283), .A2(n13282), .ZN(n13284) );
  NAND2_X2 U16627 ( .A1(n13287), .A2(n17416), .ZN(n19032) );
  NOR2_X1 U16628 ( .A1(n19059), .A2(n13285), .ZN(n19488) );
  AOI21_X1 U16629 ( .B1(n13287), .B2(n19488), .A(n13286), .ZN(n19485) );
  NOR2_X4 U16630 ( .A1(n19691), .A2(n18851), .ZN(n18893) );
  NAND2_X1 U16631 ( .A1(n19062), .A2(n19691), .ZN(n13358) );
  INV_X1 U16632 ( .A(n13289), .ZN(n13295) );
  XOR2_X1 U16633 ( .A(n13291), .B(n13290), .Z(n13294) );
  AOI21_X1 U16634 ( .B1(n13294), .B2(n13293), .A(n13292), .ZN(n17063) );
  OAI21_X1 U16635 ( .B1(n13296), .B2(n13295), .A(n17063), .ZN(n19524) );
  NOR2_X1 U16636 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n19696), .ZN(n19552) );
  NAND2_X1 U16637 ( .A1(n13359), .A2(n18635), .ZN(n13347) );
  NOR2_X1 U16638 ( .A1(n9660), .A2(n13298), .ZN(n13306) );
  NOR2_X1 U16639 ( .A1(n13306), .A2(n18236), .ZN(n13305) );
  NAND2_X1 U16640 ( .A1(n13305), .A2(n13299), .ZN(n13303) );
  NOR2_X1 U16641 ( .A1(n18229), .A2(n13303), .ZN(n13302) );
  NAND2_X1 U16642 ( .A1(n13302), .A2(n13300), .ZN(n13301) );
  NOR2_X1 U16643 ( .A1(n18222), .A2(n13301), .ZN(n13322) );
  INV_X1 U16644 ( .A(n18222), .ZN(n17287) );
  XNOR2_X1 U16645 ( .A(n13301), .B(n17287), .ZN(n18643) );
  XNOR2_X1 U16646 ( .A(n13302), .B(n18226), .ZN(n13315) );
  XOR2_X1 U16647 ( .A(n13303), .B(n18229), .Z(n13304) );
  NAND2_X1 U16648 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13304), .ZN(
        n13314) );
  XNOR2_X1 U16649 ( .A(n18985), .B(n13304), .ZN(n18667) );
  INV_X1 U16650 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18998) );
  XNOR2_X1 U16651 ( .A(n13305), .B(n18233), .ZN(n18675) );
  NAND2_X1 U16652 ( .A1(n13307), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13312) );
  XNOR2_X1 U16653 ( .A(n18241), .B(n9660), .ZN(n13308) );
  OR2_X1 U16654 ( .A1(n21354), .A2(n13308), .ZN(n13311) );
  XNOR2_X1 U16655 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n13308), .ZN(
        n18705) );
  AOI21_X1 U16656 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18247), .A(
        n10085), .ZN(n13310) );
  NOR2_X1 U16657 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18247), .ZN(
        n13309) );
  AOI221_X1 U16658 ( .B1(n10085), .B2(n18247), .C1(n13310), .C2(n19674), .A(
        n13309), .ZN(n18704) );
  NAND2_X1 U16659 ( .A1(n18705), .A2(n18704), .ZN(n18703) );
  NAND2_X1 U16660 ( .A1(n13311), .A2(n18703), .ZN(n18691) );
  NAND2_X1 U16661 ( .A1(n18675), .A2(n18676), .ZN(n18674) );
  NOR2_X1 U16662 ( .A1(n18675), .A2(n18676), .ZN(n13313) );
  AOI21_X1 U16663 ( .B1(n18998), .B2(n18674), .A(n13313), .ZN(n18666) );
  NAND2_X1 U16664 ( .A1(n18667), .A2(n18666), .ZN(n18665) );
  NAND2_X1 U16665 ( .A1(n13315), .A2(n13316), .ZN(n13317) );
  INV_X1 U16666 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13318) );
  NAND2_X1 U16667 ( .A1(n13322), .A2(n13319), .ZN(n13323) );
  INV_X1 U16668 ( .A(n13319), .ZN(n13321) );
  NAND2_X1 U16669 ( .A1(n13322), .A2(n13321), .ZN(n13320) );
  INV_X1 U16670 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18543) );
  INV_X1 U16671 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n18734) );
  NOR2_X1 U16672 ( .A1(n18734), .A2(n18367), .ZN(n17279) );
  NAND2_X1 U16673 ( .A1(n17279), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17136) );
  NAND2_X1 U16674 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18729) );
  NOR2_X1 U16675 ( .A1(n18726), .A2(n18729), .ZN(n13339) );
  INV_X1 U16676 ( .A(n18730), .ZN(n13324) );
  NAND2_X1 U16677 ( .A1(n13339), .A2(n13324), .ZN(n17262) );
  NOR4_X1 U16678 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17136), .A3(
        n17262), .A4(n21367), .ZN(n13338) );
  INV_X1 U16679 ( .A(n13339), .ZN(n18748) );
  NAND2_X1 U16680 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17281), .ZN(
        n13325) );
  AOI22_X1 U16681 ( .A1(n18786), .A2(n13338), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13325), .ZN(n13360) );
  NAND2_X1 U16682 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18628) );
  NAND2_X1 U16683 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n19045) );
  NAND2_X1 U16684 ( .A1(n19650), .A2(n19045), .ZN(n19699) );
  NAND3_X1 U16685 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17652) );
  INV_X1 U16686 ( .A(n17652), .ZN(n13327) );
  NAND2_X1 U16687 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18486) );
  INV_X1 U16688 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18472) );
  NAND2_X1 U16689 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18447) );
  NAND2_X1 U16690 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18413) );
  NAND2_X1 U16691 ( .A1(n18394), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n18375) );
  INV_X1 U16692 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18714) );
  NAND2_X1 U16693 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18376) );
  INV_X1 U16694 ( .A(n18376), .ZN(n13329) );
  INV_X1 U16695 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n17459) );
  INV_X1 U16696 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19635) );
  NAND2_X1 U16697 ( .A1(n19656), .A2(n19650), .ZN(n19659) );
  NOR2_X1 U16698 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19659), .ZN(n19708) );
  NOR2_X1 U16699 ( .A1(n19635), .A2(n19024), .ZN(n13369) );
  INV_X1 U16700 ( .A(n18375), .ZN(n18360) );
  NAND3_X1 U16701 ( .A1(n18360), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17274) );
  NOR2_X1 U16702 ( .A1(n17459), .A2(n17274), .ZN(n13333) );
  INV_X1 U16703 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19692) );
  NOR2_X1 U16704 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19692), .ZN(n18443) );
  INV_X1 U16705 ( .A(n19045), .ZN(n13332) );
  NAND2_X1 U16706 ( .A1(n19656), .A2(n19692), .ZN(n19695) );
  INV_X1 U16707 ( .A(n19671), .ZN(n19658) );
  INV_X1 U16708 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n17422) );
  NOR3_X1 U16709 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n17422), .ZN(n19108) );
  NAND2_X1 U16710 ( .A1(n13333), .A2(n18561), .ZN(n17258) );
  XOR2_X1 U16711 ( .A(n13330), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n13334) );
  NOR2_X1 U16712 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18441), .ZN(
        n17271) );
  INV_X1 U16713 ( .A(n9749), .ZN(n17423) );
  INV_X1 U16714 ( .A(n18443), .ZN(n18720) );
  OR2_X1 U16715 ( .A1(n19335), .A2(n13333), .ZN(n17275) );
  OAI211_X1 U16716 ( .C1(n17423), .C2(n18720), .A(n9585), .B(n17275), .ZN(
        n17278) );
  NOR2_X1 U16717 ( .A1(n17271), .A2(n17278), .ZN(n17257) );
  OAI22_X1 U16718 ( .A1(n17258), .A2(n13334), .B1(n17257), .B2(n13330), .ZN(
        n13335) );
  AOI211_X1 U16719 ( .C1(n18578), .C2(n17436), .A(n13369), .B(n13335), .ZN(
        n13343) );
  INV_X1 U16720 ( .A(n13336), .ZN(n18847) );
  INV_X1 U16721 ( .A(n13338), .ZN(n13367) );
  INV_X1 U16722 ( .A(n17136), .ZN(n13340) );
  NAND2_X1 U16723 ( .A1(n13339), .A2(n18860), .ZN(n18405) );
  NAND2_X1 U16724 ( .A1(n13340), .A2(n18733), .ZN(n17260) );
  OAI21_X1 U16725 ( .B1(n21367), .B2(n17260), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13341) );
  OAI21_X1 U16726 ( .B1(n18532), .B2(n13367), .A(n13341), .ZN(n13373) );
  NAND2_X1 U16727 ( .A1(n13373), .A2(n18636), .ZN(n13342) );
  AND2_X1 U16728 ( .A1(n13343), .A2(n13342), .ZN(n13344) );
  NAND2_X1 U16729 ( .A1(n13347), .A2(n13346), .ZN(P3_U2799) );
  AOI221_X1 U16730 ( .B1(n13350), .B2(n17400), .C1(n13349), .C2(n17400), .A(
        n13348), .ZN(n17066) );
  NOR2_X1 U16731 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n17397) );
  INV_X1 U16732 ( .A(n17397), .ZN(n19560) );
  OAI21_X1 U16733 ( .B1(n19062), .B2(n19691), .A(n13358), .ZN(n13351) );
  NAND2_X1 U16734 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19702) );
  OAI21_X1 U16735 ( .B1(n19690), .B2(n13351), .A(n19702), .ZN(n17398) );
  NOR2_X1 U16736 ( .A1(n19523), .A2(n17398), .ZN(n13353) );
  MUX2_X1 U16737 ( .A(n19529), .B(n13353), .S(n13352), .Z(n13354) );
  AOI21_X1 U16738 ( .B1(n13356), .B2(n13355), .A(n13354), .ZN(n13357) );
  AOI21_X2 U16739 ( .B1(n17066), .B2(n13357), .A(n19547), .ZN(n19037) );
  NAND2_X1 U16740 ( .A1(n19037), .A2(n18851), .ZN(n18994) );
  AOI21_X1 U16741 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18993) );
  NAND3_X1 U16742 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18966) );
  NOR2_X1 U16743 ( .A1(n18993), .A2(n18966), .ZN(n18949) );
  INV_X1 U16744 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18957) );
  NAND2_X1 U16745 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18948) );
  NOR2_X1 U16746 ( .A1(n18957), .A2(n18948), .ZN(n18826) );
  NAND2_X1 U16747 ( .A1(n18949), .A2(n18826), .ZN(n18846) );
  NOR2_X1 U16748 ( .A1(n18780), .A2(n18846), .ZN(n13366) );
  INV_X1 U16749 ( .A(n19512), .ZN(n19528) );
  NOR2_X1 U16750 ( .A1(n13366), .A2(n19528), .ZN(n18828) );
  AOI21_X1 U16751 ( .B1(n19512), .B2(n18726), .A(n18828), .ZN(n18728) );
  NOR2_X1 U16752 ( .A1(n19674), .A2(n18734), .ZN(n13362) );
  INV_X1 U16753 ( .A(n18826), .ZN(n18861) );
  OR3_X1 U16754 ( .A1(n21354), .A2(n13072), .A3(n18966), .ZN(n18952) );
  NOR2_X1 U16755 ( .A1(n18861), .A2(n18952), .ZN(n18888) );
  NAND2_X1 U16756 ( .A1(n9603), .A2(n18888), .ZN(n18727) );
  NOR2_X1 U16757 ( .A1(n17262), .A2(n18727), .ZN(n13361) );
  OAI21_X1 U16758 ( .B1(n19494), .B2(n13362), .A(n13361), .ZN(n13363) );
  OAI21_X1 U16759 ( .B1(n19032), .B2(n19499), .A(n13363), .ZN(n13365) );
  OAI21_X1 U16760 ( .B1(n18729), .B2(n18730), .A(n19512), .ZN(n13364) );
  NAND3_X1 U16761 ( .A1(n18728), .A2(n13365), .A3(n13364), .ZN(n17074) );
  INV_X1 U16762 ( .A(n18994), .ZN(n19031) );
  AOI22_X1 U16763 ( .A1(n19037), .A2(n17074), .B1(n19031), .B2(n17136), .ZN(
        n17138) );
  OAI211_X1 U16764 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n18994), .A(
        n17138), .B(n19027), .ZN(n13370) );
  INV_X1 U16765 ( .A(n18727), .ZN(n18784) );
  OAI21_X1 U16766 ( .B1(n19494), .B2(n19674), .A(n19501), .ZN(n19016) );
  AOI22_X1 U16767 ( .A1(n19512), .A2(n13366), .B1(n18784), .B2(n19016), .ZN(
        n18749) );
  NOR3_X1 U16768 ( .A1(n18749), .A2(n19026), .A3(n13367), .ZN(n13368) );
  AOI211_X1 U16769 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n13370), .A(
        n13369), .B(n13368), .ZN(n13371) );
  AOI21_X1 U16770 ( .B1(n13373), .B2(n18961), .A(n13372), .ZN(n13374) );
  NAND2_X1 U16771 ( .A1(n13377), .A2(n13376), .ZN(P3_U2831) );
  NOR2_X1 U16772 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13379) );
  NOR4_X1 U16773 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13378) );
  NAND4_X1 U16774 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13379), .A4(n13378), .ZN(n13391) );
  INV_X1 U16775 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21304) );
  NOR3_X1 U16776 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n21304), .ZN(n13381) );
  NOR4_X1 U16777 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13380) );
  NAND4_X1 U16778 ( .A1(n15085), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13381), .A4(
        n13380), .ZN(U214) );
  NOR4_X1 U16779 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13385) );
  NOR4_X1 U16780 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n13384) );
  NOR4_X1 U16781 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13383) );
  NOR4_X1 U16782 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13382) );
  NAND4_X1 U16783 ( .A1(n13385), .A2(n13384), .A3(n13383), .A4(n13382), .ZN(
        n13390) );
  NOR4_X1 U16784 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n13388) );
  NOR4_X1 U16785 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(
        P2_ADDRESS_REG_23__SCAN_IN), .A3(P2_ADDRESS_REG_22__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n13387) );
  NOR4_X1 U16786 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n13386) );
  INV_X1 U16787 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20570) );
  NAND4_X1 U16788 ( .A1(n13388), .A2(n13387), .A3(n13386), .A4(n20570), .ZN(
        n13389) );
  NOR2_X1 U16789 ( .A1(n16872), .A2(n13391), .ZN(n17302) );
  NAND2_X1 U16790 ( .A1(n17302), .A2(U214), .ZN(U212) );
  AND2_X1 U16791 ( .A1(n20463), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20536) );
  NAND2_X1 U16792 ( .A1(n20539), .A2(n20536), .ZN(n17248) );
  INV_X1 U16793 ( .A(n17248), .ZN(n13394) );
  NOR2_X1 U16794 ( .A1(n16825), .A2(n20463), .ZN(n13544) );
  NAND2_X1 U16795 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13544), .ZN(n17143) );
  INV_X1 U16796 ( .A(n17143), .ZN(n13479) );
  NOR3_X1 U16797 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(P2_STATE2_REG_0__SCAN_IN), .ZN(n13393) );
  NOR2_X1 U16798 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13392) );
  NOR4_X1 U16799 ( .A1(n13394), .A2(n13479), .A3(n13393), .A4(n13392), .ZN(
        P2_U3178) );
  INV_X1 U16800 ( .A(n20689), .ZN(n13396) );
  NOR2_X1 U16801 ( .A1(n20628), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19719) );
  OAI21_X1 U16802 ( .B1(P2_READREQUEST_REG_SCAN_IN), .B2(n19719), .A(n20682), 
        .ZN(n13395) );
  OAI21_X1 U16803 ( .B1(n13396), .B2(n20682), .A(n13395), .ZN(P2_U3612) );
  INV_X1 U16804 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13398) );
  NAND3_X1 U16805 ( .A1(n19715), .A2(n20686), .A3(n19972), .ZN(n13399) );
  AOI22_X1 U16806 ( .A1(n16873), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16872), .ZN(n16269) );
  INV_X1 U16807 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13397) );
  OAI21_X1 U16808 ( .B1(n20688), .B2(n20686), .A(n19715), .ZN(n13442) );
  INV_X1 U16809 ( .A(n13442), .ZN(n13402) );
  OAI222_X1 U16810 ( .A1(n13490), .A2(n13398), .B1(n13399), .B2(n16269), .C1(
        n13397), .C2(n13402), .ZN(P2_U2982) );
  INV_X1 U16811 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13498) );
  INV_X1 U16812 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n17339) );
  OR2_X1 U16813 ( .A1(n14164), .A2(n17339), .ZN(n13401) );
  NAND2_X1 U16814 ( .A1(n16872), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13400) );
  NAND2_X1 U16815 ( .A1(n13401), .A2(n13400), .ZN(n16197) );
  NAND2_X1 U16816 ( .A1(n19935), .A2(n16197), .ZN(n13408) );
  NAND2_X1 U16817 ( .A1(n19937), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13403) );
  OAI211_X1 U16818 ( .C1(n13498), .C2(n13490), .A(n13408), .B(n13403), .ZN(
        P2_U2960) );
  INV_X1 U16819 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13507) );
  INV_X1 U16820 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n21401) );
  OR2_X1 U16821 ( .A1(n16872), .A2(n21401), .ZN(n13405) );
  NAND2_X1 U16822 ( .A1(n16872), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13404) );
  NAND2_X1 U16823 ( .A1(n13405), .A2(n13404), .ZN(n16181) );
  NAND2_X1 U16824 ( .A1(n19935), .A2(n16181), .ZN(n13413) );
  NAND2_X1 U16825 ( .A1(n19937), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13406) );
  OAI211_X1 U16826 ( .C1(n13507), .C2(n13490), .A(n13413), .B(n13406), .ZN(
        P2_U2962) );
  INV_X1 U16827 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19917) );
  NAND2_X1 U16828 ( .A1(n19937), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13407) );
  OAI211_X1 U16829 ( .C1(n19917), .C2(n13490), .A(n13408), .B(n13407), .ZN(
        P2_U2975) );
  INV_X1 U16830 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19915) );
  INV_X1 U16831 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n17337) );
  OR2_X1 U16832 ( .A1(n16872), .A2(n17337), .ZN(n13410) );
  NAND2_X1 U16833 ( .A1(n16872), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13409) );
  NAND2_X1 U16834 ( .A1(n13410), .A2(n13409), .ZN(n16190) );
  NAND2_X1 U16835 ( .A1(n19935), .A2(n16190), .ZN(n13451) );
  NAND2_X1 U16836 ( .A1(n19937), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13411) );
  OAI211_X1 U16837 ( .C1(n19915), .C2(n13490), .A(n13451), .B(n13411), .ZN(
        P2_U2976) );
  INV_X1 U16838 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19913) );
  NAND2_X1 U16839 ( .A1(n19937), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13412) );
  OAI211_X1 U16840 ( .C1(n19913), .C2(n13490), .A(n13413), .B(n13412), .ZN(
        P2_U2977) );
  INV_X1 U16841 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13501) );
  INV_X1 U16842 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n17333) );
  OR2_X1 U16843 ( .A1(n16872), .A2(n17333), .ZN(n13415) );
  NAND2_X1 U16844 ( .A1(n16872), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13414) );
  NAND2_X1 U16845 ( .A1(n13415), .A2(n13414), .ZN(n16167) );
  NAND2_X1 U16846 ( .A1(n19935), .A2(n16167), .ZN(n13418) );
  NAND2_X1 U16847 ( .A1(n19937), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13416) );
  OAI211_X1 U16848 ( .C1(n13501), .C2(n13490), .A(n13418), .B(n13416), .ZN(
        P2_U2964) );
  INV_X1 U16849 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19909) );
  NAND2_X1 U16850 ( .A1(n19937), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13417) );
  OAI211_X1 U16851 ( .C1(n19909), .C2(n13490), .A(n13418), .B(n13417), .ZN(
        P2_U2979) );
  AOI22_X1 U16852 ( .A1(n19938), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n13442), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13421) );
  NAND2_X1 U16853 ( .A1(n14164), .A2(BUF2_REG_2__SCAN_IN), .ZN(n13420) );
  INV_X1 U16854 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n17348) );
  OR2_X1 U16855 ( .A1(n16872), .A2(n17348), .ZN(n13419) );
  NAND2_X1 U16856 ( .A1(n13420), .A2(n13419), .ZN(n19977) );
  NAND2_X1 U16857 ( .A1(n19935), .A2(n19977), .ZN(n13434) );
  NAND2_X1 U16858 ( .A1(n13421), .A2(n13434), .ZN(P2_U2954) );
  AOI22_X1 U16859 ( .A1(n19938), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n13442), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13425) );
  INV_X1 U16860 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13422) );
  OR2_X1 U16861 ( .A1(n14164), .A2(n13422), .ZN(n13424) );
  NAND2_X1 U16862 ( .A1(n14164), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13423) );
  NAND2_X1 U16863 ( .A1(n13424), .A2(n13423), .ZN(n16175) );
  NAND2_X1 U16864 ( .A1(n19935), .A2(n16175), .ZN(n13445) );
  NAND2_X1 U16865 ( .A1(n13425), .A2(n13445), .ZN(P2_U2963) );
  AOI22_X1 U16866 ( .A1(n19938), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n13442), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13429) );
  INV_X1 U16867 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13426) );
  OR2_X1 U16868 ( .A1(n16872), .A2(n13426), .ZN(n13428) );
  NAND2_X1 U16869 ( .A1(n16872), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13427) );
  NAND2_X1 U16870 ( .A1(n13428), .A2(n13427), .ZN(n16159) );
  NAND2_X1 U16871 ( .A1(n19935), .A2(n16159), .ZN(n13443) );
  NAND2_X1 U16872 ( .A1(n13429), .A2(n13443), .ZN(P2_U2965) );
  AOI22_X1 U16873 ( .A1(n19938), .A2(P2_EAX_REG_0__SCAN_IN), .B1(n13442), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n13432) );
  NAND2_X1 U16874 ( .A1(n14164), .A2(BUF2_REG_0__SCAN_IN), .ZN(n13431) );
  INV_X1 U16875 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n17355) );
  OR2_X1 U16876 ( .A1(n16872), .A2(n17355), .ZN(n13430) );
  NAND2_X1 U16877 ( .A1(n13431), .A2(n13430), .ZN(n16881) );
  NAND2_X1 U16878 ( .A1(n19935), .A2(n16881), .ZN(n13447) );
  NAND2_X1 U16879 ( .A1(n13432), .A2(n13447), .ZN(P2_U2967) );
  AOI22_X1 U16880 ( .A1(n19938), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n13442), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13433) );
  AOI22_X1 U16881 ( .A1(n16873), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16872), .ZN(n19897) );
  INV_X1 U16882 ( .A(n19897), .ZN(n19973) );
  NAND2_X1 U16883 ( .A1(n19935), .A2(n19973), .ZN(n13449) );
  NAND2_X1 U16884 ( .A1(n13433), .A2(n13449), .ZN(P2_U2968) );
  AOI22_X1 U16885 ( .A1(n19938), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n13442), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13435) );
  NAND2_X1 U16886 ( .A1(n13435), .A2(n13434), .ZN(P2_U2969) );
  AOI22_X1 U16887 ( .A1(n19938), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n13442), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13436) );
  AOI22_X1 U16888 ( .A1(n16873), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16872), .ZN(n19886) );
  INV_X1 U16889 ( .A(n19886), .ZN(n16913) );
  NAND2_X1 U16890 ( .A1(n19935), .A2(n16913), .ZN(n13466) );
  NAND2_X1 U16891 ( .A1(n13436), .A2(n13466), .ZN(P2_U2970) );
  AOI22_X1 U16892 ( .A1(n19938), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n13442), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n13439) );
  NAND2_X1 U16893 ( .A1(n14164), .A2(BUF2_REG_4__SCAN_IN), .ZN(n13438) );
  INV_X1 U16894 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n17344) );
  OR2_X1 U16895 ( .A1(n14164), .A2(n17344), .ZN(n13437) );
  NAND2_X1 U16896 ( .A1(n13438), .A2(n13437), .ZN(n19985) );
  NAND2_X1 U16897 ( .A1(n19935), .A2(n19985), .ZN(n13440) );
  NAND2_X1 U16898 ( .A1(n13439), .A2(n13440), .ZN(P2_U2971) );
  AOI22_X1 U16899 ( .A1(n19938), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n13442), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13441) );
  NAND2_X1 U16900 ( .A1(n13441), .A2(n13440), .ZN(P2_U2956) );
  AOI22_X1 U16901 ( .A1(n19938), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n13442), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13444) );
  NAND2_X1 U16902 ( .A1(n13444), .A2(n13443), .ZN(P2_U2980) );
  AOI22_X1 U16903 ( .A1(n19938), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n19937), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13446) );
  NAND2_X1 U16904 ( .A1(n13446), .A2(n13445), .ZN(P2_U2978) );
  AOI22_X1 U16905 ( .A1(n19938), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n19937), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13448) );
  NAND2_X1 U16906 ( .A1(n13448), .A2(n13447), .ZN(P2_U2952) );
  AOI22_X1 U16907 ( .A1(n19938), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n19937), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13450) );
  NAND2_X1 U16908 ( .A1(n13450), .A2(n13449), .ZN(P2_U2953) );
  AOI22_X1 U16909 ( .A1(n19938), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n19937), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13452) );
  NAND2_X1 U16910 ( .A1(n13452), .A2(n13451), .ZN(P2_U2961) );
  AOI22_X1 U16911 ( .A1(n19938), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n19937), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n13455) );
  NAND2_X1 U16912 ( .A1(n14164), .A2(BUF2_REG_6__SCAN_IN), .ZN(n13454) );
  INV_X1 U16913 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n21338) );
  OR2_X1 U16914 ( .A1(n14164), .A2(n21338), .ZN(n13453) );
  NAND2_X1 U16915 ( .A1(n13454), .A2(n13453), .ZN(n19994) );
  NAND2_X1 U16916 ( .A1(n19935), .A2(n19994), .ZN(n13462) );
  NAND2_X1 U16917 ( .A1(n13455), .A2(n13462), .ZN(P2_U2973) );
  AOI22_X1 U16918 ( .A1(n19938), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n19937), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n13459) );
  NAND2_X1 U16919 ( .A1(n14164), .A2(BUF2_REG_7__SCAN_IN), .ZN(n13458) );
  INV_X1 U16920 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n13456) );
  OR2_X1 U16921 ( .A1(n14164), .A2(n13456), .ZN(n13457) );
  NAND2_X1 U16922 ( .A1(n13458), .A2(n13457), .ZN(n20000) );
  NAND2_X1 U16923 ( .A1(n19935), .A2(n20000), .ZN(n13460) );
  NAND2_X1 U16924 ( .A1(n13459), .A2(n13460), .ZN(P2_U2974) );
  AOI22_X1 U16925 ( .A1(n19938), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n19937), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13461) );
  NAND2_X1 U16926 ( .A1(n13461), .A2(n13460), .ZN(P2_U2959) );
  AOI22_X1 U16927 ( .A1(n19938), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n19937), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13463) );
  NAND2_X1 U16928 ( .A1(n13463), .A2(n13462), .ZN(P2_U2958) );
  AOI22_X1 U16929 ( .A1(n19938), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n19937), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13465) );
  AOI22_X1 U16930 ( .A1(n16873), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16872), .ZN(n13464) );
  INV_X1 U16931 ( .A(n13464), .ZN(n19990) );
  NAND2_X1 U16932 ( .A1(n19935), .A2(n19990), .ZN(n13468) );
  NAND2_X1 U16933 ( .A1(n13465), .A2(n13468), .ZN(P2_U2957) );
  AOI22_X1 U16934 ( .A1(n19938), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n19937), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13467) );
  NAND2_X1 U16935 ( .A1(n13467), .A2(n13466), .ZN(P2_U2955) );
  AOI22_X1 U16936 ( .A1(n19938), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n19937), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n13469) );
  NAND2_X1 U16937 ( .A1(n13469), .A2(n13468), .ZN(P2_U2972) );
  NAND2_X1 U16938 ( .A1(n16926), .A2(n16925), .ZN(n13472) );
  INV_X1 U16939 ( .A(n16934), .ZN(n16923) );
  NAND2_X1 U16940 ( .A1(n20689), .A2(n20686), .ZN(n16932) );
  INV_X1 U16941 ( .A(n16931), .ZN(n16922) );
  NOR2_X1 U16942 ( .A1(n16932), .A2(n16922), .ZN(n13470) );
  NAND2_X1 U16943 ( .A1(n16923), .A2(n13470), .ZN(n13471) );
  NAND2_X1 U16944 ( .A1(n13472), .A2(n13471), .ZN(n13572) );
  INV_X1 U16945 ( .A(n13572), .ZN(n13478) );
  INV_X1 U16946 ( .A(n16925), .ZN(n16927) );
  NAND2_X1 U16947 ( .A1(n16927), .A2(n16924), .ZN(n13588) );
  NAND3_X1 U16948 ( .A1(n13489), .A2(n13475), .A3(n13474), .ZN(n13476) );
  NAND4_X1 U16949 ( .A1(n13478), .A2(n13477), .A3(n13588), .A4(n13476), .ZN(
        n16936) );
  NAND2_X1 U16950 ( .A1(n16936), .A2(n20542), .ZN(n13482) );
  NAND2_X1 U16951 ( .A1(n20690), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16965) );
  NAND2_X1 U16952 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(n13479), .ZN(n13480) );
  AND2_X1 U16953 ( .A1(n16965), .A2(n13480), .ZN(n13481) );
  NAND2_X1 U16954 ( .A1(n13482), .A2(n13481), .ZN(n16865) );
  INV_X1 U16955 ( .A(n13483), .ZN(n13484) );
  INV_X1 U16956 ( .A(n16951), .ZN(n13486) );
  NOR2_X1 U16957 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20631) );
  NAND3_X1 U16958 ( .A1(n16865), .A2(n13486), .A3(n20631), .ZN(n13487) );
  OAI21_X1 U16959 ( .B1(n16865), .B2(n16921), .A(n13487), .ZN(P2_U3595) );
  INV_X1 U16960 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n13496) );
  NAND2_X1 U16961 ( .A1(n13489), .A2(n13488), .ZN(n13491) );
  NAND2_X1 U16962 ( .A1(n13491), .A2(n13490), .ZN(n13492) );
  NAND2_X1 U16963 ( .A1(n20690), .A2(n13544), .ZN(n13529) );
  INV_X1 U16964 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13495) );
  INV_X1 U16965 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n13494) );
  OAI222_X1 U16966 ( .A1(n13496), .A2(n19902), .B1(n13528), .B2(n13495), .C1(
        n13529), .C2(n13494), .ZN(P2_U2933) );
  INV_X1 U16967 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n13499) );
  INV_X1 U16968 ( .A(P2_UWORD_REG_8__SCAN_IN), .ZN(n13497) );
  OAI222_X1 U16969 ( .A1(n13499), .A2(n19902), .B1(n13528), .B2(n13498), .C1(
        n13529), .C2(n13497), .ZN(P2_U2927) );
  INV_X1 U16970 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13502) );
  INV_X1 U16971 ( .A(P2_UWORD_REG_12__SCAN_IN), .ZN(n13500) );
  OAI222_X1 U16972 ( .A1(n13502), .A2(n19902), .B1(n13528), .B2(n13501), .C1(
        n13529), .C2(n13500), .ZN(P2_U2923) );
  INV_X1 U16973 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n13505) );
  INV_X1 U16974 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13504) );
  INV_X1 U16975 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13503) );
  OAI222_X1 U16976 ( .A1(n13505), .A2(n19902), .B1(n13528), .B2(n13504), .C1(
        n13529), .C2(n13503), .ZN(P2_U2935) );
  INV_X1 U16977 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n13508) );
  INV_X1 U16978 ( .A(P2_UWORD_REG_10__SCAN_IN), .ZN(n13506) );
  OAI222_X1 U16979 ( .A1(n13508), .A2(n19902), .B1(n13528), .B2(n13507), .C1(
        n13529), .C2(n13506), .ZN(P2_U2925) );
  INV_X1 U16980 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n13511) );
  INV_X1 U16981 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13510) );
  INV_X1 U16982 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n13509) );
  OAI222_X1 U16983 ( .A1(n13511), .A2(n19902), .B1(n13528), .B2(n13510), .C1(
        n13529), .C2(n13509), .ZN(P2_U2929) );
  INV_X1 U16984 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n13514) );
  INV_X1 U16985 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13513) );
  INV_X1 U16986 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n13512) );
  OAI222_X1 U16987 ( .A1(n13514), .A2(n19902), .B1(n13528), .B2(n13513), .C1(
        n13529), .C2(n13512), .ZN(P2_U2931) );
  INV_X1 U16988 ( .A(n17215), .ZN(n21212) );
  NOR2_X1 U16989 ( .A1(n21212), .A2(n11830), .ZN(n13520) );
  AOI211_X1 U16990 ( .C1(n13516), .C2(n13520), .A(n21149), .B(n13515), .ZN(
        n13517) );
  AND2_X1 U16991 ( .A1(n14757), .A2(n13517), .ZN(n13525) );
  NOR2_X1 U16992 ( .A1(n13525), .A2(n17128), .ZN(n13527) );
  INV_X1 U16993 ( .A(n13518), .ZN(n13524) );
  OAI21_X1 U16994 ( .B1(n17142), .B2(n20709), .A(n13519), .ZN(n13521) );
  AOI21_X1 U16995 ( .B1(n13521), .B2(n13520), .A(n11759), .ZN(n13522) );
  AOI21_X1 U16996 ( .B1(n13524), .B2(n13523), .A(n13522), .ZN(n13526) );
  INV_X1 U16997 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21217) );
  AOI22_X1 U16998 ( .A1(n13527), .A2(n13526), .B1(n13525), .B2(n21217), .ZN(
        P1_U3485) );
  INV_X1 U16999 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n13531) );
  AOI22_X1 U17000 ( .A1(n19899), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n20685), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13530) );
  OAI21_X1 U17001 ( .B1(n19902), .B2(n13531), .A(n13530), .ZN(P2_U2932) );
  INV_X1 U17002 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n13533) );
  AOI22_X1 U17003 ( .A1(n19899), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n20685), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13532) );
  OAI21_X1 U17004 ( .B1(n19902), .B2(n13533), .A(n13532), .ZN(P2_U2926) );
  INV_X1 U17005 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n13535) );
  AOI22_X1 U17006 ( .A1(n19899), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n20685), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13534) );
  OAI21_X1 U17007 ( .B1(n19902), .B2(n13535), .A(n13534), .ZN(P2_U2924) );
  INV_X1 U17008 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n13537) );
  AOI22_X1 U17009 ( .A1(n19899), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n20685), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13536) );
  OAI21_X1 U17010 ( .B1(n19902), .B2(n13537), .A(n13536), .ZN(P2_U2928) );
  INV_X1 U17011 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n13539) );
  AOI22_X1 U17012 ( .A1(n19899), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n20685), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13538) );
  OAI21_X1 U17013 ( .B1(n19902), .B2(n13539), .A(n13538), .ZN(P2_U2922) );
  INV_X1 U17014 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n13541) );
  AOI22_X1 U17015 ( .A1(n19899), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n20685), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13540) );
  OAI21_X1 U17016 ( .B1(n19902), .B2(n13541), .A(n13540), .ZN(P2_U2934) );
  INV_X1 U17017 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n13543) );
  AOI22_X1 U17018 ( .A1(n19899), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n20685), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13542) );
  OAI21_X1 U17019 ( .B1(n19902), .B2(n13543), .A(n13542), .ZN(P2_U2930) );
  OAI21_X1 U17020 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_2__SCAN_IN), .A(n20690), .ZN(n20695) );
  INV_X1 U17021 ( .A(n19950), .ZN(n16547) );
  XNOR2_X1 U17022 ( .A(n13548), .B(n13547), .ZN(n13652) );
  NAND2_X1 U17023 ( .A1(n13550), .A2(n13549), .ZN(n19725) );
  OR2_X1 U17024 ( .A1(n20634), .A2(n20631), .ZN(n20663) );
  NAND2_X1 U17025 ( .A1(n20663), .A2(n20690), .ZN(n13551) );
  NAND2_X1 U17026 ( .A1(n20690), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16963) );
  NAND2_X1 U17027 ( .A1(n16963), .A2(n13552), .ZN(n14341) );
  NOR2_X1 U17028 ( .A1(n16491), .A2(n20569), .ZN(n13657) );
  INV_X1 U17029 ( .A(n13657), .ZN(n13553) );
  OAI21_X1 U17030 ( .B1(n19955), .B2(n16013), .A(n13553), .ZN(n13554) );
  AOI21_X1 U17031 ( .B1(n19943), .B2(n16016), .A(n13554), .ZN(n13559) );
  NOR2_X1 U17032 ( .A1(n13556), .A2(n13555), .ZN(n13644) );
  INV_X1 U17033 ( .A(n13644), .ZN(n13557) );
  OR2_X1 U17034 ( .A1(n19725), .A2(n20688), .ZN(n16483) );
  NAND3_X1 U17035 ( .A1(n13557), .A2(n10145), .A3(n13645), .ZN(n13558) );
  OAI211_X1 U17036 ( .C1(n13652), .C2(n16550), .A(n13559), .B(n13558), .ZN(
        n13560) );
  AOI21_X1 U17037 ( .B1(n13766), .B2(n16547), .A(n13560), .ZN(n13561) );
  INV_X1 U17038 ( .A(n13561), .ZN(P2_U3012) );
  INV_X1 U17039 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n21419) );
  AND2_X1 U17040 ( .A1(n13622), .A2(n21212), .ZN(n13562) );
  NAND2_X1 U17041 ( .A1(n13600), .A2(n13563), .ZN(n20842) );
  INV_X1 U17042 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13564) );
  NOR2_X1 U17043 ( .A1(n13803), .A2(n13564), .ZN(n13565) );
  AOI21_X1 U17044 ( .B1(DATAI_15_), .B2(n13803), .A(n13565), .ZN(n15151) );
  OAI222_X1 U17045 ( .A1(n20856), .A2(n20803), .B1(n21419), .B2(n13600), .C1(
        n20842), .C2(n15151), .ZN(P1_U2967) );
  INV_X1 U17046 ( .A(n13567), .ZN(n13568) );
  XNOR2_X1 U17047 ( .A(n13566), .B(n13568), .ZN(n16779) );
  INV_X1 U17048 ( .A(n16779), .ZN(n19869) );
  INV_X1 U17049 ( .A(n10792), .ZN(n13569) );
  NOR2_X1 U17050 ( .A1(n13570), .A2(n13569), .ZN(n13571) );
  NAND2_X1 U17051 ( .A1(n16287), .A2(n11292), .ZN(n16227) );
  INV_X1 U17052 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19921) );
  INV_X1 U17053 ( .A(n16260), .ZN(n13578) );
  INV_X1 U17054 ( .A(n13575), .ZN(n13576) );
  INV_X1 U17055 ( .A(n14694), .ZN(n13577) );
  INV_X1 U17056 ( .A(n19994), .ZN(n13579) );
  OAI222_X1 U17057 ( .A1(n19869), .A2(n16275), .B1(n19921), .B2(n16287), .C1(
        n19896), .C2(n13579), .ZN(P2_U2913) );
  INV_X1 U17058 ( .A(n14344), .ZN(n13581) );
  INV_X1 U17059 ( .A(n16963), .ZN(n13580) );
  NAND2_X1 U17060 ( .A1(n13581), .A2(n13580), .ZN(n13584) );
  NAND2_X1 U17061 ( .A1(n10794), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13582) );
  AOI22_X1 U17062 ( .A1(n13865), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20634), .B2(n20667), .ZN(n13583) );
  NAND2_X1 U17063 ( .A1(n19972), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13586) );
  AND4_X1 U17064 ( .A1(n13585), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13586), 
        .A4(n20276), .ZN(n13587) );
  NAND2_X1 U17065 ( .A1(n13588), .A2(n9605), .ZN(n13589) );
  INV_X2 U17066 ( .A(n16104), .ZN(n16157) );
  NOR2_X1 U17067 ( .A1(n14344), .A2(n16157), .ZN(n13590) );
  AOI21_X1 U17068 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n16157), .A(n13590), .ZN(
        n13591) );
  OAI21_X1 U17069 ( .B1(n16907), .B2(n9716), .A(n13591), .ZN(P2_U2887) );
  OAI21_X1 U17070 ( .B1(n13592), .B2(n13595), .A(n13594), .ZN(n19852) );
  INV_X1 U17071 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19919) );
  INV_X1 U17072 ( .A(n20000), .ZN(n13596) );
  OAI222_X1 U17073 ( .A1(n19852), .A2(n16275), .B1(n19919), .B2(n16287), .C1(
        n19896), .C2(n13596), .ZN(P2_U2912) );
  NAND2_X1 U17074 ( .A1(n13803), .A2(DATAI_0_), .ZN(n13598) );
  NAND2_X1 U17075 ( .A1(n15085), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13597) );
  AND2_X1 U17076 ( .A1(n13598), .A2(n13597), .ZN(n15143) );
  INV_X1 U17077 ( .A(n15143), .ZN(n13599) );
  NAND2_X1 U17078 ( .A1(n13729), .A2(n13599), .ZN(n13732) );
  NAND2_X1 U17079 ( .A1(n13702), .A2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13601) );
  OAI211_X1 U17080 ( .C1(n20856), .C2(n15142), .A(n13732), .B(n13601), .ZN(
        P1_U2937) );
  INV_X1 U17081 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13603) );
  NAND2_X1 U17082 ( .A1(n20660), .A2(n20667), .ZN(n20212) );
  INV_X1 U17083 ( .A(n20212), .ZN(n13604) );
  NOR2_X1 U17084 ( .A1(n20313), .A2(n13604), .ZN(n20149) );
  AND2_X1 U17085 ( .A1(n20149), .A2(n20634), .ZN(n20282) );
  AOI21_X1 U17086 ( .B1(n13865), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n20282), .ZN(n13605) );
  OAI21_X1 U17087 ( .B1(n13606), .B2(n16963), .A(n13605), .ZN(n13770) );
  MUX2_X1 U17088 ( .A(n10819), .B(n16831), .S(n16104), .Z(n13608) );
  OAI21_X1 U17089 ( .B1(n20655), .B2(n9716), .A(n13608), .ZN(P2_U2886) );
  INV_X1 U17090 ( .A(n16881), .ZN(n13617) );
  INV_X1 U17091 ( .A(n13609), .ZN(n13612) );
  INV_X1 U17092 ( .A(n13610), .ZN(n13611) );
  NAND2_X1 U17093 ( .A1(n13612), .A2(n13611), .ZN(n13614) );
  AND2_X1 U17094 ( .A1(n13614), .A2(n13613), .ZN(n17235) );
  NAND2_X1 U17095 ( .A1(n20664), .A2(n17235), .ZN(n19890) );
  OAI211_X1 U17096 ( .C1(n20664), .C2(n17235), .A(n19890), .B(n19892), .ZN(
        n13616) );
  AOI22_X1 U17097 ( .A1(n19888), .A2(n17235), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19887), .ZN(n13615) );
  OAI211_X1 U17098 ( .C1(n13617), .C2(n19896), .A(n13616), .B(n13615), .ZN(
        P2_U2919) );
  NAND4_X1 U17099 ( .A1(n12561), .A2(n9601), .A3(n17210), .A4(n9737), .ZN(
        n13619) );
  OR2_X1 U17100 ( .A1(n13620), .A2(n13619), .ZN(n15671) );
  INV_X1 U17101 ( .A(n15671), .ZN(n13630) );
  XNOR2_X1 U17102 ( .A(n13621), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13627) );
  AND2_X1 U17103 ( .A1(n13622), .A2(n15020), .ZN(n17106) );
  AND2_X1 U17104 ( .A1(n13623), .A2(n17106), .ZN(n15616) );
  NOR2_X1 U17105 ( .A1(n13624), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15617) );
  INV_X1 U17106 ( .A(n13625), .ZN(n15611) );
  NOR2_X1 U17107 ( .A1(n15617), .A2(n13625), .ZN(n13631) );
  INV_X1 U17108 ( .A(n13631), .ZN(n13626) );
  AOI22_X1 U17109 ( .A1(n17084), .A2(n13627), .B1(n15616), .B2(n13626), .ZN(
        n13629) );
  NAND3_X1 U17110 ( .A1(n13630), .A2(n15613), .A3(n13631), .ZN(n13628) );
  OAI211_X1 U17111 ( .C1(n13618), .C2(n13630), .A(n13629), .B(n13628), .ZN(
        n15630) );
  INV_X1 U17112 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13790) );
  NOR2_X1 U17113 ( .A1(n17222), .A2(n13790), .ZN(n15675) );
  AOI22_X1 U17114 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20913), .B2(n13019), .ZN(
        n15673) );
  INV_X1 U17115 ( .A(n13798), .ZN(n21290) );
  AOI222_X1 U17116 ( .A1(n15630), .A2(n21291), .B1(n15675), .B2(n15673), .C1(
        n13631), .C2(n21290), .ZN(n13643) );
  INV_X1 U17117 ( .A(n12561), .ZN(n13632) );
  OAI211_X1 U17118 ( .C1(n17084), .C2(n13632), .A(n17105), .B(n17215), .ZN(
        n13633) );
  INV_X1 U17119 ( .A(n13633), .ZN(n13634) );
  MUX2_X1 U17120 ( .A(n13634), .B(n17101), .S(n17107), .Z(n13639) );
  OAI21_X1 U17121 ( .B1(n15020), .B2(n13636), .A(n13635), .ZN(n13637) );
  NAND2_X1 U17122 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17218) );
  INV_X1 U17123 ( .A(n17218), .ZN(n13799) );
  NAND2_X1 U17124 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13799), .ZN(n17223) );
  INV_X1 U17125 ( .A(n17223), .ZN(n15644) );
  AND2_X1 U17126 ( .A1(n15644), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n13640) );
  AOI21_X1 U17127 ( .B1(n15635), .B2(n9905), .A(n13640), .ZN(n17212) );
  OAI21_X1 U17128 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n21064), .A(n17212), 
        .ZN(n21294) );
  INV_X1 U17129 ( .A(n21294), .ZN(n13642) );
  NAND2_X1 U17130 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n13642), .ZN(
        n13641) );
  OAI21_X1 U17131 ( .B1(n13643), .B2(n13642), .A(n13641), .ZN(P1_U3472) );
  NOR2_X1 U17132 ( .A1(n16802), .A2(n13644), .ZN(n13646) );
  AOI22_X1 U17133 ( .A1(n13646), .A2(n13645), .B1(n17241), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13662) );
  OR2_X1 U17134 ( .A1(n13648), .A2(n13647), .ZN(n13649) );
  NAND2_X1 U17135 ( .A1(n13650), .A2(n13649), .ZN(n20645) );
  INV_X1 U17136 ( .A(n13651), .ZN(n13653) );
  OAI22_X1 U17137 ( .A1(n13654), .A2(n13653), .B1(n19970), .B2(n13652), .ZN(
        n13655) );
  NOR3_X1 U17138 ( .A1(n13657), .A2(n13656), .A3(n13655), .ZN(n13658) );
  OAI21_X1 U17139 ( .B1(n14712), .B2(n13659), .A(n13658), .ZN(n13660) );
  AOI21_X1 U17140 ( .B1(n19956), .B2(n20645), .A(n13660), .ZN(n13661) );
  OAI211_X1 U17141 ( .C1(n10868), .C2(n16782), .A(n13662), .B(n13661), .ZN(
        P2_U3044) );
  AOI22_X1 U17142 ( .A1(n15641), .A2(n15671), .B1(n13663), .B2(n13664), .ZN(
        n17082) );
  AOI22_X1 U17143 ( .A1(n21290), .A2(n13664), .B1(n13790), .B2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n13665) );
  OAI21_X1 U17144 ( .B1(n17082), .B2(n17211), .A(n13665), .ZN(n13667) );
  INV_X1 U17145 ( .A(n17084), .ZN(n15669) );
  OAI21_X1 U17146 ( .B1(n15669), .B2(n17211), .A(n21294), .ZN(n13666) );
  AOI22_X1 U17147 ( .A1(n13667), .A2(n21294), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13666), .ZN(n13668) );
  INV_X1 U17148 ( .A(n13668), .ZN(P1_U3474) );
  XNOR2_X1 U17149 ( .A(n13670), .B(n13669), .ZN(n15041) );
  NAND2_X1 U17150 ( .A1(n15301), .A2(n13671), .ZN(n13675) );
  OAI21_X1 U17151 ( .B1(n13673), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13672), .ZN(n20932) );
  NAND2_X1 U17152 ( .A1(n20916), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20937) );
  OAI21_X1 U17153 ( .B1(n20712), .B2(n20932), .A(n20937), .ZN(n13674) );
  AOI21_X1 U17154 ( .B1(n13675), .B2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n13674), .ZN(n13676) );
  OAI21_X1 U17155 ( .B1(n15041), .B2(n15382), .A(n13676), .ZN(P1_U2999) );
  INV_X1 U17156 ( .A(n13677), .ZN(n13678) );
  AOI21_X1 U17157 ( .B1(n13679), .B2(n13594), .A(n13678), .ZN(n16754) );
  INV_X1 U17158 ( .A(n16754), .ZN(n13681) );
  AOI22_X1 U17159 ( .A1(n16279), .A2(n16197), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n19887), .ZN(n13680) );
  OAI21_X1 U17160 ( .B1(n13681), .B2(n16275), .A(n13680), .ZN(P2_U2911) );
  NAND2_X1 U17161 ( .A1(n13803), .A2(DATAI_4_), .ZN(n13683) );
  NAND2_X1 U17162 ( .A1(n15085), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13682) );
  AND2_X1 U17163 ( .A1(n13683), .A2(n13682), .ZN(n15122) );
  INV_X1 U17164 ( .A(n15122), .ZN(n13684) );
  NAND2_X1 U17165 ( .A1(n13729), .A2(n13684), .ZN(n13719) );
  AOI22_X1 U17166 ( .A1(n13702), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_20__SCAN_IN), .ZN(n13685) );
  NAND2_X1 U17167 ( .A1(n13719), .A2(n13685), .ZN(P1_U2941) );
  NAND2_X1 U17168 ( .A1(n13803), .A2(DATAI_3_), .ZN(n13687) );
  NAND2_X1 U17169 ( .A1(n15085), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13686) );
  AND2_X1 U17170 ( .A1(n13687), .A2(n13686), .ZN(n15126) );
  INV_X1 U17171 ( .A(n15126), .ZN(n13688) );
  NAND2_X1 U17172 ( .A1(n13729), .A2(n13688), .ZN(n13717) );
  AOI22_X1 U17173 ( .A1(n13702), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_19__SCAN_IN), .ZN(n13689) );
  NAND2_X1 U17174 ( .A1(n13717), .A2(n13689), .ZN(P1_U2940) );
  INV_X1 U17175 ( .A(DATAI_1_), .ZN(n13691) );
  NAND2_X1 U17176 ( .A1(n15085), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13690) );
  OAI21_X1 U17177 ( .B1(n15085), .B2(n13691), .A(n13690), .ZN(n15135) );
  NAND2_X1 U17178 ( .A1(n13729), .A2(n15135), .ZN(n13711) );
  AOI22_X1 U17179 ( .A1(n13702), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_17__SCAN_IN), .ZN(n13692) );
  NAND2_X1 U17180 ( .A1(n13711), .A2(n13692), .ZN(P1_U2938) );
  NAND2_X1 U17181 ( .A1(n13803), .A2(DATAI_7_), .ZN(n13694) );
  NAND2_X1 U17182 ( .A1(n15085), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13693) );
  AND2_X1 U17183 ( .A1(n13694), .A2(n13693), .ZN(n15107) );
  INV_X1 U17184 ( .A(n15107), .ZN(n13695) );
  NAND2_X1 U17185 ( .A1(n13729), .A2(n13695), .ZN(n13723) );
  AOI22_X1 U17186 ( .A1(n13702), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_7__SCAN_IN), .ZN(n13696) );
  NAND2_X1 U17187 ( .A1(n13723), .A2(n13696), .ZN(P1_U2959) );
  INV_X1 U17188 ( .A(DATAI_8_), .ZN(n13697) );
  MUX2_X1 U17189 ( .A(n13697), .B(n17339), .S(n15085), .Z(n15103) );
  INV_X1 U17190 ( .A(n15103), .ZN(n13698) );
  NAND2_X1 U17191 ( .A1(n13729), .A2(n13698), .ZN(n13709) );
  AOI22_X1 U17192 ( .A1(n13702), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_8__SCAN_IN), .ZN(n13699) );
  NAND2_X1 U17193 ( .A1(n13709), .A2(n13699), .ZN(P1_U2960) );
  INV_X1 U17194 ( .A(DATAI_11_), .ZN(n13701) );
  NAND2_X1 U17195 ( .A1(n15085), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13700) );
  OAI21_X1 U17196 ( .B1(n15085), .B2(n13701), .A(n13700), .ZN(n15160) );
  NAND2_X1 U17197 ( .A1(n13729), .A2(n15160), .ZN(n13737) );
  AOI22_X1 U17198 ( .A1(n13702), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_27__SCAN_IN), .ZN(n13703) );
  NAND2_X1 U17199 ( .A1(n13737), .A2(n13703), .ZN(P1_U2948) );
  NAND2_X1 U17200 ( .A1(n13803), .A2(DATAI_5_), .ZN(n13705) );
  NAND2_X1 U17201 ( .A1(n15085), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13704) );
  AND2_X1 U17202 ( .A1(n13705), .A2(n13704), .ZN(n15117) );
  INV_X1 U17203 ( .A(n15117), .ZN(n13706) );
  NAND2_X1 U17204 ( .A1(n13729), .A2(n13706), .ZN(n13725) );
  AOI22_X1 U17205 ( .A1(n13702), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_5__SCAN_IN), .ZN(n13707) );
  NAND2_X1 U17206 ( .A1(n13725), .A2(n13707), .ZN(P1_U2957) );
  AOI22_X1 U17207 ( .A1(n13702), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_24__SCAN_IN), .ZN(n13708) );
  NAND2_X1 U17208 ( .A1(n13709), .A2(n13708), .ZN(P1_U2945) );
  AOI22_X1 U17209 ( .A1(n13702), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_1__SCAN_IN), .ZN(n13710) );
  NAND2_X1 U17210 ( .A1(n13711), .A2(n13710), .ZN(P1_U2953) );
  NAND2_X1 U17211 ( .A1(n13803), .A2(DATAI_6_), .ZN(n13713) );
  NAND2_X1 U17212 ( .A1(n15085), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13712) );
  AND2_X1 U17213 ( .A1(n13713), .A2(n13712), .ZN(n15112) );
  INV_X1 U17214 ( .A(n15112), .ZN(n13714) );
  NAND2_X1 U17215 ( .A1(n13729), .A2(n13714), .ZN(n13721) );
  AOI22_X1 U17216 ( .A1(n13702), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_22__SCAN_IN), .ZN(n13715) );
  NAND2_X1 U17217 ( .A1(n13721), .A2(n13715), .ZN(P1_U2943) );
  AOI22_X1 U17218 ( .A1(n13702), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_3__SCAN_IN), .ZN(n13716) );
  NAND2_X1 U17219 ( .A1(n13717), .A2(n13716), .ZN(P1_U2955) );
  AOI22_X1 U17220 ( .A1(n13702), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_4__SCAN_IN), .ZN(n13718) );
  NAND2_X1 U17221 ( .A1(n13719), .A2(n13718), .ZN(P1_U2956) );
  AOI22_X1 U17222 ( .A1(n13702), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_6__SCAN_IN), .ZN(n13720) );
  NAND2_X1 U17223 ( .A1(n13721), .A2(n13720), .ZN(P1_U2958) );
  AOI22_X1 U17224 ( .A1(n13702), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_23__SCAN_IN), .ZN(n13722) );
  NAND2_X1 U17225 ( .A1(n13723), .A2(n13722), .ZN(P1_U2944) );
  AOI22_X1 U17226 ( .A1(n13702), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_21__SCAN_IN), .ZN(n13724) );
  NAND2_X1 U17227 ( .A1(n13725), .A2(n13724), .ZN(P1_U2942) );
  NAND2_X1 U17228 ( .A1(n13803), .A2(DATAI_2_), .ZN(n13727) );
  NAND2_X1 U17229 ( .A1(n15085), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13726) );
  AND2_X1 U17230 ( .A1(n13727), .A2(n13726), .ZN(n15131) );
  INV_X1 U17231 ( .A(n15131), .ZN(n13728) );
  NAND2_X1 U17232 ( .A1(n13729), .A2(n13728), .ZN(n13734) );
  AOI22_X1 U17233 ( .A1(n13702), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_2__SCAN_IN), .ZN(n13730) );
  NAND2_X1 U17234 ( .A1(n13734), .A2(n13730), .ZN(P1_U2954) );
  AOI22_X1 U17235 ( .A1(n13702), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_0__SCAN_IN), .ZN(n13731) );
  NAND2_X1 U17236 ( .A1(n13732), .A2(n13731), .ZN(P1_U2952) );
  AOI22_X1 U17237 ( .A1(n13702), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_18__SCAN_IN), .ZN(n13733) );
  NAND2_X1 U17238 ( .A1(n13734), .A2(n13733), .ZN(P1_U2939) );
  AOI22_X1 U17239 ( .A1(n13702), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n13735), 
        .B2(P1_EAX_REG_11__SCAN_IN), .ZN(n13736) );
  NAND2_X1 U17240 ( .A1(n13737), .A2(n13736), .ZN(P1_U2963) );
  OAI21_X1 U17241 ( .B1(n13740), .B2(n13739), .A(n13738), .ZN(n20777) );
  NAND2_X1 U17242 ( .A1(n17107), .A2(n17101), .ZN(n13744) );
  OR2_X1 U17243 ( .A1(n13742), .A2(n13741), .ZN(n13743) );
  NAND2_X1 U17244 ( .A1(n13744), .A2(n13743), .ZN(n13745) );
  INV_X1 U17245 ( .A(n15070), .ZN(n20796) );
  OAI21_X1 U17246 ( .B1(n13748), .B2(n21470), .A(n13746), .ZN(n20778) );
  AOI22_X1 U17247 ( .A1(n20795), .A2(n20778), .B1(n15065), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13749) );
  OAI21_X1 U17248 ( .B1(n20777), .B2(n15067), .A(n13749), .ZN(P1_U2871) );
  NAND2_X1 U17249 ( .A1(n13750), .A2(n13790), .ZN(n13752) );
  NAND2_X1 U17250 ( .A1(n13752), .A2(n13751), .ZN(n20928) );
  INV_X1 U17251 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13753) );
  OAI222_X1 U17252 ( .A1(n20928), .A2(n15068), .B1(n15067), .B2(n15041), .C1(
        n13753), .C2(n20800), .ZN(P1_U2872) );
  INV_X1 U17253 ( .A(n13754), .ZN(n13755) );
  AOI21_X1 U17254 ( .B1(n13756), .B2(n13677), .A(n13755), .ZN(n16743) );
  INV_X1 U17255 ( .A(n16743), .ZN(n19839) );
  AOI22_X1 U17256 ( .A1(n16279), .A2(n16190), .B1(P2_EAX_REG_9__SCAN_IN), .B2(
        n19887), .ZN(n13757) );
  OAI21_X1 U17257 ( .B1(n19839), .B2(n16275), .A(n13757), .ZN(P2_U2910) );
  AND2_X1 U17258 ( .A1(n13808), .A2(n13758), .ZN(n13762) );
  INV_X1 U17259 ( .A(n13762), .ZN(n13759) );
  AND2_X1 U17260 ( .A1(n13760), .A2(n13759), .ZN(n13761) );
  NAND2_X1 U17261 ( .A1(n15144), .A2(n13763), .ZN(n15155) );
  INV_X1 U17262 ( .A(n15135), .ZN(n13828) );
  INV_X1 U17263 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20823) );
  OAI222_X1 U17264 ( .A1(n15163), .A2(n20777), .B1(n15161), .B2(n13828), .C1(
        n15150), .C2(n20823), .ZN(P1_U2903) );
  INV_X1 U17265 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20827) );
  OAI222_X1 U17266 ( .A1(n15163), .A2(n15041), .B1(n15150), .B2(n20827), .C1(
        n15143), .C2(n15161), .ZN(P1_U2904) );
  NOR2_X1 U17267 ( .A1(n20651), .A2(n20660), .ZN(n20406) );
  NAND2_X1 U17268 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20406), .ZN(
        n16868) );
  OAI21_X1 U17269 ( .B1(n20313), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n16868), .ZN(n16885) );
  NAND2_X1 U17270 ( .A1(n13865), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13764) );
  OAI21_X1 U17271 ( .B1(n20628), .B2(n16885), .A(n13764), .ZN(n13765) );
  NAND2_X1 U17272 ( .A1(n14625), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13768) );
  OAI22_X1 U17273 ( .A1(n13771), .A2(n13770), .B1(n13769), .B2(n16826), .ZN(
        n13772) );
  INV_X1 U17274 ( .A(n13772), .ZN(n13863) );
  INV_X1 U17275 ( .A(n20647), .ZN(n16848) );
  MUX2_X1 U17276 ( .A(n10868), .B(n13773), .S(n16157), .Z(n13774) );
  OAI21_X1 U17277 ( .B1(n16848), .B2(n9716), .A(n13774), .ZN(P2_U2885) );
  INV_X1 U17278 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13779) );
  NAND2_X1 U17279 ( .A1(n20801), .A2(n9581), .ZN(n14003) );
  NOR2_X1 U17280 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17218), .ZN(n13997) );
  NOR2_X4 U17281 ( .A1(n20801), .A2(n20824), .ZN(n20814) );
  AOI22_X1 U17282 ( .A1(n20824), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13778) );
  OAI21_X1 U17283 ( .B1(n13779), .B2(n14003), .A(n13778), .ZN(P1_U2909) );
  AOI22_X1 U17284 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20824), .B1(n20814), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13780) );
  OAI21_X1 U17285 ( .B1(n15073), .B2(n14003), .A(n13780), .ZN(P1_U2906) );
  INV_X1 U17286 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n20830) );
  AOI22_X1 U17287 ( .A1(n13997), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13781) );
  OAI21_X1 U17288 ( .B1(n20830), .B2(n14003), .A(n13781), .ZN(P1_U2911) );
  INV_X1 U17289 ( .A(n13879), .ZN(n13782) );
  AOI21_X1 U17290 ( .B1(n13783), .B2(n13754), .A(n13782), .ZN(n16730) );
  INV_X1 U17291 ( .A(n16730), .ZN(n19823) );
  AOI22_X1 U17292 ( .A1(n16279), .A2(n16181), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n19887), .ZN(n13784) );
  OAI21_X1 U17293 ( .B1(n19823), .B2(n16275), .A(n13784), .ZN(P2_U2909) );
  XOR2_X1 U17294 ( .A(n13785), .B(n13738), .Z(n20877) );
  INV_X1 U17295 ( .A(n20877), .ZN(n13789) );
  AOI21_X1 U17296 ( .B1(n13787), .B2(n13786), .A(n10427), .ZN(n20917) );
  AOI22_X1 U17297 ( .A1(n20795), .A2(n20917), .B1(n15065), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13788) );
  OAI21_X1 U17298 ( .B1(n13789), .B2(n15070), .A(n13788), .ZN(P1_U2870) );
  INV_X1 U17299 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20821) );
  OAI222_X1 U17300 ( .A1(n15163), .A2(n13789), .B1(n15131), .B2(n15161), .C1(
        n15150), .C2(n20821), .ZN(P1_U2902) );
  NAND2_X1 U17301 ( .A1(n20891), .A2(n13790), .ZN(n20939) );
  AOI21_X1 U17302 ( .B1(n15583), .B2(n20939), .A(n20913), .ZN(n13796) );
  OAI21_X1 U17303 ( .B1(n13792), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n13791), .ZN(n20883) );
  AOI22_X1 U17304 ( .A1(n17191), .A2(n20778), .B1(n20916), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n13794) );
  OAI211_X1 U17305 ( .C1(n20936), .C2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n15521), .B(n20913), .ZN(n13793) );
  OAI211_X1 U17306 ( .C1(n20883), .C2(n20933), .A(n13794), .B(n13793), .ZN(
        n13795) );
  OR2_X1 U17307 ( .A1(n13796), .A2(n13795), .ZN(P1_U3030) );
  NAND2_X1 U17308 ( .A1(n14190), .A2(n21136), .ZN(n13805) );
  INV_X1 U17309 ( .A(n13805), .ZN(n13801) );
  NOR2_X1 U17310 ( .A1(n13618), .A2(n13883), .ZN(n15728) );
  INV_X1 U17311 ( .A(n13797), .ZN(n14085) );
  NOR2_X1 U17312 ( .A1(n14084), .A2(n13805), .ZN(n13847) );
  AOI21_X1 U17313 ( .B1(n15728), .B2(n14085), .A(n13847), .ZN(n13806) );
  OAI21_X1 U17314 ( .B1(n15659), .B2(n20709), .A(n13806), .ZN(n13800) );
  OAI221_X1 U17315 ( .B1(n21149), .B2(n13801), .C1(n21141), .C2(n13800), .A(
        n21147), .ZN(n13802) );
  INV_X1 U17316 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13812) );
  NOR2_X2 U17317 ( .A1(n15382), .A2(n13803), .ZN(n13844) );
  AOI22_X1 U17318 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n13844), .B1(DATAI_21_), 
        .B2(n13804), .ZN(n21121) );
  INV_X1 U17319 ( .A(n21121), .ZN(n21180) );
  AOI22_X1 U17320 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n13844), .B1(DATAI_29_), 
        .B2(n13804), .ZN(n21183) );
  INV_X1 U17321 ( .A(n14013), .ZN(n15640) );
  OAI22_X1 U17322 ( .A1(n13806), .A2(n21141), .B1(n13805), .B2(n11830), .ZN(
        n13848) );
  NOR2_X1 U17323 ( .A1(n13846), .A2(n13808), .ZN(n21178) );
  AOI22_X1 U17324 ( .A1(n21179), .A2(n13848), .B1(n21178), .B2(n13847), .ZN(
        n13809) );
  OAI21_X1 U17325 ( .B1(n21183), .B2(n14193), .A(n13809), .ZN(n13810) );
  AOI21_X1 U17326 ( .B1(n15770), .B2(n21180), .A(n13810), .ZN(n13811) );
  OAI21_X1 U17327 ( .B1(n13853), .B2(n13812), .A(n13811), .ZN(P1_U3078) );
  INV_X1 U17328 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13817) );
  INV_X1 U17329 ( .A(n21191), .ZN(n21081) );
  AOI22_X1 U17330 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n13844), .B1(DATAI_30_), 
        .B2(n13804), .ZN(n21084) );
  AOI22_X1 U17331 ( .A1(n21185), .A2(n13848), .B1(n21184), .B2(n13847), .ZN(
        n13814) );
  OAI21_X1 U17332 ( .B1(n21084), .B2(n14193), .A(n13814), .ZN(n13815) );
  AOI21_X1 U17333 ( .B1(n15770), .B2(n21081), .A(n13815), .ZN(n13816) );
  OAI21_X1 U17334 ( .B1(n13853), .B2(n13817), .A(n13816), .ZN(P1_U3079) );
  INV_X1 U17335 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13822) );
  AOI22_X1 U17336 ( .A1(DATAI_16_), .A2(n13804), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n13844), .ZN(n21153) );
  INV_X1 U17337 ( .A(n21153), .ZN(n21055) );
  AOI22_X1 U17338 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n13844), .B1(DATAI_24_), 
        .B2(n13804), .ZN(n21070) );
  AOI22_X1 U17339 ( .A1(n21139), .A2(n13848), .B1(n21138), .B2(n13847), .ZN(
        n13819) );
  OAI21_X1 U17340 ( .B1(n21070), .B2(n14193), .A(n13819), .ZN(n13820) );
  AOI21_X1 U17341 ( .B1(n15770), .B2(n21055), .A(n13820), .ZN(n13821) );
  OAI21_X1 U17342 ( .B1(n13853), .B2(n13822), .A(n13821), .ZN(P1_U3073) );
  INV_X1 U17343 ( .A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13827) );
  AOI22_X1 U17344 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n13844), .B1(DATAI_19_), 
        .B2(n13804), .ZN(n21113) );
  INV_X1 U17345 ( .A(n21113), .ZN(n21168) );
  AOI22_X1 U17346 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n13844), .B1(DATAI_27_), 
        .B2(n13804), .ZN(n21171) );
  AOI22_X1 U17347 ( .A1(n21167), .A2(n13848), .B1(n21166), .B2(n13847), .ZN(
        n13824) );
  OAI21_X1 U17348 ( .B1(n21171), .B2(n14193), .A(n13824), .ZN(n13825) );
  AOI21_X1 U17349 ( .B1(n15770), .B2(n21168), .A(n13825), .ZN(n13826) );
  OAI21_X1 U17350 ( .B1(n13853), .B2(n13827), .A(n13826), .ZN(P1_U3076) );
  INV_X1 U17351 ( .A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13833) );
  AOI22_X1 U17352 ( .A1(DATAI_17_), .A2(n13804), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n13844), .ZN(n21105) );
  INV_X1 U17353 ( .A(n21105), .ZN(n21156) );
  AOI22_X1 U17354 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n13844), .B1(DATAI_25_), 
        .B2(n13804), .ZN(n21159) );
  AOI22_X1 U17355 ( .A1(n21155), .A2(n13848), .B1(n21154), .B2(n13847), .ZN(
        n13830) );
  OAI21_X1 U17356 ( .B1(n21159), .B2(n14193), .A(n13830), .ZN(n13831) );
  AOI21_X1 U17357 ( .B1(n15770), .B2(n21156), .A(n13831), .ZN(n13832) );
  OAI21_X1 U17358 ( .B1(n13853), .B2(n13833), .A(n13832), .ZN(P1_U3074) );
  AOI22_X1 U17359 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n13844), .B1(DATAI_23_), 
        .B2(n13804), .ZN(n21131) );
  INV_X1 U17360 ( .A(n21131), .ZN(n21196) );
  AOI22_X1 U17361 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n13844), .B1(DATAI_31_), 
        .B2(n13804), .ZN(n21202) );
  AOI22_X1 U17362 ( .A1(n21195), .A2(n13848), .B1(n21193), .B2(n13847), .ZN(
        n13835) );
  OAI21_X1 U17363 ( .B1(n21202), .B2(n14193), .A(n13835), .ZN(n13836) );
  AOI21_X1 U17364 ( .B1(n15770), .B2(n21196), .A(n13836), .ZN(n13837) );
  OAI21_X1 U17365 ( .B1(n13853), .B2(n13838), .A(n13837), .ZN(P1_U3080) );
  AOI22_X1 U17366 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n13844), .B1(DATAI_18_), 
        .B2(n13804), .ZN(n21109) );
  INV_X1 U17367 ( .A(n21109), .ZN(n21162) );
  AOI22_X1 U17368 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n13844), .B1(DATAI_26_), 
        .B2(n13804), .ZN(n21165) );
  NOR2_X1 U17369 ( .A1(n13846), .A2(n13839), .ZN(n21160) );
  AOI22_X1 U17370 ( .A1(n21161), .A2(n13848), .B1(n21160), .B2(n13847), .ZN(
        n13840) );
  OAI21_X1 U17371 ( .B1(n21165), .B2(n14193), .A(n13840), .ZN(n13841) );
  AOI21_X1 U17372 ( .B1(n15770), .B2(n21162), .A(n13841), .ZN(n13842) );
  OAI21_X1 U17373 ( .B1(n13853), .B2(n13843), .A(n13842), .ZN(P1_U3075) );
  AOI22_X1 U17374 ( .A1(DATAI_20_), .A2(n13804), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n13844), .ZN(n21117) );
  INV_X1 U17375 ( .A(n21117), .ZN(n21174) );
  AOI22_X1 U17376 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n13844), .B1(DATAI_28_), 
        .B2(n13804), .ZN(n21177) );
  NOR2_X1 U17377 ( .A1(n13846), .A2(n13845), .ZN(n21172) );
  AOI22_X1 U17378 ( .A1(n21173), .A2(n13848), .B1(n21172), .B2(n13847), .ZN(
        n13849) );
  OAI21_X1 U17379 ( .B1(n21177), .B2(n14193), .A(n13849), .ZN(n13850) );
  AOI21_X1 U17380 ( .B1(n15770), .B2(n21174), .A(n13850), .ZN(n13851) );
  OAI21_X1 U17381 ( .B1(n13853), .B2(n13852), .A(n13851), .ZN(P1_U3077) );
  OAI21_X1 U17382 ( .B1(n13854), .B2(n13857), .A(n13856), .ZN(n16705) );
  AOI22_X1 U17383 ( .A1(n16279), .A2(n16167), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n19887), .ZN(n13858) );
  OAI21_X1 U17384 ( .B1(n16705), .B2(n16275), .A(n13858), .ZN(P2_U2907) );
  NAND2_X1 U17385 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20643), .ZN(
        n20113) );
  INV_X1 U17386 ( .A(n20113), .ZN(n20148) );
  NAND2_X1 U17387 ( .A1(n16868), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13864) );
  AOI21_X1 U17388 ( .B1(n20216), .B2(n13864), .A(n20628), .ZN(n20345) );
  AOI21_X1 U17389 ( .B1(n13865), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n20345), .ZN(n13866) );
  INV_X1 U17390 ( .A(n14054), .ZN(n13868) );
  NAND2_X1 U17391 ( .A1(n14625), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13869) );
  INV_X1 U17392 ( .A(n13869), .ZN(n13870) );
  NAND2_X1 U17393 ( .A1(n14054), .A2(n13870), .ZN(n13925) );
  INV_X1 U17394 ( .A(n13872), .ZN(n13873) );
  NAND2_X1 U17395 ( .A1(n13873), .A2(n14056), .ZN(n13874) );
  INV_X1 U17396 ( .A(n20637), .ZN(n16864) );
  NOR2_X1 U17397 ( .A1(n13875), .A2(n16157), .ZN(n13876) );
  AOI21_X1 U17398 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n16157), .A(n13876), .ZN(
        n13877) );
  OAI21_X1 U17399 ( .B1(n16864), .B2(n9716), .A(n13877), .ZN(P2_U2884) );
  AND2_X1 U17400 ( .A1(n13879), .A2(n13878), .ZN(n13880) );
  NOR2_X1 U17401 ( .A1(n13854), .A2(n13880), .ZN(n19804) );
  INV_X1 U17402 ( .A(n19804), .ZN(n13882) );
  INV_X1 U17403 ( .A(n16175), .ZN(n13881) );
  INV_X1 U17404 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19911) );
  OAI222_X1 U17405 ( .A1(n13882), .A2(n16275), .B1(n13881), .B2(n19896), .C1(
        n19911), .C2(n16287), .ZN(P2_U2908) );
  NAND2_X1 U17406 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21135) );
  NOR2_X1 U17407 ( .A1(n21135), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13886) );
  INV_X1 U17408 ( .A(n13883), .ZN(n15633) );
  NOR2_X1 U17409 ( .A1(n13618), .A2(n15633), .ZN(n21134) );
  NOR3_X2 U17410 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n14084), .A3(
        n21135), .ZN(n13917) );
  AOI21_X1 U17411 ( .B1(n21134), .B2(n14085), .A(n13917), .ZN(n13888) );
  OAI211_X1 U17412 ( .C1(n21140), .C2(n20709), .A(n21149), .B(n13888), .ZN(
        n13884) );
  OAI211_X1 U17413 ( .C1(n21149), .C2(n13886), .A(n21147), .B(n13884), .ZN(
        n13885) );
  INV_X1 U17414 ( .A(n13886), .ZN(n13887) );
  OAI22_X1 U17415 ( .A1(n13888), .A2(n21141), .B1(n13887), .B2(n11830), .ZN(
        n13918) );
  AOI22_X1 U17416 ( .A1(n21173), .A2(n13918), .B1(n21172), .B2(n13917), .ZN(
        n13889) );
  OAI21_X1 U17417 ( .B1(n21177), .B2(n21054), .A(n13889), .ZN(n13890) );
  AOI21_X1 U17418 ( .B1(n21127), .B2(n21174), .A(n13890), .ZN(n13891) );
  OAI21_X1 U17419 ( .B1(n13923), .B2(n13892), .A(n13891), .ZN(P1_U3141) );
  INV_X1 U17420 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13896) );
  AOI22_X1 U17421 ( .A1(n21139), .A2(n13918), .B1(n21138), .B2(n13917), .ZN(
        n13893) );
  OAI21_X1 U17422 ( .B1(n21070), .B2(n21054), .A(n13893), .ZN(n13894) );
  AOI21_X1 U17423 ( .B1(n21127), .B2(n21055), .A(n13894), .ZN(n13895) );
  OAI21_X1 U17424 ( .B1(n13923), .B2(n13896), .A(n13895), .ZN(P1_U3137) );
  INV_X1 U17425 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13900) );
  AOI22_X1 U17426 ( .A1(n21179), .A2(n13918), .B1(n21178), .B2(n13917), .ZN(
        n13897) );
  OAI21_X1 U17427 ( .B1(n21183), .B2(n21054), .A(n13897), .ZN(n13898) );
  AOI21_X1 U17428 ( .B1(n21127), .B2(n21180), .A(n13898), .ZN(n13899) );
  OAI21_X1 U17429 ( .B1(n13923), .B2(n13900), .A(n13899), .ZN(P1_U3142) );
  INV_X1 U17430 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13904) );
  AOI22_X1 U17431 ( .A1(n21155), .A2(n13918), .B1(n21154), .B2(n13917), .ZN(
        n13901) );
  OAI21_X1 U17432 ( .B1(n21159), .B2(n21054), .A(n13901), .ZN(n13902) );
  AOI21_X1 U17433 ( .B1(n21127), .B2(n21156), .A(n13902), .ZN(n13903) );
  OAI21_X1 U17434 ( .B1(n13923), .B2(n13904), .A(n13903), .ZN(P1_U3138) );
  AOI22_X1 U17435 ( .A1(n21195), .A2(n13918), .B1(n21193), .B2(n13917), .ZN(
        n13905) );
  OAI21_X1 U17436 ( .B1(n21202), .B2(n21054), .A(n13905), .ZN(n13906) );
  AOI21_X1 U17437 ( .B1(n21127), .B2(n21196), .A(n13906), .ZN(n13907) );
  OAI21_X1 U17438 ( .B1(n13923), .B2(n13908), .A(n13907), .ZN(P1_U3144) );
  INV_X1 U17439 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13912) );
  AOI22_X1 U17440 ( .A1(n21161), .A2(n13918), .B1(n21160), .B2(n13917), .ZN(
        n13909) );
  OAI21_X1 U17441 ( .B1(n21165), .B2(n21054), .A(n13909), .ZN(n13910) );
  AOI21_X1 U17442 ( .B1(n21127), .B2(n21162), .A(n13910), .ZN(n13911) );
  OAI21_X1 U17443 ( .B1(n13923), .B2(n13912), .A(n13911), .ZN(P1_U3139) );
  INV_X1 U17444 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13916) );
  AOI22_X1 U17445 ( .A1(n21185), .A2(n13918), .B1(n21184), .B2(n13917), .ZN(
        n13913) );
  OAI21_X1 U17446 ( .B1(n21084), .B2(n21054), .A(n13913), .ZN(n13914) );
  AOI21_X1 U17447 ( .B1(n21127), .B2(n21081), .A(n13914), .ZN(n13915) );
  OAI21_X1 U17448 ( .B1(n13923), .B2(n13916), .A(n13915), .ZN(P1_U3143) );
  INV_X1 U17449 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13922) );
  AOI22_X1 U17450 ( .A1(n21167), .A2(n13918), .B1(n21166), .B2(n13917), .ZN(
        n13919) );
  OAI21_X1 U17451 ( .B1(n21171), .B2(n21054), .A(n13919), .ZN(n13920) );
  AOI21_X1 U17452 ( .B1(n21127), .B2(n21168), .A(n13920), .ZN(n13921) );
  OAI21_X1 U17453 ( .B1(n13923), .B2(n13922), .A(n13921), .ZN(P1_U3140) );
  NAND2_X1 U17454 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n10794), .ZN(
        n13924) );
  AND2_X1 U17455 ( .A1(n13925), .A2(n13924), .ZN(n13926) );
  NAND2_X1 U17456 ( .A1(n14625), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14103) );
  XNOR2_X1 U17457 ( .A(n14102), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13933) );
  NAND2_X1 U17458 ( .A1(n13928), .A2(n13929), .ZN(n13978) );
  OR2_X1 U17459 ( .A1(n13928), .A2(n13929), .ZN(n13930) );
  AND2_X1 U17460 ( .A1(n13978), .A2(n13930), .ZN(n16787) );
  INV_X1 U17461 ( .A(n16787), .ZN(n15980) );
  MUX2_X1 U17462 ( .A(n15980), .B(n13931), .S(n16157), .Z(n13932) );
  OAI21_X1 U17463 ( .B1(n13933), .B2(n9716), .A(n13932), .ZN(P2_U2882) );
  NAND2_X1 U17464 ( .A1(n13856), .A2(n13935), .ZN(n13936) );
  NAND2_X1 U17465 ( .A1(n13934), .A2(n13936), .ZN(n16699) );
  INV_X1 U17466 ( .A(n16159), .ZN(n13937) );
  INV_X1 U17467 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19907) );
  OAI222_X1 U17468 ( .A1(n16699), .A2(n16275), .B1(n13937), .B2(n19896), .C1(
        n19907), .C2(n16287), .ZN(P2_U2906) );
  INV_X1 U17469 ( .A(n21171), .ZN(n21110) );
  INV_X1 U17470 ( .A(n21167), .ZN(n15752) );
  INV_X1 U17471 ( .A(n13618), .ZN(n15030) );
  OR2_X1 U17472 ( .A1(n15657), .A2(n15030), .ZN(n15681) );
  INV_X1 U17473 ( .A(n15681), .ZN(n13939) );
  NOR2_X1 U17474 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n15686) );
  NAND2_X1 U17475 ( .A1(n15686), .A2(n21136), .ZN(n13943) );
  NOR2_X1 U17476 ( .A1(n14084), .A2(n13943), .ZN(n13941) );
  AOI21_X1 U17477 ( .B1(n13939), .B2(n14085), .A(n13941), .ZN(n13944) );
  OAI22_X1 U17478 ( .A1(n13944), .A2(n21141), .B1(n13943), .B2(n11830), .ZN(
        n13940) );
  INV_X1 U17479 ( .A(n21166), .ZN(n15703) );
  INV_X1 U17480 ( .A(n13941), .ZN(n13967) );
  OAI22_X1 U17481 ( .A1(n15752), .A2(n13968), .B1(n15703), .B2(n13967), .ZN(
        n13942) );
  AOI21_X1 U17482 ( .B1(n15723), .B2(n21110), .A(n13942), .ZN(n13948) );
  INV_X1 U17483 ( .A(n13943), .ZN(n13946) );
  OAI211_X1 U17484 ( .C1(n14066), .C2(n20709), .A(n21149), .B(n13944), .ZN(
        n13945) );
  NAND2_X1 U17485 ( .A1(n13970), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n13947) );
  OAI211_X1 U17486 ( .C1(n21113), .C2(n13973), .A(n13948), .B(n13947), .ZN(
        P1_U3044) );
  INV_X1 U17487 ( .A(n21084), .ZN(n21186) );
  INV_X1 U17488 ( .A(n21185), .ZN(n15764) );
  INV_X1 U17489 ( .A(n21184), .ZN(n15715) );
  OAI22_X1 U17490 ( .A1(n15764), .A2(n13968), .B1(n15715), .B2(n13967), .ZN(
        n13949) );
  AOI21_X1 U17491 ( .B1(n15723), .B2(n21186), .A(n13949), .ZN(n13951) );
  NAND2_X1 U17492 ( .A1(n13970), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n13950) );
  OAI211_X1 U17493 ( .C1(n21191), .C2(n13973), .A(n13951), .B(n13950), .ZN(
        P1_U3047) );
  INV_X1 U17494 ( .A(n21159), .ZN(n21102) );
  INV_X1 U17495 ( .A(n21155), .ZN(n15744) );
  INV_X1 U17496 ( .A(n21154), .ZN(n15695) );
  OAI22_X1 U17497 ( .A1(n15744), .A2(n13968), .B1(n15695), .B2(n13967), .ZN(
        n13952) );
  AOI21_X1 U17498 ( .B1(n15723), .B2(n21102), .A(n13952), .ZN(n13954) );
  NAND2_X1 U17499 ( .A1(n13970), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13953) );
  OAI211_X1 U17500 ( .C1(n21105), .C2(n13973), .A(n13954), .B(n13953), .ZN(
        P1_U3042) );
  INV_X1 U17501 ( .A(n21177), .ZN(n21114) );
  INV_X1 U17502 ( .A(n21172), .ZN(n15707) );
  OAI22_X1 U17503 ( .A1(n15756), .A2(n13968), .B1(n15707), .B2(n13967), .ZN(
        n13955) );
  AOI21_X1 U17504 ( .B1(n15723), .B2(n21114), .A(n13955), .ZN(n13957) );
  NAND2_X1 U17505 ( .A1(n13970), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n13956) );
  OAI211_X1 U17506 ( .C1(n21117), .C2(n13973), .A(n13957), .B(n13956), .ZN(
        P1_U3045) );
  INV_X1 U17507 ( .A(n21183), .ZN(n21118) );
  INV_X1 U17508 ( .A(n21179), .ZN(n15760) );
  INV_X1 U17509 ( .A(n21178), .ZN(n15711) );
  OAI22_X1 U17510 ( .A1(n15760), .A2(n13968), .B1(n15711), .B2(n13967), .ZN(
        n13958) );
  AOI21_X1 U17511 ( .B1(n15723), .B2(n21118), .A(n13958), .ZN(n13960) );
  NAND2_X1 U17512 ( .A1(n13970), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n13959) );
  OAI211_X1 U17513 ( .C1(n21121), .C2(n13973), .A(n13960), .B(n13959), .ZN(
        P1_U3046) );
  INV_X1 U17514 ( .A(n21070), .ZN(n21150) );
  INV_X1 U17515 ( .A(n21139), .ZN(n15740) );
  INV_X1 U17516 ( .A(n21138), .ZN(n15691) );
  OAI22_X1 U17517 ( .A1(n15740), .A2(n13968), .B1(n15691), .B2(n13967), .ZN(
        n13961) );
  AOI21_X1 U17518 ( .B1(n15723), .B2(n21150), .A(n13961), .ZN(n13963) );
  NAND2_X1 U17519 ( .A1(n13970), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13962) );
  OAI211_X1 U17520 ( .C1(n21153), .C2(n13973), .A(n13963), .B(n13962), .ZN(
        P1_U3041) );
  INV_X1 U17521 ( .A(n21165), .ZN(n21106) );
  INV_X1 U17522 ( .A(n21161), .ZN(n15748) );
  INV_X1 U17523 ( .A(n21160), .ZN(n15699) );
  OAI22_X1 U17524 ( .A1(n15748), .A2(n13968), .B1(n15699), .B2(n13967), .ZN(
        n13964) );
  AOI21_X1 U17525 ( .B1(n15723), .B2(n21106), .A(n13964), .ZN(n13966) );
  NAND2_X1 U17526 ( .A1(n13970), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n13965) );
  OAI211_X1 U17527 ( .C1(n21109), .C2(n13973), .A(n13966), .B(n13965), .ZN(
        P1_U3043) );
  INV_X1 U17528 ( .A(n21202), .ZN(n21126) );
  INV_X1 U17529 ( .A(n21195), .ZN(n15772) );
  INV_X1 U17530 ( .A(n21193), .ZN(n15721) );
  OAI22_X1 U17531 ( .A1(n15772), .A2(n13968), .B1(n15721), .B2(n13967), .ZN(
        n13969) );
  AOI21_X1 U17532 ( .B1(n15723), .B2(n21126), .A(n13969), .ZN(n13972) );
  NAND2_X1 U17533 ( .A1(n13970), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n13971) );
  OAI211_X1 U17534 ( .C1(n21131), .C2(n13973), .A(n13972), .B(n13971), .ZN(
        P1_U3048) );
  XOR2_X1 U17535 ( .A(n13974), .B(n13975), .Z(n20869) );
  INV_X1 U17536 ( .A(n20869), .ZN(n14048) );
  INV_X1 U17537 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20819) );
  OAI222_X1 U17538 ( .A1(n15163), .A2(n14048), .B1(n15161), .B2(n15126), .C1(
        n15150), .C2(n20819), .ZN(P1_U2901) );
  AND2_X1 U17539 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14057) );
  NAND2_X1 U17540 ( .A1(n14102), .A2(n14057), .ZN(n14211) );
  NAND2_X1 U17541 ( .A1(n14211), .A2(n16150), .ZN(n13983) );
  AOI21_X1 U17542 ( .B1(n14102), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13982) );
  NAND2_X1 U17543 ( .A1(n13978), .A2(n13977), .ZN(n13979) );
  NAND2_X1 U17544 ( .A1(n13976), .A2(n13979), .ZN(n19872) );
  MUX2_X1 U17545 ( .A(n19872), .B(n13980), .S(n16157), .Z(n13981) );
  OAI21_X1 U17546 ( .B1(n13983), .B2(n13982), .A(n13981), .ZN(P2_U2881) );
  INV_X1 U17547 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13985) );
  AOI22_X1 U17548 ( .A1(n13997), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13984) );
  OAI21_X1 U17549 ( .B1(n13985), .B2(n14003), .A(n13984), .ZN(P1_U2919) );
  AOI22_X1 U17550 ( .A1(n13997), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13986) );
  OAI21_X1 U17551 ( .B1(n15102), .B2(n14003), .A(n13986), .ZN(P1_U2912) );
  INV_X1 U17552 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13988) );
  AOI22_X1 U17553 ( .A1(n13997), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13987) );
  OAI21_X1 U17554 ( .B1(n13988), .B2(n14003), .A(n13987), .ZN(P1_U2913) );
  INV_X1 U17555 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13990) );
  AOI22_X1 U17556 ( .A1(n13997), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13989) );
  OAI21_X1 U17557 ( .B1(n13990), .B2(n14003), .A(n13989), .ZN(P1_U2917) );
  AOI22_X1 U17558 ( .A1(n13997), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13991) );
  OAI21_X1 U17559 ( .B1(n15116), .B2(n14003), .A(n13991), .ZN(P1_U2915) );
  INV_X1 U17560 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13993) );
  AOI22_X1 U17561 ( .A1(n13997), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13992) );
  OAI21_X1 U17562 ( .B1(n13993), .B2(n14003), .A(n13992), .ZN(P1_U2914) );
  AOI22_X1 U17563 ( .A1(n13997), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13994) );
  OAI21_X1 U17564 ( .B1(n12386), .B2(n14003), .A(n13994), .ZN(P1_U2910) );
  INV_X1 U17565 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13996) );
  AOI22_X1 U17566 ( .A1(n13997), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13995) );
  OAI21_X1 U17567 ( .B1(n13996), .B2(n14003), .A(n13995), .ZN(P1_U2916) );
  INV_X1 U17568 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13999) );
  AOI22_X1 U17569 ( .A1(n13997), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13998) );
  OAI21_X1 U17570 ( .B1(n13999), .B2(n14003), .A(n13998), .ZN(P1_U2918) );
  INV_X1 U17571 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n20840) );
  AOI22_X1 U17572 ( .A1(n20824), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n14000) );
  OAI21_X1 U17573 ( .B1(n20840), .B2(n14003), .A(n14000), .ZN(P1_U2907) );
  AOI22_X1 U17574 ( .A1(n20824), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n14001) );
  OAI21_X1 U17575 ( .B1(n15142), .B2(n14003), .A(n14001), .ZN(P1_U2920) );
  INV_X1 U17576 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n20836) );
  AOI22_X1 U17577 ( .A1(n20824), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14002) );
  OAI21_X1 U17578 ( .B1(n20836), .B2(n14003), .A(n14002), .ZN(P1_U2908) );
  INV_X1 U17579 ( .A(n15659), .ZN(n14004) );
  NAND2_X1 U17580 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n14190), .ZN(
        n15731) );
  NOR2_X1 U17581 ( .A1(n14005), .A2(n21141), .ZN(n14009) );
  INV_X1 U17582 ( .A(n14006), .ZN(n15653) );
  NAND2_X1 U17583 ( .A1(n21029), .A2(n20709), .ZN(n21057) );
  INV_X1 U17584 ( .A(n21145), .ZN(n14008) );
  OAI21_X1 U17585 ( .B1(n15653), .B2(n21141), .A(n14008), .ZN(n15652) );
  AOI211_X1 U17586 ( .C1(n15731), .C2(n21141), .A(n14009), .B(n15652), .ZN(
        n14012) );
  AND2_X1 U17587 ( .A1(n14010), .A2(n15641), .ZN(n21133) );
  NAND2_X1 U17588 ( .A1(n15728), .A2(n21133), .ZN(n14011) );
  AOI21_X1 U17589 ( .B1(n14011), .B2(n14039), .A(n21141), .ZN(n14015) );
  NAND2_X1 U17590 ( .A1(n14038), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14019) );
  INV_X1 U17591 ( .A(n15731), .ZN(n14016) );
  AOI21_X1 U17592 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14016), .A(n14015), 
        .ZN(n14040) );
  OAI22_X1 U17593 ( .A1(n15760), .A2(n14040), .B1(n15711), .B2(n14039), .ZN(
        n14017) );
  AOI21_X1 U17594 ( .B1(n14042), .B2(n21118), .A(n14017), .ZN(n14018) );
  OAI211_X1 U17595 ( .C1(n21121), .C2(n14112), .A(n14019), .B(n14018), .ZN(
        P1_U3094) );
  NAND2_X1 U17596 ( .A1(n14038), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n14022) );
  OAI22_X1 U17597 ( .A1(n15744), .A2(n14040), .B1(n15695), .B2(n14039), .ZN(
        n14020) );
  AOI21_X1 U17598 ( .B1(n14042), .B2(n21102), .A(n14020), .ZN(n14021) );
  OAI211_X1 U17599 ( .C1(n21105), .C2(n14112), .A(n14022), .B(n14021), .ZN(
        P1_U3090) );
  NAND2_X1 U17600 ( .A1(n14038), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14025) );
  OAI22_X1 U17601 ( .A1(n15772), .A2(n14040), .B1(n15721), .B2(n14039), .ZN(
        n14023) );
  AOI21_X1 U17602 ( .B1(n14042), .B2(n21126), .A(n14023), .ZN(n14024) );
  OAI211_X1 U17603 ( .C1(n21131), .C2(n14112), .A(n14025), .B(n14024), .ZN(
        P1_U3096) );
  NAND2_X1 U17604 ( .A1(n14038), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14028) );
  OAI22_X1 U17605 ( .A1(n15748), .A2(n14040), .B1(n15699), .B2(n14039), .ZN(
        n14026) );
  AOI21_X1 U17606 ( .B1(n14042), .B2(n21106), .A(n14026), .ZN(n14027) );
  OAI211_X1 U17607 ( .C1(n21109), .C2(n14112), .A(n14028), .B(n14027), .ZN(
        P1_U3091) );
  NAND2_X1 U17608 ( .A1(n14038), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n14031) );
  OAI22_X1 U17609 ( .A1(n15764), .A2(n14040), .B1(n15715), .B2(n14039), .ZN(
        n14029) );
  AOI21_X1 U17610 ( .B1(n14042), .B2(n21186), .A(n14029), .ZN(n14030) );
  OAI211_X1 U17611 ( .C1(n21191), .C2(n14112), .A(n14031), .B(n14030), .ZN(
        P1_U3095) );
  NAND2_X1 U17612 ( .A1(n14038), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n14034) );
  OAI22_X1 U17613 ( .A1(n15752), .A2(n14040), .B1(n15703), .B2(n14039), .ZN(
        n14032) );
  AOI21_X1 U17614 ( .B1(n14042), .B2(n21110), .A(n14032), .ZN(n14033) );
  OAI211_X1 U17615 ( .C1(n21113), .C2(n14112), .A(n14034), .B(n14033), .ZN(
        P1_U3092) );
  NAND2_X1 U17616 ( .A1(n14038), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14037) );
  OAI22_X1 U17617 ( .A1(n15756), .A2(n14040), .B1(n15707), .B2(n14039), .ZN(
        n14035) );
  AOI21_X1 U17618 ( .B1(n14042), .B2(n21114), .A(n14035), .ZN(n14036) );
  OAI211_X1 U17619 ( .C1(n21117), .C2(n14112), .A(n14037), .B(n14036), .ZN(
        P1_U3093) );
  NAND2_X1 U17620 ( .A1(n14038), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n14044) );
  OAI22_X1 U17621 ( .A1(n15740), .A2(n14040), .B1(n15691), .B2(n14039), .ZN(
        n14041) );
  AOI21_X1 U17622 ( .B1(n14042), .B2(n21150), .A(n14041), .ZN(n14043) );
  OAI211_X1 U17623 ( .C1(n21153), .C2(n14112), .A(n14044), .B(n14043), .ZN(
        P1_U3089) );
  AND2_X1 U17624 ( .A1(n14046), .A2(n14045), .ZN(n14047) );
  OR2_X1 U17625 ( .A1(n14047), .A2(n14169), .ZN(n20901) );
  INV_X1 U17626 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n14049) );
  OAI222_X1 U17627 ( .A1(n20901), .A2(n15068), .B1(n14049), .B2(n20800), .C1(
        n14048), .C2(n15070), .ZN(P1_U2869) );
  NOR2_X1 U17628 ( .A1(n14051), .A2(n14052), .ZN(n14053) );
  OR2_X1 U17629 ( .A1(n14050), .A2(n14053), .ZN(n16710) );
  NAND2_X1 U17630 ( .A1(n14054), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14055) );
  NAND4_X1 U17631 ( .A1(n14057), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A3(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .A4(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n14058) );
  NOR2_X1 U17632 ( .A1(n16134), .A2(n14058), .ZN(n14060) );
  AND2_X1 U17633 ( .A1(n16140), .A2(n16152), .ZN(n14059) );
  AND4_X1 U17634 ( .A1(n14060), .A2(n14059), .A3(n19972), .A4(n14212), .ZN(
        n14061) );
  AOI211_X1 U17635 ( .C1(n14063), .C2(n16136), .A(n9716), .B(n14156), .ZN(
        n14064) );
  AOI21_X1 U17636 ( .B1(P2_EBX_REG_12__SCAN_IN), .B2(n16157), .A(n14064), .ZN(
        n14065) );
  OAI21_X1 U17637 ( .B1(n16157), .B2(n16710), .A(n14065), .ZN(P2_U2875) );
  AOI21_X1 U17638 ( .B1(n14066), .B2(n21149), .A(n21145), .ZN(n14075) );
  INV_X1 U17639 ( .A(n21133), .ZN(n14067) );
  OR2_X1 U17640 ( .A1(n15681), .A2(n14067), .ZN(n14070) );
  INV_X1 U17641 ( .A(n15686), .ZN(n14068) );
  NOR2_X1 U17642 ( .A1(n14068), .A2(n21132), .ZN(n20952) );
  INV_X1 U17643 ( .A(n20952), .ZN(n14069) );
  AND2_X1 U17644 ( .A1(n14070), .A2(n14069), .ZN(n14074) );
  INV_X1 U17645 ( .A(n14074), .ZN(n14073) );
  NAND2_X1 U17646 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n15686), .ZN(
        n14218) );
  AOI21_X1 U17647 ( .B1(n21141), .B2(n14218), .A(n14071), .ZN(n14072) );
  AOI22_X1 U17648 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20954), .B1(
        n21155), .B2(n20953), .ZN(n14079) );
  AOI22_X1 U17649 ( .A1(n21154), .A2(n20952), .B1(n20951), .B2(n21102), .ZN(
        n14078) );
  OAI211_X1 U17650 ( .C1(n21105), .C2(n20972), .A(n14079), .B(n14078), .ZN(
        P1_U3058) );
  AOI22_X1 U17651 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20954), .B1(
        n21185), .B2(n20953), .ZN(n14081) );
  AOI22_X1 U17652 ( .A1(n21184), .A2(n20952), .B1(n20951), .B2(n21186), .ZN(
        n14080) );
  OAI211_X1 U17653 ( .C1(n21191), .C2(n20972), .A(n14081), .B(n14080), .ZN(
        P1_U3063) );
  AOI22_X1 U17654 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20954), .B1(
        n21167), .B2(n20953), .ZN(n14083) );
  AOI22_X1 U17655 ( .A1(n21166), .A2(n20952), .B1(n20951), .B2(n21110), .ZN(
        n14082) );
  OAI211_X1 U17656 ( .C1(n21113), .C2(n20972), .A(n14083), .B(n14082), .ZN(
        P1_U3060) );
  NAND2_X1 U17657 ( .A1(n17091), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21021) );
  NOR2_X1 U17658 ( .A1(n21021), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n14087) );
  AND2_X1 U17659 ( .A1(n13618), .A2(n15657), .ZN(n21022) );
  INV_X1 U17660 ( .A(n14087), .ZN(n14090) );
  NOR2_X1 U17661 ( .A1(n14084), .A2(n14090), .ZN(n20985) );
  AOI21_X1 U17662 ( .B1(n21022), .B2(n14085), .A(n20985), .ZN(n14091) );
  OAI211_X1 U17663 ( .C1(n21031), .C2(n20709), .A(n21149), .B(n14091), .ZN(
        n14086) );
  INV_X1 U17664 ( .A(n20988), .ZN(n14096) );
  INV_X1 U17665 ( .A(n21020), .ZN(n21012) );
  OAI22_X1 U17666 ( .A1(n14091), .A2(n21141), .B1(n14090), .B2(n11830), .ZN(
        n20986) );
  AOI22_X1 U17667 ( .A1(n21179), .A2(n20986), .B1(n21178), .B2(n20985), .ZN(
        n14092) );
  OAI21_X1 U17668 ( .B1(n21183), .B2(n14151), .A(n14092), .ZN(n14093) );
  AOI21_X1 U17669 ( .B1(n21012), .B2(n21180), .A(n14093), .ZN(n14094) );
  OAI21_X1 U17670 ( .B1(n14096), .B2(n14095), .A(n14094), .ZN(P1_U3110) );
  AOI21_X1 U17671 ( .B1(n14098), .B2(n14097), .A(n9717), .ZN(n20861) );
  INV_X1 U17672 ( .A(n20861), .ZN(n14170) );
  INV_X1 U17673 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20817) );
  OAI222_X1 U17674 ( .A1(n15163), .A2(n14170), .B1(n15161), .B2(n15122), .C1(
        n15150), .C2(n20817), .ZN(P1_U2900) );
  NOR2_X1 U17675 ( .A1(n14099), .A2(n14100), .ZN(n14101) );
  OR2_X1 U17676 ( .A1(n13928), .A2(n14101), .ZN(n19949) );
  AOI21_X1 U17677 ( .B1(n14104), .B2(n14103), .A(n14102), .ZN(n16277) );
  NAND2_X1 U17678 ( .A1(n16277), .A2(n16150), .ZN(n14106) );
  NAND2_X1 U17679 ( .A1(n16154), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n14105) );
  OAI211_X1 U17680 ( .C1(n19949), .C2(n16157), .A(n14106), .B(n14105), .ZN(
        P2_U2883) );
  XOR2_X1 U17681 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n14211), .Z(n14111)
         );
  NAND2_X1 U17682 ( .A1(n13976), .A2(n14107), .ZN(n14108) );
  NAND2_X1 U17683 ( .A1(n14208), .A2(n14108), .ZN(n19853) );
  MUX2_X1 U17684 ( .A(n19853), .B(n14109), .S(n16157), .Z(n14110) );
  OAI21_X1 U17685 ( .B1(n14111), .B2(n9716), .A(n14110), .ZN(P2_U2880) );
  NAND2_X1 U17686 ( .A1(n21022), .A2(n21060), .ZN(n14114) );
  OR2_X1 U17687 ( .A1(n21053), .A2(n21021), .ZN(n14144) );
  NAND2_X1 U17688 ( .A1(n14114), .A2(n14144), .ZN(n14117) );
  OR2_X1 U17689 ( .A1(n14120), .A2(n11830), .ZN(n20997) );
  INV_X1 U17690 ( .A(n20997), .ZN(n15683) );
  INV_X1 U17691 ( .A(n14195), .ZN(n14115) );
  INV_X1 U17692 ( .A(n20992), .ZN(n14194) );
  NOR2_X1 U17693 ( .A1(n14115), .A2(n14194), .ZN(n21061) );
  AOI22_X1 U17694 ( .A1(n14117), .A2(n21029), .B1(n15683), .B2(n21061), .ZN(
        n14145) );
  OAI22_X1 U17695 ( .A1(n15764), .A2(n14145), .B1(n15715), .B2(n14144), .ZN(
        n14116) );
  AOI21_X1 U17696 ( .B1(n14147), .B2(n21186), .A(n14116), .ZN(n14125) );
  INV_X1 U17697 ( .A(n14144), .ZN(n14123) );
  OAI21_X1 U17698 ( .B1(n20987), .B2(n14147), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14119) );
  INV_X1 U17699 ( .A(n14117), .ZN(n14118) );
  NAND2_X1 U17700 ( .A1(n14119), .A2(n14118), .ZN(n14122) );
  NAND2_X1 U17701 ( .A1(n14120), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21094) );
  NAND2_X1 U17702 ( .A1(n14121), .A2(n21094), .ZN(n14220) );
  NAND2_X1 U17703 ( .A1(n14148), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n14124) );
  OAI211_X1 U17704 ( .C1(n21191), .C2(n14151), .A(n14125), .B(n14124), .ZN(
        P1_U3103) );
  OAI22_X1 U17705 ( .A1(n15752), .A2(n14145), .B1(n15703), .B2(n14144), .ZN(
        n14126) );
  AOI21_X1 U17706 ( .B1(n14147), .B2(n21110), .A(n14126), .ZN(n14128) );
  NAND2_X1 U17707 ( .A1(n14148), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n14127) );
  OAI211_X1 U17708 ( .C1(n21113), .C2(n14151), .A(n14128), .B(n14127), .ZN(
        P1_U3100) );
  OAI22_X1 U17709 ( .A1(n15756), .A2(n14145), .B1(n15707), .B2(n14144), .ZN(
        n14129) );
  AOI21_X1 U17710 ( .B1(n14147), .B2(n21114), .A(n14129), .ZN(n14131) );
  NAND2_X1 U17711 ( .A1(n14148), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n14130) );
  OAI211_X1 U17712 ( .C1(n21117), .C2(n14151), .A(n14131), .B(n14130), .ZN(
        P1_U3101) );
  OAI22_X1 U17713 ( .A1(n15748), .A2(n14145), .B1(n15699), .B2(n14144), .ZN(
        n14132) );
  AOI21_X1 U17714 ( .B1(n14147), .B2(n21106), .A(n14132), .ZN(n14134) );
  NAND2_X1 U17715 ( .A1(n14148), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n14133) );
  OAI211_X1 U17716 ( .C1(n21109), .C2(n14151), .A(n14134), .B(n14133), .ZN(
        P1_U3099) );
  OAI22_X1 U17717 ( .A1(n15760), .A2(n14145), .B1(n15711), .B2(n14144), .ZN(
        n14135) );
  AOI21_X1 U17718 ( .B1(n14147), .B2(n21118), .A(n14135), .ZN(n14137) );
  NAND2_X1 U17719 ( .A1(n14148), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n14136) );
  OAI211_X1 U17720 ( .C1(n21121), .C2(n14151), .A(n14137), .B(n14136), .ZN(
        P1_U3102) );
  OAI22_X1 U17721 ( .A1(n15744), .A2(n14145), .B1(n15695), .B2(n14144), .ZN(
        n14138) );
  AOI21_X1 U17722 ( .B1(n14147), .B2(n21102), .A(n14138), .ZN(n14140) );
  NAND2_X1 U17723 ( .A1(n14148), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n14139) );
  OAI211_X1 U17724 ( .C1(n21105), .C2(n14151), .A(n14140), .B(n14139), .ZN(
        P1_U3098) );
  OAI22_X1 U17725 ( .A1(n15772), .A2(n14145), .B1(n15721), .B2(n14144), .ZN(
        n14141) );
  AOI21_X1 U17726 ( .B1(n14147), .B2(n21126), .A(n14141), .ZN(n14143) );
  NAND2_X1 U17727 ( .A1(n14148), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n14142) );
  OAI211_X1 U17728 ( .C1(n21131), .C2(n14151), .A(n14143), .B(n14142), .ZN(
        P1_U3104) );
  OAI22_X1 U17729 ( .A1(n15740), .A2(n14145), .B1(n15691), .B2(n14144), .ZN(
        n14146) );
  AOI21_X1 U17730 ( .B1(n14147), .B2(n21150), .A(n14146), .ZN(n14150) );
  NAND2_X1 U17731 ( .A1(n14148), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n14149) );
  OAI211_X1 U17732 ( .C1(n21153), .C2(n14151), .A(n14150), .B(n14149), .ZN(
        P1_U3097) );
  OR2_X1 U17733 ( .A1(n14050), .A2(n14152), .ZN(n14153) );
  AND2_X1 U17734 ( .A1(n9638), .A2(n14153), .ZN(n16695) );
  NAND2_X1 U17735 ( .A1(n16695), .A2(n16104), .ZN(n14158) );
  INV_X1 U17736 ( .A(n14154), .ZN(n14155) );
  OAI211_X1 U17737 ( .C1(n14156), .C2(n14155), .A(n14181), .B(n16150), .ZN(
        n14157) );
  OAI211_X1 U17738 ( .C1(n16104), .C2(n10718), .A(n14158), .B(n14157), .ZN(
        P2_U2874) );
  XNOR2_X1 U17739 ( .A(n9717), .B(n14159), .ZN(n20797) );
  INV_X1 U17740 ( .A(n20797), .ZN(n14161) );
  OAI222_X1 U17741 ( .A1(n15163), .A2(n14161), .B1(n14160), .B2(n15150), .C1(
        n15117), .C2(n15161), .ZN(P1_U2899) );
  AND2_X1 U17742 ( .A1(n13934), .A2(n14162), .ZN(n14163) );
  OR2_X1 U17743 ( .A1(n14163), .A2(n9608), .ZN(n16689) );
  INV_X1 U17744 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n15071) );
  OR2_X1 U17745 ( .A1(n14164), .A2(n15071), .ZN(n14166) );
  NAND2_X1 U17746 ( .A1(n16872), .A2(BUF2_REG_14__SCAN_IN), .ZN(n14165) );
  NAND2_X1 U17747 ( .A1(n14166), .A2(n14165), .ZN(n19934) );
  AOI22_X1 U17748 ( .A1(n16279), .A2(n19934), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19887), .ZN(n14167) );
  OAI21_X1 U17749 ( .B1(n16689), .B2(n16275), .A(n14167), .ZN(P2_U2905) );
  OAI21_X1 U17750 ( .B1(n14169), .B2(n14168), .A(n17203), .ZN(n20894) );
  OAI222_X1 U17751 ( .A1(n20894), .A2(n15068), .B1(n20800), .B2(n20768), .C1(
        n14170), .C2(n15070), .ZN(P1_U2868) );
  OR2_X1 U17752 ( .A1(n14173), .A2(n14172), .ZN(n14174) );
  NAND2_X1 U17753 ( .A1(n14171), .A2(n14174), .ZN(n20750) );
  NAND2_X1 U17754 ( .A1(n14175), .A2(n14176), .ZN(n14177) );
  AND2_X1 U17755 ( .A1(n14259), .A2(n14177), .ZN(n20746) );
  AOI22_X1 U17756 ( .A1(n20795), .A2(n20746), .B1(n15065), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n14178) );
  OAI21_X1 U17757 ( .B1(n20750), .B2(n15070), .A(n14178), .ZN(P1_U2866) );
  OR2_X1 U17758 ( .A1(n9638), .A2(n14179), .ZN(n14253) );
  NAND2_X1 U17759 ( .A1(n9638), .A2(n14179), .ZN(n14180) );
  INV_X1 U17760 ( .A(n16682), .ZN(n14187) );
  AOI21_X1 U17761 ( .B1(n14181), .B2(n14182), .A(n9716), .ZN(n14185) );
  INV_X1 U17762 ( .A(n14182), .ZN(n14183) );
  AOI22_X1 U17763 ( .A1(n14185), .A2(n14430), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n16154), .ZN(n14186) );
  OAI21_X1 U17764 ( .B1(n14187), .B2(n16154), .A(n14186), .ZN(P2_U2873) );
  OAI222_X1 U17765 ( .A1(n15163), .A2(n20750), .B1(n15112), .B2(n15161), .C1(
        n15150), .C2(n11965), .ZN(P1_U2898) );
  AOI21_X1 U17766 ( .B1(n20972), .B2(n14193), .A(n20709), .ZN(n14188) );
  AOI21_X1 U17767 ( .B1(n15728), .B2(n21060), .A(n14188), .ZN(n14189) );
  NOR2_X1 U17768 ( .A1(n14189), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n14192) );
  INV_X1 U17769 ( .A(n14190), .ZN(n14191) );
  NOR2_X1 U17770 ( .A1(n21053), .A2(n14191), .ZN(n20966) );
  NAND2_X1 U17771 ( .A1(n20969), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n14199) );
  INV_X1 U17772 ( .A(n21060), .ZN(n21092) );
  NOR2_X1 U17773 ( .A1(n21092), .A2(n21141), .ZN(n14196) );
  OR2_X1 U17774 ( .A1(n14195), .A2(n14194), .ZN(n15687) );
  INV_X1 U17775 ( .A(n15687), .ZN(n15682) );
  INV_X1 U17776 ( .A(n21094), .ZN(n15729) );
  AOI22_X1 U17777 ( .A1(n15728), .A2(n14196), .B1(n15682), .B2(n15729), .ZN(
        n20957) );
  INV_X1 U17778 ( .A(n20966), .ZN(n14203) );
  OAI22_X1 U17779 ( .A1(n15756), .A2(n20957), .B1(n15707), .B2(n14203), .ZN(
        n14197) );
  AOI21_X1 U17780 ( .B1(n20968), .B2(n21174), .A(n14197), .ZN(n14198) );
  OAI211_X1 U17781 ( .C1(n21177), .C2(n20972), .A(n14199), .B(n14198), .ZN(
        P1_U3069) );
  NAND2_X1 U17782 ( .A1(n20969), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n14202) );
  OAI22_X1 U17783 ( .A1(n15760), .A2(n20957), .B1(n15711), .B2(n14203), .ZN(
        n14200) );
  AOI21_X1 U17784 ( .B1(n20968), .B2(n21180), .A(n14200), .ZN(n14201) );
  OAI211_X1 U17785 ( .C1(n21183), .C2(n20972), .A(n14202), .B(n14201), .ZN(
        P1_U3070) );
  NAND2_X1 U17786 ( .A1(n20969), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n14206) );
  OAI22_X1 U17787 ( .A1(n15748), .A2(n20957), .B1(n15699), .B2(n14203), .ZN(
        n14204) );
  AOI21_X1 U17788 ( .B1(n20968), .B2(n21162), .A(n14204), .ZN(n14205) );
  OAI211_X1 U17789 ( .C1(n21165), .C2(n20972), .A(n14206), .B(n14205), .ZN(
        P1_U3067) );
  AND2_X1 U17790 ( .A1(n14208), .A2(n14207), .ZN(n14209) );
  OR2_X1 U17791 ( .A1(n14209), .A2(n16148), .ZN(n16756) );
  INV_X1 U17792 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14210) );
  NOR2_X1 U17793 ( .A1(n14211), .A2(n14210), .ZN(n14213) );
  NAND2_X1 U17794 ( .A1(n14213), .A2(n14212), .ZN(n16149) );
  OAI211_X1 U17795 ( .C1(n14213), .C2(n14212), .A(n16149), .B(n16150), .ZN(
        n14215) );
  NAND2_X1 U17796 ( .A1(n16154), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14214) );
  OAI211_X1 U17797 ( .C1(n16756), .C2(n16154), .A(n14215), .B(n14214), .ZN(
        P2_U2879) );
  OAI21_X1 U17798 ( .B1(n14247), .B2(n20951), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14216) );
  NAND2_X1 U17799 ( .A1(n14216), .A2(n21029), .ZN(n14223) );
  INV_X1 U17800 ( .A(n14223), .ZN(n14217) );
  NOR2_X1 U17801 ( .A1(n15681), .A2(n21060), .ZN(n14222) );
  NOR2_X1 U17802 ( .A1(n20992), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15730) );
  OR2_X1 U17803 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14218), .ZN(
        n14245) );
  OAI22_X1 U17804 ( .A1(n15703), .A2(n14245), .B1(n14244), .B2(n21113), .ZN(
        n14219) );
  AOI21_X1 U17805 ( .B1(n14247), .B2(n21110), .A(n14219), .ZN(n14225) );
  NOR2_X1 U17806 ( .A1(n15730), .A2(n11830), .ZN(n15733) );
  AOI211_X1 U17807 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n14245), .A(n15733), 
        .B(n14220), .ZN(n14221) );
  NAND2_X1 U17808 ( .A1(n14248), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n14224) );
  OAI211_X1 U17809 ( .C1(n14251), .C2(n15752), .A(n14225), .B(n14224), .ZN(
        P1_U3052) );
  OAI22_X1 U17810 ( .A1(n15711), .A2(n14245), .B1(n14244), .B2(n21121), .ZN(
        n14226) );
  AOI21_X1 U17811 ( .B1(n14247), .B2(n21118), .A(n14226), .ZN(n14228) );
  NAND2_X1 U17812 ( .A1(n14248), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n14227) );
  OAI211_X1 U17813 ( .C1(n14251), .C2(n15760), .A(n14228), .B(n14227), .ZN(
        P1_U3054) );
  OAI22_X1 U17814 ( .A1(n15715), .A2(n14245), .B1(n14244), .B2(n21191), .ZN(
        n14229) );
  AOI21_X1 U17815 ( .B1(n14247), .B2(n21186), .A(n14229), .ZN(n14231) );
  NAND2_X1 U17816 ( .A1(n14248), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n14230) );
  OAI211_X1 U17817 ( .C1(n14251), .C2(n15764), .A(n14231), .B(n14230), .ZN(
        P1_U3055) );
  OAI22_X1 U17818 ( .A1(n15699), .A2(n14245), .B1(n14244), .B2(n21109), .ZN(
        n14232) );
  AOI21_X1 U17819 ( .B1(n14247), .B2(n21106), .A(n14232), .ZN(n14234) );
  NAND2_X1 U17820 ( .A1(n14248), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n14233) );
  OAI211_X1 U17821 ( .C1(n14251), .C2(n15748), .A(n14234), .B(n14233), .ZN(
        P1_U3051) );
  OAI22_X1 U17822 ( .A1(n15707), .A2(n14245), .B1(n14244), .B2(n21117), .ZN(
        n14235) );
  AOI21_X1 U17823 ( .B1(n14247), .B2(n21114), .A(n14235), .ZN(n14237) );
  NAND2_X1 U17824 ( .A1(n14248), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n14236) );
  OAI211_X1 U17825 ( .C1(n14251), .C2(n15756), .A(n14237), .B(n14236), .ZN(
        P1_U3053) );
  OAI22_X1 U17826 ( .A1(n15695), .A2(n14245), .B1(n14244), .B2(n21105), .ZN(
        n14238) );
  AOI21_X1 U17827 ( .B1(n14247), .B2(n21102), .A(n14238), .ZN(n14240) );
  NAND2_X1 U17828 ( .A1(n14248), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n14239) );
  OAI211_X1 U17829 ( .C1(n14251), .C2(n15744), .A(n14240), .B(n14239), .ZN(
        P1_U3050) );
  OAI22_X1 U17830 ( .A1(n15691), .A2(n14245), .B1(n14244), .B2(n21153), .ZN(
        n14241) );
  AOI21_X1 U17831 ( .B1(n14247), .B2(n21150), .A(n14241), .ZN(n14243) );
  NAND2_X1 U17832 ( .A1(n14248), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n14242) );
  OAI211_X1 U17833 ( .C1(n14251), .C2(n15740), .A(n14243), .B(n14242), .ZN(
        P1_U3049) );
  OAI22_X1 U17834 ( .A1(n15721), .A2(n14245), .B1(n14244), .B2(n21131), .ZN(
        n14246) );
  AOI21_X1 U17835 ( .B1(n14247), .B2(n21126), .A(n14246), .ZN(n14250) );
  NAND2_X1 U17836 ( .A1(n14248), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n14249) );
  OAI211_X1 U17837 ( .C1(n14251), .C2(n15772), .A(n14250), .B(n14249), .ZN(
        P1_U3056) );
  AND2_X1 U17838 ( .A1(n14253), .A2(n14252), .ZN(n14255) );
  OR2_X1 U17839 ( .A1(n14255), .A2(n14254), .ZN(n19795) );
  XOR2_X1 U17840 ( .A(n14429), .B(n14430), .Z(n14256) );
  AOI22_X1 U17841 ( .A1(n14256), .A2(n16150), .B1(n16154), .B2(
        P2_EBX_REG_15__SCAN_IN), .ZN(n14257) );
  OAI21_X1 U17842 ( .B1(n19795), .B2(n16154), .A(n14257), .ZN(P2_U2872) );
  XOR2_X1 U17843 ( .A(n14258), .B(n14171), .Z(n20737) );
  INV_X1 U17844 ( .A(n20737), .ZN(n14262) );
  AOI21_X1 U17845 ( .B1(n14260), .B2(n14259), .A(n14267), .ZN(n20730) );
  AOI22_X1 U17846 ( .A1(n20730), .A2(n20795), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n15065), .ZN(n14261) );
  OAI21_X1 U17847 ( .B1(n14262), .B2(n15070), .A(n14261), .ZN(P1_U2865) );
  OAI222_X1 U17848 ( .A1(n15163), .A2(n14262), .B1(n15150), .B2(n11974), .C1(
        n15161), .C2(n15107), .ZN(P1_U2897) );
  OAI21_X1 U17849 ( .B1(n14171), .B2(n14258), .A(n14263), .ZN(n14265) );
  AND2_X1 U17850 ( .A1(n14265), .A2(n14264), .ZN(n15389) );
  INV_X1 U17851 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n21438) );
  OAI222_X1 U17852 ( .A1(n15163), .A2(n15018), .B1(n15103), .B2(n15161), .C1(
        n15150), .C2(n21438), .ZN(P1_U2896) );
  OR2_X1 U17853 ( .A1(n14267), .A2(n14266), .ZN(n14268) );
  AND2_X1 U17854 ( .A1(n14268), .A2(n14274), .ZN(n15605) );
  INV_X1 U17855 ( .A(n15605), .ZN(n14269) );
  OAI222_X1 U17856 ( .A1(n14269), .A2(n15068), .B1(n20800), .B2(n12846), .C1(
        n15018), .C2(n15070), .ZN(P1_U2864) );
  AOI21_X1 U17857 ( .B1(n14271), .B2(n14264), .A(n14270), .ZN(n14272) );
  INV_X1 U17858 ( .A(n14272), .ZN(n15381) );
  NAND2_X1 U17859 ( .A1(n14274), .A2(n14273), .ZN(n14275) );
  AND2_X1 U17860 ( .A1(n14282), .A2(n14275), .ZN(n17185) );
  AOI22_X1 U17861 ( .A1(n17185), .A2(n20795), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n15065), .ZN(n14276) );
  OAI21_X1 U17862 ( .B1(n15381), .B2(n15070), .A(n14276), .ZN(P1_U2863) );
  INV_X1 U17863 ( .A(DATAI_9_), .ZN(n14277) );
  MUX2_X1 U17864 ( .A(n14277), .B(n17337), .S(n15085), .Z(n20828) );
  INV_X1 U17865 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n14278) );
  OAI222_X1 U17866 ( .A1(n15163), .A2(n15381), .B1(n20828), .B2(n15161), .C1(
        n14278), .C2(n15150), .ZN(P1_U2895) );
  OAI21_X1 U17867 ( .B1(n14270), .B2(n14280), .A(n14279), .ZN(n17155) );
  AND2_X1 U17868 ( .A1(n14282), .A2(n14281), .ZN(n14283) );
  NOR2_X1 U17869 ( .A1(n14994), .A2(n14283), .ZN(n17151) );
  AOI22_X1 U17870 ( .A1(n17151), .A2(n20795), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n15065), .ZN(n14284) );
  OAI21_X1 U17871 ( .B1(n17155), .B2(n15070), .A(n14284), .ZN(P1_U2862) );
  INV_X1 U17872 ( .A(DATAI_10_), .ZN(n14286) );
  NAND2_X1 U17873 ( .A1(n15085), .A2(BUF1_REG_10__SCAN_IN), .ZN(n14285) );
  OAI21_X1 U17874 ( .B1(n15085), .B2(n14286), .A(n14285), .ZN(n20831) );
  AOI22_X1 U17875 ( .A1(n15155), .A2(n20831), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15154), .ZN(n14287) );
  OAI21_X1 U17876 ( .B1(n17155), .B2(n15163), .A(n14287), .ZN(P1_U2894) );
  NAND3_X1 U17877 ( .A1(n9584), .A2(n19493), .A3(n21439), .ZN(n19046) );
  NOR2_X1 U17878 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n19046), .ZN(n14288) );
  NAND3_X1 U17879 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19648)
         );
  OAI21_X1 U17880 ( .B1(n14288), .B2(n19648), .A(n19334), .ZN(n19052) );
  INV_X1 U17881 ( .A(n19052), .ZN(n14289) );
  INV_X1 U17882 ( .A(n18628), .ZN(n18693) );
  NOR2_X1 U17883 ( .A1(n18693), .A2(n19699), .ZN(n17057) );
  AOI21_X1 U17884 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n17057), .ZN(n17058) );
  NOR2_X1 U17885 ( .A1(n14289), .A2(n17058), .ZN(n14291) );
  NAND2_X1 U17886 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19195), .ZN(n19219) );
  NAND2_X1 U17887 ( .A1(n19219), .A2(n19052), .ZN(n17056) );
  OR2_X1 U17888 ( .A1(n19108), .A2(n17056), .ZN(n14290) );
  MUX2_X1 U17889 ( .A(n14291), .B(n14290), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  XNOR2_X1 U17890 ( .A(n16031), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14292) );
  XNOR2_X1 U17891 ( .A(n14337), .B(n14292), .ZN(n19957) );
  OAI21_X1 U17892 ( .B1(n14294), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n14293), .ZN(n19971) );
  NAND2_X1 U17893 ( .A1(n19941), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n19968) );
  OAI21_X1 U17894 ( .B1(n16550), .B2(n19971), .A(n19968), .ZN(n14295) );
  AOI21_X1 U17895 ( .B1(n16510), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14295), .ZN(n14296) );
  OAI21_X1 U17896 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16544), .A(
        n14296), .ZN(n14297) );
  AOI21_X1 U17897 ( .B1(n10145), .B2(n19957), .A(n14297), .ZN(n14298) );
  OAI21_X1 U17898 ( .B1(n16831), .B2(n19950), .A(n14298), .ZN(P2_U3013) );
  NAND2_X1 U17899 ( .A1(n14299), .A2(n16293), .ZN(n14304) );
  INV_X1 U17900 ( .A(n14300), .ZN(n14301) );
  NOR2_X1 U17901 ( .A1(n14302), .A2(n14301), .ZN(n14303) );
  XNOR2_X1 U17902 ( .A(n14304), .B(n14303), .ZN(n14428) );
  XNOR2_X1 U17903 ( .A(n16298), .B(n11515), .ZN(n14426) );
  NOR2_X1 U17904 ( .A1(n16491), .A2(n20616), .ZN(n14423) );
  INV_X1 U17905 ( .A(n14423), .ZN(n14308) );
  INV_X1 U17906 ( .A(n14305), .ZN(n16558) );
  AOI21_X1 U17907 ( .B1(n16558), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14307) );
  INV_X1 U17908 ( .A(n14309), .ZN(n14310) );
  OAI21_X1 U17909 ( .B1(n14701), .B2(n16782), .A(n14310), .ZN(n14311) );
  OAI21_X1 U17910 ( .B1(n14428), .B2(n16802), .A(n14312), .ZN(P2_U3016) );
  INV_X1 U17911 ( .A(n14313), .ZN(n14314) );
  AOI21_X1 U17912 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n11096), .A(
        n14315), .ZN(n14316) );
  INV_X1 U17913 ( .A(n16326), .ZN(n16334) );
  INV_X1 U17914 ( .A(n14317), .ZN(n14318) );
  NAND2_X1 U17915 ( .A1(n15795), .A2(n11096), .ZN(n14319) );
  XNOR2_X1 U17916 ( .A(n14319), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14320) );
  XNOR2_X1 U17917 ( .A(n14321), .B(n14320), .ZN(n16311) );
  INV_X1 U17918 ( .A(n14322), .ZN(n14325) );
  INV_X1 U17919 ( .A(n14323), .ZN(n14324) );
  OAI21_X1 U17920 ( .B1(n14325), .B2(n14324), .A(n15779), .ZN(n16166) );
  INV_X1 U17921 ( .A(n15775), .ZN(n14327) );
  AOI21_X1 U17922 ( .B1(n14328), .B2(n14326), .A(n14327), .ZN(n16303) );
  NAND2_X1 U17923 ( .A1(n16303), .A2(n19967), .ZN(n14334) );
  INV_X1 U17924 ( .A(n16552), .ZN(n14330) );
  NOR2_X1 U17925 ( .A1(n14330), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16568) );
  INV_X1 U17926 ( .A(n16554), .ZN(n14332) );
  INV_X1 U17927 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n15787) );
  NOR2_X1 U17928 ( .A1(n16491), .A2(n15787), .ZN(n16304) );
  NOR3_X1 U17929 ( .A1(n14330), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n14329), .ZN(n14331) );
  AOI211_X1 U17930 ( .C1(n14332), .C2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16304), .B(n14331), .ZN(n14333) );
  OAI211_X1 U17931 ( .C1(n17237), .C2(n16166), .A(n14334), .B(n14333), .ZN(
        n14335) );
  AOI21_X1 U17932 ( .B1(n16799), .B2(n16309), .A(n14335), .ZN(n14336) );
  OAI21_X1 U17933 ( .B1(n16311), .B2(n16802), .A(n14336), .ZN(P2_U3018) );
  OAI21_X1 U17934 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n16042), .A(
        n14337), .ZN(n17242) );
  INV_X1 U17935 ( .A(n17242), .ZN(n14340) );
  INV_X1 U17936 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19739) );
  NOR2_X1 U17937 ( .A1(n16491), .A2(n19739), .ZN(n17244) );
  XNOR2_X1 U17938 ( .A(n14338), .B(n19964), .ZN(n17239) );
  NOR2_X1 U17939 ( .A1(n16550), .A2(n17239), .ZN(n14339) );
  AOI211_X1 U17940 ( .C1(n10145), .C2(n14340), .A(n17244), .B(n14339), .ZN(
        n14343) );
  OAI21_X1 U17941 ( .B1(n16510), .B2(n14341), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14342) );
  OAI211_X1 U17942 ( .C1(n19950), .C2(n14344), .A(n14343), .B(n14342), .ZN(
        P2_U3014) );
  NAND2_X1 U17943 ( .A1(n14388), .A2(n14345), .ZN(n14359) );
  INV_X1 U17944 ( .A(n14346), .ZN(n14350) );
  NAND2_X1 U17945 ( .A1(n14347), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14348) );
  NAND2_X1 U17946 ( .A1(n14352), .A2(n14351), .ZN(n16425) );
  NAND2_X1 U17947 ( .A1(n16418), .A2(n16406), .ZN(n14353) );
  NOR3_X1 U17948 ( .A1(n14705), .A2(n14709), .A3(n16405), .ZN(n14356) );
  OR2_X1 U17949 ( .A1(n14356), .A2(n14355), .ZN(n14357) );
  INV_X1 U17950 ( .A(n16388), .ZN(n14358) );
  INV_X1 U17951 ( .A(n14361), .ZN(n14722) );
  OAI21_X1 U17952 ( .B1(n16394), .B2(n16650), .A(n14363), .ZN(n14364) );
  AND2_X1 U17953 ( .A1(n16112), .A2(n14365), .ZN(n14367) );
  OR2_X1 U17954 ( .A1(n14367), .A2(n14401), .ZN(n19754) );
  NOR2_X1 U17955 ( .A1(n19754), .A2(n16782), .ZN(n14379) );
  INV_X1 U17956 ( .A(n14368), .ZN(n14372) );
  NAND2_X1 U17957 ( .A1(n14369), .A2(n14370), .ZN(n14371) );
  NAND2_X1 U17958 ( .A1(n14372), .A2(n14371), .ZN(n19753) );
  INV_X1 U17959 ( .A(n16738), .ZN(n16669) );
  NOR2_X1 U17960 ( .A1(n16669), .A2(n14373), .ZN(n16639) );
  NAND2_X1 U17961 ( .A1(n16639), .A2(n16650), .ZN(n16649) );
  INV_X1 U17962 ( .A(n14373), .ZN(n14374) );
  NAND2_X1 U17963 ( .A1(n16740), .A2(n14374), .ZN(n14375) );
  NAND2_X1 U17964 ( .A1(n16685), .A2(n14375), .ZN(n16651) );
  NAND2_X1 U17965 ( .A1(n16649), .A2(n16651), .ZN(n14409) );
  NOR2_X1 U17966 ( .A1(n16491), .A2(n20596), .ZN(n14381) );
  INV_X1 U17967 ( .A(n16639), .ZN(n14406) );
  NOR3_X1 U17968 ( .A1(n14406), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n16650), .ZN(n14376) );
  AOI211_X1 U17969 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n14409), .A(
        n14381), .B(n14376), .ZN(n14377) );
  OAI21_X1 U17970 ( .B1(n17237), .B2(n19753), .A(n14377), .ZN(n14378) );
  AOI211_X1 U17971 ( .C1(n14385), .C2(n16799), .A(n14379), .B(n14378), .ZN(
        n14380) );
  OAI21_X1 U17972 ( .B1(n14387), .B2(n16802), .A(n14380), .ZN(P2_U3027) );
  AOI21_X1 U17973 ( .B1(n16510), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n14381), .ZN(n14383) );
  NAND2_X1 U17974 ( .A1(n19943), .A2(n19747), .ZN(n14382) );
  OAI211_X1 U17975 ( .C1(n19754), .C2(n19950), .A(n14383), .B(n14382), .ZN(
        n14384) );
  AOI21_X1 U17976 ( .B1(n14385), .B2(n19945), .A(n14384), .ZN(n14386) );
  INV_X1 U17977 ( .A(n14390), .ZN(n14391) );
  INV_X1 U17978 ( .A(n14392), .ZN(n16376) );
  NOR2_X1 U17979 ( .A1(n14393), .A2(n16376), .ZN(n14394) );
  XNOR2_X1 U17980 ( .A(n14395), .B(n14394), .ZN(n14420) );
  AOI21_X1 U17981 ( .B1(n14398), .B2(n14397), .A(n16385), .ZN(n14418) );
  OAI21_X1 U17982 ( .B1(n14401), .B2(n14400), .A(n14399), .ZN(n16107) );
  NOR2_X1 U17983 ( .A1(n16107), .A2(n16782), .ZN(n14412) );
  OAI21_X1 U17984 ( .B1(n14368), .B2(n14404), .A(n14403), .ZN(n16232) );
  NOR2_X1 U17985 ( .A1(n16491), .A2(n14405), .ZN(n14415) );
  NOR2_X1 U17986 ( .A1(n16638), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14407) );
  AOI211_X1 U17987 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n14407), .B(n14406), .ZN(
        n14408) );
  AOI211_X1 U17988 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n14409), .A(
        n14415), .B(n14408), .ZN(n14410) );
  OAI21_X1 U17989 ( .B1(n17237), .B2(n16232), .A(n14410), .ZN(n14411) );
  AOI211_X1 U17990 ( .C1(n14418), .C2(n16799), .A(n14412), .B(n14411), .ZN(
        n14413) );
  OAI21_X1 U17991 ( .B1(n14420), .B2(n16802), .A(n14413), .ZN(P2_U3026) );
  NOR2_X1 U17992 ( .A1(n16544), .A2(n15896), .ZN(n14414) );
  AOI211_X1 U17993 ( .C1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n16510), .A(
        n14415), .B(n14414), .ZN(n14416) );
  OAI21_X1 U17994 ( .B1(n16107), .B2(n19950), .A(n14416), .ZN(n14417) );
  AOI21_X1 U17995 ( .B1(n14418), .B2(n19945), .A(n14417), .ZN(n14419) );
  OAI21_X1 U17996 ( .B1(n14420), .B2(n16483), .A(n14419), .ZN(P2_U2994) );
  NOR2_X1 U17997 ( .A1(n16544), .A2(n14421), .ZN(n14422) );
  AOI211_X1 U17998 ( .C1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .C2(n16510), .A(
        n14423), .B(n14422), .ZN(n14424) );
  OAI21_X1 U17999 ( .B1(n14701), .B2(n19950), .A(n14424), .ZN(n14425) );
  AOI21_X1 U18000 ( .B1(n19945), .B2(n14426), .A(n14425), .ZN(n14427) );
  OAI21_X1 U18001 ( .B1(n14428), .B2(n16483), .A(n14427), .ZN(P2_U2984) );
  AOI22_X1 U18002 ( .A1(n14530), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14529), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14434) );
  AOI22_X1 U18003 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14433) );
  AOI22_X1 U18004 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n14533), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14432) );
  AOI22_X1 U18005 ( .A1(n10620), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10888), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14431) );
  NAND4_X1 U18006 ( .A1(n14434), .A2(n14433), .A3(n14432), .A4(n14431), .ZN(
        n14440) );
  AOI22_X1 U18007 ( .A1(n14478), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14438) );
  AOI22_X1 U18008 ( .A1(n10894), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9598), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14437) );
  AOI22_X1 U18009 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14436) );
  AOI22_X1 U18010 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14435) );
  NAND4_X1 U18011 ( .A1(n14438), .A2(n14437), .A3(n14436), .A4(n14435), .ZN(
        n14439) );
  OR2_X1 U18012 ( .A1(n14440), .A2(n14439), .ZN(n16126) );
  AOI22_X1 U18013 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n14530), .B1(
        n14529), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14444) );
  AOI22_X1 U18014 ( .A1(n9595), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14443) );
  AOI22_X1 U18015 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n14533), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14442) );
  AOI22_X1 U18016 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n10888), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14441) );
  NAND4_X1 U18017 ( .A1(n14444), .A2(n14443), .A3(n14442), .A4(n14441), .ZN(
        n14450) );
  AOI22_X1 U18018 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n14478), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14448) );
  AOI22_X1 U18019 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n9598), .B1(
        n10894), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14447) );
  AOI22_X1 U18020 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14446) );
  AOI22_X1 U18021 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14445) );
  NAND4_X1 U18022 ( .A1(n14448), .A2(n14447), .A3(n14446), .A4(n14445), .ZN(
        n14449) );
  NOR2_X1 U18023 ( .A1(n14450), .A2(n14449), .ZN(n16121) );
  INV_X1 U18024 ( .A(n16121), .ZN(n14451) );
  NAND2_X1 U18025 ( .A1(n14452), .A2(n14451), .ZN(n16115) );
  INV_X1 U18026 ( .A(n16115), .ZN(n16120) );
  AOI22_X1 U18027 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n14530), .B1(
        n14529), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14456) );
  AOI22_X1 U18028 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14455) );
  AOI22_X1 U18029 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n14533), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14454) );
  AOI22_X1 U18030 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n10888), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14453) );
  NAND4_X1 U18031 ( .A1(n14456), .A2(n14455), .A3(n14454), .A4(n14453), .ZN(
        n14462) );
  AOI22_X1 U18032 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n14539), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14460) );
  AOI22_X1 U18033 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n9598), .B1(
        n10894), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14459) );
  AOI22_X1 U18034 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14458) );
  AOI22_X1 U18035 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14457) );
  NAND4_X1 U18036 ( .A1(n14460), .A2(n14459), .A3(n14458), .A4(n14457), .ZN(
        n14461) );
  NOR2_X1 U18037 ( .A1(n14462), .A2(n14461), .ZN(n16116) );
  INV_X1 U18038 ( .A(n16116), .ZN(n14463) );
  AOI22_X1 U18039 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n14530), .B1(
        n14529), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14467) );
  AOI22_X1 U18040 ( .A1(n9595), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14466) );
  AOI22_X1 U18041 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n14533), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14465) );
  AOI22_X1 U18042 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n10620), .B1(
        n10888), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14464) );
  NAND4_X1 U18043 ( .A1(n14467), .A2(n14466), .A3(n14465), .A4(n14464), .ZN(
        n14473) );
  AOI22_X1 U18044 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n14539), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14471) );
  AOI22_X1 U18045 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n9597), .B1(
        n10894), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14470) );
  AOI22_X1 U18046 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14469) );
  AOI22_X1 U18047 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14468) );
  NAND4_X1 U18048 ( .A1(n14471), .A2(n14470), .A3(n14469), .A4(n14468), .ZN(
        n14472) );
  NOR2_X1 U18049 ( .A1(n14473), .A2(n14472), .ZN(n16108) );
  AOI22_X1 U18050 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n14530), .B1(
        n14529), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14477) );
  AOI22_X1 U18051 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14476) );
  AOI22_X1 U18052 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n14533), .B1(
        n10631), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14475) );
  AOI22_X1 U18053 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n10888), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14474) );
  NAND4_X1 U18054 ( .A1(n14477), .A2(n14476), .A3(n14475), .A4(n14474), .ZN(
        n14484) );
  AOI22_X1 U18055 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n14478), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14482) );
  AOI22_X1 U18056 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n9597), .B1(
        n10894), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14481) );
  AOI22_X1 U18057 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14480) );
  AOI22_X1 U18058 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14479) );
  NAND4_X1 U18059 ( .A1(n14482), .A2(n14481), .A3(n14480), .A4(n14479), .ZN(
        n14483) );
  OR2_X1 U18060 ( .A1(n14484), .A2(n14483), .ZN(n16102) );
  AOI22_X1 U18061 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n14530), .B1(
        n14529), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14488) );
  AOI22_X1 U18062 ( .A1(n9595), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14487) );
  AOI22_X1 U18063 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n14533), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14486) );
  AOI22_X1 U18064 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10888), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14485) );
  NAND4_X1 U18065 ( .A1(n14488), .A2(n14487), .A3(n14486), .A4(n14485), .ZN(
        n14494) );
  AOI22_X1 U18066 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n14539), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14492) );
  AOI22_X1 U18067 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n9598), .B1(
        n10894), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14491) );
  AOI22_X1 U18068 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14490) );
  AOI22_X1 U18069 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14489) );
  NAND4_X1 U18070 ( .A1(n14492), .A2(n14491), .A3(n14490), .A4(n14489), .ZN(
        n14493) );
  NOR2_X1 U18071 ( .A1(n14494), .A2(n14493), .ZN(n16095) );
  INV_X1 U18072 ( .A(n16095), .ZN(n14505) );
  AOI22_X1 U18073 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n14530), .B1(
        n14529), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14498) );
  AOI22_X1 U18074 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14497) );
  AOI22_X1 U18075 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n14533), .B1(
        n14532), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14496) );
  AOI22_X1 U18076 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n10888), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14495) );
  NAND4_X1 U18077 ( .A1(n14498), .A2(n14497), .A3(n14496), .A4(n14495), .ZN(
        n14504) );
  AOI22_X1 U18078 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n14539), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14502) );
  AOI22_X1 U18079 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n9597), .B1(
        n10894), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14501) );
  AOI22_X1 U18080 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n10621), .B1(
        n14541), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14500) );
  AOI22_X1 U18081 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n10622), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14499) );
  NAND4_X1 U18082 ( .A1(n14502), .A2(n14501), .A3(n14500), .A4(n14499), .ZN(
        n14503) );
  OR2_X1 U18083 ( .A1(n14504), .A2(n14503), .ZN(n16098) );
  AND2_X1 U18084 ( .A1(n14505), .A2(n16098), .ZN(n14506) );
  AND2_X1 U18085 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14508) );
  OR2_X1 U18086 ( .A1(n14508), .A2(n14507), .ZN(n14677) );
  INV_X1 U18087 ( .A(n14677), .ZN(n14647) );
  NAND2_X1 U18088 ( .A1(n14668), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n14511) );
  NAND2_X1 U18089 ( .A1(n16854), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n14510) );
  AND3_X1 U18090 ( .A1(n14647), .A2(n14511), .A3(n14510), .ZN(n14520) );
  AOI22_X1 U18091 ( .A1(n14682), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14680), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14519) );
  AOI22_X1 U18092 ( .A1(n14681), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14679), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14518) );
  INV_X1 U18093 ( .A(n14516), .ZN(n14675) );
  INV_X1 U18094 ( .A(n14675), .ZN(n14667) );
  AOI22_X1 U18095 ( .A1(n14683), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14667), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14517) );
  NAND4_X1 U18096 ( .A1(n14520), .A2(n14519), .A3(n14518), .A4(n14517), .ZN(
        n14528) );
  AOI22_X1 U18097 ( .A1(n14682), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14680), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14526) );
  NAND2_X1 U18098 ( .A1(n14668), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14522) );
  NAND2_X1 U18099 ( .A1(n16854), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n14521) );
  AND3_X1 U18100 ( .A1(n14522), .A2(n14677), .A3(n14521), .ZN(n14525) );
  AOI22_X1 U18101 ( .A1(n14681), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14679), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14524) );
  AOI22_X1 U18102 ( .A1(n14683), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14667), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14523) );
  NAND4_X1 U18103 ( .A1(n14526), .A2(n14525), .A3(n14524), .A4(n14523), .ZN(
        n14527) );
  NAND2_X1 U18104 ( .A1(n14528), .A2(n14527), .ZN(n14571) );
  AOI22_X1 U18105 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n14530), .B1(
        n14529), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14537) );
  AOI22_X1 U18106 ( .A1(n14532), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14531), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14536) );
  AOI22_X1 U18107 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n14533), .B1(
        n9595), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14535) );
  AOI22_X1 U18108 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n9597), .B1(
        n10888), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14534) );
  NAND4_X1 U18109 ( .A1(n14537), .A2(n14536), .A3(n14535), .A4(n14534), .ZN(
        n14547) );
  AOI22_X1 U18110 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n14539), .B1(
        n14538), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14545) );
  AOI22_X1 U18111 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10894), .B1(
        n10620), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14544) );
  AOI22_X1 U18112 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10621), .B1(
        n10622), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14543) );
  AOI22_X1 U18113 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14541), .B1(
        n10623), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14542) );
  NAND4_X1 U18114 ( .A1(n14545), .A2(n14544), .A3(n14543), .A4(n14542), .ZN(
        n14546) );
  NOR2_X1 U18115 ( .A1(n14547), .A2(n14546), .ZN(n14567) );
  INV_X1 U18116 ( .A(n14567), .ZN(n14564) );
  NAND2_X1 U18117 ( .A1(n14668), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n14549) );
  NAND2_X1 U18118 ( .A1(n14667), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n14548) );
  AND3_X1 U18119 ( .A1(n14647), .A2(n14549), .A3(n14548), .ZN(n14553) );
  AOI22_X1 U18120 ( .A1(n14682), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14680), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14552) );
  AOI22_X1 U18121 ( .A1(n14681), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14679), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14551) );
  AOI22_X1 U18122 ( .A1(n14683), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16854), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14550) );
  NAND4_X1 U18123 ( .A1(n14553), .A2(n14552), .A3(n14551), .A4(n14550), .ZN(
        n14562) );
  AOI22_X1 U18124 ( .A1(n14682), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14681), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14560) );
  NAND2_X1 U18125 ( .A1(n14668), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14555) );
  NAND2_X1 U18126 ( .A1(n16854), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n14554) );
  AND3_X1 U18127 ( .A1(n14555), .A2(n14677), .A3(n14554), .ZN(n14559) );
  AOI22_X1 U18128 ( .A1(n14680), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14679), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14558) );
  AOI22_X1 U18129 ( .A1(n14683), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14667), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14557) );
  NAND4_X1 U18130 ( .A1(n14560), .A2(n14559), .A3(n14558), .A4(n14557), .ZN(
        n14561) );
  NAND2_X1 U18131 ( .A1(n14562), .A2(n14561), .ZN(n16079) );
  INV_X1 U18132 ( .A(n16079), .ZN(n14563) );
  NAND2_X1 U18133 ( .A1(n14564), .A2(n14563), .ZN(n14572) );
  XOR2_X1 U18134 ( .A(n14571), .B(n14572), .Z(n14565) );
  NAND2_X1 U18135 ( .A1(n14565), .A2(n14625), .ZN(n16081) );
  NOR2_X1 U18136 ( .A1(n20688), .A2(n16079), .ZN(n14566) );
  XOR2_X1 U18137 ( .A(n14567), .B(n14566), .Z(n16080) );
  INV_X1 U18138 ( .A(n14571), .ZN(n14568) );
  NAND2_X1 U18139 ( .A1(n20688), .A2(n14568), .ZN(n16082) );
  NOR3_X1 U18140 ( .A1(n16080), .A2(n16079), .A3(n16082), .ZN(n14569) );
  AOI21_X1 U18141 ( .B1(n16094), .B2(n14570), .A(n14569), .ZN(n14604) );
  NOR2_X1 U18142 ( .A1(n14572), .A2(n14571), .ZN(n14587) );
  AOI22_X1 U18143 ( .A1(n14682), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14680), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14578) );
  NAND2_X1 U18144 ( .A1(n14668), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n14574) );
  NAND2_X1 U18145 ( .A1(n16854), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14573) );
  AND3_X1 U18146 ( .A1(n14647), .A2(n14574), .A3(n14573), .ZN(n14577) );
  AOI22_X1 U18147 ( .A1(n14681), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14679), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14576) );
  AOI22_X1 U18148 ( .A1(n14683), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14667), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14575) );
  NAND4_X1 U18149 ( .A1(n14578), .A2(n14577), .A3(n14576), .A4(n14575), .ZN(
        n14586) );
  AOI22_X1 U18150 ( .A1(n14682), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14680), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14584) );
  NAND2_X1 U18151 ( .A1(n14668), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14580) );
  NAND2_X1 U18152 ( .A1(n16854), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n14579) );
  AND3_X1 U18153 ( .A1(n14580), .A2(n14677), .A3(n14579), .ZN(n14583) );
  AOI22_X1 U18154 ( .A1(n14681), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14679), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14582) );
  AOI22_X1 U18155 ( .A1(n14683), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14667), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14581) );
  NAND4_X1 U18156 ( .A1(n14584), .A2(n14583), .A3(n14582), .A4(n14581), .ZN(
        n14585) );
  AND2_X1 U18157 ( .A1(n14586), .A2(n14585), .ZN(n14588) );
  NAND2_X1 U18158 ( .A1(n14587), .A2(n14588), .ZN(n14609) );
  OAI211_X1 U18159 ( .C1(n14587), .C2(n14588), .A(n14625), .B(n14609), .ZN(
        n14603) );
  NAND2_X1 U18160 ( .A1(n20688), .A2(n14588), .ZN(n16074) );
  NAND2_X1 U18161 ( .A1(n14668), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n14590) );
  NAND2_X1 U18162 ( .A1(n16854), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n14589) );
  AND3_X1 U18163 ( .A1(n14647), .A2(n14590), .A3(n14589), .ZN(n14594) );
  AOI22_X1 U18164 ( .A1(n14682), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14680), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14593) );
  AOI22_X1 U18165 ( .A1(n14681), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14679), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14592) );
  AOI22_X1 U18166 ( .A1(n14683), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14667), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14591) );
  NAND4_X1 U18167 ( .A1(n14594), .A2(n14593), .A3(n14592), .A4(n14591), .ZN(
        n14602) );
  AOI22_X1 U18168 ( .A1(n14682), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14680), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14600) );
  NAND2_X1 U18169 ( .A1(n14668), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14596) );
  NAND2_X1 U18170 ( .A1(n16854), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n14595) );
  AND3_X1 U18171 ( .A1(n14596), .A2(n14677), .A3(n14595), .ZN(n14599) );
  AOI22_X1 U18172 ( .A1(n14681), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14679), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14598) );
  AOI22_X1 U18173 ( .A1(n14683), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14667), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14597) );
  NAND4_X1 U18174 ( .A1(n14600), .A2(n14599), .A3(n14598), .A4(n14597), .ZN(
        n14601) );
  NAND2_X1 U18175 ( .A1(n14602), .A2(n14601), .ZN(n16066) );
  XNOR2_X1 U18176 ( .A(n14609), .B(n16066), .ZN(n14606) );
  NOR2_X1 U18177 ( .A1(n14606), .A2(n14605), .ZN(n16068) );
  NAND2_X1 U18178 ( .A1(n16065), .A2(n16068), .ZN(n14607) );
  OAI21_X1 U18179 ( .B1(n16075), .B2(n10539), .A(n14607), .ZN(n14608) );
  OR2_X1 U18180 ( .A1(n14609), .A2(n16066), .ZN(n14624) );
  INV_X1 U18181 ( .A(n14624), .ZN(n14627) );
  NAND2_X1 U18182 ( .A1(n14668), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n14611) );
  NAND2_X1 U18183 ( .A1(n16854), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14610) );
  AND3_X1 U18184 ( .A1(n14647), .A2(n14611), .A3(n14610), .ZN(n14615) );
  AOI22_X1 U18185 ( .A1(n14682), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14680), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14614) );
  AOI22_X1 U18186 ( .A1(n14683), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14679), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14613) );
  AOI22_X1 U18187 ( .A1(n14681), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14667), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14612) );
  NAND4_X1 U18188 ( .A1(n14615), .A2(n14614), .A3(n14613), .A4(n14612), .ZN(
        n14623) );
  AOI22_X1 U18189 ( .A1(n14683), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14681), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14621) );
  NAND2_X1 U18190 ( .A1(n14668), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14617) );
  NAND2_X1 U18191 ( .A1(n16854), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n14616) );
  AND3_X1 U18192 ( .A1(n14617), .A2(n14677), .A3(n14616), .ZN(n14620) );
  AOI22_X1 U18193 ( .A1(n14682), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14679), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14619) );
  INV_X1 U18194 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n21387) );
  AOI22_X1 U18195 ( .A1(n14680), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14667), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14618) );
  NAND4_X1 U18196 ( .A1(n14621), .A2(n14620), .A3(n14619), .A4(n14618), .ZN(
        n14622) );
  NAND2_X1 U18197 ( .A1(n14623), .A2(n14622), .ZN(n14630) );
  INV_X1 U18198 ( .A(n14630), .ZN(n14626) );
  OR2_X1 U18199 ( .A1(n14624), .A2(n14630), .ZN(n14660) );
  NOR2_X1 U18200 ( .A1(n19972), .A2(n14630), .ZN(n16062) );
  NAND2_X1 U18201 ( .A1(n14668), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n14632) );
  NAND2_X1 U18202 ( .A1(n16854), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n14631) );
  AND3_X1 U18203 ( .A1(n14647), .A2(n14632), .A3(n14631), .ZN(n14636) );
  AOI22_X1 U18204 ( .A1(n14682), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14680), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14635) );
  AOI22_X1 U18205 ( .A1(n14681), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14679), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14634) );
  AOI22_X1 U18206 ( .A1(n14683), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14667), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14633) );
  NAND4_X1 U18207 ( .A1(n14636), .A2(n14635), .A3(n14634), .A4(n14633), .ZN(
        n14644) );
  AOI22_X1 U18208 ( .A1(n14682), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14680), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14642) );
  NAND2_X1 U18209 ( .A1(n14668), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n14638) );
  NAND2_X1 U18210 ( .A1(n16854), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n14637) );
  AND3_X1 U18211 ( .A1(n14638), .A2(n14677), .A3(n14637), .ZN(n14641) );
  AOI22_X1 U18212 ( .A1(n14681), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14679), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14640) );
  AOI22_X1 U18213 ( .A1(n14683), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14667), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14639) );
  NAND4_X1 U18214 ( .A1(n14642), .A2(n14641), .A3(n14640), .A4(n14639), .ZN(
        n14643) );
  NAND2_X1 U18215 ( .A1(n14644), .A2(n14643), .ZN(n16056) );
  NAND2_X1 U18216 ( .A1(n14668), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n14646) );
  NAND2_X1 U18217 ( .A1(n16854), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n14645) );
  AND3_X1 U18218 ( .A1(n14647), .A2(n14646), .A3(n14645), .ZN(n14651) );
  AOI22_X1 U18219 ( .A1(n14682), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14680), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14650) );
  AOI22_X1 U18220 ( .A1(n14683), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14679), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14649) );
  AOI22_X1 U18221 ( .A1(n14681), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14667), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14648) );
  NAND4_X1 U18222 ( .A1(n14651), .A2(n14650), .A3(n14649), .A4(n14648), .ZN(
        n14659) );
  AOI22_X1 U18223 ( .A1(n14681), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14680), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14657) );
  NAND2_X1 U18224 ( .A1(n14668), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n14653) );
  NAND2_X1 U18225 ( .A1(n16854), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n14652) );
  AND3_X1 U18226 ( .A1(n14653), .A2(n14677), .A3(n14652), .ZN(n14656) );
  AOI22_X1 U18227 ( .A1(n14682), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14679), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14655) );
  AOI22_X1 U18228 ( .A1(n14683), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14667), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14654) );
  NAND4_X1 U18229 ( .A1(n14657), .A2(n14656), .A3(n14655), .A4(n14654), .ZN(
        n14658) );
  NAND2_X1 U18230 ( .A1(n14659), .A2(n14658), .ZN(n14664) );
  INV_X1 U18231 ( .A(n14660), .ZN(n16054) );
  INV_X1 U18232 ( .A(n16056), .ZN(n14661) );
  AND2_X1 U18233 ( .A1(n19972), .A2(n14661), .ZN(n14662) );
  NAND2_X1 U18234 ( .A1(n16054), .A2(n14662), .ZN(n14663) );
  NOR2_X1 U18235 ( .A1(n14663), .A2(n14664), .ZN(n14665) );
  AOI21_X1 U18236 ( .B1(n14664), .B2(n14663), .A(n14665), .ZN(n16049) );
  NAND2_X1 U18237 ( .A1(n16050), .A2(n16049), .ZN(n16051) );
  INV_X1 U18238 ( .A(n14665), .ZN(n14666) );
  NAND2_X1 U18239 ( .A1(n16051), .A2(n14666), .ZN(n14693) );
  AOI22_X1 U18240 ( .A1(n14683), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14667), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14671) );
  NAND2_X1 U18241 ( .A1(n16854), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n14670) );
  NAND2_X1 U18242 ( .A1(n14668), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14669) );
  NAND4_X1 U18243 ( .A1(n14671), .A2(n14677), .A3(n14670), .A4(n14669), .ZN(
        n14690) );
  AOI22_X1 U18244 ( .A1(n14682), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14681), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14673) );
  AOI22_X1 U18245 ( .A1(n14680), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14679), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14672) );
  NAND2_X1 U18246 ( .A1(n14673), .A2(n14672), .ZN(n14689) );
  INV_X1 U18247 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14674) );
  NOR2_X1 U18248 ( .A1(n14675), .A2(n14674), .ZN(n14676) );
  AOI211_X1 U18249 ( .C1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .C2(n14678), .A(
        n14677), .B(n14676), .ZN(n14687) );
  AOI22_X1 U18250 ( .A1(n14680), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14679), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14686) );
  AOI22_X1 U18251 ( .A1(n14682), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14681), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14685) );
  AOI22_X1 U18252 ( .A1(n14683), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16854), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14684) );
  NAND4_X1 U18253 ( .A1(n14687), .A2(n14686), .A3(n14685), .A4(n14684), .ZN(
        n14688) );
  OAI21_X1 U18254 ( .B1(n14690), .B2(n14689), .A(n14688), .ZN(n14691) );
  INV_X1 U18255 ( .A(n14691), .ZN(n14692) );
  XNOR2_X1 U18256 ( .A(n14693), .B(n14692), .ZN(n14704) );
  NAND2_X1 U18257 ( .A1(n14694), .A2(n16872), .ZN(n16264) );
  INV_X1 U18258 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n14696) );
  AOI22_X1 U18259 ( .A1(n16260), .A2(n19934), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n19887), .ZN(n14695) );
  OAI21_X1 U18260 ( .B1(n16264), .B2(n14696), .A(n14695), .ZN(n14699) );
  NOR2_X1 U18261 ( .A1(n14697), .A2(n16282), .ZN(n14698) );
  OAI21_X1 U18262 ( .B1(n14704), .B2(n16227), .A(n14700), .ZN(P2_U2889) );
  NOR2_X1 U18263 ( .A1(n14701), .A2(n16154), .ZN(n14702) );
  AOI21_X1 U18264 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n16154), .A(n14702), .ZN(
        n14703) );
  OAI21_X1 U18265 ( .B1(n14704), .B2(n9716), .A(n14703), .ZN(P2_U2857) );
  INV_X1 U18266 ( .A(n14705), .ZN(n14707) );
  AND2_X1 U18267 ( .A1(n14707), .A2(n14706), .ZN(n14711) );
  INV_X1 U18268 ( .A(n14709), .ZN(n16398) );
  INV_X1 U18269 ( .A(n16668), .ZN(n16409) );
  OR2_X1 U18270 ( .A1(n19961), .A2(n16409), .ZN(n14713) );
  NAND2_X1 U18271 ( .A1(n16740), .A2(n14713), .ZN(n16672) );
  NOR2_X1 U18272 ( .A1(n14714), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14715) );
  NOR2_X1 U18273 ( .A1(n16672), .A2(n14715), .ZN(n14716) );
  OAI21_X1 U18274 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n19961), .A(
        n16664), .ZN(n14730) );
  AOI21_X1 U18275 ( .B1(n14721), .B2(n14717), .A(n14719), .ZN(n14735) );
  INV_X1 U18276 ( .A(n14735), .ZN(n16123) );
  NAND2_X1 U18277 ( .A1(n16738), .A2(n14722), .ZN(n14723) );
  INV_X1 U18278 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14724) );
  AOI21_X1 U18279 ( .B1(n14727), .B2(n14725), .A(n14726), .ZN(n16248) );
  NOR2_X1 U18280 ( .A1(n16491), .A2(n20593), .ZN(n14732) );
  AOI21_X1 U18281 ( .B1(n16248), .B2(n19956), .A(n14732), .ZN(n14728) );
  OAI21_X1 U18282 ( .B1(n14739), .B2(n16802), .A(n14731), .ZN(P2_U3029) );
  AOI21_X1 U18283 ( .B1(n16510), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n14732), .ZN(n14733) );
  OAI21_X1 U18284 ( .B1(n16544), .B2(n15910), .A(n14733), .ZN(n14734) );
  AOI21_X1 U18285 ( .B1(n14735), .B2(n16547), .A(n14734), .ZN(n14738) );
  OAI211_X1 U18286 ( .C1(n14736), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n19945), .B(n16394), .ZN(n14737) );
  OAI211_X1 U18287 ( .C1(n14739), .C2(n16483), .A(n14738), .B(n14737), .ZN(
        P2_U2997) );
  INV_X1 U18288 ( .A(n16264), .ZN(n16203) );
  AOI22_X1 U18289 ( .A1(n16203), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19887), .ZN(n14741) );
  NAND2_X1 U18290 ( .A1(n16259), .A2(BUF1_REG_31__SCAN_IN), .ZN(n14740) );
  OAI211_X1 U18291 ( .C1(n12600), .C2(n16282), .A(n14741), .B(n14740), .ZN(
        P2_U2888) );
  NAND2_X1 U18292 ( .A1(n19943), .A2(n14742), .ZN(n14745) );
  AOI21_X1 U18293 ( .B1(n16510), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14743), .ZN(n14744) );
  AND2_X1 U18294 ( .A1(n14745), .A2(n14744), .ZN(n14746) );
  OAI21_X1 U18295 ( .B1(n14747), .B2(n19950), .A(n14746), .ZN(n14748) );
  NAND2_X1 U18296 ( .A1(n16157), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14751) );
  OAI21_X1 U18297 ( .B1(n14747), .B2(n16157), .A(n14751), .ZN(P2_U2856) );
  NAND2_X1 U18298 ( .A1(n21029), .A2(n17222), .ZN(n20706) );
  NAND2_X1 U18299 ( .A1(n14752), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n14753)
         );
  NAND3_X1 U18300 ( .A1(n14754), .A2(n20706), .A3(n14753), .ZN(P1_U2801) );
  INV_X1 U18301 ( .A(n14755), .ZN(n14759) );
  INV_X1 U18302 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n14756) );
  NAND2_X1 U18303 ( .A1(n20706), .A2(n14756), .ZN(n14758) );
  MUX2_X1 U18304 ( .A(n14759), .B(n14758), .S(n14757), .Z(P1_U3487) );
  AOI21_X1 U18305 ( .B1(n14761), .B2(n14771), .A(n14760), .ZN(n15176) );
  INV_X1 U18306 ( .A(n15176), .ZN(n15084) );
  AOI21_X1 U18307 ( .B1(n14763), .B2(n14774), .A(n14762), .ZN(n15405) );
  AOI22_X1 U18308 ( .A1(n20757), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20785), .ZN(n14764) );
  OAI21_X1 U18309 ( .B1(n15023), .B2(n15174), .A(n14764), .ZN(n14768) );
  NOR2_X1 U18310 ( .A1(n14793), .A2(n14765), .ZN(n14766) );
  MUX2_X1 U18311 ( .A(n14766), .B(n14779), .S(P1_REIP_REG_29__SCAN_IN), .Z(
        n14767) );
  OAI21_X1 U18312 ( .B1(n15084), .B2(n20749), .A(n14769), .ZN(P1_U2811) );
  INV_X1 U18313 ( .A(n14774), .ZN(n14775) );
  AOI21_X1 U18314 ( .B1(n14776), .B2(n14773), .A(n14775), .ZN(n15415) );
  INV_X1 U18315 ( .A(n15187), .ZN(n14778) );
  AOI22_X1 U18316 ( .A1(n20757), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20785), .ZN(n14777) );
  OAI21_X1 U18317 ( .B1(n15023), .B2(n14778), .A(n14777), .ZN(n14782) );
  INV_X1 U18318 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21267) );
  NOR2_X1 U18319 ( .A1(n14793), .A2(n21267), .ZN(n14780) );
  MUX2_X1 U18320 ( .A(n14780), .B(n14779), .S(P1_REIP_REG_28__SCAN_IN), .Z(
        n14781) );
  OAI21_X1 U18321 ( .B1(n15185), .B2(n20749), .A(n14783), .ZN(P1_U2812) );
  AOI21_X1 U18322 ( .B1(n14785), .B2(n14784), .A(n14770), .ZN(n15194) );
  INV_X1 U18323 ( .A(n15194), .ZN(n15093) );
  INV_X1 U18324 ( .A(n14787), .ZN(n14797) );
  NAND2_X1 U18325 ( .A1(n14786), .A2(n14797), .ZN(n14789) );
  INV_X1 U18326 ( .A(n14773), .ZN(n14788) );
  AOI22_X1 U18327 ( .A1(n20757), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20785), .ZN(n14791) );
  OAI21_X1 U18328 ( .B1(n15023), .B2(n15192), .A(n14791), .ZN(n14792) );
  AOI21_X1 U18329 ( .B1(n15424), .B2(n9580), .A(n14792), .ZN(n14795) );
  MUX2_X1 U18330 ( .A(n14793), .B(n14800), .S(P1_REIP_REG_27__SCAN_IN), .Z(
        n14794) );
  OAI211_X1 U18331 ( .C1(n15093), .C2(n20749), .A(n14795), .B(n14794), .ZN(
        P1_U2813) );
  XOR2_X1 U18332 ( .A(n14796), .B(n9606), .Z(n15203) );
  INV_X1 U18333 ( .A(n15203), .ZN(n15097) );
  OAI22_X1 U18334 ( .A1(n20781), .A2(n15050), .B1(n15201), .B2(n20762), .ZN(
        n14799) );
  XNOR2_X1 U18335 ( .A(n14786), .B(n14797), .ZN(n15427) );
  NOR2_X1 U18336 ( .A1(n15427), .A2(n20780), .ZN(n14798) );
  AOI211_X1 U18337 ( .C1(n17157), .C2(n15199), .A(n14799), .B(n14798), .ZN(
        n14803) );
  NAND3_X1 U18338 ( .A1(n14824), .A2(P1_REIP_REG_25__SCAN_IN), .A3(
        P1_REIP_REG_24__SCAN_IN), .ZN(n14801) );
  MUX2_X1 U18339 ( .A(n14801), .B(n14800), .S(P1_REIP_REG_26__SCAN_IN), .Z(
        n14802) );
  OAI211_X1 U18340 ( .C1(n15097), .C2(n20749), .A(n14803), .B(n14802), .ZN(
        P1_U2814) );
  AOI21_X1 U18341 ( .B1(n14805), .B2(n14804), .A(n9606), .ZN(n15216) );
  INV_X1 U18342 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n15212) );
  XOR2_X1 U18343 ( .A(P1_REIP_REG_25__SCAN_IN), .B(P1_REIP_REG_24__SCAN_IN), 
        .Z(n14806) );
  NAND2_X1 U18344 ( .A1(n14824), .A2(n14806), .ZN(n14812) );
  NOR2_X1 U18345 ( .A1(n9640), .A2(n14807), .ZN(n14808) );
  OR2_X1 U18346 ( .A1(n14786), .A2(n14808), .ZN(n15051) );
  INV_X1 U18347 ( .A(n15051), .ZN(n15443) );
  AOI22_X1 U18348 ( .A1(n20757), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20785), .ZN(n14809) );
  OAI21_X1 U18349 ( .B1(n12914), .B2(n15214), .A(n14809), .ZN(n14810) );
  AOI21_X1 U18350 ( .B1(n15443), .B2(n20758), .A(n14810), .ZN(n14811) );
  OAI211_X1 U18351 ( .C1(n14835), .C2(n15212), .A(n14812), .B(n14811), .ZN(
        n14813) );
  AOI21_X1 U18352 ( .B1(n15216), .B2(n12954), .A(n14813), .ZN(n14814) );
  INV_X1 U18353 ( .A(n14814), .ZN(P1_U2815) );
  OAI21_X1 U18354 ( .B1(n14815), .B2(n14816), .A(n14804), .ZN(n15222) );
  INV_X1 U18355 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21263) );
  AND2_X1 U18356 ( .A1(n14831), .A2(n14817), .ZN(n14818) );
  NOR2_X1 U18357 ( .A1(n9640), .A2(n14818), .ZN(n15455) );
  NAND2_X1 U18358 ( .A1(n15455), .A2(n20758), .ZN(n14822) );
  OR2_X1 U18359 ( .A1(n14835), .A2(n21263), .ZN(n14821) );
  AOI22_X1 U18360 ( .A1(n20757), .A2(P1_EBX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20785), .ZN(n14820) );
  NAND2_X1 U18361 ( .A1(n17157), .A2(n15225), .ZN(n14819) );
  NAND4_X1 U18362 ( .A1(n14822), .A2(n14821), .A3(n14820), .A4(n14819), .ZN(
        n14823) );
  AOI21_X1 U18363 ( .B1(n14824), .B2(n21263), .A(n14823), .ZN(n14825) );
  OAI21_X1 U18364 ( .B1(n15222), .B2(n20749), .A(n14825), .ZN(P1_U2816) );
  AOI21_X1 U18365 ( .B1(n14827), .B2(n14826), .A(n14815), .ZN(n15232) );
  INV_X1 U18366 ( .A(n15232), .ZN(n15111) );
  NAND2_X1 U18367 ( .A1(n14828), .A2(n14829), .ZN(n14830) );
  NAND2_X1 U18368 ( .A1(n14831), .A2(n14830), .ZN(n15054) );
  INV_X1 U18369 ( .A(n15054), .ZN(n15463) );
  AOI22_X1 U18370 ( .A1(n20757), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20785), .ZN(n14832) );
  OAI21_X1 U18371 ( .B1(n15023), .B2(n15230), .A(n14832), .ZN(n14833) );
  AOI21_X1 U18372 ( .B1(n15463), .B2(n9580), .A(n14833), .ZN(n14839) );
  NAND2_X1 U18373 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n14834) );
  NOR2_X1 U18374 ( .A1(n14860), .A2(n14834), .ZN(n14837) );
  INV_X1 U18375 ( .A(n14835), .ZN(n14836) );
  OAI21_X1 U18376 ( .B1(n14837), .B2(P1_REIP_REG_23__SCAN_IN), .A(n14836), 
        .ZN(n14838) );
  OAI211_X1 U18377 ( .C1(n15111), .C2(n20749), .A(n14839), .B(n14838), .ZN(
        P1_U2817) );
  XNOR2_X1 U18378 ( .A(n14840), .B(n14841), .ZN(n15243) );
  AND2_X1 U18379 ( .A1(n14842), .A2(n20729), .ZN(n14863) );
  OAI21_X1 U18380 ( .B1(n14853), .B2(n14843), .A(n14828), .ZN(n15473) );
  AOI22_X1 U18381 ( .A1(n20757), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20785), .ZN(n14845) );
  NAND2_X1 U18382 ( .A1(n17157), .A2(n15236), .ZN(n14844) );
  OAI211_X1 U18383 ( .C1(n15473), .C2(n20780), .A(n14845), .B(n14844), .ZN(
        n14848) );
  XNOR2_X1 U18384 ( .A(P1_REIP_REG_22__SCAN_IN), .B(P1_REIP_REG_21__SCAN_IN), 
        .ZN(n14846) );
  NOR2_X1 U18385 ( .A1(n14860), .A2(n14846), .ZN(n14847) );
  AOI211_X1 U18386 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(n14863), .A(n14848), 
        .B(n14847), .ZN(n14849) );
  OAI21_X1 U18387 ( .B1(n20749), .B2(n15243), .A(n14849), .ZN(P1_U2818) );
  AOI21_X1 U18388 ( .B1(n14851), .B2(n14850), .A(n14840), .ZN(n15251) );
  NAND2_X1 U18389 ( .A1(n15251), .A2(n12954), .ZN(n14859) );
  AOI22_X1 U18390 ( .A1(n20757), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20785), .ZN(n14852) );
  OAI21_X1 U18391 ( .B1(n15023), .B2(n15249), .A(n14852), .ZN(n14857) );
  INV_X1 U18392 ( .A(n14853), .ZN(n14854) );
  OAI21_X1 U18393 ( .B1(n14855), .B2(n14868), .A(n14854), .ZN(n15478) );
  NOR2_X1 U18394 ( .A1(n15478), .A2(n20780), .ZN(n14856) );
  AOI211_X1 U18395 ( .C1(n14863), .C2(P1_REIP_REG_21__SCAN_IN), .A(n14857), 
        .B(n14856), .ZN(n14858) );
  OAI211_X1 U18396 ( .C1(P1_REIP_REG_21__SCAN_IN), .C2(n14860), .A(n14859), 
        .B(n14858), .ZN(P1_U2819) );
  OAI21_X1 U18397 ( .B1(n14861), .B2(n14862), .A(n14850), .ZN(n15262) );
  INV_X1 U18398 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n15265) );
  INV_X1 U18399 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21251) );
  NOR3_X1 U18400 ( .A1(n14896), .A2(n15265), .A3(n21251), .ZN(n14864) );
  OAI21_X1 U18401 ( .B1(n14864), .B2(P1_REIP_REG_20__SCAN_IN), .A(n14863), 
        .ZN(n14872) );
  OAI22_X1 U18402 ( .A1(n20781), .A2(n15057), .B1(n15257), .B2(n20762), .ZN(
        n14870) );
  NOR2_X1 U18403 ( .A1(n14865), .A2(n14866), .ZN(n14867) );
  OR2_X1 U18404 ( .A1(n14868), .A2(n14867), .ZN(n15489) );
  NOR2_X1 U18405 ( .A1(n15489), .A2(n20780), .ZN(n14869) );
  AOI211_X1 U18406 ( .C1(n17157), .C2(n15259), .A(n14870), .B(n14869), .ZN(
        n14871) );
  OAI211_X1 U18407 ( .C1(n15262), .C2(n20749), .A(n14872), .B(n14871), .ZN(
        P1_U2820) );
  XNOR2_X1 U18408 ( .A(P1_REIP_REG_19__SCAN_IN), .B(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14888) );
  INV_X1 U18409 ( .A(n14930), .ZN(n14874) );
  NAND2_X1 U18410 ( .A1(n14928), .A2(n14916), .ZN(n14915) );
  INV_X1 U18411 ( .A(n14875), .ZN(n14889) );
  AOI21_X1 U18412 ( .B1(n14901), .B2(n14889), .A(n14876), .ZN(n14877) );
  NOR2_X1 U18413 ( .A1(n14877), .A2(n14861), .ZN(n15269) );
  NAND2_X1 U18414 ( .A1(n15269), .A2(n12954), .ZN(n14887) );
  AOI21_X1 U18415 ( .B1(n14878), .B2(n14892), .A(n14865), .ZN(n15495) );
  AOI21_X1 U18416 ( .B1(n20785), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n20772), .ZN(n14880) );
  NAND2_X1 U18417 ( .A1(n20757), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n14879) );
  OAI211_X1 U18418 ( .C1(n12914), .C2(n15267), .A(n14880), .B(n14879), .ZN(
        n14885) );
  INV_X1 U18419 ( .A(n14881), .ZN(n14883) );
  OAI21_X1 U18420 ( .B1(n14883), .B2(n14882), .A(n20729), .ZN(n14913) );
  NOR2_X1 U18421 ( .A1(n14913), .A2(n15265), .ZN(n14884) );
  AOI211_X1 U18422 ( .C1(n15495), .C2(n9580), .A(n14885), .B(n14884), .ZN(
        n14886) );
  OAI211_X1 U18423 ( .C1(n14896), .C2(n14888), .A(n14887), .B(n14886), .ZN(
        P1_U2821) );
  XNOR2_X1 U18424 ( .A(n14901), .B(n14889), .ZN(n15278) );
  INV_X1 U18425 ( .A(n14913), .ZN(n14899) );
  NAND2_X1 U18426 ( .A1(n14906), .A2(n14890), .ZN(n14891) );
  NAND2_X1 U18427 ( .A1(n14892), .A2(n14891), .ZN(n15498) );
  AOI21_X1 U18428 ( .B1(n20785), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20772), .ZN(n14893) );
  OAI21_X1 U18429 ( .B1(n20781), .B2(n15059), .A(n14893), .ZN(n14894) );
  AOI21_X1 U18430 ( .B1(n17157), .B2(n15276), .A(n14894), .ZN(n14895) );
  OAI21_X1 U18431 ( .B1(n15498), .B2(n20780), .A(n14895), .ZN(n14898) );
  NOR2_X1 U18432 ( .A1(n14896), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14897) );
  AOI211_X1 U18433 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n14899), .A(n14898), 
        .B(n14897), .ZN(n14900) );
  OAI21_X1 U18434 ( .B1(n20749), .B2(n15278), .A(n14900), .ZN(P1_U2822) );
  AOI21_X1 U18435 ( .B1(n14925), .B2(P1_REIP_REG_16__SCAN_IN), .A(
        P1_REIP_REG_17__SCAN_IN), .ZN(n14914) );
  AOI21_X1 U18436 ( .B1(n14902), .B2(n14915), .A(n14901), .ZN(n15293) );
  NAND2_X1 U18437 ( .A1(n15293), .A2(n12954), .ZN(n14912) );
  NAND2_X1 U18438 ( .A1(n14903), .A2(n14904), .ZN(n14905) );
  AND2_X1 U18439 ( .A1(n14906), .A2(n14905), .ZN(n15517) );
  OAI21_X1 U18440 ( .B1(n20762), .B2(n14907), .A(n20759), .ZN(n14908) );
  AOI21_X1 U18441 ( .B1(n20757), .B2(P1_EBX_REG_17__SCAN_IN), .A(n14908), .ZN(
        n14909) );
  OAI21_X1 U18442 ( .B1(n15023), .B2(n15291), .A(n14909), .ZN(n14910) );
  AOI21_X1 U18443 ( .B1(n15517), .B2(n9580), .A(n14910), .ZN(n14911) );
  OAI211_X1 U18444 ( .C1(n14914), .C2(n14913), .A(n14912), .B(n14911), .ZN(
        P1_U2823) );
  OAI21_X1 U18445 ( .B1(n14928), .B2(n14916), .A(n14915), .ZN(n15307) );
  INV_X1 U18446 ( .A(n15001), .ZN(n14983) );
  NOR3_X1 U18447 ( .A1(n14983), .A2(P1_REIP_REG_15__SCAN_IN), .A3(n14917), 
        .ZN(n14936) );
  AND2_X1 U18448 ( .A1(n14918), .A2(n20729), .ZN(n14944) );
  OAI21_X1 U18449 ( .B1(n14936), .B2(n14944), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n14927) );
  INV_X1 U18450 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21249) );
  OAI21_X1 U18451 ( .B1(n14919), .B2(n14920), .A(n14903), .ZN(n15529) );
  AOI21_X1 U18452 ( .B1(n20785), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20772), .ZN(n14921) );
  OAI21_X1 U18453 ( .B1(n20781), .B2(n15061), .A(n14921), .ZN(n14922) );
  AOI21_X1 U18454 ( .B1(n17157), .B2(n15303), .A(n14922), .ZN(n14923) );
  OAI21_X1 U18455 ( .B1(n20780), .B2(n15529), .A(n14923), .ZN(n14924) );
  AOI21_X1 U18456 ( .B1(n14925), .B2(n21249), .A(n14924), .ZN(n14926) );
  OAI211_X1 U18457 ( .C1(n15307), .C2(n20749), .A(n14927), .B(n14926), .ZN(
        P1_U2824) );
  INV_X1 U18458 ( .A(n14928), .ZN(n14929) );
  OAI21_X1 U18459 ( .B1(n20762), .B2(n21369), .A(n20759), .ZN(n14934) );
  INV_X1 U18460 ( .A(n14919), .ZN(n14931) );
  OAI21_X1 U18461 ( .B1(n14932), .B2(n14946), .A(n14931), .ZN(n15538) );
  NOR2_X1 U18462 ( .A1(n15538), .A2(n20780), .ZN(n14933) );
  AOI211_X1 U18463 ( .C1(P1_EBX_REG_15__SCAN_IN), .C2(n20757), .A(n14934), .B(
        n14933), .ZN(n14935) );
  OAI21_X1 U18464 ( .B1(n15315), .B2(n15023), .A(n14935), .ZN(n14937) );
  AOI211_X1 U18465 ( .C1(n14944), .C2(P1_REIP_REG_15__SCAN_IN), .A(n14937), 
        .B(n14936), .ZN(n14938) );
  OAI21_X1 U18466 ( .B1(n20749), .B2(n15319), .A(n14938), .ZN(P1_U2825) );
  NAND2_X1 U18467 ( .A1(n14939), .A2(n14940), .ZN(n14941) );
  AND2_X1 U18468 ( .A1(n14942), .A2(n14941), .ZN(n15328) );
  NOR2_X1 U18469 ( .A1(n14983), .A2(n14943), .ZN(n14945) );
  OAI21_X1 U18470 ( .B1(n14945), .B2(P1_REIP_REG_14__SCAN_IN), .A(n14944), 
        .ZN(n14952) );
  AOI21_X1 U18471 ( .B1(n14947), .B2(n14960), .A(n14946), .ZN(n15546) );
  AOI21_X1 U18472 ( .B1(n20785), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20772), .ZN(n14948) );
  OAI21_X1 U18473 ( .B1(n20781), .B2(n21352), .A(n14948), .ZN(n14950) );
  NOR2_X1 U18474 ( .A1(n15023), .A2(n15326), .ZN(n14949) );
  AOI211_X1 U18475 ( .C1(n15546), .C2(n9580), .A(n14950), .B(n14949), .ZN(
        n14951) );
  OAI211_X1 U18476 ( .C1(n15153), .C2(n20749), .A(n14952), .B(n14951), .ZN(
        P1_U2826) );
  XOR2_X1 U18477 ( .A(n14954), .B(n14279), .Z(n14990) );
  INV_X1 U18478 ( .A(n14953), .ZN(n14989) );
  INV_X1 U18479 ( .A(n14954), .ZN(n14955) );
  NOR2_X1 U18480 ( .A1(n14279), .A2(n14955), .ZN(n14973) );
  OAI21_X1 U18481 ( .B1(n14988), .B2(n14973), .A(n14972), .ZN(n14971) );
  INV_X1 U18482 ( .A(n14939), .ZN(n14956) );
  AOI21_X1 U18483 ( .B1(n14971), .B2(n14957), .A(n14956), .ZN(n15338) );
  INV_X1 U18484 ( .A(n15338), .ZN(n15157) );
  NAND2_X1 U18485 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14967) );
  INV_X1 U18486 ( .A(n14967), .ZN(n14958) );
  AOI21_X1 U18487 ( .B1(n14991), .B2(n14958), .A(n20755), .ZN(n14984) );
  INV_X1 U18488 ( .A(n14960), .ZN(n14961) );
  AOI21_X1 U18489 ( .B1(n14962), .B2(n14959), .A(n14961), .ZN(n15555) );
  NAND2_X1 U18490 ( .A1(n20757), .A2(P1_EBX_REG_13__SCAN_IN), .ZN(n14963) );
  OAI211_X1 U18491 ( .C1(n20762), .C2(n14964), .A(n14963), .B(n20759), .ZN(
        n14965) );
  AOI21_X1 U18492 ( .B1(n15555), .B2(n20758), .A(n14965), .ZN(n14966) );
  OAI21_X1 U18493 ( .B1(n15336), .B2(n15023), .A(n14966), .ZN(n14969) );
  NOR3_X1 U18494 ( .A1(n14983), .A2(P1_REIP_REG_13__SCAN_IN), .A3(n14967), 
        .ZN(n14968) );
  AOI211_X1 U18495 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(n14984), .A(n14969), 
        .B(n14968), .ZN(n14970) );
  OAI21_X1 U18496 ( .B1(n15157), .B2(n20749), .A(n14970), .ZN(P1_U2827) );
  INV_X1 U18497 ( .A(n14971), .ZN(n14975) );
  NOR3_X1 U18498 ( .A1(n14988), .A2(n14973), .A3(n14972), .ZN(n14974) );
  NOR2_X1 U18499 ( .A1(n14975), .A2(n14974), .ZN(n15351) );
  INV_X1 U18500 ( .A(n15351), .ZN(n15159) );
  OR2_X1 U18501 ( .A1(n14976), .A2(n14977), .ZN(n14978) );
  AND2_X1 U18502 ( .A1(n14959), .A2(n14978), .ZN(n15569) );
  NAND2_X1 U18503 ( .A1(n20757), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n14979) );
  OAI211_X1 U18504 ( .C1(n20762), .C2(n14980), .A(n14979), .B(n20759), .ZN(
        n14982) );
  NOR2_X1 U18505 ( .A1(n15023), .A2(n15349), .ZN(n14981) );
  AOI211_X1 U18506 ( .C1(n15569), .C2(n9580), .A(n14982), .B(n14981), .ZN(
        n14987) );
  INV_X1 U18507 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15357) );
  NOR2_X1 U18508 ( .A1(n14983), .A2(n15357), .ZN(n14985) );
  OAI21_X1 U18509 ( .B1(n14985), .B2(P1_REIP_REG_12__SCAN_IN), .A(n14984), 
        .ZN(n14986) );
  OAI211_X1 U18510 ( .C1(n15159), .C2(n20749), .A(n14987), .B(n14986), .ZN(
        P1_U2828) );
  AOI21_X1 U18511 ( .B1(n14990), .B2(n14989), .A(n14988), .ZN(n15361) );
  INV_X1 U18512 ( .A(n15361), .ZN(n15164) );
  INV_X1 U18513 ( .A(n14991), .ZN(n14992) );
  NAND2_X1 U18514 ( .A1(n14992), .A2(n20729), .ZN(n17153) );
  NOR2_X1 U18515 ( .A1(n14994), .A2(n14993), .ZN(n14995) );
  OR2_X1 U18516 ( .A1(n14976), .A2(n14995), .ZN(n15572) );
  INV_X1 U18517 ( .A(n15572), .ZN(n14996) );
  AOI22_X1 U18518 ( .A1(n14996), .A2(n20758), .B1(n20757), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n14997) );
  OAI21_X1 U18519 ( .B1(n15357), .B2(n17153), .A(n14997), .ZN(n14998) );
  AOI211_X1 U18520 ( .C1(n20785), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n14998), .B(n20772), .ZN(n14999) );
  OAI21_X1 U18521 ( .B1(n15023), .B2(n15359), .A(n14999), .ZN(n15000) );
  AOI21_X1 U18522 ( .B1(n15001), .B2(n15357), .A(n15000), .ZN(n15002) );
  OAI21_X1 U18523 ( .B1(n15164), .B2(n20749), .A(n15002), .ZN(P1_U2829) );
  INV_X1 U18524 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21237) );
  NOR3_X1 U18525 ( .A1(n15009), .A2(n20755), .A3(n21237), .ZN(n15007) );
  OAI21_X1 U18526 ( .B1(n20762), .B2(n12013), .A(n20759), .ZN(n15003) );
  AOI21_X1 U18527 ( .B1(n20757), .B2(P1_EBX_REG_9__SCAN_IN), .A(n15003), .ZN(
        n15005) );
  NAND2_X1 U18528 ( .A1(n20758), .A2(n17185), .ZN(n15004) );
  OAI211_X1 U18529 ( .C1(n12914), .C2(n15377), .A(n15005), .B(n15004), .ZN(
        n15006) );
  AOI211_X1 U18530 ( .C1(n17160), .C2(n21237), .A(n15007), .B(n15006), .ZN(
        n15008) );
  OAI21_X1 U18531 ( .B1(n20749), .B2(n15381), .A(n15008), .ZN(P1_U2831) );
  INV_X1 U18532 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21233) );
  INV_X1 U18533 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21234) );
  OAI21_X1 U18534 ( .B1(n20735), .B2(n21233), .A(n21234), .ZN(n15016) );
  NOR2_X1 U18535 ( .A1(n15009), .A2(n20755), .ZN(n15015) );
  OAI21_X1 U18536 ( .B1(n20762), .B2(n15010), .A(n20759), .ZN(n15011) );
  AOI21_X1 U18537 ( .B1(n20757), .B2(P1_EBX_REG_8__SCAN_IN), .A(n15011), .ZN(
        n15013) );
  NAND2_X1 U18538 ( .A1(n20758), .A2(n15605), .ZN(n15012) );
  OAI211_X1 U18539 ( .C1(n12914), .C2(n15387), .A(n15013), .B(n15012), .ZN(
        n15014) );
  AOI21_X1 U18540 ( .B1(n15016), .B2(n15015), .A(n15014), .ZN(n15017) );
  OAI21_X1 U18541 ( .B1(n20749), .B2(n15018), .A(n15017), .ZN(P1_U2832) );
  NAND2_X1 U18542 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n15019) );
  AOI21_X1 U18543 ( .B1(n20783), .B2(n15019), .A(n20784), .ZN(n15036) );
  INV_X1 U18544 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n21225) );
  NOR2_X1 U18545 ( .A1(n15026), .A2(n15020), .ZN(n20786) );
  AOI22_X1 U18546 ( .A1(n20757), .A2(P1_EBX_REG_3__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n20785), .ZN(n15022) );
  NAND4_X1 U18547 ( .A1(n20783), .A2(n21225), .A3(P1_REIP_REG_2__SCAN_IN), 
        .A4(P1_REIP_REG_1__SCAN_IN), .ZN(n15021) );
  OAI211_X1 U18548 ( .C1(n20780), .C2(n20901), .A(n15022), .B(n15021), .ZN(
        n15025) );
  NOR2_X1 U18549 ( .A1(n15023), .A2(n20872), .ZN(n15024) );
  AOI211_X1 U18550 ( .C1(n20786), .C2(n15657), .A(n15025), .B(n15024), .ZN(
        n15029) );
  OAI21_X1 U18551 ( .B1(n15027), .B2(n15026), .A(n20749), .ZN(n20792) );
  NAND2_X1 U18552 ( .A1(n20869), .A2(n20792), .ZN(n15028) );
  OAI211_X1 U18553 ( .C1(n15036), .C2(n21225), .A(n15029), .B(n15028), .ZN(
        P1_U2837) );
  AOI21_X1 U18554 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20783), .A(
        P1_REIP_REG_2__SCAN_IN), .ZN(n15035) );
  AOI22_X1 U18555 ( .A1(n20757), .A2(P1_EBX_REG_2__SCAN_IN), .B1(n20785), .B2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n15032) );
  AOI22_X1 U18556 ( .A1(n15030), .A2(n20786), .B1(n20758), .B2(n20917), .ZN(
        n15031) );
  OAI211_X1 U18557 ( .C1(n12914), .C2(n20880), .A(n15032), .B(n15031), .ZN(
        n15033) );
  AOI21_X1 U18558 ( .B1(n20877), .B2(n20792), .A(n15033), .ZN(n15034) );
  OAI21_X1 U18559 ( .B1(n15036), .B2(n15035), .A(n15034), .ZN(P1_U2838) );
  INV_X1 U18560 ( .A(n20792), .ZN(n15042) );
  AOI22_X1 U18561 ( .A1(n20786), .A2(n15641), .B1(n20757), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n15037) );
  OAI21_X1 U18562 ( .B1(n20780), .B2(n20928), .A(n15037), .ZN(n15038) );
  AOI21_X1 U18563 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(n20729), .A(n15038), .ZN(
        n15040) );
  OAI21_X1 U18564 ( .B1(n17157), .B2(n20785), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15039) );
  OAI211_X1 U18565 ( .C1(n15042), .C2(n15041), .A(n15040), .B(n15039), .ZN(
        P1_U2840) );
  INV_X1 U18566 ( .A(n15043), .ZN(n15045) );
  OAI22_X1 U18567 ( .A1(n15045), .A2(n15068), .B1(n20800), .B2(n15044), .ZN(
        P1_U2841) );
  AOI22_X1 U18568 ( .A1(n15397), .A2(n20795), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n15065), .ZN(n15046) );
  OAI21_X1 U18569 ( .B1(n15077), .B2(n15067), .A(n15046), .ZN(P1_U2842) );
  AOI22_X1 U18570 ( .A1(n15405), .A2(n20795), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n15065), .ZN(n15047) );
  OAI21_X1 U18571 ( .B1(n15084), .B2(n15067), .A(n15047), .ZN(P1_U2843) );
  AOI22_X1 U18572 ( .A1(n15415), .A2(n20795), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n15065), .ZN(n15048) );
  OAI21_X1 U18573 ( .B1(n15185), .B2(n15067), .A(n15048), .ZN(P1_U2844) );
  INV_X1 U18574 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n21349) );
  INV_X1 U18575 ( .A(n15424), .ZN(n15049) );
  OAI222_X1 U18576 ( .A1(n15067), .A2(n15093), .B1(n21349), .B2(n20800), .C1(
        n15049), .C2(n15068), .ZN(P1_U2845) );
  OAI222_X1 U18577 ( .A1(n15097), .A2(n15070), .B1(n15050), .B2(n20800), .C1(
        n15068), .C2(n15427), .ZN(P1_U2846) );
  INV_X1 U18578 ( .A(n15216), .ZN(n15101) );
  INV_X1 U18579 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15052) );
  OAI222_X1 U18580 ( .A1(n15067), .A2(n15101), .B1(n15052), .B2(n20800), .C1(
        n15051), .C2(n15068), .ZN(P1_U2847) );
  AOI22_X1 U18581 ( .A1(n15455), .A2(n20795), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n15065), .ZN(n15053) );
  OAI21_X1 U18582 ( .B1(n15222), .B2(n15067), .A(n15053), .ZN(P1_U2848) );
  INV_X1 U18583 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n21398) );
  OAI222_X1 U18584 ( .A1(n15111), .A2(n15070), .B1(n21398), .B2(n20800), .C1(
        n15054), .C2(n15068), .ZN(P1_U2849) );
  OAI222_X1 U18585 ( .A1(n15243), .A2(n15070), .B1(n15055), .B2(n20800), .C1(
        n15473), .C2(n15068), .ZN(P1_U2850) );
  INV_X1 U18586 ( .A(n15251), .ZN(n15121) );
  INV_X1 U18587 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15056) );
  OAI222_X1 U18588 ( .A1(n15121), .A2(n15070), .B1(n15056), .B2(n20800), .C1(
        n15478), .C2(n15068), .ZN(P1_U2851) );
  OAI222_X1 U18589 ( .A1(n15262), .A2(n15070), .B1(n15057), .B2(n20800), .C1(
        n15489), .C2(n15068), .ZN(P1_U2852) );
  INV_X1 U18590 ( .A(n15269), .ZN(n15130) );
  AOI22_X1 U18591 ( .A1(n15495), .A2(n20795), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n15065), .ZN(n15058) );
  OAI21_X1 U18592 ( .B1(n15130), .B2(n15067), .A(n15058), .ZN(P1_U2853) );
  OAI222_X1 U18593 ( .A1(n15498), .A2(n15068), .B1(n15059), .B2(n20800), .C1(
        n15278), .C2(n15067), .ZN(P1_U2854) );
  INV_X1 U18594 ( .A(n15293), .ZN(n15141) );
  AOI22_X1 U18595 ( .A1(n15517), .A2(n20795), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n15065), .ZN(n15060) );
  OAI21_X1 U18596 ( .B1(n15141), .B2(n15067), .A(n15060), .ZN(P1_U2855) );
  OAI222_X1 U18597 ( .A1(n15307), .A2(n15070), .B1(n15061), .B2(n20800), .C1(
        n15529), .C2(n15068), .ZN(P1_U2856) );
  INV_X1 U18598 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15062) );
  OAI222_X1 U18599 ( .A1(n15319), .A2(n15070), .B1(n15062), .B2(n20800), .C1(
        n15538), .C2(n15068), .ZN(P1_U2857) );
  INV_X1 U18600 ( .A(n15546), .ZN(n15063) );
  OAI222_X1 U18601 ( .A1(n15153), .A2(n15070), .B1(n21352), .B2(n20800), .C1(
        n15063), .C2(n15068), .ZN(P1_U2858) );
  AOI22_X1 U18602 ( .A1(n15555), .A2(n20795), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n15065), .ZN(n15064) );
  OAI21_X1 U18603 ( .B1(n15157), .B2(n15067), .A(n15064), .ZN(P1_U2859) );
  AOI22_X1 U18604 ( .A1(n15569), .A2(n20795), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n15065), .ZN(n15066) );
  OAI21_X1 U18605 ( .B1(n15159), .B2(n15067), .A(n15066), .ZN(P1_U2860) );
  INV_X1 U18606 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15069) );
  OAI222_X1 U18607 ( .A1(n15164), .A2(n15070), .B1(n15069), .B2(n20800), .C1(
        n15572), .C2(n15068), .ZN(P1_U2861) );
  INV_X1 U18608 ( .A(DATAI_14_), .ZN(n15072) );
  MUX2_X1 U18609 ( .A(n15072), .B(n15071), .S(n15085), .Z(n20841) );
  OAI22_X1 U18610 ( .A1(n15144), .A2(n20841), .B1(n15150), .B2(n15073), .ZN(
        n15074) );
  AOI21_X1 U18611 ( .B1(n15146), .B2(BUF1_REG_30__SCAN_IN), .A(n15074), .ZN(
        n15076) );
  NAND2_X1 U18612 ( .A1(n15147), .A2(DATAI_30_), .ZN(n15075) );
  OAI211_X1 U18613 ( .C1(n15077), .C2(n15163), .A(n15076), .B(n15075), .ZN(
        P1_U2874) );
  INV_X1 U18614 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n15081) );
  INV_X1 U18615 ( .A(n15144), .ZN(n15136) );
  INV_X1 U18616 ( .A(DATAI_13_), .ZN(n15079) );
  NAND2_X1 U18617 ( .A1(n15085), .A2(BUF1_REG_13__SCAN_IN), .ZN(n15078) );
  OAI21_X1 U18618 ( .B1(n15085), .B2(n15079), .A(n15078), .ZN(n20837) );
  AOI22_X1 U18619 ( .A1(n15136), .A2(n20837), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n15154), .ZN(n15080) );
  OAI21_X1 U18620 ( .B1(n15138), .B2(n15081), .A(n15080), .ZN(n15082) );
  AOI21_X1 U18621 ( .B1(n15147), .B2(DATAI_29_), .A(n15082), .ZN(n15083) );
  OAI21_X1 U18622 ( .B1(n15084), .B2(n15163), .A(n15083), .ZN(P1_U2875) );
  INV_X1 U18623 ( .A(DATAI_12_), .ZN(n15086) );
  MUX2_X1 U18624 ( .A(n15086), .B(n17333), .S(n15085), .Z(n20834) );
  OAI22_X1 U18625 ( .A1(n15144), .A2(n20834), .B1(n15150), .B2(n20836), .ZN(
        n15087) );
  AOI21_X1 U18626 ( .B1(n15146), .B2(BUF1_REG_28__SCAN_IN), .A(n15087), .ZN(
        n15089) );
  NAND2_X1 U18627 ( .A1(n15147), .A2(DATAI_28_), .ZN(n15088) );
  OAI211_X1 U18628 ( .C1(n15185), .C2(n15163), .A(n15089), .B(n15088), .ZN(
        P1_U2876) );
  INV_X1 U18629 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n17310) );
  AOI22_X1 U18630 ( .A1(n15136), .A2(n15160), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n15154), .ZN(n15090) );
  OAI21_X1 U18631 ( .B1(n15138), .B2(n17310), .A(n15090), .ZN(n15091) );
  AOI21_X1 U18632 ( .B1(n15147), .B2(DATAI_27_), .A(n15091), .ZN(n15092) );
  OAI21_X1 U18633 ( .B1(n15093), .B2(n15163), .A(n15092), .ZN(P1_U2877) );
  INV_X1 U18634 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n17312) );
  AOI22_X1 U18635 ( .A1(n15136), .A2(n20831), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n15154), .ZN(n15094) );
  OAI21_X1 U18636 ( .B1(n15138), .B2(n17312), .A(n15094), .ZN(n15095) );
  AOI21_X1 U18637 ( .B1(n15147), .B2(DATAI_26_), .A(n15095), .ZN(n15096) );
  OAI21_X1 U18638 ( .B1(n15097), .B2(n15163), .A(n15096), .ZN(P1_U2878) );
  OAI22_X1 U18639 ( .A1(n15144), .A2(n20828), .B1(n15150), .B2(n20830), .ZN(
        n15098) );
  AOI21_X1 U18640 ( .B1(n15146), .B2(BUF1_REG_25__SCAN_IN), .A(n15098), .ZN(
        n15100) );
  NAND2_X1 U18641 ( .A1(n15147), .A2(DATAI_25_), .ZN(n15099) );
  OAI211_X1 U18642 ( .C1(n15101), .C2(n15163), .A(n15100), .B(n15099), .ZN(
        P1_U2879) );
  OAI22_X1 U18643 ( .A1(n15144), .A2(n15103), .B1(n15150), .B2(n15102), .ZN(
        n15104) );
  AOI21_X1 U18644 ( .B1(n15146), .B2(BUF1_REG_24__SCAN_IN), .A(n15104), .ZN(
        n15106) );
  NAND2_X1 U18645 ( .A1(n15147), .A2(DATAI_24_), .ZN(n15105) );
  OAI211_X1 U18646 ( .C1(n15222), .C2(n15163), .A(n15106), .B(n15105), .ZN(
        P1_U2880) );
  OAI22_X1 U18647 ( .A1(n15144), .A2(n15107), .B1(n15150), .B2(n13988), .ZN(
        n15108) );
  AOI21_X1 U18648 ( .B1(n15146), .B2(BUF1_REG_23__SCAN_IN), .A(n15108), .ZN(
        n15110) );
  NAND2_X1 U18649 ( .A1(n15147), .A2(DATAI_23_), .ZN(n15109) );
  OAI211_X1 U18650 ( .C1(n15111), .C2(n15163), .A(n15110), .B(n15109), .ZN(
        P1_U2881) );
  OAI22_X1 U18651 ( .A1(n15144), .A2(n15112), .B1(n15150), .B2(n13993), .ZN(
        n15113) );
  AOI21_X1 U18652 ( .B1(n15146), .B2(BUF1_REG_22__SCAN_IN), .A(n15113), .ZN(
        n15115) );
  NAND2_X1 U18653 ( .A1(n15147), .A2(DATAI_22_), .ZN(n15114) );
  OAI211_X1 U18654 ( .C1(n15243), .C2(n15163), .A(n15115), .B(n15114), .ZN(
        P1_U2882) );
  OAI22_X1 U18655 ( .A1(n15144), .A2(n15117), .B1(n15150), .B2(n15116), .ZN(
        n15118) );
  AOI21_X1 U18656 ( .B1(n15146), .B2(BUF1_REG_21__SCAN_IN), .A(n15118), .ZN(
        n15120) );
  NAND2_X1 U18657 ( .A1(n15147), .A2(DATAI_21_), .ZN(n15119) );
  OAI211_X1 U18658 ( .C1(n15121), .C2(n15163), .A(n15120), .B(n15119), .ZN(
        P1_U2883) );
  OAI22_X1 U18659 ( .A1(n15144), .A2(n15122), .B1(n15150), .B2(n13996), .ZN(
        n15123) );
  AOI21_X1 U18660 ( .B1(n15146), .B2(BUF1_REG_20__SCAN_IN), .A(n15123), .ZN(
        n15125) );
  NAND2_X1 U18661 ( .A1(n15147), .A2(DATAI_20_), .ZN(n15124) );
  OAI211_X1 U18662 ( .C1(n15262), .C2(n15163), .A(n15125), .B(n15124), .ZN(
        P1_U2884) );
  OAI22_X1 U18663 ( .A1(n15144), .A2(n15126), .B1(n15150), .B2(n13990), .ZN(
        n15127) );
  AOI21_X1 U18664 ( .B1(n15146), .B2(BUF1_REG_19__SCAN_IN), .A(n15127), .ZN(
        n15129) );
  NAND2_X1 U18665 ( .A1(n15147), .A2(DATAI_19_), .ZN(n15128) );
  OAI211_X1 U18666 ( .C1(n15130), .C2(n15163), .A(n15129), .B(n15128), .ZN(
        P1_U2885) );
  OAI22_X1 U18667 ( .A1(n15144), .A2(n15131), .B1(n15150), .B2(n13999), .ZN(
        n15132) );
  AOI21_X1 U18668 ( .B1(n15146), .B2(BUF1_REG_18__SCAN_IN), .A(n15132), .ZN(
        n15134) );
  NAND2_X1 U18669 ( .A1(n15147), .A2(DATAI_18_), .ZN(n15133) );
  OAI211_X1 U18670 ( .C1(n15278), .C2(n15163), .A(n15134), .B(n15133), .ZN(
        P1_U2886) );
  INV_X1 U18671 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n21348) );
  AOI22_X1 U18672 ( .A1(n15136), .A2(n15135), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n15154), .ZN(n15137) );
  OAI21_X1 U18673 ( .B1(n15138), .B2(n21348), .A(n15137), .ZN(n15139) );
  AOI21_X1 U18674 ( .B1(n15147), .B2(DATAI_17_), .A(n15139), .ZN(n15140) );
  OAI21_X1 U18675 ( .B1(n15141), .B2(n15163), .A(n15140), .ZN(P1_U2887) );
  OAI22_X1 U18676 ( .A1(n15144), .A2(n15143), .B1(n15150), .B2(n15142), .ZN(
        n15145) );
  AOI21_X1 U18677 ( .B1(n15146), .B2(BUF1_REG_16__SCAN_IN), .A(n15145), .ZN(
        n15149) );
  NAND2_X1 U18678 ( .A1(n15147), .A2(DATAI_16_), .ZN(n15148) );
  OAI211_X1 U18679 ( .C1(n15307), .C2(n15163), .A(n15149), .B(n15148), .ZN(
        P1_U2888) );
  OAI222_X1 U18680 ( .A1(n15163), .A2(n15319), .B1(n15161), .B2(n15151), .C1(
        n20803), .C2(n15150), .ZN(P1_U2889) );
  INV_X1 U18681 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n15152) );
  OAI222_X1 U18682 ( .A1(n15153), .A2(n15163), .B1(n20841), .B2(n15161), .C1(
        n15152), .C2(n15150), .ZN(P1_U2890) );
  AOI22_X1 U18683 ( .A1(n15155), .A2(n20837), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15154), .ZN(n15156) );
  OAI21_X1 U18684 ( .B1(n15157), .B2(n15163), .A(n15156), .ZN(P1_U2891) );
  OAI222_X1 U18685 ( .A1(n15163), .A2(n15159), .B1(n20834), .B2(n15161), .C1(
        n15158), .C2(n15150), .ZN(P1_U2892) );
  INV_X1 U18686 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20808) );
  INV_X1 U18687 ( .A(n15160), .ZN(n15162) );
  OAI222_X1 U18688 ( .A1(n15164), .A2(n15163), .B1(n15150), .B2(n20808), .C1(
        n15162), .C2(n15161), .ZN(P1_U2893) );
  XNOR2_X1 U18689 ( .A(n15165), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15399) );
  NAND2_X1 U18690 ( .A1(n15166), .A2(n15304), .ZN(n15167) );
  NAND2_X1 U18691 ( .A1(n20916), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15393) );
  OAI211_X1 U18692 ( .C1(n15168), .C2(n15301), .A(n15167), .B(n15393), .ZN(
        n15169) );
  AOI21_X1 U18693 ( .B1(n15170), .B2(n20884), .A(n15169), .ZN(n15171) );
  OAI21_X1 U18694 ( .B1(n15399), .B2(n20712), .A(n15171), .ZN(P1_U2969) );
  NAND2_X1 U18695 ( .A1(n15366), .A2(n15400), .ZN(n15172) );
  NOR2_X1 U18696 ( .A1(n20893), .A2(n21272), .ZN(n15403) );
  AOI21_X1 U18697 ( .B1(n20882), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15403), .ZN(n15173) );
  OAI21_X1 U18698 ( .B1(n15174), .B2(n20881), .A(n15173), .ZN(n15175) );
  AOI21_X1 U18699 ( .B1(n15176), .B2(n20884), .A(n15175), .ZN(n15177) );
  OAI21_X1 U18700 ( .B1(n15408), .B2(n20712), .A(n15177), .ZN(P1_U2970) );
  NOR4_X1 U18701 ( .A1(n15178), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15179) );
  NAND2_X1 U18702 ( .A1(n10101), .A2(n15179), .ZN(n15182) );
  NAND3_X1 U18703 ( .A1(n15180), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15181) );
  MUX2_X1 U18704 ( .A(n15182), .B(n15181), .S(n15366), .Z(n15183) );
  XNOR2_X1 U18705 ( .A(n15183), .B(n15413), .ZN(n15417) );
  NAND2_X1 U18706 ( .A1(n20916), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15412) );
  OAI21_X1 U18707 ( .B1(n15301), .B2(n15184), .A(n15412), .ZN(n15186) );
  NAND2_X1 U18708 ( .A1(n15189), .A2(n15188), .ZN(n15190) );
  XNOR2_X1 U18709 ( .A(n15190), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15426) );
  NOR2_X1 U18710 ( .A1(n20893), .A2(n21267), .ZN(n15418) );
  AOI21_X1 U18711 ( .B1(n20882), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15418), .ZN(n15191) );
  OAI21_X1 U18712 ( .B1(n15192), .B2(n20881), .A(n15191), .ZN(n15193) );
  AOI21_X1 U18713 ( .B1(n15194), .B2(n20884), .A(n15193), .ZN(n15195) );
  OAI21_X1 U18714 ( .B1(n15426), .B2(n20712), .A(n15195), .ZN(P1_U2972) );
  OAI21_X1 U18715 ( .B1(n15228), .B2(n15430), .A(n15366), .ZN(n15196) );
  NAND2_X1 U18716 ( .A1(n15197), .A2(n15196), .ZN(n15198) );
  XNOR2_X1 U18717 ( .A(n15198), .B(n15431), .ZN(n15439) );
  NAND2_X1 U18718 ( .A1(n15199), .A2(n15304), .ZN(n15200) );
  NAND2_X1 U18719 ( .A1(n20916), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15434) );
  OAI211_X1 U18720 ( .C1(n15301), .C2(n15201), .A(n15200), .B(n15434), .ZN(
        n15202) );
  AOI21_X1 U18721 ( .B1(n15203), .B2(n20884), .A(n15202), .ZN(n15204) );
  OAI21_X1 U18722 ( .B1(n20712), .B2(n15439), .A(n15204), .ZN(P1_U2973) );
  MUX2_X1 U18723 ( .A(n15452), .B(n15205), .S(n15374), .Z(n15206) );
  INV_X1 U18724 ( .A(n15206), .ZN(n15209) );
  NAND2_X1 U18725 ( .A1(n15219), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15208) );
  NAND2_X1 U18726 ( .A1(n15209), .A2(n15208), .ZN(n15211) );
  XNOR2_X1 U18727 ( .A(n15211), .B(n15210), .ZN(n15446) );
  NOR2_X1 U18728 ( .A1(n20893), .A2(n15212), .ZN(n15441) );
  AOI21_X1 U18729 ( .B1(n20882), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15441), .ZN(n15213) );
  OAI21_X1 U18730 ( .B1(n15214), .B2(n20881), .A(n15213), .ZN(n15215) );
  AOI21_X1 U18731 ( .B1(n15216), .B2(n20884), .A(n15215), .ZN(n15217) );
  OAI21_X1 U18732 ( .B1(n20712), .B2(n15446), .A(n15217), .ZN(P1_U2974) );
  NAND2_X1 U18733 ( .A1(n15219), .A2(n15228), .ZN(n15218) );
  MUX2_X1 U18734 ( .A(n15219), .B(n15218), .S(n15374), .Z(n15220) );
  XNOR2_X1 U18735 ( .A(n15220), .B(n15452), .ZN(n15457) );
  OR2_X1 U18736 ( .A1(n20893), .A2(n21263), .ZN(n15451) );
  OAI21_X1 U18737 ( .B1(n15301), .B2(n15221), .A(n15451), .ZN(n15224) );
  NOR2_X1 U18738 ( .A1(n15222), .A2(n15382), .ZN(n15223) );
  AOI211_X1 U18739 ( .C1(n15304), .C2(n15225), .A(n15224), .B(n15223), .ZN(
        n15226) );
  OAI21_X1 U18740 ( .B1(n20712), .B2(n15457), .A(n15226), .ZN(P1_U2975) );
  XNOR2_X1 U18741 ( .A(n15366), .B(n15448), .ZN(n15227) );
  XNOR2_X1 U18742 ( .A(n15228), .B(n15227), .ZN(n15465) );
  INV_X1 U18743 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21260) );
  NOR2_X1 U18744 ( .A1(n20893), .A2(n21260), .ZN(n15458) );
  AOI21_X1 U18745 ( .B1(n20882), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15458), .ZN(n15229) );
  OAI21_X1 U18746 ( .B1(n20881), .B2(n15230), .A(n15229), .ZN(n15231) );
  AOI21_X1 U18747 ( .B1(n15232), .B2(n20884), .A(n15231), .ZN(n15233) );
  OAI21_X1 U18748 ( .B1(n15465), .B2(n20712), .A(n15233), .ZN(P1_U2976) );
  INV_X1 U18749 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21259) );
  NOR2_X1 U18750 ( .A1(n20893), .A2(n21259), .ZN(n15469) );
  INV_X1 U18751 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15234) );
  NOR2_X1 U18752 ( .A1(n15301), .A2(n15234), .ZN(n15235) );
  AOI211_X1 U18753 ( .C1(n15304), .C2(n15236), .A(n15469), .B(n15235), .ZN(
        n15242) );
  XNOR2_X1 U18754 ( .A(n15366), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15273) );
  NAND2_X1 U18755 ( .A1(n15237), .A2(n15273), .ZN(n15272) );
  NOR3_X1 U18756 ( .A1(n15272), .A2(n15244), .A3(n21379), .ZN(n15239) );
  OAI21_X1 U18757 ( .B1(n15239), .B2(n15374), .A(n15238), .ZN(n15240) );
  XNOR2_X1 U18758 ( .A(n15240), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15466) );
  NAND2_X1 U18759 ( .A1(n15466), .A2(n20887), .ZN(n15241) );
  OAI211_X1 U18760 ( .C1(n15243), .C2(n15382), .A(n15242), .B(n15241), .ZN(
        P1_U2977) );
  NOR4_X1 U18761 ( .A1(n15237), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A4(n15366), .ZN(n15255) );
  NOR3_X1 U18762 ( .A1(n15272), .A2(n15286), .A3(n15244), .ZN(n15245) );
  AOI21_X1 U18763 ( .B1(n15255), .B2(n15246), .A(n15245), .ZN(n15247) );
  XNOR2_X1 U18764 ( .A(n15247), .B(n21379), .ZN(n15482) );
  INV_X1 U18765 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21257) );
  NOR2_X1 U18766 ( .A1(n20893), .A2(n21257), .ZN(n15476) );
  AOI21_X1 U18767 ( .B1(n20882), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15476), .ZN(n15248) );
  OAI21_X1 U18768 ( .B1(n20881), .B2(n15249), .A(n15248), .ZN(n15250) );
  AOI21_X1 U18769 ( .B1(n15251), .B2(n20884), .A(n15250), .ZN(n15252) );
  OAI21_X1 U18770 ( .B1(n15482), .B2(n20712), .A(n15252), .ZN(P1_U2978) );
  NOR3_X1 U18771 ( .A1(n15272), .A2(n15374), .A3(n15253), .ZN(n15254) );
  NOR2_X1 U18772 ( .A1(n15255), .A2(n15254), .ZN(n15256) );
  XNOR2_X1 U18773 ( .A(n15256), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15483) );
  NAND2_X1 U18774 ( .A1(n15483), .A2(n20887), .ZN(n15261) );
  INV_X1 U18775 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21254) );
  NOR2_X1 U18776 ( .A1(n20893), .A2(n21254), .ZN(n15486) );
  NOR2_X1 U18777 ( .A1(n15301), .A2(n15257), .ZN(n15258) );
  AOI211_X1 U18778 ( .C1(n15304), .C2(n15259), .A(n15486), .B(n15258), .ZN(
        n15260) );
  OAI211_X1 U18779 ( .C1(n15382), .C2(n15262), .A(n15261), .B(n15260), .ZN(
        P1_U2979) );
  NOR2_X1 U18780 ( .A1(n15366), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15263) );
  MUX2_X1 U18781 ( .A(n15353), .B(n15263), .S(n15272), .Z(n15264) );
  XNOR2_X1 U18782 ( .A(n15264), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15497) );
  NOR2_X1 U18783 ( .A1(n20893), .A2(n15265), .ZN(n15490) );
  AOI21_X1 U18784 ( .B1(n20882), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15490), .ZN(n15266) );
  OAI21_X1 U18785 ( .B1(n20881), .B2(n15267), .A(n15266), .ZN(n15268) );
  AOI21_X1 U18786 ( .B1(n15269), .B2(n20884), .A(n15268), .ZN(n15270) );
  OAI21_X1 U18787 ( .B1(n20712), .B2(n15497), .A(n15270), .ZN(P1_U2980) );
  OR2_X1 U18788 ( .A1(n20893), .A2(n21251), .ZN(n15503) );
  OAI21_X1 U18789 ( .B1(n15301), .B2(n15271), .A(n15503), .ZN(n15275) );
  OAI21_X1 U18790 ( .B1(n15237), .B2(n15273), .A(n15272), .ZN(n15509) );
  NOR2_X1 U18791 ( .A1(n15509), .A2(n20712), .ZN(n15274) );
  AOI211_X1 U18792 ( .C1(n15304), .C2(n15276), .A(n15275), .B(n15274), .ZN(
        n15277) );
  OAI21_X1 U18793 ( .B1(n15278), .B2(n15382), .A(n15277), .ZN(P1_U2981) );
  OAI21_X1 U18794 ( .B1(n15385), .B2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n15383), .ZN(n15280) );
  NAND2_X1 U18795 ( .A1(n15385), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15279) );
  NAND2_X1 U18796 ( .A1(n15280), .A2(n15279), .ZN(n15376) );
  INV_X1 U18797 ( .A(n15281), .ZN(n15282) );
  OR2_X2 U18798 ( .A1(n15376), .A2(n15282), .ZN(n15363) );
  OAI21_X2 U18799 ( .B1(n15374), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15363), .ZN(n15365) );
  INV_X1 U18800 ( .A(n15283), .ZN(n15297) );
  NOR2_X1 U18801 ( .A1(n15297), .A2(n15332), .ZN(n15285) );
  AOI21_X1 U18802 ( .B1(n15365), .B2(n15285), .A(n15284), .ZN(n15288) );
  NOR2_X1 U18803 ( .A1(n15288), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15287) );
  MUX2_X1 U18804 ( .A(n15288), .B(n15287), .S(n15286), .Z(n15289) );
  XNOR2_X1 U18805 ( .A(n15289), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15519) );
  AND2_X1 U18806 ( .A1(n20916), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15516) );
  AOI21_X1 U18807 ( .B1(n20882), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15516), .ZN(n15290) );
  OAI21_X1 U18808 ( .B1(n20881), .B2(n15291), .A(n15290), .ZN(n15292) );
  AOI21_X1 U18809 ( .B1(n15293), .B2(n20884), .A(n15292), .ZN(n15294) );
  OAI21_X1 U18810 ( .B1(n15519), .B2(n20712), .A(n15294), .ZN(P1_U2982) );
  INV_X1 U18811 ( .A(n15332), .ZN(n15295) );
  OAI21_X1 U18812 ( .B1(n15365), .B2(n15296), .A(n15295), .ZN(n15308) );
  OAI21_X1 U18813 ( .B1(n15308), .B2(n15297), .A(n15311), .ZN(n15299) );
  XNOR2_X1 U18814 ( .A(n15299), .B(n15298), .ZN(n15520) );
  NAND2_X1 U18815 ( .A1(n15520), .A2(n20887), .ZN(n15306) );
  NOR2_X1 U18816 ( .A1(n20893), .A2(n21249), .ZN(n15525) );
  NOR2_X1 U18817 ( .A1(n15301), .A2(n15300), .ZN(n15302) );
  AOI211_X1 U18818 ( .C1(n15304), .C2(n15303), .A(n15525), .B(n15302), .ZN(
        n15305) );
  OAI211_X1 U18819 ( .C1(n15382), .C2(n15307), .A(n15306), .B(n15305), .ZN(
        P1_U2983) );
  INV_X1 U18820 ( .A(n15308), .ZN(n15310) );
  NAND2_X1 U18821 ( .A1(n15310), .A2(n15309), .ZN(n15314) );
  NAND2_X1 U18822 ( .A1(n15312), .A2(n15311), .ZN(n15313) );
  XNOR2_X1 U18823 ( .A(n15314), .B(n15313), .ZN(n15530) );
  NAND2_X1 U18824 ( .A1(n15530), .A2(n20887), .ZN(n15318) );
  NOR2_X1 U18825 ( .A1(n20893), .A2(n21247), .ZN(n15533) );
  NOR2_X1 U18826 ( .A1(n20881), .A2(n15315), .ZN(n15316) );
  AOI211_X1 U18827 ( .C1(n20882), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15533), .B(n15316), .ZN(n15317) );
  OAI211_X1 U18828 ( .C1(n15382), .C2(n15319), .A(n15318), .B(n15317), .ZN(
        P1_U2984) );
  INV_X1 U18829 ( .A(n15365), .ZN(n15354) );
  OAI21_X1 U18830 ( .B1(n15354), .B2(n15332), .A(n15320), .ZN(n15322) );
  NAND2_X1 U18831 ( .A1(n15322), .A2(n15321), .ZN(n15324) );
  XNOR2_X1 U18832 ( .A(n15366), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15323) );
  XNOR2_X1 U18833 ( .A(n15324), .B(n15323), .ZN(n15549) );
  INV_X1 U18834 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21244) );
  NOR2_X1 U18835 ( .A1(n20893), .A2(n21244), .ZN(n15545) );
  AOI21_X1 U18836 ( .B1(n20882), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15545), .ZN(n15325) );
  OAI21_X1 U18837 ( .B1(n20881), .B2(n15326), .A(n15325), .ZN(n15327) );
  AOI21_X1 U18838 ( .B1(n15328), .B2(n20884), .A(n15327), .ZN(n15329) );
  OAI21_X1 U18839 ( .B1(n15549), .B2(n20712), .A(n15329), .ZN(P1_U2985) );
  INV_X1 U18840 ( .A(n15330), .ZN(n15331) );
  NOR2_X1 U18841 ( .A1(n15365), .A2(n15331), .ZN(n15342) );
  OAI21_X1 U18842 ( .B1(n15342), .B2(n15332), .A(n15343), .ZN(n15333) );
  XNOR2_X1 U18843 ( .A(n15334), .B(n15333), .ZN(n15557) );
  NAND2_X1 U18844 ( .A1(n20916), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n15551) );
  NAND2_X1 U18845 ( .A1(n20882), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15335) );
  OAI211_X1 U18846 ( .C1(n20881), .C2(n15336), .A(n15551), .B(n15335), .ZN(
        n15337) );
  AOI21_X1 U18847 ( .B1(n15338), .B2(n20884), .A(n15337), .ZN(n15339) );
  OAI21_X1 U18848 ( .B1(n15557), .B2(n20712), .A(n15339), .ZN(P1_U2986) );
  INV_X1 U18849 ( .A(n15340), .ZN(n15341) );
  NOR2_X1 U18850 ( .A1(n15342), .A2(n15341), .ZN(n15346) );
  NAND2_X1 U18851 ( .A1(n15344), .A2(n15343), .ZN(n15345) );
  XNOR2_X1 U18852 ( .A(n15346), .B(n15345), .ZN(n15571) );
  INV_X1 U18853 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15347) );
  NOR2_X1 U18854 ( .A1(n20893), .A2(n15347), .ZN(n15568) );
  AOI21_X1 U18855 ( .B1(n20882), .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15568), .ZN(n15348) );
  OAI21_X1 U18856 ( .B1(n20881), .B2(n15349), .A(n15348), .ZN(n15350) );
  AOI21_X1 U18857 ( .B1(n15351), .B2(n20884), .A(n15350), .ZN(n15352) );
  OAI21_X1 U18858 ( .B1(n15571), .B2(n20712), .A(n15352), .ZN(P1_U2987) );
  NAND2_X1 U18859 ( .A1(n15374), .A2(n15364), .ZN(n15355) );
  NAND3_X1 U18860 ( .A1(n15354), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15353), .ZN(n15369) );
  OAI21_X1 U18861 ( .B1(n15363), .B2(n15355), .A(n15369), .ZN(n15356) );
  XNOR2_X1 U18862 ( .A(n15356), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15581) );
  NOR2_X1 U18863 ( .A1(n20893), .A2(n15357), .ZN(n15574) );
  AOI21_X1 U18864 ( .B1(n20882), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n15574), .ZN(n15358) );
  OAI21_X1 U18865 ( .B1(n20881), .B2(n15359), .A(n15358), .ZN(n15360) );
  AOI21_X1 U18866 ( .B1(n15361), .B2(n20884), .A(n15360), .ZN(n15362) );
  OAI21_X1 U18867 ( .B1(n15581), .B2(n20712), .A(n15362), .ZN(P1_U2988) );
  XNOR2_X1 U18868 ( .A(n15363), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15368) );
  NAND2_X1 U18869 ( .A1(n15365), .A2(n15364), .ZN(n15367) );
  MUX2_X1 U18870 ( .A(n15368), .B(n15367), .S(n15366), .Z(n15370) );
  NAND2_X1 U18871 ( .A1(n15582), .A2(n20887), .ZN(n15373) );
  INV_X1 U18872 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21238) );
  NOR2_X1 U18873 ( .A1(n20893), .A2(n21238), .ZN(n15590) );
  NOR2_X1 U18874 ( .A1(n20881), .A2(n17156), .ZN(n15371) );
  AOI211_X1 U18875 ( .C1(n20882), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15590), .B(n15371), .ZN(n15372) );
  OAI211_X1 U18876 ( .C1(n15382), .C2(n17155), .A(n15373), .B(n15372), .ZN(
        P1_U2989) );
  XNOR2_X1 U18877 ( .A(n15374), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15375) );
  XNOR2_X1 U18878 ( .A(n15376), .B(n15375), .ZN(n17187) );
  NAND2_X1 U18879 ( .A1(n17187), .A2(n20887), .ZN(n15380) );
  NOR2_X1 U18880 ( .A1(n20893), .A2(n21237), .ZN(n17184) );
  NOR2_X1 U18881 ( .A1(n20881), .A2(n15377), .ZN(n15378) );
  AOI211_X1 U18882 ( .C1(n20882), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n17184), .B(n15378), .ZN(n15379) );
  OAI211_X1 U18883 ( .C1(n15382), .C2(n15381), .A(n15380), .B(n15379), .ZN(
        P1_U2990) );
  XOR2_X1 U18884 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n15383), .Z(
        n15384) );
  XNOR2_X1 U18885 ( .A(n15385), .B(n15384), .ZN(n15610) );
  NOR2_X1 U18886 ( .A1(n20893), .A2(n21234), .ZN(n15604) );
  AOI21_X1 U18887 ( .B1(n20882), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n15604), .ZN(n15386) );
  OAI21_X1 U18888 ( .B1(n20881), .B2(n15387), .A(n15386), .ZN(n15388) );
  AOI21_X1 U18889 ( .B1(n15389), .B2(n20884), .A(n15388), .ZN(n15390) );
  OAI21_X1 U18890 ( .B1(n15610), .B2(n20712), .A(n15390), .ZN(P1_U2991) );
  INV_X1 U18891 ( .A(n15391), .ZN(n15392) );
  AOI21_X1 U18892 ( .B1(n15419), .B2(n15392), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15394) );
  OAI21_X1 U18893 ( .B1(n15395), .B2(n15394), .A(n15393), .ZN(n15396) );
  AOI21_X1 U18894 ( .B1(n15397), .B2(n17191), .A(n15396), .ZN(n15398) );
  OAI21_X1 U18895 ( .B1(n15399), .B2(n20933), .A(n15398), .ZN(P1_U3001) );
  INV_X1 U18896 ( .A(n15419), .ZN(n15401) );
  INV_X1 U18897 ( .A(n15400), .ZN(n15410) );
  NOR3_X1 U18898 ( .A1(n15401), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15410), .ZN(n15402) );
  AOI211_X1 U18899 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15404), .A(
        n15403), .B(n15402), .ZN(n15407) );
  NAND2_X1 U18900 ( .A1(n15405), .A2(n17191), .ZN(n15406) );
  NAND3_X1 U18901 ( .A1(n15419), .A2(n15410), .A3(n15409), .ZN(n15411) );
  OAI211_X1 U18902 ( .C1(n15422), .C2(n15413), .A(n15412), .B(n15411), .ZN(
        n15414) );
  AOI21_X1 U18903 ( .B1(n15415), .B2(n17191), .A(n15414), .ZN(n15416) );
  OAI21_X1 U18904 ( .B1(n15417), .B2(n20933), .A(n15416), .ZN(P1_U3003) );
  AOI21_X1 U18905 ( .B1(n15419), .B2(n15421), .A(n15418), .ZN(n15420) );
  OAI21_X1 U18906 ( .B1(n15422), .B2(n15421), .A(n15420), .ZN(n15423) );
  AOI21_X1 U18907 ( .B1(n15424), .B2(n17191), .A(n15423), .ZN(n15425) );
  OAI21_X1 U18908 ( .B1(n15426), .B2(n20933), .A(n15425), .ZN(P1_U3004) );
  INV_X1 U18909 ( .A(n15427), .ZN(n15437) );
  INV_X1 U18910 ( .A(n15428), .ZN(n15442) );
  NOR3_X1 U18911 ( .A1(n15461), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n15429), .ZN(n15440) );
  OAI21_X1 U18912 ( .B1(n15442), .B2(n15440), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15435) );
  INV_X1 U18913 ( .A(n15461), .ZN(n15449) );
  INV_X1 U18914 ( .A(n15430), .ZN(n15432) );
  NAND3_X1 U18915 ( .A1(n15449), .A2(n15432), .A3(n15431), .ZN(n15433) );
  NAND3_X1 U18916 ( .A1(n15435), .A2(n15434), .A3(n15433), .ZN(n15436) );
  AOI21_X1 U18917 ( .B1(n15437), .B2(n17191), .A(n15436), .ZN(n15438) );
  OAI21_X1 U18918 ( .B1(n15439), .B2(n20933), .A(n15438), .ZN(P1_U3005) );
  AOI211_X1 U18919 ( .C1(n15442), .C2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15441), .B(n15440), .ZN(n15445) );
  NAND2_X1 U18920 ( .A1(n15443), .A2(n17191), .ZN(n15444) );
  OAI211_X1 U18921 ( .C1(n15446), .C2(n20933), .A(n15445), .B(n15444), .ZN(
        P1_U3006) );
  AOI21_X1 U18922 ( .B1(n15448), .B2(n20910), .A(n15447), .ZN(n15453) );
  NAND3_X1 U18923 ( .A1(n15449), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n15452), .ZN(n15450) );
  OAI211_X1 U18924 ( .C1(n15453), .C2(n15452), .A(n15451), .B(n15450), .ZN(
        n15454) );
  AOI21_X1 U18925 ( .B1(n15455), .B2(n17191), .A(n15454), .ZN(n15456) );
  OAI21_X1 U18926 ( .B1(n15457), .B2(n20933), .A(n15456), .ZN(P1_U3007) );
  AOI21_X1 U18927 ( .B1(n15459), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15458), .ZN(n15460) );
  OAI21_X1 U18928 ( .B1(n15461), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15460), .ZN(n15462) );
  AOI21_X1 U18929 ( .B1(n15463), .B2(n17191), .A(n15462), .ZN(n15464) );
  OAI21_X1 U18930 ( .B1(n15465), .B2(n20933), .A(n15464), .ZN(P1_U3008) );
  NAND2_X1 U18931 ( .A1(n15466), .A2(n20922), .ZN(n15472) );
  XNOR2_X1 U18932 ( .A(n15467), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15470) );
  NOR2_X1 U18933 ( .A1(n15474), .A2(n15467), .ZN(n15468) );
  AOI211_X1 U18934 ( .C1(n15470), .C2(n15477), .A(n15469), .B(n15468), .ZN(
        n15471) );
  OAI211_X1 U18935 ( .C1(n20895), .C2(n15473), .A(n15472), .B(n15471), .ZN(
        P1_U3009) );
  NOR2_X1 U18936 ( .A1(n15474), .A2(n21379), .ZN(n15475) );
  AOI211_X1 U18937 ( .C1(n15477), .C2(n21379), .A(n15476), .B(n15475), .ZN(
        n15481) );
  INV_X1 U18938 ( .A(n15478), .ZN(n15479) );
  NAND2_X1 U18939 ( .A1(n15479), .A2(n17191), .ZN(n15480) );
  OAI211_X1 U18940 ( .C1(n15482), .C2(n20933), .A(n15481), .B(n15480), .ZN(
        P1_U3010) );
  NAND2_X1 U18941 ( .A1(n15483), .A2(n20922), .ZN(n15488) );
  XNOR2_X1 U18942 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15484) );
  NOR2_X1 U18943 ( .A1(n15493), .A2(n15484), .ZN(n15485) );
  AOI211_X1 U18944 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15491), .A(
        n15486), .B(n15485), .ZN(n15487) );
  OAI211_X1 U18945 ( .C1(n20895), .C2(n15489), .A(n15488), .B(n15487), .ZN(
        P1_U3011) );
  AOI21_X1 U18946 ( .B1(n15491), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15490), .ZN(n15492) );
  OAI21_X1 U18947 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15493), .A(
        n15492), .ZN(n15494) );
  AOI21_X1 U18948 ( .B1(n15495), .B2(n17191), .A(n15494), .ZN(n15496) );
  OAI21_X1 U18949 ( .B1(n15497), .B2(n20933), .A(n15496), .ZN(P1_U3012) );
  INV_X1 U18950 ( .A(n15498), .ZN(n15507) );
  INV_X1 U18951 ( .A(n20912), .ZN(n15600) );
  AND2_X1 U18952 ( .A1(n15542), .A2(n15559), .ZN(n15500) );
  OAI21_X1 U18953 ( .B1(n15600), .B2(n15500), .A(n15499), .ZN(n15550) );
  AOI21_X1 U18954 ( .B1(n15521), .B2(n15501), .A(n15550), .ZN(n15512) );
  NOR2_X1 U18955 ( .A1(n15512), .A2(n15502), .ZN(n15506) );
  OAI21_X1 U18956 ( .B1(n15504), .B2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15503), .ZN(n15505) );
  AOI211_X1 U18957 ( .C1(n15507), .C2(n17191), .A(n15506), .B(n15505), .ZN(
        n15508) );
  OAI21_X1 U18958 ( .B1(n15509), .B2(n20933), .A(n15508), .ZN(P1_U3013) );
  INV_X1 U18959 ( .A(n15510), .ZN(n15553) );
  NOR3_X1 U18960 ( .A1(n15553), .A2(n15522), .A3(n15511), .ZN(n15535) );
  NAND3_X1 U18961 ( .A1(n15535), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15513) );
  AOI21_X1 U18962 ( .B1(n15514), .B2(n15513), .A(n15512), .ZN(n15515) );
  AOI211_X1 U18963 ( .C1(n15517), .C2(n17191), .A(n15516), .B(n15515), .ZN(
        n15518) );
  OAI21_X1 U18964 ( .B1(n15519), .B2(n20933), .A(n15518), .ZN(P1_U3014) );
  NAND2_X1 U18965 ( .A1(n15520), .A2(n20922), .ZN(n15528) );
  XNOR2_X1 U18966 ( .A(n15534), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15526) );
  AOI21_X1 U18967 ( .B1(n15522), .B2(n15521), .A(n15550), .ZN(n15531) );
  NOR2_X1 U18968 ( .A1(n15531), .A2(n15523), .ZN(n15524) );
  AOI211_X1 U18969 ( .C1(n15535), .C2(n15526), .A(n15525), .B(n15524), .ZN(
        n15527) );
  OAI211_X1 U18970 ( .C1(n20895), .C2(n15529), .A(n15528), .B(n15527), .ZN(
        P1_U3015) );
  NAND2_X1 U18971 ( .A1(n15530), .A2(n20922), .ZN(n15537) );
  NOR2_X1 U18972 ( .A1(n15531), .A2(n15534), .ZN(n15532) );
  AOI211_X1 U18973 ( .C1(n15535), .C2(n15534), .A(n15533), .B(n15532), .ZN(
        n15536) );
  OAI211_X1 U18974 ( .C1(n20895), .C2(n15538), .A(n15537), .B(n15536), .ZN(
        P1_U3016) );
  NAND2_X1 U18975 ( .A1(n20910), .A2(n20915), .ZN(n15596) );
  INV_X1 U18976 ( .A(n20914), .ZN(n15539) );
  NAND2_X1 U18977 ( .A1(n20891), .A2(n15539), .ZN(n15540) );
  INV_X1 U18978 ( .A(n15542), .ZN(n15543) );
  NOR3_X1 U18979 ( .A1(n17200), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n15543), .ZN(n15544) );
  AOI211_X1 U18980 ( .C1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n15550), .A(
        n15545), .B(n15544), .ZN(n15548) );
  NAND2_X1 U18981 ( .A1(n15546), .A2(n17191), .ZN(n15547) );
  OAI211_X1 U18982 ( .C1(n15549), .C2(n20933), .A(n15548), .B(n15547), .ZN(
        P1_U3017) );
  NAND2_X1 U18983 ( .A1(n15550), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15552) );
  OAI211_X1 U18984 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n15553), .A(
        n15552), .B(n15551), .ZN(n15554) );
  AOI21_X1 U18985 ( .B1(n15555), .B2(n17191), .A(n15554), .ZN(n15556) );
  OAI21_X1 U18986 ( .B1(n15557), .B2(n20933), .A(n15556), .ZN(P1_U3018) );
  INV_X1 U18987 ( .A(n20891), .ZN(n20920) );
  INV_X1 U18988 ( .A(n15587), .ZN(n15558) );
  INV_X1 U18989 ( .A(n15583), .ZN(n20911) );
  AOI21_X1 U18990 ( .B1(n20891), .B2(n15558), .A(n20911), .ZN(n15598) );
  INV_X1 U18991 ( .A(n15577), .ZN(n15561) );
  INV_X1 U18992 ( .A(n15559), .ZN(n15560) );
  OAI21_X1 U18993 ( .B1(n15561), .B2(n15560), .A(n20912), .ZN(n15562) );
  OAI211_X1 U18994 ( .C1(n15563), .C2(n20920), .A(n15598), .B(n15562), .ZN(
        n15575) );
  AOI21_X1 U18995 ( .B1(n15576), .B2(n20910), .A(n15575), .ZN(n15566) );
  INV_X1 U18996 ( .A(n17200), .ZN(n15578) );
  NAND3_X1 U18997 ( .A1(n15578), .A2(n15563), .A3(n15565), .ZN(n15564) );
  OAI21_X1 U18998 ( .B1(n15566), .B2(n15565), .A(n15564), .ZN(n15567) );
  AOI211_X1 U18999 ( .C1(n17191), .C2(n15569), .A(n15568), .B(n15567), .ZN(
        n15570) );
  OAI21_X1 U19000 ( .B1(n15571), .B2(n20933), .A(n15570), .ZN(P1_U3019) );
  NOR2_X1 U19001 ( .A1(n15572), .A2(n20895), .ZN(n15573) );
  AOI211_X1 U19002 ( .C1(n15575), .C2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15574), .B(n15573), .ZN(n15580) );
  NAND3_X1 U19003 ( .A1(n15578), .A2(n15577), .A3(n15576), .ZN(n15579) );
  OAI211_X1 U19004 ( .C1(n15581), .C2(n20933), .A(n15580), .B(n15579), .ZN(
        P1_U3020) );
  INV_X1 U19005 ( .A(n15582), .ZN(n15595) );
  OAI21_X1 U19006 ( .B1(n15600), .B2(n20915), .A(n15583), .ZN(n20890) );
  NOR2_X1 U19007 ( .A1(n15584), .A2(n20890), .ZN(n15588) );
  INV_X1 U19008 ( .A(n15585), .ZN(n15586) );
  AOI21_X1 U19009 ( .B1(n15588), .B2(n15587), .A(n15586), .ZN(n17186) );
  INV_X1 U19010 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21388) );
  INV_X1 U19011 ( .A(n17196), .ZN(n15589) );
  NAND3_X1 U19012 ( .A1(n15589), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17190) );
  XNOR2_X1 U19013 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15592) );
  AOI21_X1 U19014 ( .B1(n17151), .B2(n17191), .A(n15590), .ZN(n15591) );
  OAI21_X1 U19015 ( .B1(n17190), .B2(n15592), .A(n15591), .ZN(n15593) );
  AOI21_X1 U19016 ( .B1(n17186), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n15593), .ZN(n15594) );
  OAI21_X1 U19017 ( .B1(n15595), .B2(n20933), .A(n15594), .ZN(P1_U3021) );
  INV_X1 U19018 ( .A(n15596), .ZN(n15601) );
  INV_X1 U19019 ( .A(n20892), .ZN(n15597) );
  NOR2_X1 U19020 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15597), .ZN(
        n17201) );
  AND2_X1 U19021 ( .A1(n20915), .A2(n20892), .ZN(n15599) );
  OAI21_X1 U19022 ( .B1(n15600), .B2(n15599), .A(n15598), .ZN(n17205) );
  AOI21_X1 U19023 ( .B1(n15601), .B2(n17201), .A(n17205), .ZN(n17199) );
  OAI21_X1 U19024 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15602), .A(
        n17199), .ZN(n17192) );
  NAND2_X1 U19025 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15603) );
  OAI21_X1 U19026 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n15603), .ZN(n15607) );
  AOI21_X1 U19027 ( .B1(n15605), .B2(n17191), .A(n15604), .ZN(n15606) );
  OAI21_X1 U19028 ( .B1(n17196), .B2(n15607), .A(n15606), .ZN(n15608) );
  AOI21_X1 U19029 ( .B1(n17192), .B2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n15608), .ZN(n15609) );
  OAI21_X1 U19030 ( .B1(n15610), .B2(n20933), .A(n15609), .ZN(P1_U3023) );
  NAND2_X1 U19031 ( .A1(n15657), .A2(n15671), .ZN(n15627) );
  NAND2_X1 U19032 ( .A1(n15611), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n15612) );
  NAND2_X1 U19033 ( .A1(n11767), .A2(n15612), .ZN(n21289) );
  NAND2_X1 U19034 ( .A1(n15613), .A2(n21289), .ZN(n15624) );
  XNOR2_X1 U19035 ( .A(n15615), .B(n15614), .ZN(n15622) );
  INV_X1 U19036 ( .A(n15616), .ZN(n15620) );
  INV_X1 U19037 ( .A(n15617), .ZN(n15618) );
  XNOR2_X1 U19038 ( .A(n15618), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n15619) );
  NOR2_X1 U19039 ( .A1(n15620), .A2(n15619), .ZN(n15621) );
  AOI21_X1 U19040 ( .B1(n17084), .B2(n15622), .A(n15621), .ZN(n15623) );
  OAI21_X1 U19041 ( .B1(n15671), .B2(n15624), .A(n15623), .ZN(n15625) );
  INV_X1 U19042 ( .A(n15625), .ZN(n15626) );
  NAND2_X1 U19043 ( .A1(n15627), .A2(n15626), .ZN(n21292) );
  NAND2_X1 U19044 ( .A1(n21292), .A2(n15635), .ZN(n15629) );
  INV_X1 U19045 ( .A(n15635), .ZN(n17080) );
  NAND2_X1 U19046 ( .A1(n17080), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n15628) );
  NAND2_X1 U19047 ( .A1(n15629), .A2(n15628), .ZN(n17093) );
  NOR2_X1 U19048 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n17222), .ZN(n15636) );
  AOI22_X1 U19049 ( .A1(n17093), .A2(n17222), .B1(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n15636), .ZN(n15632) );
  MUX2_X1 U19050 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n15630), .S(
        n15635), .Z(n17090) );
  AOI22_X1 U19051 ( .A1(n15636), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n17222), .B2(n17090), .ZN(n15631) );
  NOR2_X1 U19052 ( .A1(n15632), .A2(n15631), .ZN(n17117) );
  INV_X1 U19053 ( .A(n17117), .ZN(n15639) );
  XNOR2_X1 U19054 ( .A(n15634), .B(n17214), .ZN(n20769) );
  OAI21_X1 U19055 ( .B1(n20769), .B2(n17210), .A(n15635), .ZN(n15638) );
  AOI21_X1 U19056 ( .B1(n17080), .B2(n17214), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n15637) );
  AOI22_X1 U19057 ( .A1(n15638), .A2(n15637), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n15636), .ZN(n17115) );
  OAI21_X1 U19058 ( .B1(n15639), .B2(n15666), .A(n17115), .ZN(n15645) );
  NOR2_X1 U19059 ( .A1(n15645), .A2(n17218), .ZN(n17130) );
  INV_X1 U19060 ( .A(n17130), .ZN(n15643) );
  NAND2_X1 U19061 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21064), .ZN(n15649) );
  AOI22_X1 U19062 ( .A1(n15641), .A2(n15649), .B1(n15640), .B2(n21149), .ZN(
        n15642) );
  NAND2_X1 U19063 ( .A1(n15643), .A2(n15642), .ZN(n15648) );
  OAI21_X1 U19064 ( .B1(n15645), .B2(P1_FLUSH_REG_SCAN_IN), .A(n15644), .ZN(
        n15647) );
  NAND2_X1 U19065 ( .A1(n15647), .A2(n15646), .ZN(n20941) );
  MUX2_X1 U19066 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n15648), .S(
        n20941), .Z(P1_U3478) );
  INV_X1 U19067 ( .A(n15649), .ZN(n15663) );
  OAI21_X1 U19068 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14014), .A(n21145), 
        .ZN(n15650) );
  OAI21_X1 U19069 ( .B1(n15663), .B2(n21060), .A(n15650), .ZN(n15651) );
  MUX2_X1 U19070 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15651), .S(
        n20941), .Z(P1_U3477) );
  INV_X1 U19071 ( .A(n15652), .ZN(n15655) );
  AOI21_X1 U19072 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14014), .A(n15653), 
        .ZN(n15654) );
  OAI22_X1 U19073 ( .A1(n15655), .A2(n15654), .B1(n13618), .B2(n15663), .ZN(
        n15656) );
  MUX2_X1 U19074 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n15656), .S(
        n20941), .Z(P1_U3476) );
  INV_X1 U19075 ( .A(n15657), .ZN(n15664) );
  MUX2_X1 U19076 ( .A(n21140), .B(n15659), .S(n14014), .Z(n15660) );
  NAND3_X1 U19077 ( .A1(n15660), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(n21031), 
        .ZN(n15661) );
  OAI211_X1 U19078 ( .C1(n10321), .C2(P1_STATEBS16_REG_SCAN_IN), .A(n15661), 
        .B(n21149), .ZN(n15662) );
  OAI21_X1 U19079 ( .B1(n15664), .B2(n15663), .A(n15662), .ZN(n15665) );
  MUX2_X1 U19080 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n15665), .S(
        n20941), .Z(P1_U3475) );
  INV_X1 U19081 ( .A(n15666), .ZN(n15668) );
  INV_X1 U19082 ( .A(n13624), .ZN(n15667) );
  NAND2_X1 U19083 ( .A1(n15668), .A2(n15667), .ZN(n15672) );
  OAI22_X1 U19084 ( .A1(n15669), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n15672), .B2(n12120), .ZN(n15670) );
  AOI21_X1 U19085 ( .B1(n21092), .B2(n15671), .A(n15670), .ZN(n17081) );
  INV_X1 U19086 ( .A(n15672), .ZN(n15676) );
  INV_X1 U19087 ( .A(n15673), .ZN(n15674) );
  AOI22_X1 U19088 ( .A1(n21290), .A2(n15676), .B1(n15675), .B2(n15674), .ZN(
        n15677) );
  OAI21_X1 U19089 ( .B1(n17081), .B2(n17211), .A(n15677), .ZN(n15678) );
  MUX2_X1 U19090 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15678), .S(
        n21294), .Z(P1_U3473) );
  OAI21_X1 U19091 ( .B1(n15723), .B2(n21197), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15680) );
  NAND2_X1 U19092 ( .A1(n15680), .A2(n21149), .ZN(n15690) );
  INV_X1 U19093 ( .A(n15690), .ZN(n15684) );
  NOR2_X1 U19094 ( .A1(n15681), .A2(n21092), .ZN(n15689) );
  INV_X1 U19095 ( .A(n21053), .ZN(n15685) );
  NAND2_X1 U19096 ( .A1(n15686), .A2(n15685), .ZN(n15720) );
  AOI22_X1 U19097 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15687), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n15720), .ZN(n15688) );
  NAND2_X1 U19098 ( .A1(n15719), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n15694) );
  OAI22_X1 U19099 ( .A1(n15691), .A2(n15720), .B1(n21070), .B2(n21190), .ZN(
        n15692) );
  AOI21_X1 U19100 ( .B1(n15723), .B2(n21055), .A(n15692), .ZN(n15693) );
  OAI211_X1 U19101 ( .C1(n15726), .C2(n15740), .A(n15694), .B(n15693), .ZN(
        P1_U3033) );
  NAND2_X1 U19102 ( .A1(n15719), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n15698) );
  OAI22_X1 U19103 ( .A1(n15695), .A2(n15720), .B1(n21159), .B2(n21190), .ZN(
        n15696) );
  AOI21_X1 U19104 ( .B1(n15723), .B2(n21156), .A(n15696), .ZN(n15697) );
  OAI211_X1 U19105 ( .C1(n15726), .C2(n15744), .A(n15698), .B(n15697), .ZN(
        P1_U3034) );
  NAND2_X1 U19106 ( .A1(n15719), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n15702) );
  OAI22_X1 U19107 ( .A1(n15699), .A2(n15720), .B1(n21165), .B2(n21190), .ZN(
        n15700) );
  AOI21_X1 U19108 ( .B1(n15723), .B2(n21162), .A(n15700), .ZN(n15701) );
  OAI211_X1 U19109 ( .C1(n15726), .C2(n15748), .A(n15702), .B(n15701), .ZN(
        P1_U3035) );
  NAND2_X1 U19110 ( .A1(n15719), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n15706) );
  OAI22_X1 U19111 ( .A1(n15703), .A2(n15720), .B1(n21171), .B2(n21190), .ZN(
        n15704) );
  AOI21_X1 U19112 ( .B1(n15723), .B2(n21168), .A(n15704), .ZN(n15705) );
  OAI211_X1 U19113 ( .C1(n15726), .C2(n15752), .A(n15706), .B(n15705), .ZN(
        P1_U3036) );
  NAND2_X1 U19114 ( .A1(n15719), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n15710) );
  OAI22_X1 U19115 ( .A1(n15707), .A2(n15720), .B1(n21177), .B2(n21190), .ZN(
        n15708) );
  AOI21_X1 U19116 ( .B1(n15723), .B2(n21174), .A(n15708), .ZN(n15709) );
  OAI211_X1 U19117 ( .C1(n15726), .C2(n15756), .A(n15710), .B(n15709), .ZN(
        P1_U3037) );
  NAND2_X1 U19118 ( .A1(n15719), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n15714) );
  OAI22_X1 U19119 ( .A1(n15711), .A2(n15720), .B1(n21183), .B2(n21190), .ZN(
        n15712) );
  AOI21_X1 U19120 ( .B1(n15723), .B2(n21180), .A(n15712), .ZN(n15713) );
  OAI211_X1 U19121 ( .C1(n15726), .C2(n15760), .A(n15714), .B(n15713), .ZN(
        P1_U3038) );
  NAND2_X1 U19122 ( .A1(n15719), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n15718) );
  OAI22_X1 U19123 ( .A1(n15715), .A2(n15720), .B1(n21084), .B2(n21190), .ZN(
        n15716) );
  AOI21_X1 U19124 ( .B1(n15723), .B2(n21081), .A(n15716), .ZN(n15717) );
  OAI211_X1 U19125 ( .C1(n15726), .C2(n15764), .A(n15718), .B(n15717), .ZN(
        P1_U3039) );
  NAND2_X1 U19126 ( .A1(n15719), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n15725) );
  OAI22_X1 U19127 ( .A1(n15721), .A2(n15720), .B1(n21202), .B2(n21190), .ZN(
        n15722) );
  AOI21_X1 U19128 ( .B1(n15723), .B2(n21196), .A(n15722), .ZN(n15724) );
  OAI211_X1 U19129 ( .C1(n15726), .C2(n15772), .A(n15725), .B(n15724), .ZN(
        P1_U3040) );
  NAND2_X1 U19130 ( .A1(n15768), .A2(n21029), .ZN(n15727) );
  OAI21_X1 U19131 ( .B1(n15770), .B2(n15727), .A(n21057), .ZN(n15735) );
  AND2_X1 U19132 ( .A1(n15728), .A2(n21092), .ZN(n15732) );
  NOR2_X1 U19133 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15731), .ZN(
        n15766) );
  INV_X1 U19134 ( .A(n15732), .ZN(n15734) );
  AOI21_X1 U19135 ( .B1(n15735), .B2(n15734), .A(n15733), .ZN(n15736) );
  AOI22_X1 U19136 ( .A1(n21138), .A2(n15766), .B1(
        P1_INSTQUEUE_REG_6__0__SCAN_IN), .B2(n15765), .ZN(n15737) );
  OAI21_X1 U19137 ( .B1(n21153), .B2(n15768), .A(n15737), .ZN(n15738) );
  AOI21_X1 U19138 ( .B1(n15770), .B2(n21150), .A(n15738), .ZN(n15739) );
  OAI21_X1 U19139 ( .B1(n15773), .B2(n15740), .A(n15739), .ZN(P1_U3081) );
  AOI22_X1 U19140 ( .A1(n21154), .A2(n15766), .B1(
        P1_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n15765), .ZN(n15741) );
  OAI21_X1 U19141 ( .B1(n21105), .B2(n15768), .A(n15741), .ZN(n15742) );
  AOI21_X1 U19142 ( .B1(n15770), .B2(n21102), .A(n15742), .ZN(n15743) );
  OAI21_X1 U19143 ( .B1(n15773), .B2(n15744), .A(n15743), .ZN(P1_U3082) );
  AOI22_X1 U19144 ( .A1(n21160), .A2(n15766), .B1(
        P1_INSTQUEUE_REG_6__2__SCAN_IN), .B2(n15765), .ZN(n15745) );
  OAI21_X1 U19145 ( .B1(n21109), .B2(n15768), .A(n15745), .ZN(n15746) );
  AOI21_X1 U19146 ( .B1(n15770), .B2(n21106), .A(n15746), .ZN(n15747) );
  OAI21_X1 U19147 ( .B1(n15773), .B2(n15748), .A(n15747), .ZN(P1_U3083) );
  AOI22_X1 U19148 ( .A1(n21166), .A2(n15766), .B1(
        P1_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n15765), .ZN(n15749) );
  OAI21_X1 U19149 ( .B1(n21113), .B2(n15768), .A(n15749), .ZN(n15750) );
  AOI21_X1 U19150 ( .B1(n15770), .B2(n21110), .A(n15750), .ZN(n15751) );
  OAI21_X1 U19151 ( .B1(n15773), .B2(n15752), .A(n15751), .ZN(P1_U3084) );
  AOI22_X1 U19152 ( .A1(n21172), .A2(n15766), .B1(
        P1_INSTQUEUE_REG_6__4__SCAN_IN), .B2(n15765), .ZN(n15753) );
  OAI21_X1 U19153 ( .B1(n21117), .B2(n15768), .A(n15753), .ZN(n15754) );
  AOI21_X1 U19154 ( .B1(n15770), .B2(n21114), .A(n15754), .ZN(n15755) );
  OAI21_X1 U19155 ( .B1(n15773), .B2(n15756), .A(n15755), .ZN(P1_U3085) );
  AOI22_X1 U19156 ( .A1(n21178), .A2(n15766), .B1(
        P1_INSTQUEUE_REG_6__5__SCAN_IN), .B2(n15765), .ZN(n15757) );
  OAI21_X1 U19157 ( .B1(n21121), .B2(n15768), .A(n15757), .ZN(n15758) );
  AOI21_X1 U19158 ( .B1(n15770), .B2(n21118), .A(n15758), .ZN(n15759) );
  OAI21_X1 U19159 ( .B1(n15773), .B2(n15760), .A(n15759), .ZN(P1_U3086) );
  AOI22_X1 U19160 ( .A1(n21184), .A2(n15766), .B1(
        P1_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n15765), .ZN(n15761) );
  OAI21_X1 U19161 ( .B1(n21191), .B2(n15768), .A(n15761), .ZN(n15762) );
  AOI21_X1 U19162 ( .B1(n15770), .B2(n21186), .A(n15762), .ZN(n15763) );
  OAI21_X1 U19163 ( .B1(n15773), .B2(n15764), .A(n15763), .ZN(P1_U3087) );
  AOI22_X1 U19164 ( .A1(n21193), .A2(n15766), .B1(
        P1_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n15765), .ZN(n15767) );
  OAI21_X1 U19165 ( .B1(n21131), .B2(n15768), .A(n15767), .ZN(n15769) );
  AOI21_X1 U19166 ( .B1(n15770), .B2(n21126), .A(n15769), .ZN(n15771) );
  OAI21_X1 U19167 ( .B1(n15773), .B2(n15772), .A(n15771), .ZN(P1_U3088) );
  AOI21_X1 U19168 ( .B1(n15776), .B2(n15775), .A(n15774), .ZN(n15777) );
  AND2_X1 U19169 ( .A1(n15779), .A2(n15778), .ZN(n15780) );
  NOR2_X1 U19170 ( .A1(n15781), .A2(n15780), .ZN(n16559) );
  AOI22_X1 U19171 ( .A1(n19834), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19864), .ZN(n15785) );
  NAND2_X1 U19172 ( .A1(n19856), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15784) );
  NAND2_X1 U19173 ( .A1(n16303), .A2(n19768), .ZN(n15797) );
  AOI21_X1 U19174 ( .B1(n15789), .B2(n19875), .A(n16043), .ZN(n15793) );
  INV_X1 U19175 ( .A(n19834), .ZN(n19859) );
  OAI22_X1 U19176 ( .A1(n19859), .A2(n15787), .B1(n15786), .B2(n19838), .ZN(
        n15791) );
  INV_X1 U19177 ( .A(n16307), .ZN(n15788) );
  NOR3_X1 U19178 ( .A1(n15789), .A2(n15788), .A3(n16046), .ZN(n15790) );
  AOI211_X1 U19179 ( .C1(n19856), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15791), .B(n15790), .ZN(n15792) );
  OAI21_X1 U19180 ( .B1(n15793), .B2(n16307), .A(n15792), .ZN(n15794) );
  AOI21_X1 U19181 ( .B1(n15795), .B2(n19832), .A(n15794), .ZN(n15796) );
  OAI211_X1 U19182 ( .C1(n19870), .C2(n16166), .A(n15797), .B(n15796), .ZN(
        P2_U2827) );
  AND2_X1 U19183 ( .A1(n15798), .A2(n15810), .ZN(n15812) );
  OAI21_X1 U19184 ( .B1(n15812), .B2(n15799), .A(n14322), .ZN(n16572) );
  OAI21_X1 U19185 ( .B1(n15800), .B2(n15801), .A(n14326), .ZN(n16320) );
  INV_X1 U19186 ( .A(n16320), .ZN(n16574) );
  NAND2_X1 U19187 ( .A1(n16574), .A2(n19768), .ZN(n15809) );
  XOR2_X1 U19188 ( .A(n16323), .B(n15802), .Z(n15807) );
  AOI22_X1 U19189 ( .A1(n19834), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_EBX_REG_27__SCAN_IN), .B2(n19864), .ZN(n15803) );
  OAI21_X1 U19190 ( .B1(n19878), .B2(n16319), .A(n15803), .ZN(n15806) );
  NOR2_X1 U19191 ( .A1(n15804), .A2(n19860), .ZN(n15805) );
  AOI211_X1 U19192 ( .C1(n19875), .C2(n15807), .A(n15806), .B(n15805), .ZN(
        n15808) );
  OAI211_X1 U19193 ( .C1(n19870), .C2(n16572), .A(n15809), .B(n15808), .ZN(
        P2_U2828) );
  NOR2_X1 U19194 ( .A1(n15798), .A2(n15810), .ZN(n15811) );
  AOI21_X1 U19195 ( .B1(n15814), .B2(n15813), .A(n15800), .ZN(n16585) );
  NAND2_X1 U19196 ( .A1(n16585), .A2(n19768), .ZN(n15823) );
  AOI21_X1 U19197 ( .B1(n9641), .B2(n19875), .A(n16043), .ZN(n15819) );
  OAI22_X1 U19198 ( .A1(n19859), .A2(n20607), .B1(n15815), .B2(n19838), .ZN(
        n15817) );
  NOR3_X1 U19199 ( .A1(n9641), .A2(n10250), .A3(n16046), .ZN(n15816) );
  AOI211_X1 U19200 ( .C1(n19856), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15817), .B(n15816), .ZN(n15818) );
  OAI21_X1 U19201 ( .B1(n15819), .B2(n16331), .A(n15818), .ZN(n15820) );
  AOI21_X1 U19202 ( .B1(n15821), .B2(n19832), .A(n15820), .ZN(n15822) );
  OAI211_X1 U19203 ( .C1(n19870), .C2(n16583), .A(n15823), .B(n15822), .ZN(
        P2_U2829) );
  NAND2_X1 U19204 ( .A1(n15824), .A2(n15825), .ZN(n15826) );
  NAND2_X1 U19205 ( .A1(n15813), .A2(n15826), .ZN(n16591) );
  XNOR2_X1 U19206 ( .A(n15827), .B(P2_EBX_REG_25__SCAN_IN), .ZN(n15834) );
  XNOR2_X1 U19207 ( .A(n15828), .B(n16341), .ZN(n15832) );
  OAI22_X1 U19208 ( .A1(n19859), .A2(n20605), .B1(n15829), .B2(n19838), .ZN(
        n15830) );
  AOI21_X1 U19209 ( .B1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19856), .A(
        n15830), .ZN(n15831) );
  OAI21_X1 U19210 ( .B1(n15832), .B2(n20545), .A(n15831), .ZN(n15833) );
  AOI21_X1 U19211 ( .B1(n15834), .B2(n19832), .A(n15833), .ZN(n15837) );
  XOR2_X1 U19212 ( .A(n15835), .B(n9637), .Z(n16594) );
  NAND2_X1 U19213 ( .A1(n16594), .A2(n19803), .ZN(n15836) );
  OAI211_X1 U19214 ( .C1(n16591), .C2(n19871), .A(n15837), .B(n15836), .ZN(
        P2_U2830) );
  NAND2_X1 U19215 ( .A1(n15838), .A2(n15839), .ZN(n15840) );
  NAND2_X1 U19216 ( .A1(n9637), .A2(n15840), .ZN(n16605) );
  OAI21_X1 U19217 ( .B1(n15841), .B2(n15842), .A(n15824), .ZN(n16085) );
  INV_X1 U19218 ( .A(n16085), .ZN(n16607) );
  NAND2_X1 U19219 ( .A1(n16607), .A2(n19768), .ZN(n15853) );
  AOI21_X1 U19220 ( .B1(n15844), .B2(n19875), .A(n16043), .ZN(n15843) );
  NOR2_X1 U19221 ( .A1(n15843), .A2(n16350), .ZN(n15850) );
  INV_X1 U19222 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15848) );
  INV_X1 U19223 ( .A(n15844), .ZN(n15845) );
  NAND3_X1 U19224 ( .A1(n15845), .A2(n19810), .A3(n16350), .ZN(n15847) );
  AOI22_X1 U19225 ( .A1(n19834), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_EBX_REG_24__SCAN_IN), .B2(n19864), .ZN(n15846) );
  OAI211_X1 U19226 ( .C1(n19878), .C2(n15848), .A(n15847), .B(n15846), .ZN(
        n15849) );
  AOI211_X1 U19227 ( .C1(n15851), .C2(n19832), .A(n15850), .B(n15849), .ZN(
        n15852) );
  OAI211_X1 U19228 ( .C1(n19870), .C2(n16605), .A(n15853), .B(n15852), .ZN(
        P2_U2831) );
  INV_X1 U19229 ( .A(n15841), .ZN(n15855) );
  OAI21_X1 U19230 ( .B1(n15854), .B2(n15856), .A(n15855), .ZN(n16611) );
  XNOR2_X1 U19231 ( .A(n15857), .B(n16356), .ZN(n15860) );
  INV_X1 U19232 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n21449) );
  OAI22_X1 U19233 ( .A1(n19859), .A2(n20601), .B1(n21449), .B2(n19838), .ZN(
        n15858) );
  AOI21_X1 U19234 ( .B1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19856), .A(
        n15858), .ZN(n15859) );
  OAI21_X1 U19235 ( .B1(n20545), .B2(n15860), .A(n15859), .ZN(n15864) );
  OAI21_X1 U19236 ( .B1(n15861), .B2(n15862), .A(n15838), .ZN(n16612) );
  NOR2_X1 U19237 ( .A1(n16612), .A2(n19870), .ZN(n15863) );
  AOI211_X1 U19238 ( .C1(n19832), .C2(n15865), .A(n15864), .B(n15863), .ZN(
        n15866) );
  OAI21_X1 U19239 ( .B1(n16611), .B2(n19871), .A(n15866), .ZN(P2_U2832) );
  AND2_X1 U19240 ( .A1(n15884), .A2(n15869), .ZN(n15870) );
  OR2_X1 U19241 ( .A1(n15870), .A2(n15854), .ZN(n16370) );
  CLKBUF_X1 U19242 ( .A(n15871), .Z(n15872) );
  AOI21_X1 U19243 ( .B1(n15873), .B2(n15872), .A(n15861), .ZN(n16624) );
  OAI21_X1 U19244 ( .B1(n15874), .B2(n20545), .A(n19806), .ZN(n15878) );
  AOI22_X1 U19245 ( .A1(n19834), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_EBX_REG_22__SCAN_IN), .B2(n19864), .ZN(n15876) );
  INV_X1 U19246 ( .A(n15879), .ZN(n16373) );
  NAND3_X1 U19247 ( .A1(n15874), .A2(n19810), .A3(n16373), .ZN(n15875) );
  OAI211_X1 U19248 ( .C1(n19878), .C2(n10400), .A(n15876), .B(n15875), .ZN(
        n15877) );
  AOI21_X1 U19249 ( .B1(n15879), .B2(n15878), .A(n15877), .ZN(n15880) );
  OAI21_X1 U19250 ( .B1(n15881), .B2(n19860), .A(n15880), .ZN(n15882) );
  AOI21_X1 U19251 ( .B1(n16624), .B2(n19803), .A(n15882), .ZN(n15883) );
  OAI21_X1 U19252 ( .B1(n16370), .B2(n19871), .A(n15883), .ZN(P2_U2833) );
  OAI21_X1 U19253 ( .B1(n11457), .B2(n9753), .A(n15872), .ZN(n16642) );
  AOI21_X1 U19254 ( .B1(n15885), .B2(n14399), .A(n15868), .ZN(n16645) );
  NAND2_X1 U19255 ( .A1(n16645), .A2(n19768), .ZN(n15895) );
  INV_X1 U19256 ( .A(n15886), .ZN(n15887) );
  AOI221_X1 U19257 ( .B1(n10384), .B2(n15887), .C1(n16384), .C2(n15886), .A(
        n20545), .ZN(n15888) );
  AOI21_X1 U19258 ( .B1(n19834), .B2(P2_REIP_REG_21__SCAN_IN), .A(n15888), 
        .ZN(n15889) );
  OAI21_X1 U19259 ( .B1(n15890), .B2(n19838), .A(n15889), .ZN(n15893) );
  NOR2_X1 U19260 ( .A1(n15891), .A2(n19860), .ZN(n15892) );
  AOI211_X1 U19261 ( .C1(n19856), .C2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15893), .B(n15892), .ZN(n15894) );
  OAI211_X1 U19262 ( .C1(n19870), .C2(n16642), .A(n15895), .B(n15894), .ZN(
        P2_U2834) );
  INV_X1 U19263 ( .A(n16232), .ZN(n15904) );
  XNOR2_X1 U19264 ( .A(n9661), .B(P2_EBX_REG_20__SCAN_IN), .ZN(n15902) );
  AOI211_X1 U19265 ( .C1(n10234), .C2(n15897), .A(n20545), .B(n15886), .ZN(
        n15900) );
  AOI22_X1 U19266 ( .A1(n19834), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_EBX_REG_20__SCAN_IN), .B2(n19864), .ZN(n15898) );
  OAI21_X1 U19267 ( .B1(n10399), .B2(n19878), .A(n15898), .ZN(n15899) );
  AOI211_X1 U19268 ( .C1(n16043), .C2(n10234), .A(n15900), .B(n15899), .ZN(
        n15901) );
  OAI21_X1 U19269 ( .B1(n15902), .B2(n19860), .A(n15901), .ZN(n15903) );
  AOI21_X1 U19270 ( .B1(n15904), .B2(n19803), .A(n15903), .ZN(n15905) );
  OAI21_X1 U19271 ( .B1(n16107), .B2(n19871), .A(n15905), .ZN(P2_U2835) );
  NOR2_X1 U19272 ( .A1(n19806), .A2(n15910), .ZN(n15909) );
  NAND2_X1 U19273 ( .A1(n19834), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15906) );
  OAI211_X1 U19274 ( .C1(n19838), .C2(n15907), .A(n15906), .B(n16491), .ZN(
        n15908) );
  AOI211_X1 U19275 ( .C1(n19856), .C2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15909), .B(n15908), .ZN(n15913) );
  OAI211_X1 U19276 ( .C1(n15911), .C2(n15910), .A(n19810), .B(n19745), .ZN(
        n15912) );
  OAI211_X1 U19277 ( .C1(n15914), .C2(n19860), .A(n15913), .B(n15912), .ZN(
        n15915) );
  AOI21_X1 U19278 ( .B1(n16248), .B2(n19803), .A(n15915), .ZN(n15916) );
  OAI21_X1 U19279 ( .B1(n16123), .B2(n19871), .A(n15916), .ZN(P2_U2838) );
  NAND2_X1 U19280 ( .A1(n16682), .A2(n19768), .ZN(n15927) );
  NAND2_X1 U19281 ( .A1(n19866), .A2(n15917), .ZN(n15918) );
  XOR2_X1 U19282 ( .A(n16421), .B(n15918), .Z(n15925) );
  AOI21_X1 U19283 ( .B1(n19834), .B2(P2_REIP_REG_14__SCAN_IN), .A(n19941), 
        .ZN(n15920) );
  NAND2_X1 U19284 ( .A1(n19864), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15919) );
  OAI211_X1 U19285 ( .C1(n19878), .C2(n15921), .A(n15920), .B(n15919), .ZN(
        n15924) );
  NOR2_X1 U19286 ( .A1(n15922), .A2(n19860), .ZN(n15923) );
  AOI211_X1 U19287 ( .C1(n19875), .C2(n15925), .A(n15924), .B(n15923), .ZN(
        n15926) );
  OAI211_X1 U19288 ( .C1(n19870), .C2(n16689), .A(n15927), .B(n15926), .ZN(
        P2_U2841) );
  NAND2_X1 U19289 ( .A1(n16695), .A2(n19768), .ZN(n15939) );
  INV_X1 U19290 ( .A(n15928), .ZN(n15937) );
  AOI21_X1 U19291 ( .B1(n19875), .B2(n15930), .A(n16043), .ZN(n15935) );
  AOI21_X1 U19292 ( .B1(n19834), .B2(P2_REIP_REG_13__SCAN_IN), .A(n19941), 
        .ZN(n15929) );
  OAI21_X1 U19293 ( .B1(n10718), .B2(n19838), .A(n15929), .ZN(n15933) );
  INV_X1 U19294 ( .A(n16429), .ZN(n15931) );
  NOR3_X1 U19295 ( .A1(n16046), .A2(n15931), .A3(n15930), .ZN(n15932) );
  AOI211_X1 U19296 ( .C1(n19856), .C2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15933), .B(n15932), .ZN(n15934) );
  OAI21_X1 U19297 ( .B1(n15935), .B2(n16429), .A(n15934), .ZN(n15936) );
  AOI21_X1 U19298 ( .B1(n15937), .B2(n19832), .A(n15936), .ZN(n15938) );
  OAI211_X1 U19299 ( .C1(n16699), .C2(n19870), .A(n15939), .B(n15938), .ZN(
        P2_U2842) );
  INV_X1 U19300 ( .A(n16705), .ZN(n15950) );
  OAI21_X1 U19301 ( .B1(n20545), .B2(n19809), .A(n19806), .ZN(n15945) );
  AND3_X1 U19302 ( .A1(n19810), .A2(n16442), .A3(n19809), .ZN(n15944) );
  INV_X1 U19303 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15942) );
  AOI21_X1 U19304 ( .B1(n19834), .B2(P2_REIP_REG_12__SCAN_IN), .A(n19941), 
        .ZN(n15941) );
  NAND2_X1 U19305 ( .A1(n19864), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n15940) );
  OAI211_X1 U19306 ( .C1(n19878), .C2(n15942), .A(n15941), .B(n15940), .ZN(
        n15943) );
  AOI211_X1 U19307 ( .C1(n15946), .C2(n15945), .A(n15944), .B(n15943), .ZN(
        n15947) );
  OAI21_X1 U19308 ( .B1(n15948), .B2(n19860), .A(n15947), .ZN(n15949) );
  AOI21_X1 U19309 ( .B1(n15950), .B2(n19803), .A(n15949), .ZN(n15951) );
  OAI21_X1 U19310 ( .B1(n16710), .B2(n19871), .A(n15951), .ZN(P2_U2843) );
  OAI21_X1 U19311 ( .B1(n15952), .B2(n20545), .A(n19806), .ZN(n15958) );
  INV_X1 U19312 ( .A(n15952), .ZN(n15953) );
  NOR3_X1 U19313 ( .A1(n16046), .A2(n16489), .A3(n15953), .ZN(n15957) );
  AOI21_X1 U19314 ( .B1(n19834), .B2(P2_REIP_REG_8__SCAN_IN), .A(n19941), .ZN(
        n15955) );
  NAND2_X1 U19315 ( .A1(n19864), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n15954) );
  OAI211_X1 U19316 ( .C1(n19878), .C2(n16493), .A(n15955), .B(n15954), .ZN(
        n15956) );
  AOI211_X1 U19317 ( .C1(n16489), .C2(n15958), .A(n15957), .B(n15956), .ZN(
        n15959) );
  OAI21_X1 U19318 ( .B1(n15960), .B2(n19860), .A(n15959), .ZN(n15961) );
  AOI21_X1 U19319 ( .B1(n16754), .B2(n19803), .A(n15961), .ZN(n15962) );
  OAI21_X1 U19320 ( .B1(n16756), .B2(n19871), .A(n15962), .ZN(P2_U2847) );
  OR2_X1 U19321 ( .A1(n15965), .A2(n15964), .ZN(n15966) );
  NAND2_X1 U19322 ( .A1(n15963), .A2(n15966), .ZN(n16797) );
  INV_X1 U19323 ( .A(n16797), .ZN(n15978) );
  INV_X1 U19324 ( .A(n16530), .ZN(n15974) );
  INV_X1 U19325 ( .A(n15968), .ZN(n15967) );
  OAI21_X1 U19326 ( .B1(n20545), .B2(n15967), .A(n19806), .ZN(n15973) );
  NOR3_X1 U19327 ( .A1(n16046), .A2(n15968), .A3(n15974), .ZN(n15972) );
  INV_X1 U19328 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16531) );
  AOI21_X1 U19329 ( .B1(n19834), .B2(P2_REIP_REG_5__SCAN_IN), .A(n19941), .ZN(
        n15970) );
  NAND2_X1 U19330 ( .A1(n19864), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n15969) );
  OAI211_X1 U19331 ( .C1(n19878), .C2(n16531), .A(n15970), .B(n15969), .ZN(
        n15971) );
  AOI211_X1 U19332 ( .C1(n15974), .C2(n15973), .A(n15972), .B(n15971), .ZN(
        n15975) );
  OAI21_X1 U19333 ( .B1(n15976), .B2(n19860), .A(n15975), .ZN(n15977) );
  AOI21_X1 U19334 ( .B1(n15978), .B2(n19803), .A(n15977), .ZN(n15979) );
  OAI21_X1 U19335 ( .B1(n15980), .B2(n19871), .A(n15979), .ZN(P2_U2850) );
  INV_X1 U19336 ( .A(n16277), .ZN(n15995) );
  INV_X1 U19337 ( .A(n19949), .ZN(n16814) );
  XNOR2_X1 U19338 ( .A(n15981), .B(n15982), .ZN(n16809) );
  AND2_X1 U19339 ( .A1(n19866), .A2(n15983), .ZN(n15985) );
  AOI21_X1 U19340 ( .B1(n19942), .B2(n15985), .A(n20545), .ZN(n15984) );
  OAI21_X1 U19341 ( .B1(n15985), .B2(n19942), .A(n15984), .ZN(n15986) );
  INV_X1 U19342 ( .A(n15986), .ZN(n15990) );
  AOI21_X1 U19343 ( .B1(n19834), .B2(P2_REIP_REG_4__SCAN_IN), .A(n19941), .ZN(
        n15988) );
  NAND2_X1 U19344 ( .A1(n19864), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n15987) );
  OAI211_X1 U19345 ( .C1(n19878), .C2(n19954), .A(n15988), .B(n15987), .ZN(
        n15989) );
  AOI211_X1 U19346 ( .C1(n19832), .C2(n15991), .A(n15990), .B(n15989), .ZN(
        n15992) );
  OAI21_X1 U19347 ( .B1(n16809), .B2(n19870), .A(n15992), .ZN(n15993) );
  AOI21_X1 U19348 ( .B1(n16814), .B2(n19768), .A(n15993), .ZN(n15994) );
  OAI21_X1 U19349 ( .B1(n15995), .B2(n19716), .A(n15994), .ZN(P2_U2851) );
  NAND2_X1 U19350 ( .A1(n15997), .A2(n15996), .ZN(n15998) );
  NAND2_X1 U19351 ( .A1(n15981), .A2(n15998), .ZN(n17226) );
  INV_X1 U19352 ( .A(n17226), .ZN(n20635) );
  INV_X1 U19353 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n20571) );
  AOI22_X1 U19354 ( .A1(n19834), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_EBX_REG_3__SCAN_IN), .B2(n19864), .ZN(n16001) );
  NAND3_X1 U19355 ( .A1(n19810), .A2(n16543), .A3(n15999), .ZN(n16000) );
  OAI211_X1 U19356 ( .C1(n19878), .C2(n10396), .A(n16001), .B(n16000), .ZN(
        n16006) );
  AOI21_X1 U19357 ( .B1(n19875), .B2(n16002), .A(n16043), .ZN(n16004) );
  OAI22_X1 U19358 ( .A1(n16004), .A2(n16543), .B1(n16003), .B2(n19860), .ZN(
        n16005) );
  AOI211_X1 U19359 ( .C1(n20635), .C2(n19803), .A(n16006), .B(n16005), .ZN(
        n16010) );
  NAND2_X1 U19360 ( .A1(n16008), .A2(n19768), .ZN(n16009) );
  OAI211_X1 U19361 ( .C1(n16864), .C2(n19716), .A(n16010), .B(n16009), .ZN(
        P2_U2852) );
  INV_X1 U19362 ( .A(n20645), .ZN(n16020) );
  OAI21_X1 U19363 ( .B1(n20545), .B2(n16027), .A(n19806), .ZN(n16015) );
  AOI22_X1 U19364 ( .A1(n19834), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_EBX_REG_2__SCAN_IN), .B2(n19864), .ZN(n16012) );
  NAND3_X1 U19365 ( .A1(n19810), .A2(n16027), .A3(n10237), .ZN(n16011) );
  OAI211_X1 U19366 ( .C1(n19878), .C2(n16013), .A(n16012), .B(n16011), .ZN(
        n16014) );
  AOI21_X1 U19367 ( .B1(n16016), .B2(n16015), .A(n16014), .ZN(n16019) );
  NAND2_X1 U19368 ( .A1(n19832), .A2(n16017), .ZN(n16018) );
  OAI211_X1 U19369 ( .C1(n16020), .C2(n19870), .A(n16019), .B(n16018), .ZN(
        n16021) );
  AOI21_X1 U19370 ( .B1(n13766), .B2(n19768), .A(n16021), .ZN(n16022) );
  OAI21_X1 U19371 ( .B1(n16848), .B2(n19716), .A(n16022), .ZN(P2_U2853) );
  OR2_X1 U19372 ( .A1(n16024), .A2(n16023), .ZN(n16026) );
  NAND2_X1 U19373 ( .A1(n16026), .A2(n16025), .ZN(n20653) );
  NOR2_X1 U19374 ( .A1(n19806), .A2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16036) );
  OAI21_X1 U19375 ( .B1(n16028), .B2(n16823), .A(n16027), .ZN(n16029) );
  INV_X1 U19376 ( .A(n16029), .ZN(n16030) );
  NAND2_X1 U19377 ( .A1(n19866), .A2(n16030), .ZN(n16828) );
  NOR2_X1 U19378 ( .A1(n19838), .A2(n10819), .ZN(n16033) );
  OAI22_X1 U19379 ( .A1(n19859), .A2(n20567), .B1(n16031), .B2(n19860), .ZN(
        n16032) );
  AOI211_X1 U19380 ( .C1(n19856), .C2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n16033), .B(n16032), .ZN(n16034) );
  OAI21_X1 U19381 ( .B1(n20545), .B2(n16828), .A(n16034), .ZN(n16035) );
  AOI211_X1 U19382 ( .C1(n19803), .C2(n20653), .A(n16036), .B(n16035), .ZN(
        n16038) );
  NAND2_X1 U19383 ( .A1(n9927), .A2(n19768), .ZN(n16037) );
  OAI211_X1 U19384 ( .C1(n20655), .C2(n19716), .A(n16038), .B(n16037), .ZN(
        P2_U2854) );
  AOI22_X1 U19385 ( .A1(n19834), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n19803), 
        .B2(n17235), .ZN(n16039) );
  OAI21_X1 U19386 ( .B1(n16040), .B2(n19838), .A(n16039), .ZN(n16041) );
  AOI21_X1 U19387 ( .B1(n19832), .B2(n16042), .A(n16041), .ZN(n16045) );
  OAI21_X1 U19388 ( .B1(n19856), .B2(n16043), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16044) );
  OAI211_X1 U19389 ( .C1(n16823), .C2(n16046), .A(n16045), .B(n16044), .ZN(
        n16047) );
  AOI21_X1 U19390 ( .B1(n13581), .B2(n19768), .A(n16047), .ZN(n16048) );
  OAI21_X1 U19391 ( .B1(n16907), .B2(n19716), .A(n16048), .ZN(P2_U2855) );
  OR2_X1 U19392 ( .A1(n16050), .A2(n16049), .ZN(n16158) );
  NAND3_X1 U19393 ( .A1(n16158), .A2(n16051), .A3(n16150), .ZN(n16053) );
  NAND2_X1 U19394 ( .A1(n16157), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16052) );
  OAI211_X1 U19395 ( .C1(n16562), .C2(n16154), .A(n16053), .B(n16052), .ZN(
        P2_U2858) );
  NOR2_X1 U19396 ( .A1(n16055), .A2(n16054), .ZN(n16057) );
  XNOR2_X1 U19397 ( .A(n16057), .B(n16056), .ZN(n16174) );
  NAND2_X1 U19398 ( .A1(n16154), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n16059) );
  NAND2_X1 U19399 ( .A1(n16303), .A2(n16104), .ZN(n16058) );
  OAI211_X1 U19400 ( .C1(n16174), .C2(n9716), .A(n16059), .B(n16058), .ZN(
        P2_U2859) );
  OAI21_X1 U19401 ( .B1(n16060), .B2(n16062), .A(n16061), .ZN(n16180) );
  NOR2_X1 U19402 ( .A1(n16320), .A2(n16157), .ZN(n16063) );
  AOI21_X1 U19403 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n16157), .A(n16063), .ZN(
        n16064) );
  OAI21_X1 U19404 ( .B1(n16180), .B2(n9716), .A(n16064), .ZN(P2_U2860) );
  NOR2_X1 U19405 ( .A1(n16075), .A2(n16074), .ZN(n16073) );
  NOR2_X1 U19406 ( .A1(n16073), .A2(n16065), .ZN(n16070) );
  NOR2_X1 U19407 ( .A1(n19972), .A2(n16066), .ZN(n16067) );
  XNOR2_X1 U19408 ( .A(n16068), .B(n16067), .ZN(n16069) );
  XNOR2_X1 U19409 ( .A(n16070), .B(n16069), .ZN(n16188) );
  NAND2_X1 U19410 ( .A1(n16585), .A2(n16104), .ZN(n16072) );
  NAND2_X1 U19411 ( .A1(n16154), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n16071) );
  OAI211_X1 U19412 ( .C1(n16188), .C2(n9716), .A(n16072), .B(n16071), .ZN(
        P2_U2861) );
  AOI21_X1 U19413 ( .B1(n16075), .B2(n16074), .A(n16073), .ZN(n16189) );
  NAND2_X1 U19414 ( .A1(n16189), .A2(n16150), .ZN(n16077) );
  NAND2_X1 U19415 ( .A1(n16157), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n16076) );
  OAI211_X1 U19416 ( .C1(n16591), .C2(n16157), .A(n16077), .B(n16076), .ZN(
        P2_U2862) );
  XOR2_X1 U19417 ( .A(n16080), .B(n16078), .Z(n16090) );
  NOR2_X1 U19418 ( .A1(n19972), .A2(n16079), .ZN(n16089) );
  NAND2_X1 U19419 ( .A1(n16090), .A2(n16089), .ZN(n16088) );
  OAI21_X1 U19420 ( .B1(n16080), .B2(n16078), .A(n16088), .ZN(n16084) );
  XOR2_X1 U19421 ( .A(n16082), .B(n16081), .Z(n16083) );
  XNOR2_X1 U19422 ( .A(n16084), .B(n16083), .ZN(n16205) );
  NOR2_X1 U19423 ( .A1(n16085), .A2(n16157), .ZN(n16086) );
  AOI21_X1 U19424 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n16157), .A(n16086), .ZN(
        n16087) );
  OAI21_X1 U19425 ( .B1(n16205), .B2(n9716), .A(n16087), .ZN(P2_U2863) );
  OAI21_X1 U19426 ( .B1(n16090), .B2(n16089), .A(n16088), .ZN(n16211) );
  NOR2_X1 U19427 ( .A1(n16611), .A2(n16157), .ZN(n16091) );
  AOI21_X1 U19428 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n16157), .A(n16091), .ZN(
        n16092) );
  OAI21_X1 U19429 ( .B1(n9716), .B2(n16211), .A(n16092), .ZN(P2_U2864) );
  NAND2_X1 U19430 ( .A1(n16093), .A2(n16098), .ZN(n16097) );
  INV_X1 U19431 ( .A(n16078), .ZN(n16094) );
  AOI21_X1 U19432 ( .B1(n16095), .B2(n16097), .A(n16094), .ZN(n16216) );
  AOI22_X1 U19433 ( .A1(n16216), .A2(n16150), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n16154), .ZN(n16096) );
  OAI21_X1 U19434 ( .B1(n16370), .B2(n16154), .A(n16096), .ZN(P2_U2865) );
  INV_X1 U19435 ( .A(n16645), .ZN(n16101) );
  OAI21_X1 U19436 ( .B1(n16093), .B2(n16098), .A(n16097), .ZN(n16099) );
  INV_X1 U19437 ( .A(n16099), .ZN(n16223) );
  AOI22_X1 U19438 ( .A1(n16223), .A2(n16150), .B1(P2_EBX_REG_21__SCAN_IN), 
        .B2(n16157), .ZN(n16100) );
  OAI21_X1 U19439 ( .B1(n16101), .B2(n16157), .A(n16100), .ZN(P2_U2866) );
  NOR2_X1 U19440 ( .A1(n9642), .A2(n16102), .ZN(n16103) );
  OR2_X1 U19441 ( .A1(n16093), .A2(n16103), .ZN(n16228) );
  OAI22_X1 U19442 ( .A1(n16228), .A2(n9716), .B1(n16104), .B2(n10721), .ZN(
        n16105) );
  INV_X1 U19443 ( .A(n16105), .ZN(n16106) );
  OAI21_X1 U19444 ( .B1(n16107), .B2(n16154), .A(n16106), .ZN(P2_U2867) );
  AOI21_X1 U19445 ( .B1(n16108), .B2(n16113), .A(n9642), .ZN(n16237) );
  AOI22_X1 U19446 ( .A1(n16237), .A2(n16150), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n16157), .ZN(n16109) );
  OAI21_X1 U19447 ( .B1(n19754), .B2(n16154), .A(n16109), .ZN(P2_U2868) );
  NAND2_X1 U19448 ( .A1(n14720), .A2(n16110), .ZN(n16111) );
  AND2_X1 U19449 ( .A1(n16112), .A2(n16111), .ZN(n19769) );
  INV_X1 U19450 ( .A(n19769), .ZN(n16118) );
  INV_X1 U19451 ( .A(n16113), .ZN(n16114) );
  AOI21_X1 U19452 ( .B1(n16116), .B2(n16115), .A(n16114), .ZN(n16246) );
  AOI22_X1 U19453 ( .A1(n16246), .A2(n16150), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n16154), .ZN(n16117) );
  OAI21_X1 U19454 ( .B1(n16118), .B2(n16154), .A(n16117), .ZN(P2_U2869) );
  AOI21_X1 U19455 ( .B1(n16121), .B2(n16119), .A(n16120), .ZN(n16253) );
  AOI22_X1 U19456 ( .A1(n16253), .A2(n16150), .B1(P2_EBX_REG_17__SCAN_IN), 
        .B2(n16154), .ZN(n16122) );
  OAI21_X1 U19457 ( .B1(n16123), .B2(n16154), .A(n16122), .ZN(P2_U2870) );
  OR2_X1 U19458 ( .A1(n14254), .A2(n16124), .ZN(n16125) );
  NAND2_X1 U19459 ( .A1(n14717), .A2(n16125), .ZN(n19782) );
  OAI21_X1 U19460 ( .B1(n16127), .B2(n16126), .A(n16119), .ZN(n16128) );
  INV_X1 U19461 ( .A(n16128), .ZN(n16266) );
  AOI22_X1 U19462 ( .A1(n16266), .A2(n16150), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n16157), .ZN(n16129) );
  OAI21_X1 U19463 ( .B1(n19782), .B2(n16154), .A(n16129), .ZN(P2_U2871) );
  AND2_X1 U19464 ( .A1(n16130), .A2(n16131), .ZN(n16132) );
  OR2_X1 U19465 ( .A1(n16132), .A2(n14051), .ZN(n19807) );
  NOR2_X1 U19466 ( .A1(n16149), .A2(n16133), .ZN(n16141) );
  INV_X1 U19467 ( .A(n16141), .ZN(n16151) );
  OAI21_X1 U19468 ( .B1(n16151), .B2(n16135), .A(n16134), .ZN(n16137) );
  NAND3_X1 U19469 ( .A1(n16137), .A2(n16150), .A3(n16136), .ZN(n16139) );
  NAND2_X1 U19470 ( .A1(n16157), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n16138) );
  OAI211_X1 U19471 ( .C1(n19807), .C2(n16157), .A(n16139), .B(n16138), .ZN(
        P2_U2876) );
  XNOR2_X1 U19472 ( .A(n16141), .B(n16140), .ZN(n16146) );
  NAND2_X1 U19473 ( .A1(n16142), .A2(n16143), .ZN(n16144) );
  NAND2_X1 U19474 ( .A1(n16130), .A2(n16144), .ZN(n19824) );
  MUX2_X1 U19475 ( .A(n19824), .B(n19817), .S(n16157), .Z(n16145) );
  OAI21_X1 U19476 ( .B1(n16146), .B2(n9716), .A(n16145), .ZN(P2_U2877) );
  OAI21_X1 U19477 ( .B1(n16148), .B2(n16147), .A(n16142), .ZN(n19840) );
  INV_X1 U19478 ( .A(n16149), .ZN(n16153) );
  OAI211_X1 U19479 ( .C1(n16153), .C2(n16152), .A(n16151), .B(n16150), .ZN(
        n16156) );
  NAND2_X1 U19480 ( .A1(n16154), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n16155) );
  OAI211_X1 U19481 ( .C1(n19840), .C2(n16157), .A(n16156), .B(n16155), .ZN(
        P2_U2878) );
  NAND3_X1 U19482 ( .A1(n16158), .A2(n16051), .A3(n19892), .ZN(n16165) );
  INV_X1 U19483 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n16162) );
  NAND2_X1 U19484 ( .A1(n16259), .A2(BUF1_REG_29__SCAN_IN), .ZN(n16161) );
  AOI22_X1 U19485 ( .A1(n16260), .A2(n16159), .B1(n19887), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n16160) );
  OAI211_X1 U19486 ( .C1(n16162), .C2(n16264), .A(n16161), .B(n16160), .ZN(
        n16163) );
  AOI21_X1 U19487 ( .B1(n16559), .B2(n19888), .A(n16163), .ZN(n16164) );
  NAND2_X1 U19488 ( .A1(n16165), .A2(n16164), .ZN(P2_U2890) );
  INV_X1 U19489 ( .A(n16166), .ZN(n16172) );
  INV_X1 U19490 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n16170) );
  NAND2_X1 U19491 ( .A1(n16259), .A2(BUF1_REG_28__SCAN_IN), .ZN(n16169) );
  AOI22_X1 U19492 ( .A1(n16260), .A2(n16167), .B1(n19887), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n16168) );
  OAI211_X1 U19493 ( .C1(n16170), .C2(n16264), .A(n16169), .B(n16168), .ZN(
        n16171) );
  AOI21_X1 U19494 ( .B1(n16172), .B2(n19888), .A(n16171), .ZN(n16173) );
  OAI21_X1 U19495 ( .B1(n16174), .B2(n16227), .A(n16173), .ZN(P2_U2891) );
  INV_X1 U19496 ( .A(n16259), .ZN(n16200) );
  AOI22_X1 U19497 ( .A1(n16260), .A2(n16175), .B1(n19887), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n16176) );
  OAI21_X1 U19498 ( .B1(n16200), .B2(n17310), .A(n16176), .ZN(n16178) );
  NOR2_X1 U19499 ( .A1(n16572), .A2(n16282), .ZN(n16177) );
  AOI211_X1 U19500 ( .C1(n16203), .C2(BUF2_REG_27__SCAN_IN), .A(n16178), .B(
        n16177), .ZN(n16179) );
  OAI21_X1 U19501 ( .B1(n16180), .B2(n16227), .A(n16179), .ZN(P2_U2892) );
  INV_X1 U19502 ( .A(n16583), .ZN(n16186) );
  INV_X1 U19503 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n16184) );
  NAND2_X1 U19504 ( .A1(n16259), .A2(BUF1_REG_26__SCAN_IN), .ZN(n16183) );
  AOI22_X1 U19505 ( .A1(n16260), .A2(n16181), .B1(n19887), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n16182) );
  OAI211_X1 U19506 ( .C1(n16184), .C2(n16264), .A(n16183), .B(n16182), .ZN(
        n16185) );
  AOI21_X1 U19507 ( .B1(n16186), .B2(n19888), .A(n16185), .ZN(n16187) );
  OAI21_X1 U19508 ( .B1(n16188), .B2(n16227), .A(n16187), .ZN(P2_U2893) );
  INV_X1 U19509 ( .A(n16189), .ZN(n16196) );
  INV_X1 U19510 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n16193) );
  NAND2_X1 U19511 ( .A1(n16259), .A2(BUF1_REG_25__SCAN_IN), .ZN(n16192) );
  AOI22_X1 U19512 ( .A1(n16260), .A2(n16190), .B1(n19887), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n16191) );
  OAI211_X1 U19513 ( .C1(n16193), .C2(n16264), .A(n16192), .B(n16191), .ZN(
        n16194) );
  AOI21_X1 U19514 ( .B1(n16594), .B2(n19888), .A(n16194), .ZN(n16195) );
  OAI21_X1 U19515 ( .B1(n16196), .B2(n16227), .A(n16195), .ZN(P2_U2894) );
  INV_X1 U19516 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16199) );
  AOI22_X1 U19517 ( .A1(n16260), .A2(n16197), .B1(n19887), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n16198) );
  OAI21_X1 U19518 ( .B1(n16200), .B2(n16199), .A(n16198), .ZN(n16202) );
  NOR2_X1 U19519 ( .A1(n16605), .A2(n16282), .ZN(n16201) );
  AOI211_X1 U19520 ( .C1(n16203), .C2(BUF2_REG_24__SCAN_IN), .A(n16202), .B(
        n16201), .ZN(n16204) );
  OAI21_X1 U19521 ( .B1(n16205), .B2(n16227), .A(n16204), .ZN(P2_U2895) );
  INV_X1 U19522 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n16207) );
  AOI22_X1 U19523 ( .A1(n16260), .A2(n20000), .B1(n19887), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16206) );
  OAI21_X1 U19524 ( .B1(n16264), .B2(n16207), .A(n16206), .ZN(n16209) );
  NOR2_X1 U19525 ( .A1(n16612), .A2(n16282), .ZN(n16208) );
  AOI211_X1 U19526 ( .C1(BUF1_REG_23__SCAN_IN), .C2(n16259), .A(n16209), .B(
        n16208), .ZN(n16210) );
  OAI21_X1 U19527 ( .B1(n16227), .B2(n16211), .A(n16210), .ZN(P2_U2896) );
  INV_X1 U19528 ( .A(n16624), .ZN(n16218) );
  INV_X1 U19529 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n16214) );
  NAND2_X1 U19530 ( .A1(n16259), .A2(BUF1_REG_22__SCAN_IN), .ZN(n16213) );
  AOI22_X1 U19531 ( .A1(n16260), .A2(n19994), .B1(n19887), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16212) );
  OAI211_X1 U19532 ( .C1(n16264), .C2(n16214), .A(n16213), .B(n16212), .ZN(
        n16215) );
  AOI21_X1 U19533 ( .B1(n16216), .B2(n19892), .A(n16215), .ZN(n16217) );
  OAI21_X1 U19534 ( .B1(n16218), .B2(n16282), .A(n16217), .ZN(P2_U2897) );
  INV_X1 U19535 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n16221) );
  NAND2_X1 U19536 ( .A1(n16259), .A2(BUF1_REG_21__SCAN_IN), .ZN(n16220) );
  AOI22_X1 U19537 ( .A1(n16260), .A2(n19990), .B1(n19887), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n16219) );
  OAI211_X1 U19538 ( .C1(n16264), .C2(n16221), .A(n16220), .B(n16219), .ZN(
        n16222) );
  AOI21_X1 U19539 ( .B1(n16223), .B2(n19892), .A(n16222), .ZN(n16224) );
  OAI21_X1 U19540 ( .B1(n16642), .B2(n16282), .A(n16224), .ZN(P2_U2898) );
  INV_X1 U19541 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n16226) );
  AOI22_X1 U19542 ( .A1(n16260), .A2(n19985), .B1(n19887), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16225) );
  OAI21_X1 U19543 ( .B1(n16264), .B2(n16226), .A(n16225), .ZN(n16230) );
  NOR2_X1 U19544 ( .A1(n16228), .A2(n16227), .ZN(n16229) );
  AOI211_X1 U19545 ( .C1(BUF1_REG_20__SCAN_IN), .C2(n16259), .A(n16230), .B(
        n16229), .ZN(n16231) );
  OAI21_X1 U19546 ( .B1(n16232), .B2(n16282), .A(n16231), .ZN(P2_U2899) );
  INV_X1 U19547 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n16235) );
  NAND2_X1 U19548 ( .A1(n16259), .A2(BUF1_REG_19__SCAN_IN), .ZN(n16234) );
  AOI22_X1 U19549 ( .A1(n16260), .A2(n16913), .B1(n19887), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n16233) );
  OAI211_X1 U19550 ( .C1(n16264), .C2(n16235), .A(n16234), .B(n16233), .ZN(
        n16236) );
  AOI21_X1 U19551 ( .B1(n16237), .B2(n19892), .A(n16236), .ZN(n16238) );
  OAI21_X1 U19552 ( .B1(n19753), .B2(n16282), .A(n16238), .ZN(P2_U2900) );
  NAND2_X1 U19553 ( .A1(n16240), .A2(n16239), .ZN(n16241) );
  NAND2_X1 U19554 ( .A1(n14369), .A2(n16241), .ZN(n19766) );
  INV_X1 U19555 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n16244) );
  NAND2_X1 U19556 ( .A1(n16259), .A2(BUF1_REG_18__SCAN_IN), .ZN(n16243) );
  AOI22_X1 U19557 ( .A1(n16260), .A2(n19977), .B1(n19887), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16242) );
  OAI211_X1 U19558 ( .C1(n16264), .C2(n16244), .A(n16243), .B(n16242), .ZN(
        n16245) );
  AOI21_X1 U19559 ( .B1(n16246), .B2(n19892), .A(n16245), .ZN(n16247) );
  OAI21_X1 U19560 ( .B1(n16282), .B2(n19766), .A(n16247), .ZN(P2_U2901) );
  INV_X1 U19561 ( .A(n16248), .ZN(n16255) );
  INV_X1 U19562 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n16251) );
  NAND2_X1 U19563 ( .A1(n16259), .A2(BUF1_REG_17__SCAN_IN), .ZN(n16250) );
  AOI22_X1 U19564 ( .A1(n16260), .A2(n19973), .B1(n19887), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n16249) );
  OAI211_X1 U19565 ( .C1(n16264), .C2(n16251), .A(n16250), .B(n16249), .ZN(
        n16252) );
  AOI21_X1 U19566 ( .B1(n16253), .B2(n19892), .A(n16252), .ZN(n16254) );
  OAI21_X1 U19567 ( .B1(n16255), .B2(n16282), .A(n16254), .ZN(P2_U2902) );
  OR2_X1 U19568 ( .A1(n16256), .A2(n16257), .ZN(n16258) );
  AND2_X1 U19569 ( .A1(n14725), .A2(n16258), .ZN(n16659) );
  INV_X1 U19570 ( .A(n16659), .ZN(n19781) );
  INV_X1 U19571 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n16263) );
  NAND2_X1 U19572 ( .A1(n16259), .A2(BUF1_REG_16__SCAN_IN), .ZN(n16262) );
  AOI22_X1 U19573 ( .A1(n16260), .A2(n16881), .B1(n19887), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n16261) );
  OAI211_X1 U19574 ( .C1(n16264), .C2(n16263), .A(n16262), .B(n16261), .ZN(
        n16265) );
  AOI21_X1 U19575 ( .B1(n16266), .B2(n19892), .A(n16265), .ZN(n16267) );
  OAI21_X1 U19576 ( .B1(n19781), .B2(n16282), .A(n16267), .ZN(P2_U2903) );
  OAI21_X1 U19577 ( .B1(n9608), .B2(n16268), .A(n10511), .ZN(n19794) );
  OAI222_X1 U19578 ( .A1(n19794), .A2(n16275), .B1(n16287), .B2(n13398), .C1(
        n16269), .C2(n19896), .ZN(P2_U2904) );
  NOR2_X1 U19579 ( .A1(n20656), .A2(n20653), .ZN(n16270) );
  AOI21_X1 U19580 ( .B1(n20656), .B2(n20653), .A(n16270), .ZN(n19891) );
  NAND2_X1 U19581 ( .A1(n19891), .A2(n19890), .ZN(n19889) );
  INV_X1 U19582 ( .A(n16270), .ZN(n16271) );
  NAND2_X1 U19583 ( .A1(n19889), .A2(n16271), .ZN(n16284) );
  XOR2_X1 U19584 ( .A(n20645), .B(n20647), .Z(n16285) );
  NAND2_X1 U19585 ( .A1(n16284), .A2(n16285), .ZN(n16283) );
  OAI21_X1 U19586 ( .B1(n20647), .B2(n20645), .A(n16283), .ZN(n19881) );
  XNOR2_X1 U19587 ( .A(n20637), .B(n17226), .ZN(n19882) );
  NAND2_X1 U19588 ( .A1(n19881), .A2(n19882), .ZN(n19880) );
  OAI21_X1 U19589 ( .B1(n20637), .B2(n20635), .A(n19880), .ZN(n16272) );
  NAND2_X1 U19590 ( .A1(n16272), .A2(n16809), .ZN(n16276) );
  NAND3_X1 U19591 ( .A1(n16276), .A2(n19892), .A3(n16277), .ZN(n16274) );
  INV_X1 U19592 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19923) );
  AOI22_X1 U19593 ( .A1(n16279), .A2(n19990), .B1(n19887), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n16273) );
  OAI211_X1 U19594 ( .C1(n16275), .C2(n16797), .A(n16274), .B(n16273), .ZN(
        P2_U2914) );
  XOR2_X1 U19595 ( .A(n16277), .B(n16276), .Z(n16278) );
  NAND2_X1 U19596 ( .A1(n16278), .A2(n19892), .ZN(n16281) );
  AOI22_X1 U19597 ( .A1(n16279), .A2(n19985), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19887), .ZN(n16280) );
  OAI211_X1 U19598 ( .C1(n16809), .C2(n16282), .A(n16281), .B(n16280), .ZN(
        P2_U2915) );
  OAI21_X1 U19599 ( .B1(n16285), .B2(n16284), .A(n16283), .ZN(n16286) );
  NAND2_X1 U19600 ( .A1(n16286), .A2(n19892), .ZN(n16291) );
  INV_X1 U19601 ( .A(n19977), .ZN(n16288) );
  INV_X1 U19602 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n21413) );
  OAI22_X1 U19603 ( .A1(n19896), .A2(n16288), .B1(n16287), .B2(n21413), .ZN(
        n16289) );
  AOI21_X1 U19604 ( .B1(n19888), .B2(n20645), .A(n16289), .ZN(n16290) );
  NAND2_X1 U19605 ( .A1(n16291), .A2(n16290), .ZN(P2_U2917) );
  NAND2_X1 U19606 ( .A1(n16294), .A2(n16293), .ZN(n16295) );
  XOR2_X1 U19607 ( .A(n16292), .B(n16295), .Z(n16565) );
  NOR2_X1 U19608 ( .A1(n16296), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16297) );
  NOR2_X1 U19609 ( .A1(n16491), .A2(n20612), .ZN(n16556) );
  AOI21_X1 U19610 ( .B1(n16510), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16556), .ZN(n16300) );
  NAND2_X1 U19611 ( .A1(n19943), .A2(n10537), .ZN(n16299) );
  OAI211_X1 U19612 ( .C1(n16562), .C2(n19950), .A(n16300), .B(n16299), .ZN(
        n16301) );
  AOI21_X1 U19613 ( .B1(n19945), .B2(n10546), .A(n16301), .ZN(n16302) );
  OAI21_X1 U19614 ( .B1(n16565), .B2(n16483), .A(n16302), .ZN(P2_U2985) );
  NAND2_X1 U19615 ( .A1(n16303), .A2(n16547), .ZN(n16306) );
  AOI21_X1 U19616 ( .B1(n16510), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16304), .ZN(n16305) );
  OAI211_X1 U19617 ( .C1(n16544), .C2(n16307), .A(n16306), .B(n16305), .ZN(
        n16308) );
  AOI21_X1 U19618 ( .B1(n19945), .B2(n16309), .A(n16308), .ZN(n16310) );
  OAI21_X1 U19619 ( .B1(n16311), .B2(n16483), .A(n16310), .ZN(P2_U2986) );
  OAI21_X1 U19620 ( .B1(n16314), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16313), .ZN(n16577) );
  XNOR2_X1 U19621 ( .A(n16317), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16318) );
  NAND2_X1 U19622 ( .A1(n16566), .A2(n10145), .ZN(n16325) );
  NAND2_X1 U19623 ( .A1(n19941), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n16567) );
  OAI21_X1 U19624 ( .B1(n19955), .B2(n16319), .A(n16567), .ZN(n16322) );
  NOR2_X1 U19625 ( .A1(n16320), .A2(n19950), .ZN(n16321) );
  AOI211_X1 U19626 ( .C1(n19943), .C2(n16323), .A(n16322), .B(n16321), .ZN(
        n16324) );
  OAI211_X1 U19627 ( .C1(n16550), .C2(n16577), .A(n16325), .B(n16324), .ZN(
        P2_U2987) );
  NOR2_X1 U19628 ( .A1(n16491), .A2(n20607), .ZN(n16581) );
  AOI21_X1 U19629 ( .B1(n16510), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16581), .ZN(n16330) );
  OAI21_X1 U19630 ( .B1(n16544), .B2(n16331), .A(n16330), .ZN(n16332) );
  NAND2_X1 U19631 ( .A1(n16334), .A2(n16333), .ZN(n16335) );
  XNOR2_X1 U19632 ( .A(n16336), .B(n16335), .ZN(n16598) );
  NOR2_X1 U19633 ( .A1(n16491), .A2(n20605), .ZN(n16587) );
  INV_X1 U19634 ( .A(n16587), .ZN(n16337) );
  OAI21_X1 U19635 ( .B1(n19955), .B2(n16338), .A(n16337), .ZN(n16340) );
  NOR2_X1 U19636 ( .A1(n16591), .A2(n19950), .ZN(n16339) );
  AOI211_X1 U19637 ( .C1(n19943), .C2(n16341), .A(n16340), .B(n16339), .ZN(
        n16343) );
  NAND2_X1 U19638 ( .A1(n9583), .A2(n16578), .ZN(n16595) );
  NAND3_X1 U19639 ( .A1(n9645), .A2(n19945), .A3(n16595), .ZN(n16342) );
  OAI211_X1 U19640 ( .C1(n16598), .C2(n16483), .A(n16343), .B(n16342), .ZN(
        P2_U2989) );
  XNOR2_X1 U19641 ( .A(n16348), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16361) );
  NAND2_X1 U19642 ( .A1(n19941), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n16599) );
  NAND2_X1 U19643 ( .A1(n16510), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16349) );
  OAI211_X1 U19644 ( .C1(n16544), .C2(n16350), .A(n16599), .B(n16349), .ZN(
        n16352) );
  INV_X1 U19645 ( .A(n16351), .ZN(n16355) );
  OAI21_X1 U19646 ( .B1(n16630), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16355), .ZN(n16622) );
  INV_X1 U19647 ( .A(n16356), .ZN(n16360) );
  OR2_X1 U19648 ( .A1(n16491), .A2(n20601), .ZN(n16614) );
  OAI21_X1 U19649 ( .B1(n19955), .B2(n16357), .A(n16614), .ZN(n16359) );
  NOR2_X1 U19650 ( .A1(n16611), .A2(n19950), .ZN(n16358) );
  AOI211_X1 U19651 ( .C1(n16360), .C2(n19943), .A(n16359), .B(n16358), .ZN(
        n16364) );
  OR2_X1 U19652 ( .A1(n16362), .A2(n16361), .ZN(n16610) );
  NAND3_X1 U19653 ( .A1(n16610), .A2(n16609), .A3(n10145), .ZN(n16363) );
  OAI211_X1 U19654 ( .C1(n16550), .C2(n16622), .A(n16364), .B(n16363), .ZN(
        P2_U2991) );
  INV_X1 U19655 ( .A(n16365), .ZN(n16367) );
  NAND2_X1 U19656 ( .A1(n16367), .A2(n16366), .ZN(n16368) );
  XNOR2_X1 U19657 ( .A(n16369), .B(n16368), .ZN(n16634) );
  INV_X1 U19658 ( .A(n16370), .ZN(n16633) );
  INV_X1 U19659 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n16371) );
  NOR2_X1 U19660 ( .A1(n16491), .A2(n16371), .ZN(n16626) );
  AOI21_X1 U19661 ( .B1(n16510), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16626), .ZN(n16372) );
  OAI21_X1 U19662 ( .B1(n16544), .B2(n16373), .A(n16372), .ZN(n16375) );
  INV_X1 U19663 ( .A(n16353), .ZN(n16374) );
  NAND2_X1 U19664 ( .A1(n16380), .A2(n16379), .ZN(n16381) );
  XNOR2_X1 U19665 ( .A(n16382), .B(n16381), .ZN(n16647) );
  NOR2_X1 U19666 ( .A1(n16491), .A2(n20599), .ZN(n16635) );
  AOI21_X1 U19667 ( .B1(n16510), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16635), .ZN(n16383) );
  OAI21_X1 U19668 ( .B1(n16544), .B2(n16384), .A(n16383), .ZN(n16386) );
  OAI21_X1 U19669 ( .B1(n16647), .B2(n16483), .A(n16387), .ZN(P2_U2993) );
  NAND2_X1 U19670 ( .A1(n16389), .A2(n16388), .ZN(n16390) );
  XNOR2_X1 U19671 ( .A(n16391), .B(n16390), .ZN(n16657) );
  NAND2_X1 U19672 ( .A1(n19941), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n16648) );
  NAND2_X1 U19673 ( .A1(n16510), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16392) );
  OAI211_X1 U19674 ( .C1(n16544), .C2(n19760), .A(n16648), .B(n16392), .ZN(
        n16393) );
  AOI21_X1 U19675 ( .B1(n19769), .B2(n16547), .A(n16393), .ZN(n16396) );
  XNOR2_X1 U19676 ( .A(n16394), .B(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16654) );
  NAND2_X1 U19677 ( .A1(n16654), .A2(n19945), .ZN(n16395) );
  OAI211_X1 U19678 ( .C1(n16657), .C2(n16483), .A(n16396), .B(n16395), .ZN(
        P2_U2996) );
  OAI21_X1 U19679 ( .B1(n16399), .B2(n16398), .A(n16397), .ZN(n16667) );
  XNOR2_X1 U19680 ( .A(n16410), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16403) );
  NOR2_X1 U19681 ( .A1(n16491), .A2(n20591), .ZN(n16658) );
  NOR2_X1 U19682 ( .A1(n16544), .A2(n19775), .ZN(n16400) );
  AOI211_X1 U19683 ( .C1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n16510), .A(
        n16658), .B(n16400), .ZN(n16401) );
  OAI21_X1 U19684 ( .B1(n19782), .B2(n19950), .A(n16401), .ZN(n16402) );
  AOI21_X1 U19685 ( .B1(n16403), .B2(n19945), .A(n16402), .ZN(n16404) );
  OAI21_X1 U19686 ( .B1(n16667), .B2(n16483), .A(n16404), .ZN(P2_U2998) );
  NAND2_X1 U19687 ( .A1(n10301), .A2(n16406), .ZN(n16407) );
  XNOR2_X1 U19688 ( .A(n16408), .B(n16407), .ZN(n16678) );
  INV_X1 U19689 ( .A(n16410), .ZN(n16411) );
  AOI21_X1 U19690 ( .B1(n16412), .B2(n16422), .A(n16411), .ZN(n16676) );
  NOR2_X1 U19691 ( .A1(n16491), .A2(n20589), .ZN(n16671) );
  NOR2_X1 U19692 ( .A1(n19955), .A2(n19793), .ZN(n16413) );
  AOI211_X1 U19693 ( .C1(n19789), .C2(n19943), .A(n16671), .B(n16413), .ZN(
        n16414) );
  OAI21_X1 U19694 ( .B1(n19795), .B2(n19950), .A(n16414), .ZN(n16415) );
  AOI21_X1 U19695 ( .B1(n16676), .B2(n19945), .A(n16415), .ZN(n16416) );
  OAI21_X1 U19696 ( .B1(n16678), .B2(n16483), .A(n16416), .ZN(P2_U2999) );
  NAND2_X1 U19697 ( .A1(n16418), .A2(n16417), .ZN(n16419) );
  NOR2_X1 U19698 ( .A1(n16491), .A2(n20587), .ZN(n16686) );
  AOI21_X1 U19699 ( .B1(n16510), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16686), .ZN(n16420) );
  OAI21_X1 U19700 ( .B1(n16544), .B2(n16421), .A(n16420), .ZN(n16423) );
  AOI21_X1 U19701 ( .B1(n16426), .B2(n16425), .A(n16424), .ZN(n16704) );
  NOR2_X1 U19702 ( .A1(n16491), .A2(n16427), .ZN(n16696) );
  AOI21_X1 U19703 ( .B1(n16510), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16696), .ZN(n16428) );
  OAI21_X1 U19704 ( .B1(n16544), .B2(n16429), .A(n16428), .ZN(n16430) );
  AOI21_X1 U19705 ( .B1(n16695), .B2(n16547), .A(n16430), .ZN(n16433) );
  OAI211_X1 U19706 ( .C1(n16704), .C2(n16483), .A(n16433), .B(n16432), .ZN(
        P2_U3001) );
  NAND2_X1 U19707 ( .A1(n16435), .A2(n16434), .ZN(n16439) );
  XOR2_X1 U19708 ( .A(n16439), .B(n16438), .Z(n16715) );
  INV_X1 U19709 ( .A(n16710), .ZN(n16445) );
  NOR2_X1 U19710 ( .A1(n16491), .A2(n16440), .ZN(n16707) );
  AOI21_X1 U19711 ( .B1(n16510), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16707), .ZN(n16441) );
  OAI21_X1 U19712 ( .B1(n16544), .B2(n16442), .A(n16441), .ZN(n16444) );
  OAI21_X1 U19713 ( .B1(n16715), .B2(n16483), .A(n16446), .ZN(P2_U3002) );
  XNOR2_X1 U19714 ( .A(n16447), .B(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16448) );
  XNOR2_X1 U19715 ( .A(n16449), .B(n16448), .ZN(n16726) );
  INV_X1 U19716 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16465) );
  NOR2_X1 U19717 ( .A1(n16491), .A2(n20583), .ZN(n16719) );
  NOR2_X1 U19718 ( .A1(n16544), .A2(n19811), .ZN(n16452) );
  AOI211_X1 U19719 ( .C1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n16510), .A(
        n16719), .B(n16452), .ZN(n16453) );
  OAI21_X1 U19720 ( .B1(n19807), .B2(n19950), .A(n16453), .ZN(n16454) );
  AOI21_X1 U19721 ( .B1(n16724), .B2(n19945), .A(n16454), .ZN(n16455) );
  OAI21_X1 U19722 ( .B1(n16726), .B2(n16483), .A(n16455), .ZN(P2_U3003) );
  INV_X1 U19723 ( .A(n16458), .ZN(n16459) );
  OAI21_X1 U19724 ( .B1(n16505), .B2(n16460), .A(n16459), .ZN(n16475) );
  OAI21_X1 U19725 ( .B1(n16475), .B2(n16471), .A(n16472), .ZN(n16463) );
  NOR2_X1 U19726 ( .A1(n10545), .A2(n16461), .ZN(n16462) );
  XNOR2_X1 U19727 ( .A(n16463), .B(n16462), .ZN(n16737) );
  AOI21_X1 U19728 ( .B1(n16465), .B2(n16476), .A(n16464), .ZN(n16735) );
  NOR2_X1 U19729 ( .A1(n16491), .A2(n20581), .ZN(n16728) );
  NOR2_X1 U19730 ( .A1(n16544), .A2(n16466), .ZN(n16467) );
  AOI211_X1 U19731 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n16510), .A(
        n16728), .B(n16467), .ZN(n16468) );
  OAI21_X1 U19732 ( .B1(n19824), .B2(n19950), .A(n16468), .ZN(n16469) );
  AOI21_X1 U19733 ( .B1(n16735), .B2(n19945), .A(n16469), .ZN(n16470) );
  OAI21_X1 U19734 ( .B1(n16737), .B2(n16483), .A(n16470), .ZN(P2_U3004) );
  INV_X1 U19735 ( .A(n16471), .ZN(n16473) );
  NAND2_X1 U19736 ( .A1(n16473), .A2(n16472), .ZN(n16474) );
  XNOR2_X1 U19737 ( .A(n16475), .B(n16474), .ZN(n16749) );
  INV_X1 U19738 ( .A(n16476), .ZN(n16477) );
  AOI21_X1 U19739 ( .B1(n16478), .B2(n16739), .A(n16477), .ZN(n16747) );
  NOR2_X1 U19740 ( .A1(n16491), .A2(n20579), .ZN(n16742) );
  AOI21_X1 U19741 ( .B1(n16510), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16742), .ZN(n16480) );
  NAND2_X1 U19742 ( .A1(n19943), .A2(n19830), .ZN(n16479) );
  OAI211_X1 U19743 ( .C1(n19840), .C2(n19950), .A(n16480), .B(n16479), .ZN(
        n16481) );
  AOI21_X1 U19744 ( .B1(n16747), .B2(n19945), .A(n16481), .ZN(n16482) );
  OAI21_X1 U19745 ( .B1(n16749), .B2(n16483), .A(n16482), .ZN(P2_U3005) );
  INV_X1 U19746 ( .A(n16504), .ZN(n16484) );
  AOI21_X1 U19747 ( .B1(n16505), .B2(n16503), .A(n16484), .ZN(n16488) );
  NAND2_X1 U19748 ( .A1(n16486), .A2(n16485), .ZN(n16487) );
  XNOR2_X1 U19749 ( .A(n16488), .B(n16487), .ZN(n16761) );
  INV_X1 U19750 ( .A(n16756), .ZN(n16502) );
  NAND2_X1 U19751 ( .A1(n19943), .A2(n16489), .ZN(n16492) );
  OR2_X1 U19752 ( .A1(n16491), .A2(n16490), .ZN(n16751) );
  OAI211_X1 U19753 ( .C1(n16493), .C2(n19955), .A(n16492), .B(n16751), .ZN(
        n16501) );
  INV_X1 U19754 ( .A(n16494), .ZN(n16497) );
  NAND2_X1 U19755 ( .A1(n16494), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16496) );
  NAND2_X1 U19756 ( .A1(n16498), .A2(n16495), .ZN(n16507) );
  AOI22_X1 U19757 ( .A1(n16497), .A2(n16763), .B1(n16496), .B2(n16507), .ZN(
        n16499) );
  XNOR2_X1 U19758 ( .A(n16498), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16500) );
  NAND2_X1 U19759 ( .A1(n16504), .A2(n16503), .ZN(n16506) );
  XOR2_X1 U19760 ( .A(n16506), .B(n16505), .Z(n16772) );
  XNOR2_X1 U19761 ( .A(n16507), .B(n16763), .ZN(n16508) );
  XNOR2_X1 U19762 ( .A(n16494), .B(n16508), .ZN(n16770) );
  NOR2_X1 U19763 ( .A1(n16491), .A2(n20576), .ZN(n16765) );
  NOR2_X1 U19764 ( .A1(n16544), .A2(n19848), .ZN(n16509) );
  AOI211_X1 U19765 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n16510), .A(
        n16765), .B(n16509), .ZN(n16511) );
  OAI21_X1 U19766 ( .B1(n19853), .B2(n19950), .A(n16511), .ZN(n16512) );
  AOI21_X1 U19767 ( .B1(n16770), .B2(n19945), .A(n16512), .ZN(n16513) );
  OAI21_X1 U19768 ( .B1(n16772), .B2(n16483), .A(n16513), .ZN(P2_U3007) );
  XNOR2_X1 U19769 ( .A(n16515), .B(n16514), .ZN(n16786) );
  INV_X1 U19770 ( .A(n11541), .ZN(n16520) );
  NOR2_X1 U19771 ( .A1(n16520), .A2(n16517), .ZN(n16516) );
  AOI211_X1 U19772 ( .C1(n16520), .C2(n16519), .A(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n16518), .ZN(n16522) );
  NOR2_X1 U19773 ( .A1(n16522), .A2(n16521), .ZN(n16784) );
  NOR2_X1 U19774 ( .A1(n16491), .A2(n20574), .ZN(n16776) );
  INV_X1 U19775 ( .A(n16776), .ZN(n16523) );
  OAI21_X1 U19776 ( .B1(n19955), .B2(n19879), .A(n16523), .ZN(n16524) );
  AOI21_X1 U19777 ( .B1(n19943), .B2(n19868), .A(n16524), .ZN(n16525) );
  OAI21_X1 U19778 ( .B1(n19872), .B2(n19950), .A(n16525), .ZN(n16526) );
  AOI21_X1 U19779 ( .B1(n16784), .B2(n19945), .A(n16526), .ZN(n16527) );
  OAI21_X1 U19780 ( .B1(n16483), .B2(n16786), .A(n16527), .ZN(P2_U3008) );
  XNOR2_X1 U19781 ( .A(n16529), .B(n16528), .ZN(n16803) );
  NOR2_X1 U19782 ( .A1(n16544), .A2(n16530), .ZN(n16533) );
  NAND2_X1 U19783 ( .A1(n19941), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n16788) );
  OAI21_X1 U19784 ( .B1(n19955), .B2(n16531), .A(n16788), .ZN(n16532) );
  AOI211_X1 U19785 ( .C1(n16787), .C2(n16547), .A(n16533), .B(n16532), .ZN(
        n16537) );
  NAND2_X1 U19786 ( .A1(n11541), .A2(n16534), .ZN(n16535) );
  XNOR2_X1 U19787 ( .A(n11538), .B(n16535), .ZN(n16800) );
  NAND2_X1 U19788 ( .A1(n16800), .A2(n19945), .ZN(n16536) );
  OAI211_X1 U19789 ( .C1(n16803), .C2(n16483), .A(n16537), .B(n16536), .ZN(
        P2_U3009) );
  XNOR2_X1 U19790 ( .A(n16539), .B(n16538), .ZN(n17229) );
  XNOR2_X1 U19791 ( .A(n16540), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16541) );
  XNOR2_X1 U19792 ( .A(n16542), .B(n16541), .ZN(n17231) );
  NAND2_X1 U19793 ( .A1(n17231), .A2(n10145), .ZN(n16549) );
  NOR2_X1 U19794 ( .A1(n16544), .A2(n16543), .ZN(n16546) );
  NAND2_X1 U19795 ( .A1(n19941), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n17225) );
  OAI21_X1 U19796 ( .B1(n19955), .B2(n10396), .A(n17225), .ZN(n16545) );
  AOI211_X1 U19797 ( .C1(n16008), .C2(n16547), .A(n16546), .B(n16545), .ZN(
        n16548) );
  OAI211_X1 U19798 ( .C1(n17229), .C2(n16550), .A(n16549), .B(n16548), .ZN(
        P2_U3011) );
  NAND2_X1 U19799 ( .A1(n16552), .A2(n16551), .ZN(n16553) );
  AOI21_X1 U19800 ( .B1(n16554), .B2(n16553), .A(n16557), .ZN(n16555) );
  AOI211_X1 U19801 ( .C1(n16558), .C2(n16557), .A(n16556), .B(n16555), .ZN(
        n16561) );
  NAND2_X1 U19802 ( .A1(n16559), .A2(n19956), .ZN(n16560) );
  OAI211_X1 U19803 ( .C1(n16562), .C2(n16782), .A(n16561), .B(n16560), .ZN(
        n16563) );
  AOI21_X1 U19804 ( .B1(n16799), .B2(n10546), .A(n16563), .ZN(n16564) );
  OAI21_X1 U19805 ( .B1(n16565), .B2(n16802), .A(n16564), .ZN(P2_U3017) );
  INV_X1 U19806 ( .A(n16567), .ZN(n16569) );
  AOI211_X1 U19807 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n16570), .A(
        n16569), .B(n16568), .ZN(n16571) );
  OAI21_X1 U19808 ( .B1(n16572), .B2(n17237), .A(n16571), .ZN(n16573) );
  AOI21_X1 U19809 ( .B1(n16574), .B2(n19967), .A(n16573), .ZN(n16575) );
  OAI211_X1 U19810 ( .C1(n16577), .C2(n19970), .A(n16576), .B(n16575), .ZN(
        P2_U3019) );
  AOI211_X1 U19811 ( .C1(n16579), .C2(n16578), .A(n11549), .B(n16590), .ZN(
        n16580) );
  AOI211_X1 U19812 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n16588), .A(
        n16581), .B(n16580), .ZN(n16582) );
  OAI21_X1 U19813 ( .B1(n16583), .B2(n17237), .A(n16582), .ZN(n16584) );
  AOI21_X1 U19814 ( .B1(n16588), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n16587), .ZN(n16589) );
  OAI21_X1 U19815 ( .B1(n16590), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n16589), .ZN(n16593) );
  NOR2_X1 U19816 ( .A1(n16591), .A2(n16782), .ZN(n16592) );
  AOI211_X1 U19817 ( .C1(n19956), .C2(n16594), .A(n16593), .B(n16592), .ZN(
        n16597) );
  NAND3_X1 U19818 ( .A1(n9645), .A2(n16799), .A3(n16595), .ZN(n16596) );
  OAI211_X1 U19819 ( .C1(n16598), .C2(n16802), .A(n16597), .B(n16596), .ZN(
        P2_U3021) );
  INV_X1 U19820 ( .A(n16599), .ZN(n16600) );
  AOI21_X1 U19821 ( .B1(n16601), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n16600), .ZN(n16604) );
  NAND3_X1 U19822 ( .A1(n16623), .A2(n16602), .A3(n9891), .ZN(n16603) );
  OAI211_X1 U19823 ( .C1(n16605), .C2(n17237), .A(n16604), .B(n16603), .ZN(
        n16606) );
  NAND3_X1 U19824 ( .A1(n16610), .A2(n16609), .A3(n19958), .ZN(n16621) );
  INV_X1 U19825 ( .A(n16611), .ZN(n16619) );
  NOR2_X1 U19826 ( .A1(n16612), .A2(n17237), .ZN(n16618) );
  OAI211_X1 U19827 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16623), .B(n16613), .ZN(
        n16615) );
  OAI211_X1 U19828 ( .C1(n16616), .C2(n16625), .A(n16615), .B(n16614), .ZN(
        n16617) );
  AOI211_X1 U19829 ( .C1(n16619), .C2(n19967), .A(n16618), .B(n16617), .ZN(
        n16620) );
  OAI211_X1 U19830 ( .C1(n16622), .C2(n19970), .A(n16621), .B(n16620), .ZN(
        P2_U3023) );
  INV_X1 U19831 ( .A(n16623), .ZN(n16629) );
  NAND2_X1 U19832 ( .A1(n16624), .A2(n19956), .ZN(n16628) );
  INV_X1 U19833 ( .A(n16625), .ZN(n16636) );
  AOI21_X1 U19834 ( .B1(n16636), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n16626), .ZN(n16627) );
  OAI211_X1 U19835 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n16629), .A(
        n16628), .B(n16627), .ZN(n16632) );
  AOI21_X1 U19836 ( .B1(n16636), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n16635), .ZN(n16641) );
  NAND4_X1 U19837 ( .A1(n16639), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n16638), .A4(n16637), .ZN(n16640) );
  OAI211_X1 U19838 ( .C1(n16642), .C2(n17237), .A(n16641), .B(n16640), .ZN(
        n16644) );
  OAI21_X1 U19839 ( .B1(n16647), .B2(n16802), .A(n16646), .ZN(P2_U3025) );
  NOR2_X1 U19840 ( .A1(n19766), .A2(n17237), .ZN(n16653) );
  OAI211_X1 U19841 ( .C1(n16651), .C2(n16650), .A(n16649), .B(n16648), .ZN(
        n16652) );
  AOI211_X1 U19842 ( .C1(n19769), .C2(n19967), .A(n16653), .B(n16652), .ZN(
        n16656) );
  NAND2_X1 U19843 ( .A1(n16654), .A2(n16799), .ZN(n16655) );
  OAI211_X1 U19844 ( .C1(n16657), .C2(n16802), .A(n16656), .B(n16655), .ZN(
        P2_U3028) );
  AOI21_X1 U19845 ( .B1(n16659), .B2(n19956), .A(n16658), .ZN(n16660) );
  OAI21_X1 U19846 ( .B1(n19782), .B2(n16782), .A(n16660), .ZN(n16661) );
  AOI21_X1 U19847 ( .B1(n16662), .B2(n16663), .A(n16661), .ZN(n16666) );
  OAI211_X1 U19848 ( .C1(n16667), .C2(n16802), .A(n16666), .B(n16665), .ZN(
        P2_U3030) );
  NOR2_X1 U19849 ( .A1(n19795), .A2(n16782), .ZN(n16675) );
  NOR3_X1 U19850 ( .A1(n16669), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        n16668), .ZN(n16670) );
  AOI211_X1 U19851 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16672), .A(
        n16671), .B(n16670), .ZN(n16673) );
  OAI21_X1 U19852 ( .B1(n17237), .B2(n19794), .A(n16673), .ZN(n16674) );
  AOI211_X1 U19853 ( .C1(n16676), .C2(n16799), .A(n16675), .B(n16674), .ZN(
        n16677) );
  OAI21_X1 U19854 ( .B1(n16678), .B2(n16802), .A(n16677), .ZN(P2_U3031) );
  AND2_X1 U19855 ( .A1(n16738), .A2(n16683), .ZN(n16714) );
  AND2_X1 U19856 ( .A1(n16679), .A2(n10376), .ZN(n16680) );
  NOR2_X1 U19857 ( .A1(n16681), .A2(n16680), .ZN(n16692) );
  NAND2_X1 U19858 ( .A1(n16682), .A2(n19967), .ZN(n16688) );
  NAND2_X1 U19859 ( .A1(n16740), .A2(n16683), .ZN(n16684) );
  AND2_X1 U19860 ( .A1(n16685), .A2(n16684), .ZN(n16708) );
  AOI21_X1 U19861 ( .B1(n16708), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16686), .ZN(n16687) );
  OAI211_X1 U19862 ( .C1(n17237), .C2(n16689), .A(n16688), .B(n16687), .ZN(
        n16691) );
  XNOR2_X1 U19863 ( .A(n16694), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16701) );
  NAND2_X1 U19864 ( .A1(n16695), .A2(n19967), .ZN(n16698) );
  AOI21_X1 U19865 ( .B1(n16708), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n16696), .ZN(n16697) );
  OAI211_X1 U19866 ( .C1(n17237), .C2(n16699), .A(n16698), .B(n16697), .ZN(
        n16700) );
  AOI21_X1 U19867 ( .B1(n16714), .B2(n16701), .A(n16700), .ZN(n16703) );
  OAI211_X1 U19868 ( .C1(n16704), .C2(n16802), .A(n16703), .B(n16702), .ZN(
        P2_U3033) );
  NOR2_X1 U19869 ( .A1(n16705), .A2(n17237), .ZN(n16706) );
  AOI211_X1 U19870 ( .C1(n16708), .C2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n16707), .B(n16706), .ZN(n16709) );
  OAI21_X1 U19871 ( .B1(n16782), .B2(n16710), .A(n16709), .ZN(n16712) );
  NAND2_X1 U19872 ( .A1(n16738), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16727) );
  OAI21_X1 U19873 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n16716), .ZN(n16717) );
  NOR2_X1 U19874 ( .A1(n16727), .A2(n16717), .ZN(n16723) );
  OR2_X1 U19875 ( .A1(n19961), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16718) );
  NAND2_X1 U19876 ( .A1(n16740), .A2(n16718), .ZN(n16729) );
  AOI21_X1 U19877 ( .B1(n16729), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16719), .ZN(n16721) );
  NAND2_X1 U19878 ( .A1(n19804), .A2(n19956), .ZN(n16720) );
  OAI211_X1 U19879 ( .C1(n19807), .C2(n16782), .A(n16721), .B(n16720), .ZN(
        n16722) );
  AOI211_X1 U19880 ( .C1(n16724), .C2(n16799), .A(n16723), .B(n16722), .ZN(
        n16725) );
  OAI21_X1 U19881 ( .B1(n16726), .B2(n16802), .A(n16725), .ZN(P2_U3035) );
  NOR2_X1 U19882 ( .A1(n16727), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16734) );
  AOI21_X1 U19883 ( .B1(n16729), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16728), .ZN(n16732) );
  NAND2_X1 U19884 ( .A1(n16730), .A2(n19956), .ZN(n16731) );
  OAI211_X1 U19885 ( .C1(n19824), .C2(n16782), .A(n16732), .B(n16731), .ZN(
        n16733) );
  AOI211_X1 U19886 ( .C1(n16735), .C2(n16799), .A(n16734), .B(n16733), .ZN(
        n16736) );
  OAI21_X1 U19887 ( .B1(n16737), .B2(n16802), .A(n16736), .ZN(P2_U3036) );
  NAND2_X1 U19888 ( .A1(n16738), .A2(n16739), .ZN(n16745) );
  NOR2_X1 U19889 ( .A1(n16740), .A2(n16739), .ZN(n16741) );
  AOI211_X1 U19890 ( .C1(n16743), .C2(n19956), .A(n16742), .B(n16741), .ZN(
        n16744) );
  OAI211_X1 U19891 ( .C1(n19840), .C2(n16782), .A(n16745), .B(n16744), .ZN(
        n16746) );
  AOI21_X1 U19892 ( .B1(n16747), .B2(n16799), .A(n16746), .ZN(n16748) );
  OAI21_X1 U19893 ( .B1(n16749), .B2(n16802), .A(n16748), .ZN(P2_U3037) );
  XNOR2_X1 U19894 ( .A(n16763), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16760) );
  INV_X1 U19895 ( .A(n16789), .ZN(n16811) );
  NAND3_X1 U19896 ( .A1(n16811), .A2(n16790), .A3(n16775), .ZN(n16774) );
  OAI21_X1 U19897 ( .B1(n19961), .B2(n16790), .A(n16774), .ZN(n16750) );
  NOR2_X1 U19898 ( .A1(n16810), .A2(n16750), .ZN(n16773) );
  OAI21_X1 U19899 ( .B1(n16773), .B2(n16752), .A(n16751), .ZN(n16753) );
  AOI21_X1 U19900 ( .B1(n16754), .B2(n19956), .A(n16753), .ZN(n16755) );
  OAI21_X1 U19901 ( .B1(n16756), .B2(n16782), .A(n16755), .ZN(n16759) );
  NAND2_X1 U19902 ( .A1(n16762), .A2(n16763), .ZN(n16768) );
  INV_X1 U19903 ( .A(n19852), .ZN(n16766) );
  NOR2_X1 U19904 ( .A1(n16773), .A2(n16763), .ZN(n16764) );
  AOI211_X1 U19905 ( .C1(n16766), .C2(n19956), .A(n16765), .B(n16764), .ZN(
        n16767) );
  OAI211_X1 U19906 ( .C1(n19853), .C2(n16782), .A(n16768), .B(n16767), .ZN(
        n16769) );
  AOI21_X1 U19907 ( .B1(n16770), .B2(n16799), .A(n16769), .ZN(n16771) );
  OAI21_X1 U19908 ( .B1(n16772), .B2(n16802), .A(n16771), .ZN(P2_U3039) );
  INV_X1 U19909 ( .A(n16773), .ZN(n16778) );
  NAND2_X1 U19910 ( .A1(n16775), .A2(n16774), .ZN(n16777) );
  AOI21_X1 U19911 ( .B1(n16778), .B2(n16777), .A(n16776), .ZN(n16781) );
  NAND2_X1 U19912 ( .A1(n16779), .A2(n19956), .ZN(n16780) );
  OAI211_X1 U19913 ( .C1(n19872), .C2(n16782), .A(n16781), .B(n16780), .ZN(
        n16783) );
  AOI21_X1 U19914 ( .B1(n16784), .B2(n16799), .A(n16783), .ZN(n16785) );
  OAI21_X1 U19915 ( .B1(n16802), .B2(n16786), .A(n16785), .ZN(P2_U3040) );
  NAND2_X1 U19916 ( .A1(n16787), .A2(n19967), .ZN(n16796) );
  INV_X1 U19917 ( .A(n16788), .ZN(n16794) );
  AOI211_X1 U19918 ( .C1(n16792), .C2(n16791), .A(n16790), .B(n16789), .ZN(
        n16793) );
  AOI211_X1 U19919 ( .C1(n16810), .C2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n16794), .B(n16793), .ZN(n16795) );
  OAI211_X1 U19920 ( .C1(n17237), .C2(n16797), .A(n16796), .B(n16795), .ZN(
        n16798) );
  AOI21_X1 U19921 ( .B1(n16800), .B2(n16799), .A(n16798), .ZN(n16801) );
  OAI21_X1 U19922 ( .B1(n16803), .B2(n16802), .A(n16801), .ZN(P2_U3041) );
  NAND2_X1 U19923 ( .A1(n16805), .A2(n16804), .ZN(n16806) );
  XNOR2_X1 U19924 ( .A(n16806), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19946) );
  INV_X1 U19925 ( .A(n19946), .ZN(n16817) );
  INV_X1 U19926 ( .A(n16807), .ZN(n16808) );
  XNOR2_X1 U19927 ( .A(n9651), .B(n16808), .ZN(n19944) );
  NAND2_X1 U19928 ( .A1(n19944), .A2(n19958), .ZN(n16816) );
  OAI22_X1 U19929 ( .A1(n16809), .A2(n17237), .B1(n11319), .B2(n16491), .ZN(
        n16813) );
  MUX2_X1 U19930 ( .A(n16811), .B(n16810), .S(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n16812) );
  AOI211_X1 U19931 ( .C1(n16814), .C2(n19967), .A(n16813), .B(n16812), .ZN(
        n16815) );
  OAI211_X1 U19932 ( .C1(n16817), .C2(n19970), .A(n16816), .B(n16815), .ZN(
        P2_U3042) );
  INV_X1 U19933 ( .A(n17251), .ZN(n16863) );
  INV_X1 U19934 ( .A(n20631), .ZN(n20538) );
  INV_X1 U19935 ( .A(n16830), .ZN(n16862) );
  INV_X1 U19936 ( .A(n11480), .ZN(n16820) );
  NAND2_X1 U19937 ( .A1(n16820), .A2(n16819), .ZN(n16836) );
  MUX2_X1 U19938 ( .A(n16855), .B(n16836), .S(n16821), .Z(n16822) );
  AOI21_X1 U19939 ( .B1(n13581), .B2(n16862), .A(n16822), .ZN(n16938) );
  INV_X1 U19940 ( .A(n16823), .ZN(n16824) );
  MUX2_X1 U19941 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n16824), .S(
        n19866), .Z(n16829) );
  OAI222_X1 U19942 ( .A1(n16863), .A2(n16826), .B1(n20538), .B2(n16938), .C1(
        n16825), .C2(n16829), .ZN(n16827) );
  MUX2_X1 U19943 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n16827), .S(
        n16865), .Z(P2_U3601) );
  OAI21_X1 U19944 ( .B1(n19866), .B2(n19963), .A(n16828), .ZN(n16845) );
  NAND2_X1 U19945 ( .A1(n16829), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16847) );
  OR2_X1 U19946 ( .A1(n16831), .A2(n16830), .ZN(n16838) );
  INV_X1 U19947 ( .A(n16832), .ZN(n16834) );
  INV_X1 U19948 ( .A(n10566), .ZN(n16833) );
  NAND2_X1 U19949 ( .A1(n16834), .A2(n16833), .ZN(n16835) );
  AOI22_X1 U19950 ( .A1(n16836), .A2(n16835), .B1(n16855), .B2(n21312), .ZN(
        n16837) );
  NAND2_X1 U19951 ( .A1(n16838), .A2(n16837), .ZN(n16942) );
  INV_X1 U19952 ( .A(n16942), .ZN(n16839) );
  OAI222_X1 U19953 ( .A1(n16845), .A2(n16847), .B1(n20538), .B2(n16839), .C1(
        n16863), .C2(n20655), .ZN(n16840) );
  MUX2_X1 U19954 ( .A(n21340), .B(n16840), .S(n16865), .Z(P2_U3600) );
  NOR2_X1 U19955 ( .A1(n16926), .A2(n16924), .ZN(n16858) );
  NOR2_X1 U19956 ( .A1(n10567), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16857) );
  NOR2_X1 U19957 ( .A1(n16857), .A2(n16854), .ZN(n16843) );
  AOI22_X1 U19958 ( .A1(n16850), .A2(n16843), .B1(n16855), .B2(n16841), .ZN(
        n16842) );
  OAI21_X1 U19959 ( .B1(n16858), .B2(n16843), .A(n16842), .ZN(n16844) );
  AOI21_X1 U19960 ( .B1(n13766), .B2(n16862), .A(n16844), .ZN(n16939) );
  INV_X1 U19961 ( .A(n16845), .ZN(n16846) );
  OAI222_X1 U19962 ( .A1(n16848), .A2(n16863), .B1(n20538), .B2(n16939), .C1(
        n16847), .C2(n16846), .ZN(n16849) );
  MUX2_X1 U19963 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16849), .S(
        n16865), .Z(P2_U3599) );
  INV_X1 U19964 ( .A(n16850), .ZN(n16853) );
  INV_X1 U19965 ( .A(n11138), .ZN(n16851) );
  AOI21_X1 U19966 ( .B1(n16855), .B2(n16851), .A(n16857), .ZN(n16852) );
  OAI21_X1 U19967 ( .B1(n16853), .B2(n16854), .A(n16852), .ZN(n16860) );
  AOI21_X1 U19968 ( .B1(n16855), .B2(n11138), .A(n16854), .ZN(n16856) );
  OAI21_X1 U19969 ( .B1(n16858), .B2(n16857), .A(n16856), .ZN(n16859) );
  MUX2_X1 U19970 ( .A(n16860), .B(n16859), .S(n10750), .Z(n16861) );
  AOI21_X1 U19971 ( .B1(n16008), .B2(n16862), .A(n16861), .ZN(n16919) );
  OAI22_X1 U19972 ( .A1(n16864), .A2(n16863), .B1(n16919), .B2(n20538), .ZN(
        n16866) );
  MUX2_X1 U19973 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16866), .S(
        n16865), .Z(P2_U3596) );
  NOR3_X1 U19974 ( .A1(n10554), .A2(n20030), .A3(n20628), .ZN(n16867) );
  AND2_X1 U19975 ( .A1(n20634), .A2(n20687), .ZN(n20632) );
  NOR2_X1 U19976 ( .A1(n16867), .A2(n20632), .ZN(n16880) );
  INV_X1 U19977 ( .A(n16880), .ZN(n16871) );
  INV_X1 U19978 ( .A(n16868), .ZN(n16869) );
  AND2_X1 U19979 ( .A1(n16869), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20478) );
  NAND2_X1 U19980 ( .A1(n20643), .A2(n20651), .ZN(n20064) );
  NOR2_X1 U19981 ( .A1(n20212), .A2(n20064), .ZN(n19999) );
  NOR2_X1 U19982 ( .A1(n20478), .A2(n19999), .ZN(n16879) );
  INV_X1 U19983 ( .A(n20476), .ZN(n20182) );
  AOI211_X1 U19984 ( .C1(n16877), .C2(n20276), .A(n20634), .B(n19999), .ZN(
        n16870) );
  INV_X1 U19985 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16884) );
  AOI22_X1 U19986 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20002), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n20001), .ZN(n20482) );
  AOI22_X1 U19987 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20002), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20001), .ZN(n20421) );
  INV_X1 U19988 ( .A(n20030), .ZN(n16875) );
  INV_X1 U19989 ( .A(n20407), .ZN(n20468) );
  INV_X1 U19990 ( .A(n19999), .ZN(n16874) );
  OAI22_X1 U19991 ( .A1(n20421), .A2(n16875), .B1(n20468), .B2(n16874), .ZN(
        n16876) );
  AOI21_X1 U19992 ( .B1(n10554), .B2(n20408), .A(n16876), .ZN(n16883) );
  OAI21_X1 U19993 ( .B1(n16877), .B2(n19999), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16878) );
  NAND2_X1 U19994 ( .A1(n20003), .A2(n20418), .ZN(n16882) );
  OAI211_X1 U19995 ( .C1(n20006), .C2(n16884), .A(n16883), .B(n16882), .ZN(
        P2_U3048) );
  AOI21_X1 U19996 ( .B1(n16890), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n16889) );
  NOR2_X1 U19997 ( .A1(n20113), .A2(n20212), .ZN(n20107) );
  OAI21_X1 U19998 ( .B1(n20089), .B2(n20134), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n16887) );
  OR2_X1 U19999 ( .A1(n16885), .A2(n20149), .ZN(n20352) );
  INV_X1 U20000 ( .A(n20352), .ZN(n16886) );
  NAND2_X1 U20001 ( .A1(n16886), .A2(n20643), .ZN(n16893) );
  AOI21_X1 U20002 ( .B1(n16887), .B2(n16893), .A(n20182), .ZN(n16888) );
  INV_X1 U20003 ( .A(n20109), .ZN(n16899) );
  INV_X1 U20004 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16898) );
  INV_X1 U20005 ( .A(n16890), .ZN(n16891) );
  OAI21_X1 U20006 ( .B1(n16891), .B2(n20107), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16892) );
  INV_X1 U20007 ( .A(n20107), .ZN(n16895) );
  AOI22_X1 U20008 ( .A1(n20134), .A2(n20479), .B1(n20089), .B2(n20408), .ZN(
        n16894) );
  OAI21_X1 U20009 ( .B1(n20468), .B2(n16895), .A(n16894), .ZN(n16896) );
  AOI21_X1 U20010 ( .B1(n20108), .B2(n20418), .A(n16896), .ZN(n16897) );
  OAI21_X1 U20011 ( .B1(n16899), .B2(n16898), .A(n16897), .ZN(P2_U3080) );
  INV_X1 U20012 ( .A(n20114), .ZN(n16900) );
  NAND2_X1 U20013 ( .A1(n20472), .A2(n16900), .ZN(n16901) );
  NAND3_X1 U20014 ( .A1(n20660), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20346) );
  NAND2_X1 U20015 ( .A1(n16901), .A2(n20346), .ZN(n16906) );
  NOR2_X1 U20016 ( .A1(n20667), .A2(n20346), .ZN(n20410) );
  INV_X1 U20017 ( .A(n20410), .ZN(n20396) );
  NAND2_X1 U20018 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20396), .ZN(n16902) );
  OAI211_X1 U20019 ( .C1(n20410), .C2(n20276), .A(n16909), .B(n20476), .ZN(
        n16904) );
  INV_X1 U20020 ( .A(n16904), .ZN(n16905) );
  INV_X1 U20021 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16912) );
  AOI22_X1 U20022 ( .A1(n10553), .A2(n20479), .B1(n20400), .B2(n20408), .ZN(
        n16911) );
  OAI21_X1 U20023 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20346), .A(n20463), 
        .ZN(n16908) );
  NAND2_X1 U20024 ( .A1(n16909), .A2(n16908), .ZN(n20397) );
  INV_X1 U20025 ( .A(n20397), .ZN(n16915) );
  AOI22_X1 U20026 ( .A1(n16915), .A2(n20418), .B1(n20407), .B2(n20410), .ZN(
        n16910) );
  OAI211_X1 U20027 ( .C1(n20404), .C2(n16912), .A(n16911), .B(n16910), .ZN(
        P2_U3152) );
  INV_X1 U20028 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16918) );
  AOI22_X1 U20029 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20002), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20001), .ZN(n20439) );
  AOI22_X1 U20030 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n20001), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n20002), .ZN(n20503) );
  INV_X1 U20031 ( .A(n20503), .ZN(n20435) );
  AOI22_X1 U20032 ( .A1(n10553), .A2(n20500), .B1(n20400), .B2(n20435), .ZN(
        n16917) );
  AND2_X1 U20033 ( .A1(n16914), .A2(n19998), .ZN(n20434) );
  AOI22_X1 U20034 ( .A1(n16915), .A2(n20436), .B1(n20410), .B2(n20434), .ZN(
        n16916) );
  OAI211_X1 U20035 ( .C1(n20404), .C2(n16918), .A(n16917), .B(n16916), .ZN(
        P2_U3155) );
  MUX2_X1 U20036 ( .A(n10750), .B(n16919), .S(n16936), .Z(n16945) );
  MUX2_X1 U20037 ( .A(n16920), .B(n16939), .S(n16936), .Z(n16949) );
  NOR2_X1 U20038 ( .A1(n16945), .A2(n16949), .ZN(n16957) );
  NOR2_X1 U20039 ( .A1(n16936), .A2(n16921), .ZN(n16956) );
  AOI22_X1 U20040 ( .A1(n16925), .A2(n16924), .B1(n16923), .B2(n16922), .ZN(
        n16929) );
  NAND2_X1 U20041 ( .A1(n16927), .A2(n16926), .ZN(n16928) );
  NAND2_X1 U20042 ( .A1(n16929), .A2(n16928), .ZN(n20671) );
  NAND3_X1 U20043 ( .A1(n16932), .A2(n16931), .A3(n16930), .ZN(n16933) );
  NOR2_X1 U20044 ( .A1(n16934), .A2(n16933), .ZN(n19724) );
  OAI21_X1 U20045 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n19724), .ZN(n16954) );
  NAND2_X1 U20046 ( .A1(n16935), .A2(n10784), .ZN(n16953) );
  INV_X1 U20047 ( .A(n16945), .ZN(n16947) );
  AOI21_X1 U20048 ( .B1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n16938), .A(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n16943) );
  INV_X1 U20049 ( .A(n16936), .ZN(n16937) );
  AOI21_X1 U20050 ( .B1(n20313), .B2(n16938), .A(n16937), .ZN(n16941) );
  NAND2_X1 U20051 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16939), .ZN(
        n16940) );
  OAI211_X1 U20052 ( .C1(n16943), .C2(n16942), .A(n16941), .B(n16940), .ZN(
        n16944) );
  OAI21_X1 U20053 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16945), .A(
        n16944), .ZN(n16946) );
  OAI21_X1 U20054 ( .B1(n16947), .B2(n20643), .A(n16946), .ZN(n16948) );
  OAI21_X1 U20055 ( .B1(n16949), .B2(n20064), .A(n16948), .ZN(n16950) );
  NAND2_X1 U20056 ( .A1(n17144), .A2(n16950), .ZN(n16952) );
  NAND4_X1 U20057 ( .A1(n16954), .A2(n16953), .A3(n16952), .A4(n16951), .ZN(
        n16955) );
  NAND3_X1 U20058 ( .A1(n17255), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n16825), 
        .ZN(n16964) );
  NOR3_X1 U20059 ( .A1(n16960), .A2(n16959), .A3(n16958), .ZN(n16961) );
  INV_X1 U20060 ( .A(n20537), .ZN(n20540) );
  OAI211_X1 U20061 ( .C1(n20540), .C2(n20276), .A(n17143), .B(n16965), .ZN(
        P2_U3593) );
  INV_X1 U20062 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n21333) );
  INV_X1 U20063 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17599) );
  INV_X1 U20064 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17618) );
  INV_X1 U20065 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17644) );
  INV_X1 U20066 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17667) );
  INV_X1 U20067 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n18057) );
  INV_X1 U20068 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n18088) );
  NAND3_X1 U20069 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n18087) );
  NAND3_X1 U20070 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .ZN(n17807) );
  INV_X1 U20071 ( .A(n17855), .ZN(n17858) );
  NAND2_X1 U20072 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17858), .ZN(n17040) );
  INV_X1 U20073 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n17806) );
  INV_X1 U20074 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17805) );
  NOR2_X1 U20075 ( .A1(n18106), .A2(n17848), .ZN(n17849) );
  AOI22_X1 U20076 ( .A1(n18038), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16971) );
  AOI22_X1 U20077 ( .A1(n18046), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16970) );
  AOI22_X1 U20078 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17830), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16969) );
  AOI22_X1 U20079 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13253), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16968) );
  NAND4_X1 U20080 ( .A1(n16971), .A2(n16970), .A3(n16969), .A4(n16968), .ZN(
        n16977) );
  AOI22_X1 U20081 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18064), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16975) );
  AOI22_X1 U20082 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18001), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16974) );
  AOI22_X1 U20083 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18062), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16973) );
  AOI22_X1 U20084 ( .A1(n17946), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18044), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16972) );
  NAND4_X1 U20085 ( .A1(n16975), .A2(n16974), .A3(n16973), .A4(n16972), .ZN(
        n16976) );
  NOR2_X1 U20086 ( .A1(n16977), .A2(n16976), .ZN(n17844) );
  AOI22_X1 U20087 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18064), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16981) );
  AOI22_X1 U20088 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17830), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16980) );
  AOI22_X1 U20089 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n9587), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16979) );
  AOI22_X1 U20090 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16978) );
  NAND4_X1 U20091 ( .A1(n16981), .A2(n16980), .A3(n16979), .A4(n16978), .ZN(
        n16987) );
  AOI22_X1 U20092 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18038), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16985) );
  AOI22_X1 U20093 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16984) );
  AOI22_X1 U20094 ( .A1(n17946), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16983) );
  AOI22_X1 U20095 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16982) );
  NAND4_X1 U20096 ( .A1(n16985), .A2(n16984), .A3(n16983), .A4(n16982), .ZN(
        n16986) );
  NOR2_X1 U20097 ( .A1(n16987), .A2(n16986), .ZN(n17856) );
  AOI22_X1 U20098 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18044), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16991) );
  AOI22_X1 U20099 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n18065), .ZN(n16990) );
  AOI22_X1 U20100 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n9594), .ZN(n16989) );
  AOI22_X1 U20101 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18010), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n9587), .ZN(n16988) );
  NAND4_X1 U20102 ( .A1(n16991), .A2(n16990), .A3(n16989), .A4(n16988), .ZN(
        n16997) );
  AOI22_X1 U20103 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17960), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n18064), .ZN(n16995) );
  AOI22_X1 U20104 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9588), .B1(
        n17945), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16994) );
  AOI22_X1 U20105 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18001), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n18062), .ZN(n16993) );
  AOI22_X1 U20106 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n9590), .B1(
        n17946), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16992) );
  NAND4_X1 U20107 ( .A1(n16995), .A2(n16994), .A3(n16993), .A4(n16992), .ZN(
        n16996) );
  NOR2_X1 U20108 ( .A1(n16997), .A2(n16996), .ZN(n17865) );
  AOI22_X1 U20109 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18064), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17008) );
  AOI22_X1 U20110 ( .A1(n18038), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17007) );
  AOI22_X1 U20111 ( .A1(n18044), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16998) );
  OAI21_X1 U20112 ( .B1(n13197), .B2(n18061), .A(n16998), .ZN(n17005) );
  AOI22_X1 U20113 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18062), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U20114 ( .A1(n17946), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18059), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17002) );
  AOI22_X1 U20115 ( .A1(n18065), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17001) );
  AOI22_X1 U20116 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17000) );
  NAND4_X1 U20117 ( .A1(n17003), .A2(n17002), .A3(n17001), .A4(n17000), .ZN(
        n17004) );
  AOI211_X1 U20118 ( .C1(n9590), .C2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n17005), .B(n17004), .ZN(n17006) );
  NAND3_X1 U20119 ( .A1(n17008), .A2(n17007), .A3(n17006), .ZN(n17869) );
  AOI22_X1 U20120 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18064), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17018) );
  AOI22_X1 U20121 ( .A1(n18065), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17017) );
  INV_X1 U20122 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18078) );
  AOI22_X1 U20123 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18044), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17009) );
  OAI21_X1 U20124 ( .B1(n9584), .B2(n18078), .A(n17009), .ZN(n17015) );
  AOI22_X1 U20125 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17013) );
  AOI22_X1 U20126 ( .A1(n13081), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17012) );
  AOI22_X1 U20127 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17011) );
  AOI22_X1 U20128 ( .A1(n17946), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17010) );
  NAND4_X1 U20129 ( .A1(n17013), .A2(n17012), .A3(n17011), .A4(n17010), .ZN(
        n17014) );
  AOI211_X1 U20130 ( .C1(n18043), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n17015), .B(n17014), .ZN(n17016) );
  NAND3_X1 U20131 ( .A1(n17018), .A2(n17017), .A3(n17016), .ZN(n17870) );
  NAND2_X1 U20132 ( .A1(n17869), .A2(n17870), .ZN(n17868) );
  NOR2_X1 U20133 ( .A1(n17865), .A2(n17868), .ZN(n17861) );
  AOI22_X1 U20134 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20135 ( .A1(n17960), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17027) );
  AOI22_X1 U20136 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n9594), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17019) );
  OAI21_X1 U20137 ( .B1(n13197), .B2(n18100), .A(n17019), .ZN(n17025) );
  AOI22_X1 U20138 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17023) );
  AOI22_X1 U20139 ( .A1(n18044), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18064), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17022) );
  AOI22_X1 U20140 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18062), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17021) );
  AOI22_X1 U20141 ( .A1(n18065), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17020) );
  NAND4_X1 U20142 ( .A1(n17023), .A2(n17022), .A3(n17021), .A4(n17020), .ZN(
        n17024) );
  AOI211_X1 U20143 ( .C1(n18018), .C2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n17025), .B(n17024), .ZN(n17026) );
  NAND3_X1 U20144 ( .A1(n17028), .A2(n17027), .A3(n17026), .ZN(n17860) );
  NAND2_X1 U20145 ( .A1(n17861), .A2(n17860), .ZN(n17859) );
  NOR2_X1 U20146 ( .A1(n17856), .A2(n17859), .ZN(n17853) );
  AOI22_X1 U20147 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17830), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20148 ( .A1(n18044), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17037) );
  AOI22_X1 U20149 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17029) );
  OAI21_X1 U20150 ( .B1(n13197), .B2(n18092), .A(n17029), .ZN(n17035) );
  AOI22_X1 U20151 ( .A1(n18063), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U20152 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17032) );
  AOI22_X1 U20153 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9587), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17031) );
  AOI22_X1 U20154 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18038), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17030) );
  NAND4_X1 U20155 ( .A1(n17033), .A2(n17032), .A3(n17031), .A4(n17030), .ZN(
        n17034) );
  AOI211_X1 U20156 ( .C1(n18062), .C2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n17035), .B(n17034), .ZN(n17036) );
  NAND3_X1 U20157 ( .A1(n17038), .A2(n17037), .A3(n17036), .ZN(n17852) );
  NAND2_X1 U20158 ( .A1(n17853), .A2(n17852), .ZN(n17851) );
  XOR2_X1 U20159 ( .A(n17844), .B(n17851), .Z(n18122) );
  AOI22_X1 U20160 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17849), .B1(n18106), 
        .B2(n18122), .ZN(n17039) );
  OAI21_X1 U20161 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17040), .A(n17039), .ZN(
        P3_U2675) );
  AOI22_X1 U20162 ( .A1(n18063), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18062), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17052) );
  AOI22_X1 U20163 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18001), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17051) );
  INV_X1 U20164 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18086) );
  AOI22_X1 U20165 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17960), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17042) );
  OAI21_X1 U20166 ( .B1(n9592), .B2(n18086), .A(n17042), .ZN(n17049) );
  AOI22_X1 U20167 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18064), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17047) );
  AOI22_X1 U20168 ( .A1(n18065), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17046) );
  AOI22_X1 U20169 ( .A1(n17043), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17824), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17045) );
  AOI22_X1 U20170 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17044) );
  NAND4_X1 U20171 ( .A1(n17047), .A2(n17046), .A3(n17045), .A4(n17044), .ZN(
        n17048) );
  AOI211_X1 U20172 ( .C1(n17961), .C2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n17049), .B(n17048), .ZN(n17050) );
  NAND3_X1 U20173 ( .A1(n17052), .A2(n17051), .A3(n17050), .ZN(n18199) );
  INV_X1 U20174 ( .A(n18199), .ZN(n17055) );
  OAI21_X1 U20175 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17053), .A(n17983), .ZN(
        n17054) );
  AOI22_X1 U20176 ( .A1(n18106), .A2(n17055), .B1(n17054), .B2(n18101), .ZN(
        P3_U2690) );
  NAND2_X1 U20177 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19194) );
  AOI221_X1 U20178 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19194), .C1(n17057), 
        .C2(n19194), .A(n17056), .ZN(n19051) );
  NOR2_X1 U20179 ( .A1(n17058), .A2(n21428), .ZN(n17059) );
  OAI21_X1 U20180 ( .B1(n17059), .B2(n19108), .A(n19052), .ZN(n19049) );
  AOI22_X1 U20181 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19051), .B1(
        n19049), .B2(n19514), .ZN(P3_U2865) );
  NOR2_X1 U20182 ( .A1(n17061), .A2(n17060), .ZN(n17069) );
  NAND2_X1 U20183 ( .A1(n17063), .A2(n19702), .ZN(n17067) );
  NOR2_X1 U20184 ( .A1(n19691), .A2(n18305), .ZN(n19539) );
  OAI21_X1 U20185 ( .B1(n17065), .B2(n19539), .A(n19690), .ZN(n18255) );
  OAI21_X1 U20186 ( .B1(n17067), .B2(n18255), .A(n17066), .ZN(n17068) );
  NOR3_X1 U20187 ( .A1(n17069), .A2(n17147), .A3(n17068), .ZN(n19513) );
  INV_X1 U20188 ( .A(n19513), .ZN(n19534) );
  NOR2_X1 U20189 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19650), .ZN(n19055) );
  INV_X1 U20190 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n19047) );
  NOR2_X1 U20191 ( .A1(n19047), .A2(n19648), .ZN(n17070) );
  INV_X1 U20192 ( .A(n19659), .ZN(n19673) );
  AOI21_X1 U20193 ( .B1(n19493), .B2(n21439), .A(n17416), .ZN(n19530) );
  NAND3_X1 U20194 ( .A1(n19675), .A2(n19673), .A3(n19530), .ZN(n17071) );
  OAI21_X1 U20195 ( .B1(n19675), .B2(n21439), .A(n17071), .ZN(P3_U3284) );
  OAI21_X1 U20196 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n17073), .A(
        n17072), .ZN(n17285) );
  INV_X1 U20197 ( .A(n18929), .ZN(n18848) );
  AOI21_X1 U20198 ( .B1(n18848), .B2(n18734), .A(n17074), .ZN(n17289) );
  NAND2_X1 U20199 ( .A1(n19031), .A2(n18367), .ZN(n17075) );
  OAI211_X1 U20200 ( .C1(n17289), .C2(n19026), .A(n17137), .B(n17075), .ZN(
        n17076) );
  AOI22_X1 U20201 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n17076), .B1(
        n9586), .B2(P3_REIP_REG_29__SCAN_IN), .ZN(n17079) );
  NAND2_X1 U20202 ( .A1(n18222), .A2(n19525), .ZN(n18910) );
  NAND2_X1 U20203 ( .A1(n18893), .A2(n18786), .ZN(n17077) );
  OAI211_X1 U20204 ( .C1(n18532), .C2(n18910), .A(n18749), .B(n17077), .ZN(
        n18791) );
  NAND2_X1 U20205 ( .A1(n19037), .A2(n18791), .ZN(n18761) );
  NOR2_X1 U20206 ( .A1(n17262), .A2(n18761), .ZN(n18736) );
  INV_X1 U20207 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17269) );
  NAND3_X1 U20208 ( .A1(n17279), .A2(n18736), .A3(n17269), .ZN(n17078) );
  OAI211_X1 U20209 ( .C1(n17285), .C2(n18935), .A(n17079), .B(n17078), .ZN(
        P3_U2833) );
  OR2_X1 U20210 ( .A1(n17081), .A2(n17080), .ZN(n17088) );
  INV_X1 U20211 ( .A(n17082), .ZN(n17083) );
  AOI21_X1 U20212 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n17084), .A(
        n17083), .ZN(n17085) );
  AOI22_X1 U20213 ( .A1(n17088), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n17085), .B2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n17086) );
  INV_X1 U20214 ( .A(n17086), .ZN(n17087) );
  OAI21_X1 U20215 ( .B1(n17088), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n17087), .ZN(n17092) );
  OAI22_X1 U20216 ( .A1(n17092), .A2(n17091), .B1(n17089), .B2(n17093), .ZN(
        n17096) );
  AOI21_X1 U20217 ( .B1(n17092), .B2(n17091), .A(n17090), .ZN(n17095) );
  INV_X1 U20218 ( .A(n17093), .ZN(n17094) );
  OAI22_X1 U20219 ( .A1(n17096), .A2(n17095), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n17094), .ZN(n17118) );
  INV_X1 U20220 ( .A(n17097), .ZN(n17104) );
  NAND3_X1 U20221 ( .A1(n17112), .A2(n17099), .A3(n17098), .ZN(n17100) );
  MUX2_X1 U20222 ( .A(n17101), .B(n17100), .S(n17107), .Z(n17102) );
  AOI21_X1 U20223 ( .B1(n17104), .B2(n17103), .A(n17102), .ZN(n21307) );
  OR2_X1 U20224 ( .A1(n17106), .A2(n17105), .ZN(n17111) );
  INV_X1 U20225 ( .A(n17107), .ZN(n17110) );
  OAI22_X1 U20226 ( .A1(n17110), .A2(n17109), .B1(n10051), .B2(n17108), .ZN(
        n20704) );
  AOI21_X1 U20227 ( .B1(n17215), .B2(n17111), .A(n20704), .ZN(n20711) );
  INV_X1 U20228 ( .A(n17112), .ZN(n17113) );
  AOI221_X1 U20229 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(n20711), .C1(
        P1_MORE_REG_SCAN_IN), .C2(n20711), .A(n17113), .ZN(n17114) );
  NAND3_X1 U20230 ( .A1(n17115), .A2(n21307), .A3(n17114), .ZN(n17116) );
  AOI211_X1 U20231 ( .C1(n17118), .C2(n20942), .A(n17117), .B(n17116), .ZN(
        n17132) );
  INV_X1 U20232 ( .A(n17132), .ZN(n17125) );
  INV_X1 U20233 ( .A(n17119), .ZN(n17123) );
  OR3_X1 U20234 ( .A1(n17121), .A2(n17142), .A3(n17120), .ZN(n17122) );
  OAI221_X1 U20235 ( .B1(n17124), .B2(n17123), .C1(n17124), .C2(n21212), .A(
        n17122), .ZN(n17220) );
  AOI221_X1 U20236 ( .B1(n11759), .B2(n17222), .C1(n17125), .C2(n17222), .A(
        n17220), .ZN(n17127) );
  NOR2_X1 U20237 ( .A1(n17127), .A2(n11759), .ZN(n21205) );
  OAI211_X1 U20238 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n17215), .A(n21205), 
        .B(n17126), .ZN(n17221) );
  AOI21_X1 U20239 ( .B1(n17128), .B2(n21290), .A(n17127), .ZN(n17129) );
  OAI22_X1 U20240 ( .A1(n17130), .A2(n17221), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n17129), .ZN(n17131) );
  OAI21_X1 U20241 ( .B1(n17132), .B2(n20710), .A(n17131), .ZN(P1_U3161) );
  NOR2_X1 U20242 ( .A1(n17134), .A2(n17133), .ZN(n17135) );
  XNOR2_X1 U20243 ( .A(n17135), .B(n21367), .ZN(n17267) );
  NOR2_X1 U20244 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17136), .ZN(
        n17263) );
  AOI21_X1 U20245 ( .B1(n17138), .B2(n17137), .A(n21367), .ZN(n17139) );
  AOI21_X1 U20246 ( .B1(n18736), .B2(n17263), .A(n17139), .ZN(n17140) );
  NAND2_X1 U20247 ( .A1(n9586), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n17256) );
  OAI211_X1 U20248 ( .C1(n17267), .C2(n18935), .A(n17140), .B(n17256), .ZN(
        P3_U2832) );
  INV_X1 U20249 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21206) );
  NOR2_X1 U20250 ( .A1(n21206), .A2(n21217), .ZN(n21211) );
  INV_X1 U20251 ( .A(HOLD), .ZN(n20556) );
  NOR2_X1 U20252 ( .A1(n20702), .A2(n20556), .ZN(n21209) );
  NAND2_X1 U20253 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n21207) );
  OAI21_X1 U20254 ( .B1(n21211), .B2(n21209), .A(n21207), .ZN(n17141) );
  OAI211_X1 U20255 ( .C1(n17215), .C2(n20702), .A(n17142), .B(n17141), .ZN(
        P1_U3195) );
  AND2_X1 U20256 ( .A1(n20814), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  OAI221_X1 U20257 ( .B1(n11140), .B2(n17143), .C1(n20672), .C2(n17143), .A(
        n20182), .ZN(n20665) );
  NOR2_X1 U20258 ( .A1(n17144), .A2(n20665), .ZN(P2_U3047) );
  NAND2_X1 U20259 ( .A1(n17148), .A2(n10207), .ZN(n18245) );
  AOI22_X1 U20260 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18249), .B1(
        P3_EAX_REG_0__SCAN_IN), .B2(n18250), .ZN(n17150) );
  NAND2_X1 U20261 ( .A1(n19084), .A2(n10207), .ZN(n18246) );
  NOR2_X1 U20262 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18246), .ZN(n18251) );
  INV_X1 U20263 ( .A(n18251), .ZN(n17149) );
  OAI211_X1 U20264 ( .C1(n13297), .C2(n18237), .A(n17150), .B(n17149), .ZN(
        P3_U2735) );
  INV_X1 U20265 ( .A(n17151), .ZN(n17152) );
  OAI22_X1 U20266 ( .A1(n17153), .A2(n21238), .B1(n20780), .B2(n17152), .ZN(
        n17154) );
  AOI211_X1 U20267 ( .C1(n20785), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20772), .B(n17154), .ZN(n17164) );
  INV_X1 U20268 ( .A(n17155), .ZN(n17159) );
  INV_X1 U20269 ( .A(n17156), .ZN(n17158) );
  AOI22_X1 U20270 ( .A1(n17159), .A2(n12954), .B1(n17158), .B2(n17157), .ZN(
        n17163) );
  NAND3_X1 U20271 ( .A1(n17160), .A2(P1_REIP_REG_9__SCAN_IN), .A3(n21238), 
        .ZN(n17162) );
  NAND2_X1 U20272 ( .A1(n20757), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n17161) );
  NAND4_X1 U20273 ( .A1(n17164), .A2(n17163), .A3(n17162), .A4(n17161), .ZN(
        P1_U2830) );
  AOI22_X1 U20274 ( .A1(n20882), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20916), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n17170) );
  INV_X1 U20275 ( .A(n17165), .ZN(n17166) );
  AOI21_X1 U20276 ( .B1(n17168), .B2(n17167), .A(n17166), .ZN(n17193) );
  AOI22_X1 U20277 ( .A1(n17193), .A2(n20887), .B1(n20884), .B2(n20737), .ZN(
        n17169) );
  OAI211_X1 U20278 ( .C1(n20881), .C2(n20739), .A(n17170), .B(n17169), .ZN(
        P1_U2992) );
  AOI22_X1 U20279 ( .A1(n20882), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20916), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n17177) );
  NAND2_X1 U20280 ( .A1(n17172), .A2(n17171), .ZN(n17173) );
  NAND2_X1 U20281 ( .A1(n17174), .A2(n17173), .ZN(n17197) );
  INV_X1 U20282 ( .A(n20750), .ZN(n17175) );
  AOI22_X1 U20283 ( .A1(n17197), .A2(n20887), .B1(n20884), .B2(n17175), .ZN(
        n17176) );
  OAI211_X1 U20284 ( .C1(n20881), .C2(n20754), .A(n17177), .B(n17176), .ZN(
        P1_U2993) );
  AOI22_X1 U20285 ( .A1(n20882), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20916), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n17183) );
  OAI21_X1 U20286 ( .B1(n17180), .B2(n17179), .A(n17178), .ZN(n17181) );
  INV_X1 U20287 ( .A(n17181), .ZN(n17206) );
  AOI22_X1 U20288 ( .A1(n17206), .A2(n20887), .B1(n20884), .B2(n20797), .ZN(
        n17182) );
  OAI211_X1 U20289 ( .C1(n20881), .C2(n20767), .A(n17183), .B(n17182), .ZN(
        P1_U2994) );
  AOI21_X1 U20290 ( .B1(n17185), .B2(n17191), .A(n17184), .ZN(n17189) );
  AOI22_X1 U20291 ( .A1(n17187), .A2(n20922), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17186), .ZN(n17188) );
  OAI211_X1 U20292 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n17190), .A(
        n17189), .B(n17188), .ZN(P1_U3022) );
  AOI22_X1 U20293 ( .A1(n20730), .A2(n17191), .B1(n20916), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n17195) );
  AOI22_X1 U20294 ( .A1(n17193), .A2(n20922), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17192), .ZN(n17194) );
  OAI211_X1 U20295 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n17196), .A(
        n17195), .B(n17194), .ZN(P1_U3024) );
  AOI222_X1 U20296 ( .A1(n17197), .A2(n20922), .B1(n17191), .B2(n20746), .C1(
        P1_REIP_REG_6__SCAN_IN), .C2(n20916), .ZN(n17198) );
  OAI221_X1 U20297 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17200), .C1(
        n21388), .C2(n17199), .A(n17198), .ZN(P1_U3025) );
  INV_X1 U20298 ( .A(n17201), .ZN(n17209) );
  INV_X1 U20299 ( .A(n14175), .ZN(n17202) );
  AOI21_X1 U20300 ( .B1(n17204), .B2(n17203), .A(n17202), .ZN(n20794) );
  AOI22_X1 U20301 ( .A1(n17191), .A2(n20794), .B1(n20916), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n17208) );
  AOI22_X1 U20302 ( .A1(n17206), .A2(n20922), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17205), .ZN(n17207) );
  OAI211_X1 U20303 ( .C1(n20903), .C2(n17209), .A(n17208), .B(n17207), .ZN(
        P1_U3026) );
  OR4_X1 U20304 ( .A1(n20769), .A2(n17212), .A3(n17211), .A4(n17210), .ZN(
        n17213) );
  OAI21_X1 U20305 ( .B1(n21294), .B2(n17214), .A(n17213), .ZN(P1_U3468) );
  NAND4_X1 U20306 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n11830), .A4(n17215), .ZN(n17216) );
  AND2_X1 U20307 ( .A1(n17217), .A2(n17216), .ZN(n21204) );
  NAND2_X1 U20308 ( .A1(n21204), .A2(n17218), .ZN(n17219) );
  AOI22_X1 U20309 ( .A1(n17222), .A2(n17221), .B1(n17220), .B2(n17219), .ZN(
        P1_U3162) );
  OAI21_X1 U20310 ( .B1(n21205), .B2(n21064), .A(n17223), .ZN(P1_U3466) );
  INV_X1 U20311 ( .A(n17224), .ZN(n17234) );
  OAI21_X1 U20312 ( .B1(n17226), .B2(n17237), .A(n17225), .ZN(n17227) );
  AOI21_X1 U20313 ( .B1(n16008), .B2(n19967), .A(n17227), .ZN(n17228) );
  OAI21_X1 U20314 ( .B1(n17229), .B2(n19970), .A(n17228), .ZN(n17230) );
  AOI21_X1 U20315 ( .B1(n19958), .B2(n17231), .A(n17230), .ZN(n17232) );
  OAI221_X1 U20316 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17234), .C1(
        n10838), .C2(n17233), .A(n17232), .ZN(P2_U3043) );
  INV_X1 U20317 ( .A(n17235), .ZN(n17236) );
  OR2_X1 U20318 ( .A1(n17237), .A2(n17236), .ZN(n17238) );
  OAI21_X1 U20319 ( .B1(n19970), .B2(n17239), .A(n17238), .ZN(n17240) );
  INV_X1 U20320 ( .A(n17240), .ZN(n17246) );
  INV_X1 U20321 ( .A(n17241), .ZN(n19960) );
  OAI22_X1 U20322 ( .A1(n19960), .A2(n19964), .B1(n16802), .B2(n17242), .ZN(
        n17243) );
  AOI211_X1 U20323 ( .C1(n19967), .C2(n13581), .A(n17244), .B(n17243), .ZN(
        n17245) );
  OAI211_X1 U20324 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n19961), .A(
        n17246), .B(n17245), .ZN(P2_U3046) );
  NOR2_X1 U20325 ( .A1(n17247), .A2(n20463), .ZN(n20662) );
  OAI21_X1 U20326 ( .B1(n20537), .B2(n20662), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n17250) );
  AND3_X1 U20327 ( .A1(n17250), .A2(n17249), .A3(n17248), .ZN(n17254) );
  OAI21_X1 U20328 ( .B1(n17251), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n20695), 
        .ZN(n17252) );
  OAI21_X1 U20329 ( .B1(n20540), .B2(n20686), .A(n17252), .ZN(n17253) );
  OAI211_X1 U20330 ( .C1(n17255), .C2(n19723), .A(n17254), .B(n17253), .ZN(
        P2_U3176) );
  XOR2_X1 U20331 ( .A(n17270), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n17452) );
  OAI221_X1 U20332 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n17258), .C1(
        n10347), .C2(n17257), .A(n17256), .ZN(n17259) );
  AOI21_X1 U20333 ( .B1(n18578), .B2(n17452), .A(n17259), .ZN(n17266) );
  NAND2_X1 U20334 ( .A1(n18636), .A2(n17260), .ZN(n17268) );
  OAI21_X1 U20335 ( .B1(n17281), .B2(n18725), .A(n17268), .ZN(n17264) );
  INV_X1 U20336 ( .A(n18909), .ZN(n17261) );
  INV_X2 U20337 ( .A(n18636), .ZN(n18593) );
  OAI22_X2 U20338 ( .A1(n17261), .A2(n18725), .B1(n13337), .B2(n18593), .ZN(
        n18576) );
  NAND2_X2 U20339 ( .A1(n9603), .A2(n18576), .ZN(n18531) );
  NOR2_X1 U20340 ( .A1(n17262), .A2(n18531), .ZN(n18389) );
  AOI22_X1 U20341 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17264), .B1(
        n17263), .B2(n18389), .ZN(n17265) );
  OAI211_X1 U20342 ( .C1(n17267), .C2(n18609), .A(n17266), .B(n17265), .ZN(
        P3_U2800) );
  NAND2_X1 U20343 ( .A1(n17279), .A2(n18733), .ZN(n17291) );
  AOI21_X1 U20344 ( .B1(n17269), .B2(n17291), .A(n17268), .ZN(n17277) );
  NAND2_X1 U20345 ( .A1(n9586), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n17273) );
  AOI21_X1 U20346 ( .B1(n9749), .B2(n17459), .A(n17270), .ZN(n17458) );
  OAI21_X1 U20347 ( .B1(n18578), .B2(n17271), .A(n17458), .ZN(n17272) );
  OAI211_X1 U20348 ( .C1(n17275), .C2(n17274), .A(n17273), .B(n17272), .ZN(
        n17276) );
  AOI211_X1 U20349 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n17278), .A(
        n17277), .B(n17276), .ZN(n17284) );
  INV_X1 U20350 ( .A(n17279), .ZN(n17280) );
  NOR2_X1 U20351 ( .A1(n17280), .A2(n18731), .ZN(n17293) );
  NOR2_X1 U20352 ( .A1(n17281), .A2(n18725), .ZN(n17282) );
  OAI21_X1 U20353 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n17293), .A(
        n17282), .ZN(n17283) );
  OAI211_X1 U20354 ( .C1(n17285), .C2(n18609), .A(n17284), .B(n17283), .ZN(
        P3_U2801) );
  NOR2_X1 U20355 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18734), .ZN(
        n18369) );
  AOI22_X1 U20356 ( .A1(n9586), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n18736), 
        .B2(n18369), .ZN(n17299) );
  OAI21_X1 U20357 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18634), .A(
        n17286), .ZN(n18364) );
  OAI211_X1 U20358 ( .C1(n17288), .C2(n18382), .A(n19525), .B(n17287), .ZN(
        n17290) );
  OAI211_X1 U20359 ( .C1(n18363), .C2(n17290), .A(n17289), .B(n19027), .ZN(
        n17295) );
  INV_X1 U20360 ( .A(n18893), .ZN(n19527) );
  INV_X1 U20361 ( .A(n17291), .ZN(n17292) );
  OAI22_X1 U20362 ( .A1(n17293), .A2(n19527), .B1(n17292), .B2(n18910), .ZN(
        n17294) );
  OAI211_X1 U20363 ( .C1(n17295), .C2(n17294), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n19024), .ZN(n17298) );
  INV_X1 U20364 ( .A(n19035), .ZN(n19042) );
  NAND4_X1 U20365 ( .A1(n18634), .A2(n19042), .A3(n18365), .A4(n18367), .ZN(
        n17297) );
  NAND3_X1 U20366 ( .A1(n18960), .A2(n18381), .A3(n18364), .ZN(n17296) );
  NAND4_X1 U20367 ( .A1(n17299), .A2(n17298), .A3(n17297), .A4(n17296), .ZN(
        P3_U2834) );
  NOR3_X1 U20368 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n17301) );
  NOR4_X1 U20369 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17300) );
  INV_X2 U20370 ( .A(n17385), .ZN(U215) );
  NAND4_X1 U20371 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17301), .A3(n17300), .A4(
        U215), .ZN(U213) );
  INV_X1 U20372 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19898) );
  INV_X2 U20373 ( .A(U214), .ZN(n17352) );
  NOR2_X1 U20374 ( .A1(n17352), .A2(n17302), .ZN(n17304) );
  INV_X1 U20375 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n17387) );
  OAI222_X1 U20376 ( .A1(U212), .A2(n19898), .B1(n17354), .B2(n17303), .C1(
        U214), .C2(n17387), .ZN(U216) );
  AOI222_X1 U20377 ( .A1(n17351), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n17304), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n17352), .C2(P1_DATAO_REG_30__SCAN_IN), 
        .ZN(n17305) );
  INV_X1 U20378 ( .A(n17305), .ZN(U217) );
  AOI22_X1 U20379 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n17351), .ZN(n17306) );
  OAI21_X1 U20380 ( .B1(n15081), .B2(n17354), .A(n17306), .ZN(U218) );
  INV_X1 U20381 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n17308) );
  AOI22_X1 U20382 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17351), .ZN(n17307) );
  OAI21_X1 U20383 ( .B1(n17308), .B2(n17354), .A(n17307), .ZN(U219) );
  AOI22_X1 U20384 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n17351), .ZN(n17309) );
  OAI21_X1 U20385 ( .B1(n17310), .B2(n17354), .A(n17309), .ZN(U220) );
  AOI22_X1 U20386 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n17351), .ZN(n17311) );
  OAI21_X1 U20387 ( .B1(n17312), .B2(n17354), .A(n17311), .ZN(U221) );
  INV_X1 U20388 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n17314) );
  AOI22_X1 U20389 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n17351), .ZN(n17313) );
  OAI21_X1 U20390 ( .B1(n17314), .B2(n17354), .A(n17313), .ZN(U222) );
  AOI22_X1 U20391 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n17351), .ZN(n17315) );
  OAI21_X1 U20392 ( .B1(n16199), .B2(n17354), .A(n17315), .ZN(U223) );
  INV_X1 U20393 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n17317) );
  AOI22_X1 U20394 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17351), .ZN(n17316) );
  OAI21_X1 U20395 ( .B1(n17317), .B2(n17354), .A(n17316), .ZN(U224) );
  INV_X1 U20396 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n17319) );
  AOI22_X1 U20397 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n17351), .ZN(n17318) );
  OAI21_X1 U20398 ( .B1(n17319), .B2(n17354), .A(n17318), .ZN(U225) );
  INV_X1 U20399 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n17321) );
  AOI22_X1 U20400 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n17351), .ZN(n17320) );
  OAI21_X1 U20401 ( .B1(n17321), .B2(n17354), .A(n17320), .ZN(U226) );
  INV_X1 U20402 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n17323) );
  AOI22_X1 U20403 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n17351), .ZN(n17322) );
  OAI21_X1 U20404 ( .B1(n17323), .B2(n17354), .A(n17322), .ZN(U227) );
  INV_X1 U20405 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n17325) );
  AOI22_X1 U20406 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n17351), .ZN(n17324) );
  OAI21_X1 U20407 ( .B1(n17325), .B2(n17354), .A(n17324), .ZN(U228) );
  INV_X1 U20408 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n17327) );
  AOI22_X1 U20409 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n17351), .ZN(n17326) );
  OAI21_X1 U20410 ( .B1(n17327), .B2(n17354), .A(n17326), .ZN(U229) );
  AOI22_X1 U20411 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n17351), .ZN(n17328) );
  OAI21_X1 U20412 ( .B1(n21348), .B2(n17354), .A(n17328), .ZN(U230) );
  INV_X1 U20413 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n17329) );
  INV_X1 U20414 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n21448) );
  OAI222_X1 U20415 ( .A1(U212), .A2(n13505), .B1(n17354), .B2(n17329), .C1(
        U214), .C2(n21448), .ZN(U231) );
  AOI22_X1 U20416 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n17351), .ZN(n17330) );
  OAI21_X1 U20417 ( .B1(n13564), .B2(n17354), .A(n17330), .ZN(U232) );
  INV_X1 U20418 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n21370) );
  INV_X1 U20419 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n17331) );
  OAI222_X1 U20420 ( .A1(U212), .A2(n21370), .B1(n17354), .B2(n15071), .C1(
        U214), .C2(n17331), .ZN(U233) );
  AOI22_X1 U20421 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n17351), .ZN(n17332) );
  OAI21_X1 U20422 ( .B1(n13426), .B2(n17354), .A(n17332), .ZN(U234) );
  INV_X1 U20423 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n17368) );
  INV_X1 U20424 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n21433) );
  OAI222_X1 U20425 ( .A1(U212), .A2(n17368), .B1(n17354), .B2(n17333), .C1(
        U214), .C2(n21433), .ZN(U235) );
  AOI22_X1 U20426 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n17351), .ZN(n17334) );
  OAI21_X1 U20427 ( .B1(n13422), .B2(n17354), .A(n17334), .ZN(U236) );
  AOI22_X1 U20428 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n17351), .ZN(n17335) );
  OAI21_X1 U20429 ( .B1(n21401), .B2(n17354), .A(n17335), .ZN(U237) );
  AOI22_X1 U20430 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n17351), .ZN(n17336) );
  OAI21_X1 U20431 ( .B1(n17337), .B2(n17354), .A(n17336), .ZN(U238) );
  AOI22_X1 U20432 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n17351), .ZN(n17338) );
  OAI21_X1 U20433 ( .B1(n17339), .B2(n17354), .A(n17338), .ZN(U239) );
  AOI22_X1 U20434 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n17351), .ZN(n17340) );
  OAI21_X1 U20435 ( .B1(n13456), .B2(n17354), .A(n17340), .ZN(U240) );
  AOI22_X1 U20436 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n17351), .ZN(n17341) );
  OAI21_X1 U20437 ( .B1(n21338), .B2(n17354), .A(n17341), .ZN(U241) );
  INV_X1 U20438 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n21357) );
  AOI22_X1 U20439 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n17351), .ZN(n17342) );
  OAI21_X1 U20440 ( .B1(n21357), .B2(n17354), .A(n17342), .ZN(U242) );
  AOI22_X1 U20441 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n17351), .ZN(n17343) );
  OAI21_X1 U20442 ( .B1(n17344), .B2(n17354), .A(n17343), .ZN(U243) );
  INV_X1 U20443 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n17346) );
  AOI22_X1 U20444 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n17351), .ZN(n17345) );
  OAI21_X1 U20445 ( .B1(n17346), .B2(n17354), .A(n17345), .ZN(U244) );
  AOI22_X1 U20446 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n17351), .ZN(n17347) );
  OAI21_X1 U20447 ( .B1(n17348), .B2(n17354), .A(n17347), .ZN(U245) );
  INV_X1 U20448 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n17350) );
  AOI22_X1 U20449 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n17351), .ZN(n17349) );
  OAI21_X1 U20450 ( .B1(n17350), .B2(n17354), .A(n17349), .ZN(U246) );
  AOI22_X1 U20451 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n17352), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n17351), .ZN(n17353) );
  OAI21_X1 U20452 ( .B1(n17355), .B2(n17354), .A(n17353), .ZN(U247) );
  INV_X1 U20453 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n17356) );
  INV_X1 U20454 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n21451) );
  AOI22_X1 U20455 ( .A1(n17385), .A2(n17356), .B1(n21451), .B2(U215), .ZN(U251) );
  OAI22_X1 U20456 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n17385), .ZN(n17357) );
  INV_X1 U20457 ( .A(n17357), .ZN(U252) );
  INV_X1 U20458 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n17358) );
  INV_X1 U20459 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n21446) );
  AOI22_X1 U20460 ( .A1(n17385), .A2(n17358), .B1(n21446), .B2(U215), .ZN(U253) );
  INV_X1 U20461 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n17359) );
  INV_X1 U20462 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n19065) );
  AOI22_X1 U20463 ( .A1(n17385), .A2(n17359), .B1(n19065), .B2(U215), .ZN(U254) );
  INV_X1 U20464 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n17360) );
  INV_X1 U20465 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n19069) );
  AOI22_X1 U20466 ( .A1(n17385), .A2(n17360), .B1(n19069), .B2(U215), .ZN(U255) );
  INV_X1 U20467 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n17361) );
  INV_X1 U20468 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n19073) );
  AOI22_X1 U20469 ( .A1(n17385), .A2(n17361), .B1(n19073), .B2(U215), .ZN(U256) );
  INV_X1 U20470 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n17362) );
  INV_X1 U20471 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n19077) );
  AOI22_X1 U20472 ( .A1(n17385), .A2(n17362), .B1(n19077), .B2(U215), .ZN(U257) );
  INV_X1 U20473 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n17363) );
  INV_X1 U20474 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n19081) );
  AOI22_X1 U20475 ( .A1(n17383), .A2(n17363), .B1(n19081), .B2(U215), .ZN(U258) );
  INV_X1 U20476 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n17364) );
  INV_X1 U20477 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n18340) );
  AOI22_X1 U20478 ( .A1(n17383), .A2(n17364), .B1(n18340), .B2(U215), .ZN(U259) );
  INV_X1 U20479 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n17365) );
  INV_X1 U20480 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n18343) );
  AOI22_X1 U20481 ( .A1(n17383), .A2(n17365), .B1(n18343), .B2(U215), .ZN(U260) );
  INV_X1 U20482 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n17366) );
  INV_X1 U20483 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n18345) );
  AOI22_X1 U20484 ( .A1(n17385), .A2(n17366), .B1(n18345), .B2(U215), .ZN(U261) );
  OAI22_X1 U20485 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n17385), .ZN(n17367) );
  INV_X1 U20486 ( .A(n17367), .ZN(U262) );
  INV_X1 U20487 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n18349) );
  AOI22_X1 U20488 ( .A1(n17385), .A2(n17368), .B1(n18349), .B2(U215), .ZN(U263) );
  OAI22_X1 U20489 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n17385), .ZN(n17369) );
  INV_X1 U20490 ( .A(n17369), .ZN(U264) );
  INV_X1 U20491 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n21382) );
  AOI22_X1 U20492 ( .A1(n17383), .A2(n21370), .B1(n21382), .B2(U215), .ZN(U265) );
  OAI22_X1 U20493 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n17385), .ZN(n17370) );
  INV_X1 U20494 ( .A(n17370), .ZN(U266) );
  AOI22_X1 U20495 ( .A1(n17385), .A2(n13505), .B1(n16263), .B2(U215), .ZN(U267) );
  OAI22_X1 U20496 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17385), .ZN(n17371) );
  INV_X1 U20497 ( .A(n17371), .ZN(U268) );
  OAI22_X1 U20498 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17385), .ZN(n17372) );
  INV_X1 U20499 ( .A(n17372), .ZN(U269) );
  OAI22_X1 U20500 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17385), .ZN(n17373) );
  INV_X1 U20501 ( .A(n17373), .ZN(U270) );
  OAI22_X1 U20502 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17385), .ZN(n17374) );
  INV_X1 U20503 ( .A(n17374), .ZN(U271) );
  OAI22_X1 U20504 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17385), .ZN(n17375) );
  INV_X1 U20505 ( .A(n17375), .ZN(U272) );
  AOI22_X1 U20506 ( .A1(n17385), .A2(n13511), .B1(n16214), .B2(U215), .ZN(U273) );
  OAI22_X1 U20507 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17385), .ZN(n17377) );
  INV_X1 U20508 ( .A(n17377), .ZN(U274) );
  OAI22_X1 U20509 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17383), .ZN(n17378) );
  INV_X1 U20510 ( .A(n17378), .ZN(U275) );
  OAI22_X1 U20511 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17383), .ZN(n17379) );
  INV_X1 U20512 ( .A(n17379), .ZN(U276) );
  OAI22_X1 U20513 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17383), .ZN(n17380) );
  INV_X1 U20514 ( .A(n17380), .ZN(U277) );
  OAI22_X1 U20515 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17383), .ZN(n17381) );
  INV_X1 U20516 ( .A(n17381), .ZN(U278) );
  OAI22_X1 U20517 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17383), .ZN(n17382) );
  INV_X1 U20518 ( .A(n17382), .ZN(U279) );
  OAI22_X1 U20519 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17383), .ZN(n17384) );
  INV_X1 U20520 ( .A(n17384), .ZN(U280) );
  INV_X1 U20521 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19901) );
  AOI22_X1 U20522 ( .A1(n17385), .A2(n19901), .B1(n14696), .B2(U215), .ZN(U281) );
  OAI22_X1 U20523 ( .A1(U215), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n17385), .ZN(n17386) );
  INV_X1 U20524 ( .A(n17386), .ZN(U282) );
  INV_X1 U20525 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n18256) );
  AOI222_X1 U20526 ( .A1(n17387), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19898), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n18256), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n17388) );
  INV_X2 U20527 ( .A(n17390), .ZN(n17389) );
  INV_X1 U20528 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19594) );
  INV_X1 U20529 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20582) );
  AOI22_X1 U20530 ( .A1(n17389), .A2(n19594), .B1(n20582), .B2(n17390), .ZN(
        U347) );
  INV_X1 U20531 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19592) );
  INV_X1 U20532 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20580) );
  AOI22_X1 U20533 ( .A1(n17389), .A2(n19592), .B1(n20580), .B2(n17390), .ZN(
        U348) );
  INV_X1 U20534 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19590) );
  INV_X1 U20535 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20578) );
  AOI22_X1 U20536 ( .A1(n17389), .A2(n19590), .B1(n20578), .B2(n17390), .ZN(
        U349) );
  INV_X1 U20537 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19588) );
  INV_X1 U20538 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20577) );
  AOI22_X1 U20539 ( .A1(n17389), .A2(n19588), .B1(n20577), .B2(n17390), .ZN(
        U350) );
  INV_X1 U20540 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19586) );
  INV_X1 U20541 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20575) );
  AOI22_X1 U20542 ( .A1(n17389), .A2(n19586), .B1(n20575), .B2(n17390), .ZN(
        U351) );
  INV_X1 U20543 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19583) );
  INV_X1 U20544 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20573) );
  AOI22_X1 U20545 ( .A1(n17389), .A2(n19583), .B1(n20573), .B2(n17390), .ZN(
        U352) );
  INV_X1 U20546 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19582) );
  INV_X1 U20547 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20572) );
  AOI22_X1 U20548 ( .A1(n17389), .A2(n19582), .B1(n20572), .B2(n17390), .ZN(
        U353) );
  INV_X1 U20549 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19580) );
  AOI22_X1 U20550 ( .A1(n17389), .A2(n19580), .B1(n20570), .B2(n17390), .ZN(
        U354) );
  INV_X1 U20551 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19636) );
  INV_X1 U20552 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20617) );
  AOI22_X1 U20553 ( .A1(n17389), .A2(n19636), .B1(n20617), .B2(n17390), .ZN(
        U355) );
  INV_X1 U20554 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19633) );
  INV_X1 U20555 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20613) );
  AOI22_X1 U20556 ( .A1(n17389), .A2(n19633), .B1(n20613), .B2(n17390), .ZN(
        U356) );
  INV_X1 U20557 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19629) );
  INV_X1 U20558 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20611) );
  AOI22_X1 U20559 ( .A1(n17389), .A2(n19629), .B1(n20611), .B2(n17390), .ZN(
        U357) );
  INV_X1 U20560 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19628) );
  INV_X1 U20561 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20609) );
  AOI22_X1 U20562 ( .A1(n17389), .A2(n19628), .B1(n20609), .B2(n17390), .ZN(
        U358) );
  INV_X1 U20563 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19626) );
  INV_X1 U20564 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20608) );
  AOI22_X1 U20565 ( .A1(n17389), .A2(n19626), .B1(n20608), .B2(n17390), .ZN(
        U359) );
  INV_X1 U20566 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19625) );
  INV_X1 U20567 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20606) );
  AOI22_X1 U20568 ( .A1(n17389), .A2(n19625), .B1(n20606), .B2(n17390), .ZN(
        U360) );
  INV_X1 U20569 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19622) );
  INV_X1 U20570 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20604) );
  AOI22_X1 U20571 ( .A1(n17389), .A2(n19622), .B1(n20604), .B2(n17390), .ZN(
        U361) );
  INV_X1 U20572 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19620) );
  INV_X1 U20573 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20602) );
  AOI22_X1 U20574 ( .A1(n17389), .A2(n19620), .B1(n20602), .B2(n17390), .ZN(
        U362) );
  INV_X1 U20575 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19618) );
  INV_X1 U20576 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n21432) );
  AOI22_X1 U20577 ( .A1(n17389), .A2(n19618), .B1(n21432), .B2(n17390), .ZN(
        U363) );
  INV_X1 U20578 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19616) );
  INV_X1 U20579 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20600) );
  AOI22_X1 U20580 ( .A1(n17389), .A2(n19616), .B1(n20600), .B2(n17390), .ZN(
        U364) );
  INV_X1 U20581 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19578) );
  INV_X1 U20582 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20568) );
  AOI22_X1 U20583 ( .A1(n17389), .A2(n19578), .B1(n20568), .B2(n17390), .ZN(
        U365) );
  INV_X1 U20584 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19613) );
  INV_X1 U20585 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20598) );
  AOI22_X1 U20586 ( .A1(n17389), .A2(n19613), .B1(n20598), .B2(n17390), .ZN(
        U366) );
  INV_X1 U20587 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19612) );
  INV_X1 U20588 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20597) );
  AOI22_X1 U20589 ( .A1(n17389), .A2(n19612), .B1(n20597), .B2(n17390), .ZN(
        U367) );
  INV_X1 U20590 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19610) );
  INV_X1 U20591 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20595) );
  AOI22_X1 U20592 ( .A1(n17389), .A2(n19610), .B1(n20595), .B2(n17390), .ZN(
        U368) );
  INV_X1 U20593 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19608) );
  INV_X1 U20594 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n21415) );
  AOI22_X1 U20595 ( .A1(n17389), .A2(n19608), .B1(n21415), .B2(n17390), .ZN(
        U369) );
  INV_X1 U20596 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19606) );
  INV_X1 U20597 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20592) );
  AOI22_X1 U20598 ( .A1(n17389), .A2(n19606), .B1(n20592), .B2(n17390), .ZN(
        U370) );
  INV_X1 U20599 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19604) );
  INV_X1 U20600 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20590) );
  AOI22_X1 U20601 ( .A1(n17389), .A2(n19604), .B1(n20590), .B2(n17390), .ZN(
        U371) );
  INV_X1 U20602 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19601) );
  INV_X1 U20603 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20588) );
  AOI22_X1 U20604 ( .A1(n17389), .A2(n19601), .B1(n20588), .B2(n17390), .ZN(
        U372) );
  INV_X1 U20605 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19600) );
  INV_X1 U20606 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20586) );
  AOI22_X1 U20607 ( .A1(n17389), .A2(n19600), .B1(n20586), .B2(n17390), .ZN(
        U373) );
  INV_X1 U20608 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19598) );
  INV_X1 U20609 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20585) );
  AOI22_X1 U20610 ( .A1(n17389), .A2(n19598), .B1(n20585), .B2(n17390), .ZN(
        U374) );
  INV_X1 U20611 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19596) );
  INV_X1 U20612 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20584) );
  AOI22_X1 U20613 ( .A1(n17389), .A2(n19596), .B1(n20584), .B2(n17390), .ZN(
        U375) );
  INV_X1 U20614 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19576) );
  INV_X1 U20615 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20566) );
  AOI22_X1 U20616 ( .A1(n17389), .A2(n19576), .B1(n20566), .B2(n17390), .ZN(
        U376) );
  INV_X1 U20617 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n17392) );
  INV_X1 U20618 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19575) );
  NAND2_X1 U20619 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19575), .ZN(n19566) );
  INV_X1 U20620 ( .A(n19566), .ZN(n17391) );
  NOR2_X1 U20621 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n19561) );
  AOI21_X1 U20622 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(n17391), .A(n19561), 
        .ZN(n19558) );
  INV_X1 U20623 ( .A(n19558), .ZN(n19647) );
  OAI21_X1 U20624 ( .B1(n19572), .B2(n17392), .A(n19559), .ZN(P3_U2633) );
  INV_X1 U20625 ( .A(n19708), .ZN(n17395) );
  AND2_X1 U20626 ( .A1(n18305), .A2(n17400), .ZN(n17393) );
  OAI21_X1 U20627 ( .B1(n17393), .B2(n18304), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17394) );
  OAI21_X1 U20628 ( .B1(n17395), .B2(n19696), .A(n17394), .ZN(P3_U2634) );
  AOI22_X1 U20629 ( .A1(n19561), .A2(n19575), .B1(P3_D_C_N_REG_SCAN_IN), .B2(
        n19705), .ZN(n17396) );
  OAI21_X1 U20630 ( .B1(P3_CODEFETCH_REG_SCAN_IN), .B2(n19705), .A(n17396), 
        .ZN(P3_U2635) );
  OAI21_X1 U20631 ( .B1(n17397), .B2(BS16), .A(n19647), .ZN(n19645) );
  OAI21_X1 U20632 ( .B1(n19647), .B2(n17422), .A(n19645), .ZN(P3_U2636) );
  INV_X1 U20633 ( .A(n17398), .ZN(n17399) );
  AOI211_X1 U20634 ( .C1(n18305), .C2(n17400), .A(n17399), .B(n19523), .ZN(
        n19531) );
  NOR2_X1 U20635 ( .A1(n19531), .A2(n19547), .ZN(n19688) );
  OAI21_X1 U20636 ( .B1(n19688), .B2(n19047), .A(n17401), .ZN(P3_U2637) );
  NOR4_X1 U20637 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n17405) );
  NOR4_X1 U20638 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n17404) );
  NOR4_X1 U20639 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n17403) );
  NOR4_X1 U20640 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n17402) );
  NAND4_X1 U20641 ( .A1(n17405), .A2(n17404), .A3(n17403), .A4(n17402), .ZN(
        n17411) );
  NOR4_X1 U20642 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n17409) );
  AOI211_X1 U20643 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_15__SCAN_IN), .B(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17408) );
  NOR4_X1 U20644 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17407) );
  NOR4_X1 U20645 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n17406) );
  NAND4_X1 U20646 ( .A1(n17409), .A2(n17408), .A3(n17407), .A4(n17406), .ZN(
        n17410) );
  NOR2_X1 U20647 ( .A1(n17411), .A2(n17410), .ZN(n19682) );
  INV_X1 U20648 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19642) );
  NOR3_X1 U20649 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n17413) );
  OAI21_X1 U20650 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17413), .A(n19682), .ZN(
        n17412) );
  OAI21_X1 U20651 ( .B1(n19682), .B2(n19642), .A(n17412), .ZN(P3_U2638) );
  INV_X1 U20652 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19678) );
  INV_X1 U20653 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19646) );
  AOI21_X1 U20654 ( .B1(n19678), .B2(n19646), .A(n17413), .ZN(n17414) );
  INV_X1 U20655 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19639) );
  INV_X1 U20656 ( .A(n19682), .ZN(n19685) );
  AOI22_X1 U20657 ( .A1(n19682), .A2(n17414), .B1(n19639), .B2(n19685), .ZN(
        P3_U2639) );
  NAND2_X1 U20658 ( .A1(n17416), .A2(n17415), .ZN(n19522) );
  NAND3_X1 U20659 ( .A1(n19696), .A2(n19692), .A3(n17422), .ZN(n19557) );
  NOR2_X2 U20660 ( .A1(n19656), .A2(n19557), .ZN(n17753) );
  NOR2_X1 U20661 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19650), .ZN(n19388) );
  NAND2_X1 U20662 ( .A1(n19552), .A2(n19388), .ZN(n19545) );
  OAI211_X1 U20663 ( .C1(n19690), .C2(n19691), .A(n19702), .B(n17422), .ZN(
        n19540) );
  INV_X1 U20664 ( .A(n19540), .ZN(n17418) );
  AOI211_X4 U20665 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n19691), .A(n17418), .B(
        n17421), .ZN(n17800) );
  INV_X1 U20666 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19637) );
  INV_X1 U20667 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n21372) );
  INV_X1 U20668 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19623) );
  INV_X1 U20669 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19597) );
  INV_X1 U20670 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19584) );
  INV_X1 U20671 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19579) );
  NAND2_X1 U20672 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17781) );
  NOR2_X1 U20673 ( .A1(n19579), .A2(n17781), .ZN(n17747) );
  NAND2_X1 U20674 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17747), .ZN(n17730) );
  NOR2_X1 U20675 ( .A1(n19584), .A2(n17730), .ZN(n17650) );
  INV_X1 U20676 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19595) );
  INV_X1 U20677 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19593) );
  INV_X1 U20678 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19591) );
  NAND3_X1 U20679 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(P3_REIP_REG_6__SCAN_IN), .ZN(n17672) );
  NOR4_X1 U20680 ( .A1(n19595), .A2(n19593), .A3(n19591), .A4(n17672), .ZN(
        n17624) );
  NAND2_X1 U20681 ( .A1(n17650), .A2(n17624), .ZN(n17642) );
  NOR2_X1 U20682 ( .A1(n19597), .A2(n17642), .ZN(n17627) );
  NAND3_X1 U20683 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n17627), .ZN(n17528) );
  INV_X1 U20684 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19607) );
  NAND2_X1 U20685 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n17578) );
  NOR2_X1 U20686 ( .A1(n19607), .A2(n17578), .ZN(n17557) );
  NAND4_X1 U20687 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .A4(n17557), .ZN(n17536) );
  NAND2_X1 U20688 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n17537) );
  NOR3_X1 U20689 ( .A1(n17528), .A2(n17536), .A3(n17537), .ZN(n17518) );
  NAND2_X1 U20690 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n17518), .ZN(n17514) );
  NOR2_X1 U20691 ( .A1(n19623), .A2(n17514), .ZN(n17441) );
  NAND2_X1 U20692 ( .A1(n17782), .A2(n17441), .ZN(n17498) );
  INV_X1 U20693 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19624) );
  NAND4_X1 U20694 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n17476), .ZN(n17444) );
  NOR3_X1 U20695 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19637), .A3(n17444), 
        .ZN(n17419) );
  AOI21_X1 U20696 ( .B1(n17800), .B2(P3_EBX_REG_31__SCAN_IN), .A(n17419), .ZN(
        n17449) );
  NAND2_X1 U20697 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n19691), .ZN(n17420) );
  AOI211_X4 U20698 ( .C1(n17422), .C2(n19702), .A(n17421), .B(n17420), .ZN(
        n17799) );
  INV_X1 U20699 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17737) );
  NAND2_X1 U20700 ( .A1(n17745), .A2(n17737), .ZN(n17731) );
  INV_X1 U20701 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17711) );
  INV_X1 U20702 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17686) );
  INV_X1 U20703 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17663) );
  NAND2_X1 U20704 ( .A1(n17666), .A2(n17663), .ZN(n17660) );
  INV_X1 U20705 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n21373) );
  NAND2_X1 U20706 ( .A1(n17638), .A2(n21373), .ZN(n17634) );
  INV_X1 U20707 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17603) );
  INV_X1 U20708 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17953) );
  INV_X1 U20709 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17924) );
  NAND2_X1 U20710 ( .A1(n17568), .A2(n17924), .ZN(n17564) );
  INV_X1 U20711 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17901) );
  INV_X1 U20712 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17524) );
  INV_X1 U20713 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17502) );
  NAND2_X1 U20714 ( .A1(n17506), .A2(n17502), .ZN(n17501) );
  INV_X1 U20715 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17847) );
  NOR2_X1 U20716 ( .A1(n17791), .A2(n17450), .ZN(n17455) );
  INV_X1 U20717 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17814) );
  INV_X1 U20718 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17424) );
  NAND2_X1 U20719 ( .A1(n17439), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17425) );
  AOI21_X1 U20720 ( .B1(n17424), .B2(n17425), .A(n17423), .ZN(n18362) );
  OAI21_X1 U20721 ( .B1(n17439), .B2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n17425), .ZN(n18384) );
  INV_X1 U20722 ( .A(n18384), .ZN(n17479) );
  INV_X1 U20723 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17427) );
  NAND2_X1 U20724 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18433), .ZN(
        n18403) );
  INV_X1 U20725 ( .A(n18403), .ZN(n17430) );
  NAND2_X1 U20726 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17430), .ZN(
        n17428) );
  INV_X1 U20727 ( .A(n17428), .ZN(n17429) );
  NAND2_X1 U20728 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17429), .ZN(
        n17426) );
  NOR2_X1 U20729 ( .A1(n18413), .A2(n17428), .ZN(n18359) );
  AOI21_X1 U20730 ( .B1(n17427), .B2(n17426), .A(n18359), .ZN(n18404) );
  INV_X1 U20731 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18423) );
  AOI22_X1 U20732 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17429), .B1(
        n17428), .B2(n18423), .ZN(n18419) );
  INV_X1 U20733 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18435) );
  AOI21_X1 U20734 ( .B1(n18435), .B2(n18403), .A(n17429), .ZN(n18431) );
  INV_X1 U20735 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18449) );
  NOR2_X1 U20736 ( .A1(n18714), .A2(n18444), .ZN(n17433) );
  NAND2_X1 U20737 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17433), .ZN(
        n17431) );
  AOI21_X1 U20738 ( .B1(n18449), .B2(n17431), .A(n17430), .ZN(n18451) );
  XOR2_X1 U20739 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n17433), .Z(
        n18464) );
  NOR2_X1 U20740 ( .A1(n18714), .A2(n17432), .ZN(n17437) );
  INV_X1 U20741 ( .A(n17437), .ZN(n18442) );
  AOI21_X1 U20742 ( .B1(n18472), .B2(n18442), .A(n17433), .ZN(n18473) );
  NAND2_X1 U20743 ( .A1(n18562), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17435) );
  NAND2_X1 U20744 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17434), .ZN(
        n18564) );
  NOR2_X1 U20745 ( .A1(n17435), .A2(n18564), .ZN(n18521) );
  NAND2_X1 U20746 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18521), .ZN(
        n17600) );
  NOR2_X1 U20747 ( .A1(n18473), .A2(n17551), .ZN(n17550) );
  NOR2_X1 U20748 ( .A1(n17530), .A2(n17653), .ZN(n17517) );
  NOR2_X1 U20749 ( .A1(n18431), .A2(n17517), .ZN(n17516) );
  NOR2_X1 U20750 ( .A1(n17516), .A2(n17653), .ZN(n17508) );
  NOR2_X1 U20751 ( .A1(n18419), .A2(n17508), .ZN(n17507) );
  NOR2_X1 U20752 ( .A1(n17507), .A2(n17653), .ZN(n17497) );
  NOR2_X1 U20753 ( .A1(n18404), .A2(n17497), .ZN(n17496) );
  NOR2_X1 U20754 ( .A1(n17496), .A2(n17653), .ZN(n17489) );
  INV_X1 U20755 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17495) );
  INV_X1 U20756 ( .A(n18359), .ZN(n17440) );
  AOI21_X1 U20757 ( .B1(n17495), .B2(n17440), .A(n17439), .ZN(n18399) );
  NOR2_X1 U20758 ( .A1(n17488), .A2(n17653), .ZN(n17478) );
  NOR2_X1 U20759 ( .A1(n17479), .A2(n17478), .ZN(n17477) );
  NAND2_X1 U20760 ( .A1(n17436), .A2(n17753), .ZN(n17640) );
  NOR3_X1 U20761 ( .A1(n17452), .A2(n17451), .A3(n17640), .ZN(n17447) );
  NAND3_X1 U20762 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n17443) );
  NAND2_X1 U20763 ( .A1(n17788), .A2(n17801), .ZN(n17798) );
  NOR2_X1 U20764 ( .A1(n21372), .A2(n19624), .ZN(n17442) );
  OAI221_X1 U20765 ( .B1(n17788), .B2(n17442), .C1(n17788), .C2(n17441), .A(
        n17801), .ZN(n17492) );
  AOI21_X1 U20766 ( .B1(n17443), .B2(n17798), .A(n17492), .ZN(n17467) );
  NOR2_X1 U20767 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n17444), .ZN(n17454) );
  INV_X1 U20768 ( .A(n17454), .ZN(n17445) );
  AOI21_X1 U20769 ( .B1(n17467), .B2(n17445), .A(n19635), .ZN(n17446) );
  OAI211_X1 U20770 ( .C1(n13330), .C2(n17768), .A(n17449), .B(n17448), .ZN(
        P3_U2640) );
  NAND2_X1 U20771 ( .A1(n17799), .A2(n17450), .ZN(n17463) );
  OAI22_X1 U20772 ( .A1(n17467), .A2(n19637), .B1(n10347), .B2(n17768), .ZN(
        n17453) );
  INV_X1 U20773 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19632) );
  AOI211_X1 U20774 ( .C1(n17458), .C2(n17457), .A(n17456), .B(n19555), .ZN(
        n17462) );
  NAND3_X1 U20775 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n17476), .ZN(n17460) );
  OAI22_X1 U20776 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17460), .B1(n17459), 
        .B2(n17768), .ZN(n17461) );
  AOI211_X1 U20777 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n17800), .A(n17462), .B(
        n17461), .ZN(n17466) );
  INV_X1 U20778 ( .A(n17463), .ZN(n17464) );
  OAI21_X1 U20779 ( .B1(n17468), .B2(n17847), .A(n17464), .ZN(n17465) );
  OAI211_X1 U20780 ( .C1(n17467), .C2(n19632), .A(n17466), .B(n17465), .ZN(
        P3_U2642) );
  AOI22_X1 U20781 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17785), .B1(
        n17800), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n17475) );
  AOI211_X1 U20782 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17482), .A(n17468), .B(
        n17791), .ZN(n17471) );
  AOI211_X1 U20783 ( .C1(n18362), .C2(n17469), .A(n9713), .B(n19555), .ZN(
        n17470) );
  AOI211_X1 U20784 ( .C1(n17492), .C2(P3_REIP_REG_28__SCAN_IN), .A(n17471), 
        .B(n17470), .ZN(n17474) );
  NAND2_X1 U20785 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n17472) );
  OAI211_X1 U20786 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n17476), .B(n17472), .ZN(n17473) );
  NAND3_X1 U20787 ( .A1(n17475), .A2(n17474), .A3(n17473), .ZN(P3_U2643) );
  INV_X1 U20788 ( .A(n17476), .ZN(n17485) );
  AOI211_X1 U20789 ( .C1(n17479), .C2(n17478), .A(n17477), .B(n19555), .ZN(
        n17481) );
  INV_X1 U20790 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18387) );
  OAI22_X1 U20791 ( .A1(n18387), .A2(n17768), .B1(n17787), .B2(n17805), .ZN(
        n17480) );
  AOI211_X1 U20792 ( .C1(n17492), .C2(P3_REIP_REG_27__SCAN_IN), .A(n17481), 
        .B(n17480), .ZN(n17484) );
  OAI211_X1 U20793 ( .C1(n17487), .C2(n17805), .A(n17799), .B(n17482), .ZN(
        n17483) );
  OAI211_X1 U20794 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n17485), .A(n17484), 
        .B(n17483), .ZN(P3_U2644) );
  NOR3_X1 U20795 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n17498), .A3(n19624), 
        .ZN(n17486) );
  AOI21_X1 U20796 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17800), .A(n17486), .ZN(
        n17494) );
  AOI211_X1 U20797 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17501), .A(n17487), .B(
        n17791), .ZN(n17491) );
  AOI211_X1 U20798 ( .C1(n18399), .C2(n17489), .A(n17488), .B(n19555), .ZN(
        n17490) );
  AOI211_X1 U20799 ( .C1(n17492), .C2(P3_REIP_REG_26__SCAN_IN), .A(n17491), 
        .B(n17490), .ZN(n17493) );
  OAI211_X1 U20800 ( .C1(n17495), .C2(n17768), .A(n17494), .B(n17493), .ZN(
        P3_U2645) );
  NAND2_X1 U20801 ( .A1(n17782), .A2(n17514), .ZN(n17519) );
  NAND2_X1 U20802 ( .A1(n17801), .A2(n17519), .ZN(n17515) );
  AOI21_X1 U20803 ( .B1(n17782), .B2(n19623), .A(n17515), .ZN(n17505) );
  AOI211_X1 U20804 ( .C1(n18404), .C2(n17497), .A(n17496), .B(n19555), .ZN(
        n17500) );
  OAI22_X1 U20805 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n17498), .B1(n17787), 
        .B2(n17502), .ZN(n17499) );
  AOI211_X1 U20806 ( .C1(n17785), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n17500), .B(n17499), .ZN(n17504) );
  OAI211_X1 U20807 ( .C1(n17506), .C2(n17502), .A(n17799), .B(n17501), .ZN(
        n17503) );
  OAI211_X1 U20808 ( .C1(n17505), .C2(n19624), .A(n17504), .B(n17503), .ZN(
        P3_U2646) );
  NAND2_X1 U20809 ( .A1(n17782), .A2(n19623), .ZN(n17513) );
  AOI22_X1 U20810 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17785), .B1(
        n17800), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n17512) );
  AOI211_X1 U20811 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17523), .A(n17506), .B(
        n17791), .ZN(n17510) );
  AOI211_X1 U20812 ( .C1(n18419), .C2(n17508), .A(n17507), .B(n19555), .ZN(
        n17509) );
  AOI211_X1 U20813 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n17515), .A(n17510), 
        .B(n17509), .ZN(n17511) );
  OAI211_X1 U20814 ( .C1(n17514), .C2(n17513), .A(n17512), .B(n17511), .ZN(
        P3_U2647) );
  INV_X1 U20815 ( .A(n17515), .ZN(n17527) );
  INV_X1 U20816 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19619) );
  AOI211_X1 U20817 ( .C1(n18431), .C2(n17517), .A(n17516), .B(n19555), .ZN(
        n17522) );
  INV_X1 U20818 ( .A(n17518), .ZN(n17520) );
  OAI22_X1 U20819 ( .A1(n17787), .A2(n17524), .B1(n17520), .B2(n17519), .ZN(
        n17521) );
  AOI211_X1 U20820 ( .C1(n17785), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n17522), .B(n17521), .ZN(n17526) );
  OAI211_X1 U20821 ( .C1(n17532), .C2(n17524), .A(n17799), .B(n17523), .ZN(
        n17525) );
  OAI211_X1 U20822 ( .C1(n17527), .C2(n19619), .A(n17526), .B(n17525), .ZN(
        P3_U2648) );
  INV_X1 U20823 ( .A(n17801), .ZN(n17794) );
  AOI21_X1 U20824 ( .B1(n17528), .B2(n17782), .A(n17794), .ZN(n17623) );
  INV_X1 U20825 ( .A(n17623), .ZN(n17529) );
  AOI21_X1 U20826 ( .B1(n17782), .B2(n17536), .A(n17529), .ZN(n17540) );
  INV_X1 U20827 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19617) );
  AOI211_X1 U20828 ( .C1(n18451), .C2(n17531), .A(n17530), .B(n19555), .ZN(
        n17535) );
  AOI211_X1 U20829 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17544), .A(n17532), .B(
        n17791), .ZN(n17534) );
  INV_X1 U20830 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17864) );
  OAI22_X1 U20831 ( .A1(n18449), .A2(n17768), .B1(n17787), .B2(n17864), .ZN(
        n17533) );
  NOR3_X1 U20832 ( .A1(n17535), .A2(n17534), .A3(n17533), .ZN(n17539) );
  NAND4_X1 U20833 ( .A1(n17782), .A2(P3_REIP_REG_14__SCAN_IN), .A3(
        P3_REIP_REG_13__SCAN_IN), .A4(n17627), .ZN(n17590) );
  NOR2_X1 U20834 ( .A1(n17536), .A2(n17590), .ZN(n17543) );
  OAI211_X1 U20835 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(P3_REIP_REG_21__SCAN_IN), .A(n17543), .B(n17537), .ZN(n17538) );
  OAI211_X1 U20836 ( .C1(n17540), .C2(n19617), .A(n17539), .B(n17538), .ZN(
        P3_U2649) );
  AOI22_X1 U20837 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17785), .B1(
        n17800), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n17547) );
  INV_X1 U20838 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19615) );
  INV_X1 U20839 ( .A(n17540), .ZN(n17553) );
  AOI211_X1 U20840 ( .C1(n18464), .C2(n17541), .A(n9744), .B(n19555), .ZN(
        n17542) );
  AOI221_X1 U20841 ( .B1(n17543), .B2(n19615), .C1(n17553), .C2(
        P3_REIP_REG_21__SCAN_IN), .A(n17542), .ZN(n17546) );
  OAI211_X1 U20842 ( .C1(n17548), .C2(n17901), .A(n17799), .B(n17544), .ZN(
        n17545) );
  NAND3_X1 U20843 ( .A1(n17547), .A2(n17546), .A3(n17545), .ZN(P3_U2650) );
  AOI211_X1 U20844 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17564), .A(n17548), .B(
        n17791), .ZN(n17549) );
  AOI21_X1 U20845 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17800), .A(n17549), .ZN(
        n17556) );
  INV_X1 U20846 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19611) );
  INV_X1 U20847 ( .A(n17590), .ZN(n17607) );
  NAND3_X1 U20848 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n17557), .A3(n17607), 
        .ZN(n17562) );
  NOR2_X1 U20849 ( .A1(n19611), .A2(n17562), .ZN(n17554) );
  INV_X1 U20850 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19614) );
  AOI211_X1 U20851 ( .C1(n18473), .C2(n17551), .A(n17550), .B(n19555), .ZN(
        n17552) );
  AOI221_X1 U20852 ( .B1(n17554), .B2(n19614), .C1(n17553), .C2(
        P3_REIP_REG_20__SCAN_IN), .A(n17552), .ZN(n17555) );
  OAI211_X1 U20853 ( .C1(n18472), .C2(n17768), .A(n17556), .B(n17555), .ZN(
        P3_U2651) );
  AOI22_X1 U20854 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17785), .B1(
        n17800), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n17567) );
  INV_X1 U20855 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19609) );
  AND3_X1 U20856 ( .A1(n19609), .A2(n17557), .A3(n17607), .ZN(n17575) );
  OAI21_X1 U20857 ( .B1(n17557), .B2(n17788), .A(n17623), .ZN(n17582) );
  INV_X1 U20858 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17654) );
  NAND2_X1 U20859 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17654), .ZN(
        n17740) );
  NOR2_X1 U20860 ( .A1(n18485), .A2(n17740), .ZN(n17571) );
  AOI21_X1 U20861 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17571), .A(
        n17653), .ZN(n17560) );
  INV_X1 U20862 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18501) );
  INV_X1 U20863 ( .A(n18524), .ZN(n17558) );
  NAND2_X1 U20864 ( .A1(n17558), .A2(n18521), .ZN(n17591) );
  NOR2_X1 U20865 ( .A1(n10345), .A2(n17591), .ZN(n18484) );
  INV_X1 U20866 ( .A(n18484), .ZN(n17570) );
  NOR2_X1 U20867 ( .A1(n18501), .A2(n17570), .ZN(n17559) );
  OAI21_X1 U20868 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17559), .A(
        n18442), .ZN(n18488) );
  XOR2_X1 U20869 ( .A(n17560), .B(n18488), .Z(n17561) );
  OAI22_X1 U20870 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n17562), .B1(n19555), 
        .B2(n17561), .ZN(n17563) );
  AOI221_X1 U20871 ( .B1(n17575), .B2(P3_REIP_REG_19__SCAN_IN), .C1(n17582), 
        .C2(P3_REIP_REG_19__SCAN_IN), .A(n17563), .ZN(n17566) );
  OAI211_X1 U20872 ( .C1(n17568), .C2(n17924), .A(n17799), .B(n17564), .ZN(
        n17565) );
  NAND4_X1 U20873 ( .A1(n17567), .A2(n17566), .A3(n19024), .A4(n17565), .ZN(
        P3_U2652) );
  AOI211_X1 U20874 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17584), .A(n17568), .B(
        n17791), .ZN(n17569) );
  AOI211_X1 U20875 ( .C1(n17800), .C2(P3_EBX_REG_18__SCAN_IN), .A(n9586), .B(
        n17569), .ZN(n17577) );
  AOI22_X1 U20876 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17570), .B1(
        n18484), .B2(n18501), .ZN(n18498) );
  OR2_X1 U20877 ( .A1(n17571), .A2(n17653), .ZN(n17573) );
  OAI21_X1 U20878 ( .B1(n18498), .B2(n17573), .A(n17753), .ZN(n17572) );
  AOI21_X1 U20879 ( .B1(n18498), .B2(n17573), .A(n17572), .ZN(n17574) );
  AOI211_X1 U20880 ( .C1(P3_REIP_REG_18__SCAN_IN), .C2(n17582), .A(n17575), 
        .B(n17574), .ZN(n17576) );
  OAI211_X1 U20881 ( .C1(n18501), .C2(n17768), .A(n17577), .B(n17576), .ZN(
        P3_U2653) );
  AOI22_X1 U20882 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17785), .B1(
        n17800), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n17587) );
  NOR2_X1 U20883 ( .A1(n17578), .A2(n17590), .ZN(n17583) );
  AOI21_X1 U20884 ( .B1(n10345), .B2(n17591), .A(n18484), .ZN(n18512) );
  INV_X1 U20885 ( .A(n17740), .ZN(n17775) );
  AOI21_X1 U20886 ( .B1(n18508), .B2(n17775), .A(n17653), .ZN(n17580) );
  OAI21_X1 U20887 ( .B1(n18512), .B2(n17580), .A(n17753), .ZN(n17579) );
  AOI21_X1 U20888 ( .B1(n18512), .B2(n17580), .A(n17579), .ZN(n17581) );
  AOI221_X1 U20889 ( .B1(n17583), .B2(n19607), .C1(n17582), .C2(
        P3_REIP_REG_17__SCAN_IN), .A(n17581), .ZN(n17586) );
  OAI211_X1 U20890 ( .C1(n17588), .C2(n17953), .A(n17799), .B(n17584), .ZN(
        n17585) );
  NAND4_X1 U20891 ( .A1(n17587), .A2(n17586), .A3(n19024), .A4(n17585), .ZN(
        P3_U2654) );
  AOI211_X1 U20892 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17601), .A(n17588), .B(
        n17791), .ZN(n17589) );
  AOI211_X1 U20893 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n17785), .A(
        n9586), .B(n17589), .ZN(n17598) );
  OAI21_X1 U20894 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n17788), .A(n17623), 
        .ZN(n17606) );
  INV_X1 U20895 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19603) );
  NOR3_X1 U20896 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n19603), .A3(n17590), 
        .ZN(n17596) );
  INV_X1 U20897 ( .A(n17600), .ZN(n17592) );
  OAI21_X1 U20898 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17592), .A(
        n17591), .ZN(n18527) );
  INV_X1 U20899 ( .A(n17594), .ZN(n17608) );
  INV_X1 U20900 ( .A(n18527), .ZN(n17593) );
  AOI221_X1 U20901 ( .B1(n17594), .B2(n18527), .C1(n17608), .C2(n17593), .A(
        n19555), .ZN(n17595) );
  AOI211_X1 U20902 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(n17606), .A(n17596), 
        .B(n17595), .ZN(n17597) );
  OAI211_X1 U20903 ( .C1(n17787), .C2(n17599), .A(n17598), .B(n17597), .ZN(
        P3_U2655) );
  OAI21_X1 U20904 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18521), .A(
        n17600), .ZN(n18533) );
  OAI21_X1 U20905 ( .B1(n17653), .B2(n17654), .A(n17753), .ZN(n17797) );
  AOI211_X1 U20906 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17436), .A(
        n18533), .B(n17797), .ZN(n17605) );
  OAI211_X1 U20907 ( .C1(n17612), .C2(n17603), .A(n17799), .B(n17601), .ZN(
        n17602) );
  OAI211_X1 U20908 ( .C1(n17787), .C2(n17603), .A(n19024), .B(n17602), .ZN(
        n17604) );
  AOI211_X1 U20909 ( .C1(n17785), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n17605), .B(n17604), .ZN(n17611) );
  OAI21_X1 U20910 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n17607), .A(n17606), 
        .ZN(n17610) );
  NAND3_X1 U20911 ( .A1(n17753), .A2(n17608), .A3(n18533), .ZN(n17609) );
  NAND3_X1 U20912 ( .A1(n17611), .A2(n17610), .A3(n17609), .ZN(P3_U2656) );
  INV_X1 U20913 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19602) );
  NAND3_X1 U20914 ( .A1(n17782), .A2(P3_REIP_REG_13__SCAN_IN), .A3(n17627), 
        .ZN(n17622) );
  AOI211_X1 U20915 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17634), .A(n17612), .B(
        n17791), .ZN(n17620) );
  INV_X1 U20916 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17614) );
  INV_X1 U20917 ( .A(n18564), .ZN(n17613) );
  NAND2_X1 U20918 ( .A1(n18562), .A2(n17613), .ZN(n17626) );
  AOI21_X1 U20919 ( .B1(n17614), .B2(n17626), .A(n18521), .ZN(n18549) );
  OAI21_X1 U20920 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17626), .A(
        n17436), .ZN(n17628) );
  INV_X1 U20921 ( .A(n17628), .ZN(n17616) );
  INV_X1 U20922 ( .A(n18549), .ZN(n17615) );
  OAI221_X1 U20923 ( .B1(n18549), .B2(n17616), .C1(n17615), .C2(n17628), .A(
        n17753), .ZN(n17617) );
  OAI211_X1 U20924 ( .C1(n17787), .C2(n17618), .A(n19024), .B(n17617), .ZN(
        n17619) );
  AOI211_X1 U20925 ( .C1(n17785), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17620), .B(n17619), .ZN(n17621) );
  OAI221_X1 U20926 ( .B1(n17623), .B2(n19602), .C1(n17623), .C2(n17622), .A(
        n17621), .ZN(P3_U2657) );
  AOI22_X1 U20927 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17785), .B1(
        n17800), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n17637) );
  INV_X1 U20928 ( .A(n17624), .ZN(n17625) );
  NAND2_X1 U20929 ( .A1(n17650), .A2(n17801), .ZN(n17704) );
  OAI21_X1 U20930 ( .B1(n17625), .B2(n17704), .A(n17798), .ZN(n17657) );
  OAI21_X1 U20931 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n17788), .A(n17657), 
        .ZN(n17633) );
  NOR2_X1 U20932 ( .A1(n18581), .A2(n18564), .ZN(n17639) );
  OAI21_X1 U20933 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17639), .A(
        n17626), .ZN(n18565) );
  AOI211_X1 U20934 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17436), .A(
        n18565), .B(n17797), .ZN(n17632) );
  NAND2_X1 U20935 ( .A1(n17782), .A2(n17627), .ZN(n17630) );
  NAND2_X1 U20936 ( .A1(n17753), .A2(n18565), .ZN(n17629) );
  OAI22_X1 U20937 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17630), .B1(n17629), 
        .B2(n17628), .ZN(n17631) );
  AOI211_X1 U20938 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n17633), .A(n17632), 
        .B(n17631), .ZN(n17636) );
  OAI211_X1 U20939 ( .C1(n17638), .C2(n21373), .A(n17799), .B(n17634), .ZN(
        n17635) );
  NAND4_X1 U20940 ( .A1(n17637), .A2(n17636), .A3(n19024), .A4(n17635), .ZN(
        P3_U2658) );
  AOI211_X1 U20941 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17660), .A(n17638), .B(
        n17791), .ZN(n17647) );
  AOI21_X1 U20942 ( .B1(n18581), .B2(n18564), .A(n17639), .ZN(n18577) );
  INV_X1 U20943 ( .A(n17640), .ZN(n17786) );
  OAI21_X1 U20944 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18564), .A(
        n17786), .ZN(n17643) );
  NAND2_X1 U20945 ( .A1(n17782), .A2(n19597), .ZN(n17641) );
  OAI22_X1 U20946 ( .A1(n18577), .A2(n17643), .B1(n17642), .B2(n17641), .ZN(
        n17646) );
  OAI22_X1 U20947 ( .A1(n18581), .A2(n17768), .B1(n17787), .B2(n17644), .ZN(
        n17645) );
  NOR4_X1 U20948 ( .A1(n9586), .A2(n17647), .A3(n17646), .A4(n17645), .ZN(
        n17649) );
  INV_X1 U20949 ( .A(n17797), .ZN(n17718) );
  OAI211_X1 U20950 ( .C1(n18581), .C2(n17653), .A(n18577), .B(n17718), .ZN(
        n17648) );
  OAI211_X1 U20951 ( .C1(n17657), .C2(n19597), .A(n17649), .B(n17648), .ZN(
        P3_U2659) );
  NAND2_X1 U20952 ( .A1(n17782), .A2(n17650), .ZN(n17691) );
  NOR3_X1 U20953 ( .A1(n19591), .A2(n17672), .A3(n17691), .ZN(n17671) );
  AOI21_X1 U20954 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n17671), .A(
        P3_REIP_REG_11__SCAN_IN), .ZN(n17658) );
  INV_X1 U20955 ( .A(n18626), .ZN(n17651) );
  NAND2_X1 U20956 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17651), .ZN(
        n17701) );
  NOR2_X1 U20957 ( .A1(n17652), .A2(n17701), .ZN(n17665) );
  AOI21_X1 U20958 ( .B1(n17665), .B2(n17654), .A(n17653), .ZN(n17655) );
  OAI21_X1 U20959 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17665), .A(
        n18564), .ZN(n18589) );
  XOR2_X1 U20960 ( .A(n17655), .B(n18589), .Z(n17656) );
  OAI22_X1 U20961 ( .A1(n17658), .A2(n17657), .B1(n19555), .B2(n17656), .ZN(
        n17659) );
  AOI211_X1 U20962 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n17785), .A(
        n9586), .B(n17659), .ZN(n17662) );
  OAI211_X1 U20963 ( .C1(n17666), .C2(n17663), .A(n17799), .B(n17660), .ZN(
        n17661) );
  OAI211_X1 U20964 ( .C1(n17663), .C2(n17787), .A(n17662), .B(n17661), .ZN(
        P3_U2660) );
  INV_X1 U20965 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17668) );
  INV_X1 U20966 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18625) );
  NOR2_X1 U20967 ( .A1(n10338), .A2(n18625), .ZN(n18624) );
  INV_X1 U20968 ( .A(n18624), .ZN(n17664) );
  NAND2_X1 U20969 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18627), .ZN(
        n17715) );
  NOR2_X1 U20970 ( .A1(n17664), .A2(n17715), .ZN(n17693) );
  NAND2_X1 U20971 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17693), .ZN(
        n17678) );
  AOI21_X1 U20972 ( .B1(n17668), .B2(n17678), .A(n17665), .ZN(n18604) );
  OAI21_X1 U20973 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17678), .A(
        n17436), .ZN(n17681) );
  XOR2_X1 U20974 ( .A(n18604), .B(n17681), .Z(n17677) );
  AOI211_X1 U20975 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17685), .A(n17666), .B(
        n17791), .ZN(n17670) );
  OAI22_X1 U20976 ( .A1(n17668), .A2(n17768), .B1(n17787), .B2(n17667), .ZN(
        n17669) );
  NOR3_X1 U20977 ( .A1(n9586), .A2(n17670), .A3(n17669), .ZN(n17676) );
  INV_X1 U20978 ( .A(n17671), .ZN(n17674) );
  OAI21_X1 U20979 ( .B1(n17672), .B2(n17704), .A(n17798), .ZN(n17696) );
  INV_X1 U20980 ( .A(n17696), .ZN(n17684) );
  NOR3_X1 U20981 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n17672), .A3(n17691), .ZN(
        n17683) );
  NOR2_X1 U20982 ( .A1(n17684), .A2(n17683), .ZN(n17673) );
  MUX2_X1 U20983 ( .A(n17674), .B(n17673), .S(P3_REIP_REG_10__SCAN_IN), .Z(
        n17675) );
  OAI211_X1 U20984 ( .C1(n19555), .C2(n17677), .A(n17676), .B(n17675), .ZN(
        P3_U2661) );
  AOI22_X1 U20985 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17785), .B1(
        n17800), .B2(P3_EBX_REG_9__SCAN_IN), .ZN(n17689) );
  OAI21_X1 U20986 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17693), .A(
        n17678), .ZN(n18615) );
  NAND2_X1 U20987 ( .A1(n17753), .A2(n17653), .ZN(n17778) );
  INV_X1 U20988 ( .A(n18627), .ZN(n17703) );
  NOR2_X1 U20989 ( .A1(n17703), .A2(n17740), .ZN(n17679) );
  OAI221_X1 U20990 ( .B1(n18615), .B2(n18624), .C1(n18615), .C2(n17679), .A(
        n17753), .ZN(n17680) );
  AOI22_X1 U20991 ( .A1(n18615), .A2(n17681), .B1(n17778), .B2(n17680), .ZN(
        n17682) );
  AOI211_X1 U20992 ( .C1(n17684), .C2(P3_REIP_REG_9__SCAN_IN), .A(n17683), .B(
        n17682), .ZN(n17688) );
  OAI211_X1 U20993 ( .C1(n17690), .C2(n17686), .A(n17799), .B(n17685), .ZN(
        n17687) );
  NAND4_X1 U20994 ( .A1(n17689), .A2(n17688), .A3(n19024), .A4(n17687), .ZN(
        P3_U2662) );
  AOI211_X1 U20995 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17710), .A(n17690), .B(
        n17791), .ZN(n17699) );
  INV_X1 U20996 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19587) );
  INV_X1 U20997 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19585) );
  NOR2_X1 U20998 ( .A1(n19587), .A2(n19585), .ZN(n17692) );
  INV_X1 U20999 ( .A(n17691), .ZN(n17705) );
  AOI21_X1 U21000 ( .B1(n17692), .B2(n17705), .A(P3_REIP_REG_8__SCAN_IN), .ZN(
        n17697) );
  AOI21_X1 U21001 ( .B1(n18625), .B2(n17701), .A(n17693), .ZN(n18629) );
  OAI21_X1 U21002 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17701), .A(
        n17436), .ZN(n17694) );
  XOR2_X1 U21003 ( .A(n18629), .B(n17694), .Z(n17695) );
  OAI22_X1 U21004 ( .A1(n17697), .A2(n17696), .B1(n19555), .B2(n17695), .ZN(
        n17698) );
  AOI211_X1 U21005 ( .C1(n17785), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17699), .B(n17698), .ZN(n17700) );
  OAI211_X1 U21006 ( .C1(n17787), .C2(n18057), .A(n17700), .B(n19024), .ZN(
        P3_U2663) );
  INV_X1 U21007 ( .A(n17701), .ZN(n17702) );
  AOI21_X1 U21008 ( .B1(n10338), .B2(n17715), .A(n17702), .ZN(n18645) );
  OAI21_X1 U21009 ( .B1(n17703), .B2(n17740), .A(n17436), .ZN(n17726) );
  XNOR2_X1 U21010 ( .A(n18645), .B(n17726), .ZN(n17709) );
  NAND2_X1 U21011 ( .A1(n17798), .A2(n17704), .ZN(n17729) );
  NAND2_X1 U21012 ( .A1(n17705), .A2(n19585), .ZN(n17723) );
  AOI21_X1 U21013 ( .B1(n17729), .B2(n17723), .A(n19587), .ZN(n17708) );
  NAND3_X1 U21014 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n17705), .A3(n19587), 
        .ZN(n17706) );
  OAI211_X1 U21015 ( .C1(n17787), .C2(n17711), .A(n19024), .B(n17706), .ZN(
        n17707) );
  AOI211_X1 U21016 ( .C1(n17709), .C2(n17753), .A(n17708), .B(n17707), .ZN(
        n17713) );
  OAI211_X1 U21017 ( .C1(n17716), .C2(n17711), .A(n17799), .B(n17710), .ZN(
        n17712) );
  OAI211_X1 U21018 ( .C1(n17768), .C2(n10338), .A(n17713), .B(n17712), .ZN(
        P3_U2664) );
  NOR2_X1 U21019 ( .A1(n18714), .A2(n17714), .ZN(n17728) );
  OAI21_X1 U21020 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17728), .A(
        n17715), .ZN(n18657) );
  NAND2_X1 U21021 ( .A1(n17753), .A2(n18657), .ZN(n17725) );
  AOI211_X1 U21022 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17731), .A(n17716), .B(
        n17791), .ZN(n17722) );
  INV_X1 U21023 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17717) );
  OAI22_X1 U21024 ( .A1(n18652), .A2(n17768), .B1(n17787), .B2(n17717), .ZN(
        n17721) );
  OAI21_X1 U21025 ( .B1(n18652), .B2(n17653), .A(n17718), .ZN(n17719) );
  OAI22_X1 U21026 ( .A1(n19585), .A2(n17729), .B1(n18657), .B2(n17719), .ZN(
        n17720) );
  NOR4_X1 U21027 ( .A1(n9586), .A2(n17722), .A3(n17721), .A4(n17720), .ZN(
        n17724) );
  OAI211_X1 U21028 ( .C1(n17726), .C2(n17725), .A(n17724), .B(n17723), .ZN(
        P3_U2665) );
  NAND2_X1 U21029 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17727), .ZN(
        n17739) );
  AOI21_X1 U21030 ( .B1(n10337), .B2(n17739), .A(n17728), .ZN(n18669) );
  OAI21_X1 U21031 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17739), .A(
        n17436), .ZN(n17741) );
  XNOR2_X1 U21032 ( .A(n18669), .B(n17741), .ZN(n17735) );
  AOI221_X1 U21033 ( .B1(n17788), .B2(n19584), .C1(n17730), .C2(n19584), .A(
        n17729), .ZN(n17734) );
  OAI211_X1 U21034 ( .C1(n17745), .C2(n17737), .A(n17799), .B(n17731), .ZN(
        n17732) );
  OAI21_X1 U21035 ( .B1(n17768), .B2(n10337), .A(n17732), .ZN(n17733) );
  AOI211_X1 U21036 ( .C1(n17753), .C2(n17735), .A(n17734), .B(n17733), .ZN(
        n17736) );
  OAI211_X1 U21037 ( .C1(n17787), .C2(n17737), .A(n17736), .B(n19024), .ZN(
        P3_U2666) );
  NOR2_X1 U21038 ( .A1(n17747), .A2(n17788), .ZN(n17756) );
  NOR2_X1 U21039 ( .A1(n17794), .A2(n17756), .ZN(n17761) );
  INV_X1 U21040 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19581) );
  NOR2_X1 U21041 ( .A1(n18714), .A2(n17738), .ZN(n17758) );
  OAI21_X1 U21042 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17758), .A(
        n17739), .ZN(n18682) );
  INV_X1 U21043 ( .A(n18682), .ZN(n17742) );
  OR2_X1 U21044 ( .A1(n17738), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18678) );
  OAI22_X1 U21045 ( .A1(n17742), .A2(n17741), .B1(n17740), .B2(n18678), .ZN(
        n17752) );
  NOR2_X1 U21046 ( .A1(n17743), .A2(n19698), .ZN(n19712) );
  OAI21_X1 U21047 ( .B1(n18065), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n19712), .ZN(n17744) );
  OAI211_X1 U21048 ( .C1(n18682), .C2(n17778), .A(n19024), .B(n17744), .ZN(
        n17751) );
  AOI211_X1 U21049 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17764), .A(n17745), .B(
        n17791), .ZN(n17746) );
  AOI21_X1 U21050 ( .B1(n17785), .B2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n17746), .ZN(n17749) );
  NAND3_X1 U21051 ( .A1(n17782), .A2(n17747), .A3(n19581), .ZN(n17748) );
  OAI211_X1 U21052 ( .C1(n18088), .C2(n17787), .A(n17749), .B(n17748), .ZN(
        n17750) );
  AOI211_X1 U21053 ( .C1(n17753), .C2(n17752), .A(n17751), .B(n17750), .ZN(
        n17754) );
  OAI21_X1 U21054 ( .B1(n17761), .B2(n19581), .A(n17754), .ZN(P3_U2667) );
  INV_X1 U21055 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18699) );
  NOR2_X1 U21056 ( .A1(n19663), .A2(n13161), .ZN(n19495) );
  NAND2_X1 U21057 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19495), .ZN(
        n17771) );
  AOI21_X1 U21058 ( .B1(n17771), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13081), .ZN(n17755) );
  INV_X1 U21059 ( .A(n17755), .ZN(n19651) );
  INV_X1 U21060 ( .A(n17756), .ZN(n17757) );
  OAI22_X1 U21061 ( .A1(n17787), .A2(n17765), .B1(n17781), .B2(n17757), .ZN(
        n17763) );
  NAND2_X1 U21062 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17773) );
  AOI21_X1 U21063 ( .B1(n18699), .B2(n17773), .A(n17758), .ZN(n18697) );
  OAI21_X1 U21064 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17773), .A(
        n17436), .ZN(n17759) );
  XOR2_X1 U21065 ( .A(n18697), .B(n17759), .Z(n17760) );
  OAI22_X1 U21066 ( .A1(n17761), .A2(n19579), .B1(n19555), .B2(n17760), .ZN(
        n17762) );
  AOI211_X1 U21067 ( .C1(n19712), .C2(n19651), .A(n17763), .B(n17762), .ZN(
        n17767) );
  OAI211_X1 U21068 ( .C1(n17769), .C2(n17765), .A(n17799), .B(n17764), .ZN(
        n17766) );
  OAI211_X1 U21069 ( .C1(n17768), .C2(n18699), .A(n17767), .B(n17766), .ZN(
        P3_U2668) );
  OR2_X1 U21070 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), .ZN(
        n17770) );
  AOI211_X1 U21071 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17770), .A(n17769), .B(
        n17791), .ZN(n17780) );
  OAI21_X1 U21072 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17773), .ZN(n18706) );
  NAND2_X1 U21073 ( .A1(n19663), .A2(n19508), .ZN(n19497) );
  NAND2_X1 U21074 ( .A1(n19497), .A2(n17771), .ZN(n19657) );
  INV_X1 U21075 ( .A(n19657), .ZN(n17772) );
  AOI22_X1 U21076 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n17794), .B1(n17772), 
        .B2(n19712), .ZN(n17777) );
  OR2_X1 U21077 ( .A1(n17773), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17774) );
  OAI211_X1 U21078 ( .C1(n17775), .C2(n18706), .A(n17786), .B(n17774), .ZN(
        n17776) );
  OAI211_X1 U21079 ( .C1(n17778), .C2(n18706), .A(n17777), .B(n17776), .ZN(
        n17779) );
  AOI211_X1 U21080 ( .C1(n17785), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n17780), .B(n17779), .ZN(n17784) );
  OAI211_X1 U21081 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17782), .B(n17781), .ZN(n17783) );
  OAI211_X1 U21082 ( .C1(n9972), .C2(n17787), .A(n17784), .B(n17783), .ZN(
        P3_U2669) );
  AOI21_X1 U21083 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17786), .A(
        n17785), .ZN(n17796) );
  OAI22_X1 U21084 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17788), .B1(n17787), 
        .B2(n9973), .ZN(n17793) );
  NAND2_X1 U21085 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n18096) );
  OAI21_X1 U21086 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n18096), .ZN(n18104) );
  NAND2_X1 U21087 ( .A1(n17789), .A2(n19508), .ZN(n19664) );
  INV_X1 U21088 ( .A(n19712), .ZN(n17790) );
  OAI22_X1 U21089 ( .A1(n17791), .A2(n18104), .B1(n19664), .B2(n17790), .ZN(
        n17792) );
  AOI211_X1 U21090 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(n17794), .A(n17793), .B(
        n17792), .ZN(n17795) );
  OAI221_X1 U21091 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17797), .C1(
        n18714), .C2(n17796), .A(n17795), .ZN(P3_U2670) );
  AOI22_X1 U21092 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n17798), .B1(n19712), 
        .B2(n13162), .ZN(n17804) );
  OAI21_X1 U21093 ( .B1(n17800), .B2(n17799), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n17803) );
  NAND3_X1 U21094 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19659), .A3(
        n17801), .ZN(n17802) );
  NAND3_X1 U21095 ( .A1(n17804), .A2(n17803), .A3(n17802), .ZN(P3_U2671) );
  NOR2_X1 U21096 ( .A1(n17806), .A2(n17805), .ZN(n17810) );
  INV_X1 U21097 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17808) );
  NOR4_X1 U21098 ( .A1(n17847), .A2(n17808), .A3(n17887), .A4(n17807), .ZN(
        n17809) );
  NAND4_X1 U21099 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n17810), .A4(n17809), .ZN(n17813) );
  NAND2_X1 U21100 ( .A1(n18101), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17812) );
  NAND2_X1 U21101 ( .A1(n17843), .A2(n19084), .ZN(n17811) );
  OAI22_X1 U21102 ( .A1(n17843), .A2(n17812), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17811), .ZN(P3_U2672) );
  NAND2_X1 U21103 ( .A1(n17814), .A2(n17813), .ZN(n17815) );
  NAND2_X1 U21104 ( .A1(n17815), .A2(n18101), .ZN(n17842) );
  AOI22_X1 U21105 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18038), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17827) );
  AOI22_X1 U21106 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17830), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17826) );
  AOI22_X1 U21107 ( .A1(n18058), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17817) );
  OAI21_X1 U21108 ( .B1(n13197), .B2(n18078), .A(n17817), .ZN(n17823) );
  AOI22_X1 U21109 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17821) );
  AOI22_X1 U21110 ( .A1(n18063), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18064), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17820) );
  AOI22_X1 U21111 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17819) );
  AOI22_X1 U21112 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9587), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17818) );
  NAND4_X1 U21113 ( .A1(n17821), .A2(n17820), .A3(n17819), .A4(n17818), .ZN(
        n17822) );
  AOI211_X1 U21114 ( .C1(n17824), .C2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n17823), .B(n17822), .ZN(n17825) );
  NAND3_X1 U21115 ( .A1(n17827), .A2(n17826), .A3(n17825), .ZN(n17841) );
  AOI22_X1 U21116 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17839) );
  AOI22_X1 U21117 ( .A1(n18044), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17838) );
  AOI22_X1 U21118 ( .A1(n9587), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n9594), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17828) );
  OAI21_X1 U21119 ( .B1(n13197), .B2(n17829), .A(n17828), .ZN(n17836) );
  AOI22_X1 U21120 ( .A1(n13081), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17830), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17834) );
  AOI22_X1 U21121 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18062), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17833) );
  AOI22_X1 U21122 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17832) );
  AOI22_X1 U21123 ( .A1(n18018), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17945), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17831) );
  NAND4_X1 U21124 ( .A1(n17834), .A2(n17833), .A3(n17832), .A4(n17831), .ZN(
        n17835) );
  AOI211_X1 U21125 ( .C1(n9590), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n17836), .B(n17835), .ZN(n17837) );
  AND3_X1 U21126 ( .A1(n17839), .A2(n17838), .A3(n17837), .ZN(n17845) );
  NOR3_X1 U21127 ( .A1(n17845), .A2(n17844), .A3(n17851), .ZN(n17840) );
  XNOR2_X1 U21128 ( .A(n17841), .B(n17840), .ZN(n18114) );
  OAI22_X1 U21129 ( .A1(n17843), .A2(n17842), .B1(n18114), .B2(n18101), .ZN(
        P3_U2673) );
  NOR2_X1 U21130 ( .A1(n17851), .A2(n17844), .ZN(n17846) );
  XOR2_X1 U21131 ( .A(n17846), .B(n17845), .Z(n18121) );
  AOI22_X1 U21132 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17849), .B1(n17848), 
        .B2(n17847), .ZN(n17850) );
  OAI21_X1 U21133 ( .B1(n18101), .B2(n18121), .A(n17850), .ZN(P3_U2674) );
  OAI21_X1 U21134 ( .B1(n17853), .B2(n17852), .A(n17851), .ZN(n18131) );
  NAND3_X1 U21135 ( .A1(n17855), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n18101), 
        .ZN(n17854) );
  OAI221_X1 U21136 ( .B1(n17855), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n18101), 
        .C2(n18131), .A(n17854), .ZN(P3_U2676) );
  AOI21_X1 U21137 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18101), .A(n17863), .ZN(
        n17857) );
  XNOR2_X1 U21138 ( .A(n17856), .B(n17859), .ZN(n18135) );
  OAI22_X1 U21139 ( .A1(n17858), .A2(n17857), .B1(n18101), .B2(n18135), .ZN(
        P3_U2677) );
  AOI21_X1 U21140 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18101), .A(n17867), .ZN(
        n17862) );
  OAI21_X1 U21141 ( .B1(n17861), .B2(n17860), .A(n17859), .ZN(n18139) );
  OAI22_X1 U21142 ( .A1(n17863), .A2(n17862), .B1(n18101), .B2(n18139), .ZN(
        P3_U2678) );
  AOI21_X1 U21143 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18101), .A(n17872), .ZN(
        n17866) );
  XNOR2_X1 U21144 ( .A(n17865), .B(n17868), .ZN(n18145) );
  OAI22_X1 U21145 ( .A1(n17867), .A2(n17866), .B1(n18101), .B2(n18145), .ZN(
        P3_U2679) );
  AOI21_X1 U21146 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18101), .A(n17886), .ZN(
        n17871) );
  OAI21_X1 U21147 ( .B1(n17870), .B2(n17869), .A(n17868), .ZN(n18149) );
  OAI22_X1 U21148 ( .A1(n17872), .A2(n17871), .B1(n18101), .B2(n18149), .ZN(
        P3_U2680) );
  INV_X1 U21149 ( .A(n17873), .ZN(n17874) );
  AOI21_X1 U21150 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18101), .A(n17874), .ZN(
        n17885) );
  AOI22_X1 U21151 ( .A1(n13081), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17878) );
  AOI22_X1 U21152 ( .A1(n13202), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18062), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17877) );
  AOI22_X1 U21153 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17876) );
  AOI22_X1 U21154 ( .A1(n18018), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13253), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17875) );
  NAND4_X1 U21155 ( .A1(n17878), .A2(n17877), .A3(n17876), .A4(n17875), .ZN(
        n17884) );
  AOI22_X1 U21156 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17882) );
  AOI22_X1 U21157 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18065), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17881) );
  AOI22_X1 U21158 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17880) );
  AOI22_X1 U21159 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17879) );
  NAND4_X1 U21160 ( .A1(n17882), .A2(n17881), .A3(n17880), .A4(n17879), .ZN(
        n17883) );
  NOR2_X1 U21161 ( .A1(n17884), .A2(n17883), .ZN(n18151) );
  OAI22_X1 U21162 ( .A1(n17886), .A2(n17885), .B1(n18151), .B2(n18101), .ZN(
        P3_U2681) );
  NAND2_X1 U21163 ( .A1(n18101), .A2(n17887), .ZN(n17912) );
  AOI22_X1 U21164 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18065), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17898) );
  AOI22_X1 U21165 ( .A1(n18038), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17897) );
  AOI22_X1 U21166 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17888) );
  OAI21_X1 U21167 ( .B1(n9584), .B2(n18086), .A(n17888), .ZN(n17895) );
  AOI22_X1 U21168 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17893) );
  AOI22_X1 U21169 ( .A1(n17945), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17892) );
  AOI22_X1 U21170 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17891) );
  AOI22_X1 U21171 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13253), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17890) );
  NAND4_X1 U21172 ( .A1(n17893), .A2(n17892), .A3(n17891), .A4(n17890), .ZN(
        n17894) );
  AOI211_X1 U21173 ( .C1(n18018), .C2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n17895), .B(n17894), .ZN(n17896) );
  NAND3_X1 U21174 ( .A1(n17898), .A2(n17897), .A3(n17896), .ZN(n18157) );
  AOI22_X1 U21175 ( .A1(n18106), .A2(n18157), .B1(n17899), .B2(n17901), .ZN(
        n17900) );
  OAI21_X1 U21176 ( .B1(n17901), .B2(n17912), .A(n17900), .ZN(P3_U2682) );
  NOR3_X1 U21177 ( .A1(n18213), .A2(n21333), .A3(n17937), .ZN(n17925) );
  AOI21_X1 U21178 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17925), .A(
        P3_EBX_REG_20__SCAN_IN), .ZN(n17913) );
  AOI22_X1 U21179 ( .A1(n13076), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18065), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17905) );
  AOI22_X1 U21180 ( .A1(n17946), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17945), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17904) );
  AOI22_X1 U21181 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17903) );
  AOI22_X1 U21182 ( .A1(n13253), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17902) );
  NAND4_X1 U21183 ( .A1(n17905), .A2(n17904), .A3(n17903), .A4(n17902), .ZN(
        n17911) );
  AOI22_X1 U21184 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17961), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17909) );
  AOI22_X1 U21185 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17908) );
  AOI22_X1 U21186 ( .A1(n18044), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18001), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17907) );
  AOI22_X1 U21187 ( .A1(n18038), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17906) );
  NAND4_X1 U21188 ( .A1(n17909), .A2(n17908), .A3(n17907), .A4(n17906), .ZN(
        n17910) );
  NOR2_X1 U21189 ( .A1(n17911), .A2(n17910), .ZN(n18166) );
  OAI22_X1 U21190 ( .A1(n17913), .A2(n17912), .B1(n18166), .B2(n18101), .ZN(
        P3_U2683) );
  AOI22_X1 U21191 ( .A1(n17946), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17917) );
  AOI22_X1 U21192 ( .A1(n17960), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17916) );
  AOI22_X1 U21193 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17915) );
  AOI22_X1 U21194 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13253), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17914) );
  NAND4_X1 U21195 ( .A1(n17917), .A2(n17916), .A3(n17915), .A4(n17914), .ZN(
        n17923) );
  AOI22_X1 U21196 ( .A1(n18065), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18001), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17921) );
  AOI22_X1 U21197 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17920) );
  AOI22_X1 U21198 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17945), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17919) );
  AOI22_X1 U21199 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18062), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17918) );
  NAND4_X1 U21200 ( .A1(n17921), .A2(n17920), .A3(n17919), .A4(n17918), .ZN(
        n17922) );
  NOR2_X1 U21201 ( .A1(n17923), .A2(n17922), .ZN(n18170) );
  NOR2_X1 U21202 ( .A1(n18106), .A2(n9727), .ZN(n17938) );
  AOI22_X1 U21203 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17938), .B1(n17925), 
        .B2(n17924), .ZN(n17926) );
  OAI21_X1 U21204 ( .B1(n18170), .B2(n18101), .A(n17926), .ZN(P3_U2684) );
  AOI22_X1 U21205 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17930) );
  AOI22_X1 U21206 ( .A1(n13081), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18062), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17929) );
  AOI22_X1 U21207 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18065), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17928) );
  AOI22_X1 U21208 ( .A1(n13253), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17927) );
  NAND4_X1 U21209 ( .A1(n17930), .A2(n17929), .A3(n17928), .A4(n17927), .ZN(
        n17936) );
  AOI22_X1 U21210 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17934) );
  AOI22_X1 U21211 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18059), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17933) );
  AOI22_X1 U21212 ( .A1(n17946), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17932) );
  AOI22_X1 U21213 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17931) );
  NAND4_X1 U21214 ( .A1(n17934), .A2(n17933), .A3(n17932), .A4(n17931), .ZN(
        n17935) );
  NOR2_X1 U21215 ( .A1(n17936), .A2(n17935), .ZN(n18175) );
  INV_X1 U21216 ( .A(n17937), .ZN(n17939) );
  OAI21_X1 U21217 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17939), .A(n17938), .ZN(
        n17940) );
  OAI21_X1 U21218 ( .B1(n18175), .B2(n18101), .A(n17940), .ZN(P3_U2685) );
  AOI22_X1 U21219 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18046), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n18065), .ZN(n17944) );
  AOI22_X1 U21220 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n18058), .ZN(n17943) );
  AOI22_X1 U21221 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n9588), .ZN(n17942) );
  AOI22_X1 U21222 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n13253), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17941) );
  NAND4_X1 U21223 ( .A1(n17944), .A2(n17943), .A3(n17942), .A4(n17941), .ZN(
        n17952) );
  AOI22_X1 U21224 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n9594), .ZN(n17950) );
  AOI22_X1 U21225 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17945), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17949) );
  AOI22_X1 U21226 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17946), .B1(
        n17960), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17948) );
  AOI22_X1 U21227 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18044), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n18045), .ZN(n17947) );
  NAND4_X1 U21228 ( .A1(n17950), .A2(n17949), .A3(n17948), .A4(n17947), .ZN(
        n17951) );
  NOR2_X1 U21229 ( .A1(n17952), .A2(n17951), .ZN(n18181) );
  NOR2_X1 U21230 ( .A1(n18106), .A2(n17954), .ZN(n17968) );
  OAI222_X1 U21231 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n19084), .B1(
        P3_EBX_REG_17__SCAN_IN), .B2(n17954), .C1(n17968), .C2(n17953), .ZN(
        n17955) );
  OAI21_X1 U21232 ( .B1(n18181), .B2(n18101), .A(n17955), .ZN(P3_U2686) );
  AOI22_X1 U21233 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17959) );
  AOI22_X1 U21234 ( .A1(n13076), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17958) );
  AOI22_X1 U21235 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17957) );
  AOI22_X1 U21236 ( .A1(n13253), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18001), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17956) );
  NAND4_X1 U21237 ( .A1(n17959), .A2(n17958), .A3(n17957), .A4(n17956), .ZN(
        n17967) );
  AOI22_X1 U21238 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17960), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17965) );
  AOI22_X1 U21239 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17964) );
  AOI22_X1 U21240 ( .A1(n17946), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17961), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17963) );
  AOI22_X1 U21241 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18065), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17962) );
  NAND4_X1 U21242 ( .A1(n17965), .A2(n17964), .A3(n17963), .A4(n17962), .ZN(
        n17966) );
  NOR2_X1 U21243 ( .A1(n17967), .A2(n17966), .ZN(n18187) );
  INV_X1 U21244 ( .A(n17981), .ZN(n17969) );
  OAI21_X1 U21245 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17969), .A(n17968), .ZN(
        n17970) );
  OAI21_X1 U21246 ( .B1(n18187), .B2(n18101), .A(n17970), .ZN(P3_U2687) );
  AOI22_X1 U21247 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17974) );
  AOI22_X1 U21248 ( .A1(n18018), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17973) );
  AOI22_X1 U21249 ( .A1(n18058), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17972) );
  AOI22_X1 U21250 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13253), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17971) );
  NAND4_X1 U21251 ( .A1(n17974), .A2(n17973), .A3(n17972), .A4(n17971), .ZN(
        n17980) );
  AOI22_X1 U21252 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18065), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17978) );
  AOI22_X1 U21253 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18059), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17977) );
  AOI22_X1 U21254 ( .A1(n18038), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17976) );
  AOI22_X1 U21255 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18062), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17975) );
  NAND4_X1 U21256 ( .A1(n17978), .A2(n17977), .A3(n17976), .A4(n17975), .ZN(
        n17979) );
  NOR2_X1 U21257 ( .A1(n17980), .A2(n17979), .ZN(n18192) );
  OAI21_X1 U21258 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17996), .A(n17981), .ZN(
        n17982) );
  AOI22_X1 U21259 ( .A1(n18106), .A2(n18192), .B1(n17982), .B2(n18101), .ZN(
        P3_U2688) );
  INV_X1 U21260 ( .A(n17983), .ZN(n17984) );
  OAI21_X1 U21261 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17984), .A(n18101), .ZN(
        n17995) );
  AOI22_X1 U21262 ( .A1(n17946), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18065), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17988) );
  AOI22_X1 U21263 ( .A1(n18044), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17987) );
  AOI22_X1 U21264 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18026), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17986) );
  AOI22_X1 U21265 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13253), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17985) );
  NAND4_X1 U21266 ( .A1(n17988), .A2(n17987), .A3(n17986), .A4(n17985), .ZN(
        n17994) );
  AOI22_X1 U21267 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17992) );
  AOI22_X1 U21268 ( .A1(n17041), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18059), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17991) );
  AOI22_X1 U21269 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17990) );
  AOI22_X1 U21270 ( .A1(n18038), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18046), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17989) );
  NAND4_X1 U21271 ( .A1(n17992), .A2(n17991), .A3(n17990), .A4(n17989), .ZN(
        n17993) );
  NOR2_X1 U21272 ( .A1(n17994), .A2(n17993), .ZN(n18198) );
  OAI22_X1 U21273 ( .A1(n17996), .A2(n17995), .B1(n18198), .B2(n18101), .ZN(
        P3_U2689) );
  OR2_X1 U21274 ( .A1(n18213), .A2(n18022), .ZN(n18009) );
  AOI22_X1 U21275 ( .A1(n18038), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18000) );
  AOI22_X1 U21276 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17999) );
  AOI22_X1 U21277 ( .A1(n18018), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18010), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17998) );
  AOI22_X1 U21278 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13253), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17997) );
  NAND4_X1 U21279 ( .A1(n18000), .A2(n17999), .A3(n17998), .A4(n17997), .ZN(
        n18007) );
  AOI22_X1 U21280 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18065), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18005) );
  AOI22_X1 U21281 ( .A1(n18044), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18001), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18004) );
  AOI22_X1 U21282 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18003) );
  AOI22_X1 U21283 ( .A1(n13202), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n18002) );
  NAND4_X1 U21284 ( .A1(n18005), .A2(n18004), .A3(n18003), .A4(n18002), .ZN(
        n18006) );
  NOR2_X1 U21285 ( .A1(n18007), .A2(n18006), .ZN(n18204) );
  NAND3_X1 U21286 ( .A1(n18009), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n18101), 
        .ZN(n18008) );
  OAI221_X1 U21287 ( .B1(n18009), .B2(P3_EBX_REG_12__SCAN_IN), .C1(n18101), 
        .C2(n18204), .A(n18008), .ZN(P3_U2691) );
  AOI22_X1 U21288 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18021) );
  AOI22_X1 U21289 ( .A1(n18043), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18065), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18020) );
  INV_X1 U21290 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18095) );
  AOI22_X1 U21291 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18045), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18011) );
  OAI21_X1 U21292 ( .B1(n9592), .B2(n18095), .A(n18011), .ZN(n18017) );
  AOI22_X1 U21293 ( .A1(n13202), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18015) );
  AOI22_X1 U21294 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18014) );
  AOI22_X1 U21295 ( .A1(n18038), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18013) );
  AOI22_X1 U21296 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18012) );
  NAND4_X1 U21297 ( .A1(n18015), .A2(n18014), .A3(n18013), .A4(n18012), .ZN(
        n18016) );
  AOI211_X1 U21298 ( .C1(n18018), .C2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n18017), .B(n18016), .ZN(n18019) );
  NAND3_X1 U21299 ( .A1(n18021), .A2(n18020), .A3(n18019), .ZN(n18207) );
  INV_X1 U21300 ( .A(n18207), .ZN(n18024) );
  OAI21_X1 U21301 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n9746), .A(n18022), .ZN(
        n18023) );
  AOI22_X1 U21302 ( .A1(n18106), .A2(n18024), .B1(n18023), .B2(n18101), .ZN(
        P3_U2692) );
  INV_X1 U21303 ( .A(n18053), .ZN(n18025) );
  OAI21_X1 U21304 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n18025), .A(n18101), .ZN(
        n18037) );
  AOI22_X1 U21305 ( .A1(n9590), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18010), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18030) );
  AOI22_X1 U21306 ( .A1(n18026), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18029) );
  AOI22_X1 U21307 ( .A1(n13081), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18028) );
  AOI22_X1 U21308 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13253), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18027) );
  NAND4_X1 U21309 ( .A1(n18030), .A2(n18029), .A3(n18028), .A4(n18027), .ZN(
        n18036) );
  AOI22_X1 U21310 ( .A1(n13202), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18034) );
  AOI22_X1 U21311 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18065), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18033) );
  AOI22_X1 U21312 ( .A1(n18018), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18032) );
  AOI22_X1 U21313 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18031) );
  NAND4_X1 U21314 ( .A1(n18034), .A2(n18033), .A3(n18032), .A4(n18031), .ZN(
        n18035) );
  NOR2_X1 U21315 ( .A1(n18036), .A2(n18035), .ZN(n18210) );
  OAI22_X1 U21316 ( .A1(n9746), .A2(n18037), .B1(n18210), .B2(n18101), .ZN(
        P3_U2693) );
  AOI22_X1 U21317 ( .A1(n13202), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18042) );
  AOI22_X1 U21318 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n18041) );
  AOI22_X1 U21319 ( .A1(n18018), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n9594), .ZN(n18040) );
  AOI22_X1 U21320 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18038), .B1(
        n13253), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18039) );
  NAND4_X1 U21321 ( .A1(n18042), .A2(n18041), .A3(n18040), .A4(n18039), .ZN(
        n18052) );
  AOI22_X1 U21322 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18044), .B1(
        n18043), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18050) );
  AOI22_X1 U21323 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18046), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n18045), .ZN(n18049) );
  AOI22_X1 U21324 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18062), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18048) );
  AOI22_X1 U21325 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n9590), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n18065), .ZN(n18047) );
  NAND4_X1 U21326 ( .A1(n18050), .A2(n18049), .A3(n18048), .A4(n18047), .ZN(
        n18051) );
  NOR2_X1 U21327 ( .A1(n18052), .A2(n18051), .ZN(n18215) );
  OAI21_X1 U21328 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n18055), .A(n18053), .ZN(
        n18054) );
  AOI22_X1 U21329 ( .A1(n18106), .A2(n18215), .B1(n18054), .B2(n18101), .ZN(
        P3_U2694) );
  AOI21_X1 U21330 ( .B1(n18057), .B2(n18056), .A(n18055), .ZN(n18076) );
  AOI22_X1 U21331 ( .A1(n16999), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18058), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18075) );
  AOI22_X1 U21332 ( .A1(n13081), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18059), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18074) );
  AOI22_X1 U21333 ( .A1(n18010), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18060) );
  OAI21_X1 U21334 ( .B1(n9592), .B2(n18061), .A(n18060), .ZN(n18072) );
  AOI22_X1 U21335 ( .A1(n18062), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9594), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18070) );
  AOI22_X1 U21336 ( .A1(n18063), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9590), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18069) );
  AOI22_X1 U21337 ( .A1(n18065), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18064), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18068) );
  AOI22_X1 U21338 ( .A1(n9589), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18066), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18067) );
  NAND4_X1 U21339 ( .A1(n18070), .A2(n18069), .A3(n18068), .A4(n18067), .ZN(
        n18071) );
  AOI211_X1 U21340 ( .C1(n17945), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n18072), .B(n18071), .ZN(n18073) );
  NAND3_X1 U21341 ( .A1(n18075), .A2(n18074), .A3(n18073), .ZN(n18218) );
  MUX2_X1 U21342 ( .A(n18076), .B(n18218), .S(n18106), .Z(P3_U2695) );
  NAND3_X1 U21343 ( .A1(n19084), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n18080), .ZN(
        n18079) );
  NAND3_X1 U21344 ( .A1(n18079), .A2(P3_EBX_REG_7__SCAN_IN), .A3(n18101), .ZN(
        n18077) );
  OAI221_X1 U21345 ( .B1(n18079), .B2(P3_EBX_REG_7__SCAN_IN), .C1(n18101), 
        .C2(n18078), .A(n18077), .ZN(P3_U2696) );
  NAND2_X1 U21346 ( .A1(n19084), .A2(n18080), .ZN(n18082) );
  NOR2_X1 U21347 ( .A1(n18106), .A2(n18080), .ZN(n18083) );
  AOI22_X1 U21348 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18106), .B1(
        P3_EBX_REG_6__SCAN_IN), .B2(n18083), .ZN(n18081) );
  OAI21_X1 U21349 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n18082), .A(n18081), .ZN(
        P3_U2697) );
  OAI21_X1 U21350 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n18084), .A(n18083), .ZN(
        n18085) );
  OAI21_X1 U21351 ( .B1(n18101), .B2(n18086), .A(n18085), .ZN(P3_U2698) );
  INV_X1 U21352 ( .A(n18105), .ZN(n18103) );
  NAND2_X1 U21353 ( .A1(n19084), .A2(n18103), .ZN(n18108) );
  NOR2_X1 U21354 ( .A1(n18087), .A2(n18108), .ZN(n18098) );
  NAND2_X1 U21355 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n18098), .ZN(n18093) );
  OAI21_X1 U21356 ( .B1(n18106), .B2(n18088), .A(n18093), .ZN(n18089) );
  OAI21_X1 U21357 ( .B1(n18108), .B2(n18090), .A(n18089), .ZN(n18091) );
  OAI21_X1 U21358 ( .B1(n18101), .B2(n18092), .A(n18091), .ZN(P3_U2699) );
  OAI211_X1 U21359 ( .C1(n18098), .C2(P3_EBX_REG_3__SCAN_IN), .A(n18101), .B(
        n18093), .ZN(n18094) );
  OAI21_X1 U21360 ( .B1(n18101), .B2(n18095), .A(n18094), .ZN(P3_U2700) );
  INV_X1 U21361 ( .A(n18096), .ZN(n18097) );
  AOI221_X1 U21362 ( .B1(n18097), .B2(n18103), .C1(n18213), .C2(n18103), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n18099) );
  AOI211_X1 U21363 ( .C1(n18106), .C2(n18100), .A(n18099), .B(n18098), .ZN(
        P3_U2701) );
  INV_X1 U21364 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18102) );
  OAI222_X1 U21365 ( .A1(n18108), .A2(n18104), .B1(n9973), .B2(n18103), .C1(
        n18102), .C2(n18101), .ZN(P3_U2702) );
  AOI22_X1 U21366 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18106), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n18105), .ZN(n18107) );
  OAI21_X1 U21367 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n18108), .A(n18107), .ZN(
        P3_U2703) );
  INV_X1 U21368 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n18324) );
  INV_X1 U21369 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18284) );
  INV_X1 U21370 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n21358) );
  INV_X1 U21371 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18316) );
  INV_X1 U21372 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18314) );
  INV_X1 U21373 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18259) );
  NOR2_X2 U21374 ( .A1(n19078), .A2(n18177), .ZN(n18182) );
  OAI21_X1 U21375 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n18246), .A(n18117), .ZN(
        n18110) );
  AOI22_X1 U21376 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18182), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n18110), .ZN(n18111) );
  OAI21_X1 U21377 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n18112), .A(n18111), .ZN(
        P3_U2704) );
  INV_X1 U21378 ( .A(n18182), .ZN(n18150) );
  OAI22_X1 U21379 ( .A1(n18114), .A2(n18237), .B1(n14696), .B2(n18150), .ZN(
        n18115) );
  AOI21_X1 U21380 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n18183), .A(n18115), .ZN(
        n18116) );
  OAI221_X1 U21381 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n18118), .C1(n18259), 
        .C2(n18117), .A(n18116), .ZN(P3_U2705) );
  AOI22_X1 U21382 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18183), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18182), .ZN(n18120) );
  OAI211_X1 U21383 ( .C1(n18123), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18177), .B(
        n18118), .ZN(n18119) );
  OAI211_X1 U21384 ( .C1(n18242), .C2(n18121), .A(n18120), .B(n18119), .ZN(
        P3_U2706) );
  INV_X1 U21385 ( .A(n18183), .ZN(n18156) );
  AOI22_X1 U21386 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18182), .B1(n18122), .B2(
        n18248), .ZN(n18127) );
  INV_X1 U21387 ( .A(n18123), .ZN(n18124) );
  OAI211_X1 U21388 ( .C1(n18125), .C2(P3_EAX_REG_28__SCAN_IN), .A(n18177), .B(
        n18124), .ZN(n18126) );
  OAI211_X1 U21389 ( .C1(n18156), .C2(n18349), .A(n18127), .B(n18126), .ZN(
        P3_U2707) );
  AOI22_X1 U21390 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18183), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18182), .ZN(n18130) );
  OAI211_X1 U21391 ( .C1(n9720), .C2(P3_EAX_REG_27__SCAN_IN), .A(n18177), .B(
        n18128), .ZN(n18129) );
  OAI211_X1 U21392 ( .C1(n18242), .C2(n18131), .A(n18130), .B(n18129), .ZN(
        P3_U2708) );
  AOI22_X1 U21393 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18183), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18182), .ZN(n18134) );
  AOI211_X1 U21394 ( .C1(n18324), .C2(n18136), .A(n9720), .B(n18194), .ZN(
        n18132) );
  INV_X1 U21395 ( .A(n18132), .ZN(n18133) );
  OAI211_X1 U21396 ( .C1(n18135), .C2(n18242), .A(n18134), .B(n18133), .ZN(
        P3_U2709) );
  AOI22_X1 U21397 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18183), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18182), .ZN(n18138) );
  OAI211_X1 U21398 ( .C1(n18141), .C2(P3_EAX_REG_25__SCAN_IN), .A(n18177), .B(
        n18136), .ZN(n18137) );
  OAI211_X1 U21399 ( .C1(n18139), .C2(n18242), .A(n18138), .B(n18137), .ZN(
        P3_U2710) );
  AOI22_X1 U21400 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18183), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18182), .ZN(n18144) );
  INV_X1 U21401 ( .A(n18141), .ZN(n18142) );
  OAI211_X1 U21402 ( .C1(n18140), .C2(P3_EAX_REG_24__SCAN_IN), .A(n18177), .B(
        n18142), .ZN(n18143) );
  OAI211_X1 U21403 ( .C1(n18145), .C2(n18237), .A(n18144), .B(n18143), .ZN(
        P3_U2711) );
  AOI22_X1 U21404 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18183), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18182), .ZN(n18148) );
  OAI211_X1 U21405 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n9731), .A(n18177), .B(
        n18146), .ZN(n18147) );
  OAI211_X1 U21406 ( .C1(n18149), .C2(n18237), .A(n18148), .B(n18147), .ZN(
        P3_U2712) );
  INV_X1 U21407 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18310) );
  INV_X1 U21408 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18308) );
  NAND2_X1 U21409 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18171), .ZN(n18167) );
  INV_X1 U21410 ( .A(n18167), .ZN(n18163) );
  NAND2_X1 U21411 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18163), .ZN(n18162) );
  NAND2_X1 U21412 ( .A1(n18177), .A2(n18162), .ZN(n18161) );
  OAI21_X1 U21413 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18246), .A(n18161), .ZN(
        n18154) );
  NOR3_X1 U21414 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18316), .A3(n18162), .ZN(
        n18153) );
  OAI22_X1 U21415 ( .A1(n18151), .A2(n18237), .B1(n16214), .B2(n18150), .ZN(
        n18152) );
  AOI211_X1 U21416 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n18154), .A(n18153), .B(
        n18152), .ZN(n18155) );
  OAI21_X1 U21417 ( .B1(n19077), .B2(n18156), .A(n18155), .ZN(P3_U2713) );
  AOI22_X1 U21418 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18182), .B1(n18248), .B2(
        n18157), .ZN(n18160) );
  INV_X1 U21419 ( .A(n18162), .ZN(n18158) );
  AOI22_X1 U21420 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18183), .B1(n18158), .B2(
        n18316), .ZN(n18159) );
  OAI211_X1 U21421 ( .C1(n18316), .C2(n18161), .A(n18160), .B(n18159), .ZN(
        P3_U2714) );
  AOI22_X1 U21422 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18183), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n18182), .ZN(n18165) );
  OAI211_X1 U21423 ( .C1(n18163), .C2(P3_EAX_REG_20__SCAN_IN), .A(n18177), .B(
        n18162), .ZN(n18164) );
  OAI211_X1 U21424 ( .C1(n18166), .C2(n18237), .A(n18165), .B(n18164), .ZN(
        P3_U2715) );
  AOI22_X1 U21425 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18183), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18182), .ZN(n18169) );
  OAI211_X1 U21426 ( .C1(n18171), .C2(P3_EAX_REG_19__SCAN_IN), .A(n18177), .B(
        n18167), .ZN(n18168) );
  OAI211_X1 U21427 ( .C1(n18170), .C2(n18237), .A(n18169), .B(n18168), .ZN(
        P3_U2716) );
  AOI22_X1 U21428 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18183), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18182), .ZN(n18174) );
  AOI211_X1 U21429 ( .C1(n18310), .C2(n18176), .A(n18171), .B(n18194), .ZN(
        n18172) );
  INV_X1 U21430 ( .A(n18172), .ZN(n18173) );
  OAI211_X1 U21431 ( .C1(n18175), .C2(n18237), .A(n18174), .B(n18173), .ZN(
        P3_U2717) );
  AOI22_X1 U21432 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18183), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18182), .ZN(n18180) );
  INV_X1 U21433 ( .A(n18184), .ZN(n18178) );
  OAI211_X1 U21434 ( .C1(n18178), .C2(P3_EAX_REG_17__SCAN_IN), .A(n18177), .B(
        n18176), .ZN(n18179) );
  OAI211_X1 U21435 ( .C1(n18181), .C2(n18237), .A(n18180), .B(n18179), .ZN(
        P3_U2718) );
  AOI22_X1 U21436 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18183), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n18182), .ZN(n18186) );
  OAI211_X1 U21437 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n18188), .A(n18177), .B(
        n18184), .ZN(n18185) );
  OAI211_X1 U21438 ( .C1(n18187), .C2(n18237), .A(n18186), .B(n18185), .ZN(
        P3_U2719) );
  AOI21_X1 U21439 ( .B1(n21358), .B2(n18189), .A(n18188), .ZN(n18190) );
  AOI22_X1 U21440 ( .A1(n18249), .A2(BUF2_REG_15__SCAN_IN), .B1(n18190), .B2(
        n18177), .ZN(n18191) );
  OAI21_X1 U21441 ( .B1(n18192), .B2(n18237), .A(n18191), .ZN(P3_U2720) );
  INV_X1 U21442 ( .A(n18193), .ZN(n18195) );
  OAI33_X1 U21443 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n18213), .A3(n18195), 
        .B1(n10209), .B2(n18194), .B3(n18193), .ZN(n18196) );
  AOI21_X1 U21444 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n18249), .A(n18196), .ZN(
        n18197) );
  OAI21_X1 U21445 ( .B1(n18198), .B2(n18237), .A(n18197), .ZN(P3_U2721) );
  INV_X1 U21446 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18347) );
  NOR3_X1 U21447 ( .A1(n18213), .A2(n18284), .A3(n18219), .ZN(n18217) );
  NAND2_X1 U21448 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18217), .ZN(n18209) );
  NOR2_X1 U21449 ( .A1(n18347), .A2(n18209), .ZN(n18203) );
  NAND2_X1 U21450 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18203), .ZN(n18202) );
  NAND3_X1 U21451 ( .A1(n18177), .A2(P3_EAX_REG_13__SCAN_IN), .A3(n18202), 
        .ZN(n18201) );
  AOI22_X1 U21452 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18249), .B1(n18248), .B2(
        n18199), .ZN(n18200) );
  OAI211_X1 U21453 ( .C1(P3_EAX_REG_13__SCAN_IN), .C2(n18202), .A(n18201), .B(
        n18200), .ZN(P3_U2722) );
  INV_X1 U21454 ( .A(n18202), .ZN(n18206) );
  AOI21_X1 U21455 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n18177), .A(n18203), .ZN(
        n18205) );
  OAI222_X1 U21456 ( .A1(n18245), .A2(n18349), .B1(n18206), .B2(n18205), .C1(
        n18242), .C2(n18204), .ZN(P3_U2723) );
  NAND2_X1 U21457 ( .A1(n18177), .A2(n18209), .ZN(n18212) );
  AOI22_X1 U21458 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18249), .B1(n18248), .B2(
        n18207), .ZN(n18208) );
  OAI221_X1 U21459 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n18209), .C1(n18347), 
        .C2(n18212), .A(n18208), .ZN(P3_U2724) );
  NOR2_X1 U21460 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18217), .ZN(n18211) );
  OAI222_X1 U21461 ( .A1(n18245), .A2(n18345), .B1(n18212), .B2(n18211), .C1(
        n18242), .C2(n18210), .ZN(P3_U2725) );
  NOR2_X1 U21462 ( .A1(n18213), .A2(n18219), .ZN(n18214) );
  AOI21_X1 U21463 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n18177), .A(n18214), .ZN(
        n18216) );
  OAI222_X1 U21464 ( .A1(n18245), .A2(n18343), .B1(n18217), .B2(n18216), .C1(
        n18242), .C2(n18215), .ZN(P3_U2726) );
  AOI22_X1 U21465 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18249), .B1(n18248), .B2(
        n18218), .ZN(n18221) );
  OAI211_X1 U21466 ( .C1(P3_EAX_REG_8__SCAN_IN), .C2(n18224), .A(n18177), .B(
        n18219), .ZN(n18220) );
  NAND2_X1 U21467 ( .A1(n18221), .A2(n18220), .ZN(P3_U2727) );
  INV_X1 U21468 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18289) );
  INV_X1 U21469 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18294) );
  INV_X1 U21470 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18332) );
  INV_X1 U21471 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18303) );
  NOR3_X1 U21472 ( .A1(n18332), .A2(n18303), .A3(n18246), .ZN(n18240) );
  NAND2_X1 U21473 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18244), .ZN(n18232) );
  NAND2_X1 U21474 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18235), .ZN(n18225) );
  NOR2_X1 U21475 ( .A1(n18289), .A2(n18225), .ZN(n18228) );
  AOI21_X1 U21476 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n18177), .A(n18228), .ZN(
        n18223) );
  OAI222_X1 U21477 ( .A1(n18245), .A2(n19081), .B1(n18224), .B2(n18223), .C1(
        n18242), .C2(n18222), .ZN(P3_U2728) );
  INV_X1 U21478 ( .A(n18225), .ZN(n18231) );
  AOI21_X1 U21479 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n18177), .A(n18231), .ZN(
        n18227) );
  OAI222_X1 U21480 ( .A1(n19077), .A2(n18245), .B1(n18228), .B2(n18227), .C1(
        n18242), .C2(n18226), .ZN(P3_U2729) );
  AOI21_X1 U21481 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n18177), .A(n18235), .ZN(
        n18230) );
  OAI222_X1 U21482 ( .A1(n19073), .A2(n18245), .B1(n18231), .B2(n18230), .C1(
        n18242), .C2(n18229), .ZN(P3_U2730) );
  INV_X1 U21483 ( .A(n18232), .ZN(n18239) );
  AOI21_X1 U21484 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n18177), .A(n18239), .ZN(
        n18234) );
  OAI222_X1 U21485 ( .A1(n19069), .A2(n18245), .B1(n18235), .B2(n18234), .C1(
        n18237), .C2(n18233), .ZN(P3_U2731) );
  AOI21_X1 U21486 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n18177), .A(n18244), .ZN(
        n18238) );
  OAI222_X1 U21487 ( .A1(n19065), .A2(n18245), .B1(n18239), .B2(n18238), .C1(
        n18237), .C2(n18236), .ZN(P3_U2732) );
  AOI21_X1 U21488 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n18177), .A(n18240), .ZN(
        n18243) );
  OAI222_X1 U21489 ( .A1(n21446), .A2(n18245), .B1(n18244), .B2(n18243), .C1(
        n18242), .C2(n18241), .ZN(P3_U2733) );
  OR2_X1 U21490 ( .A1(n18303), .A2(n18246), .ZN(n18254) );
  AOI22_X1 U21491 ( .A1(n18249), .A2(BUF2_REG_1__SCAN_IN), .B1(n18248), .B2(
        n18247), .ZN(n18253) );
  OAI21_X1 U21492 ( .B1(n18251), .B2(n18250), .A(P3_EAX_REG_1__SCAN_IN), .ZN(
        n18252) );
  OAI211_X1 U21493 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n18254), .A(n18253), .B(
        n18252), .ZN(P3_U2734) );
  OR2_X1 U21494 ( .A1(n19656), .A2(n18720), .ZN(n18274) );
  NOR2_X1 U21495 ( .A1(n18292), .A2(n18256), .ZN(P3_U2736) );
  AOI22_X1 U21496 ( .A1(n18300), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18258) );
  OAI21_X1 U21497 ( .B1(n18259), .B2(n18272), .A(n18258), .ZN(P3_U2737) );
  INV_X1 U21498 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18328) );
  AOI22_X1 U21499 ( .A1(n18300), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18260) );
  OAI21_X1 U21500 ( .B1(n18328), .B2(n18272), .A(n18260), .ZN(P3_U2738) );
  INV_X1 U21501 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n21434) );
  AOI22_X1 U21502 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n21311), .B1(n18300), 
        .B2(P3_UWORD_REG_12__SCAN_IN), .ZN(n18261) );
  OAI21_X1 U21503 ( .B1(n18292), .B2(n21434), .A(n18261), .ZN(P3_U2739) );
  AOI22_X1 U21504 ( .A1(n18300), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18262) );
  OAI21_X1 U21505 ( .B1(n10203), .B2(n18272), .A(n18262), .ZN(P3_U2740) );
  INV_X2 U21506 ( .A(n18274), .ZN(n18300) );
  AOI22_X1 U21507 ( .A1(n18300), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18263) );
  OAI21_X1 U21508 ( .B1(n18324), .B2(n18272), .A(n18263), .ZN(P3_U2741) );
  AOI22_X1 U21509 ( .A1(n18300), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18264) );
  OAI21_X1 U21510 ( .B1(n10202), .B2(n18272), .A(n18264), .ZN(P3_U2742) );
  INV_X1 U21511 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n18321) );
  AOI22_X1 U21512 ( .A1(n18300), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18265) );
  OAI21_X1 U21513 ( .B1(n18321), .B2(n18272), .A(n18265), .ZN(P3_U2743) );
  AOI22_X1 U21514 ( .A1(n18300), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18266) );
  OAI21_X1 U21515 ( .B1(n10194), .B2(n18272), .A(n18266), .ZN(P3_U2744) );
  INV_X1 U21516 ( .A(P3_UWORD_REG_6__SCAN_IN), .ZN(n21335) );
  AOI22_X1 U21517 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n21311), .B1(n21310), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18267) );
  OAI21_X1 U21518 ( .B1(n18274), .B2(n21335), .A(n18267), .ZN(P3_U2745) );
  AOI22_X1 U21519 ( .A1(n18300), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18268) );
  OAI21_X1 U21520 ( .B1(n18316), .B2(n18272), .A(n18268), .ZN(P3_U2746) );
  AOI22_X1 U21521 ( .A1(n18300), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18269) );
  OAI21_X1 U21522 ( .B1(n18314), .B2(n18272), .A(n18269), .ZN(P3_U2747) );
  INV_X1 U21523 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18312) );
  AOI22_X1 U21524 ( .A1(n18300), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18270) );
  OAI21_X1 U21525 ( .B1(n18312), .B2(n18272), .A(n18270), .ZN(P3_U2748) );
  AOI22_X1 U21526 ( .A1(n18300), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18271) );
  OAI21_X1 U21527 ( .B1(n18310), .B2(n18272), .A(n18271), .ZN(P3_U2749) );
  INV_X1 U21528 ( .A(P3_UWORD_REG_0__SCAN_IN), .ZN(n21339) );
  AOI22_X1 U21529 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n21311), .B1(n21310), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18273) );
  OAI21_X1 U21530 ( .B1(n18274), .B2(n21339), .A(n18273), .ZN(P3_U2751) );
  AOI22_X1 U21531 ( .A1(n18300), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18275) );
  OAI21_X1 U21532 ( .B1(n21358), .B2(n18302), .A(n18275), .ZN(P3_U2752) );
  AOI22_X1 U21533 ( .A1(n18300), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18276) );
  OAI21_X1 U21534 ( .B1(n10209), .B2(n18302), .A(n18276), .ZN(P3_U2753) );
  INV_X1 U21535 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18351) );
  AOI22_X1 U21536 ( .A1(n18300), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18277) );
  OAI21_X1 U21537 ( .B1(n18351), .B2(n18302), .A(n18277), .ZN(P3_U2754) );
  INV_X1 U21538 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18279) );
  AOI22_X1 U21539 ( .A1(n18300), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18278) );
  OAI21_X1 U21540 ( .B1(n18279), .B2(n18302), .A(n18278), .ZN(P3_U2755) );
  AOI22_X1 U21541 ( .A1(n18300), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18280) );
  OAI21_X1 U21542 ( .B1(n18347), .B2(n18302), .A(n18280), .ZN(P3_U2756) );
  INV_X1 U21543 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18282) );
  AOI22_X1 U21544 ( .A1(n18300), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18281) );
  OAI21_X1 U21545 ( .B1(n18282), .B2(n18302), .A(n18281), .ZN(P3_U2757) );
  AOI22_X1 U21546 ( .A1(n18300), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18283) );
  OAI21_X1 U21547 ( .B1(n18284), .B2(n18302), .A(n18283), .ZN(P3_U2758) );
  AOI22_X1 U21548 ( .A1(n18300), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18285) );
  OAI21_X1 U21549 ( .B1(n10211), .B2(n18302), .A(n18285), .ZN(P3_U2759) );
  INV_X1 U21550 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18287) );
  AOI22_X1 U21551 ( .A1(n18300), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18286) );
  OAI21_X1 U21552 ( .B1(n18287), .B2(n18302), .A(n18286), .ZN(P3_U2760) );
  AOI22_X1 U21553 ( .A1(n18300), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18288) );
  OAI21_X1 U21554 ( .B1(n18289), .B2(n18302), .A(n18288), .ZN(P3_U2761) );
  INV_X1 U21555 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18291) );
  AOI22_X1 U21556 ( .A1(n18300), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18290) );
  OAI21_X1 U21557 ( .B1(n18291), .B2(n18302), .A(n18290), .ZN(P3_U2762) );
  INV_X2 U21558 ( .A(n18292), .ZN(n21310) );
  AOI22_X1 U21559 ( .A1(n18300), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18293) );
  OAI21_X1 U21560 ( .B1(n18294), .B2(n18302), .A(n18293), .ZN(P3_U2763) );
  INV_X1 U21561 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18296) );
  AOI22_X1 U21562 ( .A1(n18300), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18295) );
  OAI21_X1 U21563 ( .B1(n18296), .B2(n18302), .A(n18295), .ZN(P3_U2764) );
  INV_X1 U21564 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18298) );
  AOI22_X1 U21565 ( .A1(n18300), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18297) );
  OAI21_X1 U21566 ( .B1(n18298), .B2(n18302), .A(n18297), .ZN(P3_U2765) );
  AOI22_X1 U21567 ( .A1(n18300), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18299) );
  OAI21_X1 U21568 ( .B1(n18332), .B2(n18302), .A(n18299), .ZN(P3_U2766) );
  AOI22_X1 U21569 ( .A1(n18300), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n21310), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18301) );
  OAI21_X1 U21570 ( .B1(n18303), .B2(n18302), .A(n18301), .ZN(P3_U2767) );
  INV_X1 U21571 ( .A(n19702), .ZN(n19693) );
  NOR2_X2 U21572 ( .A1(n19059), .A2(n18341), .ZN(n18356) );
  NOR3_X4 U21573 ( .A1(n19691), .A2(n18305), .A3(n18304), .ZN(n18352) );
  AOI22_X1 U21574 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18356), .B1(
        P3_EAX_REG_16__SCAN_IN), .B2(n18352), .ZN(n18306) );
  OAI21_X1 U21575 ( .B1(n18318), .B2(n21339), .A(n18306), .ZN(P3_U2768) );
  AOI22_X1 U21576 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18356), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18341), .ZN(n18307) );
  OAI21_X1 U21577 ( .B1(n18308), .B2(n18358), .A(n18307), .ZN(P3_U2769) );
  AOI22_X1 U21578 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18356), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18341), .ZN(n18309) );
  OAI21_X1 U21579 ( .B1(n18310), .B2(n18358), .A(n18309), .ZN(P3_U2770) );
  AOI22_X1 U21580 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18356), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18341), .ZN(n18311) );
  OAI21_X1 U21581 ( .B1(n18312), .B2(n18358), .A(n18311), .ZN(P3_U2771) );
  AOI22_X1 U21582 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18356), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18341), .ZN(n18313) );
  OAI21_X1 U21583 ( .B1(n18314), .B2(n18358), .A(n18313), .ZN(P3_U2772) );
  AOI22_X1 U21584 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18356), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18341), .ZN(n18315) );
  OAI21_X1 U21585 ( .B1(n18316), .B2(n18358), .A(n18315), .ZN(P3_U2773) );
  AOI22_X1 U21586 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n18356), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n18352), .ZN(n18317) );
  OAI21_X1 U21587 ( .B1(n18318), .B2(n21335), .A(n18317), .ZN(P3_U2774) );
  AOI22_X1 U21588 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18356), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18341), .ZN(n18319) );
  OAI21_X1 U21589 ( .B1(n10194), .B2(n18358), .A(n18319), .ZN(P3_U2775) );
  AOI22_X1 U21590 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18356), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18341), .ZN(n18320) );
  OAI21_X1 U21591 ( .B1(n18321), .B2(n18358), .A(n18320), .ZN(P3_U2776) );
  AOI22_X1 U21592 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18356), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18341), .ZN(n18322) );
  OAI21_X1 U21593 ( .B1(n10202), .B2(n18358), .A(n18322), .ZN(P3_U2777) );
  AOI22_X1 U21594 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18356), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18341), .ZN(n18323) );
  OAI21_X1 U21595 ( .B1(n18324), .B2(n18358), .A(n18323), .ZN(P3_U2778) );
  AOI22_X1 U21596 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18356), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18341), .ZN(n18325) );
  OAI21_X1 U21597 ( .B1(n10203), .B2(n18358), .A(n18325), .ZN(P3_U2779) );
  AOI22_X1 U21598 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n18352), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18341), .ZN(n18326) );
  OAI21_X1 U21599 ( .B1(n18349), .B2(n18354), .A(n18326), .ZN(P3_U2780) );
  AOI22_X1 U21600 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18356), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18355), .ZN(n18327) );
  OAI21_X1 U21601 ( .B1(n18328), .B2(n18358), .A(n18327), .ZN(P3_U2781) );
  AOI22_X1 U21602 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n18352), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18355), .ZN(n18329) );
  OAI21_X1 U21603 ( .B1(n21382), .B2(n18354), .A(n18329), .ZN(P3_U2782) );
  AOI22_X1 U21604 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18352), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18355), .ZN(n18330) );
  OAI21_X1 U21605 ( .B1(n21451), .B2(n18354), .A(n18330), .ZN(P3_U2783) );
  AOI22_X1 U21606 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18356), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18355), .ZN(n18331) );
  OAI21_X1 U21607 ( .B1(n18332), .B2(n18358), .A(n18331), .ZN(P3_U2784) );
  AOI22_X1 U21608 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18352), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18355), .ZN(n18333) );
  OAI21_X1 U21609 ( .B1(n21446), .B2(n18354), .A(n18333), .ZN(P3_U2785) );
  AOI22_X1 U21610 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18352), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18355), .ZN(n18334) );
  OAI21_X1 U21611 ( .B1(n19065), .B2(n18354), .A(n18334), .ZN(P3_U2786) );
  AOI22_X1 U21612 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18352), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18355), .ZN(n18335) );
  OAI21_X1 U21613 ( .B1(n19069), .B2(n18354), .A(n18335), .ZN(P3_U2787) );
  AOI22_X1 U21614 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18352), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18341), .ZN(n18336) );
  OAI21_X1 U21615 ( .B1(n19073), .B2(n18354), .A(n18336), .ZN(P3_U2788) );
  AOI22_X1 U21616 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18352), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18341), .ZN(n18337) );
  OAI21_X1 U21617 ( .B1(n19077), .B2(n18354), .A(n18337), .ZN(P3_U2789) );
  AOI22_X1 U21618 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n18352), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18341), .ZN(n18338) );
  OAI21_X1 U21619 ( .B1(n19081), .B2(n18354), .A(n18338), .ZN(P3_U2790) );
  AOI22_X1 U21620 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18352), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18341), .ZN(n18339) );
  OAI21_X1 U21621 ( .B1(n18340), .B2(n18354), .A(n18339), .ZN(P3_U2791) );
  AOI22_X1 U21622 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18352), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18341), .ZN(n18342) );
  OAI21_X1 U21623 ( .B1(n18343), .B2(n18354), .A(n18342), .ZN(P3_U2792) );
  AOI22_X1 U21624 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18352), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18355), .ZN(n18344) );
  OAI21_X1 U21625 ( .B1(n18345), .B2(n18354), .A(n18344), .ZN(P3_U2793) );
  AOI22_X1 U21626 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18356), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18355), .ZN(n18346) );
  OAI21_X1 U21627 ( .B1(n18347), .B2(n18358), .A(n18346), .ZN(P3_U2794) );
  AOI22_X1 U21628 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18352), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18355), .ZN(n18348) );
  OAI21_X1 U21629 ( .B1(n18349), .B2(n18354), .A(n18348), .ZN(P3_U2795) );
  AOI22_X1 U21630 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18356), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18355), .ZN(n18350) );
  OAI21_X1 U21631 ( .B1(n18351), .B2(n18358), .A(n18350), .ZN(P3_U2796) );
  AOI22_X1 U21632 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n18352), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18355), .ZN(n18353) );
  OAI21_X1 U21633 ( .B1(n21382), .B2(n18354), .A(n18353), .ZN(P3_U2797) );
  AOI22_X1 U21634 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18356), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18355), .ZN(n18357) );
  OAI21_X1 U21635 ( .B1(n21358), .B2(n18358), .A(n18357), .ZN(P3_U2798) );
  INV_X1 U21636 ( .A(n9585), .ZN(n18673) );
  OAI22_X1 U21637 ( .A1(n18360), .A2(n18628), .B1(n18359), .B2(n18720), .ZN(
        n18361) );
  NOR2_X1 U21638 ( .A1(n18673), .A2(n18361), .ZN(n18396) );
  OAI21_X1 U21639 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18441), .A(
        n18396), .ZN(n18386) );
  AOI22_X1 U21640 ( .A1(n18578), .A2(n18362), .B1(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n18386), .ZN(n18380) );
  INV_X1 U21641 ( .A(n18363), .ZN(n18374) );
  AOI21_X1 U21642 ( .B1(n18365), .B2(n18364), .A(n18609), .ZN(n18373) );
  INV_X1 U21643 ( .A(n18731), .ZN(n18366) );
  OAI22_X1 U21644 ( .A1(n18366), .A2(n18725), .B1(n18733), .B2(n18593), .ZN(
        n18400) );
  NOR2_X1 U21645 ( .A1(n18734), .A2(n18400), .ZN(n18368) );
  AOI211_X1 U21646 ( .C1(n18725), .C2(n18593), .A(n18368), .B(n18367), .ZN(
        n18371) );
  NAND2_X1 U21647 ( .A1(n9586), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n18378) );
  NOR2_X1 U21648 ( .A1(n18523), .A2(n18375), .ZN(n18388) );
  OAI211_X1 U21649 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n18388), .B(n18376), .ZN(n18377) );
  NAND4_X1 U21650 ( .A1(n18380), .A2(n18379), .A3(n18378), .A4(n18377), .ZN(
        P3_U2802) );
  NAND2_X1 U21651 ( .A1(n9821), .A2(n18382), .ZN(n18383) );
  XNOR2_X1 U21652 ( .A(n18634), .B(n18383), .ZN(n18739) );
  INV_X1 U21653 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19627) );
  OAI22_X1 U21654 ( .A1(n19024), .A2(n19627), .B1(n18566), .B2(n18384), .ZN(
        n18385) );
  AOI221_X1 U21655 ( .B1(n18388), .B2(n18387), .C1(n18386), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n18385), .ZN(n18391) );
  AOI22_X1 U21656 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18400), .B1(
        n18389), .B2(n18734), .ZN(n18390) );
  OAI211_X1 U21657 ( .C1(n18739), .C2(n18609), .A(n18391), .B(n18390), .ZN(
        P3_U2803) );
  AOI21_X1 U21658 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n18393), .A(
        n18392), .ZN(n18743) );
  INV_X1 U21659 ( .A(n18441), .ZN(n18398) );
  AOI21_X1 U21660 ( .B1(n18394), .B2(n19427), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18395) );
  OAI22_X1 U21661 ( .A1(n18396), .A2(n18395), .B1(n19024), .B2(n21372), .ZN(
        n18397) );
  AOI221_X1 U21662 ( .B1(n18578), .B2(n18399), .C1(n18398), .C2(n18399), .A(
        n18397), .ZN(n18402) );
  NOR3_X1 U21663 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18409), .A3(
        n18729), .ZN(n18741) );
  NOR2_X1 U21664 ( .A1(n18726), .A2(n18531), .ZN(n18439) );
  AOI22_X1 U21665 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18400), .B1(
        n18741), .B2(n18439), .ZN(n18401) );
  OAI211_X1 U21666 ( .C1(n18743), .C2(n18609), .A(n18402), .B(n18401), .ZN(
        P3_U2804) );
  AND2_X1 U21667 ( .A1(n18412), .A2(n19427), .ZN(n18432) );
  AOI211_X1 U21668 ( .C1(n18443), .C2(n18403), .A(n18673), .B(n18432), .ZN(
        n18436) );
  OAI21_X1 U21669 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18441), .A(
        n18436), .ZN(n18422) );
  AOI22_X1 U21670 ( .A1(n18578), .A2(n18404), .B1(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18422), .ZN(n18416) );
  XNOR2_X1 U21671 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n18405), .ZN(
        n18758) );
  XNOR2_X1 U21672 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n18406), .ZN(
        n18760) );
  OAI21_X1 U21673 ( .B1(n10142), .B2(n18408), .A(n18407), .ZN(n18410) );
  XNOR2_X1 U21674 ( .A(n18410), .B(n18409), .ZN(n18756) );
  OAI22_X1 U21675 ( .A1(n18725), .A2(n18760), .B1(n18609), .B2(n18756), .ZN(
        n18411) );
  AOI21_X1 U21676 ( .B1(n18636), .B2(n18758), .A(n18411), .ZN(n18415) );
  NAND2_X1 U21677 ( .A1(n9586), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18754) );
  NOR2_X1 U21678 ( .A1(n18523), .A2(n18412), .ZN(n18424) );
  OAI211_X1 U21679 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n18424), .B(n18413), .ZN(n18414) );
  NAND4_X1 U21680 ( .A1(n18416), .A2(n18415), .A3(n18754), .A4(n18414), .ZN(
        P3_U2805) );
  AOI21_X1 U21681 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18418), .A(
        n18417), .ZN(n18774) );
  AOI22_X1 U21682 ( .A1(n9586), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n18578), 
        .B2(n18419), .ZN(n18420) );
  INV_X1 U21683 ( .A(n18420), .ZN(n18421) );
  AOI221_X1 U21684 ( .B1(n18424), .B2(n18423), .C1(n18422), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18421), .ZN(n18426) );
  NOR2_X1 U21685 ( .A1(n18532), .A2(n9745), .ZN(n18763) );
  NOR2_X1 U21686 ( .A1(n18859), .A2(n9745), .ZN(n18762) );
  OAI22_X1 U21687 ( .A1(n18763), .A2(n18593), .B1(n18762), .B2(n18725), .ZN(
        n18438) );
  NOR2_X1 U21688 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n9745), .ZN(
        n18771) );
  AOI22_X1 U21689 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18438), .B1(
        n18459), .B2(n18771), .ZN(n18425) );
  OAI211_X1 U21690 ( .C1(n18774), .C2(n18609), .A(n18426), .B(n18425), .ZN(
        P3_U2806) );
  AOI22_X1 U21691 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n10142), .B1(
        n18428), .B2(n18452), .ZN(n18429) );
  NAND2_X1 U21692 ( .A1(n18427), .A2(n18429), .ZN(n18430) );
  XNOR2_X1 U21693 ( .A(n18430), .B(n18767), .ZN(n18779) );
  NAND2_X2 U21694 ( .A1(n18566), .A2(n18441), .ZN(n18715) );
  AOI22_X1 U21695 ( .A1(n18433), .A2(n18432), .B1(n18431), .B2(n18715), .ZN(
        n18434) );
  NAND2_X1 U21696 ( .A1(n9586), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18778) );
  OAI211_X1 U21697 ( .C1(n18436), .C2(n18435), .A(n18434), .B(n18778), .ZN(
        n18437) );
  AOI221_X1 U21698 ( .B1(n18439), .B2(n18767), .C1(n18438), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n18437), .ZN(n18440) );
  OAI21_X1 U21699 ( .B1(n18609), .B2(n18779), .A(n18440), .ZN(P3_U2807) );
  NAND2_X1 U21700 ( .A1(n18792), .A2(n18459), .ZN(n18458) );
  NOR2_X1 U21701 ( .A1(n19024), .A2(n19617), .ZN(n18794) );
  AOI22_X1 U21702 ( .A1(n18693), .A2(n18444), .B1(n18443), .B2(n18442), .ZN(
        n18445) );
  NAND2_X1 U21703 ( .A1(n18445), .A2(n9585), .ZN(n18478) );
  AOI21_X1 U21704 ( .B1(n18398), .B2(n18472), .A(n18478), .ZN(n18460) );
  NAND2_X1 U21705 ( .A1(n18446), .A2(n18561), .ZN(n18462) );
  OAI21_X1 U21706 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n18447), .ZN(n18448) );
  OAI22_X1 U21707 ( .A1(n18460), .A2(n18449), .B1(n18462), .B2(n18448), .ZN(
        n18450) );
  AOI211_X1 U21708 ( .C1(n18451), .C2(n18578), .A(n18794), .B(n18450), .ZN(
        n18457) );
  INV_X1 U21709 ( .A(n18725), .ZN(n18713) );
  NOR2_X1 U21710 ( .A1(n18713), .A2(n18636), .ZN(n18479) );
  AOI22_X1 U21711 ( .A1(n18713), .A2(n18859), .B1(n18636), .B2(n18532), .ZN(
        n18530) );
  OAI21_X1 U21712 ( .B1(n18792), .B2(n18479), .A(n18530), .ZN(n18468) );
  INV_X1 U21713 ( .A(n18452), .ZN(n18454) );
  OAI221_X1 U21714 ( .B1(n18454), .B2(n18453), .C1(n18454), .C2(n18792), .A(
        n18427), .ZN(n18455) );
  XNOR2_X1 U21715 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n18455), .ZN(
        n18793) );
  AOI22_X1 U21716 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18468), .B1(
        n18635), .B2(n18793), .ZN(n18456) );
  OAI211_X1 U21717 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n18458), .A(
        n18457), .B(n18456), .ZN(P3_U2808) );
  NAND2_X1 U21718 ( .A1(n18803), .A2(n18800), .ZN(n18809) );
  INV_X1 U21719 ( .A(n18782), .ZN(n18799) );
  NAND2_X1 U21720 ( .A1(n18799), .A2(n18459), .ZN(n18496) );
  INV_X1 U21721 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18461) );
  NAND2_X1 U21722 ( .A1(n9586), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n18807) );
  OAI221_X1 U21723 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n18462), .C1(
        n18461), .C2(n18460), .A(n18807), .ZN(n18463) );
  AOI21_X1 U21724 ( .B1(n18578), .B2(n18464), .A(n18463), .ZN(n18470) );
  INV_X1 U21725 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18497) );
  NOR3_X1 U21726 ( .A1(n18497), .A2(n10142), .A3(n18465), .ZN(n18490) );
  INV_X1 U21727 ( .A(n18504), .ZN(n18491) );
  AOI22_X1 U21728 ( .A1(n18803), .A2(n18490), .B1(n18491), .B2(n18466), .ZN(
        n18467) );
  XNOR2_X1 U21729 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18467), .ZN(
        n18806) );
  AOI22_X1 U21730 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18468), .B1(
        n18635), .B2(n18806), .ZN(n18469) );
  OAI211_X1 U21731 ( .C1(n18809), .C2(n18496), .A(n18470), .B(n18469), .ZN(
        P3_U2809) );
  NAND2_X1 U21732 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18471), .ZN(
        n18819) );
  OAI21_X1 U21733 ( .B1(n17432), .B2(n19335), .A(n18472), .ZN(n18477) );
  INV_X1 U21734 ( .A(n18473), .ZN(n18474) );
  AOI21_X1 U21735 ( .B1(n18566), .B2(n18441), .A(n18474), .ZN(n18476) );
  NOR2_X1 U21736 ( .A1(n19024), .A2(n19614), .ZN(n18475) );
  AOI211_X1 U21737 ( .C1(n18478), .C2(n18477), .A(n18476), .B(n18475), .ZN(
        n18483) );
  NOR2_X1 U21738 ( .A1(n18782), .A2(n18480), .ZN(n18811) );
  OAI21_X1 U21739 ( .B1(n18479), .B2(n18811), .A(n18530), .ZN(n18493) );
  OAI221_X1 U21740 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18503), 
        .C1(n18480), .C2(n18490), .A(n18427), .ZN(n18481) );
  XNOR2_X1 U21741 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n18481), .ZN(
        n18810) );
  AOI22_X1 U21742 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18493), .B1(
        n18635), .B2(n18810), .ZN(n18482) );
  OAI211_X1 U21743 ( .C1(n18496), .C2(n18819), .A(n18483), .B(n18482), .ZN(
        P3_U2810) );
  AOI21_X1 U21744 ( .B1(n18693), .B2(n18485), .A(n18673), .ZN(n18509) );
  OAI21_X1 U21745 ( .B1(n18484), .B2(n18720), .A(n18509), .ZN(n18500) );
  NAND2_X1 U21746 ( .A1(n9586), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18822) );
  NOR2_X1 U21747 ( .A1(n18523), .A2(n18485), .ZN(n18502) );
  OAI211_X1 U21748 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n18502), .B(n18486), .ZN(n18487) );
  OAI211_X1 U21749 ( .C1(n18566), .C2(n18488), .A(n18822), .B(n18487), .ZN(
        n18489) );
  AOI21_X1 U21750 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18500), .A(
        n18489), .ZN(n18495) );
  AOI21_X1 U21751 ( .B1(n18503), .B2(n18491), .A(n18490), .ZN(n18492) );
  XNOR2_X1 U21752 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n18492), .ZN(
        n18820) );
  AOI22_X1 U21753 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18493), .B1(
        n18635), .B2(n18820), .ZN(n18494) );
  OAI211_X1 U21754 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18496), .A(
        n18495), .B(n18494), .ZN(P3_U2811) );
  NAND2_X1 U21755 ( .A1(n18830), .A2(n18497), .ZN(n18838) );
  NAND2_X1 U21756 ( .A1(n9586), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18836) );
  OAI21_X1 U21757 ( .B1(n18566), .B2(n18498), .A(n18836), .ZN(n18499) );
  AOI221_X1 U21758 ( .B1(n18502), .B2(n18501), .C1(n18500), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n18499), .ZN(n18507) );
  OAI21_X1 U21759 ( .B1(n18830), .B2(n18531), .A(n18530), .ZN(n18515) );
  AOI21_X1 U21760 ( .B1(n18634), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n18503), .ZN(n18505) );
  XNOR2_X1 U21761 ( .A(n18505), .B(n18504), .ZN(n18834) );
  AOI22_X1 U21762 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18515), .B1(
        n18635), .B2(n18834), .ZN(n18506) );
  OAI211_X1 U21763 ( .C1(n18531), .C2(n18838), .A(n18507), .B(n18506), .ZN(
        P3_U2812) );
  NAND2_X1 U21764 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18839), .ZN(
        n18845) );
  AOI21_X1 U21765 ( .B1(n18508), .B2(n19427), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18510) );
  OAI22_X1 U21766 ( .A1(n18510), .A2(n18509), .B1(n19024), .B2(n19607), .ZN(
        n18511) );
  AOI21_X1 U21767 ( .B1(n18512), .B2(n18715), .A(n18511), .ZN(n18517) );
  OAI21_X1 U21768 ( .B1(n18513), .B2(n18839), .A(n18514), .ZN(n18843) );
  AOI22_X1 U21769 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18515), .B1(
        n18635), .B2(n18843), .ZN(n18516) );
  OAI211_X1 U21770 ( .C1(n18531), .C2(n18845), .A(n18517), .B(n18516), .ZN(
        P3_U2813) );
  AOI21_X1 U21771 ( .B1(n18634), .B2(n18518), .A(n18519), .ZN(n18520) );
  XNOR2_X1 U21772 ( .A(n18520), .B(n18856), .ZN(n18853) );
  AOI21_X1 U21773 ( .B1(n18693), .B2(n18522), .A(n18673), .ZN(n18559) );
  OAI21_X1 U21774 ( .B1(n18521), .B2(n18720), .A(n18559), .ZN(n18535) );
  AOI22_X1 U21775 ( .A1(n9586), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18535), .ZN(n18526) );
  NOR2_X1 U21776 ( .A1(n18523), .A2(n18522), .ZN(n18537) );
  OAI211_X1 U21777 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18537), .B(n18524), .ZN(n18525) );
  OAI211_X1 U21778 ( .C1(n18566), .C2(n18527), .A(n18526), .B(n18525), .ZN(
        n18528) );
  AOI21_X1 U21779 ( .B1(n18635), .B2(n18853), .A(n18528), .ZN(n18529) );
  OAI221_X1 U21780 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18531), 
        .C1(n18856), .C2(n18530), .A(n18529), .ZN(P3_U2814) );
  NOR2_X1 U21781 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18550), .ZN(
        n18866) );
  NAND2_X1 U21782 ( .A1(n18636), .A2(n18532), .ZN(n18547) );
  INV_X1 U21783 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18536) );
  OAI22_X1 U21784 ( .A1(n19024), .A2(n19603), .B1(n18566), .B2(n18533), .ZN(
        n18534) );
  AOI221_X1 U21785 ( .B1(n18537), .B2(n18536), .C1(n18535), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n18534), .ZN(n18546) );
  NAND2_X1 U21786 ( .A1(n18538), .A2(n10142), .ZN(n18611) );
  NOR3_X1 U21787 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18605), .A3(
        n18611), .ZN(n18573) );
  NOR3_X1 U21788 ( .A1(n18903), .A2(n18876), .A3(n18539), .ZN(n18541) );
  AOI22_X1 U21789 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n10142), .B1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n21454), .ZN(n18540) );
  OAI221_X1 U21790 ( .B1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n18573), 
        .C1(n10233), .C2(n18541), .A(n18540), .ZN(n18542) );
  XNOR2_X1 U21791 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18542), .ZN(
        n18867) );
  NOR2_X1 U21792 ( .A1(n18786), .A2(n18725), .ZN(n18544) );
  NAND2_X1 U21793 ( .A1(n18554), .A2(n18543), .ZN(n18858) );
  AOI22_X1 U21794 ( .A1(n18635), .A2(n18867), .B1(n18544), .B2(n18858), .ZN(
        n18545) );
  OAI211_X1 U21795 ( .C1(n18866), .C2(n18547), .A(n18546), .B(n18545), .ZN(
        P3_U2815) );
  INV_X1 U21796 ( .A(n17434), .ZN(n18548) );
  NOR2_X1 U21797 ( .A1(n18548), .A2(n19335), .ZN(n18591) );
  AOI21_X1 U21798 ( .B1(n18562), .B2(n18591), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18558) );
  AOI22_X1 U21799 ( .A1(n9586), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n18549), 
        .B2(n18715), .ZN(n18557) );
  AOI221_X1 U21800 ( .B1(n18862), .B2(n18876), .C1(n13337), .C2(n18876), .A(
        n18550), .ZN(n18884) );
  NAND2_X1 U21801 ( .A1(n18634), .A2(n18911), .ZN(n18612) );
  NAND2_X1 U21802 ( .A1(n21454), .A2(n10233), .ZN(n18552) );
  INV_X1 U21803 ( .A(n18573), .ZN(n18551) );
  OAI22_X1 U21804 ( .A1(n18862), .A2(n18612), .B1(n18552), .B2(n18551), .ZN(
        n18553) );
  XNOR2_X1 U21805 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18553), .ZN(
        n18882) );
  INV_X1 U21806 ( .A(n18862), .ZN(n18874) );
  OAI221_X1 U21807 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18874), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18909), .A(n18554), .ZN(
        n18881) );
  OAI22_X1 U21808 ( .A1(n18882), .A2(n18609), .B1(n18725), .B2(n18881), .ZN(
        n18555) );
  AOI21_X1 U21809 ( .B1(n18636), .B2(n18884), .A(n18555), .ZN(n18556) );
  OAI211_X1 U21810 ( .C1(n18559), .C2(n18558), .A(n18557), .B(n18556), .ZN(
        P3_U2816) );
  NOR2_X1 U21811 ( .A1(n18903), .A2(n18612), .ZN(n18574) );
  AOI22_X1 U21812 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18574), .B1(
        n18573), .B2(n21454), .ZN(n18560) );
  XNOR2_X1 U21813 ( .A(n18560), .B(n10233), .ZN(n18898) );
  NAND2_X1 U21814 ( .A1(n17434), .A2(n18561), .ZN(n18582) );
  AOI211_X1 U21815 ( .C1(n18581), .C2(n18567), .A(n18562), .B(n18582), .ZN(
        n18569) );
  OAI21_X1 U21816 ( .B1(n17434), .B2(n18628), .A(n18720), .ZN(n18563) );
  AOI21_X1 U21817 ( .B1(n18564), .B2(n18563), .A(n18673), .ZN(n18580) );
  OAI22_X1 U21818 ( .A1(n18580), .A2(n18567), .B1(n18566), .B2(n18565), .ZN(
        n18568) );
  AOI211_X1 U21819 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n9586), .A(n18569), .B(
        n18568), .ZN(n18572) );
  INV_X1 U21820 ( .A(n18873), .ZN(n18899) );
  NOR2_X1 U21821 ( .A1(n18899), .A2(n13337), .ZN(n18890) );
  NAND2_X1 U21822 ( .A1(n18873), .A2(n18909), .ZN(n18892) );
  INV_X1 U21823 ( .A(n18892), .ZN(n18570) );
  OAI22_X1 U21824 ( .A1(n18890), .A2(n18593), .B1(n18570), .B2(n18725), .ZN(
        n18584) );
  NOR2_X1 U21825 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18899), .ZN(
        n18887) );
  AOI22_X1 U21826 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18584), .B1(
        n18887), .B2(n18576), .ZN(n18571) );
  OAI211_X1 U21827 ( .C1(n18898), .C2(n18609), .A(n18572), .B(n18571), .ZN(
        P3_U2817) );
  NOR2_X1 U21828 ( .A1(n18574), .A2(n18573), .ZN(n18575) );
  XNOR2_X1 U21829 ( .A(n18575), .B(n21454), .ZN(n18908) );
  INV_X1 U21830 ( .A(n18576), .ZN(n18621) );
  NOR2_X1 U21831 ( .A1(n18621), .A2(n18903), .ZN(n18585) );
  AOI22_X1 U21832 ( .A1(n9586), .A2(P3_REIP_REG_12__SCAN_IN), .B1(n18578), 
        .B2(n18577), .ZN(n18579) );
  OAI221_X1 U21833 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18582), .C1(
        n18581), .C2(n18580), .A(n18579), .ZN(n18583) );
  AOI221_X1 U21834 ( .B1(n18585), .B2(n21454), .C1(n18584), .C2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n18583), .ZN(n18586) );
  OAI21_X1 U21835 ( .B1(n18908), .B2(n18609), .A(n18586), .ZN(P3_U2818) );
  INV_X1 U21836 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18918) );
  NAND2_X1 U21837 ( .A1(n18916), .A2(n18918), .ZN(n18925) );
  INV_X1 U21838 ( .A(n18916), .ZN(n18599) );
  OAI22_X1 U21839 ( .A1(n18599), .A2(n18612), .B1(n18605), .B2(n18611), .ZN(
        n18587) );
  XNOR2_X1 U21840 ( .A(n18918), .B(n18587), .ZN(n18923) );
  NOR2_X1 U21841 ( .A1(n19024), .A2(n19595), .ZN(n18922) );
  NAND2_X1 U21842 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18588) );
  NOR3_X1 U21843 ( .A1(n17714), .A2(n18652), .A3(n19335), .ZN(n18640) );
  NAND2_X1 U21844 ( .A1(n18640), .A2(n18624), .ZN(n18600) );
  NOR2_X1 U21845 ( .A1(n18588), .A2(n18600), .ZN(n18602) );
  AOI21_X1 U21846 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18716), .A(
        n18602), .ZN(n18590) );
  OAI22_X1 U21847 ( .A1(n18591), .A2(n18590), .B1(n18707), .B2(n18589), .ZN(
        n18592) );
  AOI211_X1 U21848 ( .C1(n18635), .C2(n18923), .A(n18922), .B(n18592), .ZN(
        n18595) );
  NOR2_X1 U21849 ( .A1(n18916), .A2(n18621), .ZN(n18606) );
  OAI22_X1 U21850 ( .A1(n18911), .A2(n18593), .B1(n18725), .B2(n18909), .ZN(
        n18610) );
  OAI21_X1 U21851 ( .B1(n18606), .B2(n18610), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18594) );
  OAI211_X1 U21852 ( .C1(n18621), .C2(n18925), .A(n18595), .B(n18594), .ZN(
        P3_U2819) );
  OAI221_X1 U21853 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18611), .C1(
        n18940), .C2(n18612), .A(n18917), .ZN(n18598) );
  NAND4_X1 U21854 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18538), .A3(
        n18940), .A4(n10142), .ZN(n18597) );
  OAI211_X1 U21855 ( .C1(n18612), .C2(n18599), .A(n18598), .B(n18597), .ZN(
        n18936) );
  INV_X1 U21856 ( .A(n18600), .ZN(n18614) );
  AND2_X1 U21857 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18614), .ZN(
        n18617) );
  AOI21_X1 U21858 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18716), .A(
        n18617), .ZN(n18601) );
  OAI22_X1 U21859 ( .A1(n18602), .A2(n18601), .B1(n19024), .B2(n19593), .ZN(
        n18603) );
  AOI21_X1 U21860 ( .B1(n18604), .B2(n18715), .A(n18603), .ZN(n18608) );
  AOI22_X1 U21861 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18610), .B1(
        n18606), .B2(n18605), .ZN(n18607) );
  OAI211_X1 U21862 ( .C1(n18609), .C2(n18936), .A(n18608), .B(n18607), .ZN(
        P3_U2820) );
  INV_X1 U21863 ( .A(n18610), .ZN(n18620) );
  NAND2_X1 U21864 ( .A1(n18612), .A2(n18611), .ZN(n18613) );
  XNOR2_X1 U21865 ( .A(n18613), .B(n18940), .ZN(n18945) );
  NOR2_X1 U21866 ( .A1(n19024), .A2(n19591), .ZN(n18944) );
  AOI21_X1 U21867 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18716), .A(
        n18614), .ZN(n18616) );
  OAI22_X1 U21868 ( .A1(n18617), .A2(n18616), .B1(n18707), .B2(n18615), .ZN(
        n18618) );
  AOI211_X1 U21869 ( .C1(n18635), .C2(n18945), .A(n18944), .B(n18618), .ZN(
        n18619) );
  OAI221_X1 U21870 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18621), .C1(
        n18940), .C2(n18620), .A(n18619), .ZN(P3_U2821) );
  OAI21_X1 U21871 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18623), .A(
        n18622), .ZN(n18965) );
  AOI211_X1 U21872 ( .C1(n18626), .C2(n18625), .A(n18624), .B(n19335), .ZN(
        n18632) );
  OAI21_X1 U21873 ( .B1(n18628), .B2(n18627), .A(n9585), .ZN(n18641) );
  AOI22_X1 U21874 ( .A1(n18715), .A2(n18629), .B1(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18641), .ZN(n18630) );
  INV_X1 U21875 ( .A(n18630), .ZN(n18631) );
  AOI211_X1 U21876 ( .C1(P3_REIP_REG_8__SCAN_IN), .C2(n9586), .A(n18632), .B(
        n18631), .ZN(n18638) );
  OAI21_X1 U21877 ( .B1(n18634), .B2(n18962), .A(n18633), .ZN(n18959) );
  AOI22_X1 U21878 ( .A1(n18636), .A2(n18962), .B1(n18635), .B2(n18959), .ZN(
        n18637) );
  OAI211_X1 U21879 ( .C1(n18725), .C2(n18965), .A(n18638), .B(n18637), .ZN(
        P3_U2822) );
  NOR2_X1 U21880 ( .A1(n19024), .A2(n19587), .ZN(n18972) );
  AOI221_X1 U21881 ( .B1(n18641), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n18640), .C2(n10338), .A(n18972), .ZN(n18648) );
  AOI21_X1 U21882 ( .B1(n18643), .B2(n18642), .A(n9625), .ZN(n18644) );
  XNOR2_X1 U21883 ( .A(n18644), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18968) );
  INV_X1 U21884 ( .A(n18968), .ZN(n18646) );
  AOI22_X1 U21885 ( .A1(n18713), .A2(n18646), .B1(n18645), .B2(n18715), .ZN(
        n18647) );
  OAI211_X1 U21886 ( .C1(n18724), .C2(n18974), .A(n18648), .B(n18647), .ZN(
        P3_U2823) );
  OAI21_X1 U21887 ( .B1(n18651), .B2(n18650), .A(n18649), .ZN(n18976) );
  NOR2_X1 U21888 ( .A1(n17714), .A2(n19335), .ZN(n18653) );
  AOI22_X1 U21889 ( .A1(n9586), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n18653), .B2(
        n18652), .ZN(n18660) );
  INV_X1 U21890 ( .A(n18716), .ZN(n18654) );
  NOR2_X1 U21891 ( .A1(n18654), .A2(n18653), .ZN(n18670) );
  OAI21_X1 U21892 ( .B1(n18656), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n18655), .ZN(n18981) );
  OAI22_X1 U21893 ( .A1(n18707), .A2(n18657), .B1(n18725), .B2(n18981), .ZN(
        n18658) );
  AOI21_X1 U21894 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18670), .A(
        n18658), .ZN(n18659) );
  OAI211_X1 U21895 ( .C1(n18724), .C2(n18976), .A(n18660), .B(n18659), .ZN(
        P3_U2824) );
  OAI21_X1 U21896 ( .B1(n18663), .B2(n18662), .A(n18661), .ZN(n18664) );
  XNOR2_X1 U21897 ( .A(n18664), .B(n18985), .ZN(n18988) );
  OAI21_X1 U21898 ( .B1(n18667), .B2(n18666), .A(n18665), .ZN(n18982) );
  OAI22_X1 U21899 ( .A1(n18725), .A2(n18982), .B1(n19024), .B2(n19584), .ZN(
        n18668) );
  AOI21_X1 U21900 ( .B1(n18669), .B2(n18715), .A(n18668), .ZN(n18672) );
  OAI221_X1 U21901 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17727), .C1(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n9585), .A(n18670), .ZN(n18671)
         );
  OAI211_X1 U21902 ( .C1(n18724), .C2(n18988), .A(n18672), .B(n18671), .ZN(
        P3_U2825) );
  AOI21_X1 U21903 ( .B1(n18693), .B2(n17738), .A(n18673), .ZN(n18700) );
  OAI21_X1 U21904 ( .B1(n18676), .B2(n18675), .A(n18674), .ZN(n18677) );
  XNOR2_X1 U21905 ( .A(n18677), .B(n18998), .ZN(n19001) );
  OAI22_X1 U21906 ( .A1(n18725), .A2(n19001), .B1(n19335), .B2(n18678), .ZN(
        n18684) );
  AOI21_X1 U21907 ( .B1(n18681), .B2(n18680), .A(n18679), .ZN(n18995) );
  OAI22_X1 U21908 ( .A1(n18707), .A2(n18682), .B1(n18995), .B2(n18724), .ZN(
        n18683) );
  AOI211_X1 U21909 ( .C1(n9586), .C2(P3_REIP_REG_4__SCAN_IN), .A(n18684), .B(
        n18683), .ZN(n18685) );
  OAI21_X1 U21910 ( .B1(n18700), .B2(n18686), .A(n18685), .ZN(P3_U2826) );
  OAI21_X1 U21911 ( .B1(n18689), .B2(n18688), .A(n18687), .ZN(n19004) );
  OAI22_X1 U21912 ( .A1(n18724), .A2(n19004), .B1(n19024), .B2(n19579), .ZN(
        n18696) );
  OAI21_X1 U21913 ( .B1(n18692), .B2(n18691), .A(n18690), .ZN(n19005) );
  NAND2_X1 U21914 ( .A1(n18693), .A2(n17738), .ZN(n18694) );
  NAND2_X1 U21915 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n9585), .ZN(
        n18709) );
  OAI22_X1 U21916 ( .A1(n18725), .A2(n19005), .B1(n18694), .B2(n18709), .ZN(
        n18695) );
  AOI211_X1 U21917 ( .C1(n18697), .C2(n18715), .A(n18696), .B(n18695), .ZN(
        n18698) );
  OAI21_X1 U21918 ( .B1(n18700), .B2(n18699), .A(n18698), .ZN(P3_U2827) );
  OAI21_X1 U21919 ( .B1(n18705), .B2(n18704), .A(n18703), .ZN(n19019) );
  OAI22_X1 U21920 ( .A1(n18707), .A2(n18706), .B1(n18725), .B2(n19019), .ZN(
        n18708) );
  AOI221_X1 U21921 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18709), .C1(
        n19427), .C2(n18709), .A(n18708), .ZN(n18710) );
  NAND2_X1 U21922 ( .A1(n9586), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n19021) );
  OAI211_X1 U21923 ( .C1(n18724), .C2(n19023), .A(n18710), .B(n19021), .ZN(
        P3_U2828) );
  NAND2_X1 U21924 ( .A1(n19674), .A2(n13297), .ZN(n18712) );
  XNOR2_X1 U21925 ( .A(n18712), .B(n18711), .ZN(n19030) );
  AOI22_X1 U21926 ( .A1(n18713), .A2(n19030), .B1(n9586), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18718) );
  AOI22_X1 U21927 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18716), .B1(
        n18715), .B2(n18714), .ZN(n18717) );
  OAI211_X1 U21928 ( .C1(n18724), .C2(n19036), .A(n18718), .B(n18717), .ZN(
        P3_U2829) );
  AOI21_X1 U21929 ( .B1(n13297), .B2(n19674), .A(n18719), .ZN(n19041) );
  INV_X1 U21930 ( .A(n19041), .ZN(n19039) );
  NAND3_X1 U21931 ( .A1(n19656), .A2(n9585), .A3(n18720), .ZN(n18722) );
  AOI22_X1 U21932 ( .A1(n9586), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18722), .ZN(n18723) );
  OAI221_X1 U21933 ( .B1(n19041), .B2(n18725), .C1(n19039), .C2(n18724), .A(
        n18723), .ZN(P3_U2830) );
  AOI22_X1 U21934 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n10157), .B1(
        n9586), .B2(P3_REIP_REG_27__SCAN_IN), .ZN(n18738) );
  NOR2_X1 U21935 ( .A1(n19026), .A2(n18734), .ZN(n18735) );
  INV_X1 U21936 ( .A(n18726), .ZN(n18740) );
  NOR2_X1 U21937 ( .A1(n19494), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18989) );
  NOR2_X1 U21938 ( .A1(n18989), .A2(n18727), .ZN(n18827) );
  NOR2_X1 U21939 ( .A1(n19032), .A2(n19499), .ZN(n18990) );
  AOI21_X1 U21940 ( .B1(n18740), .B2(n18827), .A(n18990), .ZN(n18765) );
  INV_X1 U21941 ( .A(n18728), .ZN(n18766) );
  AOI211_X1 U21942 ( .C1(n18851), .C2(n18729), .A(n18765), .B(n18766), .ZN(
        n18750) );
  AOI22_X1 U21943 ( .A1(n18893), .A2(n18731), .B1(n18851), .B2(n18730), .ZN(
        n18732) );
  OAI211_X1 U21944 ( .C1(n18733), .C2(n18910), .A(n18750), .B(n18732), .ZN(
        n18742) );
  OAI22_X1 U21945 ( .A1(n18736), .A2(n18735), .B1(n18742), .B2(n18734), .ZN(
        n18737) );
  OAI211_X1 U21946 ( .C1(n18739), .C2(n18935), .A(n18738), .B(n18737), .ZN(
        P3_U2835) );
  AND2_X1 U21947 ( .A1(n18791), .A2(n18740), .ZN(n18776) );
  AOI22_X1 U21948 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18742), .B1(
        n18741), .B2(n18776), .ZN(n18747) );
  INV_X1 U21949 ( .A(n18743), .ZN(n18744) );
  AOI22_X1 U21950 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n10157), .B1(
        n18960), .B2(n18744), .ZN(n18746) );
  NAND2_X1 U21951 ( .A1(n9586), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18745) );
  OAI211_X1 U21952 ( .C1(n18747), .C2(n19026), .A(n18746), .B(n18745), .ZN(
        P3_U2836) );
  NOR2_X1 U21953 ( .A1(n18749), .A2(n18748), .ZN(n18752) );
  INV_X1 U21954 ( .A(n18750), .ZN(n18751) );
  MUX2_X1 U21955 ( .A(n18752), .B(n18751), .S(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(n18753) );
  AOI22_X1 U21956 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n10157), .B1(
        n19037), .B2(n18753), .ZN(n18755) );
  OAI211_X1 U21957 ( .C1(n18756), .C2(n18935), .A(n18755), .B(n18754), .ZN(
        n18757) );
  AOI21_X1 U21958 ( .B1(n18961), .B2(n18758), .A(n18757), .ZN(n18759) );
  OAI21_X1 U21959 ( .B1(n19006), .B2(n18760), .A(n18759), .ZN(P3_U2837) );
  INV_X1 U21960 ( .A(n18761), .ZN(n18798) );
  OAI22_X1 U21961 ( .A1(n18763), .A2(n18910), .B1(n18762), .B2(n19527), .ZN(
        n18764) );
  NOR3_X1 U21962 ( .A1(n10157), .A2(n18765), .A3(n18764), .ZN(n18769) );
  NOR2_X1 U21963 ( .A1(n18767), .A2(n18766), .ZN(n18768) );
  AOI21_X1 U21964 ( .B1(n18769), .B2(n18768), .A(n9586), .ZN(n18775) );
  AOI21_X1 U21965 ( .B1(n18954), .B2(n18769), .A(n10226), .ZN(n18770) );
  AOI22_X1 U21966 ( .A1(n18798), .A2(n18771), .B1(n18775), .B2(n18770), .ZN(
        n18773) );
  NAND2_X1 U21967 ( .A1(n9586), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18772) );
  OAI211_X1 U21968 ( .C1(n18774), .C2(n18935), .A(n18773), .B(n18772), .ZN(
        P3_U2838) );
  OAI221_X1 U21969 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18776), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n19027), .A(n18775), .ZN(
        n18777) );
  OAI211_X1 U21970 ( .C1(n18779), .C2(n18935), .A(n18778), .B(n18777), .ZN(
        P3_U2839) );
  NOR2_X1 U21971 ( .A1(n19512), .A2(n19499), .ZN(n19025) );
  NAND2_X1 U21972 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18888), .ZN(
        n18937) );
  NOR2_X1 U21973 ( .A1(n18780), .A2(n18937), .ZN(n18850) );
  AOI21_X1 U21974 ( .B1(n18799), .B2(n18850), .A(n19494), .ZN(n18781) );
  AOI211_X1 U21975 ( .C1(n19512), .C2(n18782), .A(n18828), .B(n18781), .ZN(
        n18783) );
  OAI221_X1 U21976 ( .B1(n19501), .B2(n18784), .C1(n19501), .C2(n18811), .A(
        n18783), .ZN(n18812) );
  NAND2_X1 U21977 ( .A1(n19527), .A2(n18910), .ZN(n18813) );
  INV_X1 U21978 ( .A(n18813), .ZN(n18915) );
  OAI22_X1 U21979 ( .A1(n19501), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n18792), .B2(n18915), .ZN(n18785) );
  NOR2_X1 U21980 ( .A1(n18812), .A2(n18785), .ZN(n18802) );
  INV_X1 U21981 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18787) );
  AOI211_X1 U21982 ( .C1(n19032), .C2(n18800), .A(n18787), .B(n18801), .ZN(
        n18788) );
  OAI211_X1 U21983 ( .C1(n18789), .C2(n19025), .A(n18802), .B(n18788), .ZN(
        n18790) );
  OAI221_X1 U21984 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18792), 
        .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n18791), .A(n18790), .ZN(
        n18797) );
  AOI22_X1 U21985 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n10157), .B1(
        n18960), .B2(n18793), .ZN(n18796) );
  INV_X1 U21986 ( .A(n18794), .ZN(n18795) );
  OAI211_X1 U21987 ( .C1(n19026), .C2(n18797), .A(n18796), .B(n18795), .ZN(
        P3_U2840) );
  NAND2_X1 U21988 ( .A1(n18799), .A2(n18798), .ZN(n18824) );
  NOR2_X1 U21989 ( .A1(n9586), .A2(n18800), .ZN(n18805) );
  OAI211_X1 U21990 ( .C1(n18803), .C2(n19025), .A(n18831), .B(n18802), .ZN(
        n18804) );
  AOI22_X1 U21991 ( .A1(n18960), .A2(n18806), .B1(n18805), .B2(n18804), .ZN(
        n18808) );
  OAI211_X1 U21992 ( .C1(n18809), .C2(n18824), .A(n18808), .B(n18807), .ZN(
        P3_U2841) );
  AOI22_X1 U21993 ( .A1(n9586), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18960), 
        .B2(n18810), .ZN(n18818) );
  INV_X1 U21994 ( .A(n18811), .ZN(n18814) );
  AOI21_X1 U21995 ( .B1(n18814), .B2(n18813), .A(n18812), .ZN(n18815) );
  AOI21_X1 U21996 ( .B1(n18831), .B2(n18815), .A(n9586), .ZN(n18821) );
  NOR3_X1 U21997 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n19025), .A3(
        n19692), .ZN(n18816) );
  OAI21_X1 U21998 ( .B1(n18821), .B2(n18816), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18817) );
  OAI211_X1 U21999 ( .C1(n18819), .C2(n18824), .A(n18818), .B(n18817), .ZN(
        P3_U2842) );
  AOI22_X1 U22000 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18821), .B1(
        n18960), .B2(n18820), .ZN(n18823) );
  OAI211_X1 U22001 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18824), .A(
        n18823), .B(n18822), .ZN(P3_U2843) );
  INV_X1 U22002 ( .A(n19006), .ZN(n19040) );
  INV_X1 U22003 ( .A(n18993), .ZN(n19012) );
  NOR2_X1 U22004 ( .A1(n21354), .A2(n13072), .ZN(n18992) );
  AOI22_X1 U22005 ( .A1(n19512), .A2(n19012), .B1(n18992), .B2(n19016), .ZN(
        n19003) );
  NOR3_X1 U22006 ( .A1(n19003), .A2(n19026), .A3(n19011), .ZN(n18999) );
  NAND3_X1 U22007 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n18999), .ZN(n18977) );
  INV_X1 U22008 ( .A(n18977), .ZN(n18825) );
  AOI222_X1 U22009 ( .A1(n18961), .A2(n18911), .B1(n19040), .B2(n18909), .C1(
        n18826), .C2(n18825), .ZN(n18947) );
  INV_X1 U22010 ( .A(n18947), .ZN(n18926) );
  NAND2_X1 U22011 ( .A1(n9603), .A2(n18926), .ZN(n18857) );
  AOI21_X1 U22012 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18827), .A(
        n18990), .ZN(n18833) );
  INV_X1 U22013 ( .A(n18828), .ZN(n18829) );
  AOI22_X1 U22014 ( .A1(n18830), .A2(n18829), .B1(n18915), .B2(n19528), .ZN(
        n18832) );
  AOI221_X1 U22015 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18840), 
        .C1(n18990), .C2(n18840), .A(n9586), .ZN(n18835) );
  AOI22_X1 U22016 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18835), .B1(
        n18960), .B2(n18834), .ZN(n18837) );
  OAI211_X1 U22017 ( .C1(n18857), .C2(n18838), .A(n18837), .B(n18836), .ZN(
        P3_U2844) );
  NOR2_X1 U22018 ( .A1(n19024), .A2(n19607), .ZN(n18842) );
  NOR3_X1 U22019 ( .A1(n9586), .A2(n18840), .A3(n18839), .ZN(n18841) );
  AOI211_X1 U22020 ( .C1(n18960), .C2(n18843), .A(n18842), .B(n18841), .ZN(
        n18844) );
  OAI21_X1 U22021 ( .B1(n18857), .B2(n18845), .A(n18844), .ZN(P3_U2845) );
  NOR2_X1 U22022 ( .A1(n19501), .A2(n18888), .ZN(n18928) );
  INV_X1 U22023 ( .A(n18846), .ZN(n18872) );
  NOR2_X1 U22024 ( .A1(n18872), .A2(n19528), .ZN(n18913) );
  AOI211_X1 U22025 ( .C1(n18848), .C2(n18847), .A(n18928), .B(n18913), .ZN(
        n18849) );
  OAI211_X1 U22026 ( .C1(n18850), .C2(n19494), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18849), .ZN(n18863) );
  OAI221_X1 U22027 ( .B1(n18852), .B2(n18851), .C1(n18852), .C2(n18863), .A(
        n19024), .ZN(n18855) );
  AOI22_X1 U22028 ( .A1(n9586), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18960), 
        .B2(n18853), .ZN(n18854) );
  OAI221_X1 U22029 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18857), 
        .C1(n18856), .C2(n18855), .A(n18854), .ZN(P3_U2846) );
  NAND2_X1 U22030 ( .A1(n18859), .A2(n18858), .ZN(n18871) );
  AOI22_X1 U22031 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n10157), .B1(
        n9586), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n18870) );
  OR2_X1 U22032 ( .A1(n18910), .A2(n18860), .ZN(n18865) );
  NOR4_X1 U22033 ( .A1(n19003), .A2(n18966), .A3(n18862), .A4(n18861), .ZN(
        n18879) );
  OAI221_X1 U22034 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18879), .A(n18863), .ZN(
        n18864) );
  OAI21_X1 U22035 ( .B1(n18866), .B2(n18865), .A(n18864), .ZN(n18868) );
  AOI22_X1 U22036 ( .A1(n19037), .A2(n18868), .B1(n18960), .B2(n18867), .ZN(
        n18869) );
  OAI211_X1 U22037 ( .C1(n19006), .C2(n18871), .A(n18870), .B(n18869), .ZN(
        P3_U2847) );
  AOI21_X1 U22038 ( .B1(n18873), .B2(n18872), .A(n19528), .ZN(n18877) );
  OAI22_X1 U22039 ( .A1(n19501), .A2(n18874), .B1(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n19025), .ZN(n18875) );
  NOR4_X1 U22040 ( .A1(n18877), .A2(n18928), .A3(n18876), .A4(n18875), .ZN(
        n18878) );
  OAI21_X1 U22041 ( .B1(n18899), .B2(n18937), .A(n19499), .ZN(n18894) );
  AOI21_X1 U22042 ( .B1(n18878), .B2(n18894), .A(n19026), .ZN(n18880) );
  AOI222_X1 U22043 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18880), 
        .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n10157), .C1(n18880), 
        .C2(n18879), .ZN(n18886) );
  OAI22_X1 U22044 ( .A1(n18882), .A2(n18935), .B1(n19006), .B2(n18881), .ZN(
        n18883) );
  AOI21_X1 U22045 ( .B1(n18961), .B2(n18884), .A(n18883), .ZN(n18885) );
  OAI211_X1 U22046 ( .C1(n19024), .C2(n19602), .A(n18886), .B(n18885), .ZN(
        P3_U2848) );
  AOI22_X1 U22047 ( .A1(n9586), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18887), 
        .B2(n18926), .ZN(n18897) );
  AOI21_X1 U22048 ( .B1(n19032), .B2(n18918), .A(n21454), .ZN(n18901) );
  AOI21_X1 U22049 ( .B1(n18916), .B2(n18888), .A(n19501), .ZN(n18889) );
  AOI21_X1 U22050 ( .B1(n19512), .B2(n18903), .A(n18889), .ZN(n18920) );
  OAI21_X1 U22051 ( .B1(n18890), .B2(n18910), .A(n18920), .ZN(n18891) );
  AOI211_X1 U22052 ( .C1(n18893), .C2(n18892), .A(n18913), .B(n18891), .ZN(
        n18900) );
  OAI211_X1 U22053 ( .C1(n18929), .C2(n18901), .A(n18900), .B(n18894), .ZN(
        n18895) );
  OAI211_X1 U22054 ( .C1(n19026), .C2(n18895), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n19024), .ZN(n18896) );
  OAI211_X1 U22055 ( .C1(n18898), .C2(n18935), .A(n18897), .B(n18896), .ZN(
        P3_U2849) );
  NOR2_X1 U22056 ( .A1(n18899), .A2(n18937), .ZN(n18902) );
  OAI211_X1 U22057 ( .C1(n18902), .C2(n19494), .A(n18901), .B(n18900), .ZN(
        n18905) );
  OAI22_X1 U22058 ( .A1(n18947), .A2(n18903), .B1(n21454), .B2(n19026), .ZN(
        n18904) );
  AOI22_X1 U22059 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n10157), .B1(
        n18905), .B2(n18904), .ZN(n18907) );
  NAND2_X1 U22060 ( .A1(n9586), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18906) );
  OAI211_X1 U22061 ( .C1(n18908), .C2(n18935), .A(n18907), .B(n18906), .ZN(
        P3_U2850) );
  OAI22_X1 U22062 ( .A1(n18911), .A2(n18910), .B1(n19527), .B2(n18909), .ZN(
        n18912) );
  NOR3_X1 U22063 ( .A1(n18913), .A2(n19026), .A3(n18912), .ZN(n18942) );
  OAI21_X1 U22064 ( .B1(n18940), .B2(n18937), .A(n19499), .ZN(n18914) );
  OAI211_X1 U22065 ( .C1(n18916), .C2(n18915), .A(n18942), .B(n18914), .ZN(
        n18931) );
  AOI21_X1 U22066 ( .B1(n19499), .B2(n18917), .A(n18931), .ZN(n18919) );
  AOI211_X1 U22067 ( .C1(n18920), .C2(n18919), .A(n9586), .B(n18918), .ZN(
        n18921) );
  AOI211_X1 U22068 ( .C1(n18960), .C2(n18923), .A(n18922), .B(n18921), .ZN(
        n18924) );
  OAI21_X1 U22069 ( .B1(n18947), .B2(n18925), .A(n18924), .ZN(P3_U2851) );
  NOR2_X1 U22070 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18940), .ZN(
        n18927) );
  AOI22_X1 U22071 ( .A1(n9586), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18927), 
        .B2(n18926), .ZN(n18934) );
  INV_X1 U22072 ( .A(n18928), .ZN(n18930) );
  AOI21_X1 U22073 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18930), .A(
        n18929), .ZN(n18932) );
  OAI211_X1 U22074 ( .C1(n18932), .C2(n18931), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n19024), .ZN(n18933) );
  OAI211_X1 U22075 ( .C1(n18936), .C2(n18935), .A(n18934), .B(n18933), .ZN(
        P3_U2852) );
  INV_X1 U22076 ( .A(n18937), .ZN(n18938) );
  AOI211_X1 U22077 ( .C1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n19494), .A(
        n18990), .B(n18938), .ZN(n18939) );
  AOI221_X1 U22078 ( .B1(n18948), .B2(n19032), .C1(n18952), .C2(n19032), .A(
        n18939), .ZN(n18941) );
  AOI211_X1 U22079 ( .C1(n18942), .C2(n18941), .A(n9586), .B(n18940), .ZN(
        n18943) );
  AOI211_X1 U22080 ( .C1(n18960), .C2(n18945), .A(n18944), .B(n18943), .ZN(
        n18946) );
  OAI21_X1 U22081 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18947), .A(
        n18946), .ZN(P3_U2853) );
  NOR2_X1 U22082 ( .A1(n18948), .A2(n18977), .ZN(n18958) );
  INV_X1 U22083 ( .A(n18990), .ZN(n18951) );
  NOR2_X1 U22084 ( .A1(n18949), .A2(n19528), .ZN(n18950) );
  AOI211_X1 U22085 ( .C1(n18952), .C2(n18951), .A(n18950), .B(n18989), .ZN(
        n18975) );
  OAI211_X1 U22086 ( .C1(n18954), .C2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n18975), .ZN(n18953) );
  NAND2_X1 U22087 ( .A1(n19037), .A2(n18953), .ZN(n18969) );
  OAI21_X1 U22088 ( .B1(n18954), .B2(n18969), .A(n19027), .ZN(n18956) );
  INV_X1 U22089 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19589) );
  NOR2_X1 U22090 ( .A1(n19024), .A2(n19589), .ZN(n18955) );
  AOI221_X1 U22091 ( .B1(n18958), .B2(n18957), .C1(n18956), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18955), .ZN(n18964) );
  AOI22_X1 U22092 ( .A1(n18962), .A2(n18961), .B1(n18960), .B2(n18959), .ZN(
        n18963) );
  OAI211_X1 U22093 ( .C1(n19006), .C2(n18965), .A(n18964), .B(n18963), .ZN(
        P3_U2854) );
  NOR2_X1 U22094 ( .A1(n19003), .A2(n18966), .ZN(n18967) );
  AOI21_X1 U22095 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18967), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18970) );
  OAI22_X1 U22096 ( .A1(n18970), .A2(n18969), .B1(n19006), .B2(n18968), .ZN(
        n18971) );
  AOI211_X1 U22097 ( .C1(n10157), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18972), .B(n18971), .ZN(n18973) );
  OAI21_X1 U22098 ( .B1(n19035), .B2(n18974), .A(n18973), .ZN(P3_U2855) );
  AOI21_X1 U22099 ( .B1(n19037), .B2(n18975), .A(n9586), .ZN(n18984) );
  NOR2_X1 U22100 ( .A1(n19024), .A2(n19585), .ZN(n18979) );
  OAI22_X1 U22101 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18977), .B1(
        n18976), .B2(n19035), .ZN(n18978) );
  AOI211_X1 U22102 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n18984), .A(
        n18979), .B(n18978), .ZN(n18980) );
  OAI21_X1 U22103 ( .B1(n19006), .B2(n18981), .A(n18980), .ZN(P3_U2856) );
  OAI22_X1 U22104 ( .A1(n19024), .A2(n19584), .B1(n19006), .B2(n18982), .ZN(
        n18983) );
  AOI21_X1 U22105 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18984), .A(
        n18983), .ZN(n18987) );
  NAND3_X1 U22106 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18999), .A3(
        n18985), .ZN(n18986) );
  OAI211_X1 U22107 ( .C1(n18988), .C2(n19035), .A(n18987), .B(n18986), .ZN(
        P3_U2857) );
  INV_X1 U22108 ( .A(n18989), .ZN(n18991) );
  AOI21_X1 U22109 ( .B1(n18992), .B2(n18991), .A(n18990), .ZN(n19015) );
  AOI211_X1 U22110 ( .C1(n19512), .C2(n18993), .A(n19015), .B(n19011), .ZN(
        n19002) );
  OAI21_X1 U22111 ( .B1(n19002), .B2(n18994), .A(n19027), .ZN(n18997) );
  OAI22_X1 U22112 ( .A1(n18995), .A2(n19035), .B1(n19024), .B2(n19581), .ZN(
        n18996) );
  AOI221_X1 U22113 ( .B1(n18999), .B2(n18998), .C1(n18997), .C2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n18996), .ZN(n19000) );
  OAI21_X1 U22114 ( .B1(n19006), .B2(n19001), .A(n19000), .ZN(P3_U2858) );
  AOI211_X1 U22115 ( .C1(n19003), .C2(n19011), .A(n19002), .B(n19026), .ZN(
        n19008) );
  OAI22_X1 U22116 ( .A1(n19006), .A2(n19005), .B1(n19035), .B2(n19004), .ZN(
        n19007) );
  NOR2_X1 U22117 ( .A1(n19008), .A2(n19007), .ZN(n19010) );
  NAND2_X1 U22118 ( .A1(n9586), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n19009) );
  OAI211_X1 U22119 ( .C1(n19027), .C2(n19011), .A(n19010), .B(n19009), .ZN(
        P3_U2859) );
  NOR3_X1 U22120 ( .A1(n19528), .A2(n19674), .A3(n13072), .ZN(n19014) );
  NOR2_X1 U22121 ( .A1(n19528), .A2(n19012), .ZN(n19013) );
  AOI221_X1 U22122 ( .B1(n19015), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .C1(
        n19014), .C2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n19013), .ZN(
        n19018) );
  NAND3_X1 U22123 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19016), .A3(
        n21354), .ZN(n19017) );
  OAI211_X1 U22124 ( .C1(n19019), .C2(n19527), .A(n19018), .B(n19017), .ZN(
        n19020) );
  AOI22_X1 U22125 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10157), .B1(
        n19037), .B2(n19020), .ZN(n19022) );
  OAI211_X1 U22126 ( .C1(n19035), .C2(n19023), .A(n19022), .B(n19021), .ZN(
        P3_U2860) );
  NOR2_X1 U22127 ( .A1(n19024), .A2(n19678), .ZN(n19029) );
  OR3_X1 U22128 ( .A1(n19026), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n19025), .ZN(n19043) );
  AOI21_X1 U22129 ( .B1(n19027), .B2(n19043), .A(n13072), .ZN(n19028) );
  AOI211_X1 U22130 ( .C1(n19040), .C2(n19030), .A(n19029), .B(n19028), .ZN(
        n19034) );
  OAI211_X1 U22131 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n19032), .A(
        n19031), .B(n13072), .ZN(n19033) );
  OAI211_X1 U22132 ( .C1(n19036), .C2(n19035), .A(n19034), .B(n19033), .ZN(
        P3_U2861) );
  INV_X1 U22133 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n19684) );
  AOI211_X1 U22134 ( .C1(n19501), .C2(n19037), .A(n9586), .B(n19674), .ZN(
        n19038) );
  AOI221_X1 U22135 ( .B1(n19042), .B2(n19041), .C1(n19040), .C2(n19039), .A(
        n19038), .ZN(n19044) );
  OAI211_X1 U22136 ( .C1(n19684), .C2(n19024), .A(n19044), .B(n19043), .ZN(
        P3_U2862) );
  AOI21_X1 U22137 ( .B1(n19047), .B2(n19046), .A(n19045), .ZN(n19542) );
  INV_X1 U22138 ( .A(n19219), .ZN(n19088) );
  OAI21_X1 U22139 ( .B1(n19542), .B2(n19088), .A(n19052), .ZN(n19048) );
  OAI221_X1 U22140 ( .B1(n19195), .B2(n19699), .C1(n19195), .C2(n19052), .A(
        n19048), .ZN(P3_U2863) );
  NOR2_X1 U22141 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19514), .ZN(
        n19220) );
  NOR2_X1 U22142 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19517), .ZN(
        n19286) );
  NOR2_X1 U22143 ( .A1(n19220), .A2(n19286), .ZN(n19050) );
  OAI22_X1 U22144 ( .A1(n19051), .A2(n19517), .B1(n19050), .B2(n19049), .ZN(
        P3_U2866) );
  INV_X1 U22145 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19518) );
  NOR2_X1 U22146 ( .A1(n19518), .A2(n19052), .ZN(P3_U2867) );
  NOR2_X1 U22147 ( .A1(n19514), .A2(n19517), .ZN(n19363) );
  NOR2_X1 U22148 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19195), .ZN(
        n19264) );
  NAND2_X1 U22149 ( .A1(n19363), .A2(n19264), .ZN(n19481) );
  NAND2_X1 U22150 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19427), .ZN(n19431) );
  NOR2_X1 U22151 ( .A1(n19517), .A2(n19194), .ZN(n19425) );
  NAND2_X1 U22152 ( .A1(n19195), .A2(n19425), .ZN(n19398) );
  INV_X1 U22153 ( .A(n19398), .ZN(n19416) );
  NOR2_X2 U22154 ( .A1(n19335), .A2(n16263), .ZN(n19423) );
  NOR2_X2 U22155 ( .A1(n19334), .A2(n21451), .ZN(n19422) );
  NAND2_X1 U22156 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19425), .ZN(
        n19450) );
  INV_X1 U22157 ( .A(n19450), .ZN(n19476) );
  NAND2_X1 U22158 ( .A1(n21428), .A2(n19195), .ZN(n19505) );
  NAND2_X1 U22159 ( .A1(n19514), .A2(n19517), .ZN(n19107) );
  NOR2_X2 U22160 ( .A1(n19505), .A2(n19107), .ZN(n19140) );
  NOR2_X1 U22161 ( .A1(n19476), .A2(n19140), .ZN(n19109) );
  NOR2_X1 U22162 ( .A1(n19388), .A2(n19109), .ZN(n19082) );
  AOI22_X1 U22163 ( .A1(n19416), .A2(n19423), .B1(n19422), .B2(n19082), .ZN(
        n19058) );
  INV_X1 U22164 ( .A(n19481), .ZN(n19465) );
  NOR2_X1 U22165 ( .A1(n19465), .A2(n19416), .ZN(n19390) );
  OAI21_X1 U22166 ( .B1(n19195), .B2(n19650), .A(n19394), .ZN(n19196) );
  OAI22_X1 U22167 ( .A1(n19335), .A2(n19390), .B1(n19196), .B2(n19109), .ZN(
        n19053) );
  INV_X1 U22168 ( .A(n19053), .ZN(n19085) );
  NAND2_X1 U22169 ( .A1(n19055), .A2(n19054), .ZN(n19083) );
  NOR2_X1 U22170 ( .A1(n19056), .A2(n19083), .ZN(n19428) );
  AOI22_X1 U22171 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19085), .B1(
        n19140), .B2(n19428), .ZN(n19057) );
  OAI211_X1 U22172 ( .C1(n19481), .C2(n19431), .A(n19058), .B(n19057), .ZN(
        P3_U2868) );
  NAND2_X1 U22173 ( .A1(n19427), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19437) );
  AND2_X1 U22174 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19427), .ZN(n19433) );
  AND2_X1 U22175 ( .A1(n19394), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19432) );
  AOI22_X1 U22176 ( .A1(n19465), .A2(n19433), .B1(n19082), .B2(n19432), .ZN(
        n19061) );
  NOR2_X1 U22177 ( .A1(n19059), .A2(n19083), .ZN(n19434) );
  AOI22_X1 U22178 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19085), .B1(
        n19140), .B2(n19434), .ZN(n19060) );
  OAI211_X1 U22179 ( .C1(n19398), .C2(n19437), .A(n19061), .B(n19060), .ZN(
        P3_U2869) );
  NAND2_X1 U22180 ( .A1(n19427), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19372) );
  NAND2_X1 U22181 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19427), .ZN(n19443) );
  INV_X1 U22182 ( .A(n19443), .ZN(n19369) );
  NOR2_X2 U22183 ( .A1(n19334), .A2(n21446), .ZN(n19438) );
  AOI22_X1 U22184 ( .A1(n19465), .A2(n19369), .B1(n19082), .B2(n19438), .ZN(
        n19064) );
  NOR2_X2 U22185 ( .A1(n19062), .A2(n19083), .ZN(n19440) );
  AOI22_X1 U22186 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19085), .B1(
        n19140), .B2(n19440), .ZN(n19063) );
  OAI211_X1 U22187 ( .C1(n19398), .C2(n19372), .A(n19064), .B(n19063), .ZN(
        P3_U2870) );
  NAND2_X1 U22188 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19427), .ZN(n19406) );
  AND2_X1 U22189 ( .A1(n19427), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19446) );
  NOR2_X2 U22190 ( .A1(n19334), .A2(n19065), .ZN(n19444) );
  AOI22_X1 U22191 ( .A1(n19416), .A2(n19446), .B1(n19082), .B2(n19444), .ZN(
        n19068) );
  NOR2_X1 U22192 ( .A1(n19066), .A2(n19083), .ZN(n19403) );
  AOI22_X1 U22193 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19085), .B1(
        n19140), .B2(n19403), .ZN(n19067) );
  OAI211_X1 U22194 ( .C1(n19481), .C2(n19406), .A(n19068), .B(n19067), .ZN(
        P3_U2871) );
  NAND2_X1 U22195 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19427), .ZN(n19378) );
  NAND2_X1 U22196 ( .A1(n19427), .A2(BUF2_REG_20__SCAN_IN), .ZN(n19456) );
  INV_X1 U22197 ( .A(n19456), .ZN(n19375) );
  NOR2_X2 U22198 ( .A1(n19334), .A2(n19069), .ZN(n19451) );
  AOI22_X1 U22199 ( .A1(n19416), .A2(n19375), .B1(n19082), .B2(n19451), .ZN(
        n19072) );
  NOR2_X2 U22200 ( .A1(n19070), .A2(n19083), .ZN(n19453) );
  AOI22_X1 U22201 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19085), .B1(
        n19140), .B2(n19453), .ZN(n19071) );
  OAI211_X1 U22202 ( .C1(n19481), .C2(n19378), .A(n19072), .B(n19071), .ZN(
        P3_U2872) );
  NAND2_X1 U22203 ( .A1(n19427), .A2(BUF2_REG_21__SCAN_IN), .ZN(n19462) );
  AND2_X1 U22204 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19427), .ZN(n19458) );
  NOR2_X2 U22205 ( .A1(n19334), .A2(n19073), .ZN(n19457) );
  AOI22_X1 U22206 ( .A1(n19465), .A2(n19458), .B1(n19082), .B2(n19457), .ZN(
        n19076) );
  NOR2_X2 U22207 ( .A1(n19074), .A2(n19083), .ZN(n19459) );
  AOI22_X1 U22208 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19085), .B1(
        n19140), .B2(n19459), .ZN(n19075) );
  OAI211_X1 U22209 ( .C1(n19398), .C2(n19462), .A(n19076), .B(n19075), .ZN(
        P3_U2873) );
  NAND2_X1 U22210 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19427), .ZN(n19470) );
  NOR2_X1 U22211 ( .A1(n19335), .A2(n16214), .ZN(n19464) );
  NOR2_X2 U22212 ( .A1(n19334), .A2(n19077), .ZN(n19463) );
  AOI22_X1 U22213 ( .A1(n19416), .A2(n19464), .B1(n19082), .B2(n19463), .ZN(
        n19080) );
  NOR2_X2 U22214 ( .A1(n19078), .A2(n19083), .ZN(n19466) );
  AOI22_X1 U22215 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19085), .B1(
        n19140), .B2(n19466), .ZN(n19079) );
  OAI211_X1 U22216 ( .C1(n19481), .C2(n19470), .A(n19080), .B(n19079), .ZN(
        P3_U2874) );
  NAND2_X1 U22217 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19427), .ZN(n19480) );
  NAND2_X1 U22218 ( .A1(n19427), .A2(BUF2_REG_31__SCAN_IN), .ZN(n19421) );
  INV_X1 U22219 ( .A(n19421), .ZN(n19474) );
  NOR2_X2 U22220 ( .A1(n19081), .A2(n19334), .ZN(n19472) );
  AOI22_X1 U22221 ( .A1(n19465), .A2(n19474), .B1(n19082), .B2(n19472), .ZN(
        n19087) );
  NOR2_X2 U22222 ( .A1(n19084), .A2(n19083), .ZN(n19475) );
  AOI22_X1 U22223 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19085), .B1(
        n19140), .B2(n19475), .ZN(n19086) );
  OAI211_X1 U22224 ( .C1(n19398), .C2(n19480), .A(n19087), .B(n19086), .ZN(
        P3_U2875) );
  INV_X1 U22225 ( .A(n19107), .ZN(n19129) );
  NAND2_X1 U22226 ( .A1(n19129), .A2(n19264), .ZN(n19166) );
  INV_X1 U22227 ( .A(n19431), .ZN(n19389) );
  INV_X1 U22228 ( .A(n19388), .ZN(n19550) );
  NAND2_X1 U22229 ( .A1(n21428), .A2(n19550), .ZN(n19360) );
  NOR2_X1 U22230 ( .A1(n19107), .A2(n19360), .ZN(n19103) );
  AOI22_X1 U22231 ( .A1(n19416), .A2(n19389), .B1(n19422), .B2(n19103), .ZN(
        n19090) );
  NOR2_X1 U22232 ( .A1(n19334), .A2(n19088), .ZN(n19424) );
  AND2_X1 U22233 ( .A1(n21428), .A2(n19424), .ZN(n19362) );
  AOI22_X1 U22234 ( .A1(n19427), .A2(n19425), .B1(n19129), .B2(n19362), .ZN(
        n19104) );
  AOI22_X1 U22235 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19104), .B1(
        n19476), .B2(n19423), .ZN(n19089) );
  OAI211_X1 U22236 ( .C1(n19397), .C2(n19166), .A(n19090), .B(n19089), .ZN(
        P3_U2876) );
  INV_X1 U22237 ( .A(n19437), .ZN(n19340) );
  AOI22_X1 U22238 ( .A1(n19476), .A2(n19340), .B1(n19432), .B2(n19103), .ZN(
        n19092) );
  AOI22_X1 U22239 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19104), .B1(
        n19416), .B2(n19433), .ZN(n19091) );
  OAI211_X1 U22240 ( .C1(n19343), .C2(n19166), .A(n19092), .B(n19091), .ZN(
        P3_U2877) );
  AOI22_X1 U22241 ( .A1(n19416), .A2(n19369), .B1(n19438), .B2(n19103), .ZN(
        n19094) );
  INV_X1 U22242 ( .A(n19166), .ZN(n19168) );
  AOI22_X1 U22243 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19104), .B1(
        n19440), .B2(n19168), .ZN(n19093) );
  OAI211_X1 U22244 ( .C1(n19450), .C2(n19372), .A(n19094), .B(n19093), .ZN(
        P3_U2878) );
  AOI22_X1 U22245 ( .A1(n19476), .A2(n19446), .B1(n19444), .B2(n19103), .ZN(
        n19096) );
  AOI22_X1 U22246 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19104), .B1(
        n19403), .B2(n19168), .ZN(n19095) );
  OAI211_X1 U22247 ( .C1(n19398), .C2(n19406), .A(n19096), .B(n19095), .ZN(
        P3_U2879) );
  INV_X1 U22248 ( .A(n19378), .ZN(n19452) );
  AOI22_X1 U22249 ( .A1(n19416), .A2(n19452), .B1(n19451), .B2(n19103), .ZN(
        n19098) );
  AOI22_X1 U22250 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19104), .B1(
        n19453), .B2(n19168), .ZN(n19097) );
  OAI211_X1 U22251 ( .C1(n19450), .C2(n19456), .A(n19098), .B(n19097), .ZN(
        P3_U2880) );
  AOI22_X1 U22252 ( .A1(n19416), .A2(n19458), .B1(n19457), .B2(n19103), .ZN(
        n19100) );
  AOI22_X1 U22253 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19104), .B1(
        n19459), .B2(n19168), .ZN(n19099) );
  OAI211_X1 U22254 ( .C1(n19450), .C2(n19462), .A(n19100), .B(n19099), .ZN(
        P3_U2881) );
  AOI22_X1 U22255 ( .A1(n19476), .A2(n19464), .B1(n19463), .B2(n19103), .ZN(
        n19102) );
  AOI22_X1 U22256 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19104), .B1(
        n19466), .B2(n19168), .ZN(n19101) );
  OAI211_X1 U22257 ( .C1(n19398), .C2(n19470), .A(n19102), .B(n19101), .ZN(
        P3_U2882) );
  AOI22_X1 U22258 ( .A1(n19416), .A2(n19474), .B1(n19472), .B2(n19103), .ZN(
        n19106) );
  AOI22_X1 U22259 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19104), .B1(
        n19475), .B2(n19168), .ZN(n19105) );
  OAI211_X1 U22260 ( .C1(n19450), .C2(n19480), .A(n19106), .B(n19105), .ZN(
        P3_U2883) );
  NOR2_X1 U22261 ( .A1(n21428), .A2(n19107), .ZN(n19173) );
  NAND2_X1 U22262 ( .A1(n19173), .A2(n19195), .ZN(n19193) );
  NOR2_X1 U22263 ( .A1(n19168), .A2(n19186), .ZN(n19150) );
  NOR2_X1 U22264 ( .A1(n19388), .A2(n19150), .ZN(n19125) );
  AOI22_X1 U22265 ( .A1(n19476), .A2(n19389), .B1(n19422), .B2(n19125), .ZN(
        n19112) );
  INV_X1 U22266 ( .A(n19108), .ZN(n19391) );
  OAI21_X1 U22267 ( .B1(n19109), .B2(n19391), .A(n19150), .ZN(n19110) );
  OAI211_X1 U22268 ( .C1(n19186), .C2(n19650), .A(n19394), .B(n19110), .ZN(
        n19126) );
  AOI22_X1 U22269 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19126), .B1(
        n19140), .B2(n19423), .ZN(n19111) );
  OAI211_X1 U22270 ( .C1(n19397), .C2(n19193), .A(n19112), .B(n19111), .ZN(
        P3_U2884) );
  AOI22_X1 U22271 ( .A1(n19140), .A2(n19340), .B1(n19432), .B2(n19125), .ZN(
        n19114) );
  AOI22_X1 U22272 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19126), .B1(
        n19476), .B2(n19433), .ZN(n19113) );
  OAI211_X1 U22273 ( .C1(n19343), .C2(n19193), .A(n19114), .B(n19113), .ZN(
        P3_U2885) );
  INV_X1 U22274 ( .A(n19372), .ZN(n19439) );
  AOI22_X1 U22275 ( .A1(n19140), .A2(n19439), .B1(n19438), .B2(n19125), .ZN(
        n19116) );
  AOI22_X1 U22276 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19126), .B1(
        n19440), .B2(n19186), .ZN(n19115) );
  OAI211_X1 U22277 ( .C1(n19450), .C2(n19443), .A(n19116), .B(n19115), .ZN(
        P3_U2886) );
  INV_X1 U22278 ( .A(n19403), .ZN(n19449) );
  INV_X1 U22279 ( .A(n19406), .ZN(n19445) );
  AOI22_X1 U22280 ( .A1(n19476), .A2(n19445), .B1(n19444), .B2(n19125), .ZN(
        n19118) );
  AOI22_X1 U22281 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19126), .B1(
        n19140), .B2(n19446), .ZN(n19117) );
  OAI211_X1 U22282 ( .C1(n19449), .C2(n19193), .A(n19118), .B(n19117), .ZN(
        P3_U2887) );
  INV_X1 U22283 ( .A(n19140), .ZN(n19149) );
  AOI22_X1 U22284 ( .A1(n19476), .A2(n19452), .B1(n19451), .B2(n19125), .ZN(
        n19120) );
  AOI22_X1 U22285 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19126), .B1(
        n19453), .B2(n19186), .ZN(n19119) );
  OAI211_X1 U22286 ( .C1(n19149), .C2(n19456), .A(n19120), .B(n19119), .ZN(
        P3_U2888) );
  AOI22_X1 U22287 ( .A1(n19476), .A2(n19458), .B1(n19457), .B2(n19125), .ZN(
        n19122) );
  AOI22_X1 U22288 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19126), .B1(
        n19459), .B2(n19186), .ZN(n19121) );
  OAI211_X1 U22289 ( .C1(n19149), .C2(n19462), .A(n19122), .B(n19121), .ZN(
        P3_U2889) );
  INV_X1 U22290 ( .A(n19464), .ZN(n19327) );
  INV_X1 U22291 ( .A(n19470), .ZN(n19324) );
  AOI22_X1 U22292 ( .A1(n19476), .A2(n19324), .B1(n19463), .B2(n19125), .ZN(
        n19124) );
  AOI22_X1 U22293 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19126), .B1(
        n19466), .B2(n19186), .ZN(n19123) );
  OAI211_X1 U22294 ( .C1(n19149), .C2(n19327), .A(n19124), .B(n19123), .ZN(
        P3_U2890) );
  INV_X1 U22295 ( .A(n19480), .ZN(n19415) );
  AOI22_X1 U22296 ( .A1(n19140), .A2(n19415), .B1(n19472), .B2(n19125), .ZN(
        n19128) );
  AOI22_X1 U22297 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19126), .B1(
        n19475), .B2(n19186), .ZN(n19127) );
  OAI211_X1 U22298 ( .C1(n19450), .C2(n19421), .A(n19128), .B(n19127), .ZN(
        P3_U2891) );
  NAND2_X1 U22299 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19173), .ZN(
        n19213) );
  AND2_X1 U22300 ( .A1(n19550), .A2(n19173), .ZN(n19145) );
  AOI22_X1 U22301 ( .A1(n19140), .A2(n19389), .B1(n19422), .B2(n19145), .ZN(
        n19131) );
  AOI21_X1 U22302 ( .B1(n21428), .B2(n19391), .A(n19334), .ZN(n19221) );
  OAI211_X1 U22303 ( .C1(n19215), .C2(n19650), .A(n19129), .B(n19221), .ZN(
        n19146) );
  AOI22_X1 U22304 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19146), .B1(
        n19423), .B2(n19168), .ZN(n19130) );
  OAI211_X1 U22305 ( .C1(n19397), .C2(n19213), .A(n19131), .B(n19130), .ZN(
        P3_U2892) );
  AOI22_X1 U22306 ( .A1(n19340), .A2(n19168), .B1(n19432), .B2(n19145), .ZN(
        n19133) );
  AOI22_X1 U22307 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19146), .B1(
        n19140), .B2(n19433), .ZN(n19132) );
  OAI211_X1 U22308 ( .C1(n19343), .C2(n19213), .A(n19133), .B(n19132), .ZN(
        P3_U2893) );
  AOI22_X1 U22309 ( .A1(n19140), .A2(n19369), .B1(n19438), .B2(n19145), .ZN(
        n19135) );
  AOI22_X1 U22310 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19146), .B1(
        n19440), .B2(n19215), .ZN(n19134) );
  OAI211_X1 U22311 ( .C1(n19372), .C2(n19166), .A(n19135), .B(n19134), .ZN(
        P3_U2894) );
  AOI22_X1 U22312 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19146), .B1(
        n19444), .B2(n19145), .ZN(n19137) );
  AOI22_X1 U22313 ( .A1(n19403), .A2(n19215), .B1(n19446), .B2(n19168), .ZN(
        n19136) );
  OAI211_X1 U22314 ( .C1(n19149), .C2(n19406), .A(n19137), .B(n19136), .ZN(
        P3_U2895) );
  AOI22_X1 U22315 ( .A1(n19375), .A2(n19168), .B1(n19451), .B2(n19145), .ZN(
        n19139) );
  AOI22_X1 U22316 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19146), .B1(
        n19453), .B2(n19215), .ZN(n19138) );
  OAI211_X1 U22317 ( .C1(n19149), .C2(n19378), .A(n19139), .B(n19138), .ZN(
        P3_U2896) );
  AOI22_X1 U22318 ( .A1(n19140), .A2(n19458), .B1(n19457), .B2(n19145), .ZN(
        n19142) );
  AOI22_X1 U22319 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19146), .B1(
        n19459), .B2(n19215), .ZN(n19141) );
  OAI211_X1 U22320 ( .C1(n19462), .C2(n19166), .A(n19142), .B(n19141), .ZN(
        P3_U2897) );
  AOI22_X1 U22321 ( .A1(n19463), .A2(n19145), .B1(n19464), .B2(n19168), .ZN(
        n19144) );
  AOI22_X1 U22322 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19146), .B1(
        n19466), .B2(n19215), .ZN(n19143) );
  OAI211_X1 U22323 ( .C1(n19149), .C2(n19470), .A(n19144), .B(n19143), .ZN(
        P3_U2898) );
  AOI22_X1 U22324 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19146), .B1(
        n19472), .B2(n19145), .ZN(n19148) );
  AOI22_X1 U22325 ( .A1(n19415), .A2(n19168), .B1(n19475), .B2(n19215), .ZN(
        n19147) );
  OAI211_X1 U22326 ( .C1(n19149), .C2(n19421), .A(n19148), .B(n19147), .ZN(
        P3_U2899) );
  INV_X1 U22327 ( .A(n19505), .ZN(n19333) );
  NAND2_X1 U22328 ( .A1(n19333), .A2(n19220), .ZN(n19241) );
  INV_X1 U22329 ( .A(n19241), .ZN(n19234) );
  NOR2_X1 U22330 ( .A1(n19215), .A2(n19234), .ZN(n19197) );
  NOR2_X1 U22331 ( .A1(n19388), .A2(n19197), .ZN(n19167) );
  AOI22_X1 U22332 ( .A1(n19389), .A2(n19168), .B1(n19422), .B2(n19167), .ZN(
        n19153) );
  OAI22_X1 U22333 ( .A1(n19150), .A2(n19335), .B1(n19197), .B2(n19334), .ZN(
        n19151) );
  OAI21_X1 U22334 ( .B1(n19234), .B2(n19650), .A(n19151), .ZN(n19169) );
  AOI22_X1 U22335 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19169), .B1(
        n19423), .B2(n19186), .ZN(n19152) );
  OAI211_X1 U22336 ( .C1(n19397), .C2(n19241), .A(n19153), .B(n19152), .ZN(
        P3_U2900) );
  AOI22_X1 U22337 ( .A1(n19433), .A2(n19168), .B1(n19432), .B2(n19167), .ZN(
        n19155) );
  AOI22_X1 U22338 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19169), .B1(
        n19434), .B2(n19234), .ZN(n19154) );
  OAI211_X1 U22339 ( .C1(n19437), .C2(n19193), .A(n19155), .B(n19154), .ZN(
        P3_U2901) );
  AOI22_X1 U22340 ( .A1(n19369), .A2(n19168), .B1(n19438), .B2(n19167), .ZN(
        n19157) );
  AOI22_X1 U22341 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19169), .B1(
        n19440), .B2(n19234), .ZN(n19156) );
  OAI211_X1 U22342 ( .C1(n19372), .C2(n19193), .A(n19157), .B(n19156), .ZN(
        P3_U2902) );
  AOI22_X1 U22343 ( .A1(n19445), .A2(n19168), .B1(n19444), .B2(n19167), .ZN(
        n19159) );
  AOI22_X1 U22344 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19169), .B1(
        n19446), .B2(n19186), .ZN(n19158) );
  OAI211_X1 U22345 ( .C1(n19449), .C2(n19241), .A(n19159), .B(n19158), .ZN(
        P3_U2903) );
  AOI22_X1 U22346 ( .A1(n19375), .A2(n19186), .B1(n19451), .B2(n19167), .ZN(
        n19161) );
  AOI22_X1 U22347 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19169), .B1(
        n19453), .B2(n19234), .ZN(n19160) );
  OAI211_X1 U22348 ( .C1(n19378), .C2(n19166), .A(n19161), .B(n19160), .ZN(
        P3_U2904) );
  AOI22_X1 U22349 ( .A1(n19458), .A2(n19168), .B1(n19457), .B2(n19167), .ZN(
        n19163) );
  AOI22_X1 U22350 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19169), .B1(
        n19459), .B2(n19234), .ZN(n19162) );
  OAI211_X1 U22351 ( .C1(n19462), .C2(n19193), .A(n19163), .B(n19162), .ZN(
        P3_U2905) );
  AOI22_X1 U22352 ( .A1(n19463), .A2(n19167), .B1(n19464), .B2(n19186), .ZN(
        n19165) );
  AOI22_X1 U22353 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19169), .B1(
        n19466), .B2(n19234), .ZN(n19164) );
  OAI211_X1 U22354 ( .C1(n19470), .C2(n19166), .A(n19165), .B(n19164), .ZN(
        P3_U2906) );
  AOI22_X1 U22355 ( .A1(n19474), .A2(n19168), .B1(n19472), .B2(n19167), .ZN(
        n19171) );
  AOI22_X1 U22356 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19169), .B1(
        n19475), .B2(n19234), .ZN(n19170) );
  OAI211_X1 U22357 ( .C1(n19480), .C2(n19193), .A(n19171), .B(n19170), .ZN(
        P3_U2907) );
  NAND2_X1 U22358 ( .A1(n19264), .A2(n19220), .ZN(n19258) );
  INV_X1 U22359 ( .A(n19220), .ZN(n19172) );
  NOR2_X1 U22360 ( .A1(n19360), .A2(n19172), .ZN(n19189) );
  AOI22_X1 U22361 ( .A1(n19389), .A2(n19186), .B1(n19422), .B2(n19189), .ZN(
        n19175) );
  AOI22_X1 U22362 ( .A1(n19427), .A2(n19173), .B1(n19362), .B2(n19220), .ZN(
        n19190) );
  AOI22_X1 U22363 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19190), .B1(
        n19423), .B2(n19215), .ZN(n19174) );
  OAI211_X1 U22364 ( .C1(n19397), .C2(n19258), .A(n19175), .B(n19174), .ZN(
        P3_U2908) );
  AOI22_X1 U22365 ( .A1(n19340), .A2(n19215), .B1(n19432), .B2(n19189), .ZN(
        n19177) );
  AOI22_X1 U22366 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19190), .B1(
        n19433), .B2(n19186), .ZN(n19176) );
  OAI211_X1 U22367 ( .C1(n19343), .C2(n19258), .A(n19177), .B(n19176), .ZN(
        P3_U2909) );
  AOI22_X1 U22368 ( .A1(n19369), .A2(n19186), .B1(n19438), .B2(n19189), .ZN(
        n19179) );
  AOI22_X1 U22369 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19190), .B1(
        n19440), .B2(n19260), .ZN(n19178) );
  OAI211_X1 U22370 ( .C1(n19372), .C2(n19213), .A(n19179), .B(n19178), .ZN(
        P3_U2910) );
  AOI22_X1 U22371 ( .A1(n19446), .A2(n19215), .B1(n19444), .B2(n19189), .ZN(
        n19181) );
  AOI22_X1 U22372 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19190), .B1(
        n19403), .B2(n19260), .ZN(n19180) );
  OAI211_X1 U22373 ( .C1(n19406), .C2(n19193), .A(n19181), .B(n19180), .ZN(
        P3_U2911) );
  AOI22_X1 U22374 ( .A1(n19375), .A2(n19215), .B1(n19451), .B2(n19189), .ZN(
        n19183) );
  AOI22_X1 U22375 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19190), .B1(
        n19453), .B2(n19260), .ZN(n19182) );
  OAI211_X1 U22376 ( .C1(n19378), .C2(n19193), .A(n19183), .B(n19182), .ZN(
        P3_U2912) );
  AOI22_X1 U22377 ( .A1(n19458), .A2(n19186), .B1(n19457), .B2(n19189), .ZN(
        n19185) );
  AOI22_X1 U22378 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19190), .B1(
        n19459), .B2(n19260), .ZN(n19184) );
  OAI211_X1 U22379 ( .C1(n19462), .C2(n19213), .A(n19185), .B(n19184), .ZN(
        P3_U2913) );
  AOI22_X1 U22380 ( .A1(n19324), .A2(n19186), .B1(n19463), .B2(n19189), .ZN(
        n19188) );
  AOI22_X1 U22381 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19190), .B1(
        n19466), .B2(n19260), .ZN(n19187) );
  OAI211_X1 U22382 ( .C1(n19327), .C2(n19213), .A(n19188), .B(n19187), .ZN(
        P3_U2914) );
  AOI22_X1 U22383 ( .A1(n19415), .A2(n19215), .B1(n19472), .B2(n19189), .ZN(
        n19192) );
  AOI22_X1 U22384 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19190), .B1(
        n19475), .B2(n19260), .ZN(n19191) );
  OAI211_X1 U22385 ( .C1(n19421), .C2(n19193), .A(n19192), .B(n19191), .ZN(
        P3_U2915) );
  NOR2_X1 U22386 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19194), .ZN(
        n19266) );
  NAND2_X1 U22387 ( .A1(n19266), .A2(n19195), .ZN(n19277) );
  INV_X1 U22388 ( .A(n19277), .ZN(n19282) );
  NOR2_X1 U22389 ( .A1(n19260), .A2(n19282), .ZN(n19242) );
  NOR2_X1 U22390 ( .A1(n19388), .A2(n19242), .ZN(n19214) );
  AOI22_X1 U22391 ( .A1(n19389), .A2(n19215), .B1(n19422), .B2(n19214), .ZN(
        n19200) );
  AOI221_X1 U22392 ( .B1(n19242), .B2(n19391), .C1(n19242), .C2(n19197), .A(
        n19196), .ZN(n19198) );
  INV_X1 U22393 ( .A(n19198), .ZN(n19216) );
  AOI22_X1 U22394 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19216), .B1(
        n19423), .B2(n19234), .ZN(n19199) );
  OAI211_X1 U22395 ( .C1(n19397), .C2(n19277), .A(n19200), .B(n19199), .ZN(
        P3_U2916) );
  AOI22_X1 U22396 ( .A1(n19340), .A2(n19234), .B1(n19432), .B2(n19214), .ZN(
        n19202) );
  AOI22_X1 U22397 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19216), .B1(
        n19433), .B2(n19215), .ZN(n19201) );
  OAI211_X1 U22398 ( .C1(n19343), .C2(n19277), .A(n19202), .B(n19201), .ZN(
        P3_U2917) );
  AOI22_X1 U22399 ( .A1(n19369), .A2(n19215), .B1(n19438), .B2(n19214), .ZN(
        n19204) );
  AOI22_X1 U22400 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19216), .B1(
        n19440), .B2(n19282), .ZN(n19203) );
  OAI211_X1 U22401 ( .C1(n19372), .C2(n19241), .A(n19204), .B(n19203), .ZN(
        P3_U2918) );
  AOI22_X1 U22402 ( .A1(n19445), .A2(n19215), .B1(n19444), .B2(n19214), .ZN(
        n19206) );
  AOI22_X1 U22403 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19216), .B1(
        n19446), .B2(n19234), .ZN(n19205) );
  OAI211_X1 U22404 ( .C1(n19449), .C2(n19277), .A(n19206), .B(n19205), .ZN(
        P3_U2919) );
  AOI22_X1 U22405 ( .A1(n19452), .A2(n19215), .B1(n19451), .B2(n19214), .ZN(
        n19208) );
  AOI22_X1 U22406 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19216), .B1(
        n19453), .B2(n19282), .ZN(n19207) );
  OAI211_X1 U22407 ( .C1(n19456), .C2(n19241), .A(n19208), .B(n19207), .ZN(
        P3_U2920) );
  AOI22_X1 U22408 ( .A1(n19458), .A2(n19215), .B1(n19457), .B2(n19214), .ZN(
        n19210) );
  AOI22_X1 U22409 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19216), .B1(
        n19459), .B2(n19282), .ZN(n19209) );
  OAI211_X1 U22410 ( .C1(n19462), .C2(n19241), .A(n19210), .B(n19209), .ZN(
        P3_U2921) );
  AOI22_X1 U22411 ( .A1(n19463), .A2(n19214), .B1(n19464), .B2(n19234), .ZN(
        n19212) );
  AOI22_X1 U22412 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19216), .B1(
        n19466), .B2(n19282), .ZN(n19211) );
  OAI211_X1 U22413 ( .C1(n19470), .C2(n19213), .A(n19212), .B(n19211), .ZN(
        P3_U2922) );
  AOI22_X1 U22414 ( .A1(n19474), .A2(n19215), .B1(n19472), .B2(n19214), .ZN(
        n19218) );
  AOI22_X1 U22415 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19216), .B1(
        n19475), .B2(n19282), .ZN(n19217) );
  OAI211_X1 U22416 ( .C1(n19480), .C2(n19241), .A(n19218), .B(n19217), .ZN(
        P3_U2923) );
  NAND2_X1 U22417 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19266), .ZN(
        n19297) );
  AND2_X1 U22418 ( .A1(n19550), .A2(n19266), .ZN(n19237) );
  AOI22_X1 U22419 ( .A1(n19423), .A2(n19260), .B1(n19422), .B2(n19237), .ZN(
        n19223) );
  NAND3_X1 U22420 ( .A1(n19221), .A2(n19220), .A3(n19219), .ZN(n19238) );
  AOI22_X1 U22421 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19238), .B1(
        n19389), .B2(n19234), .ZN(n19222) );
  OAI211_X1 U22422 ( .C1(n19397), .C2(n19297), .A(n19223), .B(n19222), .ZN(
        P3_U2924) );
  AOI22_X1 U22423 ( .A1(n19340), .A2(n19260), .B1(n19432), .B2(n19237), .ZN(
        n19225) );
  AOI22_X1 U22424 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19238), .B1(
        n19433), .B2(n19234), .ZN(n19224) );
  OAI211_X1 U22425 ( .C1(n19343), .C2(n19297), .A(n19225), .B(n19224), .ZN(
        P3_U2925) );
  AOI22_X1 U22426 ( .A1(n19439), .A2(n19260), .B1(n19438), .B2(n19237), .ZN(
        n19227) );
  INV_X1 U22427 ( .A(n19297), .ZN(n19305) );
  AOI22_X1 U22428 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19238), .B1(
        n19440), .B2(n19305), .ZN(n19226) );
  OAI211_X1 U22429 ( .C1(n19443), .C2(n19241), .A(n19227), .B(n19226), .ZN(
        P3_U2926) );
  AOI22_X1 U22430 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19238), .B1(
        n19444), .B2(n19237), .ZN(n19229) );
  AOI22_X1 U22431 ( .A1(n19403), .A2(n19305), .B1(n19446), .B2(n19260), .ZN(
        n19228) );
  OAI211_X1 U22432 ( .C1(n19406), .C2(n19241), .A(n19229), .B(n19228), .ZN(
        P3_U2927) );
  AOI22_X1 U22433 ( .A1(n19375), .A2(n19260), .B1(n19451), .B2(n19237), .ZN(
        n19231) );
  AOI22_X1 U22434 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19238), .B1(
        n19453), .B2(n19305), .ZN(n19230) );
  OAI211_X1 U22435 ( .C1(n19378), .C2(n19241), .A(n19231), .B(n19230), .ZN(
        P3_U2928) );
  AOI22_X1 U22436 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19238), .B1(
        n19457), .B2(n19237), .ZN(n19233) );
  AOI22_X1 U22437 ( .A1(n19459), .A2(n19305), .B1(n19458), .B2(n19234), .ZN(
        n19232) );
  OAI211_X1 U22438 ( .C1(n19462), .C2(n19258), .A(n19233), .B(n19232), .ZN(
        P3_U2929) );
  AOI22_X1 U22439 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19238), .B1(
        n19463), .B2(n19237), .ZN(n19236) );
  AOI22_X1 U22440 ( .A1(n19324), .A2(n19234), .B1(n19466), .B2(n19305), .ZN(
        n19235) );
  OAI211_X1 U22441 ( .C1(n19327), .C2(n19258), .A(n19236), .B(n19235), .ZN(
        P3_U2930) );
  AOI22_X1 U22442 ( .A1(n19415), .A2(n19260), .B1(n19472), .B2(n19237), .ZN(
        n19240) );
  AOI22_X1 U22443 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19238), .B1(
        n19475), .B2(n19305), .ZN(n19239) );
  OAI211_X1 U22444 ( .C1(n19421), .C2(n19241), .A(n19240), .B(n19239), .ZN(
        P3_U2931) );
  NAND2_X1 U22445 ( .A1(n19333), .A2(n19286), .ZN(n19317) );
  NOR2_X1 U22446 ( .A1(n19305), .A2(n19329), .ZN(n19287) );
  NOR2_X1 U22447 ( .A1(n19388), .A2(n19287), .ZN(n19259) );
  AOI22_X1 U22448 ( .A1(n19389), .A2(n19260), .B1(n19422), .B2(n19259), .ZN(
        n19245) );
  OAI21_X1 U22449 ( .B1(n19242), .B2(n19391), .A(n19287), .ZN(n19243) );
  OAI211_X1 U22450 ( .C1(n19329), .C2(n19650), .A(n19394), .B(n19243), .ZN(
        n19261) );
  AOI22_X1 U22451 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19261), .B1(
        n19423), .B2(n19282), .ZN(n19244) );
  OAI211_X1 U22452 ( .C1(n19397), .C2(n19317), .A(n19245), .B(n19244), .ZN(
        P3_U2932) );
  AOI22_X1 U22453 ( .A1(n19340), .A2(n19282), .B1(n19432), .B2(n19259), .ZN(
        n19247) );
  AOI22_X1 U22454 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19261), .B1(
        n19433), .B2(n19260), .ZN(n19246) );
  OAI211_X1 U22455 ( .C1(n19343), .C2(n19317), .A(n19247), .B(n19246), .ZN(
        P3_U2933) );
  AOI22_X1 U22456 ( .A1(n19369), .A2(n19260), .B1(n19438), .B2(n19259), .ZN(
        n19249) );
  AOI22_X1 U22457 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19261), .B1(
        n19440), .B2(n19329), .ZN(n19248) );
  OAI211_X1 U22458 ( .C1(n19372), .C2(n19277), .A(n19249), .B(n19248), .ZN(
        P3_U2934) );
  AOI22_X1 U22459 ( .A1(n19445), .A2(n19260), .B1(n19444), .B2(n19259), .ZN(
        n19251) );
  AOI22_X1 U22460 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19261), .B1(
        n19446), .B2(n19282), .ZN(n19250) );
  OAI211_X1 U22461 ( .C1(n19449), .C2(n19317), .A(n19251), .B(n19250), .ZN(
        P3_U2935) );
  AOI22_X1 U22462 ( .A1(n19375), .A2(n19282), .B1(n19451), .B2(n19259), .ZN(
        n19253) );
  AOI22_X1 U22463 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19261), .B1(
        n19453), .B2(n19329), .ZN(n19252) );
  OAI211_X1 U22464 ( .C1(n19378), .C2(n19258), .A(n19253), .B(n19252), .ZN(
        P3_U2936) );
  AOI22_X1 U22465 ( .A1(n19458), .A2(n19260), .B1(n19457), .B2(n19259), .ZN(
        n19255) );
  AOI22_X1 U22466 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19261), .B1(
        n19459), .B2(n19329), .ZN(n19254) );
  OAI211_X1 U22467 ( .C1(n19462), .C2(n19277), .A(n19255), .B(n19254), .ZN(
        P3_U2937) );
  AOI22_X1 U22468 ( .A1(n19463), .A2(n19259), .B1(n19464), .B2(n19282), .ZN(
        n19257) );
  AOI22_X1 U22469 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19261), .B1(
        n19466), .B2(n19329), .ZN(n19256) );
  OAI211_X1 U22470 ( .C1(n19470), .C2(n19258), .A(n19257), .B(n19256), .ZN(
        P3_U2938) );
  AOI22_X1 U22471 ( .A1(n19474), .A2(n19260), .B1(n19472), .B2(n19259), .ZN(
        n19263) );
  AOI22_X1 U22472 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19261), .B1(
        n19475), .B2(n19329), .ZN(n19262) );
  OAI211_X1 U22473 ( .C1(n19480), .C2(n19277), .A(n19263), .B(n19262), .ZN(
        P3_U2939) );
  NAND2_X1 U22474 ( .A1(n19264), .A2(n19286), .ZN(n19354) );
  INV_X1 U22475 ( .A(n19286), .ZN(n19265) );
  NOR2_X1 U22476 ( .A1(n19360), .A2(n19265), .ZN(n19310) );
  AOI22_X1 U22477 ( .A1(n19389), .A2(n19282), .B1(n19422), .B2(n19310), .ZN(
        n19268) );
  AOI22_X1 U22478 ( .A1(n19427), .A2(n19266), .B1(n19362), .B2(n19286), .ZN(
        n19283) );
  AOI22_X1 U22479 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19283), .B1(
        n19423), .B2(n19305), .ZN(n19267) );
  OAI211_X1 U22480 ( .C1(n19397), .C2(n19354), .A(n19268), .B(n19267), .ZN(
        P3_U2940) );
  AOI22_X1 U22481 ( .A1(n19340), .A2(n19305), .B1(n19432), .B2(n19310), .ZN(
        n19270) );
  AOI22_X1 U22482 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19283), .B1(
        n19433), .B2(n19282), .ZN(n19269) );
  OAI211_X1 U22483 ( .C1(n19343), .C2(n19354), .A(n19270), .B(n19269), .ZN(
        P3_U2941) );
  AOI22_X1 U22484 ( .A1(n19439), .A2(n19305), .B1(n19438), .B2(n19310), .ZN(
        n19272) );
  INV_X1 U22485 ( .A(n19354), .ZN(n19356) );
  AOI22_X1 U22486 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19283), .B1(
        n19440), .B2(n19356), .ZN(n19271) );
  OAI211_X1 U22487 ( .C1(n19443), .C2(n19277), .A(n19272), .B(n19271), .ZN(
        P3_U2942) );
  AOI22_X1 U22488 ( .A1(n19445), .A2(n19282), .B1(n19444), .B2(n19310), .ZN(
        n19274) );
  AOI22_X1 U22489 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19283), .B1(
        n19446), .B2(n19305), .ZN(n19273) );
  OAI211_X1 U22490 ( .C1(n19449), .C2(n19354), .A(n19274), .B(n19273), .ZN(
        P3_U2943) );
  AOI22_X1 U22491 ( .A1(n19375), .A2(n19305), .B1(n19451), .B2(n19310), .ZN(
        n19276) );
  AOI22_X1 U22492 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19283), .B1(
        n19453), .B2(n19356), .ZN(n19275) );
  OAI211_X1 U22493 ( .C1(n19378), .C2(n19277), .A(n19276), .B(n19275), .ZN(
        P3_U2944) );
  AOI22_X1 U22494 ( .A1(n19458), .A2(n19282), .B1(n19457), .B2(n19310), .ZN(
        n19279) );
  AOI22_X1 U22495 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19283), .B1(
        n19459), .B2(n19356), .ZN(n19278) );
  OAI211_X1 U22496 ( .C1(n19462), .C2(n19297), .A(n19279), .B(n19278), .ZN(
        P3_U2945) );
  AOI22_X1 U22497 ( .A1(n19324), .A2(n19282), .B1(n19463), .B2(n19310), .ZN(
        n19281) );
  AOI22_X1 U22498 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19283), .B1(
        n19466), .B2(n19356), .ZN(n19280) );
  OAI211_X1 U22499 ( .C1(n19327), .C2(n19297), .A(n19281), .B(n19280), .ZN(
        P3_U2946) );
  AOI22_X1 U22500 ( .A1(n19474), .A2(n19282), .B1(n19472), .B2(n19310), .ZN(
        n19285) );
  AOI22_X1 U22501 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19283), .B1(
        n19475), .B2(n19356), .ZN(n19284) );
  OAI211_X1 U22502 ( .C1(n19480), .C2(n19297), .A(n19285), .B(n19284), .ZN(
        P3_U2947) );
  NAND2_X1 U22503 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19286), .ZN(
        n19309) );
  NOR2_X2 U22504 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19309), .ZN(
        n19379) );
  NOR2_X1 U22505 ( .A1(n19356), .A2(n19379), .ZN(n19336) );
  NOR2_X1 U22506 ( .A1(n19388), .A2(n19336), .ZN(n19304) );
  AOI22_X1 U22507 ( .A1(n19423), .A2(n19329), .B1(n19422), .B2(n19304), .ZN(
        n19290) );
  OAI21_X1 U22508 ( .B1(n19287), .B2(n19391), .A(n19336), .ZN(n19288) );
  OAI211_X1 U22509 ( .C1(n19379), .C2(n19650), .A(n19394), .B(n19288), .ZN(
        n19306) );
  AOI22_X1 U22510 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19306), .B1(
        n19428), .B2(n19379), .ZN(n19289) );
  OAI211_X1 U22511 ( .C1(n19431), .C2(n19297), .A(n19290), .B(n19289), .ZN(
        P3_U2948) );
  INV_X1 U22512 ( .A(n19379), .ZN(n19387) );
  AOI22_X1 U22513 ( .A1(n19340), .A2(n19329), .B1(n19432), .B2(n19304), .ZN(
        n19292) );
  AOI22_X1 U22514 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19306), .B1(
        n19433), .B2(n19305), .ZN(n19291) );
  OAI211_X1 U22515 ( .C1(n19343), .C2(n19387), .A(n19292), .B(n19291), .ZN(
        P3_U2949) );
  AOI22_X1 U22516 ( .A1(n19439), .A2(n19329), .B1(n19438), .B2(n19304), .ZN(
        n19294) );
  AOI22_X1 U22517 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19306), .B1(
        n19440), .B2(n19379), .ZN(n19293) );
  OAI211_X1 U22518 ( .C1(n19443), .C2(n19297), .A(n19294), .B(n19293), .ZN(
        P3_U2950) );
  AOI22_X1 U22519 ( .A1(n19446), .A2(n19329), .B1(n19444), .B2(n19304), .ZN(
        n19296) );
  AOI22_X1 U22520 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19306), .B1(
        n19403), .B2(n19379), .ZN(n19295) );
  OAI211_X1 U22521 ( .C1(n19406), .C2(n19297), .A(n19296), .B(n19295), .ZN(
        P3_U2951) );
  AOI22_X1 U22522 ( .A1(n19452), .A2(n19305), .B1(n19451), .B2(n19304), .ZN(
        n19299) );
  AOI22_X1 U22523 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19306), .B1(
        n19453), .B2(n19379), .ZN(n19298) );
  OAI211_X1 U22524 ( .C1(n19456), .C2(n19317), .A(n19299), .B(n19298), .ZN(
        P3_U2952) );
  AOI22_X1 U22525 ( .A1(n19458), .A2(n19305), .B1(n19457), .B2(n19304), .ZN(
        n19301) );
  AOI22_X1 U22526 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19306), .B1(
        n19459), .B2(n19379), .ZN(n19300) );
  OAI211_X1 U22527 ( .C1(n19462), .C2(n19317), .A(n19301), .B(n19300), .ZN(
        P3_U2953) );
  AOI22_X1 U22528 ( .A1(n19324), .A2(n19305), .B1(n19463), .B2(n19304), .ZN(
        n19303) );
  AOI22_X1 U22529 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19306), .B1(
        n19466), .B2(n19379), .ZN(n19302) );
  OAI211_X1 U22530 ( .C1(n19327), .C2(n19317), .A(n19303), .B(n19302), .ZN(
        P3_U2954) );
  AOI22_X1 U22531 ( .A1(n19474), .A2(n19305), .B1(n19472), .B2(n19304), .ZN(
        n19308) );
  AOI22_X1 U22532 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19306), .B1(
        n19475), .B2(n19379), .ZN(n19307) );
  OAI211_X1 U22533 ( .C1(n19480), .C2(n19317), .A(n19308), .B(n19307), .ZN(
        P3_U2955) );
  INV_X1 U22534 ( .A(n19309), .ZN(n19364) );
  NAND2_X1 U22535 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19364), .ZN(
        n19420) );
  NOR2_X1 U22536 ( .A1(n19388), .A2(n19309), .ZN(n19328) );
  AOI22_X1 U22537 ( .A1(n19389), .A2(n19329), .B1(n19422), .B2(n19328), .ZN(
        n19312) );
  AOI22_X1 U22538 ( .A1(n19427), .A2(n19310), .B1(n19424), .B2(n19364), .ZN(
        n19330) );
  AOI22_X1 U22539 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19330), .B1(
        n19423), .B2(n19356), .ZN(n19311) );
  OAI211_X1 U22540 ( .C1(n19397), .C2(n19420), .A(n19312), .B(n19311), .ZN(
        P3_U2956) );
  AOI22_X1 U22541 ( .A1(n19433), .A2(n19329), .B1(n19432), .B2(n19328), .ZN(
        n19314) );
  AOI22_X1 U22542 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19330), .B1(
        n19340), .B2(n19356), .ZN(n19313) );
  OAI211_X1 U22543 ( .C1(n19343), .C2(n19420), .A(n19314), .B(n19313), .ZN(
        P3_U2957) );
  AOI22_X1 U22544 ( .A1(n19439), .A2(n19356), .B1(n19438), .B2(n19328), .ZN(
        n19316) );
  INV_X1 U22545 ( .A(n19420), .ZN(n19409) );
  AOI22_X1 U22546 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19330), .B1(
        n19440), .B2(n19409), .ZN(n19315) );
  OAI211_X1 U22547 ( .C1(n19443), .C2(n19317), .A(n19316), .B(n19315), .ZN(
        P3_U2958) );
  AOI22_X1 U22548 ( .A1(n19445), .A2(n19329), .B1(n19444), .B2(n19328), .ZN(
        n19319) );
  AOI22_X1 U22549 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19330), .B1(
        n19446), .B2(n19356), .ZN(n19318) );
  OAI211_X1 U22550 ( .C1(n19449), .C2(n19420), .A(n19319), .B(n19318), .ZN(
        P3_U2959) );
  AOI22_X1 U22551 ( .A1(n19452), .A2(n19329), .B1(n19451), .B2(n19328), .ZN(
        n19321) );
  AOI22_X1 U22552 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19330), .B1(
        n19453), .B2(n19409), .ZN(n19320) );
  OAI211_X1 U22553 ( .C1(n19456), .C2(n19354), .A(n19321), .B(n19320), .ZN(
        P3_U2960) );
  AOI22_X1 U22554 ( .A1(n19458), .A2(n19329), .B1(n19457), .B2(n19328), .ZN(
        n19323) );
  AOI22_X1 U22555 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19330), .B1(
        n19459), .B2(n19409), .ZN(n19322) );
  OAI211_X1 U22556 ( .C1(n19462), .C2(n19354), .A(n19323), .B(n19322), .ZN(
        P3_U2961) );
  AOI22_X1 U22557 ( .A1(n19324), .A2(n19329), .B1(n19463), .B2(n19328), .ZN(
        n19326) );
  AOI22_X1 U22558 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19330), .B1(
        n19466), .B2(n19409), .ZN(n19325) );
  OAI211_X1 U22559 ( .C1(n19327), .C2(n19354), .A(n19326), .B(n19325), .ZN(
        P3_U2962) );
  AOI22_X1 U22560 ( .A1(n19474), .A2(n19329), .B1(n19472), .B2(n19328), .ZN(
        n19332) );
  AOI22_X1 U22561 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19330), .B1(
        n19475), .B2(n19409), .ZN(n19331) );
  OAI211_X1 U22562 ( .C1(n19480), .C2(n19354), .A(n19332), .B(n19331), .ZN(
        P3_U2963) );
  NAND2_X1 U22563 ( .A1(n19333), .A2(n19363), .ZN(n19469) );
  INV_X1 U22564 ( .A(n19469), .ZN(n19473) );
  NOR2_X1 U22565 ( .A1(n19409), .A2(n19473), .ZN(n19392) );
  NOR2_X1 U22566 ( .A1(n19388), .A2(n19392), .ZN(n19355) );
  AOI22_X1 U22567 ( .A1(n19423), .A2(n19379), .B1(n19422), .B2(n19355), .ZN(
        n19339) );
  OAI22_X1 U22568 ( .A1(n19336), .A2(n19335), .B1(n19392), .B2(n19334), .ZN(
        n19337) );
  OAI21_X1 U22569 ( .B1(n19473), .B2(n19650), .A(n19337), .ZN(n19357) );
  AOI22_X1 U22570 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19357), .B1(
        n19389), .B2(n19356), .ZN(n19338) );
  OAI211_X1 U22571 ( .C1(n19397), .C2(n19469), .A(n19339), .B(n19338), .ZN(
        P3_U2964) );
  AOI22_X1 U22572 ( .A1(n19340), .A2(n19379), .B1(n19432), .B2(n19355), .ZN(
        n19342) );
  AOI22_X1 U22573 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19357), .B1(
        n19433), .B2(n19356), .ZN(n19341) );
  OAI211_X1 U22574 ( .C1(n19343), .C2(n19469), .A(n19342), .B(n19341), .ZN(
        P3_U2965) );
  AOI22_X1 U22575 ( .A1(n19369), .A2(n19356), .B1(n19438), .B2(n19355), .ZN(
        n19345) );
  AOI22_X1 U22576 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19357), .B1(
        n19440), .B2(n19473), .ZN(n19344) );
  OAI211_X1 U22577 ( .C1(n19372), .C2(n19387), .A(n19345), .B(n19344), .ZN(
        P3_U2966) );
  AOI22_X1 U22578 ( .A1(n19445), .A2(n19356), .B1(n19444), .B2(n19355), .ZN(
        n19347) );
  AOI22_X1 U22579 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19357), .B1(
        n19446), .B2(n19379), .ZN(n19346) );
  OAI211_X1 U22580 ( .C1(n19449), .C2(n19469), .A(n19347), .B(n19346), .ZN(
        P3_U2967) );
  AOI22_X1 U22581 ( .A1(n19375), .A2(n19379), .B1(n19451), .B2(n19355), .ZN(
        n19349) );
  AOI22_X1 U22582 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19357), .B1(
        n19453), .B2(n19473), .ZN(n19348) );
  OAI211_X1 U22583 ( .C1(n19378), .C2(n19354), .A(n19349), .B(n19348), .ZN(
        P3_U2968) );
  AOI22_X1 U22584 ( .A1(n19458), .A2(n19356), .B1(n19457), .B2(n19355), .ZN(
        n19351) );
  AOI22_X1 U22585 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19357), .B1(
        n19459), .B2(n19473), .ZN(n19350) );
  OAI211_X1 U22586 ( .C1(n19462), .C2(n19387), .A(n19351), .B(n19350), .ZN(
        P3_U2969) );
  AOI22_X1 U22587 ( .A1(n19463), .A2(n19355), .B1(n19464), .B2(n19379), .ZN(
        n19353) );
  AOI22_X1 U22588 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19357), .B1(
        n19466), .B2(n19473), .ZN(n19352) );
  OAI211_X1 U22589 ( .C1(n19470), .C2(n19354), .A(n19353), .B(n19352), .ZN(
        P3_U2970) );
  AOI22_X1 U22590 ( .A1(n19474), .A2(n19356), .B1(n19472), .B2(n19355), .ZN(
        n19359) );
  AOI22_X1 U22591 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19357), .B1(
        n19475), .B2(n19473), .ZN(n19358) );
  OAI211_X1 U22592 ( .C1(n19480), .C2(n19387), .A(n19359), .B(n19358), .ZN(
        P3_U2971) );
  INV_X1 U22593 ( .A(n19363), .ZN(n19361) );
  NOR2_X1 U22594 ( .A1(n19361), .A2(n19360), .ZN(n19426) );
  AOI22_X1 U22595 ( .A1(n19389), .A2(n19379), .B1(n19422), .B2(n19426), .ZN(
        n19366) );
  AOI22_X1 U22596 ( .A1(n19427), .A2(n19364), .B1(n19363), .B2(n19362), .ZN(
        n19384) );
  AOI22_X1 U22597 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19384), .B1(
        n19423), .B2(n19409), .ZN(n19365) );
  OAI211_X1 U22598 ( .C1(n19481), .C2(n19397), .A(n19366), .B(n19365), .ZN(
        P3_U2972) );
  AOI22_X1 U22599 ( .A1(n19433), .A2(n19379), .B1(n19432), .B2(n19426), .ZN(
        n19368) );
  AOI22_X1 U22600 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19384), .B1(
        n19465), .B2(n19434), .ZN(n19367) );
  OAI211_X1 U22601 ( .C1(n19437), .C2(n19420), .A(n19368), .B(n19367), .ZN(
        P3_U2973) );
  AOI22_X1 U22602 ( .A1(n19369), .A2(n19379), .B1(n19438), .B2(n19426), .ZN(
        n19371) );
  AOI22_X1 U22603 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19384), .B1(
        n19465), .B2(n19440), .ZN(n19370) );
  OAI211_X1 U22604 ( .C1(n19372), .C2(n19420), .A(n19371), .B(n19370), .ZN(
        P3_U2974) );
  AOI22_X1 U22605 ( .A1(n19445), .A2(n19379), .B1(n19444), .B2(n19426), .ZN(
        n19374) );
  AOI22_X1 U22606 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19384), .B1(
        n19446), .B2(n19409), .ZN(n19373) );
  OAI211_X1 U22607 ( .C1(n19481), .C2(n19449), .A(n19374), .B(n19373), .ZN(
        P3_U2975) );
  AOI22_X1 U22608 ( .A1(n19375), .A2(n19409), .B1(n19451), .B2(n19426), .ZN(
        n19377) );
  AOI22_X1 U22609 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19384), .B1(
        n19465), .B2(n19453), .ZN(n19376) );
  OAI211_X1 U22610 ( .C1(n19378), .C2(n19387), .A(n19377), .B(n19376), .ZN(
        P3_U2976) );
  AOI22_X1 U22611 ( .A1(n19458), .A2(n19379), .B1(n19457), .B2(n19426), .ZN(
        n19381) );
  AOI22_X1 U22612 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19384), .B1(
        n19465), .B2(n19459), .ZN(n19380) );
  OAI211_X1 U22613 ( .C1(n19462), .C2(n19420), .A(n19381), .B(n19380), .ZN(
        P3_U2977) );
  AOI22_X1 U22614 ( .A1(n19463), .A2(n19426), .B1(n19464), .B2(n19409), .ZN(
        n19383) );
  AOI22_X1 U22615 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19384), .B1(
        n19465), .B2(n19466), .ZN(n19382) );
  OAI211_X1 U22616 ( .C1(n19470), .C2(n19387), .A(n19383), .B(n19382), .ZN(
        P3_U2978) );
  AOI22_X1 U22617 ( .A1(n19415), .A2(n19409), .B1(n19472), .B2(n19426), .ZN(
        n19386) );
  AOI22_X1 U22618 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19384), .B1(
        n19465), .B2(n19475), .ZN(n19385) );
  OAI211_X1 U22619 ( .C1(n19421), .C2(n19387), .A(n19386), .B(n19385), .ZN(
        P3_U2979) );
  NOR2_X1 U22620 ( .A1(n19388), .A2(n19390), .ZN(n19414) );
  AOI22_X1 U22621 ( .A1(n19389), .A2(n19409), .B1(n19422), .B2(n19414), .ZN(
        n19396) );
  OAI21_X1 U22622 ( .B1(n19392), .B2(n19391), .A(n19390), .ZN(n19393) );
  OAI211_X1 U22623 ( .C1(n19416), .C2(n19650), .A(n19394), .B(n19393), .ZN(
        n19417) );
  AOI22_X1 U22624 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19417), .B1(
        n19423), .B2(n19473), .ZN(n19395) );
  OAI211_X1 U22625 ( .C1(n19398), .C2(n19397), .A(n19396), .B(n19395), .ZN(
        P3_U2980) );
  AOI22_X1 U22626 ( .A1(n19433), .A2(n19409), .B1(n19432), .B2(n19414), .ZN(
        n19400) );
  AOI22_X1 U22627 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19434), .ZN(n19399) );
  OAI211_X1 U22628 ( .C1(n19437), .C2(n19469), .A(n19400), .B(n19399), .ZN(
        P3_U2981) );
  AOI22_X1 U22629 ( .A1(n19439), .A2(n19473), .B1(n19438), .B2(n19414), .ZN(
        n19402) );
  AOI22_X1 U22630 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19440), .ZN(n19401) );
  OAI211_X1 U22631 ( .C1(n19443), .C2(n19420), .A(n19402), .B(n19401), .ZN(
        P3_U2982) );
  AOI22_X1 U22632 ( .A1(n19446), .A2(n19473), .B1(n19444), .B2(n19414), .ZN(
        n19405) );
  AOI22_X1 U22633 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19403), .ZN(n19404) );
  OAI211_X1 U22634 ( .C1(n19406), .C2(n19420), .A(n19405), .B(n19404), .ZN(
        P3_U2983) );
  AOI22_X1 U22635 ( .A1(n19452), .A2(n19409), .B1(n19451), .B2(n19414), .ZN(
        n19408) );
  AOI22_X1 U22636 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19453), .ZN(n19407) );
  OAI211_X1 U22637 ( .C1(n19456), .C2(n19469), .A(n19408), .B(n19407), .ZN(
        P3_U2984) );
  AOI22_X1 U22638 ( .A1(n19458), .A2(n19409), .B1(n19457), .B2(n19414), .ZN(
        n19411) );
  AOI22_X1 U22639 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19459), .ZN(n19410) );
  OAI211_X1 U22640 ( .C1(n19462), .C2(n19469), .A(n19411), .B(n19410), .ZN(
        P3_U2985) );
  AOI22_X1 U22641 ( .A1(n19463), .A2(n19414), .B1(n19464), .B2(n19473), .ZN(
        n19413) );
  AOI22_X1 U22642 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19466), .ZN(n19412) );
  OAI211_X1 U22643 ( .C1(n19470), .C2(n19420), .A(n19413), .B(n19412), .ZN(
        P3_U2986) );
  AOI22_X1 U22644 ( .A1(n19415), .A2(n19473), .B1(n19472), .B2(n19414), .ZN(
        n19419) );
  AOI22_X1 U22645 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19417), .B1(
        n19416), .B2(n19475), .ZN(n19418) );
  OAI211_X1 U22646 ( .C1(n19421), .C2(n19420), .A(n19419), .B(n19418), .ZN(
        P3_U2987) );
  AND2_X1 U22647 ( .A1(n19550), .A2(n19425), .ZN(n19471) );
  AOI22_X1 U22648 ( .A1(n19465), .A2(n19423), .B1(n19422), .B2(n19471), .ZN(
        n19430) );
  AOI22_X1 U22649 ( .A1(n19427), .A2(n19426), .B1(n19425), .B2(n19424), .ZN(
        n19477) );
  AOI22_X1 U22650 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19477), .B1(
        n19476), .B2(n19428), .ZN(n19429) );
  OAI211_X1 U22651 ( .C1(n19431), .C2(n19469), .A(n19430), .B(n19429), .ZN(
        P3_U2988) );
  AOI22_X1 U22652 ( .A1(n19433), .A2(n19473), .B1(n19432), .B2(n19471), .ZN(
        n19436) );
  AOI22_X1 U22653 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19477), .B1(
        n19476), .B2(n19434), .ZN(n19435) );
  OAI211_X1 U22654 ( .C1(n19481), .C2(n19437), .A(n19436), .B(n19435), .ZN(
        P3_U2989) );
  AOI22_X1 U22655 ( .A1(n19465), .A2(n19439), .B1(n19438), .B2(n19471), .ZN(
        n19442) );
  AOI22_X1 U22656 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19477), .B1(
        n19476), .B2(n19440), .ZN(n19441) );
  OAI211_X1 U22657 ( .C1(n19443), .C2(n19469), .A(n19442), .B(n19441), .ZN(
        P3_U2990) );
  AOI22_X1 U22658 ( .A1(n19445), .A2(n19473), .B1(n19444), .B2(n19471), .ZN(
        n19448) );
  AOI22_X1 U22659 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19477), .B1(
        n19465), .B2(n19446), .ZN(n19447) );
  OAI211_X1 U22660 ( .C1(n19450), .C2(n19449), .A(n19448), .B(n19447), .ZN(
        P3_U2991) );
  AOI22_X1 U22661 ( .A1(n19452), .A2(n19473), .B1(n19451), .B2(n19471), .ZN(
        n19455) );
  AOI22_X1 U22662 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19477), .B1(
        n19476), .B2(n19453), .ZN(n19454) );
  OAI211_X1 U22663 ( .C1(n19481), .C2(n19456), .A(n19455), .B(n19454), .ZN(
        P3_U2992) );
  AOI22_X1 U22664 ( .A1(n19458), .A2(n19473), .B1(n19457), .B2(n19471), .ZN(
        n19461) );
  AOI22_X1 U22665 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19477), .B1(
        n19476), .B2(n19459), .ZN(n19460) );
  OAI211_X1 U22666 ( .C1(n19481), .C2(n19462), .A(n19461), .B(n19460), .ZN(
        P3_U2993) );
  AOI22_X1 U22667 ( .A1(n19465), .A2(n19464), .B1(n19463), .B2(n19471), .ZN(
        n19468) );
  AOI22_X1 U22668 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19477), .B1(
        n19476), .B2(n19466), .ZN(n19467) );
  OAI211_X1 U22669 ( .C1(n19470), .C2(n19469), .A(n19468), .B(n19467), .ZN(
        P3_U2994) );
  AOI22_X1 U22670 ( .A1(n19474), .A2(n19473), .B1(n19472), .B2(n19471), .ZN(
        n19479) );
  AOI22_X1 U22671 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19477), .B1(
        n19476), .B2(n19475), .ZN(n19478) );
  OAI211_X1 U22672 ( .C1(n19481), .C2(n19480), .A(n19479), .B(n19478), .ZN(
        P3_U2995) );
  INV_X1 U22673 ( .A(n19482), .ZN(n19487) );
  NAND2_X1 U22674 ( .A1(n19483), .A2(n19487), .ZN(n19484) );
  NAND2_X1 U22675 ( .A1(n19485), .A2(n19484), .ZN(n19507) );
  NOR2_X1 U22676 ( .A1(n19487), .A2(n19486), .ZN(n19490) );
  INV_X1 U22677 ( .A(n19488), .ZN(n19489) );
  NAND4_X1 U22678 ( .A1(n19491), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n19490), .A4(n19489), .ZN(n19492) );
  AOI22_X1 U22679 ( .A1(n13162), .A2(n19507), .B1(n19493), .B2(n19492), .ZN(
        n19498) );
  AOI22_X1 U22680 ( .A1(n19512), .A2(n19497), .B1(n19502), .B2(n19495), .ZN(
        n19496) );
  AOI22_X1 U22681 ( .A1(n19498), .A2(n19497), .B1(n19496), .B2(n19654), .ZN(
        n19652) );
  AOI22_X1 U22682 ( .A1(n19513), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19652), .B2(n19534), .ZN(n19519) );
  NOR2_X1 U22683 ( .A1(n19500), .A2(n19499), .ZN(n19503) );
  AOI22_X1 U22684 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19501), .B1(
        n19503), .B2(n13162), .ZN(n19672) );
  NOR2_X1 U22685 ( .A1(n19672), .A2(n21428), .ZN(n19506) );
  OAI22_X1 U22686 ( .A1(n19503), .A2(n19664), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19509), .ZN(n19669) );
  OAI221_X1 U22687 ( .B1(n19669), .B2(n19672), .C1(n19669), .C2(n21428), .A(
        n19534), .ZN(n19504) );
  AOI22_X1 U22688 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19506), .B1(
        n19505), .B2(n19504), .ZN(n19515) );
  AND3_X1 U22689 ( .A1(n19508), .A2(n19507), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19511) );
  AOI221_X1 U22690 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C1(n19663), .C2(n13161), .A(
        n19509), .ZN(n19510) );
  AOI211_X1 U22691 ( .C1(n19512), .C2(n19657), .A(n19511), .B(n19510), .ZN(
        n19660) );
  INV_X1 U22692 ( .A(n19516), .ZN(n19521) );
  NAND2_X1 U22693 ( .A1(n19518), .A2(n19517), .ZN(n19520) );
  AOI21_X1 U22694 ( .B1(n19521), .B2(n19520), .A(n19519), .ZN(n19536) );
  AOI22_X1 U22695 ( .A1(n19525), .A2(n19524), .B1(n19523), .B2(n19522), .ZN(
        n19526) );
  OAI221_X1 U22696 ( .B1(n19529), .B2(n19528), .C1(n19529), .C2(n19527), .A(
        n19526), .ZN(n19689) );
  AOI221_X1 U22697 ( .B1(P3_MORE_REG_SCAN_IN), .B2(n19531), .C1(
        P3_FLUSH_REG_SCAN_IN), .C2(n19531), .A(n19530), .ZN(n19532) );
  OAI211_X1 U22698 ( .C1(n21439), .C2(n19534), .A(n19533), .B(n19532), .ZN(
        n19535) );
  AOI22_X1 U22699 ( .A1(n19671), .A2(n19537), .B1(n19693), .B2(n18300), .ZN(
        n19538) );
  INV_X1 U22700 ( .A(n19538), .ZN(n19544) );
  INV_X1 U22701 ( .A(n19539), .ZN(n19541) );
  OAI211_X1 U22702 ( .C1(n19541), .C2(n19540), .A(n19700), .B(n19548), .ZN(
        n19649) );
  OAI21_X1 U22703 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19702), .A(n19649), 
        .ZN(n19549) );
  NOR2_X1 U22704 ( .A1(n19542), .A2(n19549), .ZN(n19543) );
  MUX2_X1 U22705 ( .A(n19544), .B(n19543), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n19546) );
  OAI211_X1 U22706 ( .C1(n19548), .C2(n19547), .A(n19546), .B(n19545), .ZN(
        P3_U2996) );
  NAND2_X1 U22707 ( .A1(n19693), .A2(n18300), .ZN(n19554) );
  NAND4_X1 U22708 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n19693), .A4(n19692), .ZN(n19556) );
  INV_X1 U22709 ( .A(n19549), .ZN(n19551) );
  NAND3_X1 U22710 ( .A1(n19552), .A2(n19551), .A3(n19550), .ZN(n19553) );
  NAND4_X1 U22711 ( .A1(n19555), .A2(n19554), .A3(n19556), .A4(n19553), .ZN(
        P3_U2997) );
  AND4_X1 U22712 ( .A1(n19695), .A2(n19557), .A3(n19556), .A4(n19648), .ZN(
        P3_U2998) );
  AND2_X1 U22713 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19559), .ZN(
        P3_U2999) );
  AND2_X1 U22714 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19559), .ZN(
        P3_U3000) );
  AND2_X1 U22715 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19559), .ZN(
        P3_U3001) );
  AND2_X1 U22716 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19559), .ZN(
        P3_U3002) );
  AND2_X1 U22717 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19559), .ZN(
        P3_U3003) );
  AND2_X1 U22718 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19559), .ZN(
        P3_U3004) );
  AND2_X1 U22719 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19559), .ZN(
        P3_U3005) );
  AND2_X1 U22720 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19559), .ZN(
        P3_U3006) );
  AND2_X1 U22721 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19559), .ZN(
        P3_U3007) );
  AND2_X1 U22722 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19559), .ZN(
        P3_U3008) );
  AND2_X1 U22723 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19559), .ZN(
        P3_U3009) );
  AND2_X1 U22724 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19559), .ZN(
        P3_U3010) );
  AND2_X1 U22725 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19559), .ZN(
        P3_U3011) );
  AND2_X1 U22726 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19559), .ZN(
        P3_U3012) );
  AND2_X1 U22727 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19559), .ZN(
        P3_U3013) );
  AND2_X1 U22728 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19558), .ZN(
        P3_U3014) );
  INV_X1 U22729 ( .A(P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n21351) );
  NOR2_X1 U22730 ( .A1(n21351), .A2(n19647), .ZN(P3_U3015) );
  AND2_X1 U22731 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19558), .ZN(
        P3_U3016) );
  AND2_X1 U22732 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19558), .ZN(
        P3_U3017) );
  AND2_X1 U22733 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19558), .ZN(
        P3_U3018) );
  AND2_X1 U22734 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19558), .ZN(
        P3_U3019) );
  INV_X1 U22735 ( .A(P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n21355) );
  NOR2_X1 U22736 ( .A1(n21355), .A2(n19647), .ZN(P3_U3020) );
  AND2_X1 U22737 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19558), .ZN(P3_U3021) );
  AND2_X1 U22738 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19558), .ZN(P3_U3022) );
  AND2_X1 U22739 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19559), .ZN(P3_U3023) );
  AND2_X1 U22740 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19559), .ZN(P3_U3024) );
  AND2_X1 U22741 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19559), .ZN(P3_U3025) );
  AND2_X1 U22742 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19559), .ZN(P3_U3026) );
  AND2_X1 U22743 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19559), .ZN(P3_U3027) );
  AND2_X1 U22744 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19559), .ZN(P3_U3028) );
  INV_X1 U22745 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19563) );
  AOI21_X1 U22746 ( .B1(HOLD), .B2(n19560), .A(n19563), .ZN(n19562) );
  AOI21_X1 U22747 ( .B1(n19693), .B2(P3_STATE_REG_1__SCAN_IN), .A(n19572), 
        .ZN(n19574) );
  AOI21_X1 U22748 ( .B1(NA), .B2(n19561), .A(n19575), .ZN(n19567) );
  OAI22_X1 U22749 ( .A1(n19707), .A2(n19562), .B1(n19574), .B2(n19567), .ZN(
        P3_U3029) );
  NOR2_X1 U22750 ( .A1(n19575), .A2(n20556), .ZN(n19570) );
  NOR3_X1 U22751 ( .A1(n19570), .A2(n19572), .A3(n19563), .ZN(n19564) );
  NOR2_X1 U22752 ( .A1(n19564), .A2(n19690), .ZN(n19565) );
  NAND2_X1 U22753 ( .A1(n19693), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19568) );
  OAI211_X1 U22754 ( .C1(n20556), .C2(n19566), .A(n19565), .B(n19568), .ZN(
        P3_U3030) );
  INV_X1 U22755 ( .A(n19567), .ZN(n19573) );
  OAI22_X1 U22756 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19568), .ZN(n19569) );
  OAI22_X1 U22757 ( .A1(n19570), .A2(n19569), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19571) );
  OAI22_X1 U22758 ( .A1(n19574), .A2(n19573), .B1(n19572), .B2(n19571), .ZN(
        P3_U3031) );
  INV_X1 U22759 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19577) );
  NAND2_X1 U22760 ( .A1(n19707), .A2(n19575), .ZN(n19621) );
  CLKBUF_X1 U22761 ( .A(n19621), .Z(n19634) );
  OAI222_X1 U22762 ( .A1(n19678), .A2(n19630), .B1(n19576), .B2(n19707), .C1(
        n19577), .C2(n19634), .ZN(P3_U3032) );
  OAI222_X1 U22763 ( .A1(n19634), .A2(n19579), .B1(n19578), .B2(n19707), .C1(
        n19577), .C2(n19630), .ZN(P3_U3033) );
  OAI222_X1 U22764 ( .A1(n19621), .A2(n19581), .B1(n19580), .B2(n19707), .C1(
        n19579), .C2(n19630), .ZN(P3_U3034) );
  OAI222_X1 U22765 ( .A1(n19621), .A2(n19584), .B1(n19582), .B2(n19707), .C1(
        n19581), .C2(n19630), .ZN(P3_U3035) );
  OAI222_X1 U22766 ( .A1(n19584), .A2(n19630), .B1(n19583), .B2(n19707), .C1(
        n19585), .C2(n19634), .ZN(P3_U3036) );
  OAI222_X1 U22767 ( .A1(n19621), .A2(n19587), .B1(n19586), .B2(n19707), .C1(
        n19585), .C2(n19630), .ZN(P3_U3037) );
  OAI222_X1 U22768 ( .A1(n19621), .A2(n19589), .B1(n19588), .B2(n19707), .C1(
        n19587), .C2(n19630), .ZN(P3_U3038) );
  OAI222_X1 U22769 ( .A1(n19621), .A2(n19591), .B1(n19590), .B2(n19707), .C1(
        n19589), .C2(n19630), .ZN(P3_U3039) );
  OAI222_X1 U22770 ( .A1(n19621), .A2(n19593), .B1(n19592), .B2(n19707), .C1(
        n19591), .C2(n19630), .ZN(P3_U3040) );
  OAI222_X1 U22771 ( .A1(n19634), .A2(n19595), .B1(n19594), .B2(n19707), .C1(
        n19593), .C2(n19630), .ZN(P3_U3041) );
  OAI222_X1 U22772 ( .A1(n19634), .A2(n19597), .B1(n19596), .B2(n19707), .C1(
        n19595), .C2(n19630), .ZN(P3_U3042) );
  INV_X1 U22773 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19599) );
  OAI222_X1 U22774 ( .A1(n19634), .A2(n19599), .B1(n19598), .B2(n19707), .C1(
        n19597), .C2(n19630), .ZN(P3_U3043) );
  OAI222_X1 U22775 ( .A1(n19634), .A2(n19602), .B1(n19600), .B2(n19707), .C1(
        n19599), .C2(n19630), .ZN(P3_U3044) );
  OAI222_X1 U22776 ( .A1(n19602), .A2(n19630), .B1(n19601), .B2(n19707), .C1(
        n19603), .C2(n19634), .ZN(P3_U3045) );
  INV_X1 U22777 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19605) );
  OAI222_X1 U22778 ( .A1(n19634), .A2(n19605), .B1(n19604), .B2(n19707), .C1(
        n19603), .C2(n19630), .ZN(P3_U3046) );
  OAI222_X1 U22779 ( .A1(n19634), .A2(n19607), .B1(n19606), .B2(n19707), .C1(
        n19605), .C2(n19630), .ZN(P3_U3047) );
  OAI222_X1 U22780 ( .A1(n19621), .A2(n19609), .B1(n19608), .B2(n19707), .C1(
        n19607), .C2(n19630), .ZN(P3_U3048) );
  OAI222_X1 U22781 ( .A1(n19621), .A2(n19611), .B1(n19610), .B2(n19707), .C1(
        n19609), .C2(n19630), .ZN(P3_U3049) );
  OAI222_X1 U22782 ( .A1(n19621), .A2(n19614), .B1(n19612), .B2(n19707), .C1(
        n19611), .C2(n19630), .ZN(P3_U3050) );
  OAI222_X1 U22783 ( .A1(n19614), .A2(n19630), .B1(n19613), .B2(n19707), .C1(
        n19615), .C2(n19634), .ZN(P3_U3051) );
  OAI222_X1 U22784 ( .A1(n19621), .A2(n19617), .B1(n19616), .B2(n19707), .C1(
        n19615), .C2(n19630), .ZN(P3_U3052) );
  OAI222_X1 U22785 ( .A1(n19621), .A2(n19619), .B1(n19618), .B2(n19707), .C1(
        n19617), .C2(n19630), .ZN(P3_U3053) );
  OAI222_X1 U22786 ( .A1(n19621), .A2(n19623), .B1(n19620), .B2(n19707), .C1(
        n19619), .C2(n19630), .ZN(P3_U3054) );
  OAI222_X1 U22787 ( .A1(n19623), .A2(n19630), .B1(n19622), .B2(n19707), .C1(
        n19624), .C2(n19634), .ZN(P3_U3055) );
  OAI222_X1 U22788 ( .A1(n19634), .A2(n21372), .B1(n19625), .B2(n19707), .C1(
        n19624), .C2(n19630), .ZN(P3_U3056) );
  OAI222_X1 U22789 ( .A1(n19634), .A2(n19627), .B1(n19626), .B2(n19707), .C1(
        n21372), .C2(n19630), .ZN(P3_U3057) );
  INV_X1 U22790 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19631) );
  OAI222_X1 U22791 ( .A1(n19634), .A2(n19631), .B1(n19628), .B2(n19707), .C1(
        n19627), .C2(n19630), .ZN(P3_U3058) );
  OAI222_X1 U22792 ( .A1(n19631), .A2(n19630), .B1(n19629), .B2(n19707), .C1(
        n19632), .C2(n19634), .ZN(P3_U3059) );
  OAI222_X1 U22793 ( .A1(n19634), .A2(n19637), .B1(n19633), .B2(n19707), .C1(
        n19632), .C2(n19630), .ZN(P3_U3060) );
  OAI222_X1 U22794 ( .A1(n19630), .A2(n19637), .B1(n19636), .B2(n19707), .C1(
        n19635), .C2(n19634), .ZN(P3_U3061) );
  INV_X1 U22795 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n19638) );
  AOI22_X1 U22796 ( .A1(n19707), .A2(n19639), .B1(n19638), .B2(n19705), .ZN(
        P3_U3274) );
  INV_X1 U22797 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19680) );
  INV_X1 U22798 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n19640) );
  AOI22_X1 U22799 ( .A1(n19707), .A2(n19680), .B1(n19640), .B2(n19705), .ZN(
        P3_U3275) );
  INV_X1 U22800 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n19641) );
  AOI22_X1 U22801 ( .A1(n19707), .A2(n19642), .B1(n19641), .B2(n19705), .ZN(
        P3_U3276) );
  INV_X1 U22802 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19686) );
  INV_X1 U22803 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n19643) );
  AOI22_X1 U22804 ( .A1(n19707), .A2(n19686), .B1(n19643), .B2(n19705), .ZN(
        P3_U3277) );
  OAI21_X1 U22805 ( .B1(n19647), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19645), 
        .ZN(n19644) );
  INV_X1 U22806 ( .A(n19644), .ZN(P3_U3280) );
  OAI21_X1 U22807 ( .B1(n19647), .B2(n19646), .A(n19645), .ZN(P3_U3281) );
  OAI221_X1 U22808 ( .B1(n19650), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19650), 
        .C2(n19649), .A(n19648), .ZN(P3_U3282) );
  AOI22_X1 U22809 ( .A1(n19673), .A2(n19652), .B1(n19671), .B2(n19651), .ZN(
        n19653) );
  AOI22_X1 U22810 ( .A1(n19677), .A2(n19654), .B1(n19653), .B2(n19675), .ZN(
        P3_U3285) );
  AOI22_X1 U22811 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n19655), .B2(n13072), .ZN(
        n19665) );
  NOR2_X1 U22812 ( .A1(n19656), .A2(n19674), .ZN(n19666) );
  OAI22_X1 U22813 ( .A1(n19660), .A2(n19659), .B1(n19658), .B2(n19657), .ZN(
        n19661) );
  AOI21_X1 U22814 ( .B1(n19665), .B2(n19666), .A(n19661), .ZN(n19662) );
  AOI22_X1 U22815 ( .A1(n19677), .A2(n19663), .B1(n19662), .B2(n19675), .ZN(
        P3_U3288) );
  INV_X1 U22816 ( .A(n19664), .ZN(n19668) );
  INV_X1 U22817 ( .A(n19665), .ZN(n19667) );
  AOI222_X1 U22818 ( .A1(n19669), .A2(n19673), .B1(n19671), .B2(n19668), .C1(
        n19667), .C2(n19666), .ZN(n19670) );
  AOI22_X1 U22819 ( .A1(n19677), .A2(n13161), .B1(n19670), .B2(n19675), .ZN(
        P3_U3289) );
  AOI222_X1 U22820 ( .A1(n19674), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19673), 
        .B2(n19672), .C1(n13162), .C2(n19671), .ZN(n19676) );
  AOI22_X1 U22821 ( .A1(n19677), .A2(n13162), .B1(n19676), .B2(n19675), .ZN(
        P3_U3290) );
  AOI21_X1 U22822 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19679) );
  AOI22_X1 U22823 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19679), .B2(n19678), .ZN(n19681) );
  AOI22_X1 U22824 ( .A1(n19682), .A2(n19681), .B1(n19680), .B2(n19685), .ZN(
        P3_U3292) );
  NOR2_X1 U22825 ( .A1(n19685), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19683) );
  AOI22_X1 U22826 ( .A1(n19686), .A2(n19685), .B1(n19684), .B2(n19683), .ZN(
        P3_U3293) );
  INV_X1 U22827 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19687) );
  AOI22_X1 U22828 ( .A1(n19707), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19687), 
        .B2(n19705), .ZN(P3_U3294) );
  MUX2_X1 U22829 ( .A(P3_MORE_REG_SCAN_IN), .B(n19689), .S(n19688), .Z(
        P3_U3295) );
  OAI21_X1 U22830 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n19691), .A(n19690), 
        .ZN(n19694) );
  AOI211_X1 U22831 ( .C1(n19711), .C2(n19694), .A(n19693), .B(n19692), .ZN(
        n19697) );
  OAI21_X1 U22832 ( .B1(n19697), .B2(n19696), .A(n19695), .ZN(n19704) );
  OAI21_X1 U22833 ( .B1(n19700), .B2(n19699), .A(n19698), .ZN(n19701) );
  AOI21_X1 U22834 ( .B1(n18300), .B2(n19702), .A(n19701), .ZN(n19703) );
  MUX2_X1 U22835 ( .A(n19704), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n19703), 
        .Z(P3_U3296) );
  INV_X1 U22836 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19713) );
  INV_X1 U22837 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n19706) );
  AOI22_X1 U22838 ( .A1(n19707), .A2(n19713), .B1(n19706), .B2(n19705), .ZN(
        P3_U3297) );
  NOR2_X1 U22839 ( .A1(n19708), .A2(n19710), .ZN(n19714) );
  INV_X1 U22840 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n19709) );
  AOI22_X1 U22841 ( .A1(n19711), .A2(n19710), .B1(n19714), .B2(n19709), .ZN(
        P3_U3298) );
  AOI21_X1 U22842 ( .B1(n19714), .B2(n19713), .A(n19712), .ZN(P3_U3299) );
  AOI211_X1 U22843 ( .C1(n19716), .C2(P2_MEMORYFETCH_REG_SCAN_IN), .A(n19719), 
        .B(n19715), .ZN(n19717) );
  INV_X1 U22844 ( .A(n19717), .ZN(P2_U2814) );
  INV_X1 U22845 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n19718) );
  INV_X1 U22846 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20565) );
  NAND2_X1 U22847 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20565), .ZN(n20555) );
  INV_X1 U22848 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n21404) );
  NAND2_X1 U22849 ( .A1(n20562), .A2(n21404), .ZN(n20552) );
  OAI21_X1 U22850 ( .B1(n20562), .B2(n20555), .A(n20552), .ZN(n20627) );
  OAI21_X1 U22851 ( .B1(n20562), .B2(n19718), .A(n20546), .ZN(P2_U2815) );
  AOI22_X1 U22852 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19719), .B1(n20682), 
        .B2(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19720) );
  INV_X1 U22853 ( .A(n19720), .ZN(P2_U2816) );
  OAI21_X1 U22854 ( .B1(n21404), .B2(P2_CODEFETCH_REG_SCAN_IN), .A(n20547), 
        .ZN(n19721) );
  AOI22_X1 U22855 ( .A1(n20700), .A2(P2_D_C_N_REG_SCAN_IN), .B1(n20562), .B2(
        n19721), .ZN(n19722) );
  INV_X1 U22856 ( .A(n19722), .ZN(P2_U2817) );
  OAI21_X1 U22857 ( .B1(n20559), .B2(BS16), .A(n20627), .ZN(n20625) );
  OAI21_X1 U22858 ( .B1(n20627), .B2(n20687), .A(n20625), .ZN(P2_U2818) );
  NOR2_X1 U22859 ( .A1(n19724), .A2(n19723), .ZN(n20679) );
  OAI21_X1 U22860 ( .B1(n20679), .B2(n11140), .A(n19725), .ZN(P2_U2819) );
  NOR4_X1 U22861 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A3(P2_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n19735) );
  NOR4_X1 U22862 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n19734) );
  NOR4_X1 U22863 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(P2_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n19726) );
  INV_X1 U22864 ( .A(P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n21336) );
  INV_X1 U22865 ( .A(P2_DATAWIDTH_REG_28__SCAN_IN), .ZN(n21455) );
  NAND3_X1 U22866 ( .A1(n19726), .A2(n21336), .A3(n21455), .ZN(n19732) );
  NOR4_X1 U22867 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_19__SCAN_IN), .A3(P2_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_21__SCAN_IN), .ZN(n19730) );
  NOR4_X1 U22868 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_15__SCAN_IN), .A3(P2_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_17__SCAN_IN), .ZN(n19729) );
  NOR4_X1 U22869 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_27__SCAN_IN), .A3(P2_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19728) );
  NOR4_X1 U22870 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_23__SCAN_IN), .A3(P2_DATAWIDTH_REG_24__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_25__SCAN_IN), .ZN(n19727) );
  NAND4_X1 U22871 ( .A1(n19730), .A2(n19729), .A3(n19728), .A4(n19727), .ZN(
        n19731) );
  AOI211_X1 U22872 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19732), .B(n19731), .ZN(n19733) );
  NAND3_X1 U22873 ( .A1(n19735), .A2(n19734), .A3(n19733), .ZN(n19736) );
  NOR2_X1 U22874 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19736), .ZN(n19738) );
  INV_X1 U22875 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20623) );
  AOI22_X1 U22876 ( .A1(n19738), .A2(n19739), .B1(n19736), .B2(n20623), .ZN(
        P2_U2820) );
  INV_X1 U22877 ( .A(n19736), .ZN(n19744) );
  NOR2_X1 U22878 ( .A1(n19744), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19737)
         );
  OR4_X1 U22879 ( .A1(n19736), .A2(P2_REIP_REG_0__SCAN_IN), .A3(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A4(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19743) );
  OAI21_X1 U22880 ( .B1(n19738), .B2(n19737), .A(n19743), .ZN(P2_U2821) );
  INV_X1 U22881 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20626) );
  NAND2_X1 U22882 ( .A1(n19738), .A2(n20626), .ZN(n19742) );
  OAI21_X1 U22883 ( .B1(n19739), .B2(n20567), .A(n19744), .ZN(n19740) );
  OAI21_X1 U22884 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19744), .A(n19740), 
        .ZN(n19741) );
  OAI221_X1 U22885 ( .B1(n19742), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19742), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19741), .ZN(P2_U2822) );
  INV_X1 U22886 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20620) );
  OAI211_X1 U22887 ( .C1(n19744), .C2(n20620), .A(n19743), .B(n19742), .ZN(
        P2_U2823) );
  NAND2_X1 U22888 ( .A1(n19866), .A2(n19745), .ZN(n19759) );
  OAI21_X1 U22889 ( .B1(n10245), .B2(n19760), .A(n19759), .ZN(n19746) );
  XNOR2_X1 U22890 ( .A(n19747), .B(n19746), .ZN(n19758) );
  NAND2_X1 U22891 ( .A1(n19856), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n19749) );
  AOI21_X1 U22892 ( .B1(n19834), .B2(P2_REIP_REG_19__SCAN_IN), .A(n19941), 
        .ZN(n19748) );
  OAI211_X1 U22893 ( .C1(n19838), .C2(n19750), .A(n19749), .B(n19748), .ZN(
        n19751) );
  AOI21_X1 U22894 ( .B1(n19752), .B2(n19832), .A(n19751), .ZN(n19757) );
  OAI22_X1 U22895 ( .A1(n19754), .A2(n19871), .B1(n19753), .B2(n19870), .ZN(
        n19755) );
  INV_X1 U22896 ( .A(n19755), .ZN(n19756) );
  OAI211_X1 U22897 ( .C1(n20545), .C2(n19758), .A(n19757), .B(n19756), .ZN(
        P2_U2836) );
  XNOR2_X1 U22898 ( .A(n19760), .B(n19759), .ZN(n19772) );
  AOI21_X1 U22899 ( .B1(n19834), .B2(P2_REIP_REG_18__SCAN_IN), .A(n19941), 
        .ZN(n19761) );
  OAI21_X1 U22900 ( .B1(n19762), .B2(n19838), .A(n19761), .ZN(n19765) );
  NOR2_X1 U22901 ( .A1(n19763), .A2(n19860), .ZN(n19764) );
  AOI211_X1 U22902 ( .C1(n19856), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n19765), .B(n19764), .ZN(n19771) );
  NOR2_X1 U22903 ( .A1(n19766), .A2(n19870), .ZN(n19767) );
  AOI21_X1 U22904 ( .B1(n19769), .B2(n19768), .A(n19767), .ZN(n19770) );
  OAI211_X1 U22905 ( .C1(n20545), .C2(n19772), .A(n19771), .B(n19770), .ZN(
        P2_U2837) );
  NAND2_X1 U22906 ( .A1(n19866), .A2(n19773), .ZN(n19774) );
  XNOR2_X1 U22907 ( .A(n19775), .B(n19774), .ZN(n19786) );
  INV_X1 U22908 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n19778) );
  OAI21_X1 U22909 ( .B1(n19859), .B2(n20591), .A(n16491), .ZN(n19776) );
  AOI21_X1 U22910 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n19864), .A(n19776), .ZN(
        n19777) );
  OAI21_X1 U22911 ( .B1(n19778), .B2(n19878), .A(n19777), .ZN(n19779) );
  AOI21_X1 U22912 ( .B1(n19780), .B2(n19832), .A(n19779), .ZN(n19785) );
  OAI22_X1 U22913 ( .A1(n19782), .A2(n19871), .B1(n19781), .B2(n19870), .ZN(
        n19783) );
  INV_X1 U22914 ( .A(n19783), .ZN(n19784) );
  OAI211_X1 U22915 ( .C1(n20545), .C2(n19786), .A(n19785), .B(n19784), .ZN(
        P2_U2839) );
  NOR2_X1 U22916 ( .A1(n10245), .A2(n19787), .ZN(n19788) );
  XNOR2_X1 U22917 ( .A(n19789), .B(n19788), .ZN(n19799) );
  NAND2_X1 U22918 ( .A1(n19790), .A2(n19832), .ZN(n19792) );
  AOI21_X1 U22919 ( .B1(n19864), .B2(P2_EBX_REG_15__SCAN_IN), .A(n19941), .ZN(
        n19791) );
  OAI211_X1 U22920 ( .C1(n19878), .C2(n19793), .A(n19792), .B(n19791), .ZN(
        n19797) );
  OAI22_X1 U22921 ( .A1(n19795), .A2(n19871), .B1(n19794), .B2(n19870), .ZN(
        n19796) );
  AOI211_X1 U22922 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n19834), .A(n19797), 
        .B(n19796), .ZN(n19798) );
  OAI21_X1 U22923 ( .B1(n20545), .B2(n19799), .A(n19798), .ZN(P2_U2840) );
  AOI21_X1 U22924 ( .B1(n19834), .B2(P2_REIP_REG_11__SCAN_IN), .A(n19941), 
        .ZN(n19800) );
  OAI21_X1 U22925 ( .B1(n19801), .B2(n19838), .A(n19800), .ZN(n19802) );
  AOI21_X1 U22926 ( .B1(n19804), .B2(n19803), .A(n19802), .ZN(n19815) );
  AOI22_X1 U22927 ( .A1(n19805), .A2(n19832), .B1(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19856), .ZN(n19814) );
  OAI22_X1 U22928 ( .A1(n19807), .A2(n19871), .B1(n19806), .B2(n19811), .ZN(
        n19808) );
  INV_X1 U22929 ( .A(n19808), .ZN(n19813) );
  OAI211_X1 U22930 ( .C1(n9750), .C2(n19811), .A(n19810), .B(n19809), .ZN(
        n19812) );
  NAND4_X1 U22931 ( .A1(n19815), .A2(n19814), .A3(n19813), .A4(n19812), .ZN(
        P2_U2844) );
  AOI21_X1 U22932 ( .B1(n19834), .B2(P2_REIP_REG_10__SCAN_IN), .A(n19941), 
        .ZN(n19816) );
  OAI21_X1 U22933 ( .B1(n19817), .B2(n19838), .A(n19816), .ZN(n19818) );
  AOI21_X1 U22934 ( .B1(n19819), .B2(n19832), .A(n19818), .ZN(n19828) );
  NAND2_X1 U22935 ( .A1(n19866), .A2(n19820), .ZN(n19821) );
  XNOR2_X1 U22936 ( .A(n19822), .B(n19821), .ZN(n19826) );
  OAI22_X1 U22937 ( .A1(n19871), .A2(n19824), .B1(n19823), .B2(n19870), .ZN(
        n19825) );
  AOI21_X1 U22938 ( .B1(n19875), .B2(n19826), .A(n19825), .ZN(n19827) );
  OAI211_X1 U22939 ( .C1(n10404), .C2(n19878), .A(n19828), .B(n19827), .ZN(
        P2_U2845) );
  NOR2_X1 U22940 ( .A1(n10245), .A2(n19829), .ZN(n19831) );
  XNOR2_X1 U22941 ( .A(n19831), .B(n19830), .ZN(n19844) );
  NAND2_X1 U22942 ( .A1(n19833), .A2(n19832), .ZN(n19836) );
  AOI21_X1 U22943 ( .B1(n19834), .B2(P2_REIP_REG_9__SCAN_IN), .A(n19941), .ZN(
        n19835) );
  OAI211_X1 U22944 ( .C1(n19838), .C2(n19837), .A(n19836), .B(n19835), .ZN(
        n19842) );
  OAI22_X1 U22945 ( .A1(n19840), .A2(n19871), .B1(n19839), .B2(n19870), .ZN(
        n19841) );
  AOI211_X1 U22946 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19856), .A(
        n19842), .B(n19841), .ZN(n19843) );
  OAI21_X1 U22947 ( .B1(n20545), .B2(n19844), .A(n19843), .ZN(P2_U2846) );
  NOR2_X1 U22948 ( .A1(n10245), .A2(n19845), .ZN(n19847) );
  XOR2_X1 U22949 ( .A(n19848), .B(n19847), .Z(n19858) );
  OAI21_X1 U22950 ( .B1(n19859), .B2(n20576), .A(n16491), .ZN(n19849) );
  AOI21_X1 U22951 ( .B1(P2_EBX_REG_7__SCAN_IN), .B2(n19864), .A(n19849), .ZN(
        n19850) );
  OAI21_X1 U22952 ( .B1(n19851), .B2(n19860), .A(n19850), .ZN(n19855) );
  OAI22_X1 U22953 ( .A1(n19853), .A2(n19871), .B1(n19870), .B2(n19852), .ZN(
        n19854) );
  AOI211_X1 U22954 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19856), .A(
        n19855), .B(n19854), .ZN(n19857) );
  OAI21_X1 U22955 ( .B1(n20545), .B2(n19858), .A(n19857), .ZN(P2_U2848) );
  OAI21_X1 U22956 ( .B1(n19859), .B2(n20574), .A(n16491), .ZN(n19863) );
  NOR2_X1 U22957 ( .A1(n19861), .A2(n19860), .ZN(n19862) );
  AOI211_X1 U22958 ( .C1(n19864), .C2(P2_EBX_REG_6__SCAN_IN), .A(n19863), .B(
        n19862), .ZN(n19877) );
  NAND2_X1 U22959 ( .A1(n19866), .A2(n19865), .ZN(n19867) );
  XNOR2_X1 U22960 ( .A(n19868), .B(n19867), .ZN(n19874) );
  OAI22_X1 U22961 ( .A1(n19872), .A2(n19871), .B1(n19870), .B2(n19869), .ZN(
        n19873) );
  AOI21_X1 U22962 ( .B1(n19875), .B2(n19874), .A(n19873), .ZN(n19876) );
  OAI211_X1 U22963 ( .C1(n19879), .C2(n19878), .A(n19877), .B(n19876), .ZN(
        P2_U2849) );
  AOI22_X1 U22964 ( .A1(n20635), .A2(n19888), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19887), .ZN(n19885) );
  OAI21_X1 U22965 ( .B1(n19882), .B2(n19881), .A(n19880), .ZN(n19883) );
  NAND2_X1 U22966 ( .A1(n19883), .A2(n19892), .ZN(n19884) );
  OAI211_X1 U22967 ( .C1(n19886), .C2(n19896), .A(n19885), .B(n19884), .ZN(
        P2_U2916) );
  AOI22_X1 U22968 ( .A1(n19888), .A2(n20653), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19887), .ZN(n19895) );
  OAI21_X1 U22969 ( .B1(n19891), .B2(n19890), .A(n19889), .ZN(n19893) );
  NAND2_X1 U22970 ( .A1(n19893), .A2(n19892), .ZN(n19894) );
  OAI211_X1 U22971 ( .C1(n19897), .C2(n19896), .A(n19895), .B(n19894), .ZN(
        P2_U2918) );
  NOR2_X1 U22972 ( .A1(n19902), .A2(n19898), .ZN(P2_U2920) );
  AOI22_X1 U22973 ( .A1(n19899), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n20685), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19900) );
  OAI21_X1 U22974 ( .B1(n19902), .B2(n19901), .A(n19900), .ZN(P2_U2921) );
  AOI22_X1 U22975 ( .A1(n19931), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n20685), 
        .B2(P2_LWORD_REG_15__SCAN_IN), .ZN(n19903) );
  OAI21_X1 U22976 ( .B1(n13398), .B2(n19933), .A(n19903), .ZN(P2_U2936) );
  INV_X1 U22977 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19905) );
  AOI22_X1 U22978 ( .A1(n19931), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n20685), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19904) );
  OAI21_X1 U22979 ( .B1(n19905), .B2(n19933), .A(n19904), .ZN(P2_U2937) );
  AOI22_X1 U22980 ( .A1(n19931), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n20685), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n19906) );
  OAI21_X1 U22981 ( .B1(n19907), .B2(n19933), .A(n19906), .ZN(P2_U2938) );
  AOI22_X1 U22982 ( .A1(n19931), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n20685), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n19908) );
  OAI21_X1 U22983 ( .B1(n19909), .B2(n19933), .A(n19908), .ZN(P2_U2939) );
  AOI22_X1 U22984 ( .A1(n19931), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n20685), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n19910) );
  OAI21_X1 U22985 ( .B1(n19911), .B2(n19933), .A(n19910), .ZN(P2_U2940) );
  AOI22_X1 U22986 ( .A1(n19931), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n20685), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n19912) );
  OAI21_X1 U22987 ( .B1(n19913), .B2(n19933), .A(n19912), .ZN(P2_U2941) );
  AOI22_X1 U22988 ( .A1(n19931), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n20685), 
        .B2(P2_LWORD_REG_9__SCAN_IN), .ZN(n19914) );
  OAI21_X1 U22989 ( .B1(n19915), .B2(n19933), .A(n19914), .ZN(P2_U2942) );
  AOI22_X1 U22990 ( .A1(n19931), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n20685), 
        .B2(P2_LWORD_REG_8__SCAN_IN), .ZN(n19916) );
  OAI21_X1 U22991 ( .B1(n19917), .B2(n19933), .A(n19916), .ZN(P2_U2943) );
  AOI22_X1 U22992 ( .A1(n19931), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n20685), 
        .B2(P2_LWORD_REG_7__SCAN_IN), .ZN(n19918) );
  OAI21_X1 U22993 ( .B1(n19919), .B2(n19933), .A(n19918), .ZN(P2_U2944) );
  AOI22_X1 U22994 ( .A1(n19931), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n20685), 
        .B2(P2_LWORD_REG_6__SCAN_IN), .ZN(n19920) );
  OAI21_X1 U22995 ( .B1(n19921), .B2(n19933), .A(n19920), .ZN(P2_U2945) );
  AOI22_X1 U22996 ( .A1(n19931), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n20685), 
        .B2(P2_LWORD_REG_5__SCAN_IN), .ZN(n19922) );
  OAI21_X1 U22997 ( .B1(n19923), .B2(n19933), .A(n19922), .ZN(P2_U2946) );
  INV_X1 U22998 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19925) );
  AOI22_X1 U22999 ( .A1(n19931), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n20685), 
        .B2(P2_LWORD_REG_4__SCAN_IN), .ZN(n19924) );
  OAI21_X1 U23000 ( .B1(n19925), .B2(n19933), .A(n19924), .ZN(P2_U2947) );
  INV_X1 U23001 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19927) );
  AOI22_X1 U23002 ( .A1(n19931), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n20685), 
        .B2(P2_LWORD_REG_3__SCAN_IN), .ZN(n19926) );
  OAI21_X1 U23003 ( .B1(n19927), .B2(n19933), .A(n19926), .ZN(P2_U2948) );
  AOI22_X1 U23004 ( .A1(n19931), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n20685), 
        .B2(P2_LWORD_REG_2__SCAN_IN), .ZN(n19928) );
  OAI21_X1 U23005 ( .B1(n21413), .B2(n19933), .A(n19928), .ZN(P2_U2949) );
  INV_X1 U23006 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19930) );
  AOI22_X1 U23007 ( .A1(n19931), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n20685), 
        .B2(P2_LWORD_REG_1__SCAN_IN), .ZN(n19929) );
  OAI21_X1 U23008 ( .B1(n19930), .B2(n19933), .A(n19929), .ZN(P2_U2950) );
  AOI22_X1 U23009 ( .A1(n19931), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(n20685), 
        .B2(P2_LWORD_REG_0__SCAN_IN), .ZN(n19932) );
  OAI21_X1 U23010 ( .B1(n11282), .B2(n19933), .A(n19932), .ZN(P2_U2951) );
  AOI22_X1 U23011 ( .A1(n19938), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n19937), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19936) );
  NAND2_X1 U23012 ( .A1(n19935), .A2(n19934), .ZN(n19939) );
  NAND2_X1 U23013 ( .A1(n19936), .A2(n19939), .ZN(P2_U2966) );
  AOI22_X1 U23014 ( .A1(n19938), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n19937), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19940) );
  NAND2_X1 U23015 ( .A1(n19940), .A2(n19939), .ZN(P2_U2981) );
  AOI22_X1 U23016 ( .A1(n19943), .A2(n19942), .B1(P2_REIP_REG_4__SCAN_IN), 
        .B2(n19941), .ZN(n19953) );
  NAND2_X1 U23017 ( .A1(n19944), .A2(n10145), .ZN(n19948) );
  NAND2_X1 U23018 ( .A1(n19946), .A2(n19945), .ZN(n19947) );
  OAI211_X1 U23019 ( .C1(n19950), .C2(n19949), .A(n19948), .B(n19947), .ZN(
        n19951) );
  INV_X1 U23020 ( .A(n19951), .ZN(n19952) );
  OAI211_X1 U23021 ( .C1(n19955), .C2(n19954), .A(n19953), .B(n19952), .ZN(
        P2_U3010) );
  AOI22_X1 U23022 ( .A1(n19958), .A2(n19957), .B1(n19956), .B2(n20653), .ZN(
        n19959) );
  OAI21_X1 U23023 ( .B1(n19963), .B2(n19960), .A(n19959), .ZN(n19966) );
  AOI211_X1 U23024 ( .C1(n19964), .C2(n19963), .A(n19962), .B(n19961), .ZN(
        n19965) );
  AOI211_X1 U23025 ( .C1(n19967), .C2(n9927), .A(n19966), .B(n19965), .ZN(
        n19969) );
  OAI211_X1 U23026 ( .C1(n19971), .C2(n19970), .A(n19969), .B(n19968), .ZN(
        P2_U3045) );
  AOI22_X1 U23027 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20002), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n20001), .ZN(n20489) );
  AOI22_X1 U23028 ( .A1(n10554), .A2(n20423), .B1(n19999), .B2(n20422), .ZN(
        n19975) );
  AND2_X1 U23029 ( .A1(n20476), .A2(n19973), .ZN(n20424) );
  AOI22_X1 U23030 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20002), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20001), .ZN(n20427) );
  AOI22_X1 U23031 ( .A1(n20424), .A2(n20003), .B1(n20030), .B2(n20486), .ZN(
        n19974) );
  OAI211_X1 U23032 ( .C1(n20006), .C2(n13603), .A(n19975), .B(n19974), .ZN(
        P2_U3049) );
  INV_X1 U23033 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19980) );
  AOI22_X1 U23034 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n20001), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n20002), .ZN(n20496) );
  INV_X1 U23035 ( .A(n20496), .ZN(n20429) );
  AND2_X1 U23036 ( .A1(n19998), .A2(n19976), .ZN(n20428) );
  AOI22_X1 U23037 ( .A1(n20429), .A2(n10554), .B1(n19999), .B2(n20428), .ZN(
        n19979) );
  AND2_X1 U23038 ( .A1(n20476), .A2(n19977), .ZN(n20430) );
  AOI22_X1 U23039 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20002), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20001), .ZN(n20433) );
  AOI22_X1 U23040 ( .A1(n20430), .A2(n20003), .B1(n20030), .B2(n20493), .ZN(
        n19978) );
  OAI211_X1 U23041 ( .C1(n20006), .C2(n19980), .A(n19979), .B(n19978), .ZN(
        P2_U3050) );
  INV_X1 U23042 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19983) );
  AOI22_X1 U23043 ( .A1(n20435), .A2(n10554), .B1(n20434), .B2(n19999), .ZN(
        n19982) );
  AOI22_X1 U23044 ( .A1(n20436), .A2(n20003), .B1(n20030), .B2(n20500), .ZN(
        n19981) );
  OAI211_X1 U23045 ( .C1(n20006), .C2(n19983), .A(n19982), .B(n19981), .ZN(
        P2_U3051) );
  INV_X1 U23046 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19988) );
  AOI22_X1 U23047 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20002), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n20001), .ZN(n20510) );
  INV_X1 U23048 ( .A(n20510), .ZN(n20383) );
  AND2_X1 U23049 ( .A1(n19998), .A2(n19984), .ZN(n20440) );
  AOI22_X1 U23050 ( .A1(n20383), .A2(n10554), .B1(n19999), .B2(n20440), .ZN(
        n19987) );
  AND2_X1 U23051 ( .A1(n20476), .A2(n19985), .ZN(n20441) );
  AOI22_X1 U23052 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20002), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n20001), .ZN(n20386) );
  AOI22_X1 U23053 ( .A1(n20441), .A2(n20003), .B1(n20030), .B2(n20507), .ZN(
        n19986) );
  OAI211_X1 U23054 ( .C1(n20006), .C2(n19988), .A(n19987), .B(n19986), .ZN(
        P2_U3052) );
  INV_X1 U23055 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n19993) );
  AOI22_X1 U23056 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20002), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n20001), .ZN(n20517) );
  INV_X1 U23057 ( .A(n20517), .ZN(n20445) );
  AOI22_X1 U23058 ( .A1(n20445), .A2(n10554), .B1(n19999), .B2(n20444), .ZN(
        n19992) );
  AND2_X1 U23059 ( .A1(n20476), .A2(n19990), .ZN(n20446) );
  AOI22_X1 U23060 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20002), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n20001), .ZN(n20449) );
  AOI22_X1 U23061 ( .A1(n20446), .A2(n20003), .B1(n20030), .B2(n20514), .ZN(
        n19991) );
  OAI211_X1 U23062 ( .C1(n20006), .C2(n19993), .A(n19992), .B(n19991), .ZN(
        P2_U3053) );
  INV_X1 U23063 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19997) );
  AOI22_X1 U23064 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n20001), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n20002), .ZN(n20524) );
  INV_X1 U23065 ( .A(n20524), .ZN(n20391) );
  AND2_X1 U23066 ( .A1(n19998), .A2(n10794), .ZN(n20450) );
  AOI22_X1 U23067 ( .A1(n20391), .A2(n10554), .B1(n19999), .B2(n20450), .ZN(
        n19996) );
  AND2_X1 U23068 ( .A1(n20476), .A2(n19994), .ZN(n20451) );
  AOI22_X1 U23069 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20002), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n20001), .ZN(n20395) );
  AOI22_X1 U23070 ( .A1(n20451), .A2(n20003), .B1(n20030), .B2(n20521), .ZN(
        n19995) );
  OAI211_X1 U23071 ( .C1(n20006), .C2(n19997), .A(n19996), .B(n19995), .ZN(
        P2_U3054) );
  AOI22_X1 U23072 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20002), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n20001), .ZN(n20535) );
  INV_X1 U23073 ( .A(n20535), .ZN(n20399) );
  AND2_X1 U23074 ( .A1(n19998), .A2(n10786), .ZN(n20455) );
  AOI22_X1 U23075 ( .A1(n20399), .A2(n10554), .B1(n19999), .B2(n20455), .ZN(
        n20005) );
  AND2_X1 U23076 ( .A1(n20476), .A2(n20000), .ZN(n20458) );
  AOI22_X1 U23077 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20002), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n20001), .ZN(n20344) );
  AOI22_X1 U23078 ( .A1(n20458), .A2(n20003), .B1(n20030), .B2(n20530), .ZN(
        n20004) );
  OAI211_X1 U23079 ( .C1(n20006), .C2(n14210), .A(n20005), .B(n20004), .ZN(
        P2_U3055) );
  NOR3_X2 U23080 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20667), .A3(
        n20064), .ZN(n20028) );
  OR2_X1 U23081 ( .A1(n20064), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20009) );
  OAI21_X1 U23082 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20009), .A(n20463), 
        .ZN(n20010) );
  AOI22_X1 U23083 ( .A1(n20029), .A2(n20418), .B1(n20407), .B2(n20028), .ZN(
        n20015) );
  NOR3_X1 U23084 ( .A1(n20640), .A2(P2_STATE2_REG_3__SCAN_IN), .A3(n20247), 
        .ZN(n20013) );
  NOR3_X1 U23085 ( .A1(n20661), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(
        n20064), .ZN(n20012) );
  OAI211_X1 U23086 ( .C1(n20013), .C2(n20012), .A(n20476), .B(n20011), .ZN(
        n20031) );
  AOI22_X1 U23087 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20031), .B1(
        n20030), .B2(n20408), .ZN(n20014) );
  OAI211_X1 U23088 ( .C1(n20421), .C2(n20062), .A(n20015), .B(n20014), .ZN(
        P2_U3056) );
  AOI22_X1 U23089 ( .A1(n20029), .A2(n20424), .B1(n20422), .B2(n20028), .ZN(
        n20017) );
  AOI22_X1 U23090 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20031), .B1(
        n20030), .B2(n20423), .ZN(n20016) );
  OAI211_X1 U23091 ( .C1(n20427), .C2(n20062), .A(n20017), .B(n20016), .ZN(
        P2_U3057) );
  AOI22_X1 U23092 ( .A1(n20029), .A2(n20430), .B1(n20428), .B2(n20028), .ZN(
        n20019) );
  AOI22_X1 U23093 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20031), .B1(
        n20030), .B2(n20429), .ZN(n20018) );
  OAI211_X1 U23094 ( .C1(n20433), .C2(n20062), .A(n20019), .B(n20018), .ZN(
        P2_U3058) );
  AOI22_X1 U23095 ( .A1(n20029), .A2(n20436), .B1(n20434), .B2(n20028), .ZN(
        n20021) );
  AOI22_X1 U23096 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20031), .B1(
        n20030), .B2(n20435), .ZN(n20020) );
  OAI211_X1 U23097 ( .C1(n20439), .C2(n20062), .A(n20021), .B(n20020), .ZN(
        P2_U3059) );
  AOI22_X1 U23098 ( .A1(n20029), .A2(n20441), .B1(n20440), .B2(n20028), .ZN(
        n20023) );
  AOI22_X1 U23099 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20031), .B1(
        n20030), .B2(n20383), .ZN(n20022) );
  OAI211_X1 U23100 ( .C1(n20386), .C2(n20062), .A(n20023), .B(n20022), .ZN(
        P2_U3060) );
  AOI22_X1 U23101 ( .A1(n20029), .A2(n20446), .B1(n20444), .B2(n20028), .ZN(
        n20025) );
  AOI22_X1 U23102 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20031), .B1(
        n20030), .B2(n20445), .ZN(n20024) );
  OAI211_X1 U23103 ( .C1(n20449), .C2(n20062), .A(n20025), .B(n20024), .ZN(
        P2_U3061) );
  AOI22_X1 U23104 ( .A1(n20029), .A2(n20451), .B1(n20450), .B2(n20028), .ZN(
        n20027) );
  AOI22_X1 U23105 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20031), .B1(
        n20030), .B2(n20391), .ZN(n20026) );
  OAI211_X1 U23106 ( .C1(n20395), .C2(n20062), .A(n20027), .B(n20026), .ZN(
        P2_U3062) );
  AOI22_X1 U23107 ( .A1(n20029), .A2(n20458), .B1(n20455), .B2(n20028), .ZN(
        n20033) );
  AOI22_X1 U23108 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20031), .B1(
        n20030), .B2(n20399), .ZN(n20032) );
  OAI211_X1 U23109 ( .C1(n20344), .C2(n20062), .A(n20033), .B(n20032), .ZN(
        P2_U3063) );
  NOR3_X2 U23110 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20660), .A3(
        n20064), .ZN(n20057) );
  OAI21_X1 U23111 ( .B1(n20035), .B2(n20057), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20034) );
  INV_X1 U23112 ( .A(n20064), .ZN(n20063) );
  NAND2_X1 U23113 ( .A1(n20282), .A2(n20063), .ZN(n20039) );
  AOI22_X1 U23114 ( .A1(n20058), .A2(n20418), .B1(n20407), .B2(n20057), .ZN(
        n20044) );
  INV_X1 U23115 ( .A(n20035), .ZN(n20036) );
  AOI21_X1 U23116 ( .B1(n20036), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20042) );
  INV_X1 U23117 ( .A(n20146), .ZN(n20037) );
  INV_X1 U23118 ( .A(n20630), .ZN(n20321) );
  INV_X1 U23119 ( .A(n20062), .ZN(n20038) );
  OAI21_X1 U23120 ( .B1(n20085), .B2(n20038), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20040) );
  NAND3_X1 U23121 ( .A1(n20040), .A2(n20634), .A3(n20039), .ZN(n20041) );
  AOI22_X1 U23122 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20059), .B1(
        n20085), .B2(n20479), .ZN(n20043) );
  OAI211_X1 U23123 ( .C1(n20482), .C2(n20062), .A(n20044), .B(n20043), .ZN(
        P2_U3064) );
  AOI22_X1 U23124 ( .A1(n20058), .A2(n20424), .B1(n20422), .B2(n20057), .ZN(
        n20046) );
  AOI22_X1 U23125 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20059), .B1(
        n20085), .B2(n20486), .ZN(n20045) );
  OAI211_X1 U23126 ( .C1(n20489), .C2(n20062), .A(n20046), .B(n20045), .ZN(
        P2_U3065) );
  AOI22_X1 U23127 ( .A1(n20058), .A2(n20430), .B1(n20428), .B2(n20057), .ZN(
        n20048) );
  AOI22_X1 U23128 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20059), .B1(
        n20085), .B2(n20493), .ZN(n20047) );
  OAI211_X1 U23129 ( .C1(n20496), .C2(n20062), .A(n20048), .B(n20047), .ZN(
        P2_U3066) );
  AOI22_X1 U23130 ( .A1(n20058), .A2(n20436), .B1(n20434), .B2(n20057), .ZN(
        n20050) );
  AOI22_X1 U23131 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20059), .B1(
        n20085), .B2(n20500), .ZN(n20049) );
  OAI211_X1 U23132 ( .C1(n20503), .C2(n20062), .A(n20050), .B(n20049), .ZN(
        P2_U3067) );
  AOI22_X1 U23133 ( .A1(n20058), .A2(n20441), .B1(n20440), .B2(n20057), .ZN(
        n20052) );
  AOI22_X1 U23134 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20059), .B1(
        n20085), .B2(n20507), .ZN(n20051) );
  OAI211_X1 U23135 ( .C1(n20510), .C2(n20062), .A(n20052), .B(n20051), .ZN(
        P2_U3068) );
  AOI22_X1 U23136 ( .A1(n20058), .A2(n20446), .B1(n20444), .B2(n20057), .ZN(
        n20054) );
  AOI22_X1 U23137 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20059), .B1(
        n20085), .B2(n20514), .ZN(n20053) );
  OAI211_X1 U23138 ( .C1(n20517), .C2(n20062), .A(n20054), .B(n20053), .ZN(
        P2_U3069) );
  AOI22_X1 U23139 ( .A1(n20058), .A2(n20451), .B1(n20450), .B2(n20057), .ZN(
        n20056) );
  AOI22_X1 U23140 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20059), .B1(
        n20085), .B2(n20521), .ZN(n20055) );
  OAI211_X1 U23141 ( .C1(n20524), .C2(n20062), .A(n20056), .B(n20055), .ZN(
        P2_U3070) );
  AOI22_X1 U23142 ( .A1(n20058), .A2(n20458), .B1(n20455), .B2(n20057), .ZN(
        n20061) );
  AOI22_X1 U23143 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20059), .B1(
        n20085), .B2(n20530), .ZN(n20060) );
  OAI211_X1 U23144 ( .C1(n20535), .C2(n20062), .A(n20061), .B(n20060), .ZN(
        P2_U3071) );
  AND2_X1 U23145 ( .A1(n20313), .A2(n20063), .ZN(n20088) );
  AOI22_X1 U23146 ( .A1(n20089), .A2(n20479), .B1(n20407), .B2(n20088), .ZN(
        n20074) );
  OAI21_X1 U23147 ( .B1(n20640), .B2(n20630), .A(n20634), .ZN(n20072) );
  NOR2_X1 U23148 ( .A1(n20660), .A2(n20064), .ZN(n20068) );
  INV_X1 U23149 ( .A(n20069), .ZN(n20066) );
  INV_X1 U23150 ( .A(n20088), .ZN(n20065) );
  OAI211_X1 U23151 ( .C1(n20066), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20628), 
        .B(n20065), .ZN(n20067) );
  OAI211_X1 U23152 ( .C1(n20072), .C2(n20068), .A(n20476), .B(n20067), .ZN(
        n20091) );
  INV_X1 U23153 ( .A(n20068), .ZN(n20071) );
  OAI21_X1 U23154 ( .B1(n20069), .B2(n20088), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20070) );
  AOI22_X1 U23155 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20091), .B1(
        n20418), .B2(n20090), .ZN(n20073) );
  OAI211_X1 U23156 ( .C1(n20482), .C2(n20094), .A(n20074), .B(n20073), .ZN(
        P2_U3072) );
  AOI22_X1 U23157 ( .A1(n20085), .A2(n20423), .B1(n20088), .B2(n20422), .ZN(
        n20076) );
  AOI22_X1 U23158 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20091), .B1(
        n20424), .B2(n20090), .ZN(n20075) );
  OAI211_X1 U23159 ( .C1(n20427), .C2(n20112), .A(n20076), .B(n20075), .ZN(
        P2_U3073) );
  AOI22_X1 U23160 ( .A1(n20085), .A2(n20429), .B1(n20088), .B2(n20428), .ZN(
        n20078) );
  AOI22_X1 U23161 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20091), .B1(
        n20430), .B2(n20090), .ZN(n20077) );
  OAI211_X1 U23162 ( .C1(n20433), .C2(n20112), .A(n20078), .B(n20077), .ZN(
        P2_U3074) );
  AOI22_X1 U23163 ( .A1(n20085), .A2(n20435), .B1(n20434), .B2(n20088), .ZN(
        n20080) );
  AOI22_X1 U23164 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20091), .B1(
        n20436), .B2(n20090), .ZN(n20079) );
  OAI211_X1 U23165 ( .C1(n20439), .C2(n20112), .A(n20080), .B(n20079), .ZN(
        P2_U3075) );
  AOI22_X1 U23166 ( .A1(n20089), .A2(n20507), .B1(n20088), .B2(n20440), .ZN(
        n20082) );
  AOI22_X1 U23167 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20091), .B1(
        n20441), .B2(n20090), .ZN(n20081) );
  OAI211_X1 U23168 ( .C1(n20510), .C2(n20094), .A(n20082), .B(n20081), .ZN(
        P2_U3076) );
  AOI22_X1 U23169 ( .A1(n20089), .A2(n20514), .B1(n20088), .B2(n20444), .ZN(
        n20084) );
  AOI22_X1 U23170 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20091), .B1(
        n20446), .B2(n20090), .ZN(n20083) );
  OAI211_X1 U23171 ( .C1(n20517), .C2(n20094), .A(n20084), .B(n20083), .ZN(
        P2_U3077) );
  AOI22_X1 U23172 ( .A1(n20085), .A2(n20391), .B1(n20088), .B2(n20450), .ZN(
        n20087) );
  AOI22_X1 U23173 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20091), .B1(
        n20451), .B2(n20090), .ZN(n20086) );
  OAI211_X1 U23174 ( .C1(n20395), .C2(n20112), .A(n20087), .B(n20086), .ZN(
        P2_U3078) );
  AOI22_X1 U23175 ( .A1(n20089), .A2(n20530), .B1(n20088), .B2(n20455), .ZN(
        n20093) );
  AOI22_X1 U23176 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20091), .B1(
        n20458), .B2(n20090), .ZN(n20092) );
  OAI211_X1 U23177 ( .C1(n20535), .C2(n20094), .A(n20093), .B(n20092), .ZN(
        P2_U3079) );
  AOI22_X1 U23178 ( .A1(n20108), .A2(n20424), .B1(n20422), .B2(n20107), .ZN(
        n20096) );
  AOI22_X1 U23179 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20109), .B1(
        n20134), .B2(n20486), .ZN(n20095) );
  OAI211_X1 U23180 ( .C1(n20489), .C2(n20112), .A(n20096), .B(n20095), .ZN(
        P2_U3081) );
  AOI22_X1 U23181 ( .A1(n20108), .A2(n20430), .B1(n20428), .B2(n20107), .ZN(
        n20098) );
  AOI22_X1 U23182 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20109), .B1(
        n20134), .B2(n20493), .ZN(n20097) );
  OAI211_X1 U23183 ( .C1(n20496), .C2(n20112), .A(n20098), .B(n20097), .ZN(
        P2_U3082) );
  AOI22_X1 U23184 ( .A1(n20108), .A2(n20436), .B1(n20434), .B2(n20107), .ZN(
        n20100) );
  AOI22_X1 U23185 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20109), .B1(
        n20134), .B2(n20500), .ZN(n20099) );
  OAI211_X1 U23186 ( .C1(n20503), .C2(n20112), .A(n20100), .B(n20099), .ZN(
        P2_U3083) );
  AOI22_X1 U23187 ( .A1(n20108), .A2(n20441), .B1(n20440), .B2(n20107), .ZN(
        n20102) );
  AOI22_X1 U23188 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20109), .B1(
        n20134), .B2(n20507), .ZN(n20101) );
  OAI211_X1 U23189 ( .C1(n20510), .C2(n20112), .A(n20102), .B(n20101), .ZN(
        P2_U3084) );
  AOI22_X1 U23190 ( .A1(n20108), .A2(n20446), .B1(n20444), .B2(n20107), .ZN(
        n20104) );
  AOI22_X1 U23191 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20109), .B1(
        n20134), .B2(n20514), .ZN(n20103) );
  OAI211_X1 U23192 ( .C1(n20517), .C2(n20112), .A(n20104), .B(n20103), .ZN(
        P2_U3085) );
  AOI22_X1 U23193 ( .A1(n20108), .A2(n20451), .B1(n20450), .B2(n20107), .ZN(
        n20106) );
  AOI22_X1 U23194 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20109), .B1(
        n20134), .B2(n20521), .ZN(n20105) );
  OAI211_X1 U23195 ( .C1(n20524), .C2(n20112), .A(n20106), .B(n20105), .ZN(
        P2_U3086) );
  AOI22_X1 U23196 ( .A1(n20108), .A2(n20458), .B1(n20455), .B2(n20107), .ZN(
        n20111) );
  AOI22_X1 U23197 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20109), .B1(
        n20134), .B2(n20530), .ZN(n20110) );
  OAI211_X1 U23198 ( .C1(n20535), .C2(n20112), .A(n20111), .B(n20110), .ZN(
        P2_U3087) );
  NOR3_X2 U23199 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20667), .A3(
        n20113), .ZN(n20137) );
  AOI22_X1 U23200 ( .A1(n20147), .A2(n20479), .B1(n20407), .B2(n20137), .ZN(
        n20123) );
  OAI21_X1 U23201 ( .B1(n20640), .B2(n20114), .A(n20634), .ZN(n20121) );
  NAND2_X1 U23202 ( .A1(n20660), .A2(n20148), .ZN(n20120) );
  INV_X1 U23203 ( .A(n20120), .ZN(n20118) );
  OAI21_X1 U23204 ( .B1(n9635), .B2(n20463), .A(n20276), .ZN(n20116) );
  INV_X1 U23205 ( .A(n20137), .ZN(n20115) );
  AOI21_X1 U23206 ( .B1(n20116), .B2(n20115), .A(n20182), .ZN(n20117) );
  OAI21_X1 U23207 ( .B1(n9635), .B2(n20137), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20119) );
  AOI22_X1 U23208 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20139), .B1(
        n20418), .B2(n20138), .ZN(n20122) );
  OAI211_X1 U23209 ( .C1(n20482), .C2(n20142), .A(n20123), .B(n20122), .ZN(
        P2_U3088) );
  AOI22_X1 U23210 ( .A1(n20134), .A2(n20423), .B1(n20422), .B2(n20137), .ZN(
        n20125) );
  AOI22_X1 U23211 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20139), .B1(
        n20424), .B2(n20138), .ZN(n20124) );
  OAI211_X1 U23212 ( .C1(n20427), .C2(n20173), .A(n20125), .B(n20124), .ZN(
        P2_U3089) );
  AOI22_X1 U23213 ( .A1(n20147), .A2(n20493), .B1(n20137), .B2(n20428), .ZN(
        n20127) );
  AOI22_X1 U23214 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20139), .B1(
        n20430), .B2(n20138), .ZN(n20126) );
  OAI211_X1 U23215 ( .C1(n20496), .C2(n20142), .A(n20127), .B(n20126), .ZN(
        P2_U3090) );
  AOI22_X1 U23216 ( .A1(n20147), .A2(n20500), .B1(n20434), .B2(n20137), .ZN(
        n20129) );
  AOI22_X1 U23217 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20139), .B1(
        n20436), .B2(n20138), .ZN(n20128) );
  OAI211_X1 U23218 ( .C1(n20503), .C2(n20142), .A(n20129), .B(n20128), .ZN(
        P2_U3091) );
  AOI22_X1 U23219 ( .A1(n20147), .A2(n20507), .B1(n20137), .B2(n20440), .ZN(
        n20131) );
  AOI22_X1 U23220 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20139), .B1(
        n20441), .B2(n20138), .ZN(n20130) );
  OAI211_X1 U23221 ( .C1(n20510), .C2(n20142), .A(n20131), .B(n20130), .ZN(
        P2_U3092) );
  AOI22_X1 U23222 ( .A1(n20445), .A2(n20134), .B1(n20137), .B2(n20444), .ZN(
        n20133) );
  AOI22_X1 U23223 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20139), .B1(
        n20446), .B2(n20138), .ZN(n20132) );
  OAI211_X1 U23224 ( .C1(n20449), .C2(n20173), .A(n20133), .B(n20132), .ZN(
        P2_U3093) );
  AOI22_X1 U23225 ( .A1(n20391), .A2(n20134), .B1(n20137), .B2(n20450), .ZN(
        n20136) );
  AOI22_X1 U23226 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20139), .B1(
        n20451), .B2(n20138), .ZN(n20135) );
  OAI211_X1 U23227 ( .C1(n20395), .C2(n20173), .A(n20136), .B(n20135), .ZN(
        P2_U3094) );
  AOI22_X1 U23228 ( .A1(n20147), .A2(n20530), .B1(n20137), .B2(n20455), .ZN(
        n20141) );
  AOI22_X1 U23229 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20139), .B1(
        n20458), .B2(n20138), .ZN(n20140) );
  OAI211_X1 U23230 ( .C1(n20535), .C2(n20142), .A(n20141), .B(n20140), .ZN(
        P2_U3095) );
  NAND3_X1 U23231 ( .A1(n20149), .A2(n20148), .A3(n20276), .ZN(n20145) );
  INV_X1 U23232 ( .A(n20143), .ZN(n20144) );
  NAND2_X1 U23233 ( .A1(n20406), .A2(n20643), .ZN(n20183) );
  NOR2_X1 U23234 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20183), .ZN(
        n20168) );
  AOI22_X1 U23235 ( .A1(n20169), .A2(n20418), .B1(n20407), .B2(n20168), .ZN(
        n20155) );
  OAI21_X1 U23236 ( .B1(n20147), .B2(n20208), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20152) );
  NAND2_X1 U23237 ( .A1(n20149), .A2(n20148), .ZN(n20151) );
  AOI211_X1 U23238 ( .C1(n20152), .C2(n20151), .A(n20182), .B(n20150), .ZN(
        n20153) );
  AOI22_X1 U23239 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20170), .B1(
        n20208), .B2(n20479), .ZN(n20154) );
  OAI211_X1 U23240 ( .C1(n20482), .C2(n20173), .A(n20155), .B(n20154), .ZN(
        P2_U3096) );
  AOI22_X1 U23241 ( .A1(n20169), .A2(n20424), .B1(n20422), .B2(n20168), .ZN(
        n20157) );
  AOI22_X1 U23242 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20170), .B1(
        n20208), .B2(n20486), .ZN(n20156) );
  OAI211_X1 U23243 ( .C1(n20489), .C2(n20173), .A(n20157), .B(n20156), .ZN(
        P2_U3097) );
  AOI22_X1 U23244 ( .A1(n20169), .A2(n20430), .B1(n20428), .B2(n20168), .ZN(
        n20159) );
  AOI22_X1 U23245 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20170), .B1(
        n20208), .B2(n20493), .ZN(n20158) );
  OAI211_X1 U23246 ( .C1(n20496), .C2(n20173), .A(n20159), .B(n20158), .ZN(
        P2_U3098) );
  AOI22_X1 U23247 ( .A1(n20169), .A2(n20436), .B1(n20434), .B2(n20168), .ZN(
        n20161) );
  AOI22_X1 U23248 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20170), .B1(
        n20208), .B2(n20500), .ZN(n20160) );
  OAI211_X1 U23249 ( .C1(n20503), .C2(n20173), .A(n20161), .B(n20160), .ZN(
        P2_U3099) );
  AOI22_X1 U23250 ( .A1(n20169), .A2(n20441), .B1(n20440), .B2(n20168), .ZN(
        n20163) );
  AOI22_X1 U23251 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20170), .B1(
        n20208), .B2(n20507), .ZN(n20162) );
  OAI211_X1 U23252 ( .C1(n20510), .C2(n20173), .A(n20163), .B(n20162), .ZN(
        P2_U3100) );
  AOI22_X1 U23253 ( .A1(n20169), .A2(n20446), .B1(n20444), .B2(n20168), .ZN(
        n20165) );
  AOI22_X1 U23254 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20170), .B1(
        n20208), .B2(n20514), .ZN(n20164) );
  OAI211_X1 U23255 ( .C1(n20517), .C2(n20173), .A(n20165), .B(n20164), .ZN(
        P2_U3101) );
  AOI22_X1 U23256 ( .A1(n20169), .A2(n20451), .B1(n20450), .B2(n20168), .ZN(
        n20167) );
  AOI22_X1 U23257 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20170), .B1(
        n20208), .B2(n20521), .ZN(n20166) );
  OAI211_X1 U23258 ( .C1(n20524), .C2(n20173), .A(n20167), .B(n20166), .ZN(
        P2_U3102) );
  AOI22_X1 U23259 ( .A1(n20169), .A2(n20458), .B1(n20455), .B2(n20168), .ZN(
        n20172) );
  AOI22_X1 U23260 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20170), .B1(
        n20208), .B2(n20530), .ZN(n20171) );
  OAI211_X1 U23261 ( .C1(n20535), .C2(n20173), .A(n20172), .B(n20171), .ZN(
        P2_U3103) );
  NAND2_X1 U23262 ( .A1(n20216), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20175) );
  NOR2_X1 U23263 ( .A1(n20176), .A2(n20175), .ZN(n20181) );
  INV_X1 U23264 ( .A(n20183), .ZN(n20177) );
  AOI21_X1 U23265 ( .B1(n20276), .B2(n20177), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20178) );
  INV_X1 U23266 ( .A(n20418), .ZN(n20469) );
  OAI22_X1 U23267 ( .A1(n20206), .A2(n20469), .B1(n20216), .B2(n20468), .ZN(
        n20179) );
  INV_X1 U23268 ( .A(n20179), .ZN(n20187) );
  INV_X1 U23269 ( .A(n20640), .ZN(n20180) );
  INV_X1 U23270 ( .A(n20629), .ZN(n20471) );
  NAND2_X1 U23271 ( .A1(n20180), .A2(n20471), .ZN(n20184) );
  AOI211_X1 U23272 ( .C1(n20184), .C2(n20183), .A(n20182), .B(n20181), .ZN(
        n20185) );
  OAI21_X1 U23273 ( .B1(n20219), .B2(n20276), .A(n20185), .ZN(n20209) );
  AOI22_X1 U23274 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20209), .B1(
        n20208), .B2(n20408), .ZN(n20186) );
  OAI211_X1 U23275 ( .C1(n20421), .C2(n20242), .A(n20187), .B(n20186), .ZN(
        P2_U3104) );
  INV_X1 U23276 ( .A(n20424), .ZN(n20484) );
  INV_X1 U23277 ( .A(n20422), .ZN(n20483) );
  OAI22_X1 U23278 ( .A1(n20206), .A2(n20484), .B1(n20216), .B2(n20483), .ZN(
        n20188) );
  INV_X1 U23279 ( .A(n20188), .ZN(n20190) );
  AOI22_X1 U23280 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20209), .B1(
        n20208), .B2(n20423), .ZN(n20189) );
  OAI211_X1 U23281 ( .C1(n20427), .C2(n20242), .A(n20190), .B(n20189), .ZN(
        P2_U3105) );
  INV_X1 U23282 ( .A(n20430), .ZN(n20491) );
  INV_X1 U23283 ( .A(n20428), .ZN(n20490) );
  OAI22_X1 U23284 ( .A1(n20206), .A2(n20491), .B1(n20216), .B2(n20490), .ZN(
        n20191) );
  INV_X1 U23285 ( .A(n20191), .ZN(n20193) );
  AOI22_X1 U23286 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20209), .B1(
        n20208), .B2(n20429), .ZN(n20192) );
  OAI211_X1 U23287 ( .C1(n20433), .C2(n20242), .A(n20193), .B(n20192), .ZN(
        P2_U3106) );
  INV_X1 U23288 ( .A(n20436), .ZN(n20498) );
  INV_X1 U23289 ( .A(n20434), .ZN(n20497) );
  OAI22_X1 U23290 ( .A1(n20206), .A2(n20498), .B1(n20216), .B2(n20497), .ZN(
        n20194) );
  INV_X1 U23291 ( .A(n20194), .ZN(n20196) );
  AOI22_X1 U23292 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20209), .B1(
        n20208), .B2(n20435), .ZN(n20195) );
  OAI211_X1 U23293 ( .C1(n20439), .C2(n20242), .A(n20196), .B(n20195), .ZN(
        P2_U3107) );
  INV_X1 U23294 ( .A(n20441), .ZN(n20505) );
  INV_X1 U23295 ( .A(n20440), .ZN(n20504) );
  OAI22_X1 U23296 ( .A1(n20206), .A2(n20505), .B1(n20216), .B2(n20504), .ZN(
        n20197) );
  INV_X1 U23297 ( .A(n20197), .ZN(n20199) );
  AOI22_X1 U23298 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20209), .B1(
        n20208), .B2(n20383), .ZN(n20198) );
  OAI211_X1 U23299 ( .C1(n20386), .C2(n20242), .A(n20199), .B(n20198), .ZN(
        P2_U3108) );
  INV_X1 U23300 ( .A(n20446), .ZN(n20512) );
  INV_X1 U23301 ( .A(n20444), .ZN(n20511) );
  OAI22_X1 U23302 ( .A1(n20206), .A2(n20512), .B1(n20216), .B2(n20511), .ZN(
        n20200) );
  INV_X1 U23303 ( .A(n20200), .ZN(n20202) );
  AOI22_X1 U23304 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20209), .B1(
        n20208), .B2(n20445), .ZN(n20201) );
  OAI211_X1 U23305 ( .C1(n20449), .C2(n20242), .A(n20202), .B(n20201), .ZN(
        P2_U3109) );
  INV_X1 U23306 ( .A(n20451), .ZN(n20519) );
  INV_X1 U23307 ( .A(n20450), .ZN(n20518) );
  OAI22_X1 U23308 ( .A1(n20206), .A2(n20519), .B1(n20216), .B2(n20518), .ZN(
        n20203) );
  INV_X1 U23309 ( .A(n20203), .ZN(n20205) );
  AOI22_X1 U23310 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20209), .B1(
        n20208), .B2(n20391), .ZN(n20204) );
  OAI211_X1 U23311 ( .C1(n20395), .C2(n20242), .A(n20205), .B(n20204), .ZN(
        P2_U3110) );
  INV_X1 U23312 ( .A(n20458), .ZN(n20527) );
  INV_X1 U23313 ( .A(n20455), .ZN(n20526) );
  OAI22_X1 U23314 ( .A1(n20206), .A2(n20527), .B1(n20216), .B2(n20526), .ZN(
        n20207) );
  INV_X1 U23315 ( .A(n20207), .ZN(n20211) );
  AOI22_X1 U23316 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20209), .B1(
        n20208), .B2(n20399), .ZN(n20210) );
  OAI211_X1 U23317 ( .C1(n20344), .C2(n20242), .A(n20211), .B(n20210), .ZN(
        P2_U3111) );
  NAND2_X1 U23318 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20651), .ZN(
        n20311) );
  NOR2_X1 U23319 ( .A1(n20212), .A2(n20311), .ZN(n20237) );
  AOI22_X1 U23320 ( .A1(n10547), .A2(n20479), .B1(n20407), .B2(n20237), .ZN(
        n20224) );
  NOR3_X1 U23321 ( .A1(n10547), .A2(n20213), .A3(n20628), .ZN(n20214) );
  NOR2_X1 U23322 ( .A1(n20214), .A2(n20632), .ZN(n20222) );
  INV_X1 U23323 ( .A(n20222), .ZN(n20217) );
  AOI21_X1 U23324 ( .B1(n10921), .B2(n20276), .A(n20634), .ZN(n20215) );
  AOI21_X1 U23325 ( .B1(n20217), .B2(n20216), .A(n20215), .ZN(n20218) );
  NOR2_X1 U23326 ( .A1(n20219), .A2(n20237), .ZN(n20221) );
  OAI21_X1 U23327 ( .B1(n10921), .B2(n20237), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20220) );
  AOI22_X1 U23328 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20239), .B1(
        n20418), .B2(n20238), .ZN(n20223) );
  OAI211_X1 U23329 ( .C1(n20482), .C2(n20242), .A(n20224), .B(n20223), .ZN(
        P2_U3112) );
  AOI22_X1 U23330 ( .A1(n20486), .A2(n10547), .B1(n20422), .B2(n20237), .ZN(
        n20226) );
  AOI22_X1 U23331 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20239), .B1(
        n20238), .B2(n20424), .ZN(n20225) );
  OAI211_X1 U23332 ( .C1(n20489), .C2(n20242), .A(n20226), .B(n20225), .ZN(
        P2_U3113) );
  AOI22_X1 U23333 ( .A1(n10547), .A2(n20493), .B1(n20428), .B2(n20237), .ZN(
        n20228) );
  AOI22_X1 U23334 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20239), .B1(
        n20238), .B2(n20430), .ZN(n20227) );
  OAI211_X1 U23335 ( .C1(n20496), .C2(n20242), .A(n20228), .B(n20227), .ZN(
        P2_U3114) );
  AOI22_X1 U23336 ( .A1(n10547), .A2(n20500), .B1(n20434), .B2(n20237), .ZN(
        n20230) );
  AOI22_X1 U23337 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20239), .B1(
        n20238), .B2(n20436), .ZN(n20229) );
  OAI211_X1 U23338 ( .C1(n20503), .C2(n20242), .A(n20230), .B(n20229), .ZN(
        P2_U3115) );
  AOI22_X1 U23339 ( .A1(n10547), .A2(n20507), .B1(n20440), .B2(n20237), .ZN(
        n20232) );
  AOI22_X1 U23340 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20239), .B1(
        n20238), .B2(n20441), .ZN(n20231) );
  OAI211_X1 U23341 ( .C1(n20510), .C2(n20242), .A(n20232), .B(n20231), .ZN(
        P2_U3116) );
  AOI22_X1 U23342 ( .A1(n10547), .A2(n20514), .B1(n20444), .B2(n20237), .ZN(
        n20234) );
  AOI22_X1 U23343 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20239), .B1(
        n20238), .B2(n20446), .ZN(n20233) );
  OAI211_X1 U23344 ( .C1(n20517), .C2(n20242), .A(n20234), .B(n20233), .ZN(
        P2_U3117) );
  AOI22_X1 U23345 ( .A1(n10547), .A2(n20521), .B1(n20450), .B2(n20237), .ZN(
        n20236) );
  AOI22_X1 U23346 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20239), .B1(
        n20238), .B2(n20451), .ZN(n20235) );
  OAI211_X1 U23347 ( .C1(n20524), .C2(n20242), .A(n20236), .B(n20235), .ZN(
        P2_U3118) );
  AOI22_X1 U23348 ( .A1(n10547), .A2(n20530), .B1(n20455), .B2(n20237), .ZN(
        n20241) );
  AOI22_X1 U23349 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20239), .B1(
        n20238), .B2(n20458), .ZN(n20240) );
  OAI211_X1 U23350 ( .C1(n20535), .C2(n20242), .A(n20241), .B(n20240), .ZN(
        P2_U3119) );
  NOR2_X1 U23351 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20311), .ZN(
        n20244) );
  INV_X1 U23352 ( .A(n20244), .ZN(n20250) );
  NOR2_X1 U23353 ( .A1(n20628), .A2(n20250), .ZN(n20246) );
  INV_X1 U23354 ( .A(n20243), .ZN(n20253) );
  NAND2_X1 U23355 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20244), .ZN(
        n20252) );
  AOI21_X1 U23356 ( .B1(n20253), .B2(n20252), .A(n20463), .ZN(n20245) );
  NOR2_X1 U23357 ( .A1(n20246), .A2(n20245), .ZN(n20274) );
  INV_X1 U23358 ( .A(n20252), .ZN(n20275) );
  AOI22_X1 U23359 ( .A1(n20292), .A2(n20479), .B1(n20407), .B2(n20275), .ZN(
        n20258) );
  NAND2_X1 U23360 ( .A1(n20472), .A2(n20249), .ZN(n20251) );
  NAND2_X1 U23361 ( .A1(n20251), .A2(n20250), .ZN(n20255) );
  OAI21_X1 U23362 ( .B1(n20253), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20252), 
        .ZN(n20254) );
  MUX2_X1 U23363 ( .A(n20255), .B(n20254), .S(n20628), .Z(n20256) );
  NAND2_X1 U23364 ( .A1(n20256), .A2(n20476), .ZN(n20271) );
  AOI22_X1 U23365 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20271), .B1(
        n10547), .B2(n20408), .ZN(n20257) );
  OAI211_X1 U23366 ( .C1(n20274), .C2(n20469), .A(n20258), .B(n20257), .ZN(
        P2_U3120) );
  AOI22_X1 U23367 ( .A1(n10547), .A2(n20423), .B1(n20422), .B2(n20275), .ZN(
        n20260) );
  AOI22_X1 U23368 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20271), .B1(
        n20292), .B2(n20486), .ZN(n20259) );
  OAI211_X1 U23369 ( .C1(n20274), .C2(n20484), .A(n20260), .B(n20259), .ZN(
        P2_U3121) );
  AOI22_X1 U23370 ( .A1(n20292), .A2(n20493), .B1(n20428), .B2(n20275), .ZN(
        n20262) );
  AOI22_X1 U23371 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20271), .B1(
        n10547), .B2(n20429), .ZN(n20261) );
  OAI211_X1 U23372 ( .C1(n20274), .C2(n20491), .A(n20262), .B(n20261), .ZN(
        P2_U3122) );
  AOI22_X1 U23373 ( .A1(n20435), .A2(n10547), .B1(n20434), .B2(n20275), .ZN(
        n20264) );
  AOI22_X1 U23374 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20271), .B1(
        n20292), .B2(n20500), .ZN(n20263) );
  OAI211_X1 U23375 ( .C1(n20274), .C2(n20498), .A(n20264), .B(n20263), .ZN(
        P2_U3123) );
  AOI22_X1 U23376 ( .A1(n20292), .A2(n20507), .B1(n20440), .B2(n20275), .ZN(
        n20266) );
  AOI22_X1 U23377 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20271), .B1(
        n10547), .B2(n20383), .ZN(n20265) );
  OAI211_X1 U23378 ( .C1(n20274), .C2(n20505), .A(n20266), .B(n20265), .ZN(
        P2_U3124) );
  AOI22_X1 U23379 ( .A1(n20292), .A2(n20514), .B1(n20444), .B2(n20275), .ZN(
        n20268) );
  AOI22_X1 U23380 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20271), .B1(
        n10547), .B2(n20445), .ZN(n20267) );
  OAI211_X1 U23381 ( .C1(n20274), .C2(n20512), .A(n20268), .B(n20267), .ZN(
        P2_U3125) );
  AOI22_X1 U23382 ( .A1(n20391), .A2(n10547), .B1(n20450), .B2(n20275), .ZN(
        n20270) );
  AOI22_X1 U23383 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20271), .B1(
        n20292), .B2(n20521), .ZN(n20269) );
  OAI211_X1 U23384 ( .C1(n20274), .C2(n20519), .A(n20270), .B(n20269), .ZN(
        P2_U3126) );
  AOI22_X1 U23385 ( .A1(n20399), .A2(n10547), .B1(n20455), .B2(n20275), .ZN(
        n20273) );
  AOI22_X1 U23386 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20271), .B1(
        n20292), .B2(n20530), .ZN(n20272) );
  OAI211_X1 U23387 ( .C1(n20274), .C2(n20527), .A(n20273), .B(n20272), .ZN(
        P2_U3127) );
  AOI221_X1 U23388 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n20292), .C1(
        P2_STATEBS16_REG_SCAN_IN), .C2(n20340), .A(n20275), .ZN(n20278) );
  OAI21_X1 U23389 ( .B1(n20283), .B2(n20463), .A(n20276), .ZN(n20277) );
  OR2_X1 U23390 ( .A1(n20278), .A2(n20277), .ZN(n20280) );
  NOR2_X1 U23391 ( .A1(n20660), .A2(n20311), .ZN(n20322) );
  INV_X1 U23392 ( .A(n20322), .ZN(n20310) );
  NOR2_X1 U23393 ( .A1(n20310), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20304) );
  INV_X1 U23394 ( .A(n20304), .ZN(n20279) );
  NAND2_X1 U23395 ( .A1(n20280), .A2(n20279), .ZN(n20281) );
  INV_X1 U23396 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n20288) );
  INV_X1 U23397 ( .A(n20282), .ZN(n20285) );
  OAI21_X1 U23398 ( .B1(n20283), .B2(n20304), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20284) );
  AOI22_X1 U23399 ( .A1(n20305), .A2(n20418), .B1(n20407), .B2(n20304), .ZN(
        n20287) );
  AOI22_X1 U23400 ( .A1(n20340), .A2(n20479), .B1(n20292), .B2(n20408), .ZN(
        n20286) );
  OAI211_X1 U23401 ( .C1(n20293), .C2(n20288), .A(n20287), .B(n20286), .ZN(
        P2_U3128) );
  INV_X1 U23402 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n20291) );
  AOI22_X1 U23403 ( .A1(n20305), .A2(n20424), .B1(n20422), .B2(n20304), .ZN(
        n20290) );
  AOI22_X1 U23404 ( .A1(n20340), .A2(n20486), .B1(n20292), .B2(n20423), .ZN(
        n20289) );
  OAI211_X1 U23405 ( .C1(n20293), .C2(n20291), .A(n20290), .B(n20289), .ZN(
        P2_U3129) );
  AOI22_X1 U23406 ( .A1(n20305), .A2(n20430), .B1(n20428), .B2(n20304), .ZN(
        n20295) );
  AOI22_X1 U23407 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20306), .B1(
        n20340), .B2(n20493), .ZN(n20294) );
  OAI211_X1 U23408 ( .C1(n20496), .C2(n20248), .A(n20295), .B(n20294), .ZN(
        P2_U3130) );
  AOI22_X1 U23409 ( .A1(n20305), .A2(n20436), .B1(n20434), .B2(n20304), .ZN(
        n20297) );
  AOI22_X1 U23410 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20306), .B1(
        n20340), .B2(n20500), .ZN(n20296) );
  OAI211_X1 U23411 ( .C1(n20503), .C2(n20248), .A(n20297), .B(n20296), .ZN(
        P2_U3131) );
  AOI22_X1 U23412 ( .A1(n20305), .A2(n20441), .B1(n20440), .B2(n20304), .ZN(
        n20299) );
  AOI22_X1 U23413 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20306), .B1(
        n20340), .B2(n20507), .ZN(n20298) );
  OAI211_X1 U23414 ( .C1(n20510), .C2(n20248), .A(n20299), .B(n20298), .ZN(
        P2_U3132) );
  AOI22_X1 U23415 ( .A1(n20305), .A2(n20446), .B1(n20444), .B2(n20304), .ZN(
        n20301) );
  AOI22_X1 U23416 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20306), .B1(
        n20340), .B2(n20514), .ZN(n20300) );
  OAI211_X1 U23417 ( .C1(n20517), .C2(n20248), .A(n20301), .B(n20300), .ZN(
        P2_U3133) );
  AOI22_X1 U23418 ( .A1(n20305), .A2(n20451), .B1(n20450), .B2(n20304), .ZN(
        n20303) );
  AOI22_X1 U23419 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20306), .B1(
        n20340), .B2(n20521), .ZN(n20302) );
  OAI211_X1 U23420 ( .C1(n20524), .C2(n20248), .A(n20303), .B(n20302), .ZN(
        P2_U3134) );
  AOI22_X1 U23421 ( .A1(n20305), .A2(n20458), .B1(n20455), .B2(n20304), .ZN(
        n20308) );
  AOI22_X1 U23422 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20306), .B1(
        n20340), .B2(n20530), .ZN(n20307) );
  OAI211_X1 U23423 ( .C1(n20535), .C2(n20248), .A(n20308), .B(n20307), .ZN(
        P2_U3135) );
  OR2_X1 U23424 ( .A1(n20310), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20316) );
  INV_X1 U23425 ( .A(n20311), .ZN(n20312) );
  NAND2_X1 U23426 ( .A1(n20313), .A2(n20312), .ZN(n20317) );
  NAND2_X1 U23427 ( .A1(n20317), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20314) );
  INV_X1 U23428 ( .A(n20317), .ZN(n20338) );
  AOI22_X1 U23429 ( .A1(n20339), .A2(n20418), .B1(n20407), .B2(n20338), .ZN(
        n20324) );
  OAI21_X1 U23430 ( .B1(n20338), .B2(n20276), .A(n20476), .ZN(n20318) );
  NOR2_X1 U23431 ( .A1(n20319), .A2(n20318), .ZN(n20320) );
  AOI22_X1 U23432 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20341), .B1(
        n20340), .B2(n20408), .ZN(n20323) );
  OAI211_X1 U23433 ( .C1(n20421), .C2(n20374), .A(n20324), .B(n20323), .ZN(
        P2_U3136) );
  AOI22_X1 U23434 ( .A1(n20339), .A2(n20424), .B1(n20422), .B2(n20338), .ZN(
        n20326) );
  AOI22_X1 U23435 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20341), .B1(
        n20340), .B2(n20423), .ZN(n20325) );
  OAI211_X1 U23436 ( .C1(n20427), .C2(n20374), .A(n20326), .B(n20325), .ZN(
        P2_U3137) );
  AOI22_X1 U23437 ( .A1(n20339), .A2(n20430), .B1(n20428), .B2(n20338), .ZN(
        n20328) );
  AOI22_X1 U23438 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20341), .B1(
        n20350), .B2(n20493), .ZN(n20327) );
  OAI211_X1 U23439 ( .C1(n20496), .C2(n20337), .A(n20328), .B(n20327), .ZN(
        P2_U3138) );
  AOI22_X1 U23440 ( .A1(n20339), .A2(n20436), .B1(n20434), .B2(n20338), .ZN(
        n20330) );
  AOI22_X1 U23441 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20341), .B1(
        n20350), .B2(n20500), .ZN(n20329) );
  OAI211_X1 U23442 ( .C1(n20503), .C2(n20337), .A(n20330), .B(n20329), .ZN(
        P2_U3139) );
  AOI22_X1 U23443 ( .A1(n20339), .A2(n20441), .B1(n20440), .B2(n20338), .ZN(
        n20332) );
  AOI22_X1 U23444 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20341), .B1(
        n20340), .B2(n20383), .ZN(n20331) );
  OAI211_X1 U23445 ( .C1(n20386), .C2(n20374), .A(n20332), .B(n20331), .ZN(
        P2_U3140) );
  AOI22_X1 U23446 ( .A1(n20339), .A2(n20446), .B1(n20444), .B2(n20338), .ZN(
        n20334) );
  AOI22_X1 U23447 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20341), .B1(
        n20350), .B2(n20514), .ZN(n20333) );
  OAI211_X1 U23448 ( .C1(n20517), .C2(n20337), .A(n20334), .B(n20333), .ZN(
        P2_U3141) );
  AOI22_X1 U23449 ( .A1(n20339), .A2(n20451), .B1(n20450), .B2(n20338), .ZN(
        n20336) );
  AOI22_X1 U23450 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20341), .B1(
        n20350), .B2(n20521), .ZN(n20335) );
  OAI211_X1 U23451 ( .C1(n20524), .C2(n20337), .A(n20336), .B(n20335), .ZN(
        P2_U3142) );
  AOI22_X1 U23452 ( .A1(n20339), .A2(n20458), .B1(n20455), .B2(n20338), .ZN(
        n20343) );
  AOI22_X1 U23453 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20341), .B1(
        n20340), .B2(n20399), .ZN(n20342) );
  OAI211_X1 U23454 ( .C1(n20344), .C2(n20374), .A(n20343), .B(n20342), .ZN(
        P2_U3143) );
  INV_X1 U23455 ( .A(n20345), .ZN(n20349) );
  NOR2_X1 U23456 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20346), .ZN(
        n20369) );
  OAI21_X1 U23457 ( .B1(n20347), .B2(n20369), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20348) );
  AOI22_X1 U23458 ( .A1(n20370), .A2(n20418), .B1(n20407), .B2(n20369), .ZN(
        n20356) );
  OAI21_X1 U23459 ( .B1(n20400), .B2(n20350), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20351) );
  OAI21_X1 U23460 ( .B1(n20352), .B2(n20643), .A(n20351), .ZN(n20354) );
  NAND3_X1 U23461 ( .A1(n20354), .A2(n20476), .A3(n20353), .ZN(n20371) );
  AOI22_X1 U23462 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20371), .B1(
        n20400), .B2(n20479), .ZN(n20355) );
  OAI211_X1 U23463 ( .C1(n20482), .C2(n20374), .A(n20356), .B(n20355), .ZN(
        P2_U3144) );
  AOI22_X1 U23464 ( .A1(n20370), .A2(n20424), .B1(n20422), .B2(n20369), .ZN(
        n20358) );
  AOI22_X1 U23465 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20371), .B1(
        n20400), .B2(n20486), .ZN(n20357) );
  OAI211_X1 U23466 ( .C1(n20489), .C2(n20374), .A(n20358), .B(n20357), .ZN(
        P2_U3145) );
  AOI22_X1 U23467 ( .A1(n20370), .A2(n20430), .B1(n20428), .B2(n20369), .ZN(
        n20360) );
  AOI22_X1 U23468 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20371), .B1(
        n20400), .B2(n20493), .ZN(n20359) );
  OAI211_X1 U23469 ( .C1(n20496), .C2(n20374), .A(n20360), .B(n20359), .ZN(
        P2_U3146) );
  AOI22_X1 U23470 ( .A1(n20370), .A2(n20436), .B1(n20434), .B2(n20369), .ZN(
        n20362) );
  AOI22_X1 U23471 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20371), .B1(
        n20400), .B2(n20500), .ZN(n20361) );
  OAI211_X1 U23472 ( .C1(n20503), .C2(n20374), .A(n20362), .B(n20361), .ZN(
        P2_U3147) );
  AOI22_X1 U23473 ( .A1(n20370), .A2(n20441), .B1(n20440), .B2(n20369), .ZN(
        n20364) );
  AOI22_X1 U23474 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20371), .B1(
        n20400), .B2(n20507), .ZN(n20363) );
  OAI211_X1 U23475 ( .C1(n20510), .C2(n20374), .A(n20364), .B(n20363), .ZN(
        P2_U3148) );
  AOI22_X1 U23476 ( .A1(n20370), .A2(n20446), .B1(n20444), .B2(n20369), .ZN(
        n20366) );
  AOI22_X1 U23477 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20371), .B1(
        n20400), .B2(n20514), .ZN(n20365) );
  OAI211_X1 U23478 ( .C1(n20517), .C2(n20374), .A(n20366), .B(n20365), .ZN(
        P2_U3149) );
  AOI22_X1 U23479 ( .A1(n20370), .A2(n20451), .B1(n20450), .B2(n20369), .ZN(
        n20368) );
  AOI22_X1 U23480 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20371), .B1(
        n20400), .B2(n20521), .ZN(n20367) );
  OAI211_X1 U23481 ( .C1(n20524), .C2(n20374), .A(n20368), .B(n20367), .ZN(
        P2_U3150) );
  AOI22_X1 U23482 ( .A1(n20370), .A2(n20458), .B1(n20455), .B2(n20369), .ZN(
        n20373) );
  AOI22_X1 U23483 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20371), .B1(
        n20400), .B2(n20530), .ZN(n20372) );
  OAI211_X1 U23484 ( .C1(n20535), .C2(n20374), .A(n20373), .B(n20372), .ZN(
        P2_U3151) );
  OAI22_X1 U23485 ( .A1(n20397), .A2(n20484), .B1(n20396), .B2(n20483), .ZN(
        n20375) );
  INV_X1 U23486 ( .A(n20375), .ZN(n20377) );
  AOI22_X1 U23487 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20392), .B1(
        n20400), .B2(n20423), .ZN(n20376) );
  OAI211_X1 U23488 ( .C1(n20427), .C2(n20462), .A(n20377), .B(n20376), .ZN(
        P2_U3153) );
  INV_X1 U23489 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n20381) );
  OAI22_X1 U23490 ( .A1(n20397), .A2(n20491), .B1(n20396), .B2(n20490), .ZN(
        n20378) );
  INV_X1 U23491 ( .A(n20378), .ZN(n20380) );
  AOI22_X1 U23492 ( .A1(n10553), .A2(n20493), .B1(n20400), .B2(n20429), .ZN(
        n20379) );
  OAI211_X1 U23493 ( .C1(n20404), .C2(n20381), .A(n20380), .B(n20379), .ZN(
        P2_U3154) );
  OAI22_X1 U23494 ( .A1(n20397), .A2(n20505), .B1(n20396), .B2(n20504), .ZN(
        n20382) );
  INV_X1 U23495 ( .A(n20382), .ZN(n20385) );
  AOI22_X1 U23496 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20392), .B1(
        n20400), .B2(n20383), .ZN(n20384) );
  OAI211_X1 U23497 ( .C1(n20386), .C2(n20462), .A(n20385), .B(n20384), .ZN(
        P2_U3156) );
  OAI22_X1 U23498 ( .A1(n20397), .A2(n20512), .B1(n20396), .B2(n20511), .ZN(
        n20387) );
  INV_X1 U23499 ( .A(n20387), .ZN(n20389) );
  AOI22_X1 U23500 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20392), .B1(
        n20400), .B2(n20445), .ZN(n20388) );
  OAI211_X1 U23501 ( .C1(n20449), .C2(n20462), .A(n20389), .B(n20388), .ZN(
        P2_U3157) );
  OAI22_X1 U23502 ( .A1(n20397), .A2(n20519), .B1(n20396), .B2(n20518), .ZN(
        n20390) );
  INV_X1 U23503 ( .A(n20390), .ZN(n20394) );
  AOI22_X1 U23504 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20392), .B1(
        n20400), .B2(n20391), .ZN(n20393) );
  OAI211_X1 U23505 ( .C1(n20395), .C2(n20462), .A(n20394), .B(n20393), .ZN(
        P2_U3158) );
  INV_X1 U23506 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n20403) );
  OAI22_X1 U23507 ( .A1(n20397), .A2(n20527), .B1(n20396), .B2(n20526), .ZN(
        n20398) );
  INV_X1 U23508 ( .A(n20398), .ZN(n20402) );
  AOI22_X1 U23509 ( .A1(n10553), .A2(n20530), .B1(n20400), .B2(n20399), .ZN(
        n20401) );
  OAI211_X1 U23510 ( .C1(n20404), .C2(n20403), .A(n20402), .B(n20401), .ZN(
        P2_U3159) );
  NAND2_X1 U23511 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20406), .ZN(
        n20474) );
  NOR2_X1 U23512 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20474), .ZN(
        n20454) );
  AOI22_X1 U23513 ( .A1(n20408), .A2(n10553), .B1(n20407), .B2(n20454), .ZN(
        n20420) );
  NOR3_X1 U23514 ( .A1(n20456), .A2(n10553), .A3(n20628), .ZN(n20409) );
  NOR2_X1 U23515 ( .A1(n20409), .A2(n20632), .ZN(n20417) );
  NOR2_X1 U23516 ( .A1(n20454), .A2(n20410), .ZN(n20416) );
  INV_X1 U23517 ( .A(n20416), .ZN(n20413) );
  INV_X1 U23518 ( .A(n20454), .ZN(n20411) );
  OAI211_X1 U23519 ( .C1(n10926), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20628), 
        .B(n20411), .ZN(n20412) );
  OAI211_X1 U23520 ( .C1(n20417), .C2(n20413), .A(n20476), .B(n20412), .ZN(
        n20459) );
  INV_X1 U23521 ( .A(n10926), .ZN(n20414) );
  OAI21_X1 U23522 ( .B1(n20414), .B2(n20454), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20415) );
  AOI22_X1 U23523 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20459), .B1(
        n20418), .B2(n20457), .ZN(n20419) );
  OAI211_X1 U23524 ( .C1(n20421), .C2(n20534), .A(n20420), .B(n20419), .ZN(
        P2_U3160) );
  AOI22_X1 U23525 ( .A1(n10553), .A2(n20423), .B1(n20422), .B2(n20454), .ZN(
        n20426) );
  AOI22_X1 U23526 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20459), .B1(
        n20424), .B2(n20457), .ZN(n20425) );
  OAI211_X1 U23527 ( .C1(n20427), .C2(n20534), .A(n20426), .B(n20425), .ZN(
        P2_U3161) );
  AOI22_X1 U23528 ( .A1(n20429), .A2(n10553), .B1(n20428), .B2(n20454), .ZN(
        n20432) );
  AOI22_X1 U23529 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20459), .B1(
        n20430), .B2(n20457), .ZN(n20431) );
  OAI211_X1 U23530 ( .C1(n20433), .C2(n20534), .A(n20432), .B(n20431), .ZN(
        P2_U3162) );
  AOI22_X1 U23531 ( .A1(n20435), .A2(n10553), .B1(n20434), .B2(n20454), .ZN(
        n20438) );
  AOI22_X1 U23532 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20459), .B1(
        n20436), .B2(n20457), .ZN(n20437) );
  OAI211_X1 U23533 ( .C1(n20439), .C2(n20534), .A(n20438), .B(n20437), .ZN(
        P2_U3163) );
  AOI22_X1 U23534 ( .A1(n20456), .A2(n20507), .B1(n20440), .B2(n20454), .ZN(
        n20443) );
  AOI22_X1 U23535 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20459), .B1(
        n20441), .B2(n20457), .ZN(n20442) );
  OAI211_X1 U23536 ( .C1(n20510), .C2(n20462), .A(n20443), .B(n20442), .ZN(
        P2_U3164) );
  AOI22_X1 U23537 ( .A1(n20445), .A2(n10553), .B1(n20444), .B2(n20454), .ZN(
        n20448) );
  AOI22_X1 U23538 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20459), .B1(
        n20446), .B2(n20457), .ZN(n20447) );
  OAI211_X1 U23539 ( .C1(n20449), .C2(n20534), .A(n20448), .B(n20447), .ZN(
        P2_U3165) );
  AOI22_X1 U23540 ( .A1(n20456), .A2(n20521), .B1(n20450), .B2(n20454), .ZN(
        n20453) );
  AOI22_X1 U23541 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20459), .B1(
        n20451), .B2(n20457), .ZN(n20452) );
  OAI211_X1 U23542 ( .C1(n20524), .C2(n20462), .A(n20453), .B(n20452), .ZN(
        P2_U3166) );
  AOI22_X1 U23543 ( .A1(n20456), .A2(n20530), .B1(n20455), .B2(n20454), .ZN(
        n20461) );
  AOI22_X1 U23544 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20459), .B1(
        n20458), .B2(n20457), .ZN(n20460) );
  OAI211_X1 U23545 ( .C1(n20535), .C2(n20462), .A(n20461), .B(n20460), .ZN(
        P2_U3167) );
  OR2_X1 U23546 ( .A1(n20478), .A2(n20463), .ZN(n20464) );
  NOR2_X1 U23547 ( .A1(n20465), .A2(n20464), .ZN(n20473) );
  INV_X1 U23548 ( .A(n20474), .ZN(n20466) );
  AOI21_X1 U23549 ( .B1(n20276), .B2(n20466), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20467) );
  INV_X1 U23550 ( .A(n20478), .ZN(n20525) );
  OAI22_X1 U23551 ( .A1(n20528), .A2(n20469), .B1(n20468), .B2(n20525), .ZN(
        n20470) );
  INV_X1 U23552 ( .A(n20470), .ZN(n20481) );
  NAND2_X1 U23553 ( .A1(n20472), .A2(n20471), .ZN(n20475) );
  AOI21_X1 U23554 ( .B1(n20475), .B2(n20474), .A(n20473), .ZN(n20477) );
  OAI211_X1 U23555 ( .C1(n20478), .C2(n20276), .A(n20477), .B(n20476), .ZN(
        n20531) );
  AOI22_X1 U23556 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20531), .B1(
        n10554), .B2(n20479), .ZN(n20480) );
  OAI211_X1 U23557 ( .C1(n20482), .C2(n20534), .A(n20481), .B(n20480), .ZN(
        P2_U3168) );
  OAI22_X1 U23558 ( .A1(n20528), .A2(n20484), .B1(n20483), .B2(n20525), .ZN(
        n20485) );
  INV_X1 U23559 ( .A(n20485), .ZN(n20488) );
  AOI22_X1 U23560 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20531), .B1(
        n10554), .B2(n20486), .ZN(n20487) );
  OAI211_X1 U23561 ( .C1(n20489), .C2(n20534), .A(n20488), .B(n20487), .ZN(
        P2_U3169) );
  OAI22_X1 U23562 ( .A1(n20528), .A2(n20491), .B1(n20490), .B2(n20525), .ZN(
        n20492) );
  INV_X1 U23563 ( .A(n20492), .ZN(n20495) );
  AOI22_X1 U23564 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20531), .B1(
        n10554), .B2(n20493), .ZN(n20494) );
  OAI211_X1 U23565 ( .C1(n20496), .C2(n20534), .A(n20495), .B(n20494), .ZN(
        P2_U3170) );
  OAI22_X1 U23566 ( .A1(n20528), .A2(n20498), .B1(n20497), .B2(n20525), .ZN(
        n20499) );
  INV_X1 U23567 ( .A(n20499), .ZN(n20502) );
  AOI22_X1 U23568 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20531), .B1(
        n10554), .B2(n20500), .ZN(n20501) );
  OAI211_X1 U23569 ( .C1(n20503), .C2(n20534), .A(n20502), .B(n20501), .ZN(
        P2_U3171) );
  OAI22_X1 U23570 ( .A1(n20528), .A2(n20505), .B1(n20504), .B2(n20525), .ZN(
        n20506) );
  INV_X1 U23571 ( .A(n20506), .ZN(n20509) );
  AOI22_X1 U23572 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20531), .B1(
        n10554), .B2(n20507), .ZN(n20508) );
  OAI211_X1 U23573 ( .C1(n20510), .C2(n20534), .A(n20509), .B(n20508), .ZN(
        P2_U3172) );
  OAI22_X1 U23574 ( .A1(n20528), .A2(n20512), .B1(n20511), .B2(n20525), .ZN(
        n20513) );
  INV_X1 U23575 ( .A(n20513), .ZN(n20516) );
  AOI22_X1 U23576 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20531), .B1(
        n10554), .B2(n20514), .ZN(n20515) );
  OAI211_X1 U23577 ( .C1(n20517), .C2(n20534), .A(n20516), .B(n20515), .ZN(
        P2_U3173) );
  OAI22_X1 U23578 ( .A1(n20528), .A2(n20519), .B1(n20518), .B2(n20525), .ZN(
        n20520) );
  INV_X1 U23579 ( .A(n20520), .ZN(n20523) );
  AOI22_X1 U23580 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20531), .B1(
        n10554), .B2(n20521), .ZN(n20522) );
  OAI211_X1 U23581 ( .C1(n20524), .C2(n20534), .A(n20523), .B(n20522), .ZN(
        P2_U3174) );
  OAI22_X1 U23582 ( .A1(n20528), .A2(n20527), .B1(n20526), .B2(n20525), .ZN(
        n20529) );
  INV_X1 U23583 ( .A(n20529), .ZN(n20533) );
  AOI22_X1 U23584 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20531), .B1(
        n10554), .B2(n20530), .ZN(n20532) );
  OAI211_X1 U23585 ( .C1(n20535), .C2(n20534), .A(n20533), .B(n20532), .ZN(
        P2_U3175) );
  OAI211_X1 U23586 ( .C1(n20537), .C2(n20536), .A(n20539), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20544) );
  NOR3_X1 U23587 ( .A1(n20690), .A2(n20539), .A3(n20538), .ZN(n20541) );
  OAI21_X1 U23588 ( .B1(n20542), .B2(n20541), .A(n20540), .ZN(n20543) );
  NAND3_X1 U23589 ( .A1(n20545), .A2(n20544), .A3(n20543), .ZN(P2_U3177) );
  NOR2_X1 U23590 ( .A1(n21336), .A2(n20627), .ZN(P2_U3179) );
  AND2_X1 U23591 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20546), .ZN(
        P2_U3180) );
  AND2_X1 U23592 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20546), .ZN(
        P2_U3181) );
  NOR2_X1 U23593 ( .A1(n21455), .A2(n20627), .ZN(P2_U3182) );
  AND2_X1 U23594 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20546), .ZN(
        P2_U3183) );
  AND2_X1 U23595 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20546), .ZN(
        P2_U3184) );
  AND2_X1 U23596 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20546), .ZN(
        P2_U3185) );
  AND2_X1 U23597 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20546), .ZN(
        P2_U3186) );
  AND2_X1 U23598 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20546), .ZN(
        P2_U3187) );
  AND2_X1 U23599 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20546), .ZN(
        P2_U3188) );
  AND2_X1 U23600 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20546), .ZN(
        P2_U3189) );
  AND2_X1 U23601 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20546), .ZN(
        P2_U3190) );
  AND2_X1 U23602 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20546), .ZN(
        P2_U3191) );
  AND2_X1 U23603 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20546), .ZN(
        P2_U3192) );
  AND2_X1 U23604 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20546), .ZN(
        P2_U3193) );
  AND2_X1 U23605 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20546), .ZN(
        P2_U3194) );
  AND2_X1 U23606 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20546), .ZN(
        P2_U3195) );
  AND2_X1 U23607 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20546), .ZN(
        P2_U3196) );
  AND2_X1 U23608 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20546), .ZN(
        P2_U3197) );
  AND2_X1 U23609 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20546), .ZN(
        P2_U3198) );
  AND2_X1 U23610 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20546), .ZN(
        P2_U3199) );
  AND2_X1 U23611 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20546), .ZN(
        P2_U3200) );
  AND2_X1 U23612 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20546), .ZN(P2_U3201) );
  AND2_X1 U23613 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20546), .ZN(P2_U3202) );
  AND2_X1 U23614 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20546), .ZN(P2_U3203) );
  AND2_X1 U23615 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20546), .ZN(P2_U3204) );
  AND2_X1 U23616 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20546), .ZN(P2_U3205) );
  AND2_X1 U23617 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20546), .ZN(P2_U3206) );
  AND2_X1 U23618 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20546), .ZN(P2_U3207) );
  AND2_X1 U23619 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20546), .ZN(P2_U3208) );
  NOR2_X1 U23620 ( .A1(n20686), .A2(n21404), .ZN(n20557) );
  INV_X1 U23621 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20558) );
  NOR3_X1 U23622 ( .A1(n20557), .A2(n20558), .A3(n20562), .ZN(n20550) );
  OAI211_X1 U23623 ( .C1(HOLD), .C2(n20558), .A(n20700), .B(n20547), .ZN(
        n20549) );
  INV_X1 U23624 ( .A(NA), .ZN(n21213) );
  NOR2_X1 U23625 ( .A1(n21213), .A2(n20552), .ZN(n20564) );
  INV_X1 U23626 ( .A(n20564), .ZN(n20548) );
  OAI211_X1 U23627 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n20550), .A(n20549), 
        .B(n20548), .ZN(P2_U3209) );
  NAND2_X1 U23628 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20556), .ZN(n20551) );
  AOI21_X1 U23629 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n20551), .A(n20558), 
        .ZN(n20553) );
  AOI211_X1 U23630 ( .C1(n20553), .C2(n20552), .A(n20692), .B(n20557), .ZN(
        n20554) );
  OAI21_X1 U23631 ( .B1(n20556), .B2(n20555), .A(n20554), .ZN(P2_U3210) );
  NOR3_X1 U23632 ( .A1(HOLD), .A2(n20557), .A3(n20562), .ZN(n20563) );
  NOR2_X1 U23633 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(HOLD), .ZN(n20561)
         );
  AOI22_X1 U23634 ( .A1(n20559), .A2(n20558), .B1(n20557), .B2(n21213), .ZN(
        n20560) );
  OAI33_X1 U23635 ( .A1(n20565), .A2(n20564), .A3(n20563), .B1(n20562), .B2(
        n20561), .B3(n20560), .ZN(P2_U3211) );
  OAI222_X1 U23636 ( .A1(n20615), .A2(n20567), .B1(n20566), .B2(n20699), .C1(
        n20569), .C2(n20614), .ZN(P2_U3212) );
  OAI222_X1 U23637 ( .A1(n20615), .A2(n20569), .B1(n20568), .B2(n20699), .C1(
        n20571), .C2(n20614), .ZN(P2_U3213) );
  OAI222_X1 U23638 ( .A1(n20615), .A2(n20571), .B1(n20570), .B2(n20699), .C1(
        n11319), .C2(n20614), .ZN(P2_U3214) );
  OAI222_X1 U23639 ( .A1(n20614), .A2(n11324), .B1(n20572), .B2(n20699), .C1(
        n11319), .C2(n20615), .ZN(P2_U3215) );
  OAI222_X1 U23640 ( .A1(n20614), .A2(n20574), .B1(n20573), .B2(n20699), .C1(
        n11324), .C2(n20615), .ZN(P2_U3216) );
  OAI222_X1 U23641 ( .A1(n20614), .A2(n20576), .B1(n20575), .B2(n20699), .C1(
        n20574), .C2(n20615), .ZN(P2_U3217) );
  OAI222_X1 U23642 ( .A1(n20614), .A2(n16490), .B1(n20577), .B2(n20699), .C1(
        n20576), .C2(n20615), .ZN(P2_U3218) );
  OAI222_X1 U23643 ( .A1(n20614), .A2(n20579), .B1(n20578), .B2(n20699), .C1(
        n16490), .C2(n20615), .ZN(P2_U3219) );
  OAI222_X1 U23644 ( .A1(n20614), .A2(n20581), .B1(n20580), .B2(n20699), .C1(
        n20579), .C2(n20615), .ZN(P2_U3220) );
  OAI222_X1 U23645 ( .A1(n20614), .A2(n20583), .B1(n20582), .B2(n20699), .C1(
        n20581), .C2(n20615), .ZN(P2_U3221) );
  OAI222_X1 U23646 ( .A1(n20614), .A2(n16440), .B1(n20584), .B2(n20699), .C1(
        n20583), .C2(n20615), .ZN(P2_U3222) );
  OAI222_X1 U23647 ( .A1(n20614), .A2(n16427), .B1(n20585), .B2(n20699), .C1(
        n16440), .C2(n20615), .ZN(P2_U3223) );
  OAI222_X1 U23648 ( .A1(n20614), .A2(n20587), .B1(n20586), .B2(n20699), .C1(
        n16427), .C2(n20615), .ZN(P2_U3224) );
  OAI222_X1 U23649 ( .A1(n20614), .A2(n20589), .B1(n20588), .B2(n20699), .C1(
        n20587), .C2(n20615), .ZN(P2_U3225) );
  OAI222_X1 U23650 ( .A1(n20614), .A2(n20591), .B1(n20590), .B2(n20699), .C1(
        n20589), .C2(n20615), .ZN(P2_U3226) );
  OAI222_X1 U23651 ( .A1(n20614), .A2(n20593), .B1(n20592), .B2(n20699), .C1(
        n20591), .C2(n20615), .ZN(P2_U3227) );
  INV_X1 U23652 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20594) );
  OAI222_X1 U23653 ( .A1(n20614), .A2(n20594), .B1(n21415), .B2(n20699), .C1(
        n20593), .C2(n20615), .ZN(P2_U3228) );
  OAI222_X1 U23654 ( .A1(n20614), .A2(n20596), .B1(n20595), .B2(n20699), .C1(
        n20594), .C2(n20615), .ZN(P2_U3229) );
  OAI222_X1 U23655 ( .A1(n20614), .A2(n14405), .B1(n20597), .B2(n20699), .C1(
        n20596), .C2(n20615), .ZN(P2_U3230) );
  OAI222_X1 U23656 ( .A1(n20614), .A2(n20599), .B1(n20598), .B2(n20699), .C1(
        n14405), .C2(n20615), .ZN(P2_U3231) );
  OAI222_X1 U23657 ( .A1(n20614), .A2(n16371), .B1(n20600), .B2(n20699), .C1(
        n20599), .C2(n20615), .ZN(P2_U3232) );
  OAI222_X1 U23658 ( .A1(n20614), .A2(n20601), .B1(n21432), .B2(n20699), .C1(
        n16371), .C2(n20615), .ZN(P2_U3233) );
  INV_X1 U23659 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20603) );
  OAI222_X1 U23660 ( .A1(n20614), .A2(n20603), .B1(n20602), .B2(n20699), .C1(
        n20601), .C2(n20615), .ZN(P2_U3234) );
  OAI222_X1 U23661 ( .A1(n20614), .A2(n20605), .B1(n20604), .B2(n20699), .C1(
        n20603), .C2(n20615), .ZN(P2_U3235) );
  OAI222_X1 U23662 ( .A1(n20614), .A2(n20607), .B1(n20606), .B2(n20699), .C1(
        n20605), .C2(n20615), .ZN(P2_U3236) );
  OAI222_X1 U23663 ( .A1(n20614), .A2(n20610), .B1(n20608), .B2(n20699), .C1(
        n20607), .C2(n20615), .ZN(P2_U3237) );
  OAI222_X1 U23664 ( .A1(n20615), .A2(n20610), .B1(n20609), .B2(n20699), .C1(
        n15787), .C2(n20614), .ZN(P2_U3238) );
  OAI222_X1 U23665 ( .A1(n20614), .A2(n20612), .B1(n20611), .B2(n20699), .C1(
        n15787), .C2(n20615), .ZN(P2_U3239) );
  OAI222_X1 U23666 ( .A1(n20614), .A2(n20616), .B1(n20613), .B2(n20699), .C1(
        n20612), .C2(n20615), .ZN(P2_U3240) );
  OAI222_X1 U23667 ( .A1(n20614), .A2(n20618), .B1(n20617), .B2(n20699), .C1(
        n20616), .C2(n20615), .ZN(P2_U3241) );
  INV_X1 U23668 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20619) );
  AOI22_X1 U23669 ( .A1(n20699), .A2(n20620), .B1(n20619), .B2(n20700), .ZN(
        P2_U3585) );
  INV_X1 U23670 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21429) );
  INV_X1 U23671 ( .A(P2_BE_N_REG_2__SCAN_IN), .ZN(n20621) );
  AOI22_X1 U23672 ( .A1(n20699), .A2(n21429), .B1(n20621), .B2(n20700), .ZN(
        P2_U3586) );
  MUX2_X1 U23673 ( .A(P2_BE_N_REG_1__SCAN_IN), .B(P2_BYTEENABLE_REG_1__SCAN_IN), .S(n20699), .Z(P2_U3587) );
  INV_X1 U23674 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20622) );
  AOI22_X1 U23675 ( .A1(n20699), .A2(n20623), .B1(n20622), .B2(n20700), .ZN(
        P2_U3588) );
  OAI21_X1 U23676 ( .B1(n20627), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20625), 
        .ZN(n20624) );
  INV_X1 U23677 ( .A(n20624), .ZN(P2_U3591) );
  OAI21_X1 U23678 ( .B1(n20627), .B2(n20626), .A(n20625), .ZN(P2_U3592) );
  INV_X1 U23679 ( .A(n20665), .ZN(n20668) );
  OR2_X1 U23680 ( .A1(n20629), .A2(n20628), .ZN(n20639) );
  NAND2_X1 U23681 ( .A1(n20634), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20652) );
  OR2_X1 U23682 ( .A1(n20630), .A2(n20652), .ZN(n20649) );
  OR2_X1 U23683 ( .A1(n20632), .A2(n20631), .ZN(n20633) );
  AOI21_X1 U23684 ( .B1(n20655), .B2(n20634), .A(n20633), .ZN(n20644) );
  NAND2_X1 U23685 ( .A1(n20649), .A2(n20644), .ZN(n20636) );
  AOI22_X1 U23686 ( .A1(n20637), .A2(n20636), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20635), .ZN(n20638) );
  OAI21_X1 U23687 ( .B1(n20640), .B2(n20639), .A(n20638), .ZN(n20641) );
  INV_X1 U23688 ( .A(n20641), .ZN(n20642) );
  AOI22_X1 U23689 ( .A1(n20668), .A2(n20643), .B1(n20642), .B2(n20665), .ZN(
        P2_U3602) );
  INV_X1 U23690 ( .A(n20644), .ZN(n20646) );
  AOI22_X1 U23691 ( .A1(n20647), .A2(n20646), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20645), .ZN(n20648) );
  AND2_X1 U23692 ( .A1(n20649), .A2(n20648), .ZN(n20650) );
  AOI22_X1 U23693 ( .A1(n20668), .A2(n20651), .B1(n20650), .B2(n20665), .ZN(
        P2_U3603) );
  INV_X1 U23694 ( .A(n20652), .ZN(n20654) );
  AOI22_X1 U23695 ( .A1(n20655), .A2(n20654), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20653), .ZN(n20658) );
  NAND3_X1 U23696 ( .A1(n20656), .A2(n20663), .A3(n10551), .ZN(n20657) );
  AND2_X1 U23697 ( .A1(n20658), .A2(n20657), .ZN(n20659) );
  AOI22_X1 U23698 ( .A1(n20668), .A2(n20660), .B1(n20659), .B2(n20665), .ZN(
        P2_U3604) );
  AOI211_X1 U23699 ( .C1(n20664), .C2(n20663), .A(n20662), .B(n20661), .ZN(
        n20666) );
  AOI22_X1 U23700 ( .A1(n20668), .A2(n20667), .B1(n20666), .B2(n20665), .ZN(
        P2_U3605) );
  INV_X1 U23701 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20669) );
  AOI22_X1 U23702 ( .A1(n20699), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20669), 
        .B2(n20700), .ZN(P2_U3608) );
  INV_X1 U23703 ( .A(n20670), .ZN(n20677) );
  INV_X1 U23704 ( .A(n20671), .ZN(n20676) );
  INV_X1 U23705 ( .A(n20672), .ZN(n20673) );
  NAND2_X1 U23706 ( .A1(n20674), .A2(n20673), .ZN(n20675) );
  OAI211_X1 U23707 ( .C1(n20678), .C2(n20677), .A(n20676), .B(n20675), .ZN(
        n20680) );
  MUX2_X1 U23708 ( .A(P2_MORE_REG_SCAN_IN), .B(n20680), .S(n20679), .Z(
        P2_U3609) );
  AOI21_X1 U23709 ( .B1(n20681), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20684) );
  INV_X1 U23710 ( .A(n20682), .ZN(n20683) );
  AOI211_X1 U23711 ( .C1(n20686), .C2(n20685), .A(n20684), .B(n20683), .ZN(
        n20698) );
  NAND2_X1 U23712 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n20686), .ZN(n20694) );
  NAND2_X1 U23713 ( .A1(n20688), .A2(n20687), .ZN(n20691) );
  AOI211_X1 U23714 ( .C1(n20692), .C2(n20691), .A(n20690), .B(n20689), .ZN(
        n20693) );
  AOI21_X1 U23715 ( .B1(n20695), .B2(n20694), .A(n20693), .ZN(n20697) );
  NAND2_X1 U23716 ( .A1(n20698), .A2(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20696) );
  OAI21_X1 U23717 ( .B1(n20698), .B2(n20697), .A(n20696), .ZN(P2_U3610) );
  OAI22_X1 U23718 ( .A1(n20700), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20699), .ZN(n20701) );
  INV_X1 U23719 ( .A(n20701), .ZN(P2_U3611) );
  OAI21_X1 U23720 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20702), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n21214) );
  OR2_X2 U23721 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20702), .ZN(n21303) );
  OAI21_X1 U23722 ( .B1(n21214), .B2(P1_ADS_N_REG_SCAN_IN), .A(n21303), .ZN(
        n20703) );
  INV_X1 U23723 ( .A(n20703), .ZN(P1_U2802) );
  OAI21_X1 U23724 ( .B1(n20704), .B2(n20710), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20705) );
  OAI21_X1 U23725 ( .B1(n20706), .B2(n11759), .A(n20705), .ZN(P1_U2803) );
  NOR2_X1 U23726 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20708) );
  OAI21_X1 U23727 ( .B1(n20708), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21303), .ZN(
        n20707) );
  OAI21_X1 U23728 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21303), .A(n20707), 
        .ZN(P1_U2804) );
  AND2_X1 U23729 ( .A1(n21214), .A2(n21303), .ZN(n21288) );
  OAI21_X1 U23730 ( .B1(BS16), .B2(n20708), .A(n21288), .ZN(n21286) );
  OAI21_X1 U23731 ( .B1(n21288), .B2(n20709), .A(n21286), .ZN(P1_U2805) );
  NOR2_X1 U23732 ( .A1(n20711), .A2(n20710), .ZN(n21308) );
  INV_X1 U23733 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20713) );
  OAI21_X1 U23734 ( .B1(n21308), .B2(n20713), .A(n20712), .ZN(P1_U2806) );
  NOR4_X1 U23735 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20717) );
  NOR4_X1 U23736 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20716) );
  NOR4_X1 U23737 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20715) );
  NOR4_X1 U23738 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20714) );
  NAND4_X1 U23739 ( .A1(n20717), .A2(n20716), .A3(n20715), .A4(n20714), .ZN(
        n20723) );
  NOR4_X1 U23740 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20721) );
  AOI211_X1 U23741 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20720) );
  NOR4_X1 U23742 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20719) );
  NOR4_X1 U23743 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20718) );
  NAND4_X1 U23744 ( .A1(n20721), .A2(n20720), .A3(n20719), .A4(n20718), .ZN(
        n20722) );
  NOR2_X1 U23745 ( .A1(n20723), .A2(n20722), .ZN(n21302) );
  INV_X1 U23746 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21281) );
  NOR3_X1 U23747 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20725) );
  OAI21_X1 U23748 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20725), .A(n21302), .ZN(
        n20724) );
  OAI21_X1 U23749 ( .B1(n21302), .B2(n21281), .A(n20724), .ZN(P1_U2807) );
  INV_X1 U23750 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20726) );
  INV_X1 U23751 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21287) );
  AOI21_X1 U23752 ( .B1(n20726), .B2(n21287), .A(n20725), .ZN(n20727) );
  INV_X1 U23753 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21278) );
  INV_X1 U23754 ( .A(n21302), .ZN(n21299) );
  AOI22_X1 U23755 ( .A1(n21302), .A2(n20727), .B1(n21278), .B2(n21299), .ZN(
        P1_U2808) );
  NAND2_X1 U23756 ( .A1(n20729), .A2(n20728), .ZN(n20741) );
  INV_X1 U23757 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20732) );
  INV_X1 U23758 ( .A(n20730), .ZN(n20731) );
  OAI22_X1 U23759 ( .A1(n20732), .A2(n20781), .B1(n20780), .B2(n20731), .ZN(
        n20733) );
  AOI211_X1 U23760 ( .C1(n20785), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n20772), .B(n20733), .ZN(n20734) );
  OAI221_X1 U23761 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n20735), .C1(n21233), 
        .C2(n20741), .A(n20734), .ZN(n20736) );
  AOI21_X1 U23762 ( .B1(n12954), .B2(n20737), .A(n20736), .ZN(n20738) );
  OAI21_X1 U23763 ( .B1(n20739), .B2(n12914), .A(n20738), .ZN(P1_U2833) );
  INV_X1 U23764 ( .A(n20764), .ZN(n20740) );
  INV_X1 U23765 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21229) );
  NOR2_X1 U23766 ( .A1(n20740), .A2(n21229), .ZN(n20743) );
  INV_X1 U23767 ( .A(n20741), .ZN(n20742) );
  MUX2_X1 U23768 ( .A(n20743), .B(n20742), .S(P1_REIP_REG_6__SCAN_IN), .Z(
        n20752) );
  INV_X1 U23769 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n20744) );
  OAI21_X1 U23770 ( .B1(n20762), .B2(n20744), .A(n20759), .ZN(n20745) );
  AOI21_X1 U23771 ( .B1(n20757), .B2(P1_EBX_REG_6__SCAN_IN), .A(n20745), .ZN(
        n20748) );
  NAND2_X1 U23772 ( .A1(n20758), .A2(n20746), .ZN(n20747) );
  OAI211_X1 U23773 ( .C1(n20750), .C2(n20749), .A(n20748), .B(n20747), .ZN(
        n20751) );
  NOR2_X1 U23774 ( .A1(n20752), .A2(n20751), .ZN(n20753) );
  OAI21_X1 U23775 ( .B1(n20754), .B2(n12914), .A(n20753), .ZN(P1_U2834) );
  AOI22_X1 U23776 ( .A1(n20758), .A2(n20794), .B1(n20757), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n20760) );
  OAI211_X1 U23777 ( .C1(n20762), .C2(n20761), .A(n20760), .B(n20759), .ZN(
        n20763) );
  AOI221_X1 U23778 ( .B1(n20764), .B2(n21229), .C1(n9643), .C2(
        P1_REIP_REG_5__SCAN_IN), .A(n20763), .ZN(n20766) );
  NAND2_X1 U23779 ( .A1(n20797), .A2(n20792), .ZN(n20765) );
  OAI211_X1 U23780 ( .C1(n12914), .C2(n20767), .A(n20766), .B(n20765), .ZN(
        P1_U2835) );
  INV_X1 U23781 ( .A(n20786), .ZN(n20770) );
  OAI222_X1 U23782 ( .A1(n20894), .A2(n20780), .B1(n20770), .B2(n20769), .C1(
        n20768), .C2(n20781), .ZN(n20771) );
  AOI211_X1 U23783 ( .C1(n20785), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20772), .B(n20771), .ZN(n20776) );
  NAND2_X1 U23784 ( .A1(n21226), .A2(n20773), .ZN(n20774) );
  AOI22_X1 U23785 ( .A1(n9643), .A2(n20774), .B1(n20861), .B2(n20792), .ZN(
        n20775) );
  OAI211_X1 U23786 ( .C1(n20864), .C2(n12914), .A(n20776), .B(n20775), .ZN(
        P1_U2836) );
  INV_X1 U23787 ( .A(n20777), .ZN(n20885) );
  INV_X1 U23788 ( .A(n20778), .ZN(n20779) );
  OAI22_X1 U23789 ( .A1(n20782), .A2(n20781), .B1(n20780), .B2(n20779), .ZN(
        n20791) );
  INV_X1 U23790 ( .A(n20783), .ZN(n20789) );
  AOI22_X1 U23791 ( .A1(n20785), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20784), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n20788) );
  NAND2_X1 U23792 ( .A1(n20786), .A2(n21092), .ZN(n20787) );
  OAI211_X1 U23793 ( .C1(n20789), .C2(P1_REIP_REG_1__SCAN_IN), .A(n20788), .B(
        n20787), .ZN(n20790) );
  AOI211_X1 U23794 ( .C1(n20792), .C2(n20885), .A(n20791), .B(n20790), .ZN(
        n20793) );
  OAI21_X1 U23795 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n12914), .A(
        n20793), .ZN(P1_U2839) );
  INV_X1 U23796 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20799) );
  AOI22_X1 U23797 ( .A1(n20797), .A2(n20796), .B1(n20795), .B2(n20794), .ZN(
        n20798) );
  OAI21_X1 U23798 ( .B1(n20800), .B2(n20799), .A(n20798), .ZN(P1_U2867) );
  AOI22_X1 U23799 ( .A1(n20824), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20802) );
  OAI21_X1 U23800 ( .B1(n20803), .B2(n20826), .A(n20802), .ZN(P1_U2921) );
  AOI22_X1 U23801 ( .A1(n20824), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20804) );
  OAI21_X1 U23802 ( .B1(n15152), .B2(n20826), .A(n20804), .ZN(P1_U2922) );
  INV_X1 U23803 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20853) );
  AOI22_X1 U23804 ( .A1(n20824), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20805) );
  OAI21_X1 U23805 ( .B1(n20853), .B2(n20826), .A(n20805), .ZN(P1_U2923) );
  AOI22_X1 U23806 ( .A1(n20824), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20806) );
  OAI21_X1 U23807 ( .B1(n15158), .B2(n20826), .A(n20806), .ZN(P1_U2924) );
  AOI22_X1 U23808 ( .A1(n20824), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20807) );
  OAI21_X1 U23809 ( .B1(n20808), .B2(n20826), .A(n20807), .ZN(P1_U2925) );
  INV_X1 U23810 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20848) );
  AOI22_X1 U23811 ( .A1(n20824), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20809) );
  OAI21_X1 U23812 ( .B1(n20848), .B2(n20826), .A(n20809), .ZN(P1_U2926) );
  AOI22_X1 U23813 ( .A1(n20824), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20810) );
  OAI21_X1 U23814 ( .B1(n14278), .B2(n20826), .A(n20810), .ZN(P1_U2927) );
  AOI22_X1 U23815 ( .A1(n20824), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20811) );
  OAI21_X1 U23816 ( .B1(n21438), .B2(n20826), .A(n20811), .ZN(P1_U2928) );
  AOI22_X1 U23817 ( .A1(n20824), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20812) );
  OAI21_X1 U23818 ( .B1(n11974), .B2(n20826), .A(n20812), .ZN(P1_U2929) );
  AOI22_X1 U23819 ( .A1(n20824), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20813) );
  OAI21_X1 U23820 ( .B1(n11965), .B2(n20826), .A(n20813), .ZN(P1_U2930) );
  AOI22_X1 U23821 ( .A1(n20824), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20815) );
  OAI21_X1 U23822 ( .B1(n14160), .B2(n20826), .A(n20815), .ZN(P1_U2931) );
  AOI22_X1 U23823 ( .A1(n20824), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20816) );
  OAI21_X1 U23824 ( .B1(n20817), .B2(n20826), .A(n20816), .ZN(P1_U2932) );
  AOI22_X1 U23825 ( .A1(n20824), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20818) );
  OAI21_X1 U23826 ( .B1(n20819), .B2(n20826), .A(n20818), .ZN(P1_U2933) );
  AOI22_X1 U23827 ( .A1(n20824), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20820) );
  OAI21_X1 U23828 ( .B1(n20821), .B2(n20826), .A(n20820), .ZN(P1_U2934) );
  AOI22_X1 U23829 ( .A1(n20824), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20822) );
  OAI21_X1 U23830 ( .B1(n20823), .B2(n20826), .A(n20822), .ZN(P1_U2935) );
  AOI22_X1 U23831 ( .A1(n20824), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20814), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20825) );
  OAI21_X1 U23832 ( .B1(n20827), .B2(n20826), .A(n20825), .ZN(P1_U2936) );
  NOR2_X1 U23833 ( .A1(n20842), .A2(n20828), .ZN(n20844) );
  AOI21_X1 U23834 ( .B1(P1_UWORD_REG_9__SCAN_IN), .B2(n13702), .A(n20844), 
        .ZN(n20829) );
  OAI21_X1 U23835 ( .B1(n20830), .B2(n20856), .A(n20829), .ZN(P1_U2946) );
  INV_X1 U23836 ( .A(n20831), .ZN(n20832) );
  NOR2_X1 U23837 ( .A1(n20842), .A2(n20832), .ZN(n20846) );
  AOI21_X1 U23838 ( .B1(P1_UWORD_REG_10__SCAN_IN), .B2(n13702), .A(n20846), 
        .ZN(n20833) );
  OAI21_X1 U23839 ( .B1(n12386), .B2(n20856), .A(n20833), .ZN(P1_U2947) );
  NOR2_X1 U23840 ( .A1(n20842), .A2(n20834), .ZN(n20849) );
  AOI21_X1 U23841 ( .B1(P1_UWORD_REG_12__SCAN_IN), .B2(n13702), .A(n20849), 
        .ZN(n20835) );
  OAI21_X1 U23842 ( .B1(n20836), .B2(n20856), .A(n20835), .ZN(P1_U2949) );
  INV_X1 U23843 ( .A(n20837), .ZN(n20838) );
  NOR2_X1 U23844 ( .A1(n20842), .A2(n20838), .ZN(n20851) );
  AOI21_X1 U23845 ( .B1(P1_UWORD_REG_13__SCAN_IN), .B2(n13702), .A(n20851), 
        .ZN(n20839) );
  OAI21_X1 U23846 ( .B1(n20840), .B2(n20856), .A(n20839), .ZN(P1_U2950) );
  NOR2_X1 U23847 ( .A1(n20842), .A2(n20841), .ZN(n20854) );
  AOI21_X1 U23848 ( .B1(P1_UWORD_REG_14__SCAN_IN), .B2(n13702), .A(n20854), 
        .ZN(n20843) );
  OAI21_X1 U23849 ( .B1(n15073), .B2(n20856), .A(n20843), .ZN(P1_U2951) );
  AOI21_X1 U23850 ( .B1(P1_LWORD_REG_9__SCAN_IN), .B2(n13702), .A(n20844), 
        .ZN(n20845) );
  OAI21_X1 U23851 ( .B1(n14278), .B2(n20856), .A(n20845), .ZN(P1_U2961) );
  AOI21_X1 U23852 ( .B1(P1_LWORD_REG_10__SCAN_IN), .B2(n13702), .A(n20846), 
        .ZN(n20847) );
  OAI21_X1 U23853 ( .B1(n20848), .B2(n20856), .A(n20847), .ZN(P1_U2962) );
  AOI21_X1 U23854 ( .B1(P1_LWORD_REG_12__SCAN_IN), .B2(n13702), .A(n20849), 
        .ZN(n20850) );
  OAI21_X1 U23855 ( .B1(n15158), .B2(n20856), .A(n20850), .ZN(P1_U2964) );
  AOI21_X1 U23856 ( .B1(P1_LWORD_REG_13__SCAN_IN), .B2(n13702), .A(n20851), 
        .ZN(n20852) );
  OAI21_X1 U23857 ( .B1(n20853), .B2(n20856), .A(n20852), .ZN(P1_U2965) );
  AOI21_X1 U23858 ( .B1(P1_LWORD_REG_14__SCAN_IN), .B2(n13702), .A(n20854), 
        .ZN(n20855) );
  OAI21_X1 U23859 ( .B1(n15152), .B2(n20856), .A(n20855), .ZN(P1_U2966) );
  AOI22_X1 U23860 ( .A1(n20882), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20916), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20863) );
  OAI21_X1 U23861 ( .B1(n20859), .B2(n20858), .A(n20857), .ZN(n20860) );
  INV_X1 U23862 ( .A(n20860), .ZN(n20898) );
  AOI22_X1 U23863 ( .A1(n20884), .A2(n20861), .B1(n20898), .B2(n20887), .ZN(
        n20862) );
  OAI211_X1 U23864 ( .C1(n20881), .C2(n20864), .A(n20863), .B(n20862), .ZN(
        P1_U2995) );
  AOI22_X1 U23865 ( .A1(n20882), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20916), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n20871) );
  OAI21_X1 U23866 ( .B1(n20867), .B2(n20866), .A(n20865), .ZN(n20868) );
  INV_X1 U23867 ( .A(n20868), .ZN(n20905) );
  AOI22_X1 U23868 ( .A1(n20869), .A2(n20884), .B1(n20905), .B2(n20887), .ZN(
        n20870) );
  OAI211_X1 U23869 ( .C1(n20881), .C2(n20872), .A(n20871), .B(n20870), .ZN(
        P1_U2996) );
  AOI22_X1 U23870 ( .A1(n20882), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20916), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n20879) );
  OAI21_X1 U23871 ( .B1(n20875), .B2(n20874), .A(n20873), .ZN(n20876) );
  INV_X1 U23872 ( .A(n20876), .ZN(n20923) );
  AOI22_X1 U23873 ( .A1(n20877), .A2(n20884), .B1(n20923), .B2(n20887), .ZN(
        n20878) );
  OAI211_X1 U23874 ( .C1(n20881), .C2(n20880), .A(n20879), .B(n20878), .ZN(
        P1_U2997) );
  AOI22_X1 U23875 ( .A1(n20882), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20916), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n20889) );
  INV_X1 U23876 ( .A(n20883), .ZN(n20886) );
  AOI22_X1 U23877 ( .A1(n20887), .A2(n20886), .B1(n20885), .B2(n20884), .ZN(
        n20888) );
  OAI211_X1 U23878 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20881), .A(
        n20889), .B(n20888), .ZN(P1_U2998) );
  AOI21_X1 U23879 ( .B1(n20891), .B2(n20914), .A(n20890), .ZN(n20909) );
  AOI211_X1 U23880 ( .C1(n20900), .C2(n20908), .A(n20892), .B(n20903), .ZN(
        n20897) );
  OAI22_X1 U23881 ( .A1(n20895), .A2(n20894), .B1(n21226), .B2(n20893), .ZN(
        n20896) );
  AOI211_X1 U23882 ( .C1(n20898), .C2(n20922), .A(n20897), .B(n20896), .ZN(
        n20899) );
  OAI21_X1 U23883 ( .B1(n20909), .B2(n20900), .A(n20899), .ZN(P1_U3027) );
  INV_X1 U23884 ( .A(n20901), .ZN(n20902) );
  AOI22_X1 U23885 ( .A1(n17191), .A2(n20902), .B1(n20916), .B2(
        P1_REIP_REG_3__SCAN_IN), .ZN(n20907) );
  INV_X1 U23886 ( .A(n20903), .ZN(n20904) );
  AOI22_X1 U23887 ( .A1(n20905), .A2(n20922), .B1(n20908), .B2(n20904), .ZN(
        n20906) );
  OAI211_X1 U23888 ( .C1(n20909), .C2(n20908), .A(n20907), .B(n20906), .ZN(
        P1_U3028) );
  NAND2_X1 U23889 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20910), .ZN(
        n20927) );
  AOI21_X1 U23890 ( .B1(n20913), .B2(n20912), .A(n20911), .ZN(n20925) );
  AOI21_X1 U23891 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n20915), .A(
        n20914), .ZN(n20919) );
  AOI22_X1 U23892 ( .A1(n17191), .A2(n20917), .B1(n20916), .B2(
        P1_REIP_REG_2__SCAN_IN), .ZN(n20918) );
  OAI21_X1 U23893 ( .B1(n20920), .B2(n20919), .A(n20918), .ZN(n20921) );
  AOI21_X1 U23894 ( .B1(n20923), .B2(n20922), .A(n20921), .ZN(n20924) );
  OAI221_X1 U23895 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20927), .C1(
        n20926), .C2(n20925), .A(n20924), .ZN(P1_U3029) );
  INV_X1 U23896 ( .A(n20928), .ZN(n20929) );
  NAND2_X1 U23897 ( .A1(n17191), .A2(n20929), .ZN(n20930) );
  OAI211_X1 U23898 ( .C1(n20933), .C2(n20932), .A(n20931), .B(n20930), .ZN(
        n20934) );
  INV_X1 U23899 ( .A(n20934), .ZN(n20940) );
  OAI21_X1 U23900 ( .B1(n20936), .B2(n20935), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20938) );
  NAND4_X1 U23901 ( .A1(n20940), .A2(n20939), .A3(n20938), .A4(n20937), .ZN(
        P1_U3031) );
  NOR2_X1 U23902 ( .A1(n20942), .A2(n20941), .ZN(P1_U3032) );
  AOI22_X1 U23903 ( .A1(n21138), .A2(n20952), .B1(n20951), .B2(n21150), .ZN(
        n20944) );
  AOI22_X1 U23904 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20954), .B1(
        n21139), .B2(n20953), .ZN(n20943) );
  OAI211_X1 U23905 ( .C1(n21153), .C2(n20972), .A(n20944), .B(n20943), .ZN(
        P1_U3057) );
  AOI22_X1 U23906 ( .A1(n21160), .A2(n20952), .B1(n20951), .B2(n21106), .ZN(
        n20946) );
  AOI22_X1 U23907 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20954), .B1(
        n21161), .B2(n20953), .ZN(n20945) );
  OAI211_X1 U23908 ( .C1(n21109), .C2(n20972), .A(n20946), .B(n20945), .ZN(
        P1_U3059) );
  AOI22_X1 U23909 ( .A1(n21172), .A2(n20952), .B1(n20951), .B2(n21114), .ZN(
        n20948) );
  AOI22_X1 U23910 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20954), .B1(
        n21173), .B2(n20953), .ZN(n20947) );
  OAI211_X1 U23911 ( .C1(n21117), .C2(n20972), .A(n20948), .B(n20947), .ZN(
        P1_U3061) );
  AOI22_X1 U23912 ( .A1(n21178), .A2(n20952), .B1(n20951), .B2(n21118), .ZN(
        n20950) );
  AOI22_X1 U23913 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20954), .B1(
        n21179), .B2(n20953), .ZN(n20949) );
  OAI211_X1 U23914 ( .C1(n21121), .C2(n20972), .A(n20950), .B(n20949), .ZN(
        P1_U3062) );
  AOI22_X1 U23915 ( .A1(n21193), .A2(n20952), .B1(n20951), .B2(n21126), .ZN(
        n20956) );
  AOI22_X1 U23916 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20954), .B1(
        n21195), .B2(n20953), .ZN(n20955) );
  OAI211_X1 U23917 ( .C1(n21131), .C2(n20972), .A(n20956), .B(n20955), .ZN(
        P1_U3064) );
  INV_X1 U23918 ( .A(n20957), .ZN(n20967) );
  AOI22_X1 U23919 ( .A1(n21139), .A2(n20967), .B1(n21138), .B2(n20966), .ZN(
        n20959) );
  AOI22_X1 U23920 ( .A1(n20969), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n20968), .B2(n21055), .ZN(n20958) );
  OAI211_X1 U23921 ( .C1(n21070), .C2(n20972), .A(n20959), .B(n20958), .ZN(
        P1_U3065) );
  AOI22_X1 U23922 ( .A1(n21155), .A2(n20967), .B1(n21154), .B2(n20966), .ZN(
        n20961) );
  AOI22_X1 U23923 ( .A1(n20969), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n20968), .B2(n21156), .ZN(n20960) );
  OAI211_X1 U23924 ( .C1(n21159), .C2(n20972), .A(n20961), .B(n20960), .ZN(
        P1_U3066) );
  AOI22_X1 U23925 ( .A1(n21167), .A2(n20967), .B1(n21166), .B2(n20966), .ZN(
        n20963) );
  AOI22_X1 U23926 ( .A1(n20969), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n20968), .B2(n21168), .ZN(n20962) );
  OAI211_X1 U23927 ( .C1(n21171), .C2(n20972), .A(n20963), .B(n20962), .ZN(
        P1_U3068) );
  AOI22_X1 U23928 ( .A1(n21185), .A2(n20967), .B1(n21184), .B2(n20966), .ZN(
        n20965) );
  AOI22_X1 U23929 ( .A1(n20969), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n20968), .B2(n21081), .ZN(n20964) );
  OAI211_X1 U23930 ( .C1(n21084), .C2(n20972), .A(n20965), .B(n20964), .ZN(
        P1_U3071) );
  AOI22_X1 U23931 ( .A1(n21195), .A2(n20967), .B1(n21193), .B2(n20966), .ZN(
        n20971) );
  AOI22_X1 U23932 ( .A1(n20969), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n20968), .B2(n21196), .ZN(n20970) );
  OAI211_X1 U23933 ( .C1(n21202), .C2(n20972), .A(n20971), .B(n20970), .ZN(
        P1_U3072) );
  AOI22_X1 U23934 ( .A1(n21139), .A2(n20986), .B1(n21138), .B2(n20985), .ZN(
        n20974) );
  AOI22_X1 U23935 ( .A1(n20988), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n20987), .B2(n21150), .ZN(n20973) );
  OAI211_X1 U23936 ( .C1(n21153), .C2(n21020), .A(n20974), .B(n20973), .ZN(
        P1_U3105) );
  AOI22_X1 U23937 ( .A1(n21155), .A2(n20986), .B1(n21154), .B2(n20985), .ZN(
        n20976) );
  AOI22_X1 U23938 ( .A1(n20988), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n20987), .B2(n21102), .ZN(n20975) );
  OAI211_X1 U23939 ( .C1(n21105), .C2(n21020), .A(n20976), .B(n20975), .ZN(
        P1_U3106) );
  AOI22_X1 U23940 ( .A1(n21161), .A2(n20986), .B1(n21160), .B2(n20985), .ZN(
        n20978) );
  AOI22_X1 U23941 ( .A1(n20988), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n20987), .B2(n21106), .ZN(n20977) );
  OAI211_X1 U23942 ( .C1(n21109), .C2(n21020), .A(n20978), .B(n20977), .ZN(
        P1_U3107) );
  AOI22_X1 U23943 ( .A1(n21167), .A2(n20986), .B1(n21166), .B2(n20985), .ZN(
        n20980) );
  AOI22_X1 U23944 ( .A1(n20988), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n20987), .B2(n21110), .ZN(n20979) );
  OAI211_X1 U23945 ( .C1(n21113), .C2(n21020), .A(n20980), .B(n20979), .ZN(
        P1_U3108) );
  AOI22_X1 U23946 ( .A1(n21173), .A2(n20986), .B1(n21172), .B2(n20985), .ZN(
        n20982) );
  AOI22_X1 U23947 ( .A1(n20988), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n20987), .B2(n21114), .ZN(n20981) );
  OAI211_X1 U23948 ( .C1(n21117), .C2(n21020), .A(n20982), .B(n20981), .ZN(
        P1_U3109) );
  AOI22_X1 U23949 ( .A1(n21185), .A2(n20986), .B1(n21184), .B2(n20985), .ZN(
        n20984) );
  AOI22_X1 U23950 ( .A1(n20988), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n20987), .B2(n21186), .ZN(n20983) );
  OAI211_X1 U23951 ( .C1(n21191), .C2(n21020), .A(n20984), .B(n20983), .ZN(
        P1_U3111) );
  AOI22_X1 U23952 ( .A1(n21195), .A2(n20986), .B1(n21193), .B2(n20985), .ZN(
        n20990) );
  AOI22_X1 U23953 ( .A1(n20988), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n20987), .B2(n21126), .ZN(n20989) );
  OAI211_X1 U23954 ( .C1(n21131), .C2(n21020), .A(n20990), .B(n20989), .ZN(
        P1_U3112) );
  NOR2_X1 U23955 ( .A1(n21136), .A2(n21021), .ZN(n21028) );
  INV_X1 U23956 ( .A(n21028), .ZN(n21023) );
  NOR2_X1 U23957 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21023), .ZN(
        n21015) );
  AOI22_X1 U23958 ( .A1(n21015), .A2(n21138), .B1(n21012), .B2(n21150), .ZN(
        n21001) );
  NAND3_X1 U23959 ( .A1(n21020), .A2(n21044), .A3(n21029), .ZN(n20991) );
  NAND2_X1 U23960 ( .A1(n20991), .A2(n21057), .ZN(n20996) );
  NAND2_X1 U23961 ( .A1(n21022), .A2(n21092), .ZN(n20998) );
  OR2_X1 U23962 ( .A1(n20992), .A2(n17089), .ZN(n21093) );
  NAND2_X1 U23963 ( .A1(n21093), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21097) );
  OAI211_X1 U23964 ( .C1(n21064), .C2(n21015), .A(n21097), .B(n20993), .ZN(
        n20994) );
  AOI21_X1 U23965 ( .B1(n20996), .B2(n20998), .A(n20994), .ZN(n20995) );
  INV_X1 U23966 ( .A(n20996), .ZN(n20999) );
  AOI22_X1 U23967 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n21017), .B1(
        n21139), .B2(n21016), .ZN(n21000) );
  OAI211_X1 U23968 ( .C1(n21153), .C2(n21044), .A(n21001), .B(n21000), .ZN(
        P1_U3113) );
  AOI22_X1 U23969 ( .A1(n21015), .A2(n21154), .B1(n21049), .B2(n21156), .ZN(
        n21003) );
  AOI22_X1 U23970 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n21017), .B1(
        n21155), .B2(n21016), .ZN(n21002) );
  OAI211_X1 U23971 ( .C1(n21159), .C2(n21020), .A(n21003), .B(n21002), .ZN(
        P1_U3114) );
  AOI22_X1 U23972 ( .A1(n21015), .A2(n21160), .B1(n21049), .B2(n21162), .ZN(
        n21005) );
  AOI22_X1 U23973 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n21017), .B1(
        n21161), .B2(n21016), .ZN(n21004) );
  OAI211_X1 U23974 ( .C1(n21165), .C2(n21020), .A(n21005), .B(n21004), .ZN(
        P1_U3115) );
  AOI22_X1 U23975 ( .A1(n21015), .A2(n21166), .B1(n21049), .B2(n21168), .ZN(
        n21007) );
  AOI22_X1 U23976 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n21017), .B1(
        n21167), .B2(n21016), .ZN(n21006) );
  OAI211_X1 U23977 ( .C1(n21171), .C2(n21020), .A(n21007), .B(n21006), .ZN(
        P1_U3116) );
  AOI22_X1 U23978 ( .A1(n21015), .A2(n21172), .B1(n21049), .B2(n21174), .ZN(
        n21009) );
  AOI22_X1 U23979 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n21017), .B1(
        n21173), .B2(n21016), .ZN(n21008) );
  OAI211_X1 U23980 ( .C1(n21177), .C2(n21020), .A(n21009), .B(n21008), .ZN(
        P1_U3117) );
  AOI22_X1 U23981 ( .A1(n21015), .A2(n21178), .B1(n21049), .B2(n21180), .ZN(
        n21011) );
  AOI22_X1 U23982 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n21017), .B1(
        n21179), .B2(n21016), .ZN(n21010) );
  OAI211_X1 U23983 ( .C1(n21183), .C2(n21020), .A(n21011), .B(n21010), .ZN(
        P1_U3118) );
  AOI22_X1 U23984 ( .A1(n21015), .A2(n21184), .B1(n21012), .B2(n21186), .ZN(
        n21014) );
  AOI22_X1 U23985 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n21017), .B1(
        n21185), .B2(n21016), .ZN(n21013) );
  OAI211_X1 U23986 ( .C1(n21191), .C2(n21044), .A(n21014), .B(n21013), .ZN(
        P1_U3119) );
  AOI22_X1 U23987 ( .A1(n21015), .A2(n21193), .B1(n21049), .B2(n21196), .ZN(
        n21019) );
  AOI22_X1 U23988 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n21017), .B1(
        n21195), .B2(n21016), .ZN(n21018) );
  OAI211_X1 U23989 ( .C1(n21202), .C2(n21020), .A(n21019), .B(n21018), .ZN(
        P1_U3120) );
  NOR2_X1 U23990 ( .A1(n21132), .A2(n21021), .ZN(n21047) );
  AOI21_X1 U23991 ( .B1(n21022), .B2(n21133), .A(n21047), .ZN(n21025) );
  OAI22_X1 U23992 ( .A1(n21025), .A2(n21141), .B1(n21023), .B2(n11830), .ZN(
        n21048) );
  AOI22_X1 U23993 ( .A1(n21139), .A2(n21048), .B1(n21138), .B2(n21047), .ZN(
        n21033) );
  INV_X1 U23994 ( .A(n21031), .ZN(n21024) );
  NOR2_X1 U23995 ( .A1(n21024), .A2(n21141), .ZN(n21026) );
  OAI21_X1 U23996 ( .B1(n21145), .B2(n21026), .A(n21025), .ZN(n21027) );
  AOI22_X1 U23997 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n21050), .B1(
        n21056), .B2(n21055), .ZN(n21032) );
  OAI211_X1 U23998 ( .C1(n21070), .C2(n21044), .A(n21033), .B(n21032), .ZN(
        P1_U3121) );
  AOI22_X1 U23999 ( .A1(n21155), .A2(n21048), .B1(n21154), .B2(n21047), .ZN(
        n21035) );
  AOI22_X1 U24000 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n21050), .B1(
        n21049), .B2(n21102), .ZN(n21034) );
  OAI211_X1 U24001 ( .C1(n21105), .C2(n21090), .A(n21035), .B(n21034), .ZN(
        P1_U3122) );
  AOI22_X1 U24002 ( .A1(n21161), .A2(n21048), .B1(n21160), .B2(n21047), .ZN(
        n21037) );
  AOI22_X1 U24003 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n21050), .B1(
        n21049), .B2(n21106), .ZN(n21036) );
  OAI211_X1 U24004 ( .C1(n21109), .C2(n21090), .A(n21037), .B(n21036), .ZN(
        P1_U3123) );
  AOI22_X1 U24005 ( .A1(n21167), .A2(n21048), .B1(n21166), .B2(n21047), .ZN(
        n21039) );
  AOI22_X1 U24006 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n21050), .B1(
        n21049), .B2(n21110), .ZN(n21038) );
  OAI211_X1 U24007 ( .C1(n21113), .C2(n21090), .A(n21039), .B(n21038), .ZN(
        P1_U3124) );
  AOI22_X1 U24008 ( .A1(n21173), .A2(n21048), .B1(n21172), .B2(n21047), .ZN(
        n21041) );
  AOI22_X1 U24009 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n21050), .B1(
        n21049), .B2(n21114), .ZN(n21040) );
  OAI211_X1 U24010 ( .C1(n21117), .C2(n21090), .A(n21041), .B(n21040), .ZN(
        P1_U3125) );
  AOI22_X1 U24011 ( .A1(n21179), .A2(n21048), .B1(n21178), .B2(n21047), .ZN(
        n21043) );
  AOI22_X1 U24012 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n21050), .B1(
        n21056), .B2(n21180), .ZN(n21042) );
  OAI211_X1 U24013 ( .C1(n21183), .C2(n21044), .A(n21043), .B(n21042), .ZN(
        P1_U3126) );
  AOI22_X1 U24014 ( .A1(n21185), .A2(n21048), .B1(n21184), .B2(n21047), .ZN(
        n21046) );
  AOI22_X1 U24015 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n21050), .B1(
        n21049), .B2(n21186), .ZN(n21045) );
  OAI211_X1 U24016 ( .C1(n21191), .C2(n21090), .A(n21046), .B(n21045), .ZN(
        P1_U3127) );
  AOI22_X1 U24017 ( .A1(n21195), .A2(n21048), .B1(n21193), .B2(n21047), .ZN(
        n21052) );
  AOI22_X1 U24018 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n21050), .B1(
        n21049), .B2(n21126), .ZN(n21051) );
  OAI211_X1 U24019 ( .C1(n21131), .C2(n21090), .A(n21052), .B(n21051), .ZN(
        P1_U3128) );
  AOI22_X1 U24020 ( .A1(n21138), .A2(n10548), .B1(n21085), .B2(n21055), .ZN(
        n21069) );
  NOR3_X1 U24021 ( .A1(n21056), .A2(n21085), .A3(n21141), .ZN(n21059) );
  INV_X1 U24022 ( .A(n21057), .ZN(n21058) );
  NOR2_X1 U24023 ( .A1(n21059), .A2(n21058), .ZN(n21067) );
  INV_X1 U24024 ( .A(n21067), .ZN(n21062) );
  NAND2_X1 U24025 ( .A1(n21134), .A2(n21060), .ZN(n21066) );
  INV_X1 U24026 ( .A(n21061), .ZN(n21065) );
  AOI22_X1 U24027 ( .A1(n21062), .A2(n21066), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21065), .ZN(n21063) );
  AOI22_X1 U24028 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n21087), .B1(
        n21139), .B2(n21086), .ZN(n21068) );
  OAI211_X1 U24029 ( .C1(n21070), .C2(n21090), .A(n21069), .B(n21068), .ZN(
        P1_U3129) );
  AOI22_X1 U24030 ( .A1(n21154), .A2(n10548), .B1(n21085), .B2(n21156), .ZN(
        n21072) );
  AOI22_X1 U24031 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n21087), .B1(
        n21155), .B2(n21086), .ZN(n21071) );
  OAI211_X1 U24032 ( .C1(n21159), .C2(n21090), .A(n21072), .B(n21071), .ZN(
        P1_U3130) );
  AOI22_X1 U24033 ( .A1(n21160), .A2(n10548), .B1(n21085), .B2(n21162), .ZN(
        n21074) );
  AOI22_X1 U24034 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n21087), .B1(
        n21161), .B2(n21086), .ZN(n21073) );
  OAI211_X1 U24035 ( .C1(n21165), .C2(n21090), .A(n21074), .B(n21073), .ZN(
        P1_U3131) );
  AOI22_X1 U24036 ( .A1(n21166), .A2(n10548), .B1(n21085), .B2(n21168), .ZN(
        n21076) );
  AOI22_X1 U24037 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n21087), .B1(
        n21167), .B2(n21086), .ZN(n21075) );
  OAI211_X1 U24038 ( .C1(n21171), .C2(n21090), .A(n21076), .B(n21075), .ZN(
        P1_U3132) );
  AOI22_X1 U24039 ( .A1(n21172), .A2(n10548), .B1(n21085), .B2(n21174), .ZN(
        n21078) );
  AOI22_X1 U24040 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n21087), .B1(
        n21173), .B2(n21086), .ZN(n21077) );
  OAI211_X1 U24041 ( .C1(n21177), .C2(n21090), .A(n21078), .B(n21077), .ZN(
        P1_U3133) );
  AOI22_X1 U24042 ( .A1(n21178), .A2(n10548), .B1(n21085), .B2(n21180), .ZN(
        n21080) );
  AOI22_X1 U24043 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n21087), .B1(
        n21179), .B2(n21086), .ZN(n21079) );
  OAI211_X1 U24044 ( .C1(n21183), .C2(n21090), .A(n21080), .B(n21079), .ZN(
        P1_U3134) );
  AOI22_X1 U24045 ( .A1(n21184), .A2(n10548), .B1(n21085), .B2(n21081), .ZN(
        n21083) );
  AOI22_X1 U24046 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n21087), .B1(
        n21185), .B2(n21086), .ZN(n21082) );
  OAI211_X1 U24047 ( .C1(n21084), .C2(n21090), .A(n21083), .B(n21082), .ZN(
        P1_U3135) );
  AOI22_X1 U24048 ( .A1(n21193), .A2(n10548), .B1(n21085), .B2(n21196), .ZN(
        n21089) );
  AOI22_X1 U24049 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n21087), .B1(
        n21195), .B2(n21086), .ZN(n21088) );
  OAI211_X1 U24050 ( .C1(n21202), .C2(n21090), .A(n21089), .B(n21088), .ZN(
        P1_U3136) );
  NAND2_X1 U24051 ( .A1(n21134), .A2(n21092), .ZN(n21095) );
  OAI22_X1 U24052 ( .A1(n21095), .A2(n21141), .B1(n21094), .B2(n21093), .ZN(
        n21125) );
  NOR3_X2 U24053 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21136), .A3(
        n21135), .ZN(n21124) );
  AOI22_X1 U24054 ( .A1(n21139), .A2(n21125), .B1(n21138), .B2(n21124), .ZN(
        n21101) );
  INV_X1 U24055 ( .A(n21201), .ZN(n21187) );
  OAI21_X1 U24056 ( .B1(n21187), .B2(n21127), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21096) );
  AOI21_X1 U24057 ( .B1(n21096), .B2(n21095), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n21099) );
  AOI22_X1 U24058 ( .A1(n21128), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n21127), .B2(n21150), .ZN(n21100) );
  OAI211_X1 U24059 ( .C1(n21153), .C2(n21201), .A(n21101), .B(n21100), .ZN(
        P1_U3145) );
  AOI22_X1 U24060 ( .A1(n21155), .A2(n21125), .B1(n21154), .B2(n21124), .ZN(
        n21104) );
  AOI22_X1 U24061 ( .A1(n21128), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n21127), .B2(n21102), .ZN(n21103) );
  OAI211_X1 U24062 ( .C1(n21105), .C2(n21201), .A(n21104), .B(n21103), .ZN(
        P1_U3146) );
  AOI22_X1 U24063 ( .A1(n21161), .A2(n21125), .B1(n21160), .B2(n21124), .ZN(
        n21108) );
  AOI22_X1 U24064 ( .A1(n21128), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n21127), .B2(n21106), .ZN(n21107) );
  OAI211_X1 U24065 ( .C1(n21109), .C2(n21201), .A(n21108), .B(n21107), .ZN(
        P1_U3147) );
  AOI22_X1 U24066 ( .A1(n21167), .A2(n21125), .B1(n21166), .B2(n21124), .ZN(
        n21112) );
  AOI22_X1 U24067 ( .A1(n21128), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n21127), .B2(n21110), .ZN(n21111) );
  OAI211_X1 U24068 ( .C1(n21113), .C2(n21201), .A(n21112), .B(n21111), .ZN(
        P1_U3148) );
  AOI22_X1 U24069 ( .A1(n21173), .A2(n21125), .B1(n21172), .B2(n21124), .ZN(
        n21116) );
  AOI22_X1 U24070 ( .A1(n21128), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n21127), .B2(n21114), .ZN(n21115) );
  OAI211_X1 U24071 ( .C1(n21117), .C2(n21201), .A(n21116), .B(n21115), .ZN(
        P1_U3149) );
  AOI22_X1 U24072 ( .A1(n21179), .A2(n21125), .B1(n21178), .B2(n21124), .ZN(
        n21120) );
  AOI22_X1 U24073 ( .A1(n21128), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n21127), .B2(n21118), .ZN(n21119) );
  OAI211_X1 U24074 ( .C1(n21121), .C2(n21201), .A(n21120), .B(n21119), .ZN(
        P1_U3150) );
  AOI22_X1 U24075 ( .A1(n21185), .A2(n21125), .B1(n21184), .B2(n21124), .ZN(
        n21123) );
  AOI22_X1 U24076 ( .A1(n21128), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n21127), .B2(n21186), .ZN(n21122) );
  OAI211_X1 U24077 ( .C1(n21191), .C2(n21201), .A(n21123), .B(n21122), .ZN(
        P1_U3151) );
  AOI22_X1 U24078 ( .A1(n21195), .A2(n21125), .B1(n21193), .B2(n21124), .ZN(
        n21130) );
  AOI22_X1 U24079 ( .A1(n21128), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n21127), .B2(n21126), .ZN(n21129) );
  OAI211_X1 U24080 ( .C1(n21131), .C2(n21201), .A(n21130), .B(n21129), .ZN(
        P1_U3152) );
  NOR2_X1 U24081 ( .A1(n21132), .A2(n21135), .ZN(n21192) );
  AOI21_X1 U24082 ( .B1(n21134), .B2(n21133), .A(n21192), .ZN(n21143) );
  NOR2_X1 U24083 ( .A1(n21136), .A2(n21135), .ZN(n21148) );
  INV_X1 U24084 ( .A(n21148), .ZN(n21137) );
  OAI22_X1 U24085 ( .A1(n21143), .A2(n21141), .B1(n21137), .B2(n11830), .ZN(
        n21194) );
  AOI22_X1 U24086 ( .A1(n21139), .A2(n21194), .B1(n21138), .B2(n21192), .ZN(
        n21152) );
  INV_X1 U24087 ( .A(n21140), .ZN(n21142) );
  NOR2_X1 U24088 ( .A1(n21142), .A2(n21141), .ZN(n21144) );
  OAI21_X1 U24089 ( .B1(n21145), .B2(n21144), .A(n21143), .ZN(n21146) );
  AOI22_X1 U24090 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21198), .B1(
        n21187), .B2(n21150), .ZN(n21151) );
  OAI211_X1 U24091 ( .C1(n21153), .C2(n21190), .A(n21152), .B(n21151), .ZN(
        P1_U3153) );
  AOI22_X1 U24092 ( .A1(n21155), .A2(n21194), .B1(n21154), .B2(n21192), .ZN(
        n21158) );
  AOI22_X1 U24093 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21198), .B1(
        n21197), .B2(n21156), .ZN(n21157) );
  OAI211_X1 U24094 ( .C1(n21159), .C2(n21201), .A(n21158), .B(n21157), .ZN(
        P1_U3154) );
  AOI22_X1 U24095 ( .A1(n21161), .A2(n21194), .B1(n21160), .B2(n21192), .ZN(
        n21164) );
  AOI22_X1 U24096 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21198), .B1(
        n21197), .B2(n21162), .ZN(n21163) );
  OAI211_X1 U24097 ( .C1(n21165), .C2(n21201), .A(n21164), .B(n21163), .ZN(
        P1_U3155) );
  AOI22_X1 U24098 ( .A1(n21167), .A2(n21194), .B1(n21166), .B2(n21192), .ZN(
        n21170) );
  AOI22_X1 U24099 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21198), .B1(
        n21197), .B2(n21168), .ZN(n21169) );
  OAI211_X1 U24100 ( .C1(n21171), .C2(n21201), .A(n21170), .B(n21169), .ZN(
        P1_U3156) );
  AOI22_X1 U24101 ( .A1(n21173), .A2(n21194), .B1(n21172), .B2(n21192), .ZN(
        n21176) );
  AOI22_X1 U24102 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21198), .B1(
        n21197), .B2(n21174), .ZN(n21175) );
  OAI211_X1 U24103 ( .C1(n21177), .C2(n21201), .A(n21176), .B(n21175), .ZN(
        P1_U3157) );
  AOI22_X1 U24104 ( .A1(n21179), .A2(n21194), .B1(n21178), .B2(n21192), .ZN(
        n21182) );
  AOI22_X1 U24105 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21198), .B1(
        n21197), .B2(n21180), .ZN(n21181) );
  OAI211_X1 U24106 ( .C1(n21183), .C2(n21201), .A(n21182), .B(n21181), .ZN(
        P1_U3158) );
  AOI22_X1 U24107 ( .A1(n21185), .A2(n21194), .B1(n21184), .B2(n21192), .ZN(
        n21189) );
  AOI22_X1 U24108 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21198), .B1(
        n21187), .B2(n21186), .ZN(n21188) );
  OAI211_X1 U24109 ( .C1(n21191), .C2(n21190), .A(n21189), .B(n21188), .ZN(
        P1_U3159) );
  AOI22_X1 U24110 ( .A1(n21195), .A2(n21194), .B1(n21193), .B2(n21192), .ZN(
        n21200) );
  AOI22_X1 U24111 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21198), .B1(
        n21197), .B2(n21196), .ZN(n21199) );
  OAI211_X1 U24112 ( .C1(n21202), .C2(n21201), .A(n21200), .B(n21199), .ZN(
        P1_U3160) );
  OAI211_X1 U24113 ( .C1(n21205), .C2(n11830), .A(n21204), .B(n21203), .ZN(
        P1_U3163) );
  AND2_X1 U24114 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21284), .ZN(
        P1_U3164) );
  AND2_X1 U24115 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21284), .ZN(
        P1_U3165) );
  AND2_X1 U24116 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21284), .ZN(
        P1_U3166) );
  AND2_X1 U24117 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21284), .ZN(
        P1_U3167) );
  AND2_X1 U24118 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21284), .ZN(
        P1_U3168) );
  AND2_X1 U24119 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21284), .ZN(
        P1_U3169) );
  AND2_X1 U24120 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21284), .ZN(
        P1_U3170) );
  AND2_X1 U24121 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21284), .ZN(
        P1_U3171) );
  AND2_X1 U24122 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21284), .ZN(
        P1_U3172) );
  AND2_X1 U24123 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21284), .ZN(
        P1_U3173) );
  AND2_X1 U24124 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21284), .ZN(
        P1_U3174) );
  AND2_X1 U24125 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21284), .ZN(
        P1_U3175) );
  AND2_X1 U24126 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21284), .ZN(
        P1_U3176) );
  AND2_X1 U24127 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21284), .ZN(
        P1_U3177) );
  AND2_X1 U24128 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21284), .ZN(
        P1_U3178) );
  AND2_X1 U24129 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21284), .ZN(
        P1_U3179) );
  AND2_X1 U24130 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21284), .ZN(
        P1_U3180) );
  AND2_X1 U24131 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21284), .ZN(
        P1_U3181) );
  AND2_X1 U24132 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21284), .ZN(
        P1_U3182) );
  AND2_X1 U24133 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21284), .ZN(
        P1_U3183) );
  AND2_X1 U24134 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21284), .ZN(
        P1_U3184) );
  AND2_X1 U24135 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21284), .ZN(
        P1_U3185) );
  AND2_X1 U24136 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21284), .ZN(P1_U3186) );
  AND2_X1 U24137 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21284), .ZN(P1_U3187) );
  AND2_X1 U24138 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21284), .ZN(P1_U3188) );
  AND2_X1 U24139 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21284), .ZN(P1_U3189) );
  AND2_X1 U24140 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21284), .ZN(P1_U3190) );
  AND2_X1 U24141 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21284), .ZN(P1_U3191) );
  AND2_X1 U24142 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21284), .ZN(P1_U3192) );
  AND2_X1 U24143 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21284), .ZN(P1_U3193) );
  AOI21_X1 U24144 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21212), .A(n21206), 
        .ZN(n21221) );
  OAI211_X1 U24145 ( .C1(P1_STATE_REG_0__SCAN_IN), .C2(n21213), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .B(n21207), .ZN(n21208) );
  NOR2_X1 U24146 ( .A1(n21209), .A2(n21208), .ZN(n21210) );
  OAI22_X1 U24147 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21221), .B1(n21309), 
        .B2(n21210), .ZN(P1_U3194) );
  OAI21_X1 U24148 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n21211), .A(n21213), 
        .ZN(n21219) );
  NAND3_X1 U24149 ( .A1(n21213), .A2(n21212), .A3(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n21215) );
  NAND2_X1 U24150 ( .A1(n21215), .A2(n21214), .ZN(n21216) );
  OAI211_X1 U24151 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21217), .A(HOLD), .B(
        n21216), .ZN(n21218) );
  OAI221_X1 U24152 ( .B1(n21221), .B2(n21220), .C1(n21221), .C2(n21219), .A(
        n21218), .ZN(P1_U3196) );
  NOR2_X1 U24153 ( .A1(n21303), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n21269) );
  NAND2_X1 U24154 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21309), .ZN(n21271) );
  INV_X1 U24155 ( .A(n21271), .ZN(n21273) );
  AOI222_X1 U24156 ( .A1(n21269), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n21303), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n21273), .ZN(n21222) );
  INV_X1 U24157 ( .A(n21222), .ZN(P1_U3197) );
  AOI222_X1 U24158 ( .A1(n21273), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n21303), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n21269), .ZN(n21223) );
  INV_X1 U24159 ( .A(n21223), .ZN(P1_U3198) );
  OAI222_X1 U24160 ( .A1(n21271), .A2(n21225), .B1(n21224), .B2(n21309), .C1(
        n21226), .C2(n21275), .ZN(P1_U3199) );
  INV_X1 U24161 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n21227) );
  OAI222_X1 U24162 ( .A1(n21275), .A2(n21229), .B1(n21227), .B2(n21309), .C1(
        n21226), .C2(n21271), .ZN(P1_U3200) );
  INV_X1 U24163 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n21228) );
  INV_X1 U24164 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21230) );
  OAI222_X1 U24165 ( .A1(n21271), .A2(n21229), .B1(n21228), .B2(n21309), .C1(
        n21230), .C2(n21275), .ZN(P1_U3201) );
  INV_X1 U24166 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n21231) );
  OAI222_X1 U24167 ( .A1(n21275), .A2(n21233), .B1(n21231), .B2(n21309), .C1(
        n21230), .C2(n21271), .ZN(P1_U3202) );
  INV_X1 U24168 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n21232) );
  OAI222_X1 U24169 ( .A1(n21271), .A2(n21233), .B1(n21232), .B2(n21309), .C1(
        n21234), .C2(n21275), .ZN(P1_U3203) );
  INV_X1 U24170 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n21235) );
  OAI222_X1 U24171 ( .A1(n21275), .A2(n21237), .B1(n21235), .B2(n21309), .C1(
        n21234), .C2(n21271), .ZN(P1_U3204) );
  INV_X1 U24172 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n21236) );
  OAI222_X1 U24173 ( .A1(n21271), .A2(n21237), .B1(n21236), .B2(n21309), .C1(
        n21238), .C2(n21275), .ZN(P1_U3205) );
  INV_X1 U24174 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n21239) );
  OAI222_X1 U24175 ( .A1(n21275), .A2(n15357), .B1(n21239), .B2(n21309), .C1(
        n21238), .C2(n21271), .ZN(P1_U3206) );
  AOI22_X1 U24176 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n21303), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n21269), .ZN(n21240) );
  OAI21_X1 U24177 ( .B1(n15357), .B2(n21271), .A(n21240), .ZN(P1_U3207) );
  INV_X1 U24178 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21243) );
  AOI22_X1 U24179 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n21303), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n21273), .ZN(n21241) );
  OAI21_X1 U24180 ( .B1(n21243), .B2(n21275), .A(n21241), .ZN(P1_U3208) );
  INV_X1 U24181 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n21242) );
  OAI222_X1 U24182 ( .A1(n21271), .A2(n21243), .B1(n21242), .B2(n21309), .C1(
        n21244), .C2(n21275), .ZN(P1_U3209) );
  INV_X1 U24183 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n21245) );
  OAI222_X1 U24184 ( .A1(n21275), .A2(n21247), .B1(n21245), .B2(n21309), .C1(
        n21244), .C2(n21271), .ZN(P1_U3210) );
  INV_X1 U24185 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n21246) );
  OAI222_X1 U24186 ( .A1(n21271), .A2(n21247), .B1(n21246), .B2(n21309), .C1(
        n21249), .C2(n21275), .ZN(P1_U3211) );
  AOI22_X1 U24187 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n21303), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n21269), .ZN(n21248) );
  OAI21_X1 U24188 ( .B1(n21249), .B2(n21271), .A(n21248), .ZN(P1_U3212) );
  AOI22_X1 U24189 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n21303), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n21273), .ZN(n21250) );
  OAI21_X1 U24190 ( .B1(n21251), .B2(n21275), .A(n21250), .ZN(P1_U3213) );
  AOI222_X1 U24191 ( .A1(n21273), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n21303), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n21269), .ZN(n21252) );
  INV_X1 U24192 ( .A(n21252), .ZN(P1_U3214) );
  AOI222_X1 U24193 ( .A1(n21273), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n21303), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n21269), .ZN(n21253) );
  INV_X1 U24194 ( .A(n21253), .ZN(P1_U3215) );
  INV_X1 U24195 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n21255) );
  OAI222_X1 U24196 ( .A1(n21275), .A2(n21257), .B1(n21255), .B2(n21309), .C1(
        n21254), .C2(n21271), .ZN(P1_U3216) );
  INV_X1 U24197 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n21256) );
  OAI222_X1 U24198 ( .A1(n21271), .A2(n21257), .B1(n21256), .B2(n21309), .C1(
        n21259), .C2(n21275), .ZN(P1_U3217) );
  INV_X1 U24199 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n21258) );
  OAI222_X1 U24200 ( .A1(n21271), .A2(n21259), .B1(n21258), .B2(n21309), .C1(
        n21260), .C2(n21275), .ZN(P1_U3218) );
  INV_X1 U24201 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n21261) );
  OAI222_X1 U24202 ( .A1(n21275), .A2(n21263), .B1(n21261), .B2(n21309), .C1(
        n21260), .C2(n21271), .ZN(P1_U3219) );
  AOI22_X1 U24203 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(n21303), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(n21269), .ZN(n21262) );
  OAI21_X1 U24204 ( .B1(n21263), .B2(n21271), .A(n21262), .ZN(P1_U3220) );
  INV_X1 U24205 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21384) );
  AOI22_X1 U24206 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(n21303), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(n21273), .ZN(n21264) );
  OAI21_X1 U24207 ( .B1(n21384), .B2(n21275), .A(n21264), .ZN(P1_U3221) );
  INV_X1 U24208 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n21265) );
  OAI222_X1 U24209 ( .A1(n21275), .A2(n21267), .B1(n21265), .B2(n21309), .C1(
        n21384), .C2(n21271), .ZN(P1_U3222) );
  AOI22_X1 U24210 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(n21303), .B1(
        P1_REIP_REG_28__SCAN_IN), .B2(n21269), .ZN(n21266) );
  OAI21_X1 U24211 ( .B1(n21267), .B2(n21271), .A(n21266), .ZN(P1_U3223) );
  AOI22_X1 U24212 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(n21303), .B1(
        P1_REIP_REG_28__SCAN_IN), .B2(n21273), .ZN(n21268) );
  OAI21_X1 U24213 ( .B1(n21272), .B2(n21275), .A(n21268), .ZN(P1_U3224) );
  AOI22_X1 U24214 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(n21303), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(n21269), .ZN(n21270) );
  OAI21_X1 U24215 ( .B1(n21272), .B2(n21271), .A(n21270), .ZN(P1_U3225) );
  AOI22_X1 U24216 ( .A1(P1_ADDRESS_REG_29__SCAN_IN), .A2(n21303), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(n21273), .ZN(n21274) );
  OAI21_X1 U24217 ( .B1(n21276), .B2(n21275), .A(n21274), .ZN(P1_U3226) );
  INV_X1 U24218 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n21277) );
  AOI22_X1 U24219 ( .A1(n21309), .A2(n21278), .B1(n21277), .B2(n21303), .ZN(
        P1_U3458) );
  INV_X1 U24220 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21297) );
  INV_X1 U24221 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n21279) );
  AOI22_X1 U24222 ( .A1(n21309), .A2(n21297), .B1(n21279), .B2(n21303), .ZN(
        P1_U3459) );
  INV_X1 U24223 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n21280) );
  AOI22_X1 U24224 ( .A1(n21309), .A2(n21281), .B1(n21280), .B2(n21303), .ZN(
        P1_U3460) );
  INV_X1 U24225 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21300) );
  INV_X1 U24226 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n21282) );
  AOI22_X1 U24227 ( .A1(n21309), .A2(n21300), .B1(n21282), .B2(n21303), .ZN(
        P1_U3461) );
  INV_X1 U24228 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21285) );
  INV_X1 U24229 ( .A(n21286), .ZN(n21283) );
  AOI21_X1 U24230 ( .B1(n21285), .B2(n21284), .A(n21283), .ZN(P1_U3464) );
  OAI21_X1 U24231 ( .B1(n21288), .B2(n21287), .A(n21286), .ZN(P1_U3465) );
  AOI22_X1 U24232 ( .A1(n21292), .A2(n21291), .B1(n21290), .B2(n21289), .ZN(
        n21293) );
  INV_X1 U24233 ( .A(n21293), .ZN(n21295) );
  MUX2_X1 U24234 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n21295), .S(
        n21294), .Z(P1_U3469) );
  AOI211_X1 U24235 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_REIP_REG_1__SCAN_IN), .B(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21296) );
  AOI21_X1 U24236 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n21296), .ZN(n21298) );
  AOI22_X1 U24237 ( .A1(n21302), .A2(n21298), .B1(n21297), .B2(n21299), .ZN(
        P1_U3481) );
  NOR2_X1 U24238 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n21301) );
  AOI22_X1 U24239 ( .A1(n21302), .A2(n21301), .B1(n21300), .B2(n21299), .ZN(
        P1_U3482) );
  AOI22_X1 U24240 ( .A1(n21309), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21304), 
        .B2(n21303), .ZN(P1_U3483) );
  INV_X1 U24241 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n21306) );
  INV_X1 U24242 ( .A(n21308), .ZN(n21305) );
  AOI22_X1 U24243 ( .A1(n21308), .A2(n21307), .B1(n21306), .B2(n21305), .ZN(
        P1_U3484) );
  MUX2_X1 U24244 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n21309), .Z(P1_U3486) );
  AOI222_X1 U24245 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n21311), .B1(n18300), 
        .B2(P3_UWORD_REG_1__SCAN_IN), .C1(n21310), .C2(
        P3_DATAO_REG_17__SCAN_IN), .ZN(n21469) );
  NAND4_X1 U24246 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_31__SCAN_IN), .A3(n21428), .A4(n21335), .ZN(n21316)
         );
  NAND4_X1 U24247 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n21352), .A3(n21354), .A4(n21355), .ZN(n21315) );
  NAND4_X1 U24248 ( .A1(P1_EBX_REG_27__SCAN_IN), .A2(P1_EBX_REG_4__SCAN_IN), 
        .A3(BUF1_REG_17__SCAN_IN), .A4(P3_EBX_REG_18__SCAN_IN), .ZN(n21314) );
  NAND4_X1 U24249 ( .A1(n21312), .A2(n21338), .A3(
        P1_INSTQUEUE_REG_5__0__SCAN_IN), .A4(P3_UWORD_REG_0__SCAN_IN), .ZN(
        n21313) );
  NOR4_X1 U24250 ( .A1(n21316), .A2(n21315), .A3(n21314), .A4(n21313), .ZN(
        n21467) );
  INV_X1 U24251 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n21364) );
  NAND4_X1 U24252 ( .A1(BUF1_REG_14__SCAN_IN), .A2(BUF1_REG_5__SCAN_IN), .A3(
        n21364), .A4(n21358), .ZN(n21331) );
  NOR4_X1 U24253 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(DATAI_27_), 
        .A3(P2_DATAO_REG_14__SCAN_IN), .A4(n21367), .ZN(n21319) );
  NOR4_X1 U24254 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n21372), .A4(n21373), .ZN(
        n21318) );
  NOR3_X1 U24255 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(
        P1_REIP_REG_26__SCAN_IN), .A3(n21382), .ZN(n21317) );
  NAND4_X1 U24256 ( .A1(READY22_REG_SCAN_IN), .A2(n21319), .A3(n21318), .A4(
        n21317), .ZN(n21330) );
  NOR4_X1 U24257 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n21413), .A3(
        n21388), .A4(n13753), .ZN(n21323) );
  INV_X1 U24258 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n21416) );
  INV_X1 U24259 ( .A(P2_UWORD_REG_11__SCAN_IN), .ZN(n21420) );
  NOR4_X1 U24260 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(
        P2_ADDRESS_REG_16__SCAN_IN), .A3(n21416), .A4(n21420), .ZN(n21322) );
  NOR4_X1 U24261 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n21404), .A3(
        n21418), .A4(n21419), .ZN(n21321) );
  NOR4_X1 U24262 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_12__7__SCAN_IN), .A3(P1_EBX_REG_23__SCAN_IN), .A4(
        BUF2_REG_16__SCAN_IN), .ZN(n21320) );
  NAND4_X1 U24263 ( .A1(n21323), .A2(n21322), .A3(n21321), .A4(n21320), .ZN(
        n21329) );
  NOR4_X1 U24264 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(BUF1_REG_10__SCAN_IN), 
        .A3(P1_DATAO_REG_16__SCAN_IN), .A4(n13497), .ZN(n21327) );
  NOR4_X1 U24265 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_28__SCAN_IN), 
        .A4(n21446), .ZN(n21326) );
  NOR4_X1 U24266 ( .A1(P1_EAX_REG_8__SCAN_IN), .A2(
        P2_BYTEENABLE_REG_2__SCAN_IN), .A3(n21452), .A4(n21451), .ZN(n21325)
         );
  NOR4_X1 U24267 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(
        P1_DATAO_REG_12__SCAN_IN), .A3(P3_DATAO_REG_28__SCAN_IN), .A4(n21432), 
        .ZN(n21324) );
  NAND4_X1 U24268 ( .A1(n21327), .A2(n21326), .A3(n21325), .A4(n21324), .ZN(
        n21328) );
  NOR4_X1 U24269 ( .A1(n21331), .A2(n21330), .A3(n21329), .A4(n21328), .ZN(
        n21466) );
  AOI22_X1 U24270 ( .A1(n21333), .A2(keyinput21), .B1(n20768), .B2(keyinput46), 
        .ZN(n21332) );
  OAI221_X1 U24271 ( .B1(n21333), .B2(keyinput21), .C1(n20768), .C2(keyinput46), .A(n21332), .ZN(n21346) );
  AOI22_X1 U24272 ( .A1(n21336), .A2(keyinput6), .B1(keyinput27), .B2(n21335), 
        .ZN(n21334) );
  OAI221_X1 U24273 ( .B1(n21336), .B2(keyinput6), .C1(n21335), .C2(keyinput27), 
        .A(n21334), .ZN(n21345) );
  AOI22_X1 U24274 ( .A1(n21339), .A2(keyinput14), .B1(n21338), .B2(keyinput15), 
        .ZN(n21337) );
  OAI221_X1 U24275 ( .B1(n21339), .B2(keyinput14), .C1(n21338), .C2(keyinput15), .A(n21337), .ZN(n21344) );
  XNOR2_X1 U24276 ( .A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B(keyinput29), .ZN(
        n21342) );
  XNOR2_X1 U24277 ( .A(n21340), .B(keyinput18), .ZN(n21341) );
  NAND2_X1 U24278 ( .A1(n21342), .A2(n21341), .ZN(n21343) );
  NOR4_X1 U24279 ( .A1(n21346), .A2(n21345), .A3(n21344), .A4(n21343), .ZN(
        n21396) );
  AOI22_X1 U24280 ( .A1(n21349), .A2(keyinput16), .B1(keyinput1), .B2(n21348), 
        .ZN(n21347) );
  OAI221_X1 U24281 ( .B1(n21349), .B2(keyinput16), .C1(n21348), .C2(keyinput1), 
        .A(n21347), .ZN(n21362) );
  AOI22_X1 U24282 ( .A1(n21352), .A2(keyinput56), .B1(keyinput51), .B2(n21351), 
        .ZN(n21350) );
  OAI221_X1 U24283 ( .B1(n21352), .B2(keyinput56), .C1(n21351), .C2(keyinput51), .A(n21350), .ZN(n21361) );
  AOI22_X1 U24284 ( .A1(n21355), .A2(keyinput19), .B1(n21354), .B2(keyinput55), 
        .ZN(n21353) );
  OAI221_X1 U24285 ( .B1(n21355), .B2(keyinput19), .C1(n21354), .C2(keyinput55), .A(n21353), .ZN(n21360) );
  AOI22_X1 U24286 ( .A1(n21358), .A2(keyinput62), .B1(n21357), .B2(keyinput50), 
        .ZN(n21356) );
  OAI221_X1 U24287 ( .B1(n21358), .B2(keyinput62), .C1(n21357), .C2(keyinput50), .A(n21356), .ZN(n21359) );
  NOR4_X1 U24288 ( .A1(n21362), .A2(n21361), .A3(n21360), .A4(n21359), .ZN(
        n21395) );
  AOI22_X1 U24289 ( .A1(n15071), .A2(keyinput39), .B1(n21364), .B2(keyinput53), 
        .ZN(n21363) );
  OAI221_X1 U24290 ( .B1(n15071), .B2(keyinput39), .C1(n21364), .C2(keyinput53), .A(n21363), .ZN(n21377) );
  INV_X1 U24291 ( .A(DATAI_27_), .ZN(n21366) );
  AOI22_X1 U24292 ( .A1(n21367), .A2(keyinput22), .B1(n21366), .B2(keyinput40), 
        .ZN(n21365) );
  OAI221_X1 U24293 ( .B1(n21367), .B2(keyinput22), .C1(n21366), .C2(keyinput40), .A(n21365), .ZN(n21376) );
  AOI22_X1 U24294 ( .A1(n21370), .A2(keyinput31), .B1(n21369), .B2(keyinput45), 
        .ZN(n21368) );
  OAI221_X1 U24295 ( .B1(n21370), .B2(keyinput31), .C1(n21369), .C2(keyinput45), .A(n21368), .ZN(n21375) );
  AOI22_X1 U24296 ( .A1(n21373), .A2(keyinput44), .B1(n21372), .B2(keyinput13), 
        .ZN(n21371) );
  OAI221_X1 U24297 ( .B1(n21373), .B2(keyinput44), .C1(n21372), .C2(keyinput13), .A(n21371), .ZN(n21374) );
  NOR4_X1 U24298 ( .A1(n21377), .A2(n21376), .A3(n21375), .A4(n21374), .ZN(
        n21394) );
  AOI22_X1 U24299 ( .A1(n21379), .A2(keyinput30), .B1(n12451), .B2(keyinput24), 
        .ZN(n21378) );
  OAI221_X1 U24300 ( .B1(n21379), .B2(keyinput30), .C1(n12451), .C2(keyinput24), .A(n21378), .ZN(n21392) );
  INV_X1 U24301 ( .A(READY22_REG_SCAN_IN), .ZN(n21381) );
  AOI22_X1 U24302 ( .A1(n21382), .A2(keyinput47), .B1(keyinput60), .B2(n21381), 
        .ZN(n21380) );
  OAI221_X1 U24303 ( .B1(n21382), .B2(keyinput47), .C1(n21381), .C2(keyinput60), .A(n21380), .ZN(n21391) );
  INV_X1 U24304 ( .A(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n21385) );
  AOI22_X1 U24305 ( .A1(n21385), .A2(keyinput2), .B1(keyinput12), .B2(n21384), 
        .ZN(n21383) );
  OAI221_X1 U24306 ( .B1(n21385), .B2(keyinput2), .C1(n21384), .C2(keyinput12), 
        .A(n21383), .ZN(n21390) );
  AOI22_X1 U24307 ( .A1(n21388), .A2(keyinput37), .B1(n21387), .B2(keyinput7), 
        .ZN(n21386) );
  OAI221_X1 U24308 ( .B1(n21388), .B2(keyinput37), .C1(n21387), .C2(keyinput7), 
        .A(n21386), .ZN(n21389) );
  NOR4_X1 U24309 ( .A1(n21392), .A2(n21391), .A3(n21390), .A4(n21389), .ZN(
        n21393) );
  NAND4_X1 U24310 ( .A1(n21396), .A2(n21395), .A3(n21394), .A4(n21393), .ZN(
        n21465) );
  AOI22_X1 U24311 ( .A1(n16263), .A2(keyinput20), .B1(n21398), .B2(keyinput8), 
        .ZN(n21397) );
  OAI221_X1 U24312 ( .B1(n16263), .B2(keyinput20), .C1(n21398), .C2(keyinput8), 
        .A(n21397), .ZN(n21399) );
  INV_X1 U24313 ( .A(n21399), .ZN(n21411) );
  AOI22_X1 U24314 ( .A1(n13497), .A2(keyinput28), .B1(n21401), .B2(keyinput33), 
        .ZN(n21400) );
  OAI221_X1 U24315 ( .B1(n13497), .B2(keyinput28), .C1(n21401), .C2(keyinput33), .A(n21400), .ZN(n21402) );
  INV_X1 U24316 ( .A(n21402), .ZN(n21410) );
  INV_X1 U24317 ( .A(keyinput49), .ZN(n21403) );
  XNOR2_X1 U24318 ( .A(n21404), .B(n21403), .ZN(n21409) );
  XNOR2_X1 U24319 ( .A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B(keyinput36), .ZN(
        n21407) );
  XNOR2_X1 U24320 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B(keyinput43), .ZN(
        n21406) );
  XNOR2_X1 U24321 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B(keyinput9), .ZN(
        n21405) );
  AND3_X1 U24322 ( .A1(n21407), .A2(n21406), .A3(n21405), .ZN(n21408) );
  AND4_X1 U24323 ( .A1(n21411), .A2(n21410), .A3(n21409), .A4(n21408), .ZN(
        n21463) );
  AOI22_X1 U24324 ( .A1(n13753), .A2(keyinput35), .B1(n21413), .B2(keyinput26), 
        .ZN(n21412) );
  OAI221_X1 U24325 ( .B1(n13753), .B2(keyinput35), .C1(n21413), .C2(keyinput26), .A(n21412), .ZN(n21426) );
  AOI22_X1 U24326 ( .A1(n21416), .A2(keyinput57), .B1(keyinput3), .B2(n21415), 
        .ZN(n21414) );
  OAI221_X1 U24327 ( .B1(n21416), .B2(keyinput57), .C1(n21415), .C2(keyinput3), 
        .A(n21414), .ZN(n21425) );
  AOI22_X1 U24328 ( .A1(n21419), .A2(keyinput17), .B1(n21418), .B2(keyinput54), 
        .ZN(n21417) );
  OAI221_X1 U24329 ( .B1(n21419), .B2(keyinput17), .C1(n21418), .C2(keyinput54), .A(n21417), .ZN(n21424) );
  XOR2_X1 U24330 ( .A(n21420), .B(keyinput23), .Z(n21422) );
  XNOR2_X1 U24331 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B(keyinput52), .ZN(
        n21421) );
  NAND2_X1 U24332 ( .A1(n21422), .A2(n21421), .ZN(n21423) );
  NOR4_X1 U24333 ( .A1(n21426), .A2(n21425), .A3(n21424), .A4(n21423), .ZN(
        n21462) );
  AOI22_X1 U24334 ( .A1(n21429), .A2(keyinput5), .B1(n21428), .B2(keyinput41), 
        .ZN(n21427) );
  OAI221_X1 U24335 ( .B1(n21429), .B2(keyinput5), .C1(n21428), .C2(keyinput41), 
        .A(n21427), .ZN(n21430) );
  INV_X1 U24336 ( .A(n21430), .ZN(n21444) );
  AOI22_X1 U24337 ( .A1(n21433), .A2(keyinput38), .B1(n21432), .B2(keyinput63), 
        .ZN(n21431) );
  OAI221_X1 U24338 ( .B1(n21433), .B2(keyinput38), .C1(n21432), .C2(keyinput63), .A(n21431), .ZN(n21436) );
  XNOR2_X1 U24339 ( .A(n21434), .B(keyinput10), .ZN(n21435) );
  NOR2_X1 U24340 ( .A1(n21436), .A2(n21435), .ZN(n21443) );
  AOI22_X1 U24341 ( .A1(n21439), .A2(keyinput11), .B1(n21438), .B2(keyinput61), 
        .ZN(n21437) );
  OAI221_X1 U24342 ( .B1(n21439), .B2(keyinput11), .C1(n21438), .C2(keyinput61), .A(n21437), .ZN(n21440) );
  INV_X1 U24343 ( .A(n21440), .ZN(n21442) );
  XNOR2_X1 U24344 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B(keyinput59), .ZN(
        n21441) );
  AND4_X1 U24345 ( .A1(n21444), .A2(n21443), .A3(n21442), .A4(n21441), .ZN(
        n21461) );
  AOI22_X1 U24346 ( .A1(n21446), .A2(keyinput0), .B1(n10819), .B2(keyinput34), 
        .ZN(n21445) );
  OAI221_X1 U24347 ( .B1(n21446), .B2(keyinput0), .C1(n10819), .C2(keyinput34), 
        .A(n21445), .ZN(n21459) );
  AOI22_X1 U24348 ( .A1(n21449), .A2(keyinput25), .B1(keyinput4), .B2(n21448), 
        .ZN(n21447) );
  OAI221_X1 U24349 ( .B1(n21449), .B2(keyinput25), .C1(n21448), .C2(keyinput4), 
        .A(n21447), .ZN(n21458) );
  AOI22_X1 U24350 ( .A1(n21452), .A2(keyinput58), .B1(keyinput42), .B2(n21451), 
        .ZN(n21450) );
  OAI221_X1 U24351 ( .B1(n21452), .B2(keyinput58), .C1(n21451), .C2(keyinput42), .A(n21450), .ZN(n21457) );
  AOI22_X1 U24352 ( .A1(n21455), .A2(keyinput32), .B1(n21454), .B2(keyinput48), 
        .ZN(n21453) );
  OAI221_X1 U24353 ( .B1(n21455), .B2(keyinput32), .C1(n21454), .C2(keyinput48), .A(n21453), .ZN(n21456) );
  NOR4_X1 U24354 ( .A1(n21459), .A2(n21458), .A3(n21457), .A4(n21456), .ZN(
        n21460) );
  NAND4_X1 U24355 ( .A1(n21463), .A2(n21462), .A3(n21461), .A4(n21460), .ZN(
        n21464) );
  AOI211_X1 U24356 ( .C1(n21467), .C2(n21466), .A(n21465), .B(n21464), .ZN(
        n21468) );
  XNOR2_X1 U24357 ( .A(n21469), .B(n21468), .ZN(P3_U2750) );
  AND2_X2 U13859 ( .A1(n10566), .A2(n14507), .ZN(n10622) );
  CLKBUF_X2 U11034 ( .A(n10782), .Z(n10787) );
  CLKBUF_X1 U11043 ( .A(n16329), .Z(n9582) );
  CLKBUF_X2 U11063 ( .A(n11278), .Z(n11093) );
  CLKBUF_X1 U11077 ( .A(n10834), .Z(n11275) );
  CLKBUF_X1 U11092 ( .A(n10833), .Z(n11271) );
  CLKBUF_X1 U11109 ( .A(n13997), .Z(n20824) );
  CLKBUF_X1 U11111 ( .A(n18721), .Z(n9585) );
  NAND2_X2 U11367 ( .A1(n18628), .A2(n18721), .ZN(n18716) );
  CLKBUF_X1 U12128 ( .A(n13606), .Z(n16831) );
  AND2_X2 U12245 ( .A1(n13563), .A2(n13777), .ZN(n21470) );
endmodule

