

module b22_C_AntiSAT_k_128_4 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287;

  OR2_X1 U7208 ( .A1(n13229), .A2(n12208), .ZN(n6816) );
  INV_X2 U7209 ( .A(n14871), .ZN(n14873) );
  XNOR2_X1 U7210 ( .A(n14132), .B(n13749), .ZN(n13980) );
  NAND2_X2 U7211 ( .A1(n9351), .A2(n9350), .ZN(n13288) );
  NAND2_X1 U7212 ( .A1(n13416), .A2(n13512), .ZN(n13404) );
  OAI22_X1 U7213 ( .A1(n11892), .A2(n7286), .B1(n7287), .B2(n11890), .ZN(
        n11896) );
  NAND2_X1 U7214 ( .A1(n9265), .A2(n9264), .ZN(n13562) );
  NAND2_X1 U7215 ( .A1(n7602), .A2(SI_24_), .ZN(n7604) );
  INV_X1 U7216 ( .A(n11727), .ZN(n6663) );
  CLKBUF_X2 U7217 ( .A(n10181), .Z(n6682) );
  OAI22_X1 U7218 ( .A1(n10978), .A2(n11964), .B1(n7106), .B2(n13764), .ZN(
        n10991) );
  OR2_X1 U7219 ( .A1(n7587), .A2(n7440), .ZN(n6893) );
  NOR2_X1 U7220 ( .A1(n10889), .A2(n10900), .ZN(n10826) );
  NAND2_X1 U7221 ( .A1(n14895), .A2(n14858), .ZN(n10889) );
  NAND2_X2 U7222 ( .A1(n7838), .A2(n7837), .ZN(n11837) );
  INV_X1 U7223 ( .A(n14525), .ZN(n12981) );
  INV_X4 U7224 ( .A(n9067), .ZN(n9449) );
  NAND2_X2 U7225 ( .A1(n9078), .A2(n9077), .ZN(n11413) );
  AND4_X1 U7226 ( .A1(n8349), .A2(n8348), .A3(n8347), .A4(n8346), .ZN(n12212)
         );
  INV_X2 U7227 ( .A(n11771), .ZN(n11946) );
  NAND2_X1 U7228 ( .A1(n6794), .A2(n7557), .ZN(n7804) );
  BUF_X1 U7229 ( .A(n8298), .Z(n8342) );
  BUF_X2 U7231 ( .A(n10442), .Z(n6475) );
  BUF_X2 U7232 ( .A(n7206), .Z(n9436) );
  BUF_X2 U7233 ( .A(n7707), .Z(n8072) );
  INV_X2 U7234 ( .A(n11929), .ZN(n11771) );
  AND3_X2 U7235 ( .A1(n7265), .A2(n7264), .A3(n7204), .ZN(n14895) );
  NAND4_X2 U7236 ( .A1(n8944), .A2(n8943), .A3(n8942), .A4(n8941), .ZN(n13181)
         );
  INV_X1 U7237 ( .A(n7707), .ZN(n11760) );
  CLKBUF_X2 U7238 ( .A(n8946), .Z(n8959) );
  NAND2_X1 U7239 ( .A1(n8904), .A2(n6854), .ZN(n13589) );
  INV_X2 U7240 ( .A(n8049), .ZN(n7673) );
  MUX2_X1 U7241 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8899), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n8900) );
  NAND2_X4 U7242 ( .A1(n7650), .A2(n7649), .ZN(n14132) );
  BUF_X2 U7243 ( .A(n7538), .Z(n7417) );
  NAND2_X1 U7244 ( .A1(n9684), .A2(P3_U3151), .ZN(n6460) );
  NAND2_X1 U7245 ( .A1(n9684), .A2(P3_U3151), .ZN(n6461) );
  INV_X4 U7246 ( .A(n7417), .ZN(n9684) );
  CLKBUF_X1 U7247 ( .A(n13683), .Z(n6462) );
  NOR2_X1 U7248 ( .A1(n11941), .A2(n9791), .ZN(n13683) );
  NAND2_X1 U7249 ( .A1(n8903), .A2(n8880), .ZN(n6463) );
  AND2_X1 U7250 ( .A1(n7201), .A2(n6464), .ZN(n10817) );
  NOR2_X1 U7251 ( .A1(n13087), .A2(n14934), .ZN(n6464) );
  INV_X1 U7252 ( .A(n11032), .ZN(n6465) );
  INV_X1 U7253 ( .A(n13316), .ZN(n6466) );
  NOR2_X1 U7254 ( .A1(n13340), .A2(n13331), .ZN(n6467) );
  AND2_X1 U7255 ( .A1(n14527), .A2(n14537), .ZN(n11461) );
  NOR2_X1 U7256 ( .A1(n13340), .A2(n13331), .ZN(n13330) );
  NAND2_X1 U7257 ( .A1(n13361), .A2(n13346), .ZN(n13340) );
  INV_X1 U7258 ( .A(n14954), .ZN(n14951) );
  NAND2_X1 U7259 ( .A1(n11758), .A2(n11763), .ZN(n11929) );
  NOR2_X1 U7260 ( .A1(n15094), .A2(n7391), .ZN(n7390) );
  XNOR2_X1 U7261 ( .A(n11091), .B(n15057), .ZN(n15053) );
  NAND2_X1 U7262 ( .A1(n12743), .A2(n12728), .ZN(n8553) );
  NOR2_X1 U7263 ( .A1(n10774), .A2(n8921), .ZN(n10179) );
  INV_X1 U7264 ( .A(n12068), .ZN(n9620) );
  NAND2_X1 U7265 ( .A1(n14084), .A2(n14074), .ZN(n14069) );
  INV_X1 U7267 ( .A(n8437), .ZN(n8546) );
  CLKBUF_X2 U7268 ( .A(n9251), .Z(n9426) );
  INV_X1 U7269 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13573) );
  INV_X1 U7270 ( .A(n12132), .ZN(n12121) );
  OAI21_X1 U7271 ( .B1(n9435), .B2(n9433), .A(n9419), .ZN(n9422) );
  AND4_X1 U7273 ( .A1(n8368), .A2(n8367), .A3(n8366), .A4(n8365), .ZN(n15163)
         );
  NAND2_X1 U7274 ( .A1(n13111), .A2(n12991), .ZN(n13053) );
  NAND2_X1 U7275 ( .A1(n13623), .A2(n12057), .ZN(n13689) );
  AND4_X1 U7276 ( .A1(n7730), .A2(n7729), .A3(n7728), .A4(n7727), .ZN(n11798)
         );
  INV_X1 U7277 ( .A(n14703), .ZN(n10532) );
  INV_X1 U7278 ( .A(n15163), .ZN(n12458) );
  NAND4_X1 U7279 ( .A1(n9029), .A2(n9028), .A3(n9027), .A4(n9026), .ZN(n13177)
         );
  INV_X1 U7280 ( .A(n14951), .ZN(n14535) );
  XNOR2_X1 U7281 ( .A(n8908), .B(n8907), .ZN(n9441) );
  XOR2_X1 U7282 ( .A(n14299), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n15274) );
  INV_X1 U7283 ( .A(n9406), .ZN(n9067) );
  INV_X1 U7284 ( .A(n11344), .ZN(n11396) );
  INV_X2 U7285 ( .A(n15181), .ZN(n15190) );
  OR2_X2 U7286 ( .A1(n14653), .A2(n14648), .ZN(n14654) );
  OAI21_X2 U7287 ( .B1(n10798), .B2(n6840), .A(n6839), .ZN(n10712) );
  AOI21_X2 U7288 ( .B1(n14432), .B2(n7048), .A(n6547), .ZN(n12410) );
  AOI21_X2 U7289 ( .B1(n14117), .B2(n14745), .A(n14116), .ZN(n6798) );
  NAND2_X2 U7290 ( .A1(n12671), .A2(n12247), .ZN(n12659) );
  NAND2_X2 U7291 ( .A1(n6666), .A2(n12246), .ZN(n12671) );
  NAND2_X2 U7292 ( .A1(n11450), .A2(n11449), .ZN(n14517) );
  OAI22_X2 U7293 ( .A1(n7456), .A2(n7005), .B1(n9141), .B2(n9140), .ZN(n9158)
         );
  OR2_X2 U7294 ( .A1(n14974), .A2(n15175), .ZN(n6621) );
  NAND2_X2 U7295 ( .A1(n14007), .A2(n8106), .ZN(n13992) );
  OAI21_X2 U7297 ( .B1(n12789), .B2(n7088), .A(n7086), .ZN(n12757) );
  NAND2_X2 U7298 ( .A1(n8467), .A2(n8759), .ZN(n12789) );
  NOR2_X4 U7299 ( .A1(n11604), .A2(n14571), .ZN(n14082) );
  NOR2_X2 U7300 ( .A1(n14328), .A2(n14329), .ZN(n14332) );
  NAND2_X2 U7302 ( .A1(n6793), .A2(n7420), .ZN(n7833) );
  NAND2_X2 U7303 ( .A1(n8660), .A2(n8659), .ZN(n12602) );
  AOI21_X2 U7304 ( .B1(n11649), .B2(n11648), .A(n11647), .ZN(n11650) );
  XNOR2_X1 U7305 ( .A(n9526), .B(n6736), .ZN(n10792) );
  XNOR2_X2 U7306 ( .A(n14987), .B(n11096), .ZN(n14976) );
  OAI21_X2 U7307 ( .B1(n11111), .B2(n15259), .A(n11095), .ZN(n11096) );
  XNOR2_X2 U7308 ( .A(n12462), .B(n11040), .ZN(n15181) );
  NAND3_X1 U7309 ( .A1(n6657), .A2(n8301), .A3(n8302), .ZN(n12462) );
  NAND4_X2 U7310 ( .A1(n8894), .A2(n8893), .A3(n8892), .A4(n8891), .ZN(n9472)
         );
  AND2_X2 U7311 ( .A1(n10817), .A2(n10708), .ZN(n10724) );
  NAND2_X2 U7312 ( .A1(n7825), .A2(n7824), .ZN(n14747) );
  XNOR2_X2 U7313 ( .A(n9422), .B(n9421), .ZN(n14236) );
  NAND4_X4 U7314 ( .A1(n8938), .A2(n8937), .A3(n8936), .A4(n8935), .ZN(n13182)
         );
  XNOR2_X2 U7315 ( .A(n13288), .B(n12166), .ZN(n13283) );
  OR2_X2 U7316 ( .A1(n15053), .A2(n15098), .ZN(n6752) );
  AND3_X2 U7317 ( .A1(n7719), .A2(n7718), .A3(n7717), .ZN(n14703) );
  NAND2_X2 U7318 ( .A1(n11784), .A2(n11783), .ZN(n11956) );
  NAND2_X1 U7319 ( .A1(n7128), .A2(n7127), .ZN(n10978) );
  AND3_X2 U7320 ( .A1(n7705), .A2(n7704), .A3(n7703), .ZN(n14682) );
  OAI222_X1 U7321 ( .A1(n14258), .A2(n14246), .B1(P1_U3086), .B2(n14245), .C1(
        n14262), .C2(n14244), .ZN(P1_U3327) );
  OR3_X2 U7322 ( .A1(n13968), .A2(n7120), .A3(n13980), .ZN(n7118) );
  XNOR2_X2 U7323 ( .A(n13972), .B(n12100), .ZN(n13968) );
  BUF_X1 U7324 ( .A(n8608), .Z(n6470) );
  BUF_X4 U7325 ( .A(n8608), .Z(n6471) );
  NAND2_X1 U7326 ( .A1(n8263), .A2(n12960), .ZN(n8608) );
  OAI21_X2 U7327 ( .B1(n15007), .B2(n15263), .A(n11098), .ZN(n11099) );
  XNOR2_X2 U7328 ( .A(n12299), .B(n12297), .ZN(n12400) );
  NAND2_X2 U7329 ( .A1(n12337), .A2(n12295), .ZN(n12299) );
  OAI21_X2 U7330 ( .B1(n8384), .B2(n8162), .A(n8163), .ZN(n8396) );
  OR2_X2 U7331 ( .A1(n15012), .A2(n11125), .ZN(n6751) );
  AND2_X1 U7332 ( .A1(n13242), .A2(n12182), .ZN(n13225) );
  INV_X2 U7333 ( .A(n12182), .ZN(n13438) );
  OAI21_X2 U7334 ( .B1(n6475), .B2(n15206), .A(n6623), .ZN(n10461) );
  XNOR2_X2 U7335 ( .A(n13470), .B(n13159), .ZN(n13301) );
  NAND2_X2 U7336 ( .A1(n7891), .A2(n7890), .ZN(n14558) );
  OAI21_X2 U7337 ( .B1(n15043), .B2(n15266), .A(n15040), .ZN(n11101) );
  NAND4_X4 U7338 ( .A1(n7685), .A2(n7684), .A3(n7683), .A4(n7682), .ZN(n13772)
         );
  OAI211_X2 U7339 ( .C1(n8602), .C2(n9688), .A(n8291), .B(n8290), .ZN(n10945)
         );
  NAND2_X1 U7340 ( .A1(n7193), .A2(n7194), .ZN(n6472) );
  NAND2_X4 U7341 ( .A1(n7193), .A2(n7194), .ZN(n10181) );
  INV_X2 U7342 ( .A(n7511), .ZN(n12000) );
  XNOR2_X1 U7343 ( .A(n11837), .B(n13762), .ZN(n11966) );
  XNOR2_X2 U7344 ( .A(n8120), .B(P1_IR_REG_24__SCAN_IN), .ZN(n14260) );
  OAI21_X2 U7345 ( .B1(n8141), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8120) );
  OAI21_X2 U7346 ( .B1(n8658), .B2(n8208), .A(n8209), .ZN(n8671) );
  INV_X2 U7347 ( .A(n8069), .ZN(n11938) );
  XNOR2_X2 U7348 ( .A(n8065), .B(P1_IR_REG_20__SCAN_IN), .ZN(n8069) );
  NAND2_X2 U7349 ( .A1(n9094), .A2(n9093), .ZN(n11445) );
  NAND2_X2 U7350 ( .A1(n14240), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7505) );
  NAND2_X2 U7351 ( .A1(n15188), .A2(n10945), .ZN(n9518) );
  BUF_X1 U7352 ( .A(n8293), .Z(n8678) );
  NOR2_X2 U7353 ( .A1(n14623), .A2(n14355), .ZN(n14415) );
  BUF_X1 U7354 ( .A(n10442), .Z(n6474) );
  XNOR2_X1 U7355 ( .A(n8308), .B(n8307), .ZN(n10442) );
  AND2_X4 U7356 ( .A1(n10944), .A2(n10730), .ZN(n9650) );
  INV_X1 U7357 ( .A(n9441), .ZN(n8921) );
  OAI21_X2 U7358 ( .B1(n14347), .B2(n6769), .A(n6766), .ZN(n14622) );
  OAI21_X2 U7359 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(n14342), .A(n14341), .ZN(
        n14347) );
  OR2_X1 U7360 ( .A1(n12809), .A2(n12852), .ZN(n12812) );
  NAND2_X1 U7361 ( .A1(n6810), .A2(n6816), .ZN(n13441) );
  NAND2_X1 U7362 ( .A1(n12632), .A2(n8799), .ZN(n12615) );
  XNOR2_X1 U7363 ( .A(n9416), .B(n9415), .ZN(n13580) );
  INV_X1 U7364 ( .A(n14120), .ZN(n13950) );
  OAI21_X1 U7365 ( .B1(n8553), .B2(n7083), .A(n7081), .ZN(n12698) );
  NAND2_X1 U7366 ( .A1(n14955), .A2(n15241), .ZN(n15076) );
  INV_X4 U7367 ( .A(n12296), .ZN(n12328) );
  INV_X1 U7368 ( .A(n13087), .ZN(n7200) );
  AND2_X1 U7370 ( .A1(n11791), .A2(n11792), .ZN(n11789) );
  CLKBUF_X2 U7371 ( .A(P2_U3947), .Z(n6477) );
  NAND4_X2 U7372 ( .A1(n7711), .A2(n7710), .A3(n7709), .A4(n7708), .ZN(n13771)
         );
  CLKBUF_X2 U7373 ( .A(n9057), .Z(n6478) );
  INV_X2 U7374 ( .A(n6470), .ZN(n8699) );
  INV_X4 U7375 ( .A(n8575), .ZN(n8288) );
  INV_X2 U7376 ( .A(n9406), .ZN(n8965) );
  INV_X1 U7377 ( .A(n8262), .ZN(n12960) );
  INV_X2 U7379 ( .A(n8034), .ZN(n11759) );
  NAND2_X1 U7380 ( .A1(n8259), .A2(n8237), .ZN(n12962) );
  INV_X2 U7381 ( .A(n12523), .ZN(n12550) );
  INV_X2 U7382 ( .A(n11364), .ZN(n9442) );
  CLKBUF_X2 U7383 ( .A(n9654), .Z(n12516) );
  INV_X1 U7384 ( .A(n14564), .ZN(n14058) );
  INV_X1 U7385 ( .A(n14264), .ZN(n11939) );
  NAND2_X1 U7386 ( .A1(n14264), .A2(n14564), .ZN(n11753) );
  NAND2_X1 U7387 ( .A1(n9684), .A2(P3_U3151), .ZN(n12964) );
  NAND4_X1 U7388 ( .A1(n7292), .A2(n7289), .A3(n7503), .A4(n7504), .ZN(n7615)
         );
  BUF_X1 U7389 ( .A(n10486), .Z(n6737) );
  OR2_X1 U7390 ( .A1(n6819), .A2(n14940), .ZN(n6812) );
  NAND2_X1 U7391 ( .A1(n6800), .A2(n6500), .ZN(n14115) );
  NAND2_X1 U7392 ( .A1(n8273), .A2(n8272), .ZN(n12558) );
  AND2_X1 U7393 ( .A1(n12582), .A2(n7409), .ZN(n12569) );
  AND2_X1 U7394 ( .A1(n13238), .A2(n13237), .ZN(n13443) );
  OR2_X1 U7395 ( .A1(n13441), .A2(n14938), .ZN(n6809) );
  NAND2_X1 U7396 ( .A1(n12254), .A2(n7410), .ZN(n12582) );
  AOI21_X1 U7397 ( .B1(n13438), .B2(n14933), .A(n13437), .ZN(n13439) );
  AND2_X1 U7398 ( .A1(n8812), .A2(n8813), .ZN(n12587) );
  NAND2_X1 U7399 ( .A1(n6687), .A2(n6686), .ZN(n13250) );
  NAND2_X1 U7400 ( .A1(n13447), .A2(n12206), .ZN(n13230) );
  NAND2_X1 U7401 ( .A1(n9424), .A2(n9423), .ZN(n9430) );
  NAND2_X1 U7402 ( .A1(n6808), .A2(n7249), .ZN(n13447) );
  NAND2_X1 U7403 ( .A1(n13284), .A2(n7250), .ZN(n6808) );
  AOI21_X1 U7404 ( .B1(n7250), .B2(n7251), .A(n6686), .ZN(n7249) );
  NAND2_X1 U7405 ( .A1(n8636), .A2(n8635), .ZN(n12909) );
  NAND2_X1 U7406 ( .A1(n12385), .A2(n12384), .ZN(n12383) );
  NOR2_X1 U7407 ( .A1(n13285), .A2(n13543), .ZN(n7203) );
  NAND2_X1 U7408 ( .A1(n7425), .A2(n8046), .ZN(n9416) );
  NOR2_X1 U7409 ( .A1(n14482), .A2(n14481), .ZN(n14483) );
  NAND2_X1 U7410 ( .A1(n8013), .A2(n8012), .ZN(n14006) );
  OAI21_X1 U7411 ( .B1(n8586), .B2(n7076), .A(n7074), .ZN(n8613) );
  NAND2_X2 U7412 ( .A1(n6685), .A2(n9333), .ZN(n13470) );
  NOR2_X1 U7413 ( .A1(n13996), .A2(n14212), .ZN(n6701) );
  XNOR2_X1 U7414 ( .A(n8027), .B(n8026), .ZN(n13594) );
  OR2_X1 U7415 ( .A1(n12529), .A2(n12530), .ZN(n6675) );
  XNOR2_X1 U7416 ( .A(n14365), .B(n14366), .ZN(n14374) );
  AOI21_X1 U7417 ( .B1(n9209), .B2(n9208), .A(n9207), .ZN(n9211) );
  NAND2_X1 U7418 ( .A1(n6993), .A2(n6992), .ZN(n9209) );
  NOR2_X1 U7419 ( .A1(n12496), .A2(n12495), .ZN(n12529) );
  AOI21_X1 U7420 ( .B1(n11519), .B2(n14359), .A(n14413), .ZN(n14365) );
  NAND2_X1 U7421 ( .A1(n12150), .A2(n12149), .ZN(n13399) );
  AND2_X1 U7422 ( .A1(n7661), .A2(n7600), .ZN(n7601) );
  NAND2_X1 U7423 ( .A1(n7365), .A2(n7364), .ZN(n11603) );
  NAND2_X1 U7424 ( .A1(n7921), .A2(n11862), .ZN(n11611) );
  OAI21_X1 U7425 ( .B1(n14517), .B2(n11451), .A(n11453), .ZN(n11535) );
  NAND2_X1 U7426 ( .A1(n8096), .A2(n8095), .ZN(n11315) );
  NAND2_X1 U7427 ( .A1(n8569), .A2(n8568), .ZN(n8571) );
  NAND2_X1 U7428 ( .A1(n7593), .A2(n7437), .ZN(n7997) );
  AOI21_X1 U7429 ( .B1(n11176), .B2(P2_REG1_REG_14__SCAN_IN), .A(n11175), .ZN(
        n11279) );
  NOR2_X1 U7430 ( .A1(n11573), .A2(n14558), .ZN(n6645) );
  NAND2_X1 U7431 ( .A1(n9167), .A2(n9166), .ZN(n11727) );
  AND2_X1 U7432 ( .A1(n7226), .A2(n7225), .ZN(n14606) );
  AND2_X2 U7433 ( .A1(n11461), .A2(n11712), .ZN(n11544) );
  OR2_X1 U7434 ( .A1(n14601), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7226) );
  NAND2_X1 U7435 ( .A1(n9216), .A2(n9215), .ZN(n13409) );
  NAND2_X1 U7436 ( .A1(n12231), .A2(n12230), .ZN(n12795) );
  AOI21_X1 U7437 ( .B1(n7115), .B2(n7113), .A(n6544), .ZN(n7112) );
  NAND2_X1 U7438 ( .A1(n8498), .A2(n8497), .ZN(n14424) );
  AOI21_X1 U7439 ( .B1(n11965), .B2(n7831), .A(n7116), .ZN(n7115) );
  NAND2_X1 U7440 ( .A1(n10961), .A2(n10960), .ZN(n11028) );
  NAND2_X1 U7441 ( .A1(n13081), .A2(n10750), .ZN(n10853) );
  OR2_X1 U7442 ( .A1(n10713), .A2(n6807), .ZN(n10961) );
  OAI21_X1 U7443 ( .B1(n15108), .B2(n7385), .A(n7383), .ZN(n15078) );
  NAND2_X1 U7444 ( .A1(n10746), .A2(n10745), .ZN(n13082) );
  NAND2_X1 U7445 ( .A1(n8087), .A2(n8086), .ZN(n10592) );
  NAND2_X1 U7446 ( .A1(n10691), .A2(n10690), .ZN(n10803) );
  NAND2_X1 U7447 ( .A1(n7188), .A2(n7187), .ZN(n10746) );
  AND2_X1 U7448 ( .A1(n7214), .A2(n7213), .ZN(n15037) );
  NAND2_X1 U7449 ( .A1(n15155), .A2(n7395), .ZN(n15159) );
  INV_X2 U7450 ( .A(n15204), .ZN(n15177) );
  OR2_X1 U7451 ( .A1(n8178), .A2(n10019), .ZN(n8179) );
  AND2_X1 U7452 ( .A1(n11045), .A2(n11044), .ZN(n11047) );
  NAND2_X1 U7453 ( .A1(n7201), .A2(n7200), .ZN(n10818) );
  NOR2_X1 U7454 ( .A1(n11338), .A2(n11337), .ZN(n14954) );
  NAND2_X1 U7455 ( .A1(n7554), .A2(n7553), .ZN(n7790) );
  NAND2_X1 U7456 ( .A1(n7230), .A2(n14321), .ZN(n14322) );
  AND2_X1 U7457 ( .A1(n8740), .A2(n8741), .ZN(n15138) );
  NAND2_X1 U7458 ( .A1(n7550), .A2(n7549), .ZN(n7775) );
  XNOR2_X1 U7459 ( .A(n11089), .B(n14987), .ZN(n14974) );
  INV_X2 U7460 ( .A(n14389), .ZN(n6476) );
  INV_X1 U7461 ( .A(n15111), .ZN(n15143) );
  INV_X1 U7462 ( .A(n10945), .ZN(n10738) );
  NAND2_X1 U7463 ( .A1(n7546), .A2(n7545), .ZN(n7761) );
  AND4_X1 U7464 ( .A1(n8382), .A2(n8381), .A3(n8380), .A4(n8379), .ZN(n15111)
         );
  AND4_X2 U7465 ( .A1(n8317), .A2(n8316), .A3(n8315), .A4(n8314), .ZN(n15186)
         );
  NOR2_X1 U7466 ( .A1(n11087), .A2(n6498), .ZN(n11089) );
  AND2_X1 U7467 ( .A1(n9514), .A2(n9513), .ZN(n12948) );
  AND2_X1 U7468 ( .A1(n7216), .A2(n7215), .ZN(n11087) );
  NAND4_X1 U7469 ( .A1(n7724), .A2(n7723), .A3(n7722), .A4(n7721), .ZN(n13770)
         );
  AND3_X1 U7470 ( .A1(n7674), .A2(n7675), .A3(n7141), .ZN(n7680) );
  NAND2_X2 U7471 ( .A1(n9640), .A2(n9753), .ZN(n14667) );
  AND3_X1 U7472 ( .A1(n8963), .A2(n8962), .A3(n6859), .ZN(n10827) );
  XNOR2_X1 U7473 ( .A(n8718), .B(P3_IR_REG_22__SCAN_IN), .ZN(n10730) );
  NAND2_X1 U7474 ( .A1(n8713), .A2(n8848), .ZN(n10614) );
  AND2_X1 U7475 ( .A1(n9634), .A2(n11766), .ZN(n11344) );
  OR2_X1 U7476 ( .A1(n7992), .A2(n7706), .ZN(n7709) );
  NAND2_X1 U7477 ( .A1(n12958), .A2(n12960), .ZN(n8293) );
  AND2_X1 U7478 ( .A1(n12958), .A2(n8262), .ZN(n8298) );
  XNOR2_X1 U7479 ( .A(n8884), .B(n8883), .ZN(n8889) );
  INV_X1 U7480 ( .A(n13581), .ZN(n8890) );
  NAND2_X2 U7481 ( .A1(n11753), .A2(n10518), .ZN(n12132) );
  NAND2_X1 U7482 ( .A1(n9441), .A2(n11364), .ZN(n14859) );
  NAND2_X1 U7483 ( .A1(n8888), .A2(n8887), .ZN(n13581) );
  NAND2_X1 U7484 ( .A1(n8887), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8884) );
  NAND2_X1 U7485 ( .A1(n12000), .A2(n7512), .ZN(n7707) );
  INV_X1 U7486 ( .A(n8922), .ZN(n13213) );
  OR2_X1 U7487 ( .A1(n6748), .A2(n6724), .ZN(n8258) );
  NAND2_X2 U7488 ( .A1(n7511), .A2(n14242), .ZN(n8034) );
  CLKBUF_X1 U7489 ( .A(n11364), .Z(n6618) );
  MUX2_X1 U7490 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8886), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n8888) );
  MUX2_X1 U7491 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8236), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n8237) );
  NAND2_X1 U7492 ( .A1(n8918), .A2(n9464), .ZN(n11364) );
  NAND2_X1 U7493 ( .A1(n14260), .A2(n8140), .ZN(n9634) );
  XNOR2_X1 U7494 ( .A(n8914), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8922) );
  MUX2_X1 U7495 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8902), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n8904) );
  OR2_X1 U7496 ( .A1(n8909), .A2(n13573), .ZN(n8911) );
  MUX2_X1 U7497 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8916), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n8918) );
  OR2_X1 U7498 ( .A1(n8917), .A2(n13573), .ZN(n8908) );
  AND2_X1 U7499 ( .A1(n8063), .A2(n8141), .ZN(n14264) );
  NAND2_X1 U7500 ( .A1(n8234), .A2(n8233), .ZN(n8259) );
  OAI21_X1 U7501 ( .B1(n9685), .B2(n9700), .A(n6733), .ZN(n7548) );
  NOR2_X1 U7502 ( .A1(n9232), .A2(n7196), .ZN(n8917) );
  XNOR2_X1 U7503 ( .A(n7509), .B(n7508), .ZN(n14242) );
  OR3_X1 U7504 ( .A1(n9232), .A2(n7195), .A3(P2_IR_REG_18__SCAN_IN), .ZN(n8915) );
  NAND2_X1 U7505 ( .A1(n7615), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7612) );
  AND2_X2 U7506 ( .A1(n8412), .A2(n8225), .ZN(n8227) );
  NOR2_X2 U7507 ( .A1(n7938), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n7953) );
  NOR2_X1 U7508 ( .A1(n8337), .A2(n7404), .ZN(n8354) );
  NAND2_X1 U7509 ( .A1(n8306), .A2(n8217), .ZN(n8337) );
  OR2_X1 U7510 ( .A1(n8306), .A2(n8238), .ZN(n8308) );
  NAND2_X1 U7511 ( .A1(n8895), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8286) );
  XNOR2_X1 U7512 ( .A(n6762), .B(P1_ADDR_REG_1__SCAN_IN), .ZN(n14302) );
  NOR2_X1 U7513 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n7492) );
  INV_X1 U7514 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8883) );
  INV_X1 U7515 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13218) );
  NOR2_X2 U7516 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8306) );
  INV_X1 U7517 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8895) );
  INV_X1 U7518 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8218) );
  INV_X1 U7519 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n6762) );
  AOI21_X2 U7520 ( .B1(n12261), .B2(n15183), .A(n12260), .ZN(n12813) );
  NOR2_X2 U7521 ( .A1(n10112), .A2(n10532), .ZN(n10529) );
  INV_X1 U7522 ( .A(n8923), .ZN(n10695) );
  NAND2_X1 U7523 ( .A1(n10217), .A2(n13589), .ZN(n6479) );
  NAND2_X1 U7524 ( .A1(n10217), .A2(n13589), .ZN(n6480) );
  NAND2_X1 U7525 ( .A1(n12812), .A2(n12813), .ZN(n12891) );
  NOR2_X4 U7526 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8932) );
  NOR2_X2 U7527 ( .A1(n14069), .A2(n13621), .ZN(n7108) );
  XNOR2_X2 U7528 ( .A(n13000), .B(n13001), .ZN(n13018) );
  OAI22_X2 U7529 ( .A1(n13123), .A2(n13122), .B1(n12999), .B2(n12998), .ZN(
        n13000) );
  NOR2_X2 U7530 ( .A1(n13895), .A2(n13894), .ZN(n13893) );
  NOR2_X4 U7531 ( .A1(n13417), .A2(n13520), .ZN(n13416) );
  OR2_X2 U7532 ( .A1(n11663), .A2(n13525), .ZN(n13417) );
  NOR2_X2 U7533 ( .A1(n8961), .A2(n8960), .ZN(n9863) );
  AOI22_X2 U7534 ( .A1(n11059), .A2(n11058), .B1(n11057), .B2(n11056), .ZN(
        n11064) );
  OAI22_X2 U7535 ( .A1(n10853), .A2(n10852), .B1(n10851), .B2(n10850), .ZN(
        n11059) );
  NOR2_X4 U7536 ( .A1(n13404), .A2(n13507), .ZN(n7208) );
  AND2_X2 U7537 ( .A1(n14082), .A2(n14233), .ZN(n14084) );
  NAND2_X1 U7538 ( .A1(n9755), .A2(n9684), .ZN(n7478) );
  INV_X1 U7539 ( .A(n6612), .ZN(n6611) );
  OAI21_X1 U7540 ( .B1(n12558), .B2(n12560), .A(n8705), .ZN(n8819) );
  NAND2_X1 U7541 ( .A1(n12816), .A2(n12570), .ZN(n8822) );
  NAND2_X1 U7542 ( .A1(n6731), .A2(n7610), .ZN(n8044) );
  OAI21_X1 U7543 ( .B1(n8027), .B2(n7444), .A(n7445), .ZN(n7608) );
  INV_X1 U7544 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7291) );
  AOI21_X1 U7545 ( .B1(n7561), .B2(n7421), .A(n6558), .ZN(n7420) );
  NAND2_X1 U7546 ( .A1(n8227), .A2(n7407), .ZN(n8572) );
  AND2_X1 U7547 ( .A1(n12203), .A2(n12202), .ZN(n13284) );
  NAND2_X1 U7548 ( .A1(n7258), .A2(n7257), .ZN(n12203) );
  NOR2_X1 U7549 ( .A1(n7260), .A2(n13301), .ZN(n7257) );
  NOR2_X1 U7550 ( .A1(n7371), .A2(n13932), .ZN(n7369) );
  INV_X1 U7551 ( .A(n9052), .ZN(n6971) );
  OAI21_X1 U7552 ( .B1(n6487), .B2(n6561), .A(n8727), .ZN(n8728) );
  NAND2_X1 U7553 ( .A1(n6736), .A2(n11040), .ZN(n6735) );
  NAND2_X1 U7554 ( .A1(n6945), .A2(n11834), .ZN(n6944) );
  OAI21_X1 U7555 ( .B1(n6505), .B2(n6607), .A(n8759), .ZN(n8764) );
  NAND2_X1 U7556 ( .A1(n8761), .A2(n6608), .ZN(n6607) );
  NAND2_X1 U7557 ( .A1(n14956), .A2(n14497), .ZN(n6608) );
  INV_X1 U7558 ( .A(n9332), .ZN(n7004) );
  INV_X1 U7559 ( .A(n9315), .ZN(n7470) );
  INV_X1 U7560 ( .A(n11909), .ZN(n7285) );
  AND2_X1 U7561 ( .A1(n7285), .A2(n11911), .ZN(n7284) );
  OR2_X1 U7562 ( .A1(n11911), .A2(n7285), .ZN(n7283) );
  OR2_X1 U7563 ( .A1(n11907), .A2(n11908), .ZN(n6697) );
  OR2_X1 U7564 ( .A1(n9430), .A2(n13220), .ZN(n9459) );
  INV_X1 U7565 ( .A(n12155), .ZN(n7269) );
  NAND2_X1 U7566 ( .A1(n11924), .A2(n11923), .ZN(n6905) );
  NOR2_X1 U7567 ( .A1(n7441), .A2(SI_18_), .ZN(n7440) );
  AND2_X1 U7568 ( .A1(n7574), .A2(n7477), .ZN(n7429) );
  AND2_X1 U7569 ( .A1(n12327), .A2(n6514), .ZN(n7060) );
  INV_X1 U7570 ( .A(n8844), .ZN(n8843) );
  NOR2_X1 U7571 ( .A1(n12587), .A2(n7411), .ZN(n7410) );
  INV_X1 U7572 ( .A(n12253), .ZN(n7411) );
  OR2_X1 U7573 ( .A1(n12677), .A2(n12685), .ZN(n8791) );
  NOR2_X1 U7574 ( .A1(n12773), .A2(n8767), .ZN(n7092) );
  NOR2_X1 U7575 ( .A1(n12689), .A2(n7078), .ZN(n7077) );
  INV_X1 U7576 ( .A(n8824), .ZN(n7078) );
  NAND2_X1 U7577 ( .A1(n8585), .A2(n8823), .ZN(n8586) );
  INV_X1 U7578 ( .A(n12698), .ZN(n8585) );
  INV_X1 U7579 ( .A(n8183), .ZN(n7024) );
  INV_X1 U7580 ( .A(n7017), .ZN(n7016) );
  OAI21_X1 U7581 ( .B1(n8428), .B2(n7018), .A(n8444), .ZN(n7017) );
  INV_X1 U7582 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8220) );
  INV_X1 U7583 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8219) );
  OR2_X1 U7584 ( .A1(n7161), .A2(n6593), .ZN(n7159) );
  NOR2_X1 U7585 ( .A1(n12152), .A2(n6875), .ZN(n6874) );
  INV_X1 U7586 ( .A(n12151), .ZN(n6875) );
  NAND2_X1 U7587 ( .A1(n12186), .A2(n6536), .ZN(n6832) );
  INV_X1 U7588 ( .A(n13422), .ZN(n6833) );
  INV_X1 U7589 ( .A(n6823), .ZN(n6821) );
  INV_X1 U7590 ( .A(n10669), .ZN(n6829) );
  XNOR2_X1 U7591 ( .A(n13180), .B(n10827), .ZN(n10685) );
  NAND2_X1 U7592 ( .A1(n6849), .A2(n13250), .ZN(n13235) );
  AND2_X1 U7593 ( .A1(n12171), .A2(n13231), .ZN(n6849) );
  INV_X1 U7594 ( .A(n8878), .ZN(n6856) );
  INV_X1 U7595 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8863) );
  NAND2_X1 U7596 ( .A1(n6912), .A2(n6698), .ZN(n6911) );
  INV_X1 U7597 ( .A(n10837), .ZN(n6698) );
  INV_X1 U7598 ( .A(n7317), .ZN(n6912) );
  AOI21_X1 U7599 ( .B1(n7316), .B2(n7319), .A(n11267), .ZN(n7315) );
  AND2_X1 U7600 ( .A1(n7318), .A2(n7321), .ZN(n7316) );
  AOI21_X1 U7601 ( .B1(n11921), .B2(n11920), .A(n11919), .ZN(n11925) );
  OR2_X1 U7602 ( .A1(n14558), .A2(n12016), .ZN(n11858) );
  INV_X1 U7603 ( .A(n11756), .ZN(n8113) );
  NAND2_X1 U7604 ( .A1(n7604), .A2(n6729), .ZN(n7453) );
  OAI21_X1 U7605 ( .B1(n7601), .B2(n6895), .A(n6598), .ZN(n6730) );
  NAND2_X1 U7606 ( .A1(n7431), .A2(SI_22_), .ZN(n7597) );
  OAI21_X1 U7607 ( .B1(n7587), .B2(n6887), .A(n6889), .ZN(n7591) );
  NAND2_X1 U7608 ( .A1(n6888), .A2(n7590), .ZN(n6887) );
  INV_X1 U7609 ( .A(n6890), .ZN(n6889) );
  INV_X1 U7610 ( .A(n7440), .ZN(n6888) );
  INV_X1 U7611 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U7612 ( .A1(n7581), .A2(n7580), .ZN(n7904) );
  NAND2_X1 U7613 ( .A1(n7695), .A2(n7531), .ZN(n7534) );
  AND2_X1 U7614 ( .A1(n7694), .A2(n7530), .ZN(n7531) );
  XNOR2_X1 U7615 ( .A(n14273), .B(n7237), .ZN(n14298) );
  NAND2_X1 U7616 ( .A1(n12307), .A2(n12584), .ZN(n7064) );
  OR2_X1 U7617 ( .A1(n12428), .A2(n7065), .ZN(n7062) );
  INV_X1 U7618 ( .A(n12391), .ZN(n7041) );
  OAI21_X1 U7619 ( .B1(n7063), .B2(n7060), .A(n6483), .ZN(n7055) );
  NOR2_X1 U7620 ( .A1(n12340), .A2(n7030), .ZN(n7029) );
  INV_X1 U7621 ( .A(n12293), .ZN(n7030) );
  NAND2_X1 U7622 ( .A1(n12267), .A2(n12266), .ZN(n12271) );
  NAND2_X1 U7623 ( .A1(n6506), .A2(n6624), .ZN(n6634) );
  NOR2_X1 U7624 ( .A1(n6679), .A2(n8842), .ZN(n6678) );
  INV_X1 U7625 ( .A(n10436), .ZN(n7215) );
  INV_X1 U7626 ( .A(n15038), .ZN(n7213) );
  NAND2_X1 U7627 ( .A1(n7224), .A2(n7223), .ZN(n7222) );
  INV_X1 U7628 ( .A(n11093), .ZN(n7223) );
  NOR2_X1 U7629 ( .A1(n11587), .A2(n8455), .ZN(n6754) );
  NAND2_X1 U7630 ( .A1(n6757), .A2(n6756), .ZN(n6673) );
  NAND2_X1 U7631 ( .A1(n12494), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n6756) );
  INV_X1 U7632 ( .A(n7217), .ZN(n12532) );
  AND2_X1 U7633 ( .A1(n8656), .A2(n8655), .ZN(n12597) );
  AOI21_X1 U7634 ( .B1(n7399), .B2(n7398), .A(n6512), .ZN(n7397) );
  INV_X1 U7635 ( .A(n12248), .ZN(n7398) );
  NAND2_X1 U7636 ( .A1(n12659), .A2(n12248), .ZN(n7402) );
  NAND2_X1 U7637 ( .A1(n12245), .A2(n12244), .ZN(n12673) );
  NAND2_X1 U7638 ( .A1(n12710), .A2(n7412), .ZN(n12699) );
  AND2_X1 U7639 ( .A1(n12700), .A2(n12242), .ZN(n7412) );
  AND2_X1 U7640 ( .A1(n8780), .A2(n8782), .ZN(n12713) );
  NAND2_X1 U7641 ( .A1(n7392), .A2(n7390), .ZN(n15091) );
  OAI21_X1 U7642 ( .B1(n14955), .B2(n15241), .A(n15076), .ZN(n15094) );
  INV_X1 U7643 ( .A(n15142), .ZN(n15185) );
  INV_X1 U7644 ( .A(n10614), .ZN(n10944) );
  CLKBUF_X1 U7645 ( .A(n8336), .Z(n8684) );
  AND3_X1 U7646 ( .A1(n12946), .A2(n12948), .A3(n10632), .ZN(n10608) );
  NOR2_X2 U7647 ( .A1(n6734), .A2(n7413), .ZN(n8234) );
  NAND2_X1 U7648 ( .A1(n7414), .A2(n8240), .ZN(n7413) );
  INV_X1 U7649 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8240) );
  XNOR2_X1 U7650 ( .A(n8852), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9512) );
  NAND2_X1 U7651 ( .A1(n6497), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8852) );
  NAND3_X1 U7652 ( .A1(n7008), .A2(n11240), .A3(n7007), .ZN(n8589) );
  NAND2_X1 U7653 ( .A1(n7180), .A2(n7177), .ZN(n7176) );
  NAND2_X1 U7654 ( .A1(n7182), .A2(n7179), .ZN(n7177) );
  NAND2_X1 U7655 ( .A1(n7156), .A2(n7152), .ZN(n7151) );
  INV_X1 U7656 ( .A(n13091), .ZN(n7152) );
  NAND2_X1 U7657 ( .A1(n7189), .A2(n7190), .ZN(n7188) );
  NOR2_X1 U7658 ( .A1(n7191), .A2(n10409), .ZN(n7190) );
  NOR2_X1 U7659 ( .A1(n6538), .A2(n6990), .ZN(n6989) );
  INV_X1 U7660 ( .A(n9487), .ZN(n6990) );
  AOI21_X1 U7661 ( .B1(n13580), .B2(n9436), .A(n7484), .ZN(n12182) );
  AND2_X1 U7662 ( .A1(n13254), .A2(n13540), .ZN(n13242) );
  NAND2_X1 U7663 ( .A1(n13235), .A2(n6848), .ZN(n6847) );
  NAND2_X1 U7664 ( .A1(n13540), .A2(n13155), .ZN(n6848) );
  NOR2_X2 U7665 ( .A1(n13270), .A2(n13448), .ZN(n13254) );
  NAND2_X1 U7666 ( .A1(n6834), .A2(n6489), .ZN(n7258) );
  NAND2_X1 U7667 ( .A1(n12192), .A2(n12191), .ZN(n13358) );
  NAND2_X1 U7668 ( .A1(n13372), .A2(n7270), .ZN(n13354) );
  OR2_X1 U7669 ( .A1(n11253), .A2(n6825), .ZN(n6822) );
  NAND2_X1 U7670 ( .A1(n11021), .A2(n11020), .ZN(n11022) );
  NAND2_X1 U7671 ( .A1(n10712), .A2(n10711), .ZN(n10713) );
  INV_X1 U7672 ( .A(n6838), .ZN(n6839) );
  INV_X1 U7673 ( .A(n6842), .ZN(n6840) );
  OAI21_X1 U7674 ( .B1(n6843), .B2(n6503), .A(n10674), .ZN(n6838) );
  NAND2_X1 U7675 ( .A1(n10697), .A2(n10696), .ZN(n14860) );
  INV_X2 U7677 ( .A(n9832), .ZN(n9244) );
  INV_X1 U7678 ( .A(n7433), .ZN(n7432) );
  OAI21_X1 U7679 ( .B1(n7596), .B2(n7435), .A(n9298), .ZN(n7433) );
  NAND2_X1 U7680 ( .A1(n8913), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8914) );
  NAND2_X1 U7681 ( .A1(n11265), .A2(n7324), .ZN(n7323) );
  INV_X1 U7682 ( .A(n11266), .ZN(n7324) );
  INV_X1 U7683 ( .A(n11351), .ZN(n6917) );
  OAI22_X1 U7684 ( .A1(n9620), .A2(n10136), .B1(n14682), .B2(n11717), .ZN(
        n9623) );
  NAND3_X1 U7685 ( .A1(n7498), .A2(n7497), .A3(n7734), .ZN(n7938) );
  OAI22_X1 U7686 ( .A1(n13953), .A2(n8109), .B1(n13950), .B2(n12110), .ZN(
        n7371) );
  NOR2_X1 U7687 ( .A1(n13953), .A2(n7373), .ZN(n7372) );
  INV_X1 U7688 ( .A(n13968), .ZN(n7373) );
  NOR2_X2 U7689 ( .A1(n13962), .A2(n14120), .ZN(n13947) );
  NAND2_X1 U7690 ( .A1(n8103), .A2(n8102), .ZN(n14038) );
  AND2_X1 U7691 ( .A1(n7871), .A2(n7870), .ZN(n11839) );
  INV_X1 U7692 ( .A(n14074), .ZN(n14179) );
  NAND2_X1 U7693 ( .A1(n7423), .A2(n7424), .ZN(n9435) );
  AOI21_X1 U7694 ( .B1(n7426), .B2(n7428), .A(n6597), .ZN(n7424) );
  NAND4_X1 U7695 ( .A1(n7292), .A2(n7289), .A3(n7503), .A4(n6524), .ZN(n7507)
         );
  NAND2_X1 U7696 ( .A1(n7968), .A2(n7967), .ZN(n8064) );
  OR2_X1 U7697 ( .A1(n7833), .A2(n7832), .ZN(n6884) );
  NOR2_X1 U7698 ( .A1(n14385), .A2(n6758), .ZN(n14338) );
  AOI21_X1 U7699 ( .B1(n14386), .B2(n14387), .A(P2_ADDR_REG_10__SCAN_IN), .ZN(
        n6758) );
  AOI21_X1 U7700 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14285), .A(n14284), .ZN(
        n14339) );
  OR2_X1 U7701 ( .A1(n14607), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6783) );
  INV_X1 U7702 ( .A(n12894), .ZN(n12816) );
  NAND2_X1 U7703 ( .A1(n13002), .A2(n7143), .ZN(n7142) );
  INV_X1 U7704 ( .A(n13003), .ZN(n7143) );
  NAND2_X1 U7705 ( .A1(n12009), .A2(n12008), .ZN(n7341) );
  AND2_X1 U7706 ( .A1(n8048), .A2(n8047), .ZN(n14108) );
  NAND2_X1 U7707 ( .A1(n11775), .A2(n11929), .ZN(n11776) );
  OAI21_X1 U7708 ( .B1(n9038), .B2(n9037), .A(n6647), .ZN(n6646) );
  NOR2_X1 U7709 ( .A1(n6969), .A2(n6515), .ZN(n6647) );
  INV_X1 U7710 ( .A(n9089), .ZN(n6652) );
  AND2_X1 U7711 ( .A1(n11836), .A2(n6947), .ZN(n6946) );
  INV_X1 U7712 ( .A(n11834), .ZN(n6947) );
  NOR2_X1 U7713 ( .A1(n11830), .A2(n11833), .ZN(n7298) );
  INV_X1 U7714 ( .A(n11830), .ZN(n7297) );
  INV_X1 U7715 ( .A(n11843), .ZN(n6942) );
  AND2_X1 U7716 ( .A1(n11848), .A2(n11847), .ZN(n11853) );
  MUX2_X1 U7717 ( .A(n8729), .B(n8728), .S(n9650), .Z(n8731) );
  AND2_X1 U7718 ( .A1(n7490), .A2(n11838), .ZN(n7293) );
  INV_X1 U7719 ( .A(n9175), .ZN(n7469) );
  NOR2_X1 U7720 ( .A1(n6996), .A2(n6995), .ZN(n6994) );
  NOR2_X1 U7721 ( .A1(n9174), .A2(n9175), .ZN(n6995) );
  AND2_X1 U7722 ( .A1(n6998), .A2(n6997), .ZN(n6996) );
  INV_X1 U7723 ( .A(n9193), .ZN(n6997) );
  NAND2_X1 U7724 ( .A1(n11871), .A2(n7947), .ZN(n6951) );
  NOR2_X1 U7725 ( .A1(n11869), .A2(n11866), .ZN(n7302) );
  NOR2_X1 U7726 ( .A1(n6952), .A2(n6615), .ZN(n6614) );
  MUX2_X1 U7727 ( .A(n8764), .B(n8763), .S(n10640), .Z(n8769) );
  AND2_X1 U7728 ( .A1(n7459), .A2(n9228), .ZN(n6984) );
  AND2_X1 U7729 ( .A1(n8778), .A2(n9650), .ZN(n6631) );
  NAND2_X1 U7730 ( .A1(n6962), .A2(n11889), .ZN(n6961) );
  OAI21_X1 U7731 ( .B1(n11885), .B2(n11884), .A(n11883), .ZN(n11887) );
  NAND2_X1 U7732 ( .A1(n11888), .A2(n6963), .ZN(n6960) );
  INV_X1 U7733 ( .A(n11889), .ZN(n6963) );
  NAND2_X1 U7734 ( .A1(n11903), .A2(n6956), .ZN(n6955) );
  INV_X1 U7735 ( .A(n11902), .ZN(n6956) );
  NOR2_X1 U7736 ( .A1(n7003), .A2(n7002), .ZN(n7001) );
  NOR2_X1 U7737 ( .A1(n7470), .A2(n9316), .ZN(n7002) );
  NOR2_X1 U7738 ( .A1(n6502), .A2(n7004), .ZN(n7003) );
  OAI21_X1 U7739 ( .B1(n8797), .B2(n12609), .A(n12600), .ZN(n8810) );
  NAND2_X1 U7740 ( .A1(n7284), .A2(n7283), .ZN(n6906) );
  NOR2_X1 U7741 ( .A1(n6975), .A2(n6554), .ZN(n6974) );
  AND2_X1 U7742 ( .A1(n9365), .A2(n9363), .ZN(n6975) );
  NOR2_X1 U7743 ( .A1(n11455), .A2(n7278), .ZN(n7277) );
  INV_X1 U7744 ( .A(n11242), .ZN(n7278) );
  AND2_X1 U7745 ( .A1(n8906), .A2(n8910), .ZN(n7198) );
  NAND2_X1 U7746 ( .A1(n11757), .A2(n11756), .ZN(n11763) );
  NAND2_X1 U7747 ( .A1(n7601), .A2(n11262), .ZN(n7603) );
  INV_X1 U7748 ( .A(n6791), .ZN(n6790) );
  OAI21_X1 U7749 ( .B1(n7580), .B2(n6792), .A(n7481), .ZN(n6791) );
  INV_X1 U7750 ( .A(n7582), .ZN(n6792) );
  NAND2_X1 U7751 ( .A1(n6879), .A2(n6877), .ZN(n7430) );
  AOI21_X1 U7752 ( .B1(n6880), .B2(n6883), .A(n6878), .ZN(n6877) );
  INV_X1 U7753 ( .A(n7482), .ZN(n6878) );
  AND2_X1 U7754 ( .A1(n14959), .A2(n9551), .ZN(n9552) );
  NOR2_X1 U7755 ( .A1(n8819), .A2(n8708), .ZN(n7100) );
  OAI21_X1 U7756 ( .B1(n11587), .B2(n14509), .A(n11586), .ZN(n12468) );
  NAND2_X1 U7757 ( .A1(n6755), .A2(n6600), .ZN(n7217) );
  AOI21_X1 U7758 ( .B1(n7390), .B2(n12226), .A(n7387), .ZN(n7386) );
  INV_X1 U7759 ( .A(n15076), .ZN(n7387) );
  NOR2_X1 U7760 ( .A1(n12457), .A2(n12225), .ZN(n7391) );
  INV_X1 U7761 ( .A(n7072), .ZN(n7071) );
  OAI21_X1 U7762 ( .B1(n12217), .B2(n7073), .A(n15138), .ZN(n7072) );
  INV_X1 U7763 ( .A(n8737), .ZN(n7073) );
  INV_X1 U7764 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8232) );
  INV_X1 U7765 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7415) );
  AND2_X1 U7766 ( .A1(n7406), .A2(n7080), .ZN(n7079) );
  INV_X1 U7767 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7080) );
  NOR2_X1 U7768 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n8229) );
  AND2_X1 U7769 ( .A1(n8226), .A2(n7408), .ZN(n7407) );
  INV_X1 U7770 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7408) );
  INV_X1 U7771 ( .A(n7023), .ZN(n7022) );
  OAI21_X1 U7772 ( .B1(n8487), .B2(n7024), .A(n8185), .ZN(n7023) );
  INV_X1 U7773 ( .A(n8171), .ZN(n7018) );
  INV_X1 U7774 ( .A(n13009), .ZN(n7183) );
  INV_X1 U7775 ( .A(n11525), .ZN(n7158) );
  NAND2_X1 U7776 ( .A1(n9459), .A2(n9431), .ZN(n9432) );
  NAND2_X1 U7777 ( .A1(n9430), .A2(n9449), .ZN(n9431) );
  INV_X1 U7778 ( .A(n7256), .ZN(n6851) );
  INV_X1 U7779 ( .A(n11449), .ZN(n7276) );
  OAI21_X1 U7780 ( .B1(n7277), .B2(n7276), .A(n11451), .ZN(n7275) );
  AND2_X1 U7781 ( .A1(n10693), .A2(n10692), .ZN(n6861) );
  INV_X1 U7782 ( .A(n10810), .ZN(n7273) );
  NAND2_X1 U7783 ( .A1(n6665), .A2(n6664), .ZN(n11254) );
  INV_X1 U7784 ( .A(n11033), .ZN(n6665) );
  NAND2_X1 U7785 ( .A1(n10962), .A2(n11238), .ZN(n11033) );
  INV_X1 U7786 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6858) );
  INV_X1 U7787 ( .A(n12020), .ZN(n7336) );
  INV_X1 U7788 ( .A(n12008), .ZN(n7337) );
  NOR2_X1 U7789 ( .A1(n7338), .A2(n6932), .ZN(n6931) );
  INV_X1 U7790 ( .A(n6934), .ZN(n6932) );
  INV_X1 U7791 ( .A(n7339), .ZN(n7338) );
  NAND2_X1 U7792 ( .A1(n6931), .A2(n6936), .ZN(n6929) );
  INV_X1 U7793 ( .A(n6905), .ZN(n6903) );
  NAND2_X1 U7794 ( .A1(n6898), .A2(n11926), .ZN(n6902) );
  INV_X1 U7795 ( .A(n11923), .ZN(n6898) );
  NAND2_X1 U7796 ( .A1(n6904), .A2(n11931), .ZN(n6901) );
  NAND2_X1 U7797 ( .A1(n6905), .A2(n11933), .ZN(n6904) );
  INV_X1 U7798 ( .A(n14242), .ZN(n7512) );
  INV_X1 U7799 ( .A(n11873), .ZN(n7359) );
  OR2_X1 U7800 ( .A1(n13738), .A2(n12024), .ZN(n11862) );
  AND2_X1 U7801 ( .A1(n11964), .A2(n7350), .ZN(n7349) );
  OR2_X1 U7802 ( .A1(n11963), .A2(n7351), .ZN(n7350) );
  INV_X1 U7803 ( .A(n8090), .ZN(n7351) );
  INV_X1 U7804 ( .A(n7788), .ZN(n7132) );
  INV_X1 U7805 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n7496) );
  NAND2_X1 U7806 ( .A1(n7452), .A2(n7451), .ZN(n7450) );
  INV_X1 U7807 ( .A(n7605), .ZN(n7452) );
  NAND2_X1 U7808 ( .A1(n7603), .A2(n7645), .ZN(n6897) );
  NAND2_X1 U7809 ( .A1(n7997), .A2(n7595), .ZN(n8000) );
  NAND2_X1 U7810 ( .A1(n6806), .A2(n6805), .ZN(n7593) );
  NOR2_X1 U7811 ( .A1(n6891), .A2(n10564), .ZN(n6805) );
  INV_X1 U7812 ( .A(n7593), .ZN(n7436) );
  NAND2_X1 U7813 ( .A1(n7591), .A2(n7592), .ZN(n7437) );
  INV_X1 U7814 ( .A(n7981), .ZN(n7592) );
  NAND2_X1 U7815 ( .A1(n7441), .A2(SI_18_), .ZN(n7439) );
  NAND2_X1 U7816 ( .A1(n6626), .A2(n6625), .ZN(n7587) );
  OAI21_X1 U7817 ( .B1(n7937), .B2(n10059), .A(n7935), .ZN(n6626) );
  NAND2_X1 U7818 ( .A1(n7566), .A2(n7565), .ZN(n7832) );
  NAND2_X2 U7819 ( .A1(n6786), .A2(n6785), .ZN(n7538) );
  NAND2_X1 U7820 ( .A1(n6620), .A2(n7418), .ZN(n6786) );
  NAND2_X1 U7821 ( .A1(n7525), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n6785) );
  NAND3_X1 U7822 ( .A1(n13218), .A2(n6876), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n6620) );
  OAI21_X1 U7823 ( .B1(n14298), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6550), .ZN(
        n7236) );
  XNOR2_X1 U7824 ( .A(n7236), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n14315) );
  AOI21_X1 U7825 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n15051), .A(n14280), .ZN(
        n14330) );
  AOI21_X1 U7826 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n14283), .A(n14282), .ZN(
        n14336) );
  NOR2_X1 U7827 ( .A1(n7058), .A2(n6566), .ZN(n6483) );
  NOR2_X1 U7828 ( .A1(n6499), .A2(n7059), .ZN(n7058) );
  AND2_X1 U7829 ( .A1(n7063), .A2(n7060), .ZN(n7053) );
  AND2_X1 U7830 ( .A1(n10737), .A2(n10646), .ZN(n8825) );
  NOR2_X1 U7831 ( .A1(n8453), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8478) );
  NAND2_X1 U7832 ( .A1(n12306), .A2(n12597), .ZN(n7065) );
  AND2_X1 U7833 ( .A1(n14418), .A2(n7039), .ZN(n7038) );
  NAND2_X1 U7834 ( .A1(n12391), .A2(n7040), .ZN(n7039) );
  AND3_X1 U7835 ( .A1(n8641), .A2(n8640), .A3(n8639), .ZN(n12364) );
  NAND2_X1 U7836 ( .A1(n8698), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8280) );
  NAND2_X1 U7837 ( .A1(n6621), .A2(n6522), .ZN(n7211) );
  AND2_X1 U7838 ( .A1(n7211), .A2(n7210), .ZN(n14991) );
  INV_X1 U7839 ( .A(n14992), .ZN(n7210) );
  NAND2_X1 U7840 ( .A1(n7222), .A2(n7221), .ZN(n6622) );
  NAND2_X1 U7841 ( .A1(n11202), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7221) );
  NAND2_X1 U7842 ( .A1(n6675), .A2(n6674), .ZN(n6755) );
  INV_X1 U7843 ( .A(n14449), .ZN(n6674) );
  INV_X1 U7844 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8226) );
  XNOR2_X1 U7845 ( .A(n7217), .B(n12543), .ZN(n14464) );
  NAND2_X1 U7846 ( .A1(n12608), .A2(n12251), .ZN(n12595) );
  OR2_X1 U7847 ( .A1(n12664), .A2(n12676), .ZN(n12641) );
  INV_X1 U7848 ( .A(n7075), .ZN(n7074) );
  OAI21_X1 U7849 ( .B1(n7077), .B2(n7076), .A(n8792), .ZN(n7075) );
  INV_X1 U7850 ( .A(n12450), .ZN(n12676) );
  AND2_X1 U7851 ( .A1(n8791), .A2(n8792), .ZN(n12674) );
  NAND2_X1 U7852 ( .A1(n12699), .A2(n12243), .ZN(n12683) );
  NAND2_X1 U7853 ( .A1(n12241), .A2(n12718), .ZN(n12710) );
  NOR2_X1 U7854 ( .A1(n12718), .A2(n7085), .ZN(n7084) );
  NAND2_X1 U7855 ( .A1(n8553), .A2(n12724), .ZN(n12731) );
  INV_X1 U7856 ( .A(n7089), .ZN(n7088) );
  AOI21_X1 U7857 ( .B1(n7089), .B2(n7091), .A(n7087), .ZN(n7086) );
  AOI21_X1 U7858 ( .B1(n7092), .B2(n8766), .A(n7090), .ZN(n7089) );
  INV_X1 U7859 ( .A(n12765), .ZN(n12773) );
  NAND2_X1 U7860 ( .A1(n7095), .A2(n7094), .ZN(n7093) );
  INV_X1 U7861 ( .A(n12789), .ZN(n7095) );
  NAND2_X1 U7862 ( .A1(n7093), .A2(n7092), .ZN(n12753) );
  AND2_X1 U7863 ( .A1(n12755), .A2(n8770), .ZN(n12765) );
  NAND2_X1 U7864 ( .A1(n15078), .A2(n12227), .ZN(n14492) );
  NAND2_X1 U7865 ( .A1(n7394), .A2(n7393), .ZN(n7392) );
  INV_X1 U7866 ( .A(n15109), .ZN(n7394) );
  INV_X1 U7867 ( .A(n7391), .ZN(n7389) );
  OR2_X1 U7868 ( .A1(n8362), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8377) );
  AND2_X1 U7869 ( .A1(n8737), .A2(n8736), .ZN(n12217) );
  INV_X1 U7870 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n11309) );
  INV_X1 U7871 ( .A(n11041), .ZN(n6736) );
  NAND2_X1 U7872 ( .A1(n10864), .A2(n10863), .ZN(n10869) );
  NAND2_X1 U7873 ( .A1(n10927), .A2(n10936), .ZN(n15179) );
  AND2_X1 U7874 ( .A1(n10941), .A2(n10940), .ZN(n15169) );
  NAND2_X1 U7875 ( .A1(n8586), .A2(n7077), .ZN(n12855) );
  NAND2_X1 U7876 ( .A1(n8512), .A2(n8511), .ZN(n12875) );
  AND2_X1 U7877 ( .A1(n9587), .A2(n9650), .ZN(n15142) );
  NAND2_X1 U7878 ( .A1(n9512), .A2(n9511), .ZN(n9766) );
  AND2_X1 U7879 ( .A1(n8261), .A2(n12950), .ZN(n8262) );
  AND4_X1 U7880 ( .A1(n8224), .A2(n8223), .A3(n8222), .A4(n8447), .ZN(n8225)
         );
  NOR2_X1 U7881 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n8224) );
  AND2_X1 U7882 ( .A1(n8714), .A2(n8716), .ZN(n8712) );
  INV_X1 U7883 ( .A(n8715), .ZN(n8714) );
  NAND2_X1 U7884 ( .A1(n8712), .A2(n8711), .ZN(n8848) );
  NAND2_X1 U7885 ( .A1(n6616), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7008) );
  NAND2_X1 U7886 ( .A1(n8571), .A2(n8196), .ZN(n6616) );
  NAND2_X1 U7887 ( .A1(n8571), .A2(n6594), .ZN(n7007) );
  NOR2_X1 U7888 ( .A1(n8572), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n8710) );
  INV_X1 U7889 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8709) );
  INV_X1 U7890 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8181) );
  NAND2_X1 U7891 ( .A1(n8470), .A2(n8180), .ZN(n8488) );
  NAND2_X1 U7892 ( .A1(n8488), .A2(n8487), .ZN(n8490) );
  INV_X1 U7893 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8491) );
  AND2_X1 U7894 ( .A1(n8173), .A2(n8172), .ZN(n8444) );
  NAND2_X1 U7895 ( .A1(n8169), .A2(n8168), .ZN(n8429) );
  NAND2_X1 U7896 ( .A1(n8429), .A2(n8428), .ZN(n8431) );
  OAI21_X1 U7897 ( .B1(n8319), .B2(n7012), .A(n7010), .ZN(n8335) );
  INV_X1 U7898 ( .A(n8153), .ZN(n7012) );
  NAND2_X1 U7899 ( .A1(n8303), .A2(n8151), .ZN(n8319) );
  NAND2_X1 U7900 ( .A1(n8319), .A2(n8318), .ZN(n8321) );
  NOR2_X1 U7901 ( .A1(n13595), .A2(n13593), .ZN(n9507) );
  XNOR2_X1 U7902 ( .A(n6472), .B(n14895), .ZN(n10183) );
  OR2_X1 U7903 ( .A1(n9353), .A2(n9352), .ZN(n9369) );
  NAND2_X1 U7904 ( .A1(n6684), .A2(n11230), .ZN(n11298) );
  AOI21_X1 U7905 ( .B1(n7164), .B2(n7162), .A(n6563), .ZN(n7161) );
  INV_X1 U7906 ( .A(n11370), .ZN(n7165) );
  CLKBUF_X1 U7907 ( .A(n11229), .Z(n6684) );
  INV_X1 U7908 ( .A(n10228), .ZN(n7186) );
  NOR2_X1 U7909 ( .A1(n13092), .A2(n7154), .ZN(n7153) );
  INV_X1 U7910 ( .A(n13069), .ZN(n7154) );
  AND2_X1 U7911 ( .A1(n7151), .A2(n6582), .ZN(n7149) );
  NAND2_X1 U7912 ( .A1(n7252), .A2(n6482), .ZN(n7250) );
  NAND2_X1 U7913 ( .A1(n12205), .A2(n7253), .ZN(n7252) );
  OR2_X1 U7914 ( .A1(n13283), .A2(n7254), .ZN(n7253) );
  NAND2_X1 U7915 ( .A1(n6482), .A2(n12204), .ZN(n7251) );
  NAND2_X1 U7916 ( .A1(n13284), .A2(n13283), .ZN(n13282) );
  INV_X1 U7917 ( .A(n7262), .ZN(n7261) );
  OAI21_X1 U7918 ( .B1(n13324), .B2(n7263), .A(n12201), .ZN(n7262) );
  AND2_X1 U7919 ( .A1(n12201), .A2(n12199), .ZN(n13309) );
  NAND2_X1 U7920 ( .A1(n6834), .A2(n6835), .ZN(n13325) );
  NAND2_X1 U7921 ( .A1(n13325), .A2(n13324), .ZN(n13323) );
  AOI21_X1 U7922 ( .B1(n7271), .B2(n7267), .A(n6491), .ZN(n7266) );
  NAND2_X1 U7923 ( .A1(n6866), .A2(n6868), .ZN(n13372) );
  INV_X1 U7924 ( .A(n6872), .ZN(n6871) );
  OAI22_X1 U7925 ( .A1(n12152), .A2(n6873), .B1(n13165), .B2(n13394), .ZN(
        n6872) );
  NAND2_X1 U7926 ( .A1(n6504), .A2(n12151), .ZN(n6873) );
  NAND2_X1 U7927 ( .A1(n7242), .A2(n12188), .ZN(n7241) );
  INV_X1 U7928 ( .A(n12187), .ZN(n7242) );
  INV_X1 U7929 ( .A(n12188), .ZN(n7243) );
  NAND2_X1 U7930 ( .A1(n13403), .A2(n12187), .ZN(n7240) );
  AND2_X1 U7931 ( .A1(n6832), .A2(n6509), .ZN(n13403) );
  NAND2_X1 U7932 ( .A1(n11727), .A2(n11660), .ZN(n7256) );
  AOI21_X1 U7933 ( .B1(n11455), .B2(n6824), .A(n6517), .ZN(n6823) );
  INV_X1 U7934 ( .A(n11252), .ZN(n6824) );
  NAND2_X1 U7935 ( .A1(n11028), .A2(n11027), .ZN(n11030) );
  NOR2_X1 U7936 ( .A1(n11027), .A2(n7248), .ZN(n7247) );
  NAND2_X1 U7937 ( .A1(n10719), .A2(n10966), .ZN(n6846) );
  AND2_X1 U7938 ( .A1(n10718), .A2(n10966), .ZN(n7248) );
  OR2_X1 U7939 ( .A1(n10719), .A2(n10718), .ZN(n10967) );
  NOR2_X1 U7940 ( .A1(n10813), .A2(n6844), .ZN(n6843) );
  INV_X1 U7941 ( .A(n10673), .ZN(n6844) );
  OR2_X1 U7942 ( .A1(n10803), .A2(n10692), .ZN(n6864) );
  NAND2_X1 U7943 ( .A1(n7245), .A2(n10669), .ZN(n6830) );
  INV_X1 U7944 ( .A(n10668), .ZN(n7246) );
  OAI21_X1 U7945 ( .B1(n10874), .B2(n10667), .A(n6831), .ZN(n10892) );
  INV_X1 U7946 ( .A(n10723), .ZN(n13405) );
  OR2_X1 U7947 ( .A1(n10628), .A2(n9231), .ZN(n9235) );
  INV_X1 U7948 ( .A(n10827), .ZN(n14909) );
  AND2_X1 U7949 ( .A1(n10187), .A2(n10200), .ZN(n14874) );
  NAND2_X1 U7950 ( .A1(n6854), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8899) );
  NOR2_X1 U7951 ( .A1(n9194), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n6855) );
  NOR2_X1 U7952 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n8873) );
  NOR2_X1 U7953 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n8872) );
  AND2_X1 U7954 ( .A1(n9492), .A2(n9467), .ZN(n9833) );
  INV_X1 U7955 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8907) );
  AOI21_X1 U7956 ( .B1(n7331), .B2(n7334), .A(n7328), .ZN(n7327) );
  INV_X1 U7957 ( .A(n13697), .ZN(n7334) );
  AOI21_X1 U7958 ( .B1(n13604), .B2(n12116), .A(n12130), .ZN(n7312) );
  AND2_X1 U7959 ( .A1(n11685), .A2(n11683), .ZN(n6937) );
  NAND2_X1 U7960 ( .A1(n6910), .A2(n6914), .ZN(n11401) );
  AND2_X1 U7961 ( .A1(n6915), .A2(n11354), .ZN(n6914) );
  NAND2_X1 U7962 ( .A1(n6916), .A2(n6919), .ZN(n6915) );
  OR2_X1 U7963 ( .A1(n7853), .A2(n7852), .ZN(n7873) );
  INV_X1 U7964 ( .A(n6937), .ZN(n6936) );
  OAI22_X1 U7965 ( .A1(n9615), .A2(n9614), .B1(n10131), .B2(n11396), .ZN(n9617) );
  INV_X1 U7966 ( .A(n14197), .ZN(n13894) );
  NAND2_X1 U7967 ( .A1(n13947), .A2(n14203), .ZN(n13936) );
  AND2_X1 U7968 ( .A1(n7644), .A2(n8039), .ZN(n13953) );
  NAND2_X1 U7969 ( .A1(n13961), .A2(n13968), .ZN(n13960) );
  NAND2_X1 U7970 ( .A1(n13979), .A2(n13980), .ZN(n13978) );
  AOI21_X1 U7971 ( .B1(n7378), .B2(n14039), .A(n6546), .ZN(n7376) );
  OR2_X1 U7972 ( .A1(n14038), .A2(n14039), .ZN(n14036) );
  NOR2_X1 U7973 ( .A1(n11975), .A2(n7125), .ZN(n7124) );
  INV_X1 U7974 ( .A(n11879), .ZN(n7125) );
  AND2_X1 U7975 ( .A1(n11878), .A2(n11879), .ZN(n14051) );
  INV_X1 U7976 ( .A(n14051), .ZN(n14053) );
  AND2_X1 U7977 ( .A1(n7139), .A2(n7934), .ZN(n7138) );
  INV_X1 U7978 ( .A(n14091), .ZN(n7139) );
  OR2_X1 U7979 ( .A1(n11611), .A2(n11610), .ZN(n7140) );
  AOI21_X1 U7980 ( .B1(n7366), .B2(n11968), .A(n6549), .ZN(n7364) );
  INV_X1 U7981 ( .A(n11969), .ZN(n11467) );
  NOR2_X1 U7982 ( .A1(n11467), .A2(n7367), .ZN(n7366) );
  INV_X1 U7983 ( .A(n8099), .ZN(n7367) );
  AND2_X1 U7984 ( .A1(n8069), .A2(n11756), .ZN(n11984) );
  OR2_X1 U7985 ( .A1(n11569), .A2(n11968), .ZN(n11571) );
  AND2_X1 U7986 ( .A1(n11858), .A2(n11857), .ZN(n11968) );
  AOI21_X1 U7987 ( .B1(n7112), .B2(n7114), .A(n7110), .ZN(n7109) );
  AND2_X1 U7988 ( .A1(n14402), .A2(n14407), .ZN(n14400) );
  NAND2_X1 U7989 ( .A1(n10579), .A2(n7788), .ZN(n11011) );
  NAND2_X1 U7990 ( .A1(n10579), .A2(n7131), .ZN(n11012) );
  CLKBUF_X1 U7991 ( .A(n11006), .Z(n6683) );
  NAND2_X1 U7992 ( .A1(n7635), .A2(n7634), .ZN(n14120) );
  NAND2_X1 U7993 ( .A1(n13598), .A2(n7923), .ZN(n7650) );
  NAND2_X1 U7994 ( .A1(n7972), .A2(n7971), .ZN(n13621) );
  NAND2_X1 U7995 ( .A1(n7942), .A2(n7941), .ZN(n14088) );
  NAND2_X1 U7996 ( .A1(n8145), .A2(n14560), .ZN(n14724) );
  INV_X1 U7997 ( .A(n14664), .ZN(n14728) );
  NOR2_X1 U7998 ( .A1(n14264), .A2(n8113), .ZN(n10028) );
  OR2_X1 U7999 ( .A1(n14254), .A2(n8119), .ZN(n8121) );
  XNOR2_X1 U8000 ( .A(n9435), .B(n9434), .ZN(n11998) );
  INV_X1 U8001 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7508) );
  INV_X1 U8002 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7502) );
  NOR2_X1 U8003 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n7500) );
  NAND2_X1 U8004 ( .A1(n7953), .A2(n7952), .ZN(n8117) );
  AND2_X1 U8005 ( .A1(n7952), .A2(n6965), .ZN(n7344) );
  NAND2_X1 U8006 ( .A1(n6966), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7968) );
  AND2_X1 U8007 ( .A1(n7952), .A2(n6965), .ZN(n6964) );
  INV_X1 U8008 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7967) );
  NAND2_X1 U8009 ( .A1(n7587), .A2(n10098), .ZN(n7442) );
  INV_X1 U8010 ( .A(n7948), .ZN(n7441) );
  NAND2_X1 U8011 ( .A1(n7438), .A2(SI_18_), .ZN(n7443) );
  INV_X1 U8012 ( .A(n7587), .ZN(n7438) );
  NAND2_X1 U8013 ( .A1(n7904), .A2(n7582), .ZN(n7922) );
  OAI21_X1 U8014 ( .B1(n7833), .B2(n6883), .A(n6880), .ZN(n7862) );
  XNOR2_X1 U8015 ( .A(n7833), .B(n7832), .ZN(n9768) );
  NAND2_X1 U8016 ( .A1(n7422), .A2(n7560), .ZN(n7821) );
  NAND2_X1 U8017 ( .A1(n7804), .A2(n7558), .ZN(n7422) );
  NAND2_X1 U8018 ( .A1(n7534), .A2(n7533), .ZN(n7715) );
  AND2_X1 U8019 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n6760), .ZN(n14304) );
  NAND2_X1 U8020 ( .A1(n14382), .A2(n14381), .ZN(n7230) );
  INV_X1 U8021 ( .A(n6759), .ZN(n14318) );
  OAI21_X1 U8022 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14287), .A(n14286), .ZN(
        n14292) );
  NOR2_X1 U8023 ( .A1(n14611), .A2(n6779), .ZN(n6780) );
  OR2_X1 U8024 ( .A1(n6777), .A2(n6495), .ZN(n6773) );
  NAND3_X1 U8025 ( .A1(n9512), .A2(n8859), .A3(n8858), .ZN(n9607) );
  AOI21_X1 U8026 ( .B1(n12419), .B2(n9543), .A(n7045), .ZN(n7044) );
  NAND2_X1 U8027 ( .A1(n7057), .A2(n6499), .ZN(n6718) );
  NAND2_X1 U8028 ( .A1(n8673), .A2(n8672), .ZN(n12589) );
  NAND2_X1 U8029 ( .A1(n9530), .A2(n9529), .ZN(n10954) );
  AND4_X1 U8030 ( .A1(n8567), .A2(n8566), .A3(n8565), .A4(n8564), .ZN(n12322)
         );
  AND4_X1 U8031 ( .A1(n8597), .A2(n8596), .A3(n8595), .A4(n8594), .ZN(n12704)
         );
  NAND2_X1 U8032 ( .A1(n7047), .A2(n12280), .ZN(n14432) );
  INV_X1 U8033 ( .A(n14429), .ZN(n12280) );
  NAND2_X1 U8034 ( .A1(n10954), .A2(n6508), .ZN(n11215) );
  NOR2_X1 U8035 ( .A1(n8418), .A2(n8417), .ZN(n15241) );
  NAND2_X1 U8036 ( .A1(n6599), .A2(n9524), .ZN(n10735) );
  AND4_X1 U8037 ( .A1(n8552), .A2(n8551), .A3(n8550), .A4(n8549), .ZN(n12715)
         );
  OR2_X1 U8038 ( .A1(n12418), .A2(n12419), .ZN(n12420) );
  AND2_X1 U8039 ( .A1(n9578), .A2(n9577), .ZN(n14965) );
  AND4_X1 U8040 ( .A1(n8533), .A2(n8532), .A3(n8531), .A4(n8530), .ZN(n12439)
         );
  INV_X1 U8041 ( .A(n14971), .ZN(n14436) );
  NAND2_X1 U8042 ( .A1(n6627), .A2(n15199), .ZN(n7025) );
  AND2_X1 U8043 ( .A1(n6676), .A2(n6677), .ZN(n6694) );
  INV_X1 U8044 ( .A(n12322), .ZN(n12726) );
  INV_X1 U8045 ( .A(n14495), .ZN(n12456) );
  NAND2_X1 U8046 ( .A1(n6752), .A2(n6523), .ZN(n7224) );
  INV_X1 U8047 ( .A(n7222), .ZN(n11196) );
  XNOR2_X1 U8048 ( .A(n6622), .B(n11422), .ZN(n11197) );
  NAND2_X1 U8049 ( .A1(n7220), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7219) );
  INV_X1 U8050 ( .A(n12467), .ZN(n7220) );
  AND2_X1 U8051 ( .A1(n9660), .A2(n12516), .ZN(n15058) );
  NOR2_X1 U8052 ( .A1(n14483), .A2(n6753), .ZN(n12536) );
  NOR2_X1 U8053 ( .A1(n14470), .A2(n12534), .ZN(n6753) );
  AND2_X1 U8054 ( .A1(n9660), .A2(n9658), .ZN(n14480) );
  INV_X1 U8055 ( .A(n12813), .ZN(n6655) );
  NAND2_X1 U8056 ( .A1(n8591), .A2(n8590), .ZN(n12694) );
  NAND2_X1 U8057 ( .A1(n10866), .A2(n10865), .ZN(n15104) );
  NAND2_X1 U8058 ( .A1(n10869), .A2(n15104), .ZN(n15204) );
  AND2_X1 U8059 ( .A1(n15173), .A2(n15242), .ZN(n12695) );
  NAND2_X1 U8060 ( .A1(n7028), .A2(n8697), .ZN(n12894) );
  CLKBUF_X1 U8061 ( .A(n8238), .Z(n6724) );
  NAND2_X1 U8062 ( .A1(n13138), .A2(n13009), .ZN(n13039) );
  NAND2_X1 U8063 ( .A1(n9319), .A2(n9318), .ZN(n13476) );
  NAND2_X1 U8064 ( .A1(n9246), .A2(n9245), .ZN(n13500) );
  NAND2_X1 U8065 ( .A1(n7180), .A2(n7179), .ZN(n7178) );
  OAI21_X1 U8066 ( .B1(n7180), .B2(n13042), .A(n7176), .ZN(n7175) );
  INV_X1 U8067 ( .A(n14895), .ZN(n10677) );
  NAND2_X1 U8068 ( .A1(n13598), .A2(n9436), .ZN(n6685) );
  NAND2_X1 U8069 ( .A1(n9304), .A2(n9303), .ZN(n13331) );
  NAND2_X1 U8070 ( .A1(n9180), .A2(n9179), .ZN(n13525) );
  NAND2_X1 U8071 ( .A1(n6988), .A2(n6985), .ZN(n9491) );
  AND2_X1 U8072 ( .A1(n6989), .A2(n9429), .ZN(n6986) );
  AOI211_X1 U8073 ( .C1(n13438), .C2(n12179), .A(n14849), .B(n13225), .ZN(
        n13437) );
  OAI21_X1 U8074 ( .B1(n13011), .B2(n13072), .A(n12176), .ZN(n12177) );
  XNOR2_X1 U8075 ( .A(n6847), .B(n12173), .ZN(n12178) );
  NAND2_X1 U8076 ( .A1(n9128), .A2(n9127), .ZN(n14522) );
  AND2_X1 U8077 ( .A1(n14867), .A2(n10776), .ZN(n13425) );
  AOI21_X1 U8078 ( .B1(n13229), .B2(n6814), .A(n6811), .ZN(n6810) );
  NOR2_X1 U8079 ( .A1(n12208), .A2(n12207), .ZN(n6811) );
  AND2_X1 U8080 ( .A1(n10211), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14886) );
  INV_X1 U8081 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10627) );
  AND2_X1 U8082 ( .A1(n14254), .A2(n14250), .ZN(n8140) );
  NAND2_X1 U8083 ( .A1(n7623), .A2(n7622), .ZN(n13939) );
  NOR2_X1 U8084 ( .A1(n14546), .A2(n7340), .ZN(n7339) );
  INV_X1 U8085 ( .A(n12012), .ZN(n7340) );
  NAND2_X1 U8086 ( .A1(n7341), .A2(n12012), .ZN(n14547) );
  NAND2_X1 U8087 ( .A1(n9622), .A2(n7305), .ZN(n7304) );
  INV_X1 U8088 ( .A(n9623), .ZN(n7305) );
  NAND2_X1 U8089 ( .A1(n7617), .A2(n7616), .ZN(n13915) );
  OAI21_X1 U8090 ( .B1(n12121), .B2(n10075), .A(n10074), .ZN(n10033) );
  NAND2_X1 U8091 ( .A1(n6933), .A2(n6934), .ZN(n12009) );
  OR2_X1 U8092 ( .A1(n11650), .A2(n6936), .ZN(n6933) );
  INV_X1 U8093 ( .A(n13740), .ZN(n14550) );
  NAND2_X1 U8094 ( .A1(n9641), .A2(n14667), .ZN(n14554) );
  INV_X1 U8095 ( .A(n13934), .ZN(n6799) );
  NAND2_X1 U8096 ( .A1(n13594), .A2(n7923), .ZN(n6802) );
  AND2_X1 U8097 ( .A1(n7956), .A2(n7955), .ZN(n14074) );
  AND2_X1 U8098 ( .A1(n10520), .A2(n14564), .ZN(n14686) );
  NAND2_X1 U8099 ( .A1(n14764), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n7356) );
  INV_X1 U8100 ( .A(n14766), .ZN(n14764) );
  NAND2_X1 U8101 ( .A1(n8115), .A2(n8114), .ZN(n14107) );
  AOI21_X1 U8102 ( .B1(n13911), .B2(n14664), .A(n8077), .ZN(n8115) );
  INV_X1 U8103 ( .A(n13939), .ZN(n14203) );
  NAND2_X1 U8104 ( .A1(n7664), .A2(n7663), .ZN(n14212) );
  OR2_X1 U8105 ( .A1(n14254), .A2(n14250), .ZN(n9746) );
  INV_X1 U8106 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10629) );
  XNOR2_X1 U8107 ( .A(n14332), .B(n7229), .ZN(n14384) );
  INV_X1 U8108 ( .A(n14333), .ZN(n7229) );
  INV_X1 U8109 ( .A(n14602), .ZN(n7225) );
  INV_X1 U8110 ( .A(n6778), .ZN(n6777) );
  OAI21_X1 U8111 ( .B1(n6783), .B2(n6779), .A(n14611), .ZN(n6778) );
  OR2_X1 U8112 ( .A1(n14606), .A2(n6779), .ZN(n6774) );
  NAND2_X1 U8113 ( .A1(n14606), .A2(n6783), .ZN(n6781) );
  NAND2_X1 U8114 ( .A1(n14353), .A2(n6767), .ZN(n6766) );
  OR2_X1 U8115 ( .A1(n6771), .A2(n6770), .ZN(n6769) );
  INV_X1 U8116 ( .A(n6768), .ZN(n6767) );
  OAI21_X1 U8117 ( .B1(n14347), .B2(n6771), .A(n6768), .ZN(n14354) );
  NAND2_X1 U8118 ( .A1(n11772), .A2(n11771), .ZN(n11777) );
  NOR2_X1 U8119 ( .A1(n6501), .A2(n6971), .ZN(n6969) );
  MUX2_X1 U8120 ( .A(n11794), .B(n11793), .S(n11929), .Z(n11795) );
  NAND2_X1 U8121 ( .A1(n6970), .A2(n6535), .ZN(n9091) );
  NAND2_X1 U8122 ( .A1(n6501), .A2(n6971), .ZN(n6968) );
  NOR2_X1 U8123 ( .A1(n11816), .A2(n11819), .ZN(n7300) );
  INV_X1 U8124 ( .A(n11816), .ZN(n7299) );
  NOR2_X1 U8125 ( .A1(n7455), .A2(n7454), .ZN(n7005) );
  INV_X1 U8126 ( .A(n6575), .ZN(n6998) );
  NAND2_X1 U8127 ( .A1(n6941), .A2(n6939), .ZN(n11856) );
  AND2_X1 U8128 ( .A1(n11842), .A2(n6940), .ZN(n6939) );
  NAND2_X1 U8129 ( .A1(n6511), .A2(n6946), .ZN(n6940) );
  AND2_X1 U8130 ( .A1(n11968), .A2(n7479), .ZN(n7490) );
  NAND2_X1 U8131 ( .A1(n8751), .A2(n15094), .ZN(n6715) );
  NOR2_X1 U8132 ( .A1(n11871), .A2(n7362), .ZN(n6952) );
  NOR2_X1 U8133 ( .A1(n7301), .A2(n11868), .ZN(n6615) );
  INV_X1 U8134 ( .A(n11866), .ZN(n7301) );
  NOR2_X1 U8135 ( .A1(n7468), .A2(n7469), .ZN(n7467) );
  NOR2_X1 U8136 ( .A1(n11873), .A2(n6949), .ZN(n6948) );
  INV_X1 U8137 ( .A(n6951), .ZN(n6949) );
  OR2_X1 U8138 ( .A1(n8772), .A2(n9650), .ZN(n6609) );
  NAND2_X1 U8139 ( .A1(n6982), .A2(n6525), .ZN(n6980) );
  NAND2_X1 U8140 ( .A1(n6588), .A2(n7085), .ZN(n6628) );
  NOR2_X1 U8141 ( .A1(n11893), .A2(n11891), .ZN(n7286) );
  NAND2_X1 U8142 ( .A1(n12674), .A2(n8788), .ZN(n6749) );
  NAND2_X1 U8143 ( .A1(n9277), .A2(n6527), .ZN(n7472) );
  NAND2_X1 U8144 ( .A1(n6958), .A2(n11902), .ZN(n6957) );
  AND2_X1 U8145 ( .A1(n12565), .A2(n10640), .ZN(n6712) );
  NOR2_X1 U8146 ( .A1(n6604), .A2(n10640), .ZN(n6603) );
  INV_X1 U8147 ( .A(n8813), .ZN(n6604) );
  NAND2_X1 U8148 ( .A1(n7000), .A2(n6999), .ZN(n9347) );
  NAND2_X1 U8149 ( .A1(n11754), .A2(n11753), .ZN(n11757) );
  AND2_X1 U8150 ( .A1(n15158), .A2(n12214), .ZN(n15123) );
  NAND2_X1 U8151 ( .A1(n12461), .A2(n6719), .ZN(n8726) );
  INV_X1 U8152 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8876) );
  INV_X1 U8153 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8905) );
  INV_X1 U8154 ( .A(n10518), .ZN(n11766) );
  OAI21_X1 U8155 ( .B1(n11910), .B2(n7284), .A(n6559), .ZN(n6938) );
  INV_X1 U8156 ( .A(n7446), .ZN(n7445) );
  OAI21_X1 U8157 ( .B1(n7448), .B2(n7447), .A(SI_27_), .ZN(n7446) );
  NAND2_X1 U8158 ( .A1(n7607), .A2(n6896), .ZN(n7444) );
  NAND2_X1 U8159 ( .A1(n7645), .A2(SI_24_), .ZN(n6894) );
  NOR2_X1 U8160 ( .A1(n7630), .A2(n7449), .ZN(n7448) );
  INV_X1 U8161 ( .A(n7450), .ZN(n7449) );
  INV_X1 U8162 ( .A(n7965), .ZN(n6892) );
  OAI21_X1 U8163 ( .B1(n6488), .B2(n6891), .A(n10564), .ZN(n6890) );
  AOI21_X1 U8164 ( .B1(n7832), .B2(n7566), .A(n6886), .ZN(n6885) );
  INV_X1 U8165 ( .A(n7486), .ZN(n6886) );
  NOR2_X1 U8166 ( .A1(n7820), .A2(n7803), .ZN(n7419) );
  INV_X1 U8167 ( .A(n7560), .ZN(n7421) );
  NOR2_X1 U8168 ( .A1(n7805), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n7835) );
  NAND2_X1 U8169 ( .A1(n7417), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6733) );
  INV_X1 U8170 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n7745) );
  OAI21_X1 U8171 ( .B1(n7538), .B2(P2_DATAO_REG_3__SCAN_IN), .A(n6732), .ZN(
        n7535) );
  NAND2_X1 U8172 ( .A1(n8964), .A2(n7538), .ZN(n6732) );
  INV_X1 U8173 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6876) );
  INV_X1 U8174 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7524) );
  NOR2_X1 U8175 ( .A1(n14271), .A2(n14272), .ZN(n14273) );
  OR2_X1 U8176 ( .A1(n6508), .A2(n7050), .ZN(n7049) );
  INV_X1 U8177 ( .A(n9536), .ZN(n7050) );
  INV_X1 U8178 ( .A(n12390), .ZN(n7040) );
  NOR2_X1 U8179 ( .A1(n7041), .A2(n7036), .ZN(n7035) );
  INV_X1 U8180 ( .A(n12270), .ZN(n7036) );
  NOR2_X1 U8181 ( .A1(n8816), .A2(n7097), .ZN(n7096) );
  INV_X1 U8182 ( .A(n8822), .ZN(n7097) );
  NAND2_X1 U8183 ( .A1(n12558), .A2(n8842), .ZN(n7099) );
  NAND2_X1 U8184 ( .A1(n6681), .A2(n6680), .ZN(n6679) );
  NOR2_X1 U8185 ( .A1(n12574), .A2(n8841), .ZN(n6681) );
  NAND2_X1 U8186 ( .A1(n8306), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10432) );
  OAI21_X1 U8187 ( .B1(n14439), .B2(n12873), .A(n14440), .ZN(n12544) );
  OR2_X1 U8188 ( .A1(n12602), .A2(n12584), .ZN(n8806) );
  OR2_X1 U8189 ( .A1(n8618), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8628) );
  INV_X1 U8190 ( .A(n8786), .ZN(n7076) );
  INV_X1 U8191 ( .A(n12755), .ZN(n7090) );
  INV_X1 U8192 ( .A(n7092), .ZN(n7091) );
  NAND2_X1 U8193 ( .A1(n8434), .A2(n7384), .ZN(n14488) );
  OR2_X1 U8194 ( .A1(n12217), .A2(n15156), .ZN(n15158) );
  NAND2_X1 U8195 ( .A1(n12215), .A2(n7396), .ZN(n15156) );
  AND2_X1 U8196 ( .A1(n8726), .A2(n8727), .ZN(n11046) );
  AND2_X1 U8197 ( .A1(n6693), .A2(n12445), .ZN(n6723) );
  NOR2_X1 U8198 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n8223) );
  INV_X1 U8199 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8446) );
  OR2_X1 U8200 ( .A1(n8399), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8410) );
  INV_X1 U8201 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8385) );
  NAND2_X1 U8202 ( .A1(n8218), .A2(n7405), .ZN(n7404) );
  INV_X1 U8203 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7405) );
  NAND2_X1 U8204 ( .A1(n7403), .A2(n8218), .ZN(n8356) );
  INV_X1 U8205 ( .A(n8337), .ZN(n7403) );
  OR2_X1 U8206 ( .A1(n13038), .A2(n7183), .ZN(n7182) );
  AND2_X1 U8207 ( .A1(n9007), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9021) );
  NOR2_X1 U8208 ( .A1(n7168), .A2(n7167), .ZN(n7166) );
  INV_X1 U8209 ( .A(n11725), .ZN(n7168) );
  INV_X1 U8210 ( .A(n11728), .ZN(n7167) );
  AOI21_X1 U8211 ( .B1(n6974), .B2(n6976), .A(n6481), .ZN(n6973) );
  NOR2_X1 U8212 ( .A1(n9365), .A2(n9363), .ZN(n6976) );
  CLKBUF_X3 U8213 ( .A(n9057), .Z(n9462) );
  NAND2_X1 U8214 ( .A1(n6565), .A2(n12197), .ZN(n6835) );
  INV_X1 U8215 ( .A(n12194), .ZN(n6836) );
  NOR2_X1 U8216 ( .A1(n7268), .A2(n6869), .ZN(n6867) );
  INV_X1 U8217 ( .A(n13357), .ZN(n7272) );
  OAI21_X1 U8218 ( .B1(n9464), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9466) );
  INV_X1 U8219 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9465) );
  NAND2_X1 U8220 ( .A1(n7198), .A2(n7197), .ZN(n7196) );
  NOR2_X1 U8221 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n7197) );
  INV_X1 U8222 ( .A(n7198), .ZN(n7195) );
  OR2_X1 U8223 ( .A1(n9125), .A2(n9124), .ZN(n9142) );
  OR2_X1 U8224 ( .A1(n9125), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n9053) );
  NAND2_X1 U8225 ( .A1(n6925), .A2(n6923), .ZN(n6922) );
  INV_X1 U8226 ( .A(n13688), .ZN(n6923) );
  INV_X1 U8227 ( .A(n6925), .ZN(n6924) );
  AOI21_X1 U8228 ( .B1(n13697), .B2(n7333), .A(n7332), .ZN(n7331) );
  INV_X1 U8229 ( .A(n13612), .ZN(n7328) );
  NOR2_X1 U8230 ( .A1(n13633), .A2(n6926), .ZN(n6925) );
  INV_X1 U8231 ( .A(n12064), .ZN(n6926) );
  NAND2_X1 U8232 ( .A1(n7322), .A2(n7325), .ZN(n7319) );
  NAND2_X1 U8233 ( .A1(n7314), .A2(n11159), .ZN(n7322) );
  INV_X1 U8234 ( .A(n11158), .ZN(n7325) );
  AND2_X1 U8235 ( .A1(n13928), .A2(n8110), .ZN(n13923) );
  NOR2_X1 U8236 ( .A1(n8105), .A2(n7379), .ZN(n7378) );
  INV_X1 U8237 ( .A(n8104), .ZN(n7379) );
  INV_X1 U8238 ( .A(n11789), .ZN(n11957) );
  OR2_X1 U8239 ( .A1(n14703), .A2(n13770), .ZN(n11791) );
  NAND2_X1 U8240 ( .A1(n7205), .A2(n9684), .ZN(n7102) );
  NAND2_X1 U8241 ( .A1(n9685), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7103) );
  NAND2_X1 U8242 ( .A1(n7107), .A2(n7106), .ZN(n10995) );
  INV_X1 U8243 ( .A(n7427), .ZN(n7426) );
  OAI21_X1 U8244 ( .B1(n8043), .B2(n7428), .A(n9415), .ZN(n7427) );
  INV_X1 U8245 ( .A(n8046), .ZN(n7428) );
  NAND2_X1 U8246 ( .A1(n7604), .A2(n6897), .ZN(n8027) );
  NAND2_X1 U8247 ( .A1(n8000), .A2(n6584), .ZN(n7434) );
  AOI21_X1 U8248 ( .B1(n6790), .B2(n6792), .A(n6789), .ZN(n6788) );
  INV_X1 U8249 ( .A(n7586), .ZN(n6789) );
  NOR2_X2 U8250 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n7907) );
  NAND2_X1 U8251 ( .A1(n7430), .A2(n7574), .ZN(n7883) );
  INV_X1 U8252 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n10376) );
  AOI21_X1 U8253 ( .B1(n6885), .B2(n6882), .A(n6881), .ZN(n6880) );
  INV_X1 U8254 ( .A(n7570), .ZN(n6881) );
  INV_X1 U8255 ( .A(n7566), .ZN(n6882) );
  INV_X1 U8256 ( .A(n6885), .ZN(n6883) );
  OR2_X1 U8257 ( .A1(n7849), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n7909) );
  OR2_X1 U8258 ( .A1(n7791), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n7805) );
  INV_X1 U8259 ( .A(n7774), .ZN(n7551) );
  OR2_X1 U8260 ( .A1(n7776), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n7791) );
  XNOR2_X1 U8261 ( .A(n7552), .B(SI_7_), .ZN(n7774) );
  INV_X1 U8262 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7733) );
  NAND2_X1 U8263 ( .A1(n7538), .A2(n8147), .ZN(n6784) );
  AOI21_X1 U8264 ( .B1(n6761), .B2(n14304), .A(n7235), .ZN(n14300) );
  AND2_X1 U8265 ( .A1(n14268), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7235) );
  INV_X1 U8266 ( .A(n14302), .ZN(n6761) );
  INV_X1 U8267 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14268) );
  AND2_X1 U8268 ( .A1(n7234), .A2(n7233), .ZN(n14270) );
  NAND2_X1 U8269 ( .A1(n14269), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7233) );
  OR2_X1 U8270 ( .A1(n14300), .A2(n14301), .ZN(n7234) );
  NOR2_X1 U8271 ( .A1(n14279), .A2(n14278), .ZN(n14297) );
  OR2_X1 U8272 ( .A1(n10763), .A2(n10762), .ZN(n7303) );
  INV_X1 U8273 ( .A(n12118), .ZN(n12131) );
  INV_X1 U8274 ( .A(n12347), .ZN(n7061) );
  NOR2_X1 U8275 ( .A1(n8433), .A2(n8432), .ZN(n14964) );
  XNOR2_X1 U8276 ( .A(n12296), .B(n6719), .ZN(n9531) );
  NAND2_X1 U8277 ( .A1(n14432), .A2(n12282), .ZN(n12355) );
  NAND2_X1 U8278 ( .A1(n8249), .A2(n8248), .ZN(n8592) );
  INV_X1 U8279 ( .A(n8579), .ZN(n8249) );
  OR2_X1 U8280 ( .A1(n8592), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8605) );
  NAND2_X1 U8281 ( .A1(n15188), .A2(n10738), .ZN(n15178) );
  OR2_X1 U8282 ( .A1(n8562), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8579) );
  INV_X1 U8283 ( .A(n10929), .ZN(n6632) );
  AND2_X1 U8284 ( .A1(n8704), .A2(n8278), .ZN(n12560) );
  NOR2_X1 U8285 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10867), .ZN(n10429) );
  OR2_X1 U8286 ( .A1(n10478), .A2(n10477), .ZN(n10480) );
  NAND2_X1 U8287 ( .A1(n6602), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n10475) );
  NAND2_X1 U8288 ( .A1(n6474), .A2(n15206), .ZN(n6623) );
  NOR2_X1 U8289 ( .A1(n14991), .A2(n7209), .ZN(n11090) );
  NOR2_X1 U8290 ( .A1(n15007), .A2(n11118), .ZN(n7209) );
  INV_X1 U8291 ( .A(n6752), .ZN(n15052) );
  NOR2_X1 U8292 ( .A1(n15043), .A2(n11131), .ZN(n7212) );
  INV_X1 U8293 ( .A(n12469), .ZN(n12480) );
  NAND2_X1 U8294 ( .A1(n12470), .A2(n12471), .ZN(n12473) );
  INV_X1 U8295 ( .A(n6673), .ZN(n12527) );
  AOI22_X1 U8296 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n14470), .B1(n12546), 
        .B2(n12534), .ZN(n14481) );
  INV_X1 U8297 ( .A(n12565), .ZN(n12574) );
  NOR2_X1 U8298 ( .A1(n12565), .A2(n6746), .ZN(n7409) );
  INV_X1 U8299 ( .A(n12255), .ZN(n6746) );
  NAND2_X1 U8300 ( .A1(n12582), .A2(n6672), .ZN(n6671) );
  NAND2_X1 U8301 ( .A1(n12583), .A2(n12587), .ZN(n6672) );
  NAND2_X1 U8302 ( .A1(n12254), .A2(n12253), .ZN(n12583) );
  NOR2_X1 U8303 ( .A1(n12585), .A2(n15185), .ZN(n6669) );
  AND2_X1 U8304 ( .A1(n8806), .A2(n8807), .ZN(n12600) );
  OR2_X1 U8305 ( .A1(n8628), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8637) );
  AND2_X1 U8306 ( .A1(n12641), .A2(n12640), .ZN(n12658) );
  INV_X1 U8307 ( .A(n12674), .ZN(n12246) );
  AND4_X1 U8308 ( .A1(n8612), .A2(n8611), .A3(n8610), .A4(n8609), .ZN(n12685)
         );
  INV_X1 U8309 ( .A(n7084), .ZN(n7083) );
  AOI21_X1 U8310 ( .B1(n7084), .B2(n12729), .A(n7082), .ZN(n7081) );
  INV_X1 U8311 ( .A(n8780), .ZN(n7082) );
  OR2_X1 U8312 ( .A1(n8527), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U8313 ( .A1(n12236), .A2(n12235), .ZN(n12738) );
  NOR2_X1 U8314 ( .A1(n7487), .A2(n6528), .ZN(n7380) );
  OR2_X1 U8315 ( .A1(n14424), .A2(n12781), .ZN(n12755) );
  NAND2_X1 U8316 ( .A1(n12234), .A2(n12233), .ZN(n12780) );
  OR3_X1 U8317 ( .A1(n8435), .A2(P3_REG3_REG_10__SCAN_IN), .A3(
        P3_REG3_REG_11__SCAN_IN), .ZN(n8453) );
  AND4_X1 U8318 ( .A1(n8426), .A2(n8425), .A3(n8424), .A4(n8423), .ZN(n14495)
         );
  AOI21_X1 U8319 ( .B1(n7386), .B2(n7388), .A(n7384), .ZN(n7383) );
  INV_X1 U8320 ( .A(n7386), .ZN(n7385) );
  INV_X1 U8321 ( .A(n7390), .ZN(n7388) );
  INV_X1 U8322 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8403) );
  AND2_X1 U8323 ( .A1(n8389), .A2(n11564), .ZN(n8404) );
  CLKBUF_X1 U8324 ( .A(n15108), .Z(n15109) );
  INV_X1 U8325 ( .A(n8740), .ZN(n7069) );
  INV_X1 U8326 ( .A(n15125), .ZN(n15121) );
  NAND2_X1 U8327 ( .A1(n8342), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8316) );
  NAND3_X1 U8328 ( .A1(n9657), .A2(n9650), .A3(n6722), .ZN(n15187) );
  NAND2_X1 U8329 ( .A1(n8586), .A2(n8824), .ZN(n12690) );
  INV_X1 U8330 ( .A(n15219), .ZN(n15242) );
  INV_X1 U8331 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8233) );
  AND2_X1 U8332 ( .A1(n8227), .A2(n6574), .ZN(n8239) );
  AND2_X1 U8333 ( .A1(n8231), .A2(n7407), .ZN(n7406) );
  NOR2_X1 U8334 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n8230) );
  XNOR2_X1 U8335 ( .A(n8850), .B(n8849), .ZN(n9649) );
  OAI21_X1 U8336 ( .B1(n8848), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8850) );
  NAND2_X1 U8337 ( .A1(n8589), .A2(n8197), .ZN(n8599) );
  NAND2_X1 U8338 ( .A1(n7006), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8197) );
  AND2_X1 U8339 ( .A1(n8199), .A2(n8198), .ZN(n8598) );
  AND2_X1 U8340 ( .A1(n8194), .A2(n8193), .ZN(n8554) );
  AND2_X1 U8341 ( .A1(n8192), .A2(n8191), .ZN(n8534) );
  AOI21_X1 U8342 ( .B1(n7022), .B2(n7024), .A(n7021), .ZN(n7020) );
  INV_X1 U8343 ( .A(n8186), .ZN(n7021) );
  NAND2_X1 U8344 ( .A1(n7013), .A2(n7014), .ZN(n8464) );
  AOI21_X1 U8345 ( .B1(n7016), .B2(n7018), .A(n7015), .ZN(n7014) );
  INV_X1 U8346 ( .A(n8173), .ZN(n7015) );
  INV_X1 U8347 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8447) );
  CLKBUF_X1 U8348 ( .A(n8354), .Z(n8355) );
  NAND2_X1 U8349 ( .A1(n8305), .A2(n8304), .ZN(n8303) );
  XNOR2_X1 U8350 ( .A(n8289), .B(P3_IR_REG_1__SCAN_IN), .ZN(n10486) );
  NAND2_X1 U8351 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8289) );
  NOR2_X1 U8352 ( .A1(n7182), .A2(n7179), .ZN(n7174) );
  INV_X1 U8353 ( .A(n7181), .ZN(n7180) );
  OAI22_X1 U8354 ( .A1(n13038), .A2(n6552), .B1(n13036), .B2(n13037), .ZN(
        n7181) );
  INV_X1 U8355 ( .A(n13140), .ZN(n7184) );
  INV_X1 U8356 ( .A(n13042), .ZN(n7179) );
  INV_X1 U8357 ( .A(n6619), .ZN(n11528) );
  OR2_X1 U8358 ( .A1(n7163), .A2(n6593), .ZN(n7160) );
  OR2_X1 U8359 ( .A1(n9184), .A2(n9183), .ZN(n9199) );
  OR2_X1 U8360 ( .A1(n9059), .A2(n9058), .ZN(n9081) );
  OR2_X1 U8361 ( .A1(n11701), .A2(n11702), .ZN(n7172) );
  OR2_X1 U8362 ( .A1(n9147), .A2(n11706), .ZN(n9184) );
  OR2_X1 U8363 ( .A1(n9305), .A2(n13124), .ZN(n9322) );
  INV_X1 U8364 ( .A(n7164), .ZN(n7163) );
  CLKBUF_X1 U8365 ( .A(n12974), .Z(n11736) );
  NAND2_X1 U8366 ( .A1(n7464), .A2(n7463), .ZN(n7462) );
  INV_X1 U8367 ( .A(n9408), .ZN(n7463) );
  INV_X1 U8368 ( .A(n9409), .ZN(n7464) );
  AND2_X1 U8369 ( .A1(n6989), .A2(n9407), .ZN(n6658) );
  OAI21_X1 U8370 ( .B1(n6538), .B2(n9454), .A(n6991), .ZN(n6987) );
  INV_X1 U8371 ( .A(n9005), .ZN(n9446) );
  AOI21_X1 U8372 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n9985), .A(n9980), .ZN(
        n10068) );
  AOI21_X1 U8373 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n10050), .A(n10049), .ZN(
        n10053) );
  AOI21_X1 U8374 ( .B1(n10083), .B2(P2_REG1_REG_11__SCAN_IN), .A(n10079), .ZN(
        n10082) );
  AOI21_X1 U8375 ( .B1(n13188), .B2(P2_REG1_REG_17__SCAN_IN), .A(n13187), .ZN(
        n13198) );
  AND2_X1 U8376 ( .A1(n12207), .A2(n9471), .ZN(n13232) );
  INV_X1 U8377 ( .A(n13248), .ZN(n6687) );
  NAND2_X1 U8378 ( .A1(n13267), .A2(n13266), .ZN(n13265) );
  NAND2_X1 U8379 ( .A1(n13297), .A2(n13551), .ZN(n13285) );
  AND2_X1 U8380 ( .A1(n9392), .A2(n9370), .ZN(n13272) );
  NOR2_X2 U8381 ( .A1(n13315), .A2(n13470), .ZN(n13297) );
  OR2_X1 U8382 ( .A1(n9266), .A2(n13117), .ZN(n9282) );
  AOI21_X1 U8383 ( .B1(n6484), .B2(n7243), .A(n6542), .ZN(n7239) );
  INV_X1 U8384 ( .A(n7255), .ZN(n6852) );
  AOI21_X1 U8385 ( .B1(n7255), .B2(n6851), .A(n6526), .ZN(n6850) );
  AOI21_X1 U8386 ( .B1(n6486), .B2(n7256), .A(n6545), .ZN(n7255) );
  NAND2_X1 U8387 ( .A1(n11544), .A2(n6663), .ZN(n11663) );
  OAI21_X1 U8388 ( .B1(n11243), .B2(n7276), .A(n7274), .ZN(n11452) );
  INV_X1 U8389 ( .A(n7275), .ZN(n7274) );
  NAND2_X1 U8390 ( .A1(n7281), .A2(n11459), .ZN(n11541) );
  NOR2_X1 U8391 ( .A1(n6821), .A2(n11458), .ZN(n6820) );
  INV_X1 U8392 ( .A(n10723), .ZN(n14525) );
  OR2_X1 U8393 ( .A1(n9095), .A2(n11301), .ZN(n9132) );
  INV_X1 U8394 ( .A(n10718), .ZN(n6807) );
  AND2_X1 U8395 ( .A1(n10724), .A2(n11340), .ZN(n10962) );
  NAND2_X1 U8396 ( .A1(n6860), .A2(n6862), .ZN(n10715) );
  AOI21_X1 U8397 ( .B1(n7273), .B2(n6861), .A(n6510), .ZN(n6862) );
  NOR2_X1 U8398 ( .A1(n12173), .A2(n6815), .ZN(n6814) );
  INV_X1 U8399 ( .A(n12207), .ZN(n6815) );
  OR2_X1 U8400 ( .A1(n13242), .A2(n13241), .ZN(n13442) );
  OAI21_X1 U8401 ( .B1(n13399), .B2(n6504), .A(n12151), .ZN(n13388) );
  NAND2_X1 U8402 ( .A1(n9197), .A2(n9196), .ZN(n13520) );
  NAND2_X1 U8403 ( .A1(n10202), .A2(n10201), .ZN(n11337) );
  NOR2_X1 U8404 ( .A1(n9194), .A2(n6857), .ZN(n6853) );
  NAND2_X1 U8405 ( .A1(n8879), .A2(n6858), .ZN(n6857) );
  NAND2_X1 U8406 ( .A1(n9466), .A2(n9465), .ZN(n9492) );
  OR2_X1 U8407 ( .A1(n9142), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n9164) );
  OR2_X1 U8408 ( .A1(n9070), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n9072) );
  OR2_X1 U8409 ( .A1(n9053), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n9070) );
  NAND2_X1 U8410 ( .A1(n7417), .A2(n7527), .ZN(n8897) );
  OR2_X1 U8411 ( .A1(n7782), .A2(n7781), .ZN(n7796) );
  NAND2_X1 U8412 ( .A1(n6927), .A2(n6925), .ZN(n13632) );
  NAND2_X1 U8413 ( .A1(n13689), .A2(n13688), .ZN(n6927) );
  NOR2_X1 U8414 ( .A1(n7943), .A2(n13671), .ZN(n7957) );
  NAND2_X1 U8415 ( .A1(n12096), .A2(n13676), .ZN(n13679) );
  OR2_X1 U8416 ( .A1(n7987), .A2(n13691), .ZN(n8005) );
  AOI21_X1 U8417 ( .B1(n6935), .B2(n6937), .A(n6534), .ZN(n6934) );
  INV_X1 U8418 ( .A(n11651), .ZN(n6935) );
  NOR2_X1 U8419 ( .A1(n8005), .A2(n8004), .ZN(n8016) );
  NAND2_X1 U8420 ( .A1(n11650), .A2(n11651), .ZN(n11684) );
  NAND2_X1 U8421 ( .A1(n7319), .A2(n7318), .ZN(n7317) );
  NOR2_X1 U8422 ( .A1(n7325), .A2(n7326), .ZN(n7321) );
  AND2_X1 U8423 ( .A1(n6929), .A2(n7335), .ZN(n6928) );
  AOI21_X1 U8424 ( .B1(n7339), .B2(n7337), .A(n7336), .ZN(n7335) );
  AND2_X1 U8425 ( .A1(n6901), .A2(n6900), .ZN(n6899) );
  NAND2_X1 U8426 ( .A1(n6903), .A2(n11932), .ZN(n6900) );
  AND4_X1 U8427 ( .A1(n7920), .A2(n7919), .A3(n7918), .A4(n7917), .ZN(n12024)
         );
  AND4_X1 U8428 ( .A1(n7899), .A2(n7898), .A3(n7897), .A4(n7896), .ZN(n12016)
         );
  AND4_X1 U8429 ( .A1(n7880), .A2(n7879), .A3(n7878), .A4(n7877), .ZN(n11840)
         );
  AND4_X1 U8430 ( .A1(n7859), .A2(n7858), .A3(n7857), .A4(n7856), .ZN(n11841)
         );
  NAND2_X1 U8431 ( .A1(n13923), .A2(n13922), .ZN(n13921) );
  OAI21_X1 U8432 ( .B1(n13923), .B2(n13922), .A(n13921), .ZN(n14113) );
  NAND2_X1 U8433 ( .A1(n6741), .A2(n7117), .ZN(n13952) );
  AND2_X1 U8434 ( .A1(n7118), .A2(n6579), .ZN(n7117) );
  NAND2_X1 U8435 ( .A1(n7119), .A2(n6742), .ZN(n6741) );
  NAND2_X1 U8436 ( .A1(n13952), .A2(n13953), .ZN(n13951) );
  INV_X1 U8437 ( .A(n13980), .ZN(n7352) );
  OAI21_X1 U8438 ( .B1(n14006), .B2(n14009), .A(n8023), .ZN(n13994) );
  NAND2_X1 U8439 ( .A1(n13994), .A2(n13995), .ZN(n13993) );
  NAND2_X1 U8440 ( .A1(n7123), .A2(n7121), .ZN(n14022) );
  AOI21_X1 U8441 ( .B1(n7124), .B2(n14053), .A(n7122), .ZN(n7121) );
  INV_X1 U8442 ( .A(n7996), .ZN(n7122) );
  NAND2_X1 U8443 ( .A1(n7360), .A2(n7358), .ZN(n14052) );
  AOI21_X1 U8444 ( .B1(n7361), .B2(n11870), .A(n7359), .ZN(n7358) );
  NOR2_X1 U8445 ( .A1(n11874), .A2(n7362), .ZN(n7361) );
  NAND2_X1 U8446 ( .A1(n7137), .A2(n7136), .ZN(n14066) );
  AOI21_X1 U8447 ( .B1(n7138), .B2(n11610), .A(n6548), .ZN(n7136) );
  NAND2_X1 U8448 ( .A1(n11574), .A2(n11858), .ZN(n11468) );
  NOR2_X1 U8449 ( .A1(n7873), .A2(n7872), .ZN(n7892) );
  INV_X1 U8450 ( .A(n7831), .ZN(n7113) );
  INV_X1 U8451 ( .A(n7115), .ZN(n7114) );
  NAND2_X1 U8452 ( .A1(n8094), .A2(n8093), .ZN(n14390) );
  NAND2_X1 U8453 ( .A1(n7347), .A2(n7346), .ZN(n10994) );
  AOI21_X1 U8454 ( .B1(n7349), .B2(n7351), .A(n6541), .ZN(n7346) );
  OR2_X1 U8455 ( .A1(n7796), .A2(n7795), .ZN(n7813) );
  NOR2_X1 U8456 ( .A1(n7813), .A2(n9790), .ZN(n7839) );
  INV_X1 U8457 ( .A(n7129), .ZN(n7128) );
  OAI21_X1 U8458 ( .B1(n11960), .B2(n7130), .A(n7802), .ZN(n7129) );
  NAND2_X1 U8459 ( .A1(n7133), .A2(n11960), .ZN(n10579) );
  NOR2_X2 U8460 ( .A1(n14654), .A2(n14725), .ZN(n11008) );
  NAND2_X1 U8461 ( .A1(n6700), .A2(n6699), .ZN(n14653) );
  NAND2_X1 U8462 ( .A1(n8085), .A2(n8084), .ZN(n14642) );
  INV_X1 U8463 ( .A(n11959), .ZN(n14643) );
  NAND2_X1 U8464 ( .A1(n11774), .A2(n7693), .ZN(n10116) );
  INV_X1 U8465 ( .A(n11773), .ZN(n7692) );
  NAND2_X1 U8466 ( .A1(n7680), .A2(n7679), .ZN(n11773) );
  INV_X1 U8467 ( .A(n7108), .ZN(n14042) );
  OR2_X1 U8468 ( .A1(n11754), .A2(n8069), .ZN(n14721) );
  OR2_X1 U8469 ( .A1(n10527), .A2(n14058), .ZN(n14700) );
  NAND2_X1 U8470 ( .A1(n8068), .A2(n11928), .ZN(n14664) );
  NAND2_X1 U8471 ( .A1(n8044), .A2(n8043), .ZN(n7425) );
  XNOR2_X1 U8472 ( .A(n8044), .B(n8043), .ZN(n13583) );
  AND2_X1 U8473 ( .A1(n7633), .A2(n7632), .ZN(n13591) );
  NAND2_X1 U8474 ( .A1(n7453), .A2(n7450), .ZN(n7631) );
  AND2_X1 U8475 ( .A1(n7648), .A2(n7647), .ZN(n13598) );
  NAND2_X1 U8476 ( .A1(n7604), .A2(n6743), .ZN(n7648) );
  INV_X1 U8477 ( .A(n6897), .ZN(n6743) );
  XNOR2_X1 U8478 ( .A(n8142), .B(P1_IR_REG_23__SCAN_IN), .ZN(n9756) );
  AND2_X1 U8479 ( .A1(n7434), .A2(n7597), .ZN(n9297) );
  NOR2_X1 U8480 ( .A1(n7343), .A2(n7345), .ZN(n7342) );
  NAND2_X1 U8481 ( .A1(n7344), .A2(n8066), .ZN(n7343) );
  OR2_X1 U8482 ( .A1(n8062), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n8141) );
  NAND2_X1 U8483 ( .A1(n8064), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8065) );
  AND2_X1 U8484 ( .A1(n7984), .A2(n7983), .ZN(n11214) );
  OR2_X1 U8485 ( .A1(n7437), .A2(n7436), .ZN(n7984) );
  NAND2_X1 U8486 ( .A1(n7593), .A2(n7591), .ZN(n7982) );
  NAND2_X1 U8487 ( .A1(n6893), .A2(n7439), .ZN(n7966) );
  AND2_X1 U8488 ( .A1(n7888), .A2(n7868), .ZN(n10169) );
  NAND2_X1 U8489 ( .A1(n7538), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7416) );
  NAND2_X1 U8490 ( .A1(n7687), .A2(n7686), .ZN(n7695) );
  INV_X1 U8491 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n7806) );
  INV_X1 U8492 ( .A(n14304), .ZN(n14303) );
  XNOR2_X1 U8493 ( .A(n14270), .B(n7232), .ZN(n14311) );
  OAI21_X1 U8494 ( .B1(n15275), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6531), .ZN(
        n6759) );
  NOR2_X1 U8495 ( .A1(n14275), .A2(n14274), .ZN(n14319) );
  AND2_X1 U8496 ( .A1(n7236), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n14275) );
  INV_X1 U8497 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14324) );
  NAND2_X1 U8498 ( .A1(n6763), .A2(n14325), .ZN(n14326) );
  NAND2_X1 U8499 ( .A1(n15280), .A2(n15279), .ZN(n6763) );
  OAI21_X1 U8500 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n15075), .A(n14281), .ZN(
        n14295) );
  INV_X1 U8501 ( .A(n14353), .ZN(n6770) );
  OR2_X1 U8502 ( .A1(n14348), .A2(n7227), .ZN(n6768) );
  AND2_X1 U8503 ( .A1(n14348), .A2(n7227), .ZN(n6771) );
  NAND2_X1 U8504 ( .A1(n7303), .A2(n10836), .ZN(n7314) );
  XNOR2_X1 U8505 ( .A(n7303), .B(n10836), .ZN(n10764) );
  INV_X1 U8506 ( .A(n7037), .ZN(n14419) );
  AOI21_X1 U8507 ( .B1(n12392), .B2(n12390), .A(n7041), .ZN(n7037) );
  NAND2_X1 U8508 ( .A1(n12329), .A2(n6483), .ZN(n7056) );
  OAI21_X1 U8509 ( .B1(n7063), .B2(n6483), .A(n7055), .ZN(n7054) );
  INV_X1 U8510 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n11564) );
  NAND2_X1 U8511 ( .A1(n12383), .A2(n12293), .ZN(n12339) );
  NAND2_X1 U8512 ( .A1(n8604), .A2(n8603), .ZN(n12677) );
  AND4_X1 U8513 ( .A1(n8485), .A2(n8484), .A3(n8483), .A4(n8482), .ZN(n12798)
         );
  NAND2_X1 U8514 ( .A1(n8647), .A2(n8646), .ZN(n12829) );
  AND2_X1 U8515 ( .A1(n10954), .A2(n9533), .ZN(n11216) );
  NOR2_X1 U8516 ( .A1(n12375), .A2(n7032), .ZN(n7031) );
  INV_X1 U8517 ( .A(n9547), .ZN(n7032) );
  NAND2_X1 U8518 ( .A1(n11561), .A2(n9547), .ZN(n12376) );
  NAND2_X1 U8519 ( .A1(n12271), .A2(n12270), .ZN(n12392) );
  NAND2_X1 U8520 ( .A1(n8617), .A2(n8616), .ZN(n12664) );
  AND4_X1 U8521 ( .A1(n8460), .A2(n8459), .A3(n8458), .A4(n8457), .ZN(n14496)
         );
  AND2_X1 U8522 ( .A1(n9585), .A2(n9584), .ZN(n14971) );
  AND2_X1 U8523 ( .A1(n6518), .A2(n12282), .ZN(n7048) );
  AND2_X1 U8524 ( .A1(n8681), .A2(n8680), .ZN(n12598) );
  INV_X1 U8525 ( .A(n7065), .ZN(n7052) );
  AND2_X1 U8526 ( .A1(n12947), .A2(n9607), .ZN(n10866) );
  INV_X1 U8527 ( .A(n12597), .ZN(n12447) );
  INV_X1 U8528 ( .A(n12704), .ZN(n12452) );
  INV_X1 U8529 ( .A(n12715), .ZN(n12739) );
  INV_X1 U8530 ( .A(n14496), .ZN(n12455) );
  OR2_X1 U8531 ( .A1(n6471), .A2(n10867), .ZN(n8282) );
  INV_X1 U8532 ( .A(n7216), .ZN(n10437) );
  INV_X1 U8533 ( .A(n6621), .ZN(n14973) );
  INV_X1 U8534 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15010) );
  INV_X1 U8535 ( .A(n7211), .ZN(n14993) );
  INV_X1 U8536 ( .A(n6751), .ZN(n15011) );
  INV_X1 U8537 ( .A(n7214), .ZN(n15039) );
  INV_X1 U8538 ( .A(n6622), .ZN(n11416) );
  XNOR2_X1 U8539 ( .A(n12464), .B(n12480), .ZN(n11585) );
  NOR2_X1 U8540 ( .A1(n11585), .A2(n8480), .ZN(n12465) );
  INV_X1 U8541 ( .A(n6755), .ZN(n14451) );
  INV_X1 U8542 ( .A(n6675), .ZN(n14450) );
  NAND2_X1 U8543 ( .A1(n8227), .A2(n8226), .ZN(n8538) );
  NAND2_X1 U8544 ( .A1(n6670), .A2(n6667), .ZN(n12821) );
  NOR2_X1 U8545 ( .A1(n6669), .A2(n6668), .ZN(n6667) );
  NAND2_X1 U8546 ( .A1(n6671), .A2(n15183), .ZN(n6670) );
  NOR2_X1 U8547 ( .A1(n12584), .A2(n15187), .ZN(n6668) );
  AND2_X1 U8548 ( .A1(n12612), .A2(n12611), .ZN(n12832) );
  NAND2_X1 U8549 ( .A1(n7402), .A2(n7399), .ZN(n12647) );
  NAND2_X1 U8550 ( .A1(n8627), .A2(n8626), .ZN(n12654) );
  NAND2_X1 U8551 ( .A1(n12855), .A2(n8786), .ZN(n12670) );
  AND2_X1 U8552 ( .A1(n12710), .A2(n12242), .ZN(n12701) );
  NAND2_X1 U8553 ( .A1(n12731), .A2(n8781), .ZN(n12717) );
  AND2_X1 U8554 ( .A1(n7381), .A2(n7382), .ZN(n12750) );
  NAND2_X1 U8555 ( .A1(n7093), .A2(n8765), .ZN(n12774) );
  NAND2_X1 U8556 ( .A1(n7392), .A2(n7389), .ZN(n15093) );
  INV_X1 U8557 ( .A(n12695), .ZN(n15100) );
  NAND2_X1 U8558 ( .A1(n7070), .A2(n8737), .ZN(n15136) );
  NAND2_X1 U8559 ( .A1(n15153), .A2(n12217), .ZN(n7070) );
  INV_X1 U8560 ( .A(n15104), .ZN(n15203) );
  INV_X1 U8561 ( .A(n8706), .ZN(n12890) );
  INV_X1 U8562 ( .A(n12589), .ZN(n12901) );
  INV_X1 U8563 ( .A(n12602), .ZN(n12905) );
  NAND2_X1 U8564 ( .A1(n8578), .A2(n8577), .ZN(n12931) );
  NAND2_X1 U8565 ( .A1(n6717), .A2(n6716), .ZN(n9514) );
  INV_X1 U8566 ( .A(n9766), .ZN(n6717) );
  AND2_X1 U8567 ( .A1(n9649), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12947) );
  INV_X1 U8568 ( .A(n8263), .ZN(n12958) );
  OR2_X1 U8569 ( .A1(n8694), .A2(n8693), .ZN(n8696) );
  XNOR2_X1 U8570 ( .A(n8683), .B(n8682), .ZN(n12961) );
  INV_X1 U8571 ( .A(n9659), .ZN(n9654) );
  NAND2_X1 U8572 ( .A1(n8857), .A2(n6497), .ZN(n11368) );
  NAND2_X1 U8573 ( .A1(n8848), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8718) );
  NAND2_X1 U8574 ( .A1(n7043), .A2(n7042), .ZN(n8713) );
  NAND2_X1 U8575 ( .A1(n8711), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7042) );
  OAI21_X1 U8576 ( .B1(n8712), .B2(n6724), .A(P3_IR_REG_21__SCAN_IN), .ZN(
        n7043) );
  XNOR2_X1 U8577 ( .A(n8717), .B(n8716), .ZN(n10563) );
  NAND2_X1 U8578 ( .A1(n7008), .A2(n7007), .ZN(n8587) );
  INV_X1 U8579 ( .A(SI_17_), .ZN(n10059) );
  INV_X1 U8580 ( .A(n14456), .ZN(n12543) );
  INV_X1 U8581 ( .A(SI_16_), .ZN(n10023) );
  INV_X1 U8582 ( .A(SI_15_), .ZN(n9961) );
  NAND2_X1 U8583 ( .A1(n8490), .A2(n8183), .ZN(n8507) );
  INV_X1 U8584 ( .A(SI_14_), .ZN(n9772) );
  XNOR2_X1 U8585 ( .A(n8494), .B(n8493), .ZN(n12494) );
  INV_X1 U8586 ( .A(SI_13_), .ZN(n9745) );
  INV_X1 U8587 ( .A(SI_12_), .ZN(n9728) );
  INV_X1 U8588 ( .A(SI_11_), .ZN(n9719) );
  NAND2_X1 U8589 ( .A1(n8431), .A2(n8171), .ZN(n8445) );
  NAND2_X1 U8590 ( .A1(n8153), .A2(n8321), .ZN(n8333) );
  NAND2_X1 U8591 ( .A1(n11298), .A2(n11297), .ZN(n11372) );
  NAND2_X1 U8592 ( .A1(n9279), .A2(n9278), .ZN(n13488) );
  NAND2_X1 U8593 ( .A1(n7146), .A2(n7151), .ZN(n13094) );
  AND2_X1 U8594 ( .A1(n10573), .A2(n7192), .ZN(n7187) );
  OAI21_X1 U8595 ( .B1(n6684), .B2(n7163), .A(n7161), .ZN(n11526) );
  INV_X1 U8596 ( .A(n7189), .ZN(n10410) );
  AND2_X1 U8597 ( .A1(n10207), .A2(n14865), .ZN(n13137) );
  NOR2_X1 U8598 ( .A1(n7155), .A2(n7148), .ZN(n7147) );
  INV_X1 U8599 ( .A(n7149), .ZN(n7148) );
  AND2_X1 U8600 ( .A1(n10215), .A2(n10204), .ZN(n13129) );
  AND2_X1 U8601 ( .A1(n10215), .A2(n10214), .ZN(n13097) );
  NAND2_X1 U8602 ( .A1(n13004), .A2(n6660), .ZN(n6659) );
  NAND2_X1 U8603 ( .A1(n13061), .A2(n13060), .ZN(n6661) );
  INV_X1 U8604 ( .A(n13005), .ZN(n6660) );
  AND2_X1 U8605 ( .A1(n6650), .A2(n11672), .ZN(n6649) );
  OR2_X1 U8606 ( .A1(n10179), .A2(n9503), .ZN(n6650) );
  AOI21_X1 U8607 ( .B1(n10648), .B2(P2_REG1_REG_13__SCAN_IN), .A(n10647), .ZN(
        n10651) );
  NOR2_X1 U8608 ( .A1(n11281), .A2(n11280), .ZN(n11283) );
  OAI21_X1 U8609 ( .B1(n13284), .B2(n7251), .A(n7250), .ZN(n13261) );
  NAND2_X1 U8610 ( .A1(n13282), .A2(n12204), .ZN(n13264) );
  NAND2_X1 U8611 ( .A1(n7258), .A2(n7259), .ZN(n13296) );
  NAND2_X1 U8612 ( .A1(n13323), .A2(n12198), .ZN(n13308) );
  NAND2_X1 U8613 ( .A1(n6837), .A2(n12194), .ZN(n13348) );
  OR2_X1 U8614 ( .A1(n13358), .A2(n12193), .ZN(n6837) );
  NAND2_X1 U8615 ( .A1(n13354), .A2(n12155), .ZN(n13337) );
  NAND2_X1 U8616 ( .A1(n13372), .A2(n12154), .ZN(n13352) );
  NAND2_X1 U8617 ( .A1(n6866), .A2(n6871), .ZN(n13370) );
  NAND2_X1 U8618 ( .A1(n7240), .A2(n12188), .ZN(n13385) );
  OAI21_X1 U8619 ( .B1(n13403), .B2(n7243), .A(n6484), .ZN(n13384) );
  OAI21_X1 U8620 ( .B1(n11659), .B2(n6486), .A(n7256), .ZN(n12146) );
  NAND2_X1 U8621 ( .A1(n6822), .A2(n6823), .ZN(n14524) );
  NAND2_X1 U8622 ( .A1(n11243), .A2(n11242), .ZN(n11245) );
  NAND2_X1 U8623 ( .A1(n11253), .A2(n11252), .ZN(n11456) );
  NAND2_X1 U8624 ( .A1(n10967), .A2(n10966), .ZN(n10969) );
  NAND2_X1 U8625 ( .A1(n6841), .A2(n6842), .ZN(n10675) );
  NAND2_X1 U8626 ( .A1(n10798), .A2(n6843), .ZN(n6841) );
  NAND2_X1 U8627 ( .A1(n6845), .A2(n10673), .ZN(n10811) );
  OR2_X1 U8628 ( .A1(n10798), .A2(n10672), .ZN(n6845) );
  NAND2_X1 U8629 ( .A1(n6864), .A2(n6863), .ZN(n10812) );
  OAI21_X1 U8630 ( .B1(n7245), .B2(n6828), .A(n10669), .ZN(n14848) );
  NOR2_X1 U8631 ( .A1(n10892), .A2(n7246), .ZN(n6828) );
  NAND2_X1 U8632 ( .A1(n9437), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6859) );
  INV_X1 U8633 ( .A(n13420), .ZN(n14846) );
  INV_X1 U8634 ( .A(n13425), .ZN(n14855) );
  NAND2_X1 U8635 ( .A1(n9244), .A2(n9859), .ZN(n7264) );
  NAND2_X1 U8636 ( .A1(n9437), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7265) );
  NAND2_X1 U8637 ( .A1(n7206), .A2(n7205), .ZN(n7204) );
  NAND2_X1 U8638 ( .A1(n14871), .A2(n10780), .ZN(n13420) );
  NAND2_X1 U8639 ( .A1(n14886), .A2(n10208), .ZN(n14865) );
  NAND2_X1 U8640 ( .A1(n9146), .A2(n9145), .ZN(n11696) );
  OAI22_X1 U8641 ( .A1(n10064), .A2(n9832), .B1(n9741), .B2(n7199), .ZN(n9076)
         );
  AND2_X1 U8642 ( .A1(n9439), .A2(n9438), .ZN(n13536) );
  INV_X1 U8643 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6818) );
  INV_X1 U8644 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6641) );
  INV_X1 U8645 ( .A(n13288), .ZN(n13551) );
  NAND2_X1 U8646 ( .A1(n9111), .A2(n9110), .ZN(n11457) );
  INV_X1 U8647 ( .A(n14882), .ZN(n14879) );
  INV_X1 U8648 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8881) );
  NAND2_X1 U8649 ( .A1(n9498), .A2(n8901), .ZN(n13593) );
  NAND2_X1 U8650 ( .A1(n9496), .A2(n6592), .ZN(n13595) );
  XNOR2_X1 U8651 ( .A(n9493), .B(P2_IR_REG_24__SCAN_IN), .ZN(n13597) );
  NAND2_X1 U8652 ( .A1(n9492), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9493) );
  AND2_X1 U8653 ( .A1(n8912), .A2(n8906), .ZN(n8909) );
  INV_X1 U8654 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10508) );
  INV_X1 U8655 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10127) );
  INV_X1 U8656 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9916) );
  INV_X1 U8657 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9741) );
  INV_X1 U8658 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9732) );
  INV_X1 U8659 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9726) );
  INV_X1 U8660 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9702) );
  INV_X1 U8661 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9683) );
  INV_X1 U8662 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9677) );
  NOR2_X2 U8663 ( .A1(n8947), .A2(n8959), .ZN(n14787) );
  NAND2_X1 U8664 ( .A1(n6921), .A2(n7323), .ZN(n11352) );
  NAND2_X1 U8665 ( .A1(n13720), .A2(n12117), .ZN(n6909) );
  NAND2_X1 U8666 ( .A1(n7330), .A2(n13697), .ZN(n13699) );
  NAND2_X1 U8667 ( .A1(n13632), .A2(n13696), .ZN(n7330) );
  NAND2_X1 U8668 ( .A1(n11481), .A2(n6519), .ZN(n11649) );
  NOR2_X1 U8669 ( .A1(n7308), .A2(n12137), .ZN(n7307) );
  INV_X1 U8670 ( .A(n7312), .ZN(n7308) );
  OAI21_X1 U8671 ( .B1(n12137), .B2(n7312), .A(n7310), .ZN(n7309) );
  OAI21_X1 U8672 ( .B1(n12137), .B2(n13604), .A(n7312), .ZN(n7310) );
  NAND2_X1 U8673 ( .A1(n13604), .A2(n12137), .ZN(n7311) );
  NAND2_X1 U8674 ( .A1(n6913), .A2(n6916), .ZN(n11353) );
  NAND2_X1 U8675 ( .A1(n6921), .A2(n6918), .ZN(n6913) );
  NAND2_X1 U8676 ( .A1(n6927), .A2(n12064), .ZN(n13634) );
  AND2_X2 U8677 ( .A1(n7851), .A2(n7850), .ZN(n14407) );
  NAND2_X1 U8678 ( .A1(n11684), .A2(n6937), .ZN(n11716) );
  INV_X1 U8679 ( .A(n9616), .ZN(n9618) );
  AOI21_X1 U8680 ( .B1(n10837), .B2(n7320), .A(n7317), .ZN(n11268) );
  INV_X1 U8681 ( .A(n7321), .ZN(n7320) );
  XNOR2_X1 U8682 ( .A(n12027), .B(n12025), .ZN(n13732) );
  NAND2_X1 U8683 ( .A1(n9638), .A2(n9627), .ZN(n13740) );
  OR2_X1 U8684 ( .A1(n7932), .A2(n7931), .ZN(n13757) );
  OR2_X1 U8685 ( .A1(n7707), .A2(n7681), .ZN(n7682) );
  INV_X1 U8686 ( .A(n8070), .ZN(n13916) );
  INV_X1 U8687 ( .A(n7371), .ZN(n7368) );
  NOR2_X1 U8688 ( .A1(n7375), .A2(n7374), .ZN(n13946) );
  INV_X1 U8689 ( .A(n8109), .ZN(n7374) );
  INV_X1 U8690 ( .A(n13960), .ZN(n7375) );
  NAND2_X1 U8691 ( .A1(n13978), .A2(n8025), .ZN(n13967) );
  NAND2_X1 U8692 ( .A1(n14036), .A2(n8104), .ZN(n14020) );
  NAND2_X1 U8693 ( .A1(n7126), .A2(n7124), .ZN(n14034) );
  AND2_X1 U8694 ( .A1(n7126), .A2(n11879), .ZN(n14035) );
  OR2_X1 U8695 ( .A1(n14054), .A2(n14053), .ZN(n7126) );
  NAND2_X1 U8696 ( .A1(n7363), .A2(n6553), .ZN(n14075) );
  OR2_X1 U8697 ( .A1(n14081), .A2(n11870), .ZN(n7363) );
  NAND2_X1 U8698 ( .A1(n7140), .A2(n7138), .ZN(n14093) );
  NAND2_X1 U8699 ( .A1(n7140), .A2(n7934), .ZN(n14092) );
  NAND2_X1 U8700 ( .A1(n7926), .A2(n7925), .ZN(n14571) );
  NAND2_X1 U8701 ( .A1(n7912), .A2(n7911), .ZN(n13738) );
  NAND2_X1 U8702 ( .A1(n11571), .A2(n7366), .ZN(n11469) );
  INV_X1 U8703 ( .A(n11839), .ZN(n14585) );
  NAND2_X1 U8704 ( .A1(n7348), .A2(n8090), .ZN(n10977) );
  NAND2_X1 U8705 ( .A1(n6683), .A2(n11963), .ZN(n7348) );
  OR2_X1 U8706 ( .A1(n7478), .A2(n9690), .ZN(n7705) );
  INV_X1 U8707 ( .A(n14683), .ZN(n14398) );
  NAND2_X1 U8708 ( .A1(n14764), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6708) );
  AND2_X1 U8709 ( .A1(n11752), .A2(n11751), .ZN(n14197) );
  NAND2_X1 U8710 ( .A1(n14265), .A2(n9755), .ZN(n14217) );
  NAND2_X1 U8711 ( .A1(n8003), .A2(n8002), .ZN(n14220) );
  INV_X1 U8712 ( .A(n14088), .ZN(n14233) );
  OR2_X1 U8713 ( .A1(n9756), .A2(P1_U3086), .ZN(n9747) );
  NAND2_X1 U8714 ( .A1(n7507), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7509) );
  AND2_X1 U8715 ( .A1(n8124), .A2(n8123), .ZN(n14250) );
  XNOR2_X1 U8716 ( .A(n8118), .B(P1_IR_REG_25__SCAN_IN), .ZN(n14254) );
  AND2_X1 U8717 ( .A1(n7662), .A2(n7661), .ZN(n11692) );
  XNOR2_X1 U8718 ( .A(n8067), .B(n8066), .ZN(n11756) );
  OR2_X1 U8719 ( .A1(n7968), .A2(n7967), .ZN(n7969) );
  NAND2_X1 U8720 ( .A1(n6564), .A2(n7443), .ZN(n7951) );
  INV_X1 U8721 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10236) );
  INV_X1 U8722 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10125) );
  INV_X1 U8723 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10019) );
  INV_X1 U8724 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9769) );
  INV_X1 U8725 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9750) );
  INV_X1 U8726 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9743) );
  INV_X1 U8727 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9734) );
  INV_X1 U8728 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9724) );
  INV_X1 U8729 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9698) );
  XNOR2_X1 U8730 ( .A(n6759), .B(P2_ADDR_REG_6__SCAN_IN), .ZN(n14382) );
  XNOR2_X1 U8731 ( .A(n14322), .B(n6764), .ZN(n15280) );
  INV_X1 U8732 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6764) );
  XNOR2_X1 U8733 ( .A(n14326), .B(n14327), .ZN(n14383) );
  NAND2_X1 U8734 ( .A1(n7228), .A2(n14334), .ZN(n14386) );
  NAND2_X1 U8735 ( .A1(n14384), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7228) );
  NOR2_X1 U8736 ( .A1(n14386), .A2(n14387), .ZN(n14385) );
  AND2_X1 U8737 ( .A1(n14338), .A2(n14337), .ZN(n14601) );
  NAND2_X1 U8738 ( .A1(n6772), .A2(n6775), .ZN(n14616) );
  NOR2_X1 U8739 ( .A1(n6780), .A2(n14613), .ZN(n6776) );
  INV_X1 U8740 ( .A(n7314), .ZN(n7475) );
  NAND2_X1 U8741 ( .A1(n12420), .A2(n9543), .ZN(n11502) );
  XNOR2_X1 U8742 ( .A(n6718), .B(n7059), .ZN(n12312) );
  NAND2_X1 U8743 ( .A1(n11215), .A2(n9536), .ZN(n11308) );
  NAND2_X1 U8744 ( .A1(n10735), .A2(n9525), .ZN(n10791) );
  INV_X1 U8745 ( .A(n7224), .ZN(n11094) );
  AND2_X1 U8746 ( .A1(n12556), .A2(n6726), .ZN(n6725) );
  OR2_X1 U8747 ( .A1(n12557), .A2(n15067), .ZN(n6726) );
  AOI21_X1 U8748 ( .B1(n12894), .B2(n12695), .A(n12265), .ZN(n6656) );
  NAND2_X1 U8749 ( .A1(n6655), .A2(n15204), .ZN(n6654) );
  OAI21_X1 U8750 ( .B1(n12814), .B2(n15270), .A(n6744), .ZN(P3_U3488) );
  INV_X1 U8751 ( .A(n6745), .ZN(n6744) );
  OAI22_X1 U8752 ( .A1(n12816), .A2(n12884), .B1(n15269), .B2(n12815), .ZN(
        n6745) );
  AOI21_X1 U8753 ( .B1(n6693), .B2(n6692), .A(n6691), .ZN(n6690) );
  NOR2_X1 U8754 ( .A1(n15269), .A2(n12820), .ZN(n6691) );
  AOI21_X1 U8755 ( .B1(n12894), .B2(n12910), .A(n6596), .ZN(n6721) );
  AOI21_X1 U8756 ( .B1(n6693), .B2(n12910), .A(n6689), .ZN(n6688) );
  NOR2_X1 U8757 ( .A1(n15253), .A2(n12896), .ZN(n6689) );
  NAND2_X1 U8758 ( .A1(n9502), .A2(n6649), .ZN(n6648) );
  INV_X1 U8759 ( .A(n7279), .ZN(n12210) );
  OAI21_X1 U8760 ( .B1(n13441), .B2(n13425), .A(n7280), .ZN(n7279) );
  AOI21_X1 U8761 ( .B1(n13437), .B2(n14854), .A(n12209), .ZN(n7280) );
  NAND2_X1 U8762 ( .A1(n9430), .A2(n13497), .ZN(n6662) );
  NAND2_X1 U8763 ( .A1(n14942), .A2(n14921), .ZN(n6813) );
  NAND2_X1 U8764 ( .A1(n7341), .A2(n7339), .ZN(n14549) );
  NAND2_X1 U8765 ( .A1(n11945), .A2(n14162), .ZN(n6747) );
  INV_X1 U8766 ( .A(n7355), .ZN(n7354) );
  OAI21_X1 U8767 ( .B1(n14108), .B2(n14190), .A(n7356), .ZN(n7355) );
  NAND2_X1 U8768 ( .A1(n6709), .A2(n6706), .ZN(P1_U3556) );
  INV_X1 U8769 ( .A(n6707), .ZN(n6706) );
  NAND2_X1 U8770 ( .A1(n14198), .A2(n14766), .ZN(n6709) );
  OAI21_X1 U8771 ( .B1(n14199), .B2(n14190), .A(n6708), .ZN(n6707) );
  NAND2_X1 U8772 ( .A1(n14764), .A2(n14118), .ZN(n6795) );
  AOI21_X1 U8773 ( .B1(n11945), .B2(n14221), .A(n6703), .ZN(n6702) );
  NOR2_X1 U8774 ( .A1(n14756), .A2(n14192), .ZN(n6703) );
  AOI21_X1 U8775 ( .B1(n14755), .B2(P1_REG0_REG_29__SCAN_IN), .A(n6543), .ZN(
        n7134) );
  NAND2_X1 U8776 ( .A1(n6705), .A2(n6540), .ZN(P1_U3524) );
  NAND2_X1 U8777 ( .A1(n14198), .A2(n14756), .ZN(n6705) );
  NAND2_X1 U8778 ( .A1(n14755), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6704) );
  NAND2_X1 U8779 ( .A1(n14606), .A2(n14607), .ZN(n14605) );
  NAND2_X1 U8780 ( .A1(n6781), .A2(n6782), .ZN(n14612) );
  NAND2_X1 U8781 ( .A1(n6774), .A2(n6777), .ZN(n14610) );
  AND2_X1 U8782 ( .A1(n14347), .A2(n14348), .ZN(n14620) );
  NOR2_X1 U8783 ( .A1(n14347), .A2(n14348), .ZN(n14619) );
  XNOR2_X1 U8784 ( .A(n6765), .B(n6513), .ZN(SUB_1596_U4) );
  OAI21_X1 U8785 ( .B1(n14374), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6521), .ZN(
        n6765) );
  INV_X1 U8786 ( .A(n8310), .ZN(n8476) );
  NAND2_X1 U8787 ( .A1(n9389), .A2(n9388), .ZN(n12172) );
  INV_X1 U8788 ( .A(n12172), .ZN(n13540) );
  AND2_X1 U8789 ( .A1(n7466), .A2(n6494), .ZN(n6481) );
  OR2_X1 U8790 ( .A1(n13543), .A2(n13157), .ZN(n6482) );
  AND2_X1 U8791 ( .A1(n13387), .A2(n7241), .ZN(n6484) );
  INV_X1 U8792 ( .A(n12327), .ZN(n7059) );
  INV_X1 U8793 ( .A(n12643), .ZN(n7401) );
  AND2_X1 U8794 ( .A1(n11806), .A2(n6967), .ZN(n6485) );
  INV_X1 U8795 ( .A(n11829), .ZN(n7106) );
  AND2_X1 U8796 ( .A1(n6663), .A2(n13169), .ZN(n6486) );
  INV_X1 U8797 ( .A(n11501), .ZN(n7045) );
  AND3_X1 U8798 ( .A1(n8725), .A2(n9518), .A3(n15190), .ZN(n6487) );
  NAND2_X1 U8799 ( .A1(n14607), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6782) );
  INV_X1 U8800 ( .A(n6782), .ZN(n6779) );
  AND2_X1 U8801 ( .A1(n7439), .A2(n6892), .ZN(n6488) );
  INV_X1 U8802 ( .A(n12576), .ZN(n12897) );
  INV_X1 U8803 ( .A(n12897), .ZN(n6693) );
  INV_X1 U8804 ( .A(n8766), .ZN(n7094) );
  NAND2_X1 U8805 ( .A1(n8978), .A2(n8977), .ZN(n14850) );
  INV_X1 U8806 ( .A(n14850), .ZN(n14917) );
  AND2_X1 U8807 ( .A1(n6562), .A2(n6835), .ZN(n6489) );
  INV_X1 U8808 ( .A(n11893), .ZN(n7287) );
  INV_X1 U8809 ( .A(n7268), .ZN(n7267) );
  OR2_X1 U8810 ( .A1(n12157), .A2(n7269), .ZN(n7268) );
  NAND2_X1 U8811 ( .A1(n7953), .A2(n6583), .ZN(n6490) );
  NOR2_X1 U8812 ( .A1(n13488), .A2(n12156), .ZN(n6491) );
  INV_X1 U8813 ( .A(n9430), .ZN(n13532) );
  AND2_X1 U8814 ( .A1(n9437), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6492) );
  INV_X1 U8815 ( .A(n11945), .ZN(n14193) );
  NAND2_X1 U8816 ( .A1(n11937), .A2(n11936), .ZN(n11945) );
  AND2_X1 U8817 ( .A1(n9193), .A2(n6575), .ZN(n6493) );
  AND2_X1 U8818 ( .A1(n9377), .A2(n9376), .ZN(n6494) );
  AND2_X1 U8819 ( .A1(n6783), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6495) );
  AND2_X1 U8820 ( .A1(n7470), .A2(n9316), .ZN(n6496) );
  INV_X1 U8821 ( .A(n8781), .ZN(n7085) );
  INV_X1 U8822 ( .A(n13696), .ZN(n7333) );
  INV_X1 U8823 ( .A(n8026), .ZN(n6896) );
  INV_X1 U8824 ( .A(n7645), .ZN(n6895) );
  INV_X1 U8825 ( .A(n11804), .ZN(n6699) );
  OR2_X1 U8826 ( .A1(n6734), .A2(P3_IR_REG_25__SCAN_IN), .ZN(n6497) );
  INV_X1 U8827 ( .A(n8602), .ZN(n8336) );
  INV_X1 U8828 ( .A(n13260), .ZN(n6686) );
  INV_X1 U8829 ( .A(n14391), .ZN(n7110) );
  AND2_X1 U8830 ( .A1(n11088), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6498) );
  AND2_X1 U8831 ( .A1(n7062), .A2(n7064), .ZN(n6499) );
  AND2_X1 U8832 ( .A1(n6801), .A2(n6799), .ZN(n6500) );
  INV_X1 U8833 ( .A(n6854), .ZN(n8903) );
  XOR2_X1 U8834 ( .A(n13044), .B(n13438), .Z(n12208) );
  INV_X1 U8835 ( .A(n12208), .ZN(n12173) );
  INV_X1 U8836 ( .A(n13604), .ZN(n7313) );
  INV_X1 U8837 ( .A(n13092), .ZN(n7156) );
  AND2_X1 U8838 ( .A1(n9051), .A2(n9050), .ZN(n6501) );
  AND2_X1 U8839 ( .A1(n9331), .A2(n9330), .ZN(n6502) );
  AND2_X2 U8840 ( .A1(n12118), .A2(n14674), .ZN(n12068) );
  INV_X2 U8841 ( .A(n12068), .ZN(n9615) );
  NOR2_X1 U8842 ( .A1(n14934), .A2(n13177), .ZN(n6503) );
  AND2_X1 U8843 ( .A1(n13409), .A2(n13075), .ZN(n6504) );
  AND2_X1 U8844 ( .A1(n8756), .A2(n8755), .ZN(n6505) );
  INV_X1 U8845 ( .A(n11327), .ZN(n6719) );
  AND2_X1 U8846 ( .A1(n8844), .A2(n7099), .ZN(n6506) );
  NOR2_X1 U8847 ( .A1(n13968), .A2(n7120), .ZN(n7119) );
  NOR2_X1 U8848 ( .A1(n9232), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n8912) );
  AND2_X1 U8849 ( .A1(n10614), .A2(n10638), .ZN(n6507) );
  AND2_X1 U8850 ( .A1(n9533), .A2(n11217), .ZN(n6508) );
  NAND2_X1 U8851 ( .A1(n13520), .A2(n13167), .ZN(n6509) );
  AND2_X1 U8852 ( .A1(n14934), .A2(n10698), .ZN(n6510) );
  AND2_X1 U8853 ( .A1(n6944), .A2(n6942), .ZN(n6511) );
  AND2_X1 U8854 ( .A1(n12654), .A2(n12449), .ZN(n6512) );
  XOR2_X1 U8855 ( .A(n14373), .B(n14372), .Z(n6513) );
  NOR2_X1 U8856 ( .A1(n12428), .A2(n7061), .ZN(n6514) );
  AND2_X1 U8857 ( .A1(n9036), .A2(n9035), .ZN(n6515) );
  INV_X1 U8858 ( .A(n15083), .ZN(n7384) );
  OR2_X1 U8859 ( .A1(n14199), .A2(n14232), .ZN(n6516) );
  AND2_X1 U8860 ( .A1(n11457), .A2(n13172), .ZN(n6517) );
  NOR2_X1 U8861 ( .A1(n12354), .A2(n12285), .ZN(n6518) );
  OR2_X1 U8862 ( .A1(n8373), .A2(n8372), .ZN(n11120) );
  OR2_X1 U8863 ( .A1(n11482), .A2(n11483), .ZN(n6519) );
  AND2_X1 U8864 ( .A1(n7049), .A2(n11307), .ZN(n6520) );
  OR2_X1 U8865 ( .A1(n14365), .A2(n14366), .ZN(n6521) );
  OR2_X1 U8866 ( .A1(n14987), .A2(n11089), .ZN(n6522) );
  OR2_X1 U8867 ( .A1(n15057), .A2(n11091), .ZN(n6523) );
  INV_X1 U8868 ( .A(n9174), .ZN(n7468) );
  AND2_X1 U8869 ( .A1(n7504), .A2(n7611), .ZN(n6524) );
  AND2_X1 U8870 ( .A1(n9242), .A2(n9241), .ZN(n6525) );
  AND2_X1 U8871 ( .A1(n13525), .A2(n13073), .ZN(n6526) );
  AND2_X1 U8872 ( .A1(n9275), .A2(n9274), .ZN(n6527) );
  INV_X1 U8873 ( .A(n12264), .ZN(n6680) );
  NOR2_X1 U8874 ( .A1(n12875), .A2(n12769), .ZN(n6528) );
  INV_X1 U8875 ( .A(n12198), .ZN(n7263) );
  INV_X1 U8876 ( .A(n12226), .ZN(n7393) );
  INV_X1 U8877 ( .A(n11975), .ZN(n14039) );
  INV_X1 U8878 ( .A(n11836), .ZN(n6945) );
  AND2_X1 U8879 ( .A1(n12731), .A2(n7084), .ZN(n6529) );
  OR2_X1 U8880 ( .A1(n8575), .A2(SI_2_), .ZN(n6530) );
  OR2_X1 U8881 ( .A1(n14317), .A2(n14316), .ZN(n6531) );
  INV_X1 U8882 ( .A(n12204), .ZN(n7254) );
  AOI21_X1 U8883 ( .B1(n6777), .B2(n6779), .A(n6776), .ZN(n6775) );
  OR2_X1 U8884 ( .A1(n9122), .A2(n9121), .ZN(n6532) );
  OR2_X1 U8885 ( .A1(n9295), .A2(n9294), .ZN(n6533) );
  AND2_X1 U8886 ( .A1(n11715), .A2(n11714), .ZN(n6534) );
  OR2_X1 U8887 ( .A1(n9068), .A2(n9069), .ZN(n6535) );
  INV_X1 U8888 ( .A(n7260), .ZN(n7259) );
  NOR2_X1 U8889 ( .A1(n7261), .A2(n12200), .ZN(n7260) );
  AND2_X1 U8890 ( .A1(n12185), .A2(n6833), .ZN(n6536) );
  AND2_X1 U8891 ( .A1(n13978), .A2(n7119), .ZN(n6537) );
  AND2_X1 U8892 ( .A1(n9458), .A2(n9457), .ZN(n6538) );
  NOR2_X1 U8893 ( .A1(n15138), .A2(n12222), .ZN(n6539) );
  AND2_X1 U8894 ( .A1(n6516), .A2(n6704), .ZN(n6540) );
  NOR2_X1 U8895 ( .A1(n11829), .A2(n13764), .ZN(n6541) );
  NOR2_X1 U8896 ( .A1(n13507), .A2(n13165), .ZN(n6542) );
  NOR2_X1 U8897 ( .A1(n14108), .A2(n14232), .ZN(n6543) );
  NAND2_X1 U8898 ( .A1(n6479), .A2(n9685), .ZN(n9231) );
  INV_X1 U8899 ( .A(n9231), .ZN(n7206) );
  NOR2_X1 U8900 ( .A1(n11837), .A2(n11641), .ZN(n6544) );
  NOR2_X1 U8901 ( .A1(n13525), .A2(n13073), .ZN(n6545) );
  NOR2_X1 U8902 ( .A1(n14220), .A2(n13752), .ZN(n6546) );
  NOR2_X1 U8903 ( .A1(n12285), .A2(n12408), .ZN(n6547) );
  NOR2_X1 U8904 ( .A1(n14088), .A2(n13712), .ZN(n6548) );
  NOR2_X1 U8905 ( .A1(n13738), .A2(n13758), .ZN(n6549) );
  INV_X1 U8906 ( .A(n6919), .ZN(n6918) );
  NAND2_X1 U8907 ( .A1(n6920), .A2(n7323), .ZN(n6919) );
  OR2_X1 U8908 ( .A1(n14273), .A2(n7237), .ZN(n6550) );
  AND2_X1 U8909 ( .A1(n8232), .A2(n7415), .ZN(n7414) );
  INV_X1 U8910 ( .A(n12329), .ZN(n7063) );
  AND2_X1 U8911 ( .A1(n7402), .A2(n12249), .ZN(n6551) );
  AND2_X1 U8912 ( .A1(n8263), .A2(n8262), .ZN(n8310) );
  OR2_X1 U8913 ( .A1(n7184), .A2(n7183), .ZN(n6552) );
  NAND2_X1 U8914 ( .A1(n14088), .A2(n13756), .ZN(n6553) );
  INV_X1 U8915 ( .A(n6553), .ZN(n7362) );
  NOR2_X1 U8916 ( .A1(n7466), .A2(n6494), .ZN(n6554) );
  OR2_X1 U8917 ( .A1(n9091), .A2(n9090), .ZN(n6555) );
  AND3_X1 U8918 ( .A1(n8795), .A2(n8794), .A3(n12643), .ZN(n6556) );
  NAND4_X1 U8919 ( .A1(n7292), .A2(n7503), .A3(n7734), .A4(n7476), .ZN(n6557)
         );
  INV_X1 U8920 ( .A(n6869), .ZN(n6868) );
  NAND2_X1 U8921 ( .A1(n13379), .A2(n6871), .ZN(n6869) );
  AND2_X1 U8922 ( .A1(n7562), .A2(SI_10_), .ZN(n6558) );
  AND2_X1 U8923 ( .A1(n11915), .A2(n7283), .ZN(n6559) );
  INV_X1 U8924 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8879) );
  OR2_X1 U8925 ( .A1(n7474), .A2(n7473), .ZN(n6560) );
  NAND2_X1 U8926 ( .A1(n8726), .A2(n6735), .ZN(n6561) );
  INV_X1 U8927 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9700) );
  INV_X1 U8928 ( .A(n7400), .ZN(n7399) );
  NAND2_X1 U8929 ( .A1(n7401), .A2(n12249), .ZN(n7400) );
  XNOR2_X1 U8930 ( .A(n11445), .B(n6682), .ZN(n11369) );
  AND2_X1 U8931 ( .A1(n12199), .A2(n12198), .ZN(n6562) );
  INV_X1 U8932 ( .A(n7271), .ZN(n7270) );
  NAND2_X1 U8933 ( .A1(n7272), .A2(n12154), .ZN(n7271) );
  AND2_X1 U8934 ( .A1(n11369), .A2(n7165), .ZN(n6563) );
  AND2_X1 U8935 ( .A1(n7442), .A2(n7441), .ZN(n6564) );
  INV_X1 U8936 ( .A(n8060), .ZN(n7345) );
  NOR2_X2 U8937 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n8060) );
  NAND2_X1 U8938 ( .A1(n7986), .A2(n7985), .ZN(n14043) );
  INV_X1 U8939 ( .A(n14043), .ZN(n14165) );
  OR2_X1 U8940 ( .A1(n12195), .A2(n6836), .ZN(n6565) );
  MUX2_X1 U8941 ( .A(n14132), .B(n13749), .S(n11946), .Z(n11903) );
  INV_X1 U8942 ( .A(n11903), .ZN(n6958) );
  INV_X1 U8943 ( .A(n11805), .ZN(n6967) );
  AND2_X1 U8944 ( .A1(n12326), .A2(n12598), .ZN(n6566) );
  OR2_X1 U8945 ( .A1(n12809), .A2(n12805), .ZN(n6567) );
  OR2_X1 U8946 ( .A1(n11126), .A2(n11090), .ZN(n6568) );
  OR2_X1 U8947 ( .A1(n9277), .A2(n6527), .ZN(n6569) );
  AND2_X1 U8948 ( .A1(n15110), .A2(n8747), .ZN(n6570) );
  AND2_X1 U8949 ( .A1(n7331), .A2(n6922), .ZN(n6571) );
  AND2_X1 U8950 ( .A1(n7488), .A2(n12233), .ZN(n6572) );
  AND2_X1 U8951 ( .A1(n8814), .A2(n8813), .ZN(n6573) );
  INV_X1 U8952 ( .A(n7131), .ZN(n7130) );
  NOR2_X1 U8953 ( .A1(n11963), .A2(n7132), .ZN(n7131) );
  AND2_X1 U8954 ( .A1(n7079), .A2(n7414), .ZN(n6574) );
  AND2_X1 U8955 ( .A1(n9191), .A2(n9190), .ZN(n6575) );
  AND2_X1 U8956 ( .A1(n6484), .A2(n6509), .ZN(n6576) );
  OR2_X1 U8957 ( .A1(n11932), .A2(n11931), .ZN(n6577) );
  AND2_X1 U8958 ( .A1(n8793), .A2(n12658), .ZN(n6578) );
  NAND2_X1 U8959 ( .A1(n13972), .A2(n12100), .ZN(n6579) );
  AND2_X1 U8960 ( .A1(n6502), .A2(n7004), .ZN(n6580) );
  NAND2_X1 U8961 ( .A1(n6917), .A2(n6920), .ZN(n6916) );
  OR2_X1 U8962 ( .A1(n7246), .A2(n6829), .ZN(n6581) );
  NAND2_X1 U8963 ( .A1(n12980), .A2(n12979), .ZN(n6582) );
  INV_X1 U8964 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6965) );
  INV_X1 U8965 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7232) );
  AND2_X1 U8966 ( .A1(n8060), .A2(n7344), .ZN(n6583) );
  XNOR2_X1 U8967 ( .A(n8241), .B(P3_IR_REG_27__SCAN_IN), .ZN(n9659) );
  NAND2_X1 U8968 ( .A1(n6911), .A2(n7315), .ZN(n6921) );
  INV_X1 U8969 ( .A(n13611), .ZN(n7332) );
  INV_X1 U8970 ( .A(n8965), .ZN(n9118) );
  INV_X1 U8971 ( .A(n8227), .ZN(n8522) );
  NAND2_X1 U8972 ( .A1(n8667), .A2(n8666), .ZN(n12446) );
  INV_X1 U8973 ( .A(n12446), .ZN(n12584) );
  AND2_X1 U8974 ( .A1(n7596), .A2(n7435), .ZN(n6584) );
  NOR2_X1 U8975 ( .A1(n12465), .A2(n12466), .ZN(n6585) );
  AND2_X1 U8976 ( .A1(n11571), .A2(n8099), .ZN(n6586) );
  INV_X1 U8977 ( .A(n7590), .ZN(n6891) );
  INV_X1 U8978 ( .A(n7208), .ZN(n13392) );
  INV_X1 U8979 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7237) );
  AND2_X1 U8980 ( .A1(n7146), .A2(n7149), .ZN(n6587) );
  NAND4_X1 U8981 ( .A1(n8823), .A2(n9650), .A3(n8780), .A4(n8779), .ZN(n6588)
         );
  INV_X1 U8982 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8964) );
  NAND2_X1 U8983 ( .A1(n8696), .A2(n8695), .ZN(n6589) );
  AND4_X1 U8984 ( .A1(n8443), .A2(n8442), .A3(n8441), .A4(n8440), .ZN(n12797)
         );
  INV_X1 U8985 ( .A(n12797), .ZN(n14956) );
  INV_X1 U8986 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8711) );
  AND2_X1 U8987 ( .A1(n7169), .A2(n11725), .ZN(n6590) );
  INV_X1 U8988 ( .A(n7487), .ZN(n7382) );
  INV_X1 U8989 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10368) );
  INV_X1 U8990 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10020) );
  NAND2_X2 U8991 ( .A1(n10773), .A2(n14865), .ZN(n14871) );
  INV_X1 U8992 ( .A(n11455), .ZN(n6825) );
  INV_X1 U8993 ( .A(n12884), .ZN(n6692) );
  INV_X1 U8994 ( .A(SI_18_), .ZN(n10098) );
  INV_X1 U8995 ( .A(n12754), .ZN(n7087) );
  NOR2_X1 U8996 ( .A1(n10837), .A2(n7475), .ZN(n6591) );
  AND2_X1 U8997 ( .A1(n7273), .A2(n10693), .ZN(n6863) );
  INV_X2 U8998 ( .A(n9650), .ZN(n10640) );
  INV_X1 U8999 ( .A(n11587), .ZN(n11589) );
  OR2_X1 U9000 ( .A1(n8878), .A2(n9194), .ZN(n6592) );
  INV_X1 U9001 ( .A(n13500), .ZN(n7207) );
  AND2_X1 U9002 ( .A1(n11374), .A2(n11373), .ZN(n6593) );
  AND2_X1 U9003 ( .A1(n8196), .A2(n7009), .ZN(n6594) );
  NAND2_X1 U9004 ( .A1(n11008), .A2(n14735), .ZN(n11007) );
  INV_X1 U9005 ( .A(n11007), .ZN(n7107) );
  AND2_X1 U9006 ( .A1(n6864), .A2(n10693), .ZN(n6595) );
  NOR2_X1 U9007 ( .A1(n15253), .A2(n12892), .ZN(n6596) );
  AND2_X1 U9008 ( .A1(n9417), .A2(n12959), .ZN(n6597) );
  AND2_X1 U9009 ( .A1(n6896), .A2(n6894), .ZN(n6598) );
  INV_X1 U9010 ( .A(n7607), .ZN(n7447) );
  INV_X1 U9011 ( .A(n15253), .ZN(n15252) );
  INV_X1 U9012 ( .A(n11445), .ZN(n6664) );
  AND2_X1 U9013 ( .A1(n9574), .A2(n10866), .ZN(n14960) );
  AND2_X2 U9014 ( .A1(n10517), .A2(n10025), .ZN(n14756) );
  INV_X1 U9015 ( .A(n14439), .ZN(n12538) );
  INV_X1 U9016 ( .A(n15183), .ZN(n15130) );
  NAND2_X1 U9017 ( .A1(n10930), .A2(n10929), .ZN(n15183) );
  AND2_X1 U9018 ( .A1(n9525), .A2(n9521), .ZN(n6599) );
  INV_X1 U9019 ( .A(n14753), .ZN(n14588) );
  INV_X1 U9020 ( .A(n14673), .ZN(n6700) );
  INV_X1 U9021 ( .A(n14851), .ZN(n7202) );
  AND2_X1 U9022 ( .A1(n10563), .A2(n12550), .ZN(n15199) );
  NAND2_X1 U9023 ( .A1(n7202), .A2(n14917), .ZN(n14852) );
  INV_X1 U9024 ( .A(n14852), .ZN(n7201) );
  OR2_X1 U9025 ( .A1(n14439), .A2(n12531), .ZN(n6600) );
  AND2_X1 U9026 ( .A1(n7188), .A2(n7192), .ZN(n6601) );
  XNOR2_X1 U9027 ( .A(n8574), .B(n8709), .ZN(n12523) );
  INV_X1 U9028 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n6716) );
  INV_X1 U9029 ( .A(n14470), .ZN(n12546) );
  INV_X1 U9030 ( .A(n8889), .ZN(n13577) );
  INV_X1 U9031 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7227) );
  AND2_X1 U9032 ( .A1(n10431), .A2(n10432), .ZN(n6602) );
  INV_X1 U9033 ( .A(SI_25_), .ZN(n7451) );
  INV_X1 U9034 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7231) );
  INV_X1 U9035 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6760) );
  NAND3_X1 U9036 ( .A1(n8815), .A2(n8814), .A3(n6603), .ZN(n6714) );
  AOI211_X1 U9037 ( .C1(n8769), .C2(n7489), .A(n8768), .B(n12773), .ZN(n6610)
         );
  NOR2_X1 U9038 ( .A1(n8790), .A2(n8789), .ZN(n6750) );
  NOR3_X1 U9039 ( .A1(n8731), .A2(n8730), .A3(n12213), .ZN(n8735) );
  AOI21_X1 U9040 ( .B1(n15076), .B2(n8753), .A(n8752), .ZN(n8754) );
  OAI211_X1 U9041 ( .C1(n8744), .C2(n8743), .A(n15121), .B(n8742), .ZN(n8748)
         );
  NAND2_X1 U9042 ( .A1(n8722), .A2(n8721), .ZN(n6613) );
  OAI21_X2 U9043 ( .B1(n8683), .B2(n8214), .A(n8215), .ZN(n8694) );
  OAI21_X2 U9044 ( .B1(n8615), .B2(n8614), .A(n8200), .ZN(n8625) );
  INV_X1 U9045 ( .A(n8819), .ZN(n8845) );
  NAND2_X1 U9046 ( .A1(n8149), .A2(n8148), .ZN(n8305) );
  NAND2_X1 U9047 ( .A1(n6710), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8470) );
  NAND2_X1 U9048 ( .A1(n6605), .A2(n8851), .ZN(n8862) );
  NAND3_X1 U9049 ( .A1(n6694), .A2(n6636), .A3(n7025), .ZN(n6605) );
  NAND2_X1 U9050 ( .A1(n8398), .A2(n8165), .ZN(n8416) );
  NAND2_X1 U9051 ( .A1(n12558), .A2(n12560), .ZN(n8844) );
  NAND2_X1 U9052 ( .A1(n8177), .A2(n8176), .ZN(n8178) );
  OAI21_X1 U9053 ( .B1(n8634), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n8206), .ZN(
        n8645) );
  NAND2_X1 U9054 ( .A1(n6606), .A2(n8821), .ZN(n8818) );
  NAND3_X1 U9055 ( .A1(n6714), .A2(n6711), .A3(n8811), .ZN(n6606) );
  NAND2_X1 U9056 ( .A1(n6613), .A2(n6611), .ZN(n8725) );
  OAI211_X1 U9057 ( .C1(n8810), .C2(n8809), .A(n12587), .B(n8808), .ZN(n8815)
         );
  NAND2_X1 U9058 ( .A1(n8796), .A2(n6556), .ZN(n8797) );
  OAI21_X1 U9059 ( .B1(n6610), .B2(n8773), .A(n6609), .ZN(n8776) );
  OAI21_X1 U9060 ( .B1(n10733), .B2(n10944), .A(n9518), .ZN(n6612) );
  NAND2_X1 U9061 ( .A1(n8710), .A2(n8709), .ZN(n8715) );
  NAND2_X1 U9062 ( .A1(n7027), .A2(n8212), .ZN(n8683) );
  NAND2_X1 U9063 ( .A1(n8686), .A2(n8685), .ZN(n12576) );
  OAI21_X1 U9064 ( .B1(n8645), .B2(n8644), .A(n8207), .ZN(n8658) );
  NAND2_X1 U9065 ( .A1(n8206), .A2(n8205), .ZN(n8634) );
  NAND2_X1 U9066 ( .A1(n8396), .A2(n8395), .ZN(n8398) );
  NAND2_X1 U9067 ( .A1(n8601), .A2(n8199), .ZN(n8615) );
  NAND2_X1 U9068 ( .A1(n8847), .A2(n10937), .ZN(n6677) );
  OAI21_X1 U9069 ( .B1(n11867), .B2(n7302), .A(n6614), .ZN(n6950) );
  NAND3_X1 U9070 ( .A1(n11901), .A2(n11900), .A3(n6955), .ZN(n6954) );
  OAI21_X1 U9071 ( .B1(n11952), .B2(n11951), .A(n6617), .ZN(n11997) );
  NAND2_X1 U9072 ( .A1(n11952), .A2(n11950), .ZN(n6617) );
  NAND2_X1 U9073 ( .A1(n8695), .A2(n8216), .ZN(n8269) );
  NAND2_X1 U9074 ( .A1(n8599), .A2(n8598), .ZN(n8601) );
  NAND2_X1 U9075 ( .A1(n6884), .A2(n7566), .ZN(n7848) );
  NAND2_X1 U9076 ( .A1(n6953), .A2(n11872), .ZN(n11877) );
  NAND2_X1 U9077 ( .A1(n12588), .A2(n12587), .ZN(n12586) );
  NAND2_X1 U9078 ( .A1(n7066), .A2(n7396), .ZN(n11326) );
  AND3_X1 U9079 ( .A1(n8297), .A2(n8295), .A3(n8296), .ZN(n6720) );
  NAND2_X1 U9080 ( .A1(n15191), .A2(n15190), .ZN(n15193) );
  NAND2_X1 U9081 ( .A1(n12893), .A2(n6721), .ZN(P3_U3456) );
  NAND2_X1 U9082 ( .A1(n7185), .A2(n7186), .ZN(n7189) );
  AOI21_X2 U9083 ( .B1(n13029), .B2(n13025), .A(n13027), .ZN(n13112) );
  NOR2_X1 U9084 ( .A1(n10225), .A2(n10224), .ZN(n10229) );
  OAI21_X1 U9085 ( .B1(n11229), .B2(n7160), .A(n7157), .ZN(n6619) );
  INV_X1 U9086 ( .A(n11230), .ZN(n7162) );
  XNOR2_X1 U9087 ( .A(n7540), .B(SI_4_), .ZN(n7731) );
  NAND2_X1 U9088 ( .A1(n7937), .A2(n10059), .ZN(n6625) );
  INV_X1 U9089 ( .A(n13131), .ZN(n7155) );
  NAND2_X1 U9090 ( .A1(n7443), .A2(n7442), .ZN(n7949) );
  NAND2_X1 U9091 ( .A1(n7633), .A2(n7607), .ZN(n7621) );
  XNOR2_X1 U9092 ( .A(n12996), .B(n12997), .ZN(n13123) );
  NAND2_X1 U9093 ( .A1(n8092), .A2(n8091), .ZN(n11188) );
  NAND2_X2 U9094 ( .A1(n13961), .A2(n7372), .ZN(n7370) );
  NAND2_X1 U9095 ( .A1(n14107), .A2(n14756), .ZN(n7135) );
  NAND2_X1 U9096 ( .A1(n14107), .A2(n14766), .ZN(n7357) );
  NAND2_X2 U9097 ( .A1(n8098), .A2(n8097), .ZN(n11569) );
  NAND2_X2 U9098 ( .A1(n8101), .A2(n8100), .ZN(n14081) );
  NOR2_X1 U9099 ( .A1(n14115), .A2(n6797), .ZN(n14200) );
  OAI22_X2 U9100 ( .A1(n11954), .A2(n10128), .B1(n13772), .B2(n11778), .ZN(
        n10111) );
  NAND2_X1 U9101 ( .A1(n7370), .A2(n7369), .ZN(n13928) );
  NAND2_X1 U9102 ( .A1(n7353), .A2(n7352), .ZN(n13975) );
  INV_X2 U9103 ( .A(n7680), .ZN(n10135) );
  INV_X1 U9104 ( .A(n7507), .ZN(n7506) );
  NAND2_X1 U9105 ( .A1(n8083), .A2(n8082), .ZN(n10509) );
  NAND2_X1 U9106 ( .A1(n8089), .A2(n8088), .ZN(n11006) );
  NAND2_X1 U9107 ( .A1(n8353), .A2(n8157), .ZN(n8370) );
  NAND2_X1 U9108 ( .A1(n8694), .A2(n8693), .ZN(n8695) );
  NAND2_X1 U9109 ( .A1(n8535), .A2(n8534), .ZN(n8537) );
  OAI22_X1 U9110 ( .A1(n8269), .A2(n8268), .B1(P1_DATAO_REG_30__SCAN_IN), .B2(
        n11999), .ZN(n8271) );
  NAND2_X1 U9111 ( .A1(n8537), .A2(n8192), .ZN(n8555) );
  NAND2_X1 U9112 ( .A1(n8370), .A2(n8158), .ZN(n8160) );
  NAND2_X1 U9113 ( .A1(n6635), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8206) );
  NAND2_X1 U9114 ( .A1(n15106), .A2(n8749), .ZN(n15089) );
  XNOR2_X1 U9115 ( .A(n6634), .B(n12550), .ZN(n6633) );
  NAND2_X1 U9116 ( .A1(n7067), .A2(n7068), .ZN(n15122) );
  INV_X1 U9117 ( .A(n6730), .ZN(n6729) );
  NAND2_X1 U9118 ( .A1(n7609), .A2(n11559), .ZN(n6731) );
  NAND2_X1 U9119 ( .A1(n11575), .A2(n11968), .ZN(n11574) );
  NAND2_X1 U9120 ( .A1(n7861), .A2(n7860), .ZN(n11316) );
  INV_X1 U9121 ( .A(n13979), .ZN(n6742) );
  NAND2_X1 U9122 ( .A1(n7135), .A2(n7134), .ZN(P1_U3525) );
  NAND2_X1 U9123 ( .A1(n7357), .A2(n7354), .ZN(P1_U3557) );
  NAND2_X2 U9124 ( .A1(n7964), .A2(n7963), .ZN(n14054) );
  NOR2_X1 U9125 ( .A1(n10492), .A2(n8313), .ZN(n10491) );
  NOR2_X2 U9126 ( .A1(n15037), .A2(n7212), .ZN(n11091) );
  OAI21_X1 U9127 ( .B1(n10435), .B2(n10445), .A(n10434), .ZN(n10492) );
  NOR2_X1 U9128 ( .A1(n11584), .A2(n6754), .ZN(n12464) );
  NOR2_X1 U9129 ( .A1(n11418), .A2(n11417), .ZN(n11420) );
  NAND2_X1 U9130 ( .A1(n7101), .A2(n7100), .ZN(n6624) );
  NAND2_X1 U9131 ( .A1(n6751), .A2(n6568), .ZN(n7214) );
  OAI21_X1 U9132 ( .B1(n11585), .B2(n7219), .A(n7218), .ZN(n12493) );
  NAND2_X1 U9133 ( .A1(n10435), .A2(n10445), .ZN(n10434) );
  NAND2_X1 U9134 ( .A1(n6728), .A2(n10434), .ZN(n7216) );
  NAND2_X1 U9135 ( .A1(n6633), .A2(n6632), .ZN(n6636) );
  INV_X1 U9136 ( .A(n8025), .ZN(n7120) );
  NAND2_X1 U9137 ( .A1(n13935), .A2(n14664), .ZN(n6801) );
  INV_X1 U9138 ( .A(n8847), .ZN(n6627) );
  NAND2_X1 U9139 ( .A1(n6629), .A2(n6628), .ZN(n8784) );
  NAND2_X1 U9140 ( .A1(n6630), .A2(n12724), .ZN(n6629) );
  OR2_X1 U9141 ( .A1(n8777), .A2(n6631), .ZN(n6630) );
  NAND4_X2 U9142 ( .A1(n8280), .A2(n8281), .A3(n8282), .A4(n8279), .ZN(n10737)
         );
  AOI21_X1 U9143 ( .B1(n8748), .B2(n6570), .A(n6715), .ZN(n8752) );
  INV_X1 U9144 ( .A(n8204), .ZN(n6635) );
  NAND2_X1 U9145 ( .A1(n8557), .A2(n8194), .ZN(n8569) );
  NOR2_X2 U9146 ( .A1(n10737), .A2(n10646), .ZN(n10935) );
  INV_X1 U9147 ( .A(n6798), .ZN(n6797) );
  NAND2_X1 U9148 ( .A1(n15193), .A2(n8723), .ZN(n11039) );
  AOI21_X2 U9149 ( .B1(n13932), .B2(n13930), .A(n13929), .ZN(n14114) );
  NAND2_X1 U9150 ( .A1(n8179), .A2(n8180), .ZN(n8468) );
  NAND2_X1 U9151 ( .A1(n10688), .A2(n10687), .ZN(n14840) );
  NAND2_X1 U9152 ( .A1(n13265), .A2(n12169), .ZN(n13248) );
  NAND2_X1 U9153 ( .A1(n12160), .A2(n12159), .ZN(n13310) );
  NAND2_X1 U9154 ( .A1(n13413), .A2(n12147), .ZN(n12150) );
  XNOR2_X1 U9155 ( .A(n6909), .B(n7313), .ZN(n13610) );
  OAI21_X1 U9156 ( .B1(n10099), .B2(n10100), .A(n7304), .ZN(n9628) );
  NAND2_X1 U9157 ( .A1(n8160), .A2(n8159), .ZN(n8384) );
  AND2_X4 U9158 ( .A1(n9634), .A2(n10518), .ZN(n12118) );
  NAND2_X1 U9159 ( .A1(n6637), .A2(n12432), .ZN(P3_U3180) );
  NAND2_X1 U9160 ( .A1(n6638), .A2(n14960), .ZN(n6637) );
  XNOR2_X1 U9161 ( .A(n12427), .B(n12428), .ZN(n6638) );
  NAND2_X1 U9162 ( .A1(n6639), .A2(n10792), .ZN(n9528) );
  NAND2_X1 U9163 ( .A1(n9525), .A2(n7033), .ZN(n6639) );
  NAND2_X1 U9164 ( .A1(n11561), .A2(n7031), .ZN(n14958) );
  NAND2_X1 U9165 ( .A1(n7542), .A2(n7541), .ZN(n7742) );
  MUX2_X2 U9166 ( .A(n14101), .B(n14191), .S(n14766), .Z(n14102) );
  NAND2_X1 U9167 ( .A1(n6642), .A2(n6640), .ZN(n13539) );
  NAND2_X1 U9168 ( .A1(n14940), .A2(n6641), .ZN(n6640) );
  OR2_X1 U9169 ( .A1(n13538), .A2(n14940), .ZN(n6642) );
  NAND2_X1 U9170 ( .A1(n6644), .A2(n6643), .ZN(n13445) );
  NAND2_X1 U9171 ( .A1(n14951), .A2(n9398), .ZN(n6643) );
  OR2_X1 U9172 ( .A1(n13538), .A2(n14951), .ZN(n6644) );
  INV_X1 U9173 ( .A(n6645), .ZN(n11470) );
  NAND2_X1 U9174 ( .A1(n10529), .A2(n14708), .ZN(n14673) );
  NAND2_X1 U9175 ( .A1(n7104), .A2(n9755), .ZN(n7105) );
  AND2_X1 U9176 ( .A1(n10131), .A2(n10130), .ZN(n10133) );
  INV_X1 U9177 ( .A(n6701), .ZN(n13997) );
  NOR2_X2 U9178 ( .A1(n13936), .A2(n13915), .ZN(n8070) );
  INV_X1 U9179 ( .A(n9692), .ZN(n7205) );
  AOI21_X2 U9180 ( .B1(n12613), .B2(n8669), .A(n8668), .ZN(n12588) );
  NAND3_X1 U9181 ( .A1(n6560), .A2(n6646), .A3(n6968), .ZN(n6970) );
  NAND4_X1 U9182 ( .A1(n9505), .A2(n6648), .A3(n9504), .A4(n9506), .ZN(
        P2_U3328) );
  NAND2_X2 U9183 ( .A1(n12615), .A2(n12614), .ZN(n12613) );
  INV_X1 U9184 ( .A(n9211), .ZN(n7461) );
  NAND2_X1 U9185 ( .A1(n6555), .A2(n6651), .ZN(n9105) );
  NAND2_X1 U9186 ( .A1(n6653), .A2(n6652), .ZN(n6651) );
  NAND2_X1 U9187 ( .A1(n9091), .A2(n9090), .ZN(n6653) );
  XNOR2_X1 U9188 ( .A(n6695), .B(n6680), .ZN(n12809) );
  NAND3_X1 U9189 ( .A1(n6567), .A2(n6656), .A3(n6654), .ZN(P3_U3204) );
  AND2_X1 U9190 ( .A1(n8300), .A2(n8299), .ZN(n6657) );
  NAND3_X1 U9191 ( .A1(n7465), .A2(n7462), .A3(n6658), .ZN(n6988) );
  NAND2_X1 U9192 ( .A1(n13112), .A2(n13113), .ZN(n13111) );
  NAND2_X2 U9193 ( .A1(n6661), .A2(n6659), .ZN(n13141) );
  NOR2_X1 U9194 ( .A1(n11371), .A2(n11296), .ZN(n7164) );
  AOI22_X2 U9195 ( .A1(n12974), .A2(n12973), .B1(n12972), .B2(n12971), .ZN(
        n13070) );
  AND2_X4 U9196 ( .A1(n6480), .A2(n9684), .ZN(n9437) );
  NAND2_X1 U9197 ( .A1(n13432), .A2(n6662), .ZN(P2_U3530) );
  NOR2_X4 U9198 ( .A1(n13374), .A2(n13562), .ZN(n13361) );
  INV_X1 U9199 ( .A(n12673), .ZN(n6666) );
  INV_X1 U9200 ( .A(n10491), .ZN(n6728) );
  XNOR2_X2 U9201 ( .A(n6673), .B(n12540), .ZN(n12495) );
  NAND2_X1 U9202 ( .A1(n7026), .A2(n6507), .ZN(n6676) );
  NAND3_X1 U9203 ( .A1(n8844), .A2(n8845), .A3(n6678), .ZN(n8846) );
  NAND2_X1 U9204 ( .A1(n8203), .A2(n8202), .ZN(n8204) );
  XNOR2_X1 U9205 ( .A(n8271), .B(n8270), .ZN(n12949) );
  NAND2_X1 U9206 ( .A1(n8625), .A2(n8624), .ZN(n8203) );
  NAND2_X1 U9207 ( .A1(n6713), .A2(n6712), .ZN(n6711) );
  INV_X1 U9208 ( .A(n10229), .ZN(n7185) );
  NAND2_X1 U9209 ( .A1(n11228), .A2(n11227), .ZN(n11229) );
  NOR2_X1 U9210 ( .A1(n10184), .A2(n10185), .ZN(n10225) );
  NAND2_X1 U9211 ( .A1(n6853), .A2(n6856), .ZN(n6854) );
  OAI21_X1 U9212 ( .B1(n13053), .B2(n13052), .A(n12995), .ZN(n12996) );
  NAND2_X1 U9213 ( .A1(n7370), .A2(n7368), .ZN(n13930) );
  NAND2_X1 U9214 ( .A1(n13130), .A2(n12985), .ZN(n13029) );
  NAND2_X1 U9215 ( .A1(n14200), .A2(n14766), .ZN(n6796) );
  NAND2_X1 U9216 ( .A1(n6796), .A2(n6795), .ZN(n14119) );
  INV_X1 U9217 ( .A(n7601), .ZN(n7602) );
  NAND2_X1 U9218 ( .A1(n13302), .A2(n13301), .ZN(n12165) );
  NAND2_X1 U9219 ( .A1(n7603), .A2(n7604), .ZN(n7646) );
  OAI21_X1 U9220 ( .B1(n12895), .B2(n15252), .A(n6688), .ZN(P3_U3455) );
  OAI21_X1 U9221 ( .B1(n12895), .B2(n15270), .A(n6690), .ZN(P3_U3487) );
  NAND2_X1 U9222 ( .A1(n7098), .A2(n8811), .ZN(n6695) );
  NAND2_X1 U9223 ( .A1(n7098), .A2(n7096), .ZN(n7101) );
  NAND2_X1 U9224 ( .A1(n7150), .A2(n7147), .ZN(n13130) );
  NOR2_X2 U9225 ( .A1(n14996), .A2(n14995), .ZN(n14994) );
  NAND2_X1 U9226 ( .A1(n6696), .A2(n6899), .ZN(n7288) );
  NAND3_X1 U9227 ( .A1(n11925), .A2(n6902), .A3(n6577), .ZN(n6696) );
  NAND2_X1 U9228 ( .A1(n11910), .A2(n7283), .ZN(n7282) );
  NAND2_X1 U9229 ( .A1(n11906), .A2(n6697), .ZN(n11910) );
  NAND2_X1 U9230 ( .A1(n6950), .A2(n6948), .ZN(n6953) );
  OAI22_X1 U9231 ( .A1(n11807), .A2(n6485), .B1(n11806), .B2(n6967), .ZN(
        n11810) );
  INV_X1 U9232 ( .A(n11757), .ZN(n11755) );
  OAI22_X1 U9233 ( .A1(n11817), .A2(n7300), .B1(n11818), .B2(n7299), .ZN(
        n11823) );
  NAND2_X1 U9234 ( .A1(n11896), .A2(n11897), .ZN(n11895) );
  NAND2_X1 U9235 ( .A1(n11916), .A2(n6938), .ZN(n11918) );
  NAND2_X1 U9236 ( .A1(n7294), .A2(n7293), .ZN(n7295) );
  NAND2_X1 U9237 ( .A1(n6943), .A2(n6944), .ZN(n11844) );
  NAND2_X1 U9238 ( .A1(n7329), .A2(n7327), .ZN(n13613) );
  NAND2_X1 U9239 ( .A1(n6930), .A2(n6928), .ZN(n12027) );
  NOR2_X2 U9240 ( .A1(n10764), .A2(n10765), .ZN(n10837) );
  NOR2_X1 U9241 ( .A1(n9628), .A2(n9629), .ZN(n10763) );
  NAND2_X1 U9242 ( .A1(n14400), .A2(n11839), .ZN(n11573) );
  NOR2_X2 U9243 ( .A1(n14132), .A2(n13997), .ZN(n13984) );
  NAND2_X1 U9244 ( .A1(n7108), .A2(n14165), .ZN(n14040) );
  OAI21_X1 U9245 ( .B1(n14191), .B2(n14755), .A(n6702), .ZN(P1_U3527) );
  OR2_X1 U9246 ( .A1(n14111), .A2(n14728), .ZN(n6740) );
  NAND2_X1 U9247 ( .A1(n13931), .A2(n8040), .ZN(n13914) );
  OAI21_X1 U9248 ( .B1(n13992), .B2(n13995), .A(n8107), .ZN(n13977) );
  NAND3_X1 U9249 ( .A1(n6738), .A2(n14112), .A3(n6740), .ZN(n14198) );
  NAND2_X1 U9250 ( .A1(n6739), .A2(n14753), .ZN(n6738) );
  NAND2_X1 U9251 ( .A1(n8081), .A2(n8080), .ZN(n14672) );
  NAND2_X1 U9252 ( .A1(n7377), .A2(n7376), .ZN(n14008) );
  INV_X1 U9253 ( .A(n13977), .ZN(n7353) );
  NAND2_X1 U9254 ( .A1(n7019), .A2(n7020), .ZN(n8521) );
  INV_X1 U9255 ( .A(n8468), .ZN(n6710) );
  NAND2_X1 U9256 ( .A1(n8211), .A2(n8210), .ZN(n7027) );
  INV_X1 U9257 ( .A(n7011), .ZN(n7010) );
  NAND2_X1 U9258 ( .A1(n8815), .A2(n8812), .ZN(n6713) );
  NAND2_X2 U9259 ( .A1(n8227), .A2(n7079), .ZN(n6734) );
  NAND2_X1 U9260 ( .A1(n7046), .A2(n7044), .ZN(n11500) );
  NAND2_X1 U9261 ( .A1(n7034), .A2(n7038), .ZN(n14417) );
  INV_X1 U9262 ( .A(n14430), .ZN(n7047) );
  AND2_X2 U9263 ( .A1(n9517), .A2(n9516), .ZN(n12296) );
  NAND2_X2 U9264 ( .A1(n6720), .A2(n8294), .ZN(n12463) );
  NAND2_X1 U9265 ( .A1(n9552), .A2(n9553), .ZN(n9596) );
  NAND2_X1 U9266 ( .A1(n12410), .A2(n12288), .ZN(n12320) );
  NAND2_X1 U9267 ( .A1(n14958), .A2(n9549), .ZN(n14959) );
  OAI21_X1 U9268 ( .B1(n10954), .B2(n7050), .A(n6520), .ZN(n9540) );
  NOR2_X1 U9269 ( .A1(n12569), .A2(n6723), .ZN(n12256) );
  OAI21_X2 U9270 ( .B1(n12659), .B2(n7400), .A(n7397), .ZN(n12622) );
  AND2_X1 U9271 ( .A1(n15161), .A2(n15154), .ZN(n7395) );
  NOR2_X2 U9272 ( .A1(n14465), .A2(n12533), .ZN(n14482) );
  NAND2_X1 U9273 ( .A1(n6727), .A2(n6725), .ZN(P3_U3201) );
  NAND2_X1 U9274 ( .A1(n12537), .A2(n14480), .ZN(n6727) );
  AND2_X1 U9275 ( .A1(n7714), .A2(n7533), .ZN(n6804) );
  NAND2_X1 U9276 ( .A1(n6787), .A2(n6788), .ZN(n7937) );
  INV_X1 U9277 ( .A(n9491), .ZN(n9502) );
  NOR2_X1 U9278 ( .A1(n6987), .A2(n6986), .ZN(n6985) );
  INV_X1 U9279 ( .A(n9463), .ZN(n6991) );
  INV_X1 U9280 ( .A(n14113), .ZN(n6739) );
  INV_X1 U9281 ( .A(n7203), .ZN(n13270) );
  NAND2_X1 U9282 ( .A1(n8901), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8902) );
  OAI211_X1 U9283 ( .C1(n13441), .C2(n6813), .A(n6812), .B(n6817), .ZN(
        P2_U3496) );
  NAND2_X4 U9284 ( .A1(n14245), .A2(n14247), .ZN(n9755) );
  NAND2_X2 U9285 ( .A1(n7614), .A2(n7615), .ZN(n14247) );
  XNOR2_X1 U9286 ( .A(n13893), .B(n14193), .ZN(n13888) );
  INV_X1 U9287 ( .A(n7478), .ZN(n11934) );
  OR2_X2 U9288 ( .A1(n12576), .A2(n12585), .ZN(n8811) );
  XNOR2_X1 U9289 ( .A(n8846), .B(n12550), .ZN(n7026) );
  NAND2_X4 U9290 ( .A1(n12962), .A2(n9654), .ZN(n9652) );
  NAND2_X1 U9291 ( .A1(n12586), .A2(n6573), .ZN(n7098) );
  INV_X1 U9292 ( .A(n15186), .ZN(n12461) );
  NAND2_X1 U9293 ( .A1(n12745), .A2(n12744), .ZN(n12743) );
  NAND2_X1 U9294 ( .A1(n7144), .A2(n7142), .ZN(n13061) );
  INV_X1 U9295 ( .A(n6748), .ZN(n12950) );
  OAI21_X1 U9296 ( .B1(n6750), .B2(n6749), .A(n6578), .ZN(n8796) );
  NAND2_X1 U9297 ( .A1(n10459), .A2(n10433), .ZN(n10435) );
  NAND2_X1 U9298 ( .A1(n10475), .A2(n10432), .ZN(n10460) );
  XNOR2_X1 U9299 ( .A(n11090), .B(n11126), .ZN(n15012) );
  INV_X1 U9300 ( .A(n12493), .ZN(n6757) );
  NAND2_X1 U9301 ( .A1(n12466), .A2(n7220), .ZN(n7218) );
  NAND2_X1 U9302 ( .A1(n6893), .A2(n6488), .ZN(n6806) );
  INV_X8 U9303 ( .A(n9684), .ZN(n9685) );
  NAND2_X1 U9304 ( .A1(n8335), .A2(n8155), .ZN(n8351) );
  NOR2_X2 U9305 ( .A1(n11254), .A2(n11457), .ZN(n14527) );
  NOR2_X2 U9306 ( .A1(n13219), .A2(n12981), .ZN(n13430) );
  NAND2_X1 U9307 ( .A1(n14102), .A2(n6747), .ZN(P1_U3559) );
  AND2_X2 U9308 ( .A1(n11190), .A2(n14593), .ZN(n14402) );
  NAND2_X1 U9309 ( .A1(n14024), .A2(n14217), .ZN(n13996) );
  NAND2_X4 U9310 ( .A1(n9685), .A2(n9755), .ZN(n11750) );
  NOR2_X2 U9311 ( .A1(n8259), .A2(P3_IR_REG_29__SCAN_IN), .ZN(n6748) );
  AOI21_X2 U9312 ( .B1(n8820), .B2(n8845), .A(n8843), .ZN(n8847) );
  NAND2_X1 U9313 ( .A1(n14606), .A2(n6773), .ZN(n6772) );
  XNOR2_X1 U9314 ( .A(n7528), .B(SI_1_), .ZN(n7687) );
  OAI21_X1 U9315 ( .B1(n7538), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n6784), .ZN(
        n7528) );
  NAND2_X1 U9316 ( .A1(n7581), .A2(n6790), .ZN(n6787) );
  NAND2_X1 U9317 ( .A1(n7419), .A2(n7804), .ZN(n6793) );
  NAND2_X1 U9318 ( .A1(n7790), .A2(n7555), .ZN(n6794) );
  OR2_X2 U9319 ( .A1(n14114), .A2(n14700), .ZN(n6800) );
  NAND2_X2 U9320 ( .A1(n6802), .A2(n8028), .ZN(n13972) );
  NAND2_X1 U9321 ( .A1(n6803), .A2(n7537), .ZN(n7732) );
  NAND2_X1 U9322 ( .A1(n6804), .A2(n7534), .ZN(n6803) );
  NAND2_X1 U9323 ( .A1(n6809), .A2(n6819), .ZN(n13537) );
  OR2_X1 U9324 ( .A1(n14942), .A2(n6818), .ZN(n6817) );
  AND2_X2 U9325 ( .A1(n13440), .A2(n13439), .ZN(n6819) );
  NAND2_X1 U9326 ( .A1(n6822), .A2(n6820), .ZN(n7281) );
  NAND2_X1 U9327 ( .A1(n6830), .A2(n6826), .ZN(n10671) );
  INV_X1 U9328 ( .A(n6827), .ZN(n6826) );
  OAI21_X1 U9329 ( .B1(n6581), .B2(n10892), .A(n14847), .ZN(n6827) );
  OR2_X1 U9330 ( .A1(n10677), .A2(n13182), .ZN(n6831) );
  NAND2_X1 U9331 ( .A1(n6832), .A2(n6576), .ZN(n7238) );
  NAND2_X1 U9332 ( .A1(n12186), .A2(n12185), .ZN(n13423) );
  OR3_X2 U9333 ( .A1(n13358), .A2(n12196), .A3(n12193), .ZN(n6834) );
  AOI21_X1 U9334 ( .B1(n6843), .B2(n10672), .A(n6503), .ZN(n6842) );
  NAND2_X2 U9335 ( .A1(n11022), .A2(n11031), .ZN(n11243) );
  NAND2_X1 U9336 ( .A1(n6846), .A2(n7247), .ZN(n11021) );
  OAI21_X1 U9337 ( .B1(n11659), .B2(n6852), .A(n6850), .ZN(n13413) );
  NAND2_X1 U9338 ( .A1(n6856), .A2(n6855), .ZN(n8901) );
  NAND2_X1 U9339 ( .A1(n10803), .A2(n6863), .ZN(n6860) );
  NAND2_X1 U9340 ( .A1(n13399), .A2(n6874), .ZN(n6870) );
  NAND2_X1 U9341 ( .A1(n6870), .A2(n6867), .ZN(n6865) );
  NAND2_X1 U9342 ( .A1(n6865), .A2(n7266), .ZN(n13327) );
  CLKBUF_X1 U9343 ( .A(n6870), .Z(n6866) );
  MUX2_X1 U9344 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n9684), .Z(n7552) );
  NAND2_X1 U9345 ( .A1(n7833), .A2(n6880), .ZN(n6879) );
  NAND3_X1 U9346 ( .A1(n7282), .A2(n11914), .A3(n6906), .ZN(n11913) );
  AND2_X2 U9347 ( .A1(n6907), .A2(n7502), .ZN(n7476) );
  NOR2_X2 U9348 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n6907) );
  INV_X1 U9349 ( .A(n6908), .ZN(n7141) );
  OAI22_X1 U9350 ( .A1(n7707), .A2(n9760), .B1(n8053), .B2(n10595), .ZN(n6908)
         );
  NAND2_X4 U9351 ( .A1(n7512), .A2(n7511), .ZN(n8053) );
  NAND2_X2 U9352 ( .A1(n13721), .A2(n13722), .ZN(n13720) );
  NAND3_X1 U9353 ( .A1(n7289), .A2(n7503), .A3(n7292), .ZN(n8123) );
  NAND3_X1 U9354 ( .A1(n6911), .A2(n7315), .A3(n6916), .ZN(n6910) );
  NAND2_X1 U9355 ( .A1(n11349), .A2(n11350), .ZN(n6920) );
  OAI21_X1 U9356 ( .B1(n13689), .B2(n6924), .A(n6571), .ZN(n7329) );
  NAND2_X1 U9357 ( .A1(n11650), .A2(n6931), .ZN(n6930) );
  OR2_X1 U9358 ( .A1(n11835), .A2(n6946), .ZN(n6943) );
  NAND2_X1 U9359 ( .A1(n11835), .A2(n6511), .ZN(n6941) );
  NAND2_X1 U9360 ( .A1(n6950), .A2(n6951), .ZN(n11875) );
  NAND2_X1 U9361 ( .A1(n6954), .A2(n6957), .ZN(n11907) );
  NAND3_X1 U9362 ( .A1(n11887), .A2(n11886), .A3(n6961), .ZN(n6959) );
  NAND2_X1 U9363 ( .A1(n6959), .A2(n6960), .ZN(n11892) );
  INV_X1 U9364 ( .A(n11888), .ZN(n6962) );
  NAND2_X1 U9365 ( .A1(n7953), .A2(n6964), .ZN(n6966) );
  MUX2_X1 U9366 ( .A(n11804), .B(n13768), .S(n11771), .Z(n11805) );
  NAND2_X1 U9367 ( .A1(n9364), .A2(n6974), .ZN(n6972) );
  NAND2_X1 U9368 ( .A1(n6972), .A2(n6973), .ZN(n9409) );
  NAND2_X1 U9369 ( .A1(n6977), .A2(n6980), .ZN(n9260) );
  NAND2_X1 U9370 ( .A1(n6979), .A2(n6978), .ZN(n6977) );
  AOI21_X1 U9371 ( .B1(n6983), .B2(n7460), .A(n6981), .ZN(n6978) );
  NAND2_X1 U9372 ( .A1(n6984), .A2(n7458), .ZN(n6979) );
  NOR2_X1 U9373 ( .A1(n6982), .A2(n6525), .ZN(n6981) );
  INV_X1 U9374 ( .A(n9243), .ZN(n6982) );
  AND2_X1 U9375 ( .A1(n7461), .A2(n9230), .ZN(n6983) );
  AOI21_X1 U9376 ( .B1(n6994), .B2(n7467), .A(n6493), .ZN(n6992) );
  NAND2_X1 U9377 ( .A1(n9176), .A2(n6994), .ZN(n6993) );
  AOI21_X1 U9378 ( .B1(n7001), .B2(n6496), .A(n6580), .ZN(n6999) );
  NAND2_X1 U9379 ( .A1(n9317), .A2(n7001), .ZN(n7000) );
  NAND2_X1 U9380 ( .A1(n9158), .A2(n9159), .ZN(n9157) );
  XNOR2_X1 U9381 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8287) );
  NAND2_X1 U9382 ( .A1(n8571), .A2(n8196), .ZN(n7006) );
  INV_X1 U9383 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7009) );
  OAI21_X1 U9384 ( .B1(n8318), .B2(n7012), .A(n8332), .ZN(n7011) );
  NAND2_X1 U9385 ( .A1(n8429), .A2(n7016), .ZN(n7013) );
  NAND2_X1 U9386 ( .A1(n8488), .A2(n7022), .ZN(n7019) );
  NAND3_X1 U9387 ( .A1(n8696), .A2(n8695), .A3(n8684), .ZN(n7028) );
  NAND2_X1 U9388 ( .A1(n12383), .A2(n7029), .ZN(n12337) );
  NAND2_X1 U9389 ( .A1(n9524), .A2(n9521), .ZN(n7033) );
  NAND2_X1 U9390 ( .A1(n12271), .A2(n7035), .ZN(n7034) );
  NAND2_X1 U9391 ( .A1(n12418), .A2(n9543), .ZN(n7046) );
  NAND2_X1 U9392 ( .A1(n12346), .A2(n7053), .ZN(n7051) );
  OAI211_X1 U9393 ( .C1(n12346), .C2(n7056), .A(n7054), .B(n7051), .ZN(n12330)
         );
  NAND2_X1 U9394 ( .A1(n12346), .A2(n6514), .ZN(n7057) );
  AOI21_X1 U9395 ( .B1(n12346), .B2(n12347), .A(n7052), .ZN(n12427) );
  OAI21_X1 U9396 ( .B1(n7396), .B2(n7066), .A(n11326), .ZN(n15224) );
  NAND2_X1 U9397 ( .A1(n8327), .A2(n8727), .ZN(n7066) );
  NAND2_X1 U9398 ( .A1(n15153), .A2(n7071), .ZN(n7067) );
  AOI21_X1 U9399 ( .B1(n7071), .B2(n7073), .A(n7069), .ZN(n7068) );
  NAND2_X1 U9400 ( .A1(n8227), .A2(n7406), .ZN(n8853) );
  AND2_X1 U9401 ( .A1(n12586), .A2(n8813), .ZN(n12575) );
  NAND2_X1 U9402 ( .A1(n7103), .A2(n7102), .ZN(n7104) );
  AND2_X2 U9403 ( .A1(n7691), .A2(n7105), .ZN(n10131) );
  OR2_X2 U9404 ( .A1(n11470), .A2(n13738), .ZN(n11604) );
  NOR2_X2 U9405 ( .A1(n10995), .A2(n14747), .ZN(n11190) );
  NOR2_X2 U9406 ( .A1(n14040), .A2(n14220), .ZN(n14024) );
  OAI21_X1 U9407 ( .B1(n10991), .B2(n7114), .A(n7112), .ZN(n14392) );
  NAND2_X1 U9408 ( .A1(n7111), .A2(n7109), .ZN(n7861) );
  NAND2_X1 U9409 ( .A1(n10991), .A2(n7112), .ZN(n7111) );
  OAI21_X1 U9410 ( .B1(n10991), .B2(n11965), .A(n7831), .ZN(n11183) );
  INV_X1 U9411 ( .A(n11966), .ZN(n7116) );
  NAND2_X1 U9412 ( .A1(n14054), .A2(n7124), .ZN(n7123) );
  INV_X1 U9413 ( .A(n10581), .ZN(n7133) );
  NAND2_X1 U9414 ( .A1(n10581), .A2(n7131), .ZN(n7127) );
  NAND2_X1 U9415 ( .A1(n11611), .A2(n7138), .ZN(n7137) );
  OAI21_X1 U9416 ( .B1(n14644), .B2(n7773), .A(n7772), .ZN(n10581) );
  NAND2_X1 U9417 ( .A1(n11563), .A2(n11562), .ZN(n11561) );
  NAND2_X1 U9418 ( .A1(n11500), .A2(n9544), .ZN(n11563) );
  NAND2_X1 U9419 ( .A1(n14417), .A2(n12276), .ZN(n12436) );
  NAND2_X1 U9420 ( .A1(n7713), .A2(n11784), .ZN(n10533) );
  NAND2_X1 U9421 ( .A1(n11326), .A2(n8341), .ZN(n15153) );
  NAND2_X1 U9422 ( .A1(n8613), .A2(n8791), .ZN(n12639) );
  OR2_X1 U9423 ( .A1(n9107), .A2(n9106), .ZN(n9122) );
  OR2_X1 U9424 ( .A1(n9349), .A2(n9348), .ZN(n9364) );
  NAND2_X1 U9425 ( .A1(n7457), .A2(n6532), .ZN(n7456) );
  OAI21_X1 U9426 ( .B1(n9491), .B2(n14864), .A(n9490), .ZN(n9505) );
  NAND2_X1 U9427 ( .A1(n9296), .A2(n6533), .ZN(n9317) );
  NAND2_X1 U9428 ( .A1(n15178), .A2(n12296), .ZN(n9520) );
  AND2_X4 U9429 ( .A1(n7700), .A2(n7491), .ZN(n7734) );
  OR2_X2 U9430 ( .A1(n14682), .A2(n13771), .ZN(n11784) );
  OR2_X1 U9431 ( .A1(n7673), .A2(n7672), .ZN(n7674) );
  NAND2_X1 U9432 ( .A1(n13103), .A2(n13102), .ZN(n7144) );
  OAI21_X2 U9433 ( .B1(n13018), .B2(n13017), .A(n7145), .ZN(n13103) );
  NAND2_X1 U9434 ( .A1(n13000), .A2(n13001), .ZN(n7145) );
  NAND2_X1 U9435 ( .A1(n13070), .A2(n7153), .ZN(n7150) );
  CLKBUF_X1 U9436 ( .A(n7150), .Z(n7146) );
  NAND2_X1 U9437 ( .A1(n13070), .A2(n13069), .ZN(n13068) );
  AND2_X1 U9438 ( .A1(n7159), .A2(n7158), .ZN(n7157) );
  NAND2_X1 U9439 ( .A1(n11700), .A2(n7170), .ZN(n7169) );
  NAND2_X1 U9440 ( .A1(n7169), .A2(n7166), .ZN(n12974) );
  NAND2_X1 U9441 ( .A1(n11700), .A2(n7172), .ZN(n11703) );
  INV_X1 U9442 ( .A(n7169), .ZN(n11726) );
  NOR2_X1 U9443 ( .A1(n11704), .A2(n7171), .ZN(n7170) );
  INV_X1 U9444 ( .A(n7172), .ZN(n7171) );
  NAND2_X1 U9445 ( .A1(n13141), .A2(n7174), .ZN(n7173) );
  OAI211_X1 U9446 ( .C1(n13141), .C2(n7178), .A(n7175), .B(n7173), .ZN(n13043)
         );
  OR2_X2 U9447 ( .A1(n13141), .A2(n13140), .ZN(n13138) );
  NOR2_X1 U9448 ( .A1(n10410), .A2(n10409), .ZN(n10570) );
  INV_X1 U9449 ( .A(n10569), .ZN(n7191) );
  NAND2_X1 U9450 ( .A1(n10567), .A2(n10568), .ZN(n7192) );
  AOI21_X1 U9451 ( .B1(n10179), .B2(n13213), .A(n8924), .ZN(n7193) );
  NAND2_X1 U9452 ( .A1(n10180), .A2(n13213), .ZN(n7194) );
  OAI21_X1 U9453 ( .B1(n10180), .B2(n10179), .A(n13213), .ZN(n14925) );
  INV_X1 U9454 ( .A(n9437), .ZN(n7199) );
  NAND2_X2 U9455 ( .A1(n7208), .A2(n7207), .ZN(n13374) );
  NOR2_X2 U9456 ( .A1(n14464), .A2(n8547), .ZN(n14465) );
  NAND2_X1 U9457 ( .A1(n7238), .A2(n7239), .ZN(n13380) );
  NAND2_X1 U9458 ( .A1(n7244), .A2(n10668), .ZN(n10825) );
  NAND2_X1 U9459 ( .A1(n10892), .A2(n10893), .ZN(n7244) );
  OAI21_X1 U9460 ( .B1(n10893), .B2(n7246), .A(n10685), .ZN(n7245) );
  NAND2_X1 U9461 ( .A1(n10717), .A2(n10716), .ZN(n10719) );
  NAND2_X1 U9462 ( .A1(n11243), .A2(n7277), .ZN(n11450) );
  OAI21_X2 U9463 ( .B1(n13310), .B2(n12161), .A(n12163), .ZN(n13302) );
  NAND2_X1 U9464 ( .A1(n10671), .A2(n10670), .ZN(n10798) );
  OAI21_X2 U9465 ( .B1(n11541), .B2(n11540), .A(n11542), .ZN(n11667) );
  NAND2_X1 U9466 ( .A1(n7288), .A2(n11982), .ZN(n11952) );
  AND2_X2 U9467 ( .A1(n7290), .A2(n7734), .ZN(n7289) );
  AND2_X2 U9468 ( .A1(n7476), .A2(n7291), .ZN(n7290) );
  AND2_X2 U9469 ( .A1(n7498), .A2(n7497), .ZN(n7292) );
  NAND2_X1 U9470 ( .A1(n11856), .A2(n7490), .ZN(n7296) );
  NAND2_X1 U9471 ( .A1(n11844), .A2(n11843), .ZN(n7294) );
  NAND3_X1 U9472 ( .A1(n7296), .A2(n7295), .A3(n11861), .ZN(n11865) );
  NAND2_X1 U9473 ( .A1(n11810), .A2(n11811), .ZN(n11809) );
  OAI22_X1 U9474 ( .A1(n11831), .A2(n7298), .B1(n11832), .B2(n7297), .ZN(
        n11835) );
  NAND2_X1 U9475 ( .A1(n11823), .A2(n11824), .ZN(n11822) );
  INV_X2 U9476 ( .A(n11750), .ZN(n11935) );
  NAND2_X1 U9477 ( .A1(n13720), .A2(n7307), .ZN(n7306) );
  OAI211_X1 U9478 ( .C1(n13720), .C2(n7311), .A(n7309), .B(n7306), .ZN(n12145)
         );
  NAND2_X1 U9479 ( .A1(n7475), .A2(n7326), .ZN(n7318) );
  INV_X1 U9480 ( .A(n11159), .ZN(n7326) );
  NAND2_X1 U9481 ( .A1(n7953), .A2(n7342), .ZN(n8062) );
  NOR2_X4 U9482 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n7700) );
  NAND2_X1 U9483 ( .A1(n11006), .A2(n7349), .ZN(n7347) );
  NAND2_X1 U9484 ( .A1(n14081), .A2(n7361), .ZN(n7360) );
  NAND2_X1 U9485 ( .A1(n11569), .A2(n7366), .ZN(n7365) );
  NAND2_X1 U9486 ( .A1(n14038), .A2(n7378), .ZN(n7377) );
  NAND2_X2 U9487 ( .A1(n8826), .A2(n9518), .ZN(n10936) );
  NAND2_X2 U9488 ( .A1(n12463), .A2(n10738), .ZN(n8826) );
  NAND2_X1 U9489 ( .A1(n7381), .A2(n7380), .ZN(n12236) );
  NAND2_X1 U9490 ( .A1(n12234), .A2(n6572), .ZN(n7381) );
  NAND3_X1 U9491 ( .A1(n6539), .A2(n15123), .A3(n15159), .ZN(n12224) );
  OR2_X2 U9492 ( .A1(n11047), .A2(n11046), .ZN(n15155) );
  INV_X1 U9493 ( .A(n12213), .ZN(n7396) );
  AND2_X2 U9494 ( .A1(n8354), .A2(n8221), .ZN(n8412) );
  NAND2_X1 U9495 ( .A1(n12582), .A2(n12255), .ZN(n12566) );
  NAND2_X1 U9496 ( .A1(n12683), .A2(n12689), .ZN(n12245) );
  INV_X1 U9497 ( .A(n8234), .ZN(n8235) );
  OAI21_X1 U9498 ( .B1(n7538), .B2(n9691), .A(n7416), .ZN(n7697) );
  INV_X1 U9499 ( .A(n7538), .ZN(n8014) );
  MUX2_X1 U9500 ( .A(n9698), .B(n9683), .S(n7417), .Z(n7543) );
  INV_X1 U9501 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7418) );
  NAND2_X1 U9502 ( .A1(n8044), .A2(n7426), .ZN(n7423) );
  NAND2_X1 U9503 ( .A1(n7430), .A2(n7429), .ZN(n7581) );
  NAND2_X1 U9504 ( .A1(n8000), .A2(n7596), .ZN(n7431) );
  OAI211_X1 U9505 ( .C1(n8000), .C2(n7435), .A(n7434), .B(n7432), .ZN(n9302)
         );
  INV_X1 U9506 ( .A(SI_22_), .ZN(n7435) );
  NAND2_X1 U9507 ( .A1(n7453), .A2(n7448), .ZN(n7633) );
  INV_X1 U9508 ( .A(n9141), .ZN(n7454) );
  INV_X1 U9509 ( .A(n9140), .ZN(n7455) );
  INV_X1 U9510 ( .A(n9120), .ZN(n7457) );
  NAND2_X1 U9511 ( .A1(n9210), .A2(n9229), .ZN(n7458) );
  NAND2_X1 U9512 ( .A1(n9211), .A2(n9229), .ZN(n7459) );
  INV_X1 U9513 ( .A(n9210), .ZN(n7460) );
  NAND2_X1 U9514 ( .A1(n9411), .A2(n9410), .ZN(n7465) );
  INV_X1 U9515 ( .A(n9378), .ZN(n7466) );
  NAND2_X1 U9516 ( .A1(n7471), .A2(n7472), .ZN(n9295) );
  NAND3_X1 U9517 ( .A1(n9263), .A2(n9262), .A3(n6569), .ZN(n7471) );
  INV_X1 U9518 ( .A(n9069), .ZN(n7473) );
  INV_X1 U9519 ( .A(n9068), .ZN(n7474) );
  NAND2_X1 U9520 ( .A1(n11770), .A2(n11769), .ZN(n11772) );
  INV_X1 U9521 ( .A(n13972), .ZN(n14208) );
  INV_X1 U9522 ( .A(n10953), .ZN(n9530) );
  NAND2_X1 U9523 ( .A1(n9518), .A2(n12328), .ZN(n9519) );
  XNOR2_X1 U9524 ( .A(n9613), .B(n12132), .ZN(n9616) );
  NAND2_X1 U9525 ( .A1(n8862), .A2(n8861), .ZN(P3_U3296) );
  AND2_X2 U9526 ( .A1(n13975), .A2(n8108), .ZN(n13961) );
  INV_X1 U9527 ( .A(n7953), .ZN(n7939) );
  OR2_X1 U9528 ( .A1(n8239), .A2(n6724), .ZN(n8241) );
  NOR2_X1 U9529 ( .A1(n11918), .A2(n11917), .ZN(n11919) );
  OR2_X2 U9530 ( .A1(n10131), .A2(n13772), .ZN(n11774) );
  AOI222_X1 U9531 ( .A1(n14850), .A2(n14846), .B1(P2_REG2_REG_4__SCAN_IN), 
        .B2(n14873), .C1(n14845), .C2(n14844), .ZN(n14857) );
  AND2_X2 U9532 ( .A1(n8932), .A2(n8870), .ZN(n8946) );
  INV_X1 U9533 ( .A(n10900), .ZN(n14903) );
  NAND2_X1 U9534 ( .A1(n8965), .A2(n10900), .ZN(n8951) );
  AOI22_X1 U9535 ( .A1(n8965), .A2(n13181), .B1(n9118), .B2(n10900), .ZN(n8956) );
  AOI22_X1 U9536 ( .A1(n9067), .A2(n13182), .B1(n9118), .B2(n10677), .ZN(n8952) );
  NAND2_X1 U9537 ( .A1(n8930), .A2(n8929), .ZN(n8954) );
  OAI21_X1 U9538 ( .B1(n13075), .B2(n9406), .A(n9227), .ZN(n9228) );
  NAND2_X1 U9539 ( .A1(n13181), .A2(n9406), .ZN(n8950) );
  AND2_X2 U9540 ( .A1(n12947), .A2(n9608), .ZN(P3_U3897) );
  OR2_X1 U9541 ( .A1(n7885), .A2(SI_14_), .ZN(n7477) );
  AND2_X1 U9542 ( .A1(n11855), .A2(n11854), .ZN(n7479) );
  AND3_X1 U9543 ( .A1(n8905), .A2(n8876), .A3(n8875), .ZN(n7480) );
  AND2_X1 U9544 ( .A1(n7586), .A2(n7585), .ZN(n7481) );
  AND2_X1 U9545 ( .A1(n7574), .A2(n7573), .ZN(n7482) );
  AND2_X1 U9546 ( .A1(n10218), .A2(n9499), .ZN(n13142) );
  INV_X1 U9547 ( .A(n13142), .ZN(n13072) );
  AND2_X1 U9548 ( .A1(n9401), .A2(n9400), .ZN(n13011) );
  INV_X2 U9549 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U9550 ( .A1(n14424), .A2(n12274), .ZN(n7483) );
  INV_X1 U9551 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14234) );
  AND2_X1 U9552 ( .A1(n14871), .A2(n13213), .ZN(n14854) );
  AND2_X1 U9553 ( .A1(n9437), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7484) );
  NAND2_X1 U9554 ( .A1(n13903), .A2(n14667), .ZN(n14389) );
  AND2_X1 U9555 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7485) );
  INV_X1 U9556 ( .A(n10130), .ZN(n7679) );
  AND2_X1 U9557 ( .A1(n7570), .A2(n7569), .ZN(n7486) );
  NOR2_X1 U9558 ( .A1(n7483), .A2(n12767), .ZN(n7487) );
  NOR2_X1 U9559 ( .A1(n12763), .A2(n7483), .ZN(n7488) );
  NOR2_X1 U9560 ( .A1(n8766), .A2(n8767), .ZN(n7489) );
  INV_X2 U9561 ( .A(n14940), .ZN(n14942) );
  CLKBUF_X2 U9562 ( .A(P1_U4016), .Z(n13788) );
  NAND2_X1 U9563 ( .A1(n8965), .A2(n14909), .ZN(n8971) );
  AOI22_X1 U9564 ( .A1(n8965), .A2(n13180), .B1(n9118), .B2(n14909), .ZN(n8988) );
  NAND2_X1 U9565 ( .A1(n8956), .A2(n8955), .ZN(n8973) );
  OAI21_X1 U9566 ( .B1(n14917), .B2(n9406), .A(n8986), .ZN(n8994) );
  NAND2_X1 U9567 ( .A1(n11777), .A2(n11776), .ZN(n11782) );
  NAND2_X1 U9568 ( .A1(n11826), .A2(n11825), .ZN(n11827) );
  INV_X1 U9569 ( .A(n9159), .ZN(n9160) );
  INV_X1 U9570 ( .A(n9229), .ZN(n9230) );
  NAND2_X1 U9571 ( .A1(n11899), .A2(n11898), .ZN(n11900) );
  OAI21_X1 U9572 ( .B1(n12166), .B2(n9449), .A(n9362), .ZN(n9363) );
  INV_X1 U9573 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8875) );
  INV_X1 U9574 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8222) );
  INV_X1 U9575 ( .A(n8605), .ZN(n8251) );
  INV_X1 U9576 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8228) );
  AND4_X1 U9577 ( .A1(n10376), .A2(n8220), .A3(n8385), .A4(n8219), .ZN(n8221)
         );
  INV_X1 U9578 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8880) );
  INV_X1 U9579 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8906) );
  INV_X1 U9580 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7523) );
  NAND2_X1 U9581 ( .A1(n8251), .A2(n8250), .ZN(n8618) );
  INV_X1 U9582 ( .A(n12852), .ZN(n12811) );
  AND4_X1 U9583 ( .A1(n8230), .A2(n8229), .A3(n8228), .A4(n8711), .ZN(n8231)
         );
  INV_X1 U9584 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9058) );
  INV_X1 U9585 ( .A(P2_B_REG_SCAN_IN), .ZN(n12174) );
  INV_X1 U9586 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8870) );
  AND2_X1 U9587 ( .A1(n10761), .A2(n10760), .ZN(n10762) );
  INV_X1 U9588 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7795) );
  INV_X1 U9589 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7852) );
  INV_X1 U9590 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7499) );
  INV_X1 U9591 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14269) );
  INV_X1 U9592 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8477) );
  INV_X1 U9593 ( .A(n14968), .ZN(n14420) );
  OR2_X1 U9594 ( .A1(n8661), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8674) );
  INV_X1 U9595 ( .A(n8806), .ZN(n8668) );
  INV_X1 U9596 ( .A(n10563), .ZN(n10638) );
  INV_X1 U9597 ( .A(n12948), .ZN(n10862) );
  INV_X1 U9598 ( .A(n12217), .ZN(n15161) );
  INV_X1 U9599 ( .A(n10730), .ZN(n12810) );
  OR2_X1 U9600 ( .A1(n8461), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n8471) );
  NOR2_X1 U9601 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8217) );
  INV_X1 U9602 ( .A(n12983), .ZN(n12984) );
  OR2_X1 U9603 ( .A1(n9369), .A2(n9368), .ZN(n9392) );
  INV_X1 U9604 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9236) );
  AND2_X1 U9605 ( .A1(n8921), .A2(n9442), .ZN(n10218) );
  AND2_X1 U9606 ( .A1(n8923), .A2(n8922), .ZN(n9468) );
  INV_X1 U9607 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9000) );
  INV_X1 U9608 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7872) );
  AND2_X1 U9609 ( .A1(n11646), .A2(n11645), .ZN(n11647) );
  INV_X1 U9610 ( .A(n7665), .ZN(n7652) );
  OR2_X1 U9611 ( .A1(n7974), .A2(n7973), .ZN(n7987) );
  AND2_X1 U9612 ( .A1(n10917), .A2(n10916), .ZN(n10919) );
  OR2_X1 U9613 ( .A1(n7927), .A2(n10912), .ZN(n7943) );
  INV_X1 U9614 ( .A(n13711), .ZN(n13725) );
  OR2_X1 U9615 ( .A1(n9735), .A2(P1_D_REG_1__SCAN_IN), .ZN(n8144) );
  INV_X1 U9616 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7504) );
  INV_X1 U9617 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n7491) );
  INV_X1 U9618 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14283) );
  INV_X1 U9619 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14343) );
  INV_X1 U9620 ( .A(n10952), .ZN(n9529) );
  OR2_X1 U9621 ( .A1(n8687), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8689) );
  NAND2_X1 U9622 ( .A1(n9520), .A2(n9519), .ZN(n9525) );
  NAND2_X1 U9623 ( .A1(n14420), .A2(n15145), .ZN(n12414) );
  AND2_X1 U9624 ( .A1(n10563), .A2(n12523), .ZN(n10937) );
  INV_X1 U9625 ( .A(n8689), .ZN(n12262) );
  INV_X1 U9626 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14291) );
  AND2_X1 U9627 ( .A1(n9664), .A2(n9653), .ZN(n9660) );
  AND2_X1 U9628 ( .A1(n8704), .A2(n8267), .ZN(n12259) );
  INV_X1 U9629 ( .A(n12713), .ZN(n12718) );
  OR2_X1 U9630 ( .A1(n9766), .A2(n9569), .ZN(n10632) );
  NAND2_X1 U9631 ( .A1(n12891), .A2(n15253), .ZN(n12893) );
  NAND2_X1 U9632 ( .A1(n14490), .A2(n8758), .ZN(n12793) );
  AND2_X1 U9633 ( .A1(n8749), .A2(n8750), .ZN(n15110) );
  AND2_X1 U9634 ( .A1(n15169), .A2(n12838), .ZN(n12852) );
  NAND2_X1 U9635 ( .A1(n12810), .A2(n10614), .ZN(n15219) );
  INV_X1 U9636 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8849) );
  AND2_X1 U9637 ( .A1(n8196), .A2(n8195), .ZN(n8568) );
  AND2_X1 U9638 ( .A1(n8183), .A2(n8182), .ZN(n8487) );
  INV_X1 U9639 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n11301) );
  NAND2_X1 U9640 ( .A1(n12982), .A2(n12984), .ZN(n12985) );
  NOR2_X1 U9641 ( .A1(n10209), .A2(n14883), .ZN(n10215) );
  OR2_X1 U9642 ( .A1(n13239), .A2(n9395), .ZN(n9401) );
  OR2_X1 U9643 ( .A1(n9237), .A2(n9236), .ZN(n9249) );
  INV_X1 U9644 ( .A(n9837), .ZN(n9855) );
  INV_X1 U9645 ( .A(n12189), .ZN(n13387) );
  AND2_X1 U9646 ( .A1(n10206), .A2(n9468), .ZN(n10208) );
  OR2_X1 U9647 ( .A1(n14859), .A2(n8923), .ZN(n10205) );
  INV_X1 U9648 ( .A(n14860), .ZN(n13368) );
  INV_X1 U9649 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8910) );
  INV_X1 U9650 ( .A(n13764), .ZN(n11398) );
  INV_X1 U9651 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n10912) );
  INV_X1 U9652 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13691) );
  INV_X1 U9653 ( .A(n8053), .ZN(n8022) );
  INV_X1 U9654 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9790) );
  INV_X1 U9655 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n13671) );
  NAND2_X1 U9656 ( .A1(n14264), .A2(n8113), .ZN(n11941) );
  INV_X1 U9657 ( .A(n13745), .ZN(n12134) );
  AND2_X1 U9658 ( .A1(n7947), .A2(n6553), .ZN(n14091) );
  INV_X1 U9659 ( .A(n11958), .ZN(n10513) );
  INV_X1 U9660 ( .A(n14686), .ZN(n14090) );
  AND2_X1 U9661 ( .A1(n8126), .A2(n9736), .ZN(n9643) );
  INV_X1 U9662 ( .A(n14674), .ZN(n14655) );
  NAND2_X2 U9663 ( .A1(n10028), .A2(n11938), .ZN(n14674) );
  OR2_X1 U9664 ( .A1(n14674), .A2(n14564), .ZN(n9639) );
  OAI22_X1 U9665 ( .A1(n14319), .A2(n14276), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n15010), .ZN(n14277) );
  AOI22_X1 U9666 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14289), .B1(n14292), 
        .B2(n14288), .ZN(n14345) );
  OR2_X1 U9667 ( .A1(n10866), .A2(n8851), .ZN(n9664) );
  OR2_X1 U9668 ( .A1(n8499), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8513) );
  NAND2_X1 U9669 ( .A1(n10630), .A2(n10632), .ZN(n10611) );
  INV_X1 U9670 ( .A(n10886), .ZN(n8851) );
  OR2_X1 U9671 ( .A1(n14460), .A2(n14459), .ZN(n14461) );
  MUX2_X1 U9672 ( .A(n9660), .B(P3_U3897), .S(n12257), .Z(n15056) );
  INV_X1 U9673 ( .A(n15187), .ZN(n15145) );
  INV_X1 U9674 ( .A(n12805), .ZN(n15086) );
  NOR2_X1 U9675 ( .A1(n10869), .A2(n15199), .ZN(n15173) );
  AND2_X1 U9676 ( .A1(n10642), .A2(n10641), .ZN(n10643) );
  INV_X1 U9677 ( .A(n12838), .ZN(n15243) );
  AND2_X1 U9678 ( .A1(n15253), .A2(n15242), .ZN(n12910) );
  INV_X1 U9679 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8716) );
  INV_X1 U9680 ( .A(n11139), .ZN(n15057) );
  INV_X1 U9681 ( .A(n11115), .ZN(n14987) );
  INV_X1 U9682 ( .A(n13097), .ZN(n13147) );
  INV_X1 U9683 ( .A(n13137), .ZN(n13149) );
  INV_X1 U9684 ( .A(n9006), .ZN(n9395) );
  AND2_X1 U9685 ( .A1(n9855), .A2(n10217), .ZN(n14798) );
  INV_X1 U9686 ( .A(n14803), .ZN(n14811) );
  NAND2_X1 U9687 ( .A1(n9855), .A2(n9854), .ZN(n14803) );
  AND2_X1 U9688 ( .A1(n9855), .A2(n9839), .ZN(n14820) );
  INV_X1 U9689 ( .A(n13486), .ZN(n13497) );
  NAND2_X1 U9690 ( .A1(n10205), .A2(n10203), .ZN(n14933) );
  AND2_X1 U9691 ( .A1(n14925), .A2(n10666), .ZN(n14938) );
  INV_X1 U9692 ( .A(n14938), .ZN(n14921) );
  OR2_X1 U9693 ( .A1(n10770), .A2(n10705), .ZN(n11338) );
  INV_X1 U9694 ( .A(n13593), .ZN(n10200) );
  NOR2_X1 U9695 ( .A1(n9685), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13585) );
  AND2_X1 U9696 ( .A1(n7892), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7913) );
  AND2_X1 U9697 ( .A1(n10026), .A2(n10516), .ZN(n14552) );
  INV_X1 U9698 ( .A(n14557), .ZN(n13734) );
  NAND2_X1 U9699 ( .A1(n9626), .A2(n9791), .ZN(n13711) );
  AND2_X1 U9700 ( .A1(n7980), .A2(n7979), .ZN(n13714) );
  AND3_X1 U9701 ( .A1(n7962), .A2(n7961), .A3(n7960), .ZN(n13668) );
  INV_X1 U9702 ( .A(n14245), .ZN(n9791) );
  OR2_X1 U9703 ( .A1(n9792), .A2(n9786), .ZN(n14627) );
  INV_X1 U9704 ( .A(n14636), .ZN(n13855) );
  AND2_X1 U9705 ( .A1(n9763), .A2(n14247), .ZN(n14631) );
  NAND2_X1 U9706 ( .A1(n11939), .A2(n11984), .ZN(n14560) );
  INV_X1 U9707 ( .A(n11978), .ZN(n13932) );
  INV_X1 U9708 ( .A(n14407), .ZN(n14399) );
  INV_X1 U9709 ( .A(n14050), .ZN(n14055) );
  AND3_X1 U9710 ( .A1(n9644), .A2(n9643), .A3(n9642), .ZN(n10026) );
  AND3_X1 U9711 ( .A1(n14188), .A2(n14187), .A3(n14186), .ZN(n14230) );
  AND2_X1 U9712 ( .A1(n11571), .A2(n11570), .ZN(n14566) );
  INV_X1 U9713 ( .A(n14700), .ZN(n14732) );
  NAND2_X1 U9714 ( .A1(n14700), .A2(n14721), .ZN(n14753) );
  INV_X1 U9715 ( .A(n14721), .ZN(n14745) );
  AND2_X1 U9716 ( .A1(n9634), .A2(n9738), .ZN(n9753) );
  INV_X1 U9717 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7611) );
  INV_X1 U9718 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8066) );
  AND2_X1 U9719 ( .A1(n7810), .A2(n7822), .ZN(n9900) );
  NOR2_X1 U9720 ( .A1(n9685), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14235) );
  AND2_X1 U9721 ( .A1(n9664), .A2(n9663), .ZN(n15025) );
  OR2_X1 U9722 ( .A1(n10611), .A2(n9588), .ZN(n14968) );
  INV_X1 U9723 ( .A(n14960), .ZN(n12433) );
  INV_X1 U9724 ( .A(n12598), .ZN(n12571) );
  OAI211_X1 U9725 ( .C1(n6473), .C2(n12913), .A(n8631), .B(n8630), .ZN(n12449)
         );
  INV_X1 U9726 ( .A(n12439), .ZN(n12751) );
  INV_X1 U9727 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n14990) );
  INV_X1 U9728 ( .A(n15025), .ZN(n15074) );
  NAND2_X1 U9729 ( .A1(P3_U3897), .A2(n12962), .ZN(n15067) );
  AND2_X1 U9730 ( .A1(n12625), .A2(n12624), .ZN(n12835) );
  NAND2_X1 U9731 ( .A1(n15204), .A2(n15148), .ZN(n12805) );
  AND2_X1 U9732 ( .A1(n15080), .A2(n15079), .ZN(n15248) );
  OR2_X1 U9733 ( .A1(n10859), .A2(n10643), .ZN(n15270) );
  INV_X1 U9734 ( .A(n12558), .ZN(n12887) );
  INV_X1 U9735 ( .A(n12694), .ZN(n12927) );
  AND2_X2 U9736 ( .A1(n10612), .A2(n10866), .ZN(n15253) );
  NAND2_X1 U9737 ( .A1(n12947), .A2(n9766), .ZN(n9767) );
  INV_X1 U9738 ( .A(n12964), .ZN(n10884) );
  INV_X1 U9739 ( .A(n12528), .ZN(n12540) );
  INV_X1 U9740 ( .A(n15043), .ZN(n11133) );
  INV_X1 U9741 ( .A(n14522), .ZN(n14537) );
  INV_X1 U9742 ( .A(n11696), .ZN(n11712) );
  INV_X1 U9743 ( .A(n13129), .ZN(n13151) );
  INV_X1 U9744 ( .A(n13011), .ZN(n13155) );
  INV_X1 U9745 ( .A(n14818), .ZN(n11524) );
  INV_X1 U9746 ( .A(n14854), .ZN(n14833) );
  NAND2_X1 U9747 ( .A1(n14535), .A2(n14933), .ZN(n13486) );
  OR2_X1 U9748 ( .A1(n11338), .A2(n10706), .ZN(n14940) );
  INV_X1 U9749 ( .A(n14886), .ZN(n14883) );
  NOR2_X1 U9750 ( .A1(n14874), .A2(n14883), .ZN(n14882) );
  INV_X1 U9751 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10237) );
  INV_X1 U9752 ( .A(n11820), .ZN(n14735) );
  NAND2_X1 U9753 ( .A1(n10035), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14557) );
  INV_X1 U9754 ( .A(n11837), .ZN(n14593) );
  INV_X1 U9755 ( .A(n14554), .ZN(n13730) );
  OAI21_X1 U9756 ( .B1(n14044), .B2(n8053), .A(n7994), .ZN(n13753) );
  INV_X1 U9757 ( .A(n11841), .ZN(n13761) );
  INV_X1 U9758 ( .A(n14631), .ZN(n13860) );
  INV_X1 U9759 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14641) );
  OR2_X1 U9760 ( .A1(n6476), .A2(n14560), .ZN(n14683) );
  OR2_X1 U9761 ( .A1(n6476), .A2(n11942), .ZN(n13988) );
  OR2_X1 U9762 ( .A1(n6476), .A2(n14728), .ZN(n14050) );
  OR2_X1 U9763 ( .A1(n6476), .A2(n10527), .ZN(n14077) );
  NAND2_X1 U9764 ( .A1(n14766), .A2(n14724), .ZN(n14190) );
  AND2_X2 U9765 ( .A1(n10026), .A2(n10025), .ZN(n14766) );
  INV_X1 U9766 ( .A(n13915), .ZN(n14199) );
  INV_X1 U9767 ( .A(n13621), .ZN(n14227) );
  INV_X1 U9768 ( .A(n14756), .ZN(n14755) );
  INV_X1 U9769 ( .A(n9747), .ZN(n9738) );
  INV_X1 U9770 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14246) );
  INV_X1 U9771 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10506) );
  INV_X1 U9772 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9919) );
  NAND2_X1 U9773 ( .A1(n9685), .A2(P1_U3086), .ZN(n14258) );
  OR4_X1 U9774 ( .A1(n9606), .A2(n9605), .A3(n9604), .A4(n9603), .ZN(P3_U3164)
         );
  OR4_X1 U9775 ( .A1(n9595), .A2(n9594), .A3(n9593), .A4(n9592), .ZN(P3_U3176)
         );
  NOR2_X1 U9776 ( .A1(P2_U3088), .A2(n9836), .ZN(P2_U3947) );
  NOR2_X1 U9777 ( .A1(n9634), .A2(n9747), .ZN(P1_U4016) );
  NOR2_X1 U9778 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n7495) );
  NOR2_X1 U9779 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n7494) );
  NOR2_X1 U9780 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n7493) );
  AND4_X2 U9781 ( .A1(n7495), .A2(n7494), .A3(n7493), .A4(n7492), .ZN(n7498)
         );
  AND4_X2 U9782 ( .A1(n7907), .A2(n7496), .A3(n7733), .A4(n7745), .ZN(n7497)
         );
  NOR2_X1 U9783 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n7501) );
  NAND4_X1 U9784 ( .A1(n8060), .A2(n7501), .A3(n7500), .A4(n7499), .ZN(n8116)
         );
  INV_X1 U9785 ( .A(n8116), .ZN(n7503) );
  NAND2_X1 U9786 ( .A1(n7506), .A2(n7508), .ZN(n14240) );
  XNOR2_X2 U9787 ( .A(n7505), .B(P1_IR_REG_30__SCAN_IN), .ZN(n7511) );
  NAND2_X1 U9788 ( .A1(n11760), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n7522) );
  AND2_X4 U9789 ( .A1(n12000), .A2(n14242), .ZN(n8049) );
  INV_X1 U9790 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n7510) );
  OR2_X1 U9791 ( .A1(n7992), .A2(n7510), .ZN(n7521) );
  NAND2_X1 U9792 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n7751) );
  INV_X1 U9793 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7750) );
  NOR2_X1 U9794 ( .A1(n7751), .A2(n7750), .ZN(n7765) );
  NAND2_X1 U9795 ( .A1(n7765), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7782) );
  INV_X1 U9796 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7781) );
  AND2_X1 U9797 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n7513) );
  NAND2_X1 U9798 ( .A1(n7839), .A2(n7513), .ZN(n7853) );
  NAND2_X1 U9799 ( .A1(n7913), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7927) );
  NAND2_X1 U9800 ( .A1(n7957), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7974) );
  INV_X1 U9801 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7973) );
  INV_X1 U9802 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8004) );
  NAND2_X1 U9803 ( .A1(n8016), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8017) );
  INV_X1 U9804 ( .A(n8017), .ZN(n7666) );
  NAND2_X1 U9805 ( .A1(n7666), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7665) );
  NAND2_X1 U9806 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n7652), .ZN(n8030) );
  INV_X1 U9807 ( .A(n8030), .ZN(n7514) );
  NAND2_X1 U9808 ( .A1(n7514), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8032) );
  INV_X1 U9809 ( .A(n8032), .ZN(n7515) );
  NAND2_X1 U9810 ( .A1(n7515), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n7638) );
  INV_X1 U9811 ( .A(n7638), .ZN(n7516) );
  NAND2_X1 U9812 ( .A1(n7516), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8051) );
  INV_X1 U9813 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7517) );
  XNOR2_X1 U9814 ( .A(n8051), .B(n7517), .ZN(n13918) );
  OR2_X1 U9815 ( .A1(n8053), .A2(n13918), .ZN(n7520) );
  INV_X1 U9816 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n7518) );
  OR2_X1 U9817 ( .A1(n8034), .A2(n7518), .ZN(n7519) );
  NAND4_X1 U9818 ( .A1(n7522), .A2(n7521), .A3(n7520), .A4(n7519), .ZN(n13745)
         );
  INV_X1 U9819 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9693) );
  INV_X1 U9820 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8147) );
  NAND3_X1 U9821 ( .A1(n7524), .A2(n7523), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7525) );
  AND2_X1 U9822 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n7526) );
  NAND2_X1 U9823 ( .A1(n8014), .A2(n7526), .ZN(n7678) );
  AND2_X1 U9824 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7527) );
  NAND2_X1 U9825 ( .A1(n7678), .A2(n8897), .ZN(n7686) );
  INV_X1 U9826 ( .A(n7528), .ZN(n7529) );
  NAND2_X1 U9827 ( .A1(n7529), .A2(SI_1_), .ZN(n7694) );
  NAND2_X1 U9828 ( .A1(n7697), .A2(SI_2_), .ZN(n7530) );
  INV_X1 U9829 ( .A(n7697), .ZN(n7532) );
  INV_X1 U9830 ( .A(SI_2_), .ZN(n7696) );
  NAND2_X1 U9831 ( .A1(n7532), .A2(n7696), .ZN(n7533) );
  INV_X1 U9832 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9678) );
  XNOR2_X1 U9833 ( .A(n7535), .B(SI_3_), .ZN(n7714) );
  INV_X1 U9834 ( .A(n7535), .ZN(n7536) );
  NAND2_X1 U9835 ( .A1(n7536), .A2(SI_3_), .ZN(n7537) );
  MUX2_X1 U9836 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n7417), .Z(n7540) );
  INV_X1 U9837 ( .A(n7731), .ZN(n7539) );
  NAND2_X1 U9838 ( .A1(n7732), .A2(n7539), .ZN(n7542) );
  NAND2_X1 U9839 ( .A1(n7540), .A2(SI_4_), .ZN(n7541) );
  XNOR2_X1 U9840 ( .A(n7543), .B(SI_5_), .ZN(n7740) );
  NAND2_X1 U9841 ( .A1(n7742), .A2(n7740), .ZN(n7546) );
  INV_X1 U9842 ( .A(n7543), .ZN(n7544) );
  NAND2_X1 U9843 ( .A1(n7544), .A2(SI_5_), .ZN(n7545) );
  XNOR2_X1 U9844 ( .A(n7548), .B(SI_6_), .ZN(n7760) );
  INV_X1 U9845 ( .A(n7760), .ZN(n7547) );
  NAND2_X1 U9846 ( .A1(n7761), .A2(n7547), .ZN(n7550) );
  NAND2_X1 U9847 ( .A1(n7548), .A2(SI_6_), .ZN(n7549) );
  NAND2_X1 U9848 ( .A1(n7775), .A2(n7551), .ZN(n7554) );
  NAND2_X1 U9849 ( .A1(n7552), .A2(SI_7_), .ZN(n7553) );
  MUX2_X1 U9850 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9685), .Z(n7556) );
  XNOR2_X1 U9851 ( .A(n7556), .B(SI_8_), .ZN(n7789) );
  INV_X1 U9852 ( .A(n7789), .ZN(n7555) );
  NAND2_X1 U9853 ( .A1(n7556), .A2(SI_8_), .ZN(n7557) );
  MUX2_X1 U9854 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9685), .Z(n7559) );
  XNOR2_X1 U9855 ( .A(n7559), .B(SI_9_), .ZN(n7803) );
  INV_X1 U9856 ( .A(n7803), .ZN(n7558) );
  NAND2_X1 U9857 ( .A1(n7559), .A2(SI_9_), .ZN(n7560) );
  MUX2_X1 U9858 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9685), .Z(n7562) );
  XNOR2_X1 U9859 ( .A(n7562), .B(SI_10_), .ZN(n7820) );
  INV_X1 U9860 ( .A(n7820), .ZN(n7561) );
  MUX2_X1 U9861 ( .A(n9769), .B(n10368), .S(n9685), .Z(n7563) );
  NAND2_X1 U9862 ( .A1(n7563), .A2(n9719), .ZN(n7566) );
  INV_X1 U9863 ( .A(n7563), .ZN(n7564) );
  NAND2_X1 U9864 ( .A1(n7564), .A2(SI_11_), .ZN(n7565) );
  MUX2_X1 U9865 ( .A(n9919), .B(n9916), .S(n9685), .Z(n7567) );
  NAND2_X1 U9866 ( .A1(n7567), .A2(n9728), .ZN(n7570) );
  INV_X1 U9867 ( .A(n7567), .ZN(n7568) );
  NAND2_X1 U9868 ( .A1(n7568), .A2(SI_12_), .ZN(n7569) );
  MUX2_X1 U9869 ( .A(n10019), .B(n10020), .S(n9685), .Z(n7571) );
  NAND2_X1 U9870 ( .A1(n7571), .A2(n9745), .ZN(n7574) );
  INV_X1 U9871 ( .A(n7571), .ZN(n7572) );
  NAND2_X1 U9872 ( .A1(n7572), .A2(SI_13_), .ZN(n7573) );
  MUX2_X1 U9873 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9685), .Z(n7885) );
  MUX2_X1 U9874 ( .A(n10125), .B(n10127), .S(n9685), .Z(n7575) );
  NAND2_X1 U9875 ( .A1(n7575), .A2(n9961), .ZN(n7582) );
  INV_X1 U9876 ( .A(n7575), .ZN(n7576) );
  NAND2_X1 U9877 ( .A1(n7576), .A2(SI_15_), .ZN(n7577) );
  NAND2_X1 U9878 ( .A1(n7582), .A2(n7577), .ZN(n7900) );
  INV_X1 U9879 ( .A(n7885), .ZN(n7578) );
  NOR2_X1 U9880 ( .A1(n7578), .A2(n9772), .ZN(n7579) );
  NOR2_X1 U9881 ( .A1(n7900), .A2(n7579), .ZN(n7580) );
  MUX2_X1 U9882 ( .A(n10236), .B(n10237), .S(n9685), .Z(n7583) );
  NAND2_X1 U9883 ( .A1(n7583), .A2(n10023), .ZN(n7586) );
  INV_X1 U9884 ( .A(n7583), .ZN(n7584) );
  NAND2_X1 U9885 ( .A1(n7584), .A2(SI_16_), .ZN(n7585) );
  MUX2_X1 U9886 ( .A(n10506), .B(n10508), .S(n9685), .Z(n7935) );
  MUX2_X1 U9887 ( .A(n10629), .B(n10627), .S(n9685), .Z(n7948) );
  MUX2_X1 U9888 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9685), .Z(n7588) );
  XNOR2_X1 U9889 ( .A(n7588), .B(SI_19_), .ZN(n7965) );
  INV_X1 U9890 ( .A(n7588), .ZN(n7589) );
  INV_X1 U9891 ( .A(SI_19_), .ZN(n10109) );
  NAND2_X1 U9892 ( .A1(n7589), .A2(n10109), .ZN(n7590) );
  INV_X1 U9893 ( .A(SI_20_), .ZN(n10564) );
  INV_X1 U9894 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11240) );
  MUX2_X1 U9895 ( .A(n11240), .B(n7009), .S(n9685), .Z(n7981) );
  MUX2_X1 U9896 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9685), .Z(n7594) );
  NAND2_X1 U9897 ( .A1(n7594), .A2(SI_21_), .ZN(n7596) );
  OAI21_X1 U9898 ( .B1(SI_21_), .B2(n7594), .A(n7596), .ZN(n7998) );
  INV_X1 U9899 ( .A(n7998), .ZN(n7595) );
  MUX2_X1 U9900 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9685), .Z(n9298) );
  NAND2_X1 U9901 ( .A1(n9302), .A2(n7597), .ZN(n7658) );
  MUX2_X1 U9902 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9685), .Z(n7598) );
  NAND2_X1 U9903 ( .A1(n7598), .A2(SI_23_), .ZN(n7600) );
  OAI21_X1 U9904 ( .B1(SI_23_), .B2(n7598), .A(n7600), .ZN(n7659) );
  INV_X1 U9905 ( .A(n7659), .ZN(n7599) );
  NAND2_X1 U9906 ( .A1(n7658), .A2(n7599), .ZN(n7661) );
  MUX2_X1 U9907 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9685), .Z(n7645) );
  MUX2_X1 U9908 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n9685), .Z(n7605) );
  XNOR2_X1 U9909 ( .A(n7605), .B(SI_25_), .ZN(n8026) );
  MUX2_X1 U9910 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n9685), .Z(n7606) );
  NAND2_X1 U9911 ( .A1(n7606), .A2(SI_26_), .ZN(n7607) );
  OAI21_X1 U9912 ( .B1(SI_26_), .B2(n7606), .A(n7607), .ZN(n7630) );
  INV_X1 U9913 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14249) );
  INV_X1 U9914 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13590) );
  MUX2_X1 U9915 ( .A(n14249), .B(n13590), .S(n9685), .Z(n7618) );
  NAND2_X1 U9916 ( .A1(n7608), .A2(n7618), .ZN(n7610) );
  INV_X1 U9917 ( .A(n7621), .ZN(n7609) );
  INV_X1 U9918 ( .A(SI_27_), .ZN(n11559) );
  INV_X1 U9919 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8213) );
  MUX2_X1 U9920 ( .A(n14246), .B(n8213), .S(n9685), .Z(n8045) );
  XNOR2_X1 U9921 ( .A(n8045), .B(SI_28_), .ZN(n8043) );
  XNOR2_X2 U9922 ( .A(n7612), .B(n7611), .ZN(n14245) );
  NAND2_X1 U9923 ( .A1(n8123), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7613) );
  MUX2_X1 U9924 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7613), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n7614) );
  NAND2_X1 U9925 ( .A1(n13583), .A2(n7923), .ZN(n7617) );
  OR2_X1 U9926 ( .A1(n11750), .A2(n14246), .ZN(n7616) );
  INV_X1 U9927 ( .A(n7618), .ZN(n7619) );
  XNOR2_X1 U9928 ( .A(n7619), .B(SI_27_), .ZN(n7620) );
  XNOR2_X1 U9929 ( .A(n7621), .B(n7620), .ZN(n13588) );
  INV_X2 U9930 ( .A(n7478), .ZN(n7923) );
  NAND2_X1 U9931 ( .A1(n13588), .A2(n7923), .ZN(n7623) );
  OR2_X1 U9932 ( .A1(n11750), .A2(n14249), .ZN(n7622) );
  NAND2_X1 U9933 ( .A1(n11760), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n7629) );
  INV_X1 U9934 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n13941) );
  OR2_X1 U9935 ( .A1(n8034), .A2(n13941), .ZN(n7628) );
  INV_X1 U9936 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7624) );
  NAND2_X1 U9937 ( .A1(n7638), .A2(n7624), .ZN(n7625) );
  NAND2_X1 U9938 ( .A1(n8051), .A2(n7625), .ZN(n13940) );
  OR2_X1 U9939 ( .A1(n8053), .A2(n13940), .ZN(n7627) );
  INV_X1 U9940 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n14201) );
  OR2_X1 U9941 ( .A1(n7992), .A2(n14201), .ZN(n7626) );
  NAND4_X1 U9942 ( .A1(n7629), .A2(n7628), .A3(n7627), .A4(n7626), .ZN(n13746)
         );
  INV_X1 U9943 ( .A(n13746), .ZN(n12123) );
  XNOR2_X1 U9944 ( .A(n13939), .B(n12123), .ZN(n11978) );
  NAND2_X1 U9945 ( .A1(n7631), .A2(n7630), .ZN(n7632) );
  NAND2_X1 U9946 ( .A1(n13591), .A2(n7923), .ZN(n7635) );
  INV_X1 U9947 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14251) );
  OR2_X1 U9948 ( .A1(n11750), .A2(n14251), .ZN(n7634) );
  NAND2_X1 U9949 ( .A1(n8049), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n7643) );
  INV_X1 U9950 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n7636) );
  OR2_X1 U9951 ( .A1(n8072), .A2(n7636), .ZN(n7642) );
  INV_X1 U9952 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13726) );
  NAND2_X1 U9953 ( .A1(n8032), .A2(n13726), .ZN(n7637) );
  NAND2_X1 U9954 ( .A1(n7638), .A2(n7637), .ZN(n13724) );
  OR2_X1 U9955 ( .A1(n8053), .A2(n13724), .ZN(n7641) );
  INV_X1 U9956 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n7639) );
  OR2_X1 U9957 ( .A1(n8034), .A2(n7639), .ZN(n7640) );
  NAND4_X1 U9958 ( .A1(n7643), .A2(n7642), .A3(n7641), .A4(n7640), .ZN(n13747)
         );
  NAND2_X1 U9959 ( .A1(n13950), .A2(n13747), .ZN(n7644) );
  INV_X1 U9960 ( .A(n13747), .ZN(n12110) );
  NAND2_X1 U9961 ( .A1(n14120), .A2(n12110), .ZN(n8039) );
  NAND2_X1 U9962 ( .A1(n7646), .A2(n6895), .ZN(n7647) );
  NAND2_X1 U9963 ( .A1(n11935), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7649) );
  NAND2_X1 U9964 ( .A1(n8049), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7657) );
  INV_X1 U9965 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n7651) );
  OR2_X1 U9966 ( .A1(n8072), .A2(n7651), .ZN(n7656) );
  OAI21_X1 U9967 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n7652), .A(n8030), .ZN(
        n13682) );
  OR2_X1 U9968 ( .A1(n8053), .A2(n13682), .ZN(n7655) );
  INV_X1 U9969 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n7653) );
  OR2_X1 U9970 ( .A1(n8034), .A2(n7653), .ZN(n7654) );
  NAND4_X1 U9971 ( .A1(n7657), .A2(n7656), .A3(n7655), .A4(n7654), .ZN(n13749)
         );
  INV_X1 U9972 ( .A(n7658), .ZN(n7660) );
  NAND2_X1 U9973 ( .A1(n7660), .A2(n7659), .ZN(n7662) );
  NAND2_X1 U9974 ( .A1(n11692), .A2(n7923), .ZN(n7664) );
  INV_X1 U9975 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11695) );
  OR2_X1 U9976 ( .A1(n11750), .A2(n11695), .ZN(n7663) );
  NAND2_X1 U9977 ( .A1(n11760), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n7671) );
  INV_X1 U9978 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10390) );
  OR2_X1 U9979 ( .A1(n7992), .A2(n10390), .ZN(n7670) );
  OAI21_X1 U9980 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n7666), .A(n7665), .ZN(
        n14001) );
  OR2_X1 U9981 ( .A1(n8053), .A2(n14001), .ZN(n7669) );
  INV_X1 U9982 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n7667) );
  OR2_X1 U9983 ( .A1(n8034), .A2(n7667), .ZN(n7668) );
  NAND4_X1 U9984 ( .A1(n7671), .A2(n7670), .A3(n7669), .A4(n7668), .ZN(n13750)
         );
  XNOR2_X1 U9985 ( .A(n14212), .B(n13750), .ZN(n13995) );
  NAND2_X1 U9986 ( .A1(n11759), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7675) );
  INV_X1 U9987 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9760) );
  INV_X1 U9988 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10595) );
  INV_X1 U9989 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7672) );
  INV_X1 U9990 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n13785) );
  INV_X1 U9991 ( .A(SI_0_), .ZN(n7676) );
  INV_X1 U9992 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8283) );
  OAI21_X1 U9993 ( .B1(n9685), .B2(n7676), .A(n8283), .ZN(n7677) );
  NAND2_X1 U9994 ( .A1(n7678), .A2(n7677), .ZN(n14266) );
  MUX2_X1 U9995 ( .A(n13785), .B(n14266), .S(n9755), .Z(n10130) );
  NAND2_X1 U9996 ( .A1(n8049), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n7685) );
  INV_X1 U9997 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10539) );
  OR2_X1 U9998 ( .A1(n8053), .A2(n10539), .ZN(n7684) );
  INV_X1 U9999 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9775) );
  OR2_X1 U10000 ( .A1(n8034), .A2(n9775), .ZN(n7683) );
  INV_X1 U10001 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7681) );
  XNOR2_X1 U10002 ( .A(n7687), .B(n7686), .ZN(n9692) );
  INV_X2 U10003 ( .A(n9755), .ZN(n7970) );
  NAND2_X1 U10004 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n7688) );
  MUX2_X1 U10005 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7688), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n7690) );
  INV_X1 U10006 ( .A(n7700), .ZN(n7689) );
  NAND2_X1 U10007 ( .A1(n7690), .A2(n7689), .ZN(n9796) );
  INV_X1 U10008 ( .A(n9796), .ZN(n13778) );
  NAND2_X1 U10009 ( .A1(n7970), .A2(n13778), .ZN(n7691) );
  NAND2_X1 U10010 ( .A1(n13772), .A2(n10131), .ZN(n11769) );
  NAND2_X1 U10011 ( .A1(n7692), .A2(n11769), .ZN(n7693) );
  NAND2_X1 U10012 ( .A1(n7695), .A2(n7694), .ZN(n7699) );
  XNOR2_X1 U10013 ( .A(n7697), .B(n7696), .ZN(n7698) );
  XNOR2_X1 U10014 ( .A(n7699), .B(n7698), .ZN(n9690) );
  NOR2_X1 U10015 ( .A1(n7700), .A2(n7806), .ZN(n7701) );
  MUX2_X1 U10016 ( .A(n7806), .B(n7701), .S(P1_IR_REG_2__SCAN_IN), .Z(n7702)
         );
  NOR2_X1 U10017 ( .A1(n7702), .A2(n7734), .ZN(n13792) );
  NAND2_X1 U10018 ( .A1(n7970), .A2(n13792), .ZN(n7704) );
  INV_X1 U10019 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9691) );
  OR2_X1 U10020 ( .A1(n11750), .A2(n9691), .ZN(n7703) );
  NAND2_X1 U10021 ( .A1(n11759), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7711) );
  INV_X1 U10022 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n13790) );
  OR2_X1 U10023 ( .A1(n8053), .A2(n13790), .ZN(n7710) );
  INV_X1 U10024 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7706) );
  INV_X1 U10025 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9795) );
  OR2_X1 U10026 ( .A1(n7707), .A2(n9795), .ZN(n7708) );
  NAND2_X1 U10027 ( .A1(n13771), .A2(n14682), .ZN(n11783) );
  INV_X1 U10028 ( .A(n11956), .ZN(n7712) );
  NAND2_X1 U10029 ( .A1(n10116), .A2(n7712), .ZN(n7713) );
  XNOR2_X1 U10030 ( .A(n7715), .B(n7714), .ZN(n9672) );
  NAND2_X1 U10031 ( .A1(n11934), .A2(n9672), .ZN(n7719) );
  OR2_X1 U10032 ( .A1(n11750), .A2(n9678), .ZN(n7718) );
  OR2_X1 U10033 ( .A1(n7734), .A2(n7806), .ZN(n7716) );
  XNOR2_X1 U10034 ( .A(n7716), .B(P1_IR_REG_3__SCAN_IN), .ZN(n13809) );
  NAND2_X1 U10035 ( .A1(n7970), .A2(n13809), .ZN(n7717) );
  NAND2_X1 U10036 ( .A1(n11760), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7724) );
  OR2_X1 U10037 ( .A1(n8053), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n7723) );
  INV_X1 U10038 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10536) );
  OR2_X1 U10039 ( .A1(n8034), .A2(n10536), .ZN(n7722) );
  INV_X1 U10040 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7720) );
  OR2_X1 U10041 ( .A1(n7992), .A2(n7720), .ZN(n7721) );
  NAND2_X1 U10042 ( .A1(n13770), .A2(n14703), .ZN(n11792) );
  NAND2_X1 U10043 ( .A1(n10533), .A2(n11789), .ZN(n7725) );
  NAND2_X1 U10044 ( .A1(n7725), .A2(n11791), .ZN(n14660) );
  NAND2_X1 U10045 ( .A1(n8049), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n7730) );
  INV_X1 U10046 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7726) );
  OR2_X1 U10047 ( .A1(n8072), .A2(n7726), .ZN(n7729) );
  OAI21_X1 U10048 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n7751), .ZN(n14666) );
  OR2_X1 U10049 ( .A1(n8053), .A2(n14666), .ZN(n7728) );
  INV_X1 U10050 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9780) );
  OR2_X1 U10051 ( .A1(n8034), .A2(n9780), .ZN(n7727) );
  INV_X1 U10052 ( .A(n11798), .ZN(n13769) );
  XNOR2_X1 U10053 ( .A(n7732), .B(n7731), .ZN(n9676) );
  NAND2_X1 U10054 ( .A1(n9676), .A2(n7923), .ZN(n7737) );
  NAND2_X1 U10055 ( .A1(n7734), .A2(n7733), .ZN(n7743) );
  NAND2_X1 U10056 ( .A1(n7743), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7735) );
  XNOR2_X1 U10057 ( .A(n7735), .B(P1_IR_REG_4__SCAN_IN), .ZN(n13820) );
  AOI22_X1 U10058 ( .A1(n11935), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n7970), 
        .B2(n13820), .ZN(n7736) );
  AND2_X2 U10059 ( .A1(n7737), .A2(n7736), .ZN(n14708) );
  XNOR2_X1 U10060 ( .A(n13769), .B(n14708), .ZN(n14671) );
  INV_X1 U10061 ( .A(n14671), .ZN(n14661) );
  NAND2_X1 U10062 ( .A1(n14660), .A2(n14661), .ZN(n7739) );
  INV_X1 U10063 ( .A(n14708), .ZN(n14676) );
  NAND2_X1 U10064 ( .A1(n11798), .A2(n14676), .ZN(n7738) );
  NAND2_X1 U10065 ( .A1(n7739), .A2(n7738), .ZN(n10512) );
  INV_X1 U10066 ( .A(n7740), .ZN(n7741) );
  XNOR2_X1 U10067 ( .A(n7742), .B(n7741), .ZN(n9681) );
  NAND2_X1 U10068 ( .A1(n9681), .A2(n7923), .ZN(n7749) );
  NOR2_X1 U10069 ( .A1(n7743), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n7746) );
  OR2_X1 U10070 ( .A1(n7746), .A2(n7806), .ZN(n7744) );
  MUX2_X1 U10071 ( .A(P1_IR_REG_31__SCAN_IN), .B(n7744), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n7747) );
  NAND2_X1 U10072 ( .A1(n7746), .A2(n7745), .ZN(n7776) );
  AND2_X1 U10073 ( .A1(n7747), .A2(n7776), .ZN(n9801) );
  AOI22_X1 U10074 ( .A1(n11935), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7970), 
        .B2(n9801), .ZN(n7748) );
  NAND2_X1 U10075 ( .A1(n7749), .A2(n7748), .ZN(n11804) );
  NAND2_X1 U10076 ( .A1(n8049), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n7756) );
  INV_X1 U10077 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9802) );
  OR2_X1 U10078 ( .A1(n8072), .A2(n9802), .ZN(n7755) );
  INV_X1 U10079 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9783) );
  OR2_X1 U10080 ( .A1(n8034), .A2(n9783), .ZN(n7754) );
  AND2_X1 U10081 ( .A1(n7751), .A2(n7750), .ZN(n7752) );
  OR2_X1 U10082 ( .A1(n7752), .A2(n7765), .ZN(n10844) );
  OR2_X1 U10083 ( .A1(n8053), .A2(n10844), .ZN(n7753) );
  NAND4_X1 U10084 ( .A1(n7756), .A2(n7755), .A3(n7754), .A4(n7753), .ZN(n13768) );
  XNOR2_X1 U10085 ( .A(n11804), .B(n13768), .ZN(n11958) );
  NAND2_X1 U10086 ( .A1(n10512), .A2(n11958), .ZN(n7759) );
  INV_X1 U10087 ( .A(n13768), .ZN(n7757) );
  NAND2_X1 U10088 ( .A1(n11804), .A2(n7757), .ZN(n7758) );
  NAND2_X1 U10089 ( .A1(n7759), .A2(n7758), .ZN(n14644) );
  XNOR2_X1 U10090 ( .A(n7761), .B(n7760), .ZN(n9699) );
  NAND2_X1 U10091 ( .A1(n9699), .A2(n7923), .ZN(n7764) );
  NAND2_X1 U10092 ( .A1(n7776), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7762) );
  XNOR2_X1 U10093 ( .A(n7762), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9805) );
  AOI22_X1 U10094 ( .A1(n11935), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7970), 
        .B2(n9805), .ZN(n7763) );
  NAND2_X1 U10095 ( .A1(n7764), .A2(n7763), .ZN(n14648) );
  NAND2_X1 U10096 ( .A1(n8049), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n7770) );
  INV_X1 U10097 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9804) );
  OR2_X1 U10098 ( .A1(n8072), .A2(n9804), .ZN(n7769) );
  OR2_X1 U10099 ( .A1(n7765), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7766) );
  NAND2_X1 U10100 ( .A1(n7782), .A2(n7766), .ZN(n14649) );
  OR2_X1 U10101 ( .A1(n8053), .A2(n14649), .ZN(n7768) );
  INV_X1 U10102 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9784) );
  OR2_X1 U10103 ( .A1(n8034), .A2(n9784), .ZN(n7767) );
  NAND4_X1 U10104 ( .A1(n7770), .A2(n7769), .A3(n7768), .A4(n7767), .ZN(n13767) );
  INV_X1 U10105 ( .A(n13767), .ZN(n7771) );
  AND2_X1 U10106 ( .A1(n14648), .A2(n7771), .ZN(n7773) );
  OR2_X1 U10107 ( .A1(n14648), .A2(n7771), .ZN(n7772) );
  XNOR2_X1 U10108 ( .A(n7775), .B(n7774), .ZN(n9723) );
  NAND2_X1 U10109 ( .A1(n9723), .A2(n7923), .ZN(n7779) );
  NAND2_X1 U10110 ( .A1(n7791), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7777) );
  XNOR2_X1 U10111 ( .A(n7777), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9808) );
  AOI22_X1 U10112 ( .A1(n11935), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7970), 
        .B2(n9808), .ZN(n7778) );
  NAND2_X1 U10113 ( .A1(n7779), .A2(n7778), .ZN(n14725) );
  NAND2_X1 U10114 ( .A1(n11760), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7787) );
  INV_X1 U10115 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7780) );
  OR2_X1 U10116 ( .A1(n7673), .A2(n7780), .ZN(n7786) );
  NAND2_X1 U10117 ( .A1(n7782), .A2(n7781), .ZN(n7783) );
  NAND2_X1 U10118 ( .A1(n7796), .A2(n7783), .ZN(n11274) );
  OR2_X1 U10119 ( .A1(n8053), .A2(n11274), .ZN(n7785) );
  INV_X1 U10120 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10587) );
  OR2_X1 U10121 ( .A1(n8034), .A2(n10587), .ZN(n7784) );
  NAND4_X1 U10122 ( .A1(n7787), .A2(n7786), .A3(n7785), .A4(n7784), .ZN(n13766) );
  XNOR2_X1 U10123 ( .A(n14725), .B(n13766), .ZN(n11960) );
  INV_X1 U10124 ( .A(n11960), .ZN(n10582) );
  INV_X1 U10125 ( .A(n13766), .ZN(n11269) );
  NAND2_X1 U10126 ( .A1(n14725), .A2(n11269), .ZN(n7788) );
  XNOR2_X1 U10127 ( .A(n7790), .B(n7789), .ZN(n9730) );
  NAND2_X1 U10128 ( .A1(n9730), .A2(n7923), .ZN(n7794) );
  NAND2_X1 U10129 ( .A1(n7805), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7792) );
  XNOR2_X1 U10130 ( .A(n7792), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9811) );
  AOI22_X1 U10131 ( .A1(n11935), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7970), 
        .B2(n9811), .ZN(n7793) );
  NAND2_X1 U10132 ( .A1(n7794), .A2(n7793), .ZN(n11820) );
  NAND2_X1 U10133 ( .A1(n8049), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7801) );
  INV_X1 U10134 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9810) );
  OR2_X1 U10135 ( .A1(n8072), .A2(n9810), .ZN(n7800) );
  NAND2_X1 U10136 ( .A1(n7796), .A2(n7795), .ZN(n7797) );
  NAND2_X1 U10137 ( .A1(n7813), .A2(n7797), .ZN(n11009) );
  OR2_X1 U10138 ( .A1(n8053), .A2(n11009), .ZN(n7799) );
  INV_X1 U10139 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9785) );
  OR2_X1 U10140 ( .A1(n8034), .A2(n9785), .ZN(n7798) );
  NAND4_X1 U10141 ( .A1(n7801), .A2(n7800), .A3(n7799), .A4(n7798), .ZN(n13765) );
  INV_X1 U10142 ( .A(n13765), .ZN(n11345) );
  XNOR2_X1 U10143 ( .A(n11820), .B(n11345), .ZN(n11963) );
  OR2_X1 U10144 ( .A1(n11820), .A2(n11345), .ZN(n7802) );
  XNOR2_X1 U10145 ( .A(n7804), .B(n7803), .ZN(n9740) );
  NAND2_X1 U10146 ( .A1(n9740), .A2(n7923), .ZN(n7812) );
  NOR2_X1 U10147 ( .A1(n7835), .A2(n7806), .ZN(n7807) );
  NAND2_X1 U10148 ( .A1(n7807), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n7810) );
  INV_X1 U10149 ( .A(n7807), .ZN(n7809) );
  INV_X1 U10150 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n7808) );
  NAND2_X1 U10151 ( .A1(n7809), .A2(n7808), .ZN(n7822) );
  AOI22_X1 U10152 ( .A1(n9900), .A2(n7970), .B1(n11935), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n7811) );
  NAND2_X1 U10153 ( .A1(n7812), .A2(n7811), .ZN(n11829) );
  NAND2_X1 U10154 ( .A1(n8049), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7819) );
  INV_X1 U10155 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9794) );
  OR2_X1 U10156 ( .A1(n8072), .A2(n9794), .ZN(n7818) );
  INV_X1 U10157 ( .A(n7839), .ZN(n7815) );
  NAND2_X1 U10158 ( .A1(n7813), .A2(n9790), .ZN(n7814) );
  NAND2_X1 U10159 ( .A1(n7815), .A2(n7814), .ZN(n11407) );
  OR2_X1 U10160 ( .A1(n8053), .A2(n11407), .ZN(n7817) );
  INV_X1 U10161 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10983) );
  OR2_X1 U10162 ( .A1(n8034), .A2(n10983), .ZN(n7816) );
  NAND4_X1 U10163 ( .A1(n7819), .A2(n7818), .A3(n7817), .A4(n7816), .ZN(n13764) );
  XNOR2_X1 U10164 ( .A(n11829), .B(n11398), .ZN(n11964) );
  XNOR2_X1 U10165 ( .A(n7821), .B(n7820), .ZN(n9749) );
  NAND2_X1 U10166 ( .A1(n9749), .A2(n7923), .ZN(n7825) );
  NAND2_X1 U10167 ( .A1(n7822), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7823) );
  XNOR2_X1 U10168 ( .A(n7823), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9904) );
  AOI22_X1 U10169 ( .A1(n9904), .A2(n7970), .B1(n11935), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n7824) );
  NAND2_X1 U10170 ( .A1(n11760), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7830) );
  INV_X1 U10171 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11000) );
  OR2_X1 U10172 ( .A1(n8034), .A2(n11000), .ZN(n7829) );
  XNOR2_X1 U10173 ( .A(n7839), .B(P1_REG3_REG_10__SCAN_IN), .ZN(n11491) );
  OR2_X1 U10174 ( .A1(n8053), .A2(n11491), .ZN(n7828) );
  INV_X1 U10175 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7826) );
  OR2_X1 U10176 ( .A1(n7673), .A2(n7826), .ZN(n7827) );
  NAND4_X1 U10177 ( .A1(n7830), .A2(n7829), .A3(n7828), .A4(n7827), .ZN(n13763) );
  INV_X1 U10178 ( .A(n13763), .ZN(n11484) );
  XNOR2_X1 U10179 ( .A(n14747), .B(n11484), .ZN(n11965) );
  OR2_X1 U10180 ( .A1(n14747), .A2(n11484), .ZN(n7831) );
  NAND2_X1 U10181 ( .A1(n9768), .A2(n7923), .ZN(n7838) );
  NOR2_X1 U10182 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n7834) );
  NAND2_X1 U10183 ( .A1(n7835), .A2(n7834), .ZN(n7849) );
  NAND2_X1 U10184 ( .A1(n7849), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7836) );
  XNOR2_X1 U10185 ( .A(n7836), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U10186 ( .A1(n10148), .A2(n7970), .B1(n11935), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n7837) );
  NAND2_X1 U10187 ( .A1(n11759), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7847) );
  INV_X1 U10188 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9906) );
  OR2_X1 U10189 ( .A1(n8072), .A2(n9906), .ZN(n7846) );
  NAND2_X1 U10190 ( .A1(n7839), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7841) );
  INV_X1 U10191 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7840) );
  NAND2_X1 U10192 ( .A1(n7841), .A2(n7840), .ZN(n7842) );
  NAND2_X1 U10193 ( .A1(n7842), .A2(n7853), .ZN(n11653) );
  OR2_X1 U10194 ( .A1(n8053), .A2(n11653), .ZN(n7845) );
  INV_X1 U10195 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7843) );
  OR2_X1 U10196 ( .A1(n7992), .A2(n7843), .ZN(n7844) );
  NAND4_X1 U10197 ( .A1(n7847), .A2(n7846), .A3(n7845), .A4(n7844), .ZN(n13762) );
  INV_X1 U10198 ( .A(n13762), .ZN(n11641) );
  XNOR2_X1 U10199 ( .A(n7848), .B(n7486), .ZN(n9915) );
  NAND2_X1 U10200 ( .A1(n9915), .A2(n7923), .ZN(n7851) );
  NAND2_X1 U10201 ( .A1(n7909), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7864) );
  XNOR2_X1 U10202 ( .A(n7864), .B(P1_IR_REG_12__SCAN_IN), .ZN(n13854) );
  AOI22_X1 U10203 ( .A1(n13854), .A2(n7970), .B1(n11935), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n7850) );
  NAND2_X1 U10204 ( .A1(n11759), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7859) );
  INV_X1 U10205 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10151) );
  OR2_X1 U10206 ( .A1(n8072), .A2(n10151), .ZN(n7858) );
  NAND2_X1 U10207 ( .A1(n7853), .A2(n7852), .ZN(n7854) );
  NAND2_X1 U10208 ( .A1(n7873), .A2(n7854), .ZN(n14396) );
  OR2_X1 U10209 ( .A1(n8053), .A2(n14396), .ZN(n7857) );
  INV_X1 U10210 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7855) );
  OR2_X1 U10211 ( .A1(n7673), .A2(n7855), .ZN(n7856) );
  XNOR2_X1 U10212 ( .A(n14399), .B(n13761), .ZN(n14391) );
  NAND2_X1 U10213 ( .A1(n14407), .A2(n13761), .ZN(n7860) );
  XNOR2_X1 U10214 ( .A(n7862), .B(n7482), .ZN(n10018) );
  NAND2_X1 U10215 ( .A1(n10018), .A2(n7923), .ZN(n7871) );
  INV_X1 U10216 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n7863) );
  NAND2_X1 U10217 ( .A1(n7864), .A2(n7863), .ZN(n7865) );
  NAND2_X1 U10218 ( .A1(n7865), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7867) );
  INV_X1 U10219 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n7866) );
  NAND2_X1 U10220 ( .A1(n7867), .A2(n7866), .ZN(n7888) );
  OR2_X1 U10221 ( .A1(n7867), .A2(n7866), .ZN(n7868) );
  NOR2_X1 U10222 ( .A1(n11750), .A2(n10019), .ZN(n7869) );
  AOI21_X1 U10223 ( .B1(n10169), .B2(n7970), .A(n7869), .ZN(n7870) );
  NAND2_X1 U10224 ( .A1(n11760), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7880) );
  INV_X1 U10225 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11321) );
  OR2_X1 U10226 ( .A1(n8034), .A2(n11321), .ZN(n7879) );
  INV_X1 U10227 ( .A(n7892), .ZN(n7875) );
  NAND2_X1 U10228 ( .A1(n7873), .A2(n7872), .ZN(n7874) );
  NAND2_X1 U10229 ( .A1(n7875), .A2(n7874), .ZN(n11721) );
  OR2_X1 U10230 ( .A1(n8053), .A2(n11721), .ZN(n7878) );
  INV_X1 U10231 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7876) );
  OR2_X1 U10232 ( .A1(n7992), .A2(n7876), .ZN(n7877) );
  XNOR2_X1 U10233 ( .A(n14585), .B(n11840), .ZN(n11970) );
  INV_X1 U10234 ( .A(n11970), .ZN(n11314) );
  NAND2_X1 U10235 ( .A1(n11316), .A2(n11314), .ZN(n7882) );
  INV_X1 U10236 ( .A(n11840), .ZN(n13760) );
  NAND2_X1 U10237 ( .A1(n11839), .A2(n13760), .ZN(n7881) );
  NAND2_X1 U10238 ( .A1(n7882), .A2(n7881), .ZN(n11575) );
  NAND2_X1 U10239 ( .A1(n7883), .A2(n9772), .ZN(n7901) );
  OR2_X1 U10240 ( .A1(n7883), .A2(n9772), .ZN(n7884) );
  NAND2_X1 U10241 ( .A1(n7901), .A2(n7884), .ZN(n7886) );
  OR2_X1 U10242 ( .A1(n7886), .A2(n7885), .ZN(n7903) );
  NAND2_X1 U10243 ( .A1(n7886), .A2(n7885), .ZN(n7887) );
  NAND2_X1 U10244 ( .A1(n7903), .A2(n7887), .ZN(n10239) );
  NAND2_X1 U10245 ( .A1(n10239), .A2(n7923), .ZN(n7891) );
  NAND2_X1 U10246 ( .A1(n7888), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7889) );
  XNOR2_X1 U10247 ( .A(n7889), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U10248 ( .A1(n10915), .A2(n7970), .B1(n11935), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n7890) );
  NOR2_X1 U10249 ( .A1(n7892), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7893) );
  OR2_X1 U10250 ( .A1(n7913), .A2(n7893), .ZN(n14559) );
  INV_X1 U10251 ( .A(n14559), .ZN(n7894) );
  NAND2_X1 U10252 ( .A1(n8022), .A2(n7894), .ZN(n7899) );
  INV_X1 U10253 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10172) );
  OR2_X1 U10254 ( .A1(n8072), .A2(n10172), .ZN(n7898) );
  INV_X1 U10255 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10905) );
  OR2_X1 U10256 ( .A1(n8034), .A2(n10905), .ZN(n7897) );
  INV_X1 U10257 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n7895) );
  OR2_X1 U10258 ( .A1(n7673), .A2(n7895), .ZN(n7896) );
  NAND2_X1 U10259 ( .A1(n14558), .A2(n12016), .ZN(n11857) );
  AND2_X1 U10260 ( .A1(n7901), .A2(n7900), .ZN(n7902) );
  NAND2_X1 U10261 ( .A1(n7903), .A2(n7902), .ZN(n7905) );
  NAND2_X1 U10262 ( .A1(n7905), .A2(n7904), .ZN(n10124) );
  NAND2_X1 U10263 ( .A1(n10124), .A2(n7923), .ZN(n7912) );
  INV_X1 U10264 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n7906) );
  NAND2_X1 U10265 ( .A1(n7907), .A2(n7906), .ZN(n7908) );
  OAI21_X1 U10266 ( .B1(n7909), .B2(n7908), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n7910) );
  XNOR2_X1 U10267 ( .A(n7910), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10918) );
  AOI22_X1 U10268 ( .A1(n10918), .A2(n7970), .B1(n11935), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n7911) );
  OR2_X1 U10269 ( .A1(n7913), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7914) );
  AND2_X1 U10270 ( .A1(n7927), .A2(n7914), .ZN(n13733) );
  NAND2_X1 U10271 ( .A1(n8022), .A2(n13733), .ZN(n7920) );
  INV_X1 U10272 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7915) );
  OR2_X1 U10273 ( .A1(n7992), .A2(n7915), .ZN(n7919) );
  INV_X1 U10274 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7916) );
  OR2_X1 U10275 ( .A1(n8072), .A2(n7916), .ZN(n7918) );
  INV_X1 U10276 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11475) );
  OR2_X1 U10277 ( .A1(n8034), .A2(n11475), .ZN(n7917) );
  NAND2_X1 U10278 ( .A1(n13738), .A2(n12024), .ZN(n11863) );
  NAND2_X1 U10279 ( .A1(n11862), .A2(n11863), .ZN(n11969) );
  NAND2_X1 U10280 ( .A1(n11468), .A2(n11467), .ZN(n7921) );
  XNOR2_X1 U10281 ( .A(n7922), .B(n7481), .ZN(n10235) );
  NAND2_X1 U10282 ( .A1(n10235), .A2(n7923), .ZN(n7926) );
  NAND2_X1 U10283 ( .A1(n7938), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7924) );
  XNOR2_X1 U10284 ( .A(n7924), .B(P1_IR_REG_16__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U10285 ( .A1(n11935), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7970), 
        .B2(n11615), .ZN(n7925) );
  NAND2_X1 U10286 ( .A1(n7927), .A2(n10912), .ZN(n7928) );
  NAND2_X1 U10287 ( .A1(n7943), .A2(n7928), .ZN(n13655) );
  OAI22_X1 U10288 ( .A1(n13655), .A2(n8053), .B1(n8034), .B2(n11627), .ZN(
        n7932) );
  INV_X1 U10289 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U10290 ( .A1(n11760), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n7929) );
  OAI21_X1 U10291 ( .B1(n7930), .B2(n7673), .A(n7929), .ZN(n7931) );
  XNOR2_X1 U10292 ( .A(n14571), .B(n13757), .ZN(n11972) );
  INV_X1 U10293 ( .A(n11972), .ZN(n11610) );
  INV_X1 U10294 ( .A(n13757), .ZN(n7933) );
  NAND2_X1 U10295 ( .A1(n14571), .A2(n7933), .ZN(n7934) );
  XNOR2_X1 U10296 ( .A(n7935), .B(SI_17_), .ZN(n7936) );
  XNOR2_X1 U10297 ( .A(n7937), .B(n7936), .ZN(n10505) );
  NAND2_X1 U10298 ( .A1(n10505), .A2(n7923), .ZN(n7942) );
  NAND2_X1 U10299 ( .A1(n7939), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7940) );
  XNOR2_X1 U10300 ( .A(n7940), .B(P1_IR_REG_17__SCAN_IN), .ZN(n11623) );
  AOI22_X1 U10301 ( .A1(n11935), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7970), 
        .B2(n11623), .ZN(n7941) );
  AND2_X1 U10302 ( .A1(n7943), .A2(n13671), .ZN(n7944) );
  OR2_X1 U10303 ( .A1(n7944), .A2(n7957), .ZN(n14085) );
  AOI22_X1 U10304 ( .A1(n8049), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n11760), 
        .B2(P1_REG1_REG_17__SCAN_IN), .ZN(n7946) );
  NAND2_X1 U10305 ( .A1(n11759), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7945) );
  OAI211_X1 U10306 ( .C1(n14085), .C2(n8053), .A(n7946), .B(n7945), .ZN(n13756) );
  NOR2_X1 U10307 ( .A1(n14088), .A2(n13756), .ZN(n11870) );
  INV_X1 U10308 ( .A(n11870), .ZN(n7947) );
  INV_X1 U10309 ( .A(n13756), .ZN(n13712) );
  NAND2_X1 U10310 ( .A1(n7949), .A2(n7948), .ZN(n7950) );
  NAND2_X1 U10311 ( .A1(n7951), .A2(n7950), .ZN(n10628) );
  OR2_X1 U10312 ( .A1(n10628), .A2(n7478), .ZN(n7956) );
  NAND2_X1 U10313 ( .A1(n8117), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7954) );
  XNOR2_X1 U10314 ( .A(n7954), .B(P1_IR_REG_18__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U10315 ( .A1(n11935), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7970), 
        .B2(n11629), .ZN(n7955) );
  OR2_X1 U10316 ( .A1(n7957), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n7958) );
  AND2_X1 U10317 ( .A1(n7974), .A2(n7958), .ZN(n14072) );
  NAND2_X1 U10318 ( .A1(n14072), .A2(n8022), .ZN(n7962) );
  AOI22_X1 U10319 ( .A1(n8049), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n11760), 
        .B2(P1_REG1_REG_18__SCAN_IN), .ZN(n7961) );
  INV_X1 U10320 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n7959) );
  OR2_X1 U10321 ( .A1(n8034), .A2(n7959), .ZN(n7960) );
  INV_X1 U10322 ( .A(n13668), .ZN(n13755) );
  XNOR2_X1 U10323 ( .A(n14179), .B(n13755), .ZN(n14076) );
  NAND2_X1 U10324 ( .A1(n14066), .A2(n14076), .ZN(n7964) );
  NAND2_X1 U10325 ( .A1(n14074), .A2(n13755), .ZN(n7963) );
  XNOR2_X1 U10326 ( .A(n7966), .B(n7965), .ZN(n10787) );
  NAND2_X1 U10327 ( .A1(n10787), .A2(n7923), .ZN(n7972) );
  NAND2_X2 U10328 ( .A1(n8064), .A2(n7969), .ZN(n14564) );
  AOI22_X1 U10329 ( .A1(n11935), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14058), 
        .B2(n7970), .ZN(n7971) );
  NAND2_X1 U10330 ( .A1(n7974), .A2(n7973), .ZN(n7975) );
  NAND2_X1 U10331 ( .A1(n7987), .A2(n7975), .ZN(n14059) );
  OR2_X1 U10332 ( .A1(n14059), .A2(n8053), .ZN(n7980) );
  INV_X1 U10333 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14176) );
  NAND2_X1 U10334 ( .A1(n11759), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n7977) );
  NAND2_X1 U10335 ( .A1(n8049), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n7976) );
  OAI211_X1 U10336 ( .C1(n8072), .C2(n14176), .A(n7977), .B(n7976), .ZN(n7978)
         );
  INV_X1 U10337 ( .A(n7978), .ZN(n7979) );
  OR2_X1 U10338 ( .A1(n13621), .A2(n13714), .ZN(n11878) );
  NAND2_X1 U10339 ( .A1(n13621), .A2(n13714), .ZN(n11879) );
  NAND2_X1 U10340 ( .A1(n7982), .A2(n7981), .ZN(n7983) );
  NAND2_X1 U10341 ( .A1(n11214), .A2(n7923), .ZN(n7986) );
  OR2_X1 U10342 ( .A1(n11750), .A2(n11240), .ZN(n7985) );
  NAND2_X1 U10343 ( .A1(n7987), .A2(n13691), .ZN(n7988) );
  NAND2_X1 U10344 ( .A1(n8005), .A2(n7988), .ZN(n14044) );
  INV_X1 U10345 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n7991) );
  NAND2_X1 U10346 ( .A1(n11760), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n7990) );
  NAND2_X1 U10347 ( .A1(n11759), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n7989) );
  OAI211_X1 U10348 ( .C1(n7992), .C2(n7991), .A(n7990), .B(n7989), .ZN(n7993)
         );
  INV_X1 U10349 ( .A(n7993), .ZN(n7994) );
  NAND2_X1 U10350 ( .A1(n14165), .A2(n13753), .ZN(n7996) );
  INV_X1 U10351 ( .A(n13753), .ZN(n12058) );
  NAND2_X1 U10352 ( .A1(n14043), .A2(n12058), .ZN(n7995) );
  NAND2_X1 U10353 ( .A1(n7996), .A2(n7995), .ZN(n11975) );
  INV_X1 U10354 ( .A(n7997), .ZN(n7999) );
  NAND2_X1 U10355 ( .A1(n7999), .A2(n7998), .ZN(n8001) );
  AND2_X1 U10356 ( .A1(n8001), .A2(n8000), .ZN(n11363) );
  NAND2_X1 U10357 ( .A1(n11363), .A2(n7923), .ZN(n8003) );
  INV_X1 U10358 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11391) );
  OR2_X1 U10359 ( .A1(n11750), .A2(n11391), .ZN(n8002) );
  AND2_X1 U10360 ( .A1(n8005), .A2(n8004), .ZN(n8006) );
  OR2_X1 U10361 ( .A1(n8006), .A2(n8016), .ZN(n14026) );
  INV_X1 U10362 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10259) );
  NAND2_X1 U10363 ( .A1(n11759), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8008) );
  NAND2_X1 U10364 ( .A1(n8049), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8007) );
  OAI211_X1 U10365 ( .C1(n8072), .C2(n10259), .A(n8008), .B(n8007), .ZN(n8009)
         );
  INV_X1 U10366 ( .A(n8009), .ZN(n8010) );
  OAI21_X1 U10367 ( .B1(n14026), .B2(n8053), .A(n8010), .ZN(n13752) );
  INV_X1 U10368 ( .A(n13752), .ZN(n8011) );
  XNOR2_X1 U10369 ( .A(n14220), .B(n8011), .ZN(n14021) );
  INV_X1 U10370 ( .A(n14021), .ZN(n8105) );
  NAND2_X1 U10371 ( .A1(n14022), .A2(n8105), .ZN(n8013) );
  OR2_X1 U10372 ( .A1(n14220), .A2(n8011), .ZN(n8012) );
  NAND2_X1 U10373 ( .A1(n9297), .A2(n8014), .ZN(n8015) );
  XNOR2_X1 U10374 ( .A(n8015), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14265) );
  OR2_X1 U10375 ( .A1(n8016), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8018) );
  AND2_X1 U10376 ( .A1(n8018), .A2(n8017), .ZN(n14012) );
  INV_X1 U10377 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n14215) );
  NAND2_X1 U10378 ( .A1(n11759), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8020) );
  NAND2_X1 U10379 ( .A1(n11760), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8019) );
  OAI211_X1 U10380 ( .C1(n7673), .C2(n14215), .A(n8020), .B(n8019), .ZN(n8021)
         );
  AOI21_X1 U10381 ( .B1(n14012), .B2(n8022), .A(n8021), .ZN(n13635) );
  INV_X1 U10382 ( .A(n13635), .ZN(n13751) );
  XNOR2_X1 U10383 ( .A(n14217), .B(n13751), .ZN(n14009) );
  OR2_X1 U10384 ( .A1(n14217), .A2(n13751), .ZN(n8023) );
  INV_X1 U10385 ( .A(n13750), .ZN(n12083) );
  NAND2_X1 U10386 ( .A1(n14212), .A2(n12083), .ZN(n8024) );
  AND2_X2 U10387 ( .A1(n13993), .A2(n8024), .ZN(n13979) );
  INV_X1 U10388 ( .A(n13749), .ZN(n12091) );
  OR2_X1 U10389 ( .A1(n14132), .A2(n12091), .ZN(n8025) );
  INV_X1 U10390 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14257) );
  OR2_X1 U10391 ( .A1(n11750), .A2(n14257), .ZN(n8028) );
  NAND2_X1 U10392 ( .A1(n8049), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8038) );
  INV_X1 U10393 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n14129) );
  OR2_X1 U10394 ( .A1(n8072), .A2(n14129), .ZN(n8037) );
  INV_X1 U10395 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8029) );
  NAND2_X1 U10396 ( .A1(n8030), .A2(n8029), .ZN(n8031) );
  NAND2_X1 U10397 ( .A1(n8032), .A2(n8031), .ZN(n13965) );
  OR2_X1 U10398 ( .A1(n8053), .A2(n13965), .ZN(n8036) );
  INV_X1 U10399 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n8033) );
  OR2_X1 U10400 ( .A1(n8034), .A2(n8033), .ZN(n8035) );
  NAND4_X1 U10401 ( .A1(n8038), .A2(n8037), .A3(n8036), .A4(n8035), .ZN(n13748) );
  INV_X1 U10402 ( .A(n13748), .ZN(n12100) );
  NAND2_X1 U10403 ( .A1(n13951), .A2(n8039), .ZN(n13933) );
  NAND2_X1 U10404 ( .A1(n13932), .A2(n13933), .ZN(n13931) );
  NAND2_X1 U10405 ( .A1(n13939), .A2(n12123), .ZN(n8040) );
  OAI21_X1 U10406 ( .B1(n12134), .B2(n13915), .A(n13914), .ZN(n8042) );
  NAND2_X1 U10407 ( .A1(n13915), .A2(n12134), .ZN(n8041) );
  NAND2_X1 U10408 ( .A1(n8042), .A2(n8041), .ZN(n8059) );
  INV_X1 U10409 ( .A(SI_28_), .ZN(n12965) );
  NAND2_X1 U10410 ( .A1(n8045), .A2(n12965), .ZN(n8046) );
  INV_X1 U10411 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14243) );
  INV_X1 U10412 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13582) );
  MUX2_X1 U10413 ( .A(n14243), .B(n13582), .S(n9685), .Z(n9417) );
  XNOR2_X1 U10414 ( .A(n9417), .B(SI_29_), .ZN(n9415) );
  NAND2_X1 U10415 ( .A1(n13580), .A2(n7923), .ZN(n8048) );
  NAND2_X1 U10416 ( .A1(n11935), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8047) );
  INV_X1 U10417 ( .A(n14108), .ZN(n11922) );
  NAND2_X1 U10418 ( .A1(n8049), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8058) );
  INV_X1 U10419 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8050) );
  OR2_X1 U10420 ( .A1(n8072), .A2(n8050), .ZN(n8057) );
  INV_X1 U10421 ( .A(n8051), .ZN(n8052) );
  NAND2_X1 U10422 ( .A1(n8052), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n13901) );
  OR2_X1 U10423 ( .A1(n8053), .A2(n13901), .ZN(n8056) );
  INV_X1 U10424 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8054) );
  OR2_X1 U10425 ( .A1(n8034), .A2(n8054), .ZN(n8055) );
  AND4_X1 U10426 ( .A1(n8058), .A2(n8057), .A3(n8056), .A4(n8055), .ZN(n12138)
         );
  INV_X1 U10427 ( .A(n12138), .ZN(n13744) );
  XNOR2_X1 U10428 ( .A(n11922), .B(n13744), .ZN(n11980) );
  XNOR2_X1 U10429 ( .A(n8059), .B(n11980), .ZN(n13911) );
  NAND2_X1 U10430 ( .A1(n8062), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8061) );
  MUX2_X1 U10431 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8061), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n8063) );
  NAND2_X1 U10432 ( .A1(n14264), .A2(n14058), .ZN(n8068) );
  NAND2_X1 U10433 ( .A1(n6490), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8067) );
  NAND2_X1 U10434 ( .A1(n8069), .A2(n8113), .ZN(n11928) );
  NAND2_X1 U10435 ( .A1(n10133), .A2(n14682), .ZN(n10112) );
  NAND2_X1 U10436 ( .A1(n14208), .A2(n13984), .ZN(n13962) );
  NAND2_X1 U10437 ( .A1(n14108), .A2(n8070), .ZN(n13895) );
  OAI211_X1 U10438 ( .C1(n14108), .C2(n8070), .A(n14655), .B(n13895), .ZN(
        n13908) );
  INV_X1 U10439 ( .A(n14247), .ZN(n11990) );
  NAND2_X1 U10440 ( .A1(n11990), .A2(P1_B_REG_SCAN_IN), .ZN(n8071) );
  NAND2_X1 U10441 ( .A1(n6462), .A2(n8071), .ZN(n13890) );
  INV_X1 U10442 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n14105) );
  OR2_X1 U10443 ( .A1(n8072), .A2(n14105), .ZN(n8076) );
  INV_X1 U10444 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n8073) );
  OR2_X1 U10445 ( .A1(n8034), .A2(n8073), .ZN(n8075) );
  INV_X1 U10446 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14195) );
  OR2_X1 U10447 ( .A1(n7673), .A2(n14195), .ZN(n8074) );
  AND3_X1 U10448 ( .A1(n8076), .A2(n8075), .A3(n8074), .ZN(n11927) );
  OR2_X1 U10449 ( .A1(n13890), .A2(n11927), .ZN(n13902) );
  INV_X1 U10450 ( .A(n11941), .ZN(n9626) );
  NAND2_X1 U10451 ( .A1(n13725), .A2(n13745), .ZN(n13904) );
  NAND3_X1 U10452 ( .A1(n13908), .A2(n13902), .A3(n13904), .ZN(n8077) );
  AND2_X2 U10453 ( .A1(n11774), .A2(n11769), .ZN(n11954) );
  AND2_X1 U10454 ( .A1(n10135), .A2(n7679), .ZN(n10128) );
  INV_X1 U10455 ( .A(n10131), .ZN(n11778) );
  NAND2_X1 U10456 ( .A1(n10111), .A2(n11956), .ZN(n8079) );
  INV_X1 U10457 ( .A(n14682), .ZN(n10114) );
  OR2_X1 U10458 ( .A1(n10114), .A2(n13771), .ZN(n8078) );
  NAND2_X1 U10459 ( .A1(n8079), .A2(n8078), .ZN(n10528) );
  NAND2_X1 U10460 ( .A1(n10528), .A2(n11957), .ZN(n8081) );
  OR2_X1 U10461 ( .A1(n10532), .A2(n13770), .ZN(n8080) );
  NAND2_X1 U10462 ( .A1(n14672), .A2(n14671), .ZN(n8083) );
  NAND2_X1 U10463 ( .A1(n11798), .A2(n14708), .ZN(n8082) );
  NAND2_X1 U10464 ( .A1(n10509), .A2(n10513), .ZN(n8085) );
  OR2_X1 U10465 ( .A1(n11804), .A2(n13768), .ZN(n8084) );
  XNOR2_X1 U10466 ( .A(n14648), .B(n13767), .ZN(n11959) );
  NAND2_X1 U10467 ( .A1(n14642), .A2(n14643), .ZN(n8087) );
  OR2_X1 U10468 ( .A1(n14648), .A2(n13767), .ZN(n8086) );
  NAND2_X1 U10469 ( .A1(n10592), .A2(n10582), .ZN(n8089) );
  OR2_X1 U10470 ( .A1(n14725), .A2(n13766), .ZN(n8088) );
  OR2_X1 U10471 ( .A1(n11820), .A2(n13765), .ZN(n8090) );
  NAND2_X1 U10472 ( .A1(n10994), .A2(n11965), .ZN(n8092) );
  OR2_X1 U10473 ( .A1(n14747), .A2(n13763), .ZN(n8091) );
  NAND2_X1 U10474 ( .A1(n11188), .A2(n7116), .ZN(n8094) );
  OR2_X1 U10475 ( .A1(n11837), .A2(n13762), .ZN(n8093) );
  NAND2_X1 U10476 ( .A1(n14390), .A2(n7110), .ZN(n8096) );
  NAND2_X1 U10477 ( .A1(n14407), .A2(n11841), .ZN(n8095) );
  NAND2_X1 U10478 ( .A1(n11315), .A2(n11970), .ZN(n8098) );
  NAND2_X1 U10479 ( .A1(n11839), .A2(n11840), .ZN(n8097) );
  INV_X1 U10480 ( .A(n12016), .ZN(n13759) );
  NAND2_X1 U10481 ( .A1(n14558), .A2(n13759), .ZN(n8099) );
  INV_X1 U10482 ( .A(n12024), .ZN(n13758) );
  NAND2_X1 U10483 ( .A1(n11603), .A2(n11610), .ZN(n8101) );
  OR2_X1 U10484 ( .A1(n14571), .A2(n13757), .ZN(n8100) );
  AND2_X1 U10485 ( .A1(n14179), .A2(n13755), .ZN(n11874) );
  OR2_X1 U10486 ( .A1(n14179), .A2(n13755), .ZN(n11873) );
  NAND2_X1 U10487 ( .A1(n14052), .A2(n14053), .ZN(n8103) );
  INV_X1 U10488 ( .A(n13714), .ZN(n13754) );
  OR2_X1 U10489 ( .A1(n13621), .A2(n13754), .ZN(n8102) );
  NAND2_X1 U10490 ( .A1(n14043), .A2(n13753), .ZN(n8104) );
  NAND2_X1 U10491 ( .A1(n14009), .A2(n14008), .ZN(n14007) );
  NAND2_X1 U10492 ( .A1(n14217), .A2(n13635), .ZN(n8106) );
  NAND2_X1 U10493 ( .A1(n14212), .A2(n13750), .ZN(n8107) );
  OR2_X1 U10494 ( .A1(n14132), .A2(n13749), .ZN(n8108) );
  NAND2_X1 U10495 ( .A1(n13972), .A2(n13748), .ZN(n8109) );
  OR2_X1 U10496 ( .A1(n13939), .A2(n13746), .ZN(n8110) );
  XNOR2_X1 U10497 ( .A(n13915), .B(n12134), .ZN(n13922) );
  NAND2_X1 U10498 ( .A1(n13915), .A2(n13745), .ZN(n8111) );
  NAND2_X1 U10499 ( .A1(n13921), .A2(n8111), .ZN(n8112) );
  XNOR2_X1 U10500 ( .A(n8112), .B(n11980), .ZN(n13900) );
  NAND2_X2 U10501 ( .A1(n11938), .A2(n8113), .ZN(n10518) );
  OAI21_X1 U10502 ( .B1(n11753), .B2(n10518), .A(n12132), .ZN(n10527) );
  NAND2_X1 U10503 ( .A1(n11939), .A2(n14058), .ZN(n11754) );
  NAND2_X1 U10504 ( .A1(n13900), .A2(n14753), .ZN(n8114) );
  OAI21_X1 U10505 ( .B1(n8117), .B2(n8116), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8118) );
  INV_X1 U10506 ( .A(P1_B_REG_SCAN_IN), .ZN(n8119) );
  MUX2_X1 U10507 ( .A(n8121), .B(P1_B_REG_SCAN_IN), .S(n14260), .Z(n8125) );
  NAND2_X1 U10508 ( .A1(n6557), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8122) );
  MUX2_X1 U10509 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8122), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n8124) );
  NAND2_X1 U10510 ( .A1(n8125), .A2(n14250), .ZN(n9735) );
  OR2_X1 U10511 ( .A1(n9735), .A2(P1_D_REG_0__SCAN_IN), .ZN(n8126) );
  OR2_X1 U10512 ( .A1(n14260), .A2(n14250), .ZN(n9736) );
  NAND2_X1 U10513 ( .A1(n11938), .A2(n14564), .ZN(n8127) );
  NAND2_X1 U10514 ( .A1(n9626), .A2(n8127), .ZN(n9642) );
  INV_X1 U10515 ( .A(n9642), .ZN(n8128) );
  NOR2_X1 U10516 ( .A1(n9643), .A2(n8128), .ZN(n8143) );
  NOR2_X1 U10517 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .ZN(
        n8132) );
  NOR4_X1 U10518 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n8131) );
  NOR4_X1 U10519 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n8130) );
  NOR4_X1 U10520 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n8129) );
  NAND4_X1 U10521 ( .A1(n8132), .A2(n8131), .A3(n8130), .A4(n8129), .ZN(n8138)
         );
  NOR4_X1 U10522 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n8136) );
  NOR4_X1 U10523 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n8135) );
  NOR4_X1 U10524 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n8134) );
  NOR4_X1 U10525 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n8133) );
  NAND4_X1 U10526 ( .A1(n8136), .A2(n8135), .A3(n8134), .A4(n8133), .ZN(n8137)
         );
  NOR2_X1 U10527 ( .A1(n8138), .A2(n8137), .ZN(n8139) );
  OR2_X1 U10528 ( .A1(n9735), .A2(n8139), .ZN(n9630) );
  NAND2_X1 U10529 ( .A1(n8141), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8142) );
  AND2_X1 U10530 ( .A1(n9630), .A2(n9753), .ZN(n9644) );
  AND2_X1 U10531 ( .A1(n8143), .A2(n9644), .ZN(n10517) );
  NAND2_X1 U10532 ( .A1(n8144), .A2(n9746), .ZN(n9624) );
  AND2_X1 U10533 ( .A1(n9624), .A2(n9639), .ZN(n10025) );
  NAND2_X1 U10534 ( .A1(n10028), .A2(n14058), .ZN(n8145) );
  NAND2_X1 U10535 ( .A1(n14756), .A2(n14724), .ZN(n14232) );
  INV_X4 U10536 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U10537 ( .A(n8286), .ZN(n8146) );
  NAND2_X1 U10538 ( .A1(n8146), .A2(n8287), .ZN(n8149) );
  NAND2_X1 U10539 ( .A1(n8147), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8148) );
  INV_X1 U10540 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9675) );
  NAND2_X1 U10541 ( .A1(n9675), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8151) );
  NAND2_X1 U10542 ( .A1(n9691), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8150) );
  AND2_X1 U10543 ( .A1(n8151), .A2(n8150), .ZN(n8304) );
  NAND2_X1 U10544 ( .A1(n8964), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8153) );
  NAND2_X1 U10545 ( .A1(n9678), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8152) );
  AND2_X1 U10546 ( .A1(n8153), .A2(n8152), .ZN(n8318) );
  NAND2_X1 U10547 ( .A1(n9677), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8155) );
  INV_X1 U10548 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9696) );
  NAND2_X1 U10549 ( .A1(n9696), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8154) );
  AND2_X1 U10550 ( .A1(n8155), .A2(n8154), .ZN(n8332) );
  NAND2_X1 U10551 ( .A1(n9683), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8157) );
  NAND2_X1 U10552 ( .A1(n9698), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8156) );
  AND2_X1 U10553 ( .A1(n8157), .A2(n8156), .ZN(n8350) );
  NAND2_X1 U10554 ( .A1(n8351), .A2(n8350), .ZN(n8353) );
  NAND2_X1 U10555 ( .A1(n9700), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8158) );
  NAND2_X1 U10556 ( .A1(n9702), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8159) );
  NAND2_X1 U10557 ( .A1(n9724), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8163) );
  NAND2_X1 U10558 ( .A1(n9726), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8161) );
  AND2_X1 U10559 ( .A1(n8163), .A2(n8161), .ZN(n8383) );
  INV_X1 U10560 ( .A(n8383), .ZN(n8162) );
  NAND2_X1 U10561 ( .A1(n9734), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U10562 ( .A1(n9732), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8164) );
  AND2_X1 U10563 ( .A1(n8165), .A2(n8164), .ZN(n8395) );
  NAND2_X1 U10564 ( .A1(n9743), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U10565 ( .A1(n9741), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8166) );
  NAND2_X1 U10566 ( .A1(n8168), .A2(n8166), .ZN(n8415) );
  INV_X1 U10567 ( .A(n8415), .ZN(n8167) );
  NAND2_X1 U10568 ( .A1(n8416), .A2(n8167), .ZN(n8169) );
  NAND2_X1 U10569 ( .A1(n9750), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8171) );
  INV_X1 U10570 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U10571 ( .A1(n9752), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8170) );
  AND2_X1 U10572 ( .A1(n8171), .A2(n8170), .ZN(n8428) );
  NAND2_X1 U10573 ( .A1(n9769), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8173) );
  NAND2_X1 U10574 ( .A1(n10368), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8172) );
  NAND2_X1 U10575 ( .A1(n9919), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8176) );
  NAND2_X1 U10576 ( .A1(n9916), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8174) );
  NAND2_X1 U10577 ( .A1(n8176), .A2(n8174), .ZN(n8463) );
  INV_X1 U10578 ( .A(n8463), .ZN(n8175) );
  NAND2_X1 U10579 ( .A1(n8464), .A2(n8175), .ZN(n8177) );
  NAND2_X1 U10580 ( .A1(n8178), .A2(n10019), .ZN(n8180) );
  NAND2_X1 U10581 ( .A1(n8181), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8183) );
  INV_X1 U10582 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10106) );
  NAND2_X1 U10583 ( .A1(n10106), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8182) );
  NAND2_X1 U10584 ( .A1(n10125), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8186) );
  NAND2_X1 U10585 ( .A1(n10127), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8184) );
  NAND2_X1 U10586 ( .A1(n8186), .A2(n8184), .ZN(n8506) );
  INV_X1 U10587 ( .A(n8506), .ZN(n8185) );
  NAND2_X1 U10588 ( .A1(n10236), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8189) );
  NAND2_X1 U10589 ( .A1(n10237), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8187) );
  NAND2_X1 U10590 ( .A1(n8189), .A2(n8187), .ZN(n8520) );
  INV_X1 U10591 ( .A(n8520), .ZN(n8188) );
  NAND2_X1 U10592 ( .A1(n8521), .A2(n8188), .ZN(n8190) );
  NAND2_X1 U10593 ( .A1(n8190), .A2(n8189), .ZN(n8535) );
  NAND2_X1 U10594 ( .A1(n10506), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8192) );
  NAND2_X1 U10595 ( .A1(n10508), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8191) );
  NAND2_X1 U10596 ( .A1(n10629), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8194) );
  NAND2_X1 U10597 ( .A1(n10627), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8193) );
  NAND2_X1 U10598 ( .A1(n8555), .A2(n8554), .ZN(n8557) );
  INV_X1 U10599 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10790) );
  NAND2_X1 U10600 ( .A1(n10790), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8196) );
  INV_X1 U10601 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10788) );
  NAND2_X1 U10602 ( .A1(n10788), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8195) );
  NAND2_X1 U10603 ( .A1(n11391), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8199) );
  INV_X1 U10604 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11365) );
  NAND2_X1 U10605 ( .A1(n11365), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8198) );
  INV_X1 U10606 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11677) );
  XNOR2_X1 U10607 ( .A(n11677), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8614) );
  NAND2_X1 U10608 ( .A1(n11677), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8200) );
  XNOR2_X1 U10609 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8624) );
  INV_X1 U10610 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8201) );
  NAND2_X1 U10611 ( .A1(n8201), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8202) );
  INV_X1 U10612 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13600) );
  NAND2_X1 U10613 ( .A1(n8204), .A2(n13600), .ZN(n8205) );
  INV_X1 U10614 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13596) );
  XNOR2_X1 U10615 ( .A(n13596), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8644) );
  NAND2_X1 U10616 ( .A1(n13596), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8207) );
  INV_X1 U10617 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13592) );
  AND2_X1 U10618 ( .A1(n13592), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8208) );
  NAND2_X1 U10619 ( .A1(n14251), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8209) );
  INV_X1 U10620 ( .A(n8671), .ZN(n8211) );
  NAND2_X1 U10621 ( .A1(n14249), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8210) );
  NAND2_X1 U10622 ( .A1(n13590), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8212) );
  AND2_X1 U10623 ( .A1(n8213), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8214) );
  NAND2_X1 U10624 ( .A1(n14246), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8215) );
  XNOR2_X1 U10625 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n8693) );
  NAND2_X1 U10626 ( .A1(n14243), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8216) );
  INV_X1 U10627 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n11999) );
  XNOR2_X1 U10628 ( .A(n11999), .B(P1_DATAO_REG_30__SCAN_IN), .ZN(n8268) );
  XNOR2_X1 U10629 ( .A(n8269), .B(n8268), .ZN(n12955) );
  NAND2_X1 U10630 ( .A1(n8235), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8236) );
  INV_X1 U10631 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8238) );
  NAND2_X2 U10632 ( .A1(n9652), .A2(n9684), .ZN(n8602) );
  NAND2_X1 U10633 ( .A1(n12955), .A2(n8684), .ZN(n8243) );
  NAND2_X4 U10634 ( .A1(n9652), .A2(n9685), .ZN(n8575) );
  NAND2_X1 U10635 ( .A1(n8288), .A2(SI_30_), .ZN(n8242) );
  NAND2_X1 U10636 ( .A1(n8243), .A2(n8242), .ZN(n8706) );
  NOR2_X1 U10637 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8343) );
  NAND2_X1 U10638 ( .A1(n8343), .A2(n11309), .ZN(n8362) );
  NOR2_X1 U10639 ( .A1(n8377), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8389) );
  NAND2_X1 U10640 ( .A1(n8404), .A2(n8403), .ZN(n8435) );
  NAND2_X1 U10641 ( .A1(n8478), .A2(n8477), .ZN(n8499) );
  INV_X1 U10642 ( .A(n8513), .ZN(n8245) );
  INV_X1 U10643 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8244) );
  NAND2_X1 U10644 ( .A1(n8245), .A2(n8244), .ZN(n8527) );
  INV_X1 U10645 ( .A(n8544), .ZN(n8247) );
  INV_X1 U10646 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8246) );
  NAND2_X1 U10647 ( .A1(n8247), .A2(n8246), .ZN(n8562) );
  INV_X1 U10648 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8248) );
  INV_X1 U10649 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8250) );
  INV_X1 U10650 ( .A(n8637), .ZN(n8253) );
  INV_X1 U10651 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8252) );
  NAND2_X1 U10652 ( .A1(n8253), .A2(n8252), .ZN(n8648) );
  INV_X1 U10653 ( .A(n8648), .ZN(n8255) );
  INV_X1 U10654 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8254) );
  NAND2_X1 U10655 ( .A1(n8255), .A2(n8254), .ZN(n8661) );
  INV_X1 U10656 ( .A(n8674), .ZN(n8257) );
  INV_X1 U10657 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8256) );
  NAND2_X1 U10658 ( .A1(n8257), .A2(n8256), .ZN(n8687) );
  XNOR2_X2 U10659 ( .A(n8258), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U10660 ( .A1(n8259), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8260) );
  MUX2_X1 U10661 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8260), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n8261) );
  NAND2_X1 U10663 ( .A1(n12262), .A2(n6469), .ZN(n8704) );
  INV_X1 U10664 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n10387) );
  NAND2_X1 U10665 ( .A1(n8546), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8265) );
  NAND2_X1 U10666 ( .A1(n8699), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8264) );
  OAI211_X1 U10667 ( .C1(n10387), .C2(n6473), .A(n8265), .B(n8264), .ZN(n8266)
         );
  INV_X1 U10668 ( .A(n8266), .ZN(n8267) );
  NOR2_X1 U10669 ( .A1(n8706), .A2(n12259), .ZN(n8842) );
  XNOR2_X1 U10670 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n8270) );
  NAND2_X1 U10671 ( .A1(n12949), .A2(n8684), .ZN(n8273) );
  NAND2_X1 U10672 ( .A1(n8288), .A2(SI_31_), .ZN(n8272) );
  INV_X1 U10673 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n10392) );
  NAND2_X1 U10674 ( .A1(n8342), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n8276) );
  INV_X1 U10675 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n8274) );
  OR2_X1 U10676 ( .A1(n6471), .A2(n8274), .ZN(n8275) );
  OAI211_X1 U10677 ( .C1(n10392), .C2(n6473), .A(n8276), .B(n8275), .ZN(n8277)
         );
  INV_X1 U10678 ( .A(n8277), .ZN(n8278) );
  INV_X1 U10679 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10867) );
  NAND2_X1 U10680 ( .A1(n8310), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8281) );
  INV_X2 U10681 ( .A(n8293), .ZN(n8698) );
  NAND2_X1 U10682 ( .A1(n8298), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8279) );
  NAND2_X1 U10683 ( .A1(n8283), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8284) );
  NAND2_X1 U10684 ( .A1(n8286), .A2(n8284), .ZN(n8285) );
  MUX2_X1 U10685 ( .A(n8285), .B(SI_0_), .S(n9685), .Z(n12967) );
  MUX2_X1 U10686 ( .A(P3_IR_REG_0__SCAN_IN), .B(n12967), .S(n9652), .Z(n10870)
         );
  INV_X1 U10687 ( .A(n10870), .ZN(n10646) );
  XNOR2_X1 U10688 ( .A(n8287), .B(n8286), .ZN(n9688) );
  NAND2_X1 U10689 ( .A1(n8288), .A2(SI_1_), .ZN(n8291) );
  INV_X1 U10690 ( .A(n9652), .ZN(n8449) );
  NAND2_X1 U10691 ( .A1(n8449), .A2(n6737), .ZN(n8290) );
  NAND2_X1 U10692 ( .A1(n8310), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8297) );
  NAND2_X1 U10693 ( .A1(n8298), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8296) );
  INV_X1 U10694 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8292) );
  OR2_X1 U10695 ( .A1(n8293), .A2(n8292), .ZN(n8295) );
  INV_X1 U10696 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10949) );
  OR2_X1 U10697 ( .A1(n6470), .A2(n10949), .ZN(n8294) );
  NAND2_X1 U10698 ( .A1(n10935), .A2(n8826), .ZN(n9523) );
  NAND2_X1 U10699 ( .A1(n9523), .A2(n9518), .ZN(n15191) );
  NAND2_X1 U10700 ( .A1(n8699), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8302) );
  NAND2_X1 U10701 ( .A1(n8310), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8301) );
  NAND2_X1 U10702 ( .A1(n8698), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8300) );
  NAND2_X1 U10703 ( .A1(n8298), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8299) );
  OAI21_X1 U10704 ( .B1(n8305), .B2(n8304), .A(n8303), .ZN(n9703) );
  INV_X1 U10705 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8307) );
  NAND2_X1 U10706 ( .A1(n8449), .A2(n6475), .ZN(n8309) );
  OAI211_X1 U10707 ( .C1(n8602), .C2(n9703), .A(n6530), .B(n8309), .ZN(n11040)
         );
  INV_X1 U10708 ( .A(n12462), .ZN(n11041) );
  INV_X1 U10709 ( .A(n11040), .ZN(n15198) );
  NAND2_X1 U10710 ( .A1(n11041), .A2(n15198), .ZN(n8723) );
  INV_X1 U10711 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n8311) );
  NAND2_X1 U10712 ( .A1(n8310), .A2(n8311), .ZN(n8317) );
  INV_X1 U10713 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n8312) );
  OR2_X1 U10714 ( .A1(n8293), .A2(n8312), .ZN(n8315) );
  INV_X1 U10715 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n8313) );
  OR2_X1 U10716 ( .A1(n6471), .A2(n8313), .ZN(n8314) );
  OR2_X1 U10717 ( .A1(n8319), .A2(n8318), .ZN(n8320) );
  NAND2_X1 U10718 ( .A1(n8321), .A2(n8320), .ZN(n9713) );
  NOR3_X1 U10719 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n8322) );
  INV_X1 U10720 ( .A(n8322), .ZN(n8323) );
  NAND2_X1 U10721 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n8323), .ZN(n8324) );
  XNOR2_X1 U10722 ( .A(n8324), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10502) );
  OAI22_X1 U10723 ( .A1(n8602), .A2(n9713), .B1(n10502), .B2(n6722), .ZN(n8326) );
  NOR2_X1 U10724 ( .A1(n8575), .A2(SI_3_), .ZN(n8325) );
  NOR2_X2 U10725 ( .A1(n8326), .A2(n8325), .ZN(n11327) );
  NAND2_X1 U10726 ( .A1(n15186), .A2(n11327), .ZN(n8727) );
  NAND2_X1 U10727 ( .A1(n11039), .A2(n11046), .ZN(n8327) );
  INV_X1 U10728 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11332) );
  OR2_X1 U10729 ( .A1(n6471), .A2(n11332), .ZN(n8331) );
  NAND2_X1 U10730 ( .A1(n8298), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8330) );
  OR2_X1 U10731 ( .A1(n7485), .A2(n8343), .ZN(n11333) );
  NAND2_X1 U10732 ( .A1(n8310), .A2(n11333), .ZN(n8329) );
  NAND2_X1 U10733 ( .A1(n8698), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8328) );
  NAND4_X1 U10734 ( .A1(n8331), .A2(n8330), .A3(n8329), .A4(n8328), .ZN(n12460) );
  OR2_X1 U10735 ( .A1(n8333), .A2(n8332), .ZN(n8334) );
  AND2_X1 U10736 ( .A1(n8335), .A2(n8334), .ZN(n9718) );
  NAND2_X1 U10737 ( .A1(n8336), .A2(n9718), .ZN(n8340) );
  NAND2_X1 U10738 ( .A1(n8337), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8338) );
  XNOR2_X1 U10739 ( .A(n8338), .B(n8218), .ZN(n11088) );
  NAND2_X1 U10740 ( .A1(n8449), .A2(n11088), .ZN(n8339) );
  OAI211_X1 U10741 ( .C1(SI_4_), .C2(n8575), .A(n8340), .B(n8339), .ZN(n9534)
         );
  XNOR2_X1 U10742 ( .A(n12460), .B(n9534), .ZN(n12213) );
  INV_X1 U10743 ( .A(n12460), .ZN(n15164) );
  INV_X1 U10744 ( .A(n9534), .ZN(n15223) );
  NAND2_X1 U10745 ( .A1(n15164), .A2(n15223), .ZN(n8341) );
  NAND2_X1 U10746 ( .A1(n8342), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8349) );
  OR2_X1 U10747 ( .A1(n8343), .A2(n11309), .ZN(n8344) );
  NAND2_X1 U10748 ( .A1(n8362), .A2(n8344), .ZN(n15172) );
  NAND2_X1 U10749 ( .A1(n8529), .A2(n15172), .ZN(n8348) );
  INV_X1 U10750 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15175) );
  OR2_X1 U10751 ( .A1(n6471), .A2(n15175), .ZN(n8347) );
  INV_X1 U10752 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n8345) );
  OR2_X1 U10753 ( .A1(n8678), .A2(n8345), .ZN(n8346) );
  OR2_X1 U10754 ( .A1(n8351), .A2(n8350), .ZN(n8352) );
  NAND2_X1 U10755 ( .A1(n8353), .A2(n8352), .ZN(n9709) );
  INV_X1 U10756 ( .A(n8355), .ZN(n8359) );
  NAND2_X1 U10757 ( .A1(n8356), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8357) );
  MUX2_X1 U10758 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8357), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8358) );
  NAND2_X1 U10759 ( .A1(n8359), .A2(n8358), .ZN(n11115) );
  OAI22_X1 U10760 ( .A1(n8602), .A2(n9709), .B1(n14987), .B2(n6722), .ZN(n8361) );
  NOR2_X1 U10761 ( .A1(n8575), .A2(SI_5_), .ZN(n8360) );
  NOR2_X1 U10762 ( .A1(n8361), .A2(n8360), .ZN(n15171) );
  NAND2_X1 U10763 ( .A1(n12212), .A2(n15171), .ZN(n8737) );
  INV_X1 U10764 ( .A(n12212), .ZN(n15144) );
  INV_X1 U10765 ( .A(n15171), .ZN(n12211) );
  NAND2_X1 U10766 ( .A1(n15144), .A2(n12211), .ZN(n8736) );
  NAND2_X1 U10767 ( .A1(n8342), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U10768 ( .A1(n8362), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8363) );
  NAND2_X1 U10769 ( .A1(n8377), .A2(n8363), .ZN(n15150) );
  NAND2_X1 U10770 ( .A1(n8529), .A2(n15150), .ZN(n8367) );
  INV_X1 U10771 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11118) );
  OR2_X1 U10772 ( .A1(n6471), .A2(n11118), .ZN(n8366) );
  INV_X1 U10773 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8364) );
  OR2_X1 U10774 ( .A1(n8678), .A2(n8364), .ZN(n8365) );
  XNOR2_X1 U10775 ( .A(n9702), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8369) );
  XNOR2_X1 U10776 ( .A(n8370), .B(n8369), .ZN(n9722) );
  NAND2_X1 U10777 ( .A1(n8288), .A2(SI_6_), .ZN(n8375) );
  NOR2_X1 U10778 ( .A1(n8355), .A2(n6724), .ZN(n8371) );
  MUX2_X1 U10779 ( .A(n6724), .B(n8371), .S(P3_IR_REG_6__SCAN_IN), .Z(n8373)
         );
  NAND2_X1 U10780 ( .A1(n8355), .A2(n10376), .ZN(n8399) );
  INV_X1 U10781 ( .A(n8399), .ZN(n8372) );
  INV_X1 U10782 ( .A(n11120), .ZN(n15007) );
  NAND2_X1 U10783 ( .A1(n8449), .A2(n15007), .ZN(n8374) );
  OAI211_X1 U10784 ( .C1(n9722), .C2(n8602), .A(n8375), .B(n8374), .ZN(n15149)
         );
  NAND2_X1 U10785 ( .A1(n15163), .A2(n15149), .ZN(n8740) );
  INV_X1 U10786 ( .A(n15149), .ZN(n8376) );
  NAND2_X1 U10787 ( .A1(n12458), .A2(n8376), .ZN(n8741) );
  NAND2_X1 U10788 ( .A1(n8342), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8382) );
  XNOR2_X1 U10789 ( .A(n8377), .B(P3_REG3_REG_7__SCAN_IN), .ZN(n15133) );
  NAND2_X1 U10790 ( .A1(n8529), .A2(n15133), .ZN(n8381) );
  INV_X1 U10791 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11125) );
  OR2_X1 U10792 ( .A1(n6471), .A2(n11125), .ZN(n8380) );
  INV_X1 U10793 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n8378) );
  OR2_X1 U10794 ( .A1(n8678), .A2(n8378), .ZN(n8379) );
  XNOR2_X1 U10795 ( .A(n8384), .B(n8383), .ZN(n9705) );
  NAND2_X1 U10796 ( .A1(n8399), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8386) );
  XNOR2_X1 U10797 ( .A(n8386), .B(n8385), .ZN(n15021) );
  INV_X1 U10798 ( .A(n15021), .ZN(n11126) );
  OAI22_X1 U10799 ( .A1(n8602), .A2(n9705), .B1(n11126), .B2(n6722), .ZN(n8388) );
  NOR2_X1 U10800 ( .A1(n8575), .A2(SI_7_), .ZN(n8387) );
  NOR2_X1 U10801 ( .A1(n8388), .A2(n8387), .ZN(n12218) );
  NAND2_X1 U10802 ( .A1(n15111), .A2(n12218), .ZN(n8745) );
  INV_X1 U10803 ( .A(n12218), .ZN(n15132) );
  NAND2_X1 U10804 ( .A1(n15143), .A2(n15132), .ZN(n8746) );
  NAND2_X1 U10805 ( .A1(n8745), .A2(n8746), .ZN(n15125) );
  NAND2_X1 U10806 ( .A1(n15122), .A2(n15121), .ZN(n15120) );
  NAND2_X1 U10807 ( .A1(n15120), .A2(n8745), .ZN(n15107) );
  INV_X1 U10808 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11131) );
  OR2_X1 U10809 ( .A1(n6471), .A2(n11131), .ZN(n8394) );
  NAND2_X1 U10810 ( .A1(n8698), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8393) );
  NOR2_X1 U10811 ( .A1(n8389), .A2(n11564), .ZN(n8390) );
  OR2_X1 U10812 ( .A1(n8404), .A2(n8390), .ZN(n15117) );
  NAND2_X1 U10813 ( .A1(n8529), .A2(n15117), .ZN(n8392) );
  NAND2_X1 U10814 ( .A1(n8342), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8391) );
  NAND4_X1 U10815 ( .A1(n8394), .A2(n8393), .A3(n8392), .A4(n8391), .ZN(n12457) );
  INV_X1 U10816 ( .A(n12457), .ZN(n15127) );
  OR2_X1 U10817 ( .A1(n8396), .A2(n8395), .ZN(n8397) );
  NAND2_X1 U10818 ( .A1(n8398), .A2(n8397), .ZN(n9712) );
  NAND2_X1 U10819 ( .A1(n8288), .A2(SI_8_), .ZN(n8402) );
  NAND2_X1 U10820 ( .A1(n8410), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8400) );
  XNOR2_X1 U10821 ( .A(n8400), .B(P3_IR_REG_8__SCAN_IN), .ZN(n15043) );
  NAND2_X1 U10822 ( .A1(n8449), .A2(n15043), .ZN(n8401) );
  OAI211_X1 U10823 ( .C1(n8602), .C2(n9712), .A(n8402), .B(n8401), .ZN(n12225)
         );
  NAND2_X1 U10824 ( .A1(n15127), .A2(n12225), .ZN(n8749) );
  INV_X1 U10825 ( .A(n12225), .ZN(n15116) );
  NAND2_X1 U10826 ( .A1(n12457), .A2(n15116), .ZN(n8750) );
  NAND2_X1 U10827 ( .A1(n15107), .A2(n15110), .ZN(n15106) );
  OR2_X1 U10828 ( .A1(n8404), .A2(n8403), .ZN(n8405) );
  AND2_X1 U10829 ( .A1(n8435), .A2(n8405), .ZN(n15105) );
  INV_X1 U10830 ( .A(n15105), .ZN(n12378) );
  NAND2_X1 U10831 ( .A1(n8529), .A2(n12378), .ZN(n8409) );
  INV_X1 U10832 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15098) );
  OR2_X1 U10833 ( .A1(n6471), .A2(n15098), .ZN(n8408) );
  NAND2_X1 U10834 ( .A1(n8698), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8407) );
  NAND2_X1 U10835 ( .A1(n8342), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8406) );
  NAND4_X1 U10836 ( .A1(n8409), .A2(n8408), .A3(n8407), .A4(n8406), .ZN(n14955) );
  OAI21_X1 U10837 ( .B1(n8410), .B2(P3_IR_REG_8__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8411) );
  MUX2_X1 U10838 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8411), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n8414) );
  INV_X1 U10839 ( .A(n8412), .ZN(n8413) );
  NAND2_X1 U10840 ( .A1(n8414), .A2(n8413), .ZN(n11139) );
  OAI22_X1 U10841 ( .A1(n8575), .A2(SI_9_), .B1(n15057), .B2(n6722), .ZN(n8418) );
  XNOR2_X1 U10842 ( .A(n8416), .B(n8415), .ZN(n9707) );
  NOR2_X1 U10843 ( .A1(n8602), .A2(n9707), .ZN(n8417) );
  INV_X1 U10844 ( .A(n15241), .ZN(n15099) );
  NAND2_X1 U10845 ( .A1(n14955), .A2(n15099), .ZN(n8419) );
  NAND2_X1 U10846 ( .A1(n15089), .A2(n8419), .ZN(n8421) );
  INV_X1 U10847 ( .A(n14955), .ZN(n15112) );
  NAND2_X1 U10848 ( .A1(n15112), .A2(n15241), .ZN(n8420) );
  NAND2_X1 U10849 ( .A1(n8421), .A2(n8420), .ZN(n15084) );
  INV_X1 U10850 ( .A(n15084), .ZN(n8434) );
  XNOR2_X1 U10851 ( .A(n8435), .B(P3_REG3_REG_10__SCAN_IN), .ZN(n15081) );
  NAND2_X1 U10852 ( .A1(n8529), .A2(n15081), .ZN(n8426) );
  NAND2_X1 U10853 ( .A1(n8342), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8425) );
  INV_X1 U10854 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11143) );
  OR2_X1 U10855 ( .A1(n6471), .A2(n11143), .ZN(n8424) );
  INV_X1 U10856 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n8422) );
  OR2_X1 U10857 ( .A1(n6473), .A2(n8422), .ZN(n8423) );
  OR2_X1 U10858 ( .A1(n8412), .A2(n6724), .ZN(n8427) );
  XNOR2_X1 U10859 ( .A(n8427), .B(n8446), .ZN(n11202) );
  INV_X1 U10860 ( .A(n11202), .ZN(n11144) );
  OAI22_X1 U10861 ( .A1(n8575), .A2(SI_10_), .B1(n11144), .B2(n6722), .ZN(
        n8433) );
  OR2_X1 U10862 ( .A1(n8429), .A2(n8428), .ZN(n8430) );
  AND2_X1 U10863 ( .A1(n8431), .A2(n8430), .ZN(n9715) );
  NOR2_X1 U10864 ( .A1(n8602), .A2(n9715), .ZN(n8432) );
  NAND2_X1 U10865 ( .A1(n14495), .A2(n14964), .ZN(n8755) );
  INV_X1 U10866 ( .A(n14964), .ZN(n15085) );
  NAND2_X1 U10867 ( .A1(n12456), .A2(n15085), .ZN(n8757) );
  NAND2_X1 U10868 ( .A1(n8755), .A2(n8757), .ZN(n15083) );
  OAI21_X1 U10869 ( .B1(n8435), .B2(P3_REG3_REG_10__SCAN_IN), .A(
        P3_REG3_REG_11__SCAN_IN), .ZN(n8436) );
  NAND2_X1 U10870 ( .A1(n8436), .A2(n8453), .ZN(n14498) );
  NAND2_X1 U10871 ( .A1(n6469), .A2(n14498), .ZN(n8443) );
  INV_X1 U10872 ( .A(n8342), .ZN(n8437) );
  NAND2_X1 U10873 ( .A1(n8546), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8442) );
  INV_X1 U10874 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n8438) );
  OR2_X1 U10875 ( .A1(n6471), .A2(n8438), .ZN(n8441) );
  INV_X1 U10876 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n8439) );
  OR2_X1 U10877 ( .A1(n6473), .A2(n8439), .ZN(n8440) );
  XNOR2_X1 U10878 ( .A(n8445), .B(n8444), .ZN(n9720) );
  NAND2_X1 U10879 ( .A1(n8684), .A2(n9720), .ZN(n8451) );
  NAND2_X1 U10880 ( .A1(n8412), .A2(n8446), .ZN(n8461) );
  NAND2_X1 U10881 ( .A1(n8461), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8448) );
  XNOR2_X1 U10882 ( .A(n8448), .B(n8447), .ZN(n11422) );
  NAND2_X1 U10883 ( .A1(n8449), .A2(n11422), .ZN(n8450) );
  OAI211_X1 U10884 ( .C1(SI_11_), .C2(n8575), .A(n8451), .B(n8450), .ZN(n14497) );
  INV_X1 U10885 ( .A(n14497), .ZN(n12229) );
  XNOR2_X1 U10886 ( .A(n14956), .B(n12229), .ZN(n14493) );
  AND2_X1 U10887 ( .A1(n14493), .A2(n8757), .ZN(n8452) );
  NAND2_X1 U10888 ( .A1(n14488), .A2(n8452), .ZN(n14490) );
  NAND2_X1 U10889 ( .A1(n12797), .A2(n12229), .ZN(n8758) );
  AND2_X1 U10890 ( .A1(n8453), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8454) );
  OR2_X1 U10891 ( .A1(n8454), .A2(n8478), .ZN(n9601) );
  NAND2_X1 U10892 ( .A1(n6469), .A2(n9601), .ZN(n8460) );
  NAND2_X1 U10893 ( .A1(n8546), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8459) );
  INV_X1 U10894 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n8455) );
  OR2_X1 U10895 ( .A1(n6471), .A2(n8455), .ZN(n8458) );
  INV_X1 U10896 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n8456) );
  OR2_X1 U10897 ( .A1(n6473), .A2(n8456), .ZN(n8457) );
  NAND2_X1 U10898 ( .A1(n8471), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8462) );
  XNOR2_X1 U10899 ( .A(n8462), .B(P3_IR_REG_12__SCAN_IN), .ZN(n11587) );
  XNOR2_X1 U10900 ( .A(n8464), .B(n8463), .ZN(n9727) );
  NAND2_X1 U10901 ( .A1(n9727), .A2(n8684), .ZN(n8466) );
  NAND2_X1 U10902 ( .A1(n8288), .A2(SI_12_), .ZN(n8465) );
  OAI211_X1 U10903 ( .C1(n6722), .C2(n11589), .A(n8466), .B(n8465), .ZN(n12232) );
  NAND2_X1 U10904 ( .A1(n14496), .A2(n12232), .ZN(n8759) );
  INV_X1 U10905 ( .A(n12232), .ZN(n12799) );
  NAND2_X1 U10906 ( .A1(n12455), .A2(n12799), .ZN(n8761) );
  NAND2_X1 U10907 ( .A1(n8759), .A2(n8761), .ZN(n12794) );
  INV_X1 U10908 ( .A(n12794), .ZN(n12792) );
  NAND2_X1 U10909 ( .A1(n12793), .A2(n12792), .ZN(n8467) );
  NAND2_X1 U10910 ( .A1(n8468), .A2(n10020), .ZN(n8469) );
  NAND2_X1 U10911 ( .A1(n8470), .A2(n8469), .ZN(n9744) );
  NAND2_X1 U10912 ( .A1(n9744), .A2(n8684), .ZN(n8475) );
  NOR2_X1 U10913 ( .A1(n8471), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n8492) );
  OR2_X1 U10914 ( .A1(n8492), .A2(n6724), .ZN(n8472) );
  XNOR2_X1 U10915 ( .A(n8472), .B(n8491), .ZN(n12469) );
  OAI22_X1 U10916 ( .A1(n8575), .A2(SI_13_), .B1(n12480), .B2(n6722), .ZN(
        n8473) );
  INV_X1 U10917 ( .A(n8473), .ZN(n8474) );
  NAND2_X1 U10918 ( .A1(n8475), .A2(n8474), .ZN(n12785) );
  INV_X1 U10919 ( .A(n12785), .ZN(n8486) );
  INV_X1 U10920 ( .A(n8476), .ZN(n8529) );
  OR2_X1 U10921 ( .A1(n8478), .A2(n8477), .ZN(n8479) );
  NAND2_X1 U10922 ( .A1(n8499), .A2(n8479), .ZN(n12786) );
  NAND2_X1 U10923 ( .A1(n6469), .A2(n12786), .ZN(n8485) );
  NAND2_X1 U10924 ( .A1(n8546), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8484) );
  INV_X1 U10925 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n8480) );
  OR2_X1 U10926 ( .A1(n6471), .A2(n8480), .ZN(n8483) );
  INV_X1 U10927 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n8481) );
  OR2_X1 U10928 ( .A1(n6473), .A2(n8481), .ZN(n8482) );
  AND2_X1 U10929 ( .A1(n8486), .A2(n12798), .ZN(n8766) );
  INV_X1 U10930 ( .A(n12798), .ZN(n12454) );
  NAND2_X1 U10931 ( .A1(n12785), .A2(n12454), .ZN(n8765) );
  OR2_X1 U10932 ( .A1(n8488), .A2(n8487), .ZN(n8489) );
  NAND2_X1 U10933 ( .A1(n8490), .A2(n8489), .ZN(n9771) );
  NAND2_X1 U10934 ( .A1(n9771), .A2(n8684), .ZN(n8498) );
  NAND2_X1 U10935 ( .A1(n8492), .A2(n8491), .ZN(n8508) );
  NAND2_X1 U10936 ( .A1(n8508), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8494) );
  INV_X1 U10937 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8493) );
  INV_X1 U10938 ( .A(n12494), .ZN(n8495) );
  OAI22_X1 U10939 ( .A1(n8575), .A2(SI_14_), .B1(n8495), .B2(n6722), .ZN(n8496) );
  INV_X1 U10940 ( .A(n8496), .ZN(n8497) );
  NAND2_X1 U10941 ( .A1(n8699), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8505) );
  NAND2_X1 U10942 ( .A1(n8499), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8500) );
  AND2_X1 U10943 ( .A1(n8513), .A2(n8500), .ZN(n14428) );
  INV_X1 U10944 ( .A(n14428), .ZN(n12776) );
  NAND2_X1 U10945 ( .A1(n6469), .A2(n12776), .ZN(n8504) );
  NAND2_X1 U10946 ( .A1(n8698), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8503) );
  NAND2_X1 U10947 ( .A1(n8546), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8502) );
  NAND4_X1 U10948 ( .A1(n8505), .A2(n8504), .A3(n8503), .A4(n8502), .ZN(n12781) );
  NAND2_X1 U10949 ( .A1(n14424), .A2(n12781), .ZN(n8770) );
  XNOR2_X1 U10950 ( .A(n8507), .B(n8506), .ZN(n9960) );
  NAND2_X1 U10951 ( .A1(n9960), .A2(n8684), .ZN(n8512) );
  OAI21_X1 U10952 ( .B1(n8508), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8509) );
  XNOR2_X1 U10953 ( .A(n8509), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12528) );
  OAI22_X1 U10954 ( .A1(n8575), .A2(n9961), .B1(n6722), .B2(n12540), .ZN(n8510) );
  INV_X1 U10955 ( .A(n8510), .ZN(n8511) );
  INV_X1 U10956 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12496) );
  OR2_X1 U10957 ( .A1(n6471), .A2(n12496), .ZN(n8518) );
  NAND2_X1 U10958 ( .A1(n8698), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8517) );
  NAND2_X1 U10959 ( .A1(n8513), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8514) );
  NAND2_X1 U10960 ( .A1(n8527), .A2(n8514), .ZN(n12758) );
  NAND2_X1 U10961 ( .A1(n6469), .A2(n12758), .ZN(n8516) );
  NAND2_X1 U10962 ( .A1(n8546), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8515) );
  NAND4_X1 U10963 ( .A1(n8518), .A2(n8517), .A3(n8516), .A4(n8515), .ZN(n12769) );
  XNOR2_X1 U10964 ( .A(n12875), .B(n12769), .ZN(n12754) );
  INV_X1 U10965 ( .A(n12769), .ZN(n8519) );
  NAND2_X1 U10966 ( .A1(n12875), .A2(n8519), .ZN(n8774) );
  NAND2_X1 U10967 ( .A1(n12757), .A2(n8774), .ZN(n12745) );
  XNOR2_X1 U10968 ( .A(n8521), .B(n8520), .ZN(n10022) );
  NAND2_X1 U10969 ( .A1(n10022), .A2(n8684), .ZN(n8526) );
  NAND2_X1 U10970 ( .A1(n8522), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8523) );
  XNOR2_X1 U10971 ( .A(n8523), .B(P3_IR_REG_16__SCAN_IN), .ZN(n14439) );
  OAI22_X1 U10972 ( .A1(n8575), .A2(n10023), .B1(n6722), .B2(n12538), .ZN(
        n8524) );
  INV_X1 U10973 ( .A(n8524), .ZN(n8525) );
  NAND2_X1 U10974 ( .A1(n8526), .A2(n8525), .ZN(n14434) );
  NAND2_X1 U10975 ( .A1(n8546), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U10976 ( .A1(n8527), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U10977 ( .A1(n8544), .A2(n8528), .ZN(n14435) );
  NAND2_X1 U10978 ( .A1(n6469), .A2(n14435), .ZN(n8532) );
  INV_X1 U10979 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12531) );
  OR2_X1 U10980 ( .A1(n6471), .A2(n12531), .ZN(n8531) );
  INV_X1 U10981 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12938) );
  OR2_X1 U10982 ( .A1(n6473), .A2(n12938), .ZN(n8530) );
  OR2_X1 U10983 ( .A1(n14434), .A2(n12439), .ZN(n8719) );
  NAND2_X1 U10984 ( .A1(n14434), .A2(n12439), .ZN(n12728) );
  NAND2_X1 U10985 ( .A1(n8719), .A2(n12728), .ZN(n12737) );
  INV_X1 U10986 ( .A(n12737), .ZN(n12744) );
  OR2_X1 U10987 ( .A1(n8535), .A2(n8534), .ZN(n8536) );
  NAND2_X1 U10988 ( .A1(n8537), .A2(n8536), .ZN(n10058) );
  OR2_X1 U10989 ( .A1(n10058), .A2(n8602), .ZN(n8543) );
  NAND2_X1 U10990 ( .A1(n8538), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8539) );
  MUX2_X1 U10991 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8539), .S(
        P3_IR_REG_17__SCAN_IN), .Z(n8540) );
  AND2_X1 U10992 ( .A1(n8540), .A2(n8572), .ZN(n14456) );
  OAI22_X1 U10993 ( .A1(n8575), .A2(n10059), .B1(n6722), .B2(n12543), .ZN(
        n8541) );
  INV_X1 U10994 ( .A(n8541), .ZN(n8542) );
  NAND2_X1 U10995 ( .A1(n8543), .A2(n8542), .ZN(n12867) );
  NAND2_X1 U10996 ( .A1(n8544), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U10997 ( .A1(n8562), .A2(n8545), .ZN(n12732) );
  NAND2_X1 U10998 ( .A1(n6469), .A2(n12732), .ZN(n8552) );
  NAND2_X1 U10999 ( .A1(n8546), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8551) );
  INV_X1 U11000 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n8547) );
  OR2_X1 U11001 ( .A1(n6471), .A2(n8547), .ZN(n8550) );
  INV_X1 U11002 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n8548) );
  OR2_X1 U11003 ( .A1(n6473), .A2(n8548), .ZN(n8549) );
  XNOR2_X1 U11004 ( .A(n12867), .B(n12715), .ZN(n12729) );
  INV_X1 U11005 ( .A(n12729), .ZN(n12724) );
  NAND2_X1 U11006 ( .A1(n12867), .A2(n12715), .ZN(n8781) );
  OR2_X1 U11007 ( .A1(n8555), .A2(n8554), .ZN(n8556) );
  NAND2_X1 U11008 ( .A1(n8557), .A2(n8556), .ZN(n10097) );
  OR2_X1 U11009 ( .A1(n10097), .A2(n8602), .ZN(n8561) );
  NAND2_X1 U11010 ( .A1(n8572), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8558) );
  XNOR2_X1 U11011 ( .A(n8558), .B(P3_IR_REG_18__SCAN_IN), .ZN(n14470) );
  OAI22_X1 U11012 ( .A1(n8575), .A2(n10098), .B1(n6722), .B2(n12546), .ZN(
        n8559) );
  INV_X1 U11013 ( .A(n8559), .ZN(n8560) );
  NAND2_X1 U11014 ( .A1(n8561), .A2(n8560), .ZN(n12407) );
  NAND2_X1 U11015 ( .A1(n8546), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8567) );
  NAND2_X1 U11016 ( .A1(n8562), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8563) );
  NAND2_X1 U11017 ( .A1(n8579), .A2(n8563), .ZN(n12719) );
  NAND2_X1 U11018 ( .A1(n6469), .A2(n12719), .ZN(n8566) );
  INV_X1 U11019 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12534) );
  OR2_X1 U11020 ( .A1(n6471), .A2(n12534), .ZN(n8565) );
  INV_X1 U11021 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12933) );
  OR2_X1 U11022 ( .A1(n6473), .A2(n12933), .ZN(n8564) );
  OR2_X1 U11023 ( .A1(n12407), .A2(n12322), .ZN(n8780) );
  NAND2_X1 U11024 ( .A1(n12407), .A2(n12322), .ZN(n8782) );
  OR2_X1 U11025 ( .A1(n8569), .A2(n8568), .ZN(n8570) );
  NAND2_X1 U11026 ( .A1(n8571), .A2(n8570), .ZN(n10110) );
  NAND2_X1 U11027 ( .A1(n10110), .A2(n8684), .ZN(n8578) );
  INV_X1 U11028 ( .A(n8710), .ZN(n8573) );
  NAND2_X1 U11029 ( .A1(n8573), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8574) );
  OAI22_X1 U11030 ( .A1(n8575), .A2(SI_19_), .B1(n12550), .B2(n6722), .ZN(
        n8576) );
  INV_X1 U11031 ( .A(n8576), .ZN(n8577) );
  NAND2_X1 U11032 ( .A1(n8699), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8584) );
  NAND2_X1 U11033 ( .A1(n8698), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8583) );
  NAND2_X1 U11034 ( .A1(n8579), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8580) );
  NAND2_X1 U11035 ( .A1(n8592), .A2(n8580), .ZN(n12705) );
  NAND2_X1 U11036 ( .A1(n6469), .A2(n12705), .ZN(n8582) );
  NAND2_X1 U11037 ( .A1(n8546), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8581) );
  NAND4_X1 U11038 ( .A1(n8584), .A2(n8583), .A3(n8582), .A4(n8581), .ZN(n12453) );
  NAND2_X1 U11039 ( .A1(n12931), .A2(n12453), .ZN(n8823) );
  OR2_X1 U11040 ( .A1(n12931), .A2(n12453), .ZN(n8824) );
  NAND2_X1 U11041 ( .A1(n8587), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U11042 ( .A1(n8589), .A2(n8588), .ZN(n10565) );
  OR2_X1 U11043 ( .A1(n10565), .A2(n8602), .ZN(n8591) );
  NAND2_X1 U11044 ( .A1(n8288), .A2(SI_20_), .ZN(n8590) );
  NAND2_X1 U11045 ( .A1(n8546), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U11046 ( .A1(n8592), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8593) );
  NAND2_X1 U11047 ( .A1(n8605), .A2(n8593), .ZN(n12686) );
  NAND2_X1 U11048 ( .A1(n6469), .A2(n12686), .ZN(n8596) );
  INV_X1 U11049 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12688) );
  OR2_X1 U11050 ( .A1(n6471), .A2(n12688), .ZN(n8595) );
  INV_X1 U11051 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12925) );
  OR2_X1 U11052 ( .A1(n6473), .A2(n12925), .ZN(n8594) );
  XNOR2_X1 U11053 ( .A(n12694), .B(n12704), .ZN(n12689) );
  OR2_X1 U11054 ( .A1(n12694), .A2(n12704), .ZN(n8786) );
  OR2_X1 U11055 ( .A1(n8599), .A2(n8598), .ZN(n8600) );
  NAND2_X1 U11056 ( .A1(n8601), .A2(n8600), .ZN(n10616) );
  OR2_X1 U11057 ( .A1(n10616), .A2(n8602), .ZN(n8604) );
  NAND2_X1 U11058 ( .A1(n8288), .A2(SI_21_), .ZN(n8603) );
  NAND2_X1 U11059 ( .A1(n8546), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8612) );
  NAND2_X1 U11060 ( .A1(n8605), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8606) );
  NAND2_X1 U11061 ( .A1(n8618), .A2(n8606), .ZN(n12678) );
  NAND2_X1 U11062 ( .A1(n6469), .A2(n12678), .ZN(n8611) );
  INV_X1 U11063 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n8607) );
  OR2_X1 U11064 ( .A1(n6471), .A2(n8607), .ZN(n8610) );
  INV_X1 U11065 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12921) );
  OR2_X1 U11066 ( .A1(n6473), .A2(n12921), .ZN(n8609) );
  NAND2_X1 U11067 ( .A1(n12677), .A2(n12685), .ZN(n8792) );
  XNOR2_X1 U11068 ( .A(n8615), .B(n8614), .ZN(n10729) );
  NAND2_X1 U11069 ( .A1(n10729), .A2(n8684), .ZN(n8617) );
  NAND2_X1 U11070 ( .A1(n8288), .A2(SI_22_), .ZN(n8616) );
  NAND2_X1 U11071 ( .A1(n8618), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8619) );
  NAND2_X1 U11072 ( .A1(n8628), .A2(n8619), .ZN(n12665) );
  NAND2_X1 U11073 ( .A1(n12665), .A2(n6469), .ZN(n8623) );
  NAND2_X1 U11074 ( .A1(n8546), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8622) );
  NAND2_X1 U11075 ( .A1(n8699), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8621) );
  NAND2_X1 U11076 ( .A1(n8698), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8620) );
  NAND4_X1 U11077 ( .A1(n8623), .A2(n8622), .A3(n8621), .A4(n8620), .ZN(n12450) );
  NAND2_X1 U11078 ( .A1(n12664), .A2(n12676), .ZN(n12640) );
  XNOR2_X1 U11079 ( .A(n8625), .B(n8624), .ZN(n10885) );
  NAND2_X1 U11080 ( .A1(n10885), .A2(n8684), .ZN(n8627) );
  NAND2_X1 U11081 ( .A1(n8288), .A2(SI_23_), .ZN(n8626) );
  INV_X1 U11082 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12913) );
  NAND2_X1 U11083 ( .A1(n8628), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U11084 ( .A1(n8637), .A2(n8629), .ZN(n12313) );
  NAND2_X1 U11085 ( .A1(n12313), .A2(n6469), .ZN(n8631) );
  AOI22_X1 U11086 ( .A1(n8546), .A2(P3_REG1_REG_23__SCAN_IN), .B1(n8699), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n8630) );
  XNOR2_X1 U11087 ( .A(n12654), .B(n12449), .ZN(n12643) );
  AND2_X1 U11088 ( .A1(n12640), .A2(n12643), .ZN(n8632) );
  NAND2_X1 U11089 ( .A1(n12639), .A2(n8632), .ZN(n12627) );
  INV_X1 U11090 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8633) );
  XNOR2_X1 U11091 ( .A(n8634), .B(n8633), .ZN(n11261) );
  NAND2_X1 U11092 ( .A1(n11261), .A2(n8684), .ZN(n8636) );
  NAND2_X1 U11093 ( .A1(n8288), .A2(SI_24_), .ZN(n8635) );
  NAND2_X1 U11094 ( .A1(n8637), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U11095 ( .A1(n8648), .A2(n8638), .ZN(n12634) );
  NAND2_X1 U11096 ( .A1(n12634), .A2(n6469), .ZN(n8641) );
  AOI22_X1 U11097 ( .A1(n8546), .A2(P3_REG1_REG_24__SCAN_IN), .B1(n8699), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n8640) );
  NAND2_X1 U11098 ( .A1(n8698), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8639) );
  NAND2_X1 U11099 ( .A1(n12909), .A2(n12364), .ZN(n8799) );
  OR2_X1 U11100 ( .A1(n12909), .A2(n12364), .ZN(n8642) );
  NAND2_X1 U11101 ( .A1(n8799), .A2(n8642), .ZN(n12630) );
  INV_X1 U11102 ( .A(n12449), .ZN(n12401) );
  NOR2_X1 U11103 ( .A1(n12654), .A2(n12401), .ZN(n12628) );
  NOR2_X1 U11104 ( .A1(n12630), .A2(n12628), .ZN(n8798) );
  OR2_X1 U11105 ( .A1(n7401), .A2(n12641), .ZN(n12626) );
  AND2_X1 U11106 ( .A1(n8798), .A2(n12626), .ZN(n8643) );
  NAND2_X1 U11107 ( .A1(n12627), .A2(n8643), .ZN(n12632) );
  XNOR2_X1 U11108 ( .A(n8645), .B(n8644), .ZN(n11366) );
  NAND2_X1 U11109 ( .A1(n11366), .A2(n8684), .ZN(n8647) );
  NAND2_X1 U11110 ( .A1(n8288), .A2(SI_25_), .ZN(n8646) );
  NAND2_X1 U11111 ( .A1(n8648), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8649) );
  NAND2_X1 U11112 ( .A1(n8661), .A2(n8649), .ZN(n12616) );
  NAND2_X1 U11113 ( .A1(n12616), .A2(n6469), .ZN(n8656) );
  INV_X1 U11114 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U11115 ( .A1(n8546), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8652) );
  NAND2_X1 U11116 ( .A1(n8699), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8651) );
  OAI211_X1 U11117 ( .C1(n8653), .C2(n6473), .A(n8652), .B(n8651), .ZN(n8654)
         );
  INV_X1 U11118 ( .A(n8654), .ZN(n8655) );
  OR2_X1 U11119 ( .A1(n12829), .A2(n12597), .ZN(n8803) );
  NAND2_X1 U11120 ( .A1(n12829), .A2(n12597), .ZN(n12599) );
  NAND2_X1 U11121 ( .A1(n8803), .A2(n12599), .ZN(n12609) );
  INV_X1 U11122 ( .A(n12609), .ZN(n12614) );
  XNOR2_X1 U11123 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .ZN(n8657) );
  XNOR2_X1 U11124 ( .A(n8658), .B(n8657), .ZN(n11496) );
  NAND2_X1 U11125 ( .A1(n11496), .A2(n8684), .ZN(n8660) );
  NAND2_X1 U11126 ( .A1(n8288), .A2(SI_26_), .ZN(n8659) );
  NAND2_X1 U11127 ( .A1(n8661), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8662) );
  NAND2_X1 U11128 ( .A1(n8674), .A2(n8662), .ZN(n12603) );
  NAND2_X1 U11129 ( .A1(n12603), .A2(n6469), .ZN(n8667) );
  INV_X1 U11130 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12903) );
  NAND2_X1 U11131 ( .A1(n8546), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8664) );
  NAND2_X1 U11132 ( .A1(n8699), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8663) );
  OAI211_X1 U11133 ( .C1(n12903), .C2(n6473), .A(n8664), .B(n8663), .ZN(n8665)
         );
  INV_X1 U11134 ( .A(n8665), .ZN(n8666) );
  NAND2_X1 U11135 ( .A1(n12602), .A2(n12584), .ZN(n8807) );
  AND2_X1 U11136 ( .A1(n12599), .A2(n8807), .ZN(n8669) );
  XNOR2_X1 U11137 ( .A(n13590), .B(P2_DATAO_REG_27__SCAN_IN), .ZN(n8670) );
  XNOR2_X1 U11138 ( .A(n8671), .B(n8670), .ZN(n11558) );
  NAND2_X1 U11139 ( .A1(n11558), .A2(n8684), .ZN(n8673) );
  NAND2_X1 U11140 ( .A1(n8288), .A2(SI_27_), .ZN(n8672) );
  NAND2_X1 U11141 ( .A1(n8674), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U11142 ( .A1(n8687), .A2(n8675), .ZN(n12590) );
  NAND2_X1 U11143 ( .A1(n12590), .A2(n6469), .ZN(n8681) );
  INV_X1 U11144 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12899) );
  NAND2_X1 U11145 ( .A1(n8699), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8677) );
  NAND2_X1 U11146 ( .A1(n8546), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8676) );
  OAI211_X1 U11147 ( .C1(n12899), .C2(n6473), .A(n8677), .B(n8676), .ZN(n8679)
         );
  INV_X1 U11148 ( .A(n8679), .ZN(n8680) );
  OR2_X1 U11149 ( .A1(n12589), .A2(n12598), .ZN(n8812) );
  NAND2_X1 U11150 ( .A1(n12589), .A2(n12598), .ZN(n8813) );
  XNOR2_X1 U11151 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .ZN(n8682) );
  NAND2_X1 U11152 ( .A1(n12961), .A2(n8684), .ZN(n8686) );
  NAND2_X1 U11153 ( .A1(n8288), .A2(SI_28_), .ZN(n8685) );
  NAND2_X1 U11154 ( .A1(n8687), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8688) );
  NAND2_X1 U11155 ( .A1(n8689), .A2(n8688), .ZN(n12577) );
  INV_X1 U11156 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12896) );
  NAND2_X1 U11157 ( .A1(n8699), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U11158 ( .A1(n8546), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8690) );
  OAI211_X1 U11159 ( .C1(n12896), .C2(n6473), .A(n8691), .B(n8690), .ZN(n8692)
         );
  AOI21_X1 U11160 ( .B1(n12577), .B2(n6469), .A(n8692), .ZN(n12585) );
  NAND2_X1 U11161 ( .A1(n12576), .A2(n12585), .ZN(n8814) );
  INV_X1 U11162 ( .A(n8811), .ZN(n8816) );
  NAND2_X1 U11163 ( .A1(n8288), .A2(SI_29_), .ZN(n8697) );
  INV_X1 U11164 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n12815) );
  NAND2_X1 U11165 ( .A1(n8698), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8701) );
  NAND2_X1 U11166 ( .A1(n8699), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8700) );
  OAI211_X1 U11167 ( .C1(n12815), .C2(n8437), .A(n8701), .B(n8700), .ZN(n8702)
         );
  INV_X1 U11168 ( .A(n8702), .ZN(n8703) );
  NAND2_X1 U11169 ( .A1(n8704), .A2(n8703), .ZN(n12570) );
  NAND2_X1 U11170 ( .A1(n8706), .A2(n12259), .ZN(n8705) );
  INV_X1 U11171 ( .A(n12560), .ZN(n12444) );
  INV_X1 U11172 ( .A(n12570), .ZN(n8707) );
  NAND2_X1 U11173 ( .A1(n12894), .A2(n8707), .ZN(n8821) );
  OAI21_X1 U11174 ( .B1(n12890), .B2(n12444), .A(n8821), .ZN(n8708) );
  NAND2_X1 U11175 ( .A1(n8715), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8717) );
  NAND2_X1 U11176 ( .A1(n10944), .A2(n10638), .ZN(n10929) );
  INV_X1 U11177 ( .A(n8719), .ZN(n8778) );
  MUX2_X1 U11178 ( .A(n15241), .B(n14955), .S(n10640), .Z(n8753) );
  INV_X1 U11179 ( .A(n10935), .ZN(n10733) );
  OAI21_X1 U11180 ( .B1(n8825), .B2(n10614), .A(n10640), .ZN(n8722) );
  INV_X1 U11181 ( .A(n8825), .ZN(n8720) );
  NAND3_X1 U11182 ( .A1(n8826), .A2(n8720), .A3(n10730), .ZN(n8721) );
  NAND3_X1 U11183 ( .A1(n8725), .A2(n15190), .A3(n8826), .ZN(n8724) );
  AND3_X1 U11184 ( .A1(n8724), .A2(n8727), .A3(n8723), .ZN(n8729) );
  NOR3_X1 U11185 ( .A1(n15186), .A2(n11327), .A3(n9650), .ZN(n8730) );
  NOR2_X1 U11186 ( .A1(n9534), .A2(n9650), .ZN(n8733) );
  NOR2_X1 U11187 ( .A1(n15223), .A2(n10640), .ZN(n8732) );
  MUX2_X1 U11188 ( .A(n8733), .B(n8732), .S(n12460), .Z(n8734) );
  NOR3_X1 U11189 ( .A1(n8735), .A2(n8734), .A3(n15161), .ZN(n8744) );
  NAND2_X1 U11190 ( .A1(n8741), .A2(n8736), .ZN(n8739) );
  NAND2_X1 U11191 ( .A1(n8740), .A2(n8737), .ZN(n8738) );
  MUX2_X1 U11192 ( .A(n8739), .B(n8738), .S(n9650), .Z(n8743) );
  MUX2_X1 U11193 ( .A(n8741), .B(n8740), .S(n10640), .Z(n8742) );
  MUX2_X1 U11194 ( .A(n8746), .B(n8745), .S(n9650), .Z(n8747) );
  MUX2_X1 U11195 ( .A(n8750), .B(n8749), .S(n10640), .Z(n8751) );
  OAI21_X1 U11196 ( .B1(n8754), .B2(n15083), .A(n14493), .ZN(n8760) );
  INV_X1 U11197 ( .A(n8760), .ZN(n8756) );
  INV_X1 U11198 ( .A(n8757), .ZN(n14489) );
  OAI211_X1 U11199 ( .C1(n8760), .C2(n14489), .A(n8759), .B(n8758), .ZN(n8762)
         );
  NAND2_X1 U11200 ( .A1(n8762), .A2(n8761), .ZN(n8763) );
  INV_X1 U11201 ( .A(n8765), .ZN(n8767) );
  MUX2_X1 U11202 ( .A(n8767), .B(n8766), .S(n9650), .Z(n8768) );
  MUX2_X1 U11203 ( .A(n8770), .B(n12755), .S(n10640), .Z(n8771) );
  NAND2_X1 U11204 ( .A1(n12754), .A2(n8771), .ZN(n8773) );
  INV_X1 U11205 ( .A(n12875), .ZN(n12760) );
  AOI21_X1 U11206 ( .B1(n12760), .B2(n12769), .A(n8778), .ZN(n8772) );
  AOI21_X1 U11207 ( .B1(n12728), .B2(n8774), .A(n10640), .ZN(n8775) );
  AOI21_X1 U11208 ( .B1(n8776), .B2(n12728), .A(n8775), .ZN(n8777) );
  INV_X1 U11209 ( .A(n12867), .ZN(n12734) );
  NAND3_X1 U11210 ( .A1(n8782), .A2(n12734), .A3(n12739), .ZN(n8779) );
  NAND3_X1 U11211 ( .A1(n8824), .A2(n8782), .A3(n10640), .ZN(n8783) );
  AOI22_X1 U11212 ( .A1(n8784), .A2(n12713), .B1(n6588), .B2(n8783), .ZN(n8790) );
  INV_X1 U11213 ( .A(n12689), .ZN(n8836) );
  MUX2_X1 U11214 ( .A(n8823), .B(n8824), .S(n9650), .Z(n8785) );
  NAND2_X1 U11215 ( .A1(n8836), .A2(n8785), .ZN(n8789) );
  NAND2_X1 U11216 ( .A1(n12694), .A2(n12704), .ZN(n8787) );
  MUX2_X1 U11217 ( .A(n8787), .B(n8786), .S(n9650), .Z(n8788) );
  MUX2_X1 U11218 ( .A(n8792), .B(n8791), .S(n10640), .Z(n8793) );
  INV_X1 U11219 ( .A(n12630), .ZN(n8795) );
  MUX2_X1 U11220 ( .A(n12640), .B(n12641), .S(n9650), .Z(n8794) );
  INV_X1 U11221 ( .A(n8798), .ZN(n8802) );
  XNOR2_X1 U11222 ( .A(n8799), .B(n10640), .ZN(n8801) );
  INV_X1 U11223 ( .A(n12654), .ZN(n12915) );
  NOR4_X1 U11224 ( .A1(n12630), .A2(n12915), .A3(n12449), .A4(n10640), .ZN(
        n8800) );
  AOI21_X1 U11225 ( .B1(n8802), .B2(n8801), .A(n8800), .ZN(n8805) );
  MUX2_X1 U11226 ( .A(n12599), .B(n8803), .S(n10640), .Z(n8804) );
  OAI21_X1 U11227 ( .B1(n8805), .B2(n12609), .A(n8804), .ZN(n8809) );
  MUX2_X1 U11228 ( .A(n8807), .B(n8806), .S(n9650), .Z(n8808) );
  AND2_X2 U11229 ( .A1(n8811), .A2(n8814), .ZN(n12565) );
  INV_X1 U11230 ( .A(n8842), .ZN(n8817) );
  NAND3_X1 U11231 ( .A1(n8818), .A2(n8822), .A3(n8817), .ZN(n8820) );
  INV_X1 U11232 ( .A(n15199), .ZN(n10946) );
  NAND2_X1 U11233 ( .A1(n8822), .A2(n8821), .ZN(n12264) );
  INV_X1 U11234 ( .A(n12658), .ZN(n12663) );
  NAND2_X1 U11235 ( .A1(n8824), .A2(n8823), .ZN(n12700) );
  NOR2_X1 U11236 ( .A1(n10935), .A2(n8825), .ZN(n10602) );
  NAND4_X1 U11237 ( .A1(n10602), .A2(n11046), .A3(n15138), .A4(n15110), .ZN(
        n8829) );
  INV_X1 U11238 ( .A(n10936), .ZN(n8827) );
  NAND3_X1 U11239 ( .A1(n8827), .A2(n15121), .A3(n12217), .ZN(n8828) );
  NOR2_X1 U11240 ( .A1(n8829), .A2(n8828), .ZN(n8831) );
  AND3_X1 U11241 ( .A1(n7384), .A2(n7396), .A3(n15094), .ZN(n8830) );
  AND4_X1 U11242 ( .A1(n8831), .A2(n15190), .A3(n12792), .A4(n8830), .ZN(n8832) );
  NAND4_X1 U11243 ( .A1(n8832), .A2(n12765), .A3(n14493), .A4(n7489), .ZN(
        n8833) );
  NOR2_X1 U11244 ( .A1(n12737), .A2(n8833), .ZN(n8834) );
  NAND4_X1 U11245 ( .A1(n12713), .A2(n8834), .A3(n12724), .A4(n12754), .ZN(
        n8835) );
  NOR2_X1 U11246 ( .A1(n12700), .A2(n8835), .ZN(n8837) );
  NAND3_X1 U11247 ( .A1(n12674), .A2(n8837), .A3(n8836), .ZN(n8838) );
  OR4_X1 U11248 ( .A1(n12630), .A2(n7401), .A3(n12663), .A4(n8838), .ZN(n8839)
         );
  NOR2_X1 U11249 ( .A1(n12609), .A2(n8839), .ZN(n8840) );
  NAND3_X1 U11250 ( .A1(n12587), .A2(n12600), .A3(n8840), .ZN(n8841) );
  OR2_X1 U11251 ( .A1(n9649), .A2(P3_U3151), .ZN(n10886) );
  INV_X1 U11252 ( .A(n12962), .ZN(n12257) );
  NAND2_X1 U11253 ( .A1(n12257), .A2(n9659), .ZN(n9657) );
  NAND2_X1 U11254 ( .A1(n8853), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8854) );
  MUX2_X1 U11255 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8854), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8855) );
  NAND2_X1 U11256 ( .A1(n8855), .A2(n6734), .ZN(n11264) );
  INV_X1 U11257 ( .A(n11264), .ZN(n8859) );
  NAND2_X1 U11258 ( .A1(n6734), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8856) );
  MUX2_X1 U11259 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8856), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8857) );
  INV_X1 U11260 ( .A(n11368), .ZN(n8858) );
  NAND4_X1 U11261 ( .A1(n15145), .A2(n10937), .A3(n12257), .A4(n10866), .ZN(
        n8860) );
  OAI211_X1 U11262 ( .C1(n10730), .C2(n10886), .A(n8860), .B(P3_B_REG_SCAN_IN), 
        .ZN(n8861) );
  NOR2_X1 U11263 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n8866) );
  NOR2_X2 U11264 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n8865) );
  NOR2_X2 U11265 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), 
        .ZN(n8864) );
  AND4_X2 U11266 ( .A1(n8866), .A2(n8865), .A3(n8864), .A4(n8863), .ZN(n8871)
         );
  NOR2_X2 U11267 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n8869) );
  NOR2_X2 U11268 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8868) );
  NOR2_X2 U11269 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8867) );
  AND3_X2 U11270 ( .A1(n8869), .A2(n8868), .A3(n8867), .ZN(n9123) );
  NAND3_X2 U11271 ( .A1(n8871), .A2(n9123), .A3(n8946), .ZN(n9194) );
  NOR2_X1 U11272 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n8874) );
  NAND4_X1 U11273 ( .A1(n8874), .A2(n8873), .A3(n8872), .A4(n8906), .ZN(n9494)
         );
  INV_X1 U11274 ( .A(n9494), .ZN(n8877) );
  NAND2_X1 U11275 ( .A1(n8877), .A2(n7480), .ZN(n8878) );
  NAND2_X1 U11276 ( .A1(n8903), .A2(n8880), .ZN(n8885) );
  INV_X1 U11277 ( .A(n8885), .ZN(n8882) );
  NAND2_X1 U11278 ( .A1(n8882), .A2(n8881), .ZN(n8887) );
  NAND2_X1 U11279 ( .A1(n8885), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8886) );
  AND2_X2 U11280 ( .A1(n8889), .A2(n13581), .ZN(n9251) );
  NAND2_X1 U11281 ( .A1(n9251), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8894) );
  AND2_X4 U11282 ( .A1(n8889), .A2(n8890), .ZN(n9005) );
  NAND2_X1 U11283 ( .A1(n9005), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8893) );
  AND2_X4 U11284 ( .A1(n13577), .A2(n8890), .ZN(n9006) );
  NAND2_X1 U11285 ( .A1(n9006), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8892) );
  AND2_X2 U11286 ( .A1(n13577), .A2(n13581), .ZN(n9011) );
  NAND2_X1 U11287 ( .A1(n9011), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8891) );
  INV_X1 U11288 ( .A(n9472), .ZN(n10216) );
  INV_X1 U11289 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9840) );
  NAND2_X1 U11290 ( .A1(n9685), .A2(SI_0_), .ZN(n8896) );
  NAND2_X1 U11291 ( .A1(n8896), .A2(n8895), .ZN(n8898) );
  NAND2_X1 U11292 ( .A1(n8898), .A2(n8897), .ZN(n13602) );
  NAND2_X2 U11293 ( .A1(n8900), .A2(n6463), .ZN(n10217) );
  MUX2_X1 U11294 ( .A(n9840), .B(n13602), .S(n9832), .Z(n14858) );
  NAND2_X1 U11295 ( .A1(n10216), .A2(n14858), .ZN(n9473) );
  NOR2_X2 U11296 ( .A1(n9194), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n9212) );
  NAND2_X1 U11297 ( .A1(n9212), .A2(n8905), .ZN(n9232) );
  XNOR2_X2 U11298 ( .A(n8911), .B(n8910), .ZN(n8923) );
  INV_X1 U11299 ( .A(n8912), .ZN(n8913) );
  NAND2_X1 U11300 ( .A1(n9441), .A2(n9468), .ZN(n10666) );
  NAND2_X1 U11301 ( .A1(n8915), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8916) );
  INV_X1 U11302 ( .A(n8917), .ZN(n9464) );
  OR2_X4 U11303 ( .A1(n10666), .A2(n6618), .ZN(n9406) );
  NAND2_X1 U11304 ( .A1(n9472), .A2(n9406), .ZN(n8927) );
  INV_X1 U11305 ( .A(n14858), .ZN(n8919) );
  NAND2_X1 U11306 ( .A1(n8965), .A2(n8919), .ZN(n8920) );
  NAND3_X1 U11307 ( .A1(n9473), .A2(n8927), .A3(n8920), .ZN(n8926) );
  NAND2_X1 U11308 ( .A1(n9442), .A2(n8923), .ZN(n10774) );
  INV_X1 U11309 ( .A(n10774), .ZN(n8924) );
  OAI21_X1 U11310 ( .B1(n8921), .B2(n13213), .A(n8924), .ZN(n8925) );
  NAND2_X1 U11311 ( .A1(n8926), .A2(n8925), .ZN(n8930) );
  INV_X1 U11312 ( .A(n8927), .ZN(n8928) );
  NAND2_X1 U11313 ( .A1(n8928), .A2(n14858), .ZN(n8929) );
  INV_X1 U11314 ( .A(n9840), .ZN(n14767) );
  NAND2_X1 U11315 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n14767), .ZN(n8931) );
  MUX2_X1 U11316 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8931), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8934) );
  INV_X1 U11317 ( .A(n8932), .ZN(n8933) );
  NAND2_X1 U11318 ( .A1(n8934), .A2(n8933), .ZN(n9857) );
  INV_X1 U11319 ( .A(n9857), .ZN(n9859) );
  OR2_X1 U11320 ( .A1(n9406), .A2(n14895), .ZN(n8940) );
  NAND2_X1 U11321 ( .A1(n9006), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8938) );
  NAND2_X1 U11322 ( .A1(n9005), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8937) );
  NAND2_X1 U11323 ( .A1(n9011), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8936) );
  NAND2_X1 U11324 ( .A1(n9251), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8935) );
  NAND2_X1 U11325 ( .A1(n13182), .A2(n9406), .ZN(n8939) );
  NAND2_X1 U11326 ( .A1(n8940), .A2(n8939), .ZN(n8953) );
  NAND2_X1 U11327 ( .A1(n9006), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8944) );
  NAND2_X1 U11328 ( .A1(n9005), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8943) );
  NAND2_X1 U11329 ( .A1(n9425), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8942) );
  NAND2_X1 U11330 ( .A1(n9251), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8941) );
  NAND2_X1 U11331 ( .A1(n9437), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8949) );
  NOR2_X1 U11332 ( .A1(n8932), .A2(n13573), .ZN(n8945) );
  MUX2_X1 U11333 ( .A(n13573), .B(n8945), .S(P2_IR_REG_2__SCAN_IN), .Z(n8947)
         );
  NAND2_X1 U11334 ( .A1(n9244), .A2(n14787), .ZN(n8948) );
  NAND2_X1 U11336 ( .A1(n8951), .A2(n8950), .ZN(n8955) );
  OAI22_X1 U11337 ( .A1(n8954), .A2(n8953), .B1(n8956), .B2(n8955), .ZN(n8975)
         );
  AOI21_X1 U11338 ( .B1(n8954), .B2(n8953), .A(n8952), .ZN(n8974) );
  NAND2_X1 U11339 ( .A1(n7206), .A2(n9672), .ZN(n8963) );
  NOR2_X1 U11340 ( .A1(n8959), .A2(n13573), .ZN(n8957) );
  MUX2_X1 U11341 ( .A(n13573), .B(n8957), .S(P2_IR_REG_3__SCAN_IN), .Z(n8961)
         );
  INV_X1 U11342 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8958) );
  NAND2_X1 U11343 ( .A1(n8959), .A2(n8958), .ZN(n8998) );
  INV_X1 U11344 ( .A(n8998), .ZN(n8960) );
  NAND2_X1 U11345 ( .A1(n9244), .A2(n9863), .ZN(n8962) );
  INV_X1 U11346 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8980) );
  NAND2_X1 U11347 ( .A1(n9006), .A2(n8980), .ZN(n8969) );
  NAND2_X1 U11348 ( .A1(n9005), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8968) );
  NAND2_X1 U11349 ( .A1(n9011), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8967) );
  NAND2_X1 U11350 ( .A1(n9251), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8966) );
  NAND4_X1 U11351 ( .A1(n8969), .A2(n8968), .A3(n8967), .A4(n8966), .ZN(n13180) );
  NAND2_X1 U11352 ( .A1(n13180), .A2(n9406), .ZN(n8970) );
  NAND2_X1 U11353 ( .A1(n8971), .A2(n8970), .ZN(n8987) );
  NAND2_X1 U11354 ( .A1(n8987), .A2(n8988), .ZN(n8972) );
  OAI211_X1 U11355 ( .C1(n8975), .C2(n8974), .A(n8973), .B(n8972), .ZN(n8993)
         );
  NAND2_X1 U11356 ( .A1(n9676), .A2(n7206), .ZN(n8978) );
  NAND2_X1 U11357 ( .A1(n8998), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8976) );
  XNOR2_X1 U11358 ( .A(n8976), .B(P2_IR_REG_4__SCAN_IN), .ZN(n9937) );
  AOI22_X1 U11359 ( .A1(n9437), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n9244), .B2(
        n9937), .ZN(n8977) );
  NAND2_X1 U11360 ( .A1(n9005), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8985) );
  INV_X1 U11361 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8979) );
  NAND2_X1 U11362 ( .A1(n8980), .A2(n8979), .ZN(n8981) );
  NAND2_X1 U11363 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9009) );
  AND2_X1 U11364 ( .A1(n8981), .A2(n9009), .ZN(n14845) );
  NAND2_X1 U11365 ( .A1(n9006), .A2(n14845), .ZN(n8984) );
  NAND2_X1 U11366 ( .A1(n9251), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8983) );
  NAND2_X1 U11367 ( .A1(n9443), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8982) );
  NAND4_X1 U11368 ( .A1(n8985), .A2(n8984), .A3(n8983), .A4(n8982), .ZN(n13179) );
  NAND2_X1 U11369 ( .A1(n13179), .A2(n9118), .ZN(n8986) );
  INV_X1 U11370 ( .A(n9406), .ZN(n9057) );
  AOI22_X1 U11371 ( .A1(n9057), .A2(n13179), .B1(n9406), .B2(n14850), .ZN(
        n8995) );
  OR2_X1 U11372 ( .A1(n8994), .A2(n8995), .ZN(n8992) );
  INV_X1 U11373 ( .A(n8987), .ZN(n8990) );
  INV_X1 U11374 ( .A(n8988), .ZN(n8989) );
  NAND2_X1 U11375 ( .A1(n8990), .A2(n8989), .ZN(n8991) );
  NAND3_X1 U11376 ( .A1(n8993), .A2(n8992), .A3(n8991), .ZN(n8997) );
  NAND2_X1 U11377 ( .A1(n8995), .A2(n8994), .ZN(n8996) );
  NAND2_X1 U11378 ( .A1(n8997), .A2(n8996), .ZN(n9034) );
  NAND2_X1 U11379 ( .A1(n9681), .A2(n9436), .ZN(n9004) );
  NOR2_X1 U11380 ( .A1(n8998), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n9001) );
  OR2_X1 U11381 ( .A1(n9001), .A2(n13573), .ZN(n8999) );
  MUX2_X1 U11382 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8999), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n9002) );
  NAND2_X1 U11383 ( .A1(n9001), .A2(n9000), .ZN(n9125) );
  AND2_X1 U11384 ( .A1(n9002), .A2(n9125), .ZN(n14817) );
  AOI22_X1 U11385 ( .A1(n9437), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9244), .B2(
        n14817), .ZN(n9003) );
  NAND2_X1 U11386 ( .A1(n9004), .A2(n9003), .ZN(n13087) );
  NAND2_X1 U11387 ( .A1(n6478), .A2(n13087), .ZN(n9017) );
  NAND2_X1 U11388 ( .A1(n9005), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9015) );
  INV_X1 U11389 ( .A(n9009), .ZN(n9007) );
  INV_X1 U11390 ( .A(n9021), .ZN(n9023) );
  INV_X1 U11391 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9008) );
  NAND2_X1 U11392 ( .A1(n9009), .A2(n9008), .ZN(n9010) );
  AND2_X1 U11393 ( .A1(n9023), .A2(n9010), .ZN(n13086) );
  NAND2_X1 U11394 ( .A1(n9006), .A2(n13086), .ZN(n9014) );
  NAND2_X1 U11395 ( .A1(n9426), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9013) );
  INV_X2 U11396 ( .A(n9011), .ZN(n9025) );
  INV_X2 U11397 ( .A(n9025), .ZN(n9425) );
  NAND2_X1 U11398 ( .A1(n9425), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9012) );
  NAND4_X1 U11399 ( .A1(n9015), .A2(n9014), .A3(n9013), .A4(n9012), .ZN(n13178) );
  NAND2_X1 U11400 ( .A1(n13178), .A2(n9449), .ZN(n9016) );
  NAND2_X1 U11401 ( .A1(n9017), .A2(n9016), .ZN(n9033) );
  NAND2_X1 U11402 ( .A1(n9699), .A2(n9436), .ZN(n9020) );
  NAND2_X1 U11403 ( .A1(n9125), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9018) );
  XNOR2_X1 U11404 ( .A(n9018), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9884) );
  AOI22_X1 U11405 ( .A1(n9437), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9244), .B2(
        n9884), .ZN(n9019) );
  NAND2_X1 U11406 ( .A1(n9020), .A2(n9019), .ZN(n14934) );
  NAND2_X1 U11407 ( .A1(n9005), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9029) );
  NAND2_X1 U11408 ( .A1(n9021), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9044) );
  INV_X1 U11409 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9022) );
  NAND2_X1 U11410 ( .A1(n9023), .A2(n9022), .ZN(n9024) );
  AND2_X1 U11411 ( .A1(n9044), .A2(n9024), .ZN(n10819) );
  NAND2_X1 U11412 ( .A1(n9006), .A2(n10819), .ZN(n9028) );
  NAND2_X1 U11413 ( .A1(n9251), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9027) );
  INV_X2 U11414 ( .A(n9025), .ZN(n9443) );
  NAND2_X1 U11415 ( .A1(n9443), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9026) );
  AOI22_X1 U11416 ( .A1(n14934), .A2(n9449), .B1(n6478), .B2(n13177), .ZN(
        n9036) );
  NAND2_X1 U11417 ( .A1(n14934), .A2(n9057), .ZN(n9031) );
  NAND2_X1 U11418 ( .A1(n13177), .A2(n9449), .ZN(n9030) );
  NAND2_X1 U11419 ( .A1(n9031), .A2(n9030), .ZN(n9035) );
  OAI22_X1 U11420 ( .A1(n9034), .A2(n9033), .B1(n9036), .B2(n9035), .ZN(n9038)
         );
  AOI22_X1 U11421 ( .A1(n6478), .A2(n13178), .B1(n13087), .B2(n9449), .ZN(
        n9032) );
  AOI21_X1 U11422 ( .B1(n9034), .B2(n9033), .A(n9032), .ZN(n9037) );
  NAND2_X1 U11423 ( .A1(n9723), .A2(n9436), .ZN(n9041) );
  NAND2_X1 U11424 ( .A1(n9053), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9039) );
  XNOR2_X1 U11425 ( .A(n9039), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9920) );
  AOI22_X1 U11426 ( .A1(n9437), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9244), .B2(
        n9920), .ZN(n9040) );
  NAND2_X1 U11427 ( .A1(n9041), .A2(n9040), .ZN(n14831) );
  NAND2_X1 U11428 ( .A1(n14831), .A2(n6478), .ZN(n9051) );
  NAND2_X1 U11429 ( .A1(n9005), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9049) );
  INV_X1 U11430 ( .A(n9044), .ZN(n9042) );
  NAND2_X1 U11431 ( .A1(n9042), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9059) );
  INV_X1 U11432 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9043) );
  NAND2_X1 U11433 ( .A1(n9044), .A2(n9043), .ZN(n9045) );
  AND2_X1 U11434 ( .A1(n9059), .A2(n9045), .ZN(n14827) );
  NAND2_X1 U11435 ( .A1(n9006), .A2(n14827), .ZN(n9048) );
  NAND2_X1 U11436 ( .A1(n9426), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U11437 ( .A1(n9425), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9046) );
  NAND4_X1 U11438 ( .A1(n9049), .A2(n9048), .A3(n9047), .A4(n9046), .ZN(n13176) );
  NAND2_X1 U11439 ( .A1(n13176), .A2(n9449), .ZN(n9050) );
  AOI22_X1 U11440 ( .A1(n14831), .A2(n9449), .B1(n6478), .B2(n13176), .ZN(
        n9052) );
  NAND2_X1 U11441 ( .A1(n9730), .A2(n9436), .ZN(n9056) );
  NAND2_X1 U11442 ( .A1(n9070), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9054) );
  XNOR2_X1 U11443 ( .A(n9054), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9985) );
  AOI22_X1 U11444 ( .A1(n9437), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9244), .B2(
        n9985), .ZN(n9055) );
  NAND2_X1 U11445 ( .A1(n9056), .A2(n9055), .ZN(n11060) );
  NAND2_X1 U11446 ( .A1(n11060), .A2(n9449), .ZN(n9066) );
  NAND2_X1 U11447 ( .A1(n9005), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9064) );
  NAND2_X1 U11448 ( .A1(n9059), .A2(n9058), .ZN(n9060) );
  AND2_X1 U11449 ( .A1(n9081), .A2(n9060), .ZN(n10781) );
  NAND2_X1 U11450 ( .A1(n9006), .A2(n10781), .ZN(n9063) );
  NAND2_X1 U11451 ( .A1(n9426), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9062) );
  NAND2_X1 U11452 ( .A1(n9425), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9061) );
  NAND4_X1 U11453 ( .A1(n9064), .A2(n9063), .A3(n9062), .A4(n9061), .ZN(n13175) );
  NAND2_X1 U11454 ( .A1(n9462), .A2(n13175), .ZN(n9065) );
  NAND2_X1 U11455 ( .A1(n9066), .A2(n9065), .ZN(n9069) );
  AOI22_X1 U11456 ( .A1(n11060), .A2(n9462), .B1(n9449), .B2(n13175), .ZN(
        n9068) );
  NAND2_X1 U11457 ( .A1(n9740), .A2(n9436), .ZN(n9078) );
  NAND2_X1 U11458 ( .A1(n9072), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9071) );
  MUX2_X1 U11459 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9071), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n9075) );
  INV_X1 U11460 ( .A(n9072), .ZN(n9074) );
  INV_X1 U11461 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9073) );
  NAND2_X1 U11462 ( .A1(n9074), .A2(n9073), .ZN(n9108) );
  NAND2_X1 U11463 ( .A1(n9075), .A2(n9108), .ZN(n10064) );
  INV_X1 U11464 ( .A(n9076), .ZN(n9077) );
  NAND2_X1 U11465 ( .A1(n11413), .A2(n9462), .ZN(n9088) );
  NAND2_X1 U11466 ( .A1(n9005), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n9086) );
  INV_X1 U11467 ( .A(n9081), .ZN(n9079) );
  NAND2_X1 U11468 ( .A1(n9079), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n9095) );
  INV_X1 U11469 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9080) );
  NAND2_X1 U11470 ( .A1(n9081), .A2(n9080), .ZN(n9082) );
  AND2_X1 U11471 ( .A1(n9095), .A2(n9082), .ZN(n11235) );
  NAND2_X1 U11472 ( .A1(n9006), .A2(n11235), .ZN(n9085) );
  NAND2_X1 U11473 ( .A1(n9426), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U11474 ( .A1(n9425), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9083) );
  NAND4_X1 U11475 ( .A1(n9086), .A2(n9085), .A3(n9084), .A4(n9083), .ZN(n13174) );
  NAND2_X1 U11476 ( .A1(n13174), .A2(n9449), .ZN(n9087) );
  NAND2_X1 U11477 ( .A1(n9088), .A2(n9087), .ZN(n9090) );
  AOI22_X1 U11478 ( .A1(n11413), .A2(n9449), .B1(n9462), .B2(n13174), .ZN(
        n9089) );
  NAND2_X1 U11479 ( .A1(n9749), .A2(n9436), .ZN(n9094) );
  NAND2_X1 U11480 ( .A1(n9108), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9092) );
  XNOR2_X1 U11481 ( .A(n9092), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10050) );
  AOI22_X1 U11482 ( .A1(n10050), .A2(n9244), .B1(n9437), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n9093) );
  NAND2_X1 U11483 ( .A1(n11445), .A2(n9449), .ZN(n9102) );
  NAND2_X1 U11484 ( .A1(n9005), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9100) );
  NAND2_X1 U11485 ( .A1(n9095), .A2(n11301), .ZN(n9096) );
  AND2_X1 U11486 ( .A1(n9132), .A2(n9096), .ZN(n11304) );
  NAND2_X1 U11487 ( .A1(n9006), .A2(n11304), .ZN(n9099) );
  NAND2_X1 U11488 ( .A1(n9426), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9098) );
  NAND2_X1 U11489 ( .A1(n9425), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9097) );
  NAND4_X1 U11490 ( .A1(n9100), .A2(n9099), .A3(n9098), .A4(n9097), .ZN(n13173) );
  NAND2_X1 U11491 ( .A1(n9462), .A2(n13173), .ZN(n9101) );
  NAND2_X1 U11492 ( .A1(n9102), .A2(n9101), .ZN(n9104) );
  AOI22_X1 U11493 ( .A1(n11445), .A2(n9462), .B1(n9449), .B2(n13173), .ZN(
        n9103) );
  AOI21_X1 U11494 ( .B1(n9105), .B2(n9104), .A(n9103), .ZN(n9107) );
  NOR2_X1 U11495 ( .A1(n9105), .A2(n9104), .ZN(n9106) );
  NAND2_X1 U11496 ( .A1(n9768), .A2(n9436), .ZN(n9111) );
  OAI21_X1 U11497 ( .B1(n9108), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9109) );
  XNOR2_X1 U11498 ( .A(n9109), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10083) );
  AOI21_X1 U11499 ( .B1(n10083), .B2(n9244), .A(n6492), .ZN(n9110) );
  NAND2_X1 U11500 ( .A1(n11457), .A2(n9462), .ZN(n9117) );
  XNOR2_X1 U11501 ( .A(n9132), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n11376) );
  NAND2_X1 U11502 ( .A1(n9006), .A2(n11376), .ZN(n9115) );
  NAND2_X1 U11503 ( .A1(n9005), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9114) );
  NAND2_X1 U11504 ( .A1(n9426), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n9113) );
  NAND2_X1 U11505 ( .A1(n9443), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9112) );
  NAND4_X1 U11506 ( .A1(n9115), .A2(n9114), .A3(n9113), .A4(n9112), .ZN(n13172) );
  NAND2_X1 U11507 ( .A1(n13172), .A2(n9449), .ZN(n9116) );
  NAND2_X1 U11508 ( .A1(n9117), .A2(n9116), .ZN(n9121) );
  AOI22_X1 U11509 ( .A1(n11457), .A2(n9449), .B1(n9462), .B2(n13172), .ZN(
        n9119) );
  AOI21_X1 U11510 ( .B1(n9122), .B2(n9121), .A(n9119), .ZN(n9120) );
  NAND2_X1 U11511 ( .A1(n9915), .A2(n9436), .ZN(n9128) );
  INV_X1 U11512 ( .A(n9123), .ZN(n9124) );
  NAND2_X1 U11513 ( .A1(n9142), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9126) );
  XNOR2_X1 U11514 ( .A(n9126), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U11515 ( .A1(n9437), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9244), 
        .B2(n10556), .ZN(n9127) );
  NAND2_X1 U11516 ( .A1(n14522), .A2(n9449), .ZN(n9139) );
  NAND2_X1 U11517 ( .A1(n9005), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n9137) );
  INV_X1 U11518 ( .A(n9132), .ZN(n9130) );
  AND2_X1 U11519 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n9129) );
  NAND2_X1 U11520 ( .A1(n9130), .A2(n9129), .ZN(n9147) );
  INV_X1 U11521 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n11380) );
  INV_X1 U11522 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9131) );
  OAI21_X1 U11523 ( .B1(n9132), .B2(n11380), .A(n9131), .ZN(n9133) );
  AND2_X1 U11524 ( .A1(n9147), .A2(n9133), .ZN(n14521) );
  NAND2_X1 U11525 ( .A1(n9006), .A2(n14521), .ZN(n9136) );
  NAND2_X1 U11526 ( .A1(n9426), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9135) );
  NAND2_X1 U11527 ( .A1(n9443), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n9134) );
  NAND4_X1 U11528 ( .A1(n9137), .A2(n9136), .A3(n9135), .A4(n9134), .ZN(n13171) );
  NAND2_X1 U11529 ( .A1(n9462), .A2(n13171), .ZN(n9138) );
  NAND2_X1 U11530 ( .A1(n9139), .A2(n9138), .ZN(n9141) );
  AOI22_X1 U11531 ( .A1(n14522), .A2(n9462), .B1(n9449), .B2(n13171), .ZN(
        n9140) );
  NAND2_X1 U11532 ( .A1(n10018), .A2(n9436), .ZN(n9146) );
  NAND2_X1 U11533 ( .A1(n9164), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9144) );
  INV_X1 U11534 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n9143) );
  XNOR2_X1 U11535 ( .A(n9144), .B(n9143), .ZN(n10656) );
  INV_X1 U11536 ( .A(n10656), .ZN(n10648) );
  AOI22_X1 U11537 ( .A1(n9437), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n9244), 
        .B2(n10648), .ZN(n9145) );
  NAND2_X1 U11538 ( .A1(n11696), .A2(n9462), .ZN(n9154) );
  NAND2_X1 U11539 ( .A1(n9005), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9152) );
  INV_X1 U11540 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11706) );
  NAND2_X1 U11541 ( .A1(n9147), .A2(n11706), .ZN(n9148) );
  AND2_X1 U11542 ( .A1(n9184), .A2(n9148), .ZN(n11709) );
  NAND2_X1 U11543 ( .A1(n9006), .A2(n11709), .ZN(n9151) );
  NAND2_X1 U11544 ( .A1(n9426), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n9150) );
  NAND2_X1 U11545 ( .A1(n9443), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9149) );
  NAND4_X1 U11546 ( .A1(n9152), .A2(n9151), .A3(n9150), .A4(n9149), .ZN(n13170) );
  NAND2_X1 U11547 ( .A1(n13170), .A2(n9449), .ZN(n9153) );
  NAND2_X1 U11548 ( .A1(n9154), .A2(n9153), .ZN(n9159) );
  INV_X1 U11549 ( .A(n13170), .ZN(n11536) );
  NAND2_X1 U11550 ( .A1(n11696), .A2(n9449), .ZN(n9155) );
  OAI21_X1 U11551 ( .B1(n11536), .B2(n9406), .A(n9155), .ZN(n9156) );
  NAND2_X1 U11552 ( .A1(n9157), .A2(n9156), .ZN(n9163) );
  INV_X1 U11553 ( .A(n9158), .ZN(n9161) );
  NAND2_X1 U11554 ( .A1(n9161), .A2(n9160), .ZN(n9162) );
  NAND2_X1 U11555 ( .A1(n9163), .A2(n9162), .ZN(n9176) );
  NAND2_X1 U11556 ( .A1(n10239), .A2(n9436), .ZN(n9167) );
  OR2_X1 U11557 ( .A1(n9164), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n9177) );
  NAND2_X1 U11558 ( .A1(n9177), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9165) );
  XNOR2_X1 U11559 ( .A(n9165), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11176) );
  AOI22_X1 U11560 ( .A1(n9437), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n11176), 
        .B2(n9244), .ZN(n9166) );
  NAND2_X1 U11561 ( .A1(n11727), .A2(n9449), .ZN(n9173) );
  NAND2_X1 U11562 ( .A1(n9005), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n9171) );
  XNOR2_X1 U11563 ( .A(n9184), .B(P2_REG3_REG_14__SCAN_IN), .ZN(n11733) );
  NAND2_X1 U11564 ( .A1(n9006), .A2(n11733), .ZN(n9170) );
  NAND2_X1 U11565 ( .A1(n9426), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n9169) );
  NAND2_X1 U11566 ( .A1(n9443), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n9168) );
  NAND4_X1 U11567 ( .A1(n9171), .A2(n9170), .A3(n9169), .A4(n9168), .ZN(n13169) );
  NAND2_X1 U11568 ( .A1(n9462), .A2(n13169), .ZN(n9172) );
  NAND2_X1 U11569 ( .A1(n9173), .A2(n9172), .ZN(n9175) );
  AOI22_X1 U11570 ( .A1(n11727), .A2(n9462), .B1(n9449), .B2(n13169), .ZN(
        n9174) );
  NAND2_X1 U11571 ( .A1(n10124), .A2(n9436), .ZN(n9180) );
  OAI21_X1 U11572 ( .B1(n9177), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9178) );
  XNOR2_X1 U11573 ( .A(n9178), .B(P2_IR_REG_15__SCAN_IN), .ZN(n11285) );
  AOI22_X1 U11574 ( .A1(n9244), .A2(n11285), .B1(n9437), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n9179) );
  NAND2_X1 U11575 ( .A1(n13525), .A2(n9462), .ZN(n9191) );
  INV_X1 U11576 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9182) );
  INV_X1 U11577 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9181) );
  OAI21_X1 U11578 ( .B1(n9184), .B2(n9182), .A(n9181), .ZN(n9185) );
  NAND2_X1 U11579 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .ZN(n9183) );
  AND2_X1 U11580 ( .A1(n9185), .A2(n9199), .ZN(n11743) );
  NAND2_X1 U11581 ( .A1(n9006), .A2(n11743), .ZN(n9189) );
  NAND2_X1 U11582 ( .A1(n9005), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n9188) );
  NAND2_X1 U11583 ( .A1(n9426), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n9187) );
  NAND2_X1 U11584 ( .A1(n9425), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n9186) );
  NAND4_X1 U11585 ( .A1(n9189), .A2(n9188), .A3(n9187), .A4(n9186), .ZN(n13168) );
  NAND2_X1 U11586 ( .A1(n13168), .A2(n9449), .ZN(n9190) );
  INV_X1 U11587 ( .A(n13168), .ZN(n13073) );
  NAND2_X1 U11588 ( .A1(n13525), .A2(n9449), .ZN(n9192) );
  OAI21_X1 U11589 ( .B1(n13073), .B2(n9406), .A(n9192), .ZN(n9193) );
  NAND2_X1 U11590 ( .A1(n10235), .A2(n9436), .ZN(n9197) );
  NAND2_X1 U11591 ( .A1(n9194), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9195) );
  XNOR2_X1 U11592 ( .A(n9195), .B(P2_IR_REG_16__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U11593 ( .A1(n9437), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n9244), 
        .B2(n11508), .ZN(n9196) );
  NAND2_X1 U11594 ( .A1(n13520), .A2(n9449), .ZN(n9206) );
  NAND2_X1 U11595 ( .A1(n9005), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n9204) );
  INV_X1 U11596 ( .A(n9199), .ZN(n9198) );
  NAND2_X1 U11597 ( .A1(n9198), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9221) );
  INV_X1 U11598 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n13076) );
  NAND2_X1 U11599 ( .A1(n9199), .A2(n13076), .ZN(n9200) );
  AND2_X1 U11600 ( .A1(n9221), .A2(n9200), .ZN(n13418) );
  NAND2_X1 U11601 ( .A1(n13418), .A2(n9006), .ZN(n9203) );
  NAND2_X1 U11602 ( .A1(n9426), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n9202) );
  NAND2_X1 U11603 ( .A1(n9443), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9201) );
  NAND4_X1 U11604 ( .A1(n9204), .A2(n9203), .A3(n9202), .A4(n9201), .ZN(n13167) );
  NAND2_X1 U11605 ( .A1(n9462), .A2(n13167), .ZN(n9205) );
  NAND2_X1 U11606 ( .A1(n9206), .A2(n9205), .ZN(n9208) );
  AOI22_X1 U11607 ( .A1(n13520), .A2(n9462), .B1(n9449), .B2(n13167), .ZN(
        n9207) );
  NOR2_X1 U11608 ( .A1(n9209), .A2(n9208), .ZN(n9210) );
  NAND2_X1 U11609 ( .A1(n10505), .A2(n9436), .ZN(n9216) );
  INV_X1 U11610 ( .A(n9212), .ZN(n9213) );
  NAND2_X1 U11611 ( .A1(n9213), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9214) );
  XNOR2_X1 U11612 ( .A(n9214), .B(P2_IR_REG_17__SCAN_IN), .ZN(n13188) );
  AOI22_X1 U11613 ( .A1(n9437), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n9244), 
        .B2(n13188), .ZN(n9215) );
  NAND2_X1 U11614 ( .A1(n13409), .A2(n9462), .ZN(n9226) );
  INV_X1 U11615 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13407) );
  NAND2_X1 U11616 ( .A1(n9005), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n9218) );
  NAND2_X1 U11617 ( .A1(n9426), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n9217) );
  AND2_X1 U11618 ( .A1(n9218), .A2(n9217), .ZN(n9224) );
  INV_X1 U11619 ( .A(n9221), .ZN(n9219) );
  NAND2_X1 U11620 ( .A1(n9219), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9237) );
  INV_X1 U11621 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9220) );
  NAND2_X1 U11622 ( .A1(n9221), .A2(n9220), .ZN(n9222) );
  NAND2_X1 U11623 ( .A1(n9237), .A2(n9222), .ZN(n13406) );
  OR2_X1 U11624 ( .A1(n9395), .A2(n13406), .ZN(n9223) );
  OAI211_X1 U11625 ( .C1(n9025), .C2(n13407), .A(n9224), .B(n9223), .ZN(n13166) );
  NAND2_X1 U11626 ( .A1(n13166), .A2(n9449), .ZN(n9225) );
  NAND2_X1 U11627 ( .A1(n9226), .A2(n9225), .ZN(n9229) );
  INV_X1 U11628 ( .A(n13166), .ZN(n13075) );
  NAND2_X1 U11629 ( .A1(n13409), .A2(n9449), .ZN(n9227) );
  NAND2_X1 U11630 ( .A1(n9232), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9233) );
  XNOR2_X1 U11631 ( .A(n9233), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13204) );
  AOI22_X1 U11632 ( .A1(n9437), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n9244), 
        .B2(n13204), .ZN(n9234) );
  NAND2_X2 U11633 ( .A1(n9235), .A2(n9234), .ZN(n13507) );
  NAND2_X1 U11634 ( .A1(n13507), .A2(n9449), .ZN(n9242) );
  NAND2_X1 U11635 ( .A1(n9237), .A2(n9236), .ZN(n9238) );
  NAND2_X1 U11636 ( .A1(n9249), .A2(n9238), .ZN(n13390) );
  AOI22_X1 U11637 ( .A1(n9005), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n9251), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n9240) );
  NAND2_X1 U11638 ( .A1(n9443), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9239) );
  OAI211_X1 U11639 ( .C1(n13390), .C2(n9395), .A(n9240), .B(n9239), .ZN(n13165) );
  NAND2_X1 U11640 ( .A1(n13165), .A2(n9462), .ZN(n9241) );
  AOI22_X1 U11641 ( .A1(n13507), .A2(n9462), .B1(n9449), .B2(n13165), .ZN(
        n9243) );
  NAND2_X1 U11642 ( .A1(n10787), .A2(n9436), .ZN(n9246) );
  AOI22_X1 U11643 ( .A1(n9437), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9244), 
        .B2(n8922), .ZN(n9245) );
  NAND2_X1 U11644 ( .A1(n13500), .A2(n9462), .ZN(n9256) );
  INV_X1 U11645 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9254) );
  INV_X1 U11646 ( .A(n9249), .ZN(n9247) );
  NAND2_X1 U11647 ( .A1(n9247), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9266) );
  INV_X1 U11648 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9248) );
  NAND2_X1 U11649 ( .A1(n9249), .A2(n9248), .ZN(n9250) );
  NAND2_X1 U11650 ( .A1(n9266), .A2(n9250), .ZN(n13376) );
  OR2_X1 U11651 ( .A1(n13376), .A2(n9395), .ZN(n9253) );
  AOI22_X1 U11652 ( .A1(n9005), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n9251), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n9252) );
  OAI211_X1 U11653 ( .C1(n9025), .C2(n9254), .A(n9253), .B(n9252), .ZN(n13164)
         );
  NAND2_X1 U11654 ( .A1(n13164), .A2(n9449), .ZN(n9255) );
  NAND2_X1 U11655 ( .A1(n9256), .A2(n9255), .ZN(n9259) );
  AOI22_X1 U11656 ( .A1(n13500), .A2(n9449), .B1(n9462), .B2(n13164), .ZN(
        n9257) );
  AOI21_X1 U11657 ( .B1(n9260), .B2(n9259), .A(n9257), .ZN(n9258) );
  INV_X1 U11658 ( .A(n9258), .ZN(n9263) );
  NOR2_X1 U11659 ( .A1(n9260), .A2(n9259), .ZN(n9261) );
  INV_X1 U11660 ( .A(n9261), .ZN(n9262) );
  NAND2_X1 U11661 ( .A1(n11214), .A2(n9436), .ZN(n9265) );
  NAND2_X1 U11662 ( .A1(n9437), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9264) );
  NAND2_X1 U11663 ( .A1(n13562), .A2(n9449), .ZN(n9275) );
  INV_X1 U11664 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13117) );
  NAND2_X1 U11665 ( .A1(n9266), .A2(n13117), .ZN(n9267) );
  AND2_X1 U11666 ( .A1(n9282), .A2(n9267), .ZN(n13362) );
  NAND2_X1 U11667 ( .A1(n13362), .A2(n9006), .ZN(n9273) );
  INV_X1 U11668 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9270) );
  NAND2_X1 U11669 ( .A1(n9426), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9269) );
  NAND2_X1 U11670 ( .A1(n9425), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9268) );
  OAI211_X1 U11671 ( .C1(n9270), .C2(n9446), .A(n9269), .B(n9268), .ZN(n9271)
         );
  INV_X1 U11672 ( .A(n9271), .ZN(n9272) );
  NAND2_X1 U11673 ( .A1(n9273), .A2(n9272), .ZN(n13163) );
  NAND2_X1 U11674 ( .A1(n13163), .A2(n9462), .ZN(n9274) );
  INV_X1 U11675 ( .A(n13163), .ZN(n13031) );
  NAND2_X1 U11676 ( .A1(n13562), .A2(n9462), .ZN(n9276) );
  OAI21_X1 U11677 ( .B1(n6478), .B2(n13031), .A(n9276), .ZN(n9277) );
  NAND2_X1 U11678 ( .A1(n11363), .A2(n9436), .ZN(n9279) );
  NAND2_X1 U11679 ( .A1(n9437), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n9278) );
  NAND2_X1 U11680 ( .A1(n13488), .A2(n9462), .ZN(n9291) );
  INV_X1 U11681 ( .A(n9282), .ZN(n9280) );
  NAND2_X1 U11682 ( .A1(n9280), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n9305) );
  INV_X1 U11683 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9281) );
  NAND2_X1 U11684 ( .A1(n9282), .A2(n9281), .ZN(n9283) );
  NAND2_X1 U11685 ( .A1(n9305), .A2(n9283), .ZN(n13343) );
  OR2_X1 U11686 ( .A1(n13343), .A2(n9395), .ZN(n9289) );
  INV_X1 U11687 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9286) );
  NAND2_X1 U11688 ( .A1(n9426), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9285) );
  NAND2_X1 U11689 ( .A1(n9443), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9284) );
  OAI211_X1 U11690 ( .C1(n9446), .C2(n9286), .A(n9285), .B(n9284), .ZN(n9287)
         );
  INV_X1 U11691 ( .A(n9287), .ZN(n9288) );
  NAND2_X1 U11692 ( .A1(n9289), .A2(n9288), .ZN(n13162) );
  NAND2_X1 U11693 ( .A1(n13162), .A2(n9449), .ZN(n9290) );
  NAND2_X1 U11694 ( .A1(n9291), .A2(n9290), .ZN(n9294) );
  AOI22_X1 U11695 ( .A1(n13488), .A2(n9449), .B1(n9462), .B2(n13162), .ZN(
        n9292) );
  AOI21_X1 U11696 ( .B1(n9295), .B2(n9294), .A(n9292), .ZN(n9293) );
  INV_X1 U11697 ( .A(n9293), .ZN(n9296) );
  INV_X1 U11698 ( .A(n9297), .ZN(n9300) );
  INV_X1 U11699 ( .A(n9298), .ZN(n9299) );
  NAND2_X1 U11700 ( .A1(n9300), .A2(n9299), .ZN(n9301) );
  AND2_X1 U11701 ( .A1(n9302), .A2(n9301), .ZN(n11675) );
  NAND2_X1 U11702 ( .A1(n11675), .A2(n9436), .ZN(n9304) );
  NAND2_X1 U11703 ( .A1(n9437), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9303) );
  NAND2_X1 U11704 ( .A1(n13331), .A2(n9449), .ZN(n9313) );
  INV_X1 U11705 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13124) );
  NAND2_X1 U11706 ( .A1(n9305), .A2(n13124), .ZN(n9306) );
  AND2_X1 U11707 ( .A1(n9322), .A2(n9306), .ZN(n13332) );
  NAND2_X1 U11708 ( .A1(n13332), .A2(n9006), .ZN(n9311) );
  INV_X1 U11709 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n13484) );
  NAND2_X1 U11710 ( .A1(n9425), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9308) );
  NAND2_X1 U11711 ( .A1(n9426), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9307) );
  OAI211_X1 U11712 ( .C1(n9446), .C2(n13484), .A(n9308), .B(n9307), .ZN(n9309)
         );
  INV_X1 U11713 ( .A(n9309), .ZN(n9310) );
  NAND2_X1 U11714 ( .A1(n9311), .A2(n9310), .ZN(n13161) );
  NAND2_X1 U11715 ( .A1(n13161), .A2(n9462), .ZN(n9312) );
  NAND2_X1 U11716 ( .A1(n9313), .A2(n9312), .ZN(n9316) );
  INV_X1 U11717 ( .A(n13161), .ZN(n12158) );
  NAND2_X1 U11718 ( .A1(n13331), .A2(n9462), .ZN(n9314) );
  OAI21_X1 U11719 ( .B1(n6478), .B2(n12158), .A(n9314), .ZN(n9315) );
  NAND2_X1 U11720 ( .A1(n11692), .A2(n9436), .ZN(n9319) );
  NAND2_X1 U11721 ( .A1(n9437), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9318) );
  NAND2_X1 U11722 ( .A1(n13476), .A2(n9462), .ZN(n9331) );
  INV_X1 U11723 ( .A(n9322), .ZN(n9320) );
  NAND2_X1 U11724 ( .A1(n9320), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n9335) );
  INV_X1 U11725 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9321) );
  NAND2_X1 U11726 ( .A1(n9322), .A2(n9321), .ZN(n9323) );
  NAND2_X1 U11727 ( .A1(n9335), .A2(n9323), .ZN(n13313) );
  OR2_X1 U11728 ( .A1(n13313), .A2(n9395), .ZN(n9329) );
  INV_X1 U11729 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9326) );
  NAND2_X1 U11730 ( .A1(n9443), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9325) );
  NAND2_X1 U11731 ( .A1(n9426), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9324) );
  OAI211_X1 U11732 ( .C1(n9446), .C2(n9326), .A(n9325), .B(n9324), .ZN(n9327)
         );
  INV_X1 U11733 ( .A(n9327), .ZN(n9328) );
  NAND2_X1 U11734 ( .A1(n9329), .A2(n9328), .ZN(n13160) );
  NAND2_X1 U11735 ( .A1(n13160), .A2(n9449), .ZN(n9330) );
  AOI22_X1 U11736 ( .A1(n13476), .A2(n9449), .B1(n9462), .B2(n13160), .ZN(
        n9332) );
  NAND2_X1 U11737 ( .A1(n9437), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9333) );
  NAND2_X1 U11738 ( .A1(n13470), .A2(n9449), .ZN(n9344) );
  INV_X1 U11739 ( .A(n9335), .ZN(n9334) );
  NAND2_X1 U11740 ( .A1(n9334), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n9353) );
  INV_X1 U11741 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13106) );
  NAND2_X1 U11742 ( .A1(n9335), .A2(n13106), .ZN(n9336) );
  NAND2_X1 U11743 ( .A1(n9353), .A2(n9336), .ZN(n13304) );
  OR2_X1 U11744 ( .A1(n13304), .A2(n9395), .ZN(n9342) );
  INV_X1 U11745 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9339) );
  NAND2_X1 U11746 ( .A1(n9425), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9338) );
  NAND2_X1 U11747 ( .A1(n9426), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9337) );
  OAI211_X1 U11748 ( .C1(n9446), .C2(n9339), .A(n9338), .B(n9337), .ZN(n9340)
         );
  INV_X1 U11749 ( .A(n9340), .ZN(n9341) );
  NAND2_X1 U11750 ( .A1(n9342), .A2(n9341), .ZN(n13159) );
  NAND2_X1 U11751 ( .A1(n13159), .A2(n6478), .ZN(n9343) );
  NAND2_X1 U11752 ( .A1(n9344), .A2(n9343), .ZN(n9346) );
  AOI22_X1 U11753 ( .A1(n13470), .A2(n6478), .B1(n9449), .B2(n13159), .ZN(
        n9345) );
  AOI21_X1 U11754 ( .B1(n9347), .B2(n9346), .A(n9345), .ZN(n9349) );
  NOR2_X1 U11755 ( .A1(n9347), .A2(n9346), .ZN(n9348) );
  NAND2_X1 U11756 ( .A1(n13594), .A2(n9436), .ZN(n9351) );
  NAND2_X1 U11757 ( .A1(n9437), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9350) );
  INV_X1 U11758 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9352) );
  NAND2_X1 U11759 ( .A1(n9353), .A2(n9352), .ZN(n9354) );
  NAND2_X1 U11760 ( .A1(n9369), .A2(n9354), .ZN(n13289) );
  OR2_X1 U11761 ( .A1(n13289), .A2(n9395), .ZN(n9359) );
  INV_X1 U11762 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13465) );
  NAND2_X1 U11763 ( .A1(n9443), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9356) );
  NAND2_X1 U11764 ( .A1(n9426), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9355) );
  OAI211_X1 U11765 ( .C1(n9446), .C2(n13465), .A(n9356), .B(n9355), .ZN(n9357)
         );
  INV_X1 U11766 ( .A(n9357), .ZN(n9358) );
  NAND2_X1 U11767 ( .A1(n9359), .A2(n9358), .ZN(n13158) );
  AND2_X1 U11768 ( .A1(n13158), .A2(n9449), .ZN(n9361) );
  AOI21_X1 U11769 ( .B1(n13288), .B2(n6478), .A(n9361), .ZN(n9365) );
  INV_X1 U11770 ( .A(n13158), .ZN(n12166) );
  NAND2_X1 U11771 ( .A1(n13288), .A2(n9449), .ZN(n9362) );
  NAND2_X1 U11772 ( .A1(n13591), .A2(n9436), .ZN(n9367) );
  NAND2_X1 U11773 ( .A1(n9437), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9366) );
  NAND2_X2 U11774 ( .A1(n9367), .A2(n9366), .ZN(n13543) );
  NAND2_X1 U11775 ( .A1(n13543), .A2(n9449), .ZN(n9377) );
  INV_X1 U11776 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9368) );
  NAND2_X1 U11777 ( .A1(n9369), .A2(n9368), .ZN(n9370) );
  NAND2_X1 U11778 ( .A1(n13272), .A2(n9006), .ZN(n9375) );
  INV_X1 U11779 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n10260) );
  NAND2_X1 U11780 ( .A1(n9425), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9372) );
  NAND2_X1 U11781 ( .A1(n9426), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9371) );
  OAI211_X1 U11782 ( .C1(n9446), .C2(n10260), .A(n9372), .B(n9371), .ZN(n9373)
         );
  INV_X1 U11783 ( .A(n9373), .ZN(n9374) );
  NAND2_X1 U11784 ( .A1(n9375), .A2(n9374), .ZN(n13157) );
  NAND2_X1 U11785 ( .A1(n13157), .A2(n9462), .ZN(n9376) );
  AOI22_X1 U11786 ( .A1(n13543), .A2(n9462), .B1(n9449), .B2(n13157), .ZN(
        n9378) );
  NAND2_X1 U11787 ( .A1(n13588), .A2(n9436), .ZN(n9380) );
  NAND2_X1 U11788 ( .A1(n9437), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9379) );
  NAND2_X2 U11789 ( .A1(n9380), .A2(n9379), .ZN(n13448) );
  NAND2_X1 U11790 ( .A1(n13448), .A2(n9462), .ZN(n9387) );
  XNOR2_X1 U11791 ( .A(n9392), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n13256) );
  NAND2_X1 U11792 ( .A1(n13256), .A2(n9006), .ZN(n9385) );
  INV_X1 U11793 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n13454) );
  NAND2_X1 U11794 ( .A1(n9426), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9382) );
  NAND2_X1 U11795 ( .A1(n9443), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9381) );
  OAI211_X1 U11796 ( .C1(n9446), .C2(n13454), .A(n9382), .B(n9381), .ZN(n9383)
         );
  INV_X1 U11797 ( .A(n9383), .ZN(n9384) );
  NAND2_X1 U11798 ( .A1(n9385), .A2(n9384), .ZN(n13156) );
  NAND2_X1 U11799 ( .A1(n13156), .A2(n9449), .ZN(n9386) );
  NAND2_X1 U11800 ( .A1(n9387), .A2(n9386), .ZN(n9408) );
  NAND2_X1 U11801 ( .A1(n9409), .A2(n9408), .ZN(n9411) );
  INV_X1 U11802 ( .A(n13448), .ZN(n13010) );
  INV_X1 U11803 ( .A(n13156), .ZN(n12170) );
  OAI22_X1 U11804 ( .A1(n13010), .A2(n6478), .B1(n12170), .B2(n9406), .ZN(
        n9410) );
  NAND2_X1 U11805 ( .A1(n13583), .A2(n9436), .ZN(n9389) );
  NAND2_X1 U11806 ( .A1(n9437), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9388) );
  NAND2_X1 U11807 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n9390) );
  NOR2_X1 U11808 ( .A1(n9392), .A2(n9390), .ZN(n12180) );
  INV_X1 U11809 ( .A(n12180), .ZN(n9394) );
  INV_X1 U11810 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9391) );
  INV_X1 U11811 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n13047) );
  OAI21_X1 U11812 ( .B1(n9392), .B2(n9391), .A(n13047), .ZN(n9393) );
  NAND2_X1 U11813 ( .A1(n9394), .A2(n9393), .ZN(n13239) );
  INV_X1 U11814 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9398) );
  NAND2_X1 U11815 ( .A1(n9425), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9397) );
  NAND2_X1 U11816 ( .A1(n9426), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9396) );
  OAI211_X1 U11817 ( .C1(n9446), .C2(n9398), .A(n9397), .B(n9396), .ZN(n9399)
         );
  INV_X1 U11818 ( .A(n9399), .ZN(n9400) );
  AOI22_X1 U11819 ( .A1(n12172), .A2(n6478), .B1(n9449), .B2(n13155), .ZN(
        n9413) );
  OAI22_X1 U11820 ( .A1(n13540), .A2(n6478), .B1(n13011), .B2(n9406), .ZN(
        n9412) );
  INV_X1 U11821 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9404) );
  NAND2_X1 U11822 ( .A1(n9443), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9403) );
  NAND2_X1 U11823 ( .A1(n9426), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9402) );
  OAI211_X1 U11824 ( .C1(n9446), .C2(n9404), .A(n9403), .B(n9402), .ZN(n9405)
         );
  AOI21_X1 U11825 ( .B1(n12180), .B2(n9006), .A(n9405), .ZN(n13044) );
  INV_X1 U11826 ( .A(n13044), .ZN(n13154) );
  AOI22_X1 U11827 ( .A1(n13438), .A2(n9449), .B1(n6478), .B2(n13154), .ZN(
        n9451) );
  OAI22_X1 U11828 ( .A1(n12182), .A2(n9449), .B1(n6478), .B2(n13044), .ZN(
        n9450) );
  NOR2_X1 U11829 ( .A1(n9451), .A2(n9450), .ZN(n9414) );
  AOI21_X1 U11830 ( .B1(n9413), .B2(n9412), .A(n9414), .ZN(n9407) );
  NOR3_X1 U11831 ( .A1(n9414), .A2(n9413), .A3(n9412), .ZN(n9429) );
  INV_X1 U11832 ( .A(SI_29_), .ZN(n12959) );
  MUX2_X1 U11833 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9685), .Z(n9418) );
  XNOR2_X1 U11834 ( .A(n9418), .B(SI_30_), .ZN(n9433) );
  NAND2_X1 U11835 ( .A1(n9418), .A2(SI_30_), .ZN(n9419) );
  MUX2_X1 U11836 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9685), .Z(n9420) );
  XNOR2_X1 U11837 ( .A(n9420), .B(SI_31_), .ZN(n9421) );
  NAND2_X1 U11838 ( .A1(n14236), .A2(n9436), .ZN(n9424) );
  NAND2_X1 U11839 ( .A1(n9437), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9423) );
  INV_X1 U11840 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13431) );
  NAND2_X1 U11841 ( .A1(n9425), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9428) );
  NAND2_X1 U11842 ( .A1(n9426), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9427) );
  OAI211_X1 U11843 ( .C1(n9446), .C2(n13431), .A(n9428), .B(n9427), .ZN(n13220) );
  XNOR2_X1 U11844 ( .A(n9430), .B(n13220), .ZN(n9487) );
  INV_X1 U11845 ( .A(n13220), .ZN(n9440) );
  AOI21_X1 U11846 ( .B1(n6478), .B2(n13220), .A(n9432), .ZN(n9453) );
  INV_X1 U11847 ( .A(n9433), .ZN(n9434) );
  NAND2_X1 U11848 ( .A1(n11998), .A2(n9436), .ZN(n9439) );
  NAND2_X1 U11849 ( .A1(n9437), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9438) );
  NOR2_X1 U11850 ( .A1(n9440), .A2(n6478), .ZN(n9461) );
  NAND2_X1 U11851 ( .A1(n8923), .A2(n13213), .ZN(n10210) );
  OAI211_X1 U11852 ( .C1(n9441), .C2(n10695), .A(n9442), .B(n10210), .ZN(n9447) );
  INV_X1 U11853 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13435) );
  NAND2_X1 U11854 ( .A1(n9443), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9445) );
  NAND2_X1 U11855 ( .A1(n9426), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9444) );
  OAI211_X1 U11856 ( .C1(n9446), .C2(n13435), .A(n9445), .B(n9444), .ZN(n13153) );
  OAI21_X1 U11857 ( .B1(n9461), .B2(n9447), .A(n13153), .ZN(n9448) );
  OAI21_X1 U11858 ( .B1(n13536), .B2(n9449), .A(n9448), .ZN(n9456) );
  INV_X1 U11859 ( .A(n13536), .ZN(n9484) );
  AOI22_X1 U11860 ( .A1(n9484), .A2(n9449), .B1(n9462), .B2(n13153), .ZN(n9455) );
  AOI22_X1 U11861 ( .A1(n9456), .A2(n9455), .B1(n9451), .B2(n9450), .ZN(n9452)
         );
  OR2_X1 U11862 ( .A1(n9453), .A2(n9452), .ZN(n9454) );
  INV_X1 U11863 ( .A(n9455), .ZN(n9458) );
  INV_X1 U11864 ( .A(n9456), .ZN(n9457) );
  INV_X1 U11865 ( .A(n9459), .ZN(n9460) );
  AOI211_X1 U11866 ( .C1(n9462), .C2(n9430), .A(n9461), .B(n9460), .ZN(n9463)
         );
  OR2_X1 U11867 ( .A1(n9466), .A2(n9465), .ZN(n9467) );
  AND2_X1 U11868 ( .A1(n9833), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11672) );
  INV_X1 U11869 ( .A(n9468), .ZN(n14864) );
  NAND2_X1 U11870 ( .A1(n10695), .A2(n8922), .ZN(n9469) );
  OAI22_X1 U11871 ( .A1(n9441), .A2(n14864), .B1(n6618), .B2(n9469), .ZN(n9470) );
  NAND3_X1 U11872 ( .A1(n9491), .A2(n11672), .A3(n9470), .ZN(n9506) );
  NAND2_X1 U11873 ( .A1(n12172), .A2(n13155), .ZN(n12207) );
  OR2_X1 U11874 ( .A1(n12172), .A2(n13155), .ZN(n9471) );
  XNOR2_X1 U11875 ( .A(n13448), .B(n12170), .ZN(n13260) );
  XNOR2_X1 U11876 ( .A(n13543), .B(n13157), .ZN(n13266) );
  OR2_X1 U11877 ( .A1(n13476), .A2(n13160), .ZN(n12201) );
  NAND2_X1 U11878 ( .A1(n13476), .A2(n13160), .ZN(n12199) );
  XNOR2_X1 U11879 ( .A(n13562), .B(n13031), .ZN(n13357) );
  NOR2_X1 U11880 ( .A1(n13488), .A2(n13162), .ZN(n12196) );
  AND2_X1 U11881 ( .A1(n13488), .A2(n13162), .ZN(n12195) );
  NOR2_X1 U11882 ( .A1(n12196), .A2(n12195), .ZN(n13347) );
  XNOR2_X1 U11883 ( .A(n13500), .B(n13164), .ZN(n13379) );
  OR2_X1 U11884 ( .A1(n13409), .A2(n13166), .ZN(n12188) );
  NAND2_X1 U11885 ( .A1(n13409), .A2(n13166), .ZN(n12187) );
  AND2_X1 U11886 ( .A1(n12188), .A2(n12187), .ZN(n13402) );
  XNOR2_X1 U11887 ( .A(n13525), .B(n13073), .ZN(n12183) );
  XNOR2_X1 U11888 ( .A(n11727), .B(n13169), .ZN(n11543) );
  INV_X1 U11889 ( .A(n13172), .ZN(n11448) );
  XNOR2_X1 U11890 ( .A(n11457), .B(n11448), .ZN(n11455) );
  INV_X1 U11891 ( .A(n13173), .ZN(n11241) );
  XNOR2_X1 U11892 ( .A(n11445), .B(n11241), .ZN(n11250) );
  INV_X1 U11893 ( .A(n13174), .ZN(n11019) );
  XNOR2_X1 U11894 ( .A(n11413), .B(n11019), .ZN(n11027) );
  INV_X1 U11895 ( .A(n13175), .ZN(n10965) );
  XNOR2_X1 U11896 ( .A(n11060), .B(n10965), .ZN(n10718) );
  XNOR2_X1 U11897 ( .A(n14831), .B(n13176), .ZN(n10694) );
  NAND2_X1 U11898 ( .A1(n9472), .A2(n8919), .ZN(n12002) );
  NAND2_X1 U11899 ( .A1(n9473), .A2(n12002), .ZN(n14887) );
  XNOR2_X2 U11900 ( .A(n13182), .B(n10677), .ZN(n10874) );
  XNOR2_X1 U11901 ( .A(n13181), .B(n10900), .ZN(n10681) );
  NAND4_X1 U11902 ( .A1(n14887), .A2(n10695), .A3(n10874), .A4(n10681), .ZN(
        n9474) );
  XNOR2_X1 U11903 ( .A(n13179), .B(n14917), .ZN(n14847) );
  NOR3_X1 U11904 ( .A1(n9474), .A2(n14847), .A3(n10685), .ZN(n9475) );
  XNOR2_X1 U11905 ( .A(n14934), .B(n13177), .ZN(n10813) );
  XNOR2_X1 U11906 ( .A(n13087), .B(n13178), .ZN(n10802) );
  NAND4_X1 U11907 ( .A1(n10694), .A2(n9475), .A3(n10813), .A4(n10802), .ZN(
        n9476) );
  OR4_X1 U11908 ( .A1(n11250), .A2(n11027), .A3(n10718), .A4(n9476), .ZN(n9477) );
  NOR2_X1 U11909 ( .A1(n11455), .A2(n9477), .ZN(n9478) );
  XNOR2_X1 U11910 ( .A(n11696), .B(n13170), .ZN(n11534) );
  XNOR2_X1 U11911 ( .A(n14522), .B(n13171), .ZN(n14523) );
  NAND4_X1 U11912 ( .A1(n11543), .A2(n9478), .A3(n11534), .A4(n14523), .ZN(
        n9479) );
  NOR3_X1 U11913 ( .A1(n13402), .A2(n12183), .A3(n9479), .ZN(n9480) );
  XNOR2_X1 U11914 ( .A(n13507), .B(n13165), .ZN(n12189) );
  XNOR2_X1 U11915 ( .A(n13520), .B(n13167), .ZN(n13422) );
  NAND4_X1 U11916 ( .A1(n13379), .A2(n9480), .A3(n12189), .A4(n13422), .ZN(
        n9481) );
  NOR4_X1 U11917 ( .A1(n13309), .A2(n13357), .A3(n13347), .A4(n9481), .ZN(
        n9482) );
  XNOR2_X1 U11918 ( .A(n13331), .B(n13161), .ZN(n13326) );
  NAND4_X1 U11919 ( .A1(n13266), .A2(n9482), .A3(n13301), .A4(n13326), .ZN(
        n9483) );
  NOR4_X1 U11920 ( .A1(n13232), .A2(n13260), .A3(n13283), .A4(n9483), .ZN(
        n9486) );
  XNOR2_X1 U11921 ( .A(n9484), .B(n13153), .ZN(n9485) );
  NAND4_X1 U11922 ( .A1(n9487), .A2(n9486), .A3(n9485), .A4(n12208), .ZN(n9488) );
  XOR2_X1 U11923 ( .A(n9488), .B(n8922), .Z(n9489) );
  INV_X1 U11924 ( .A(n11672), .ZN(n9501) );
  NOR3_X1 U11925 ( .A1(n9489), .A2(n9442), .A3(n9501), .ZN(n9490) );
  OAI21_X1 U11926 ( .B1(n9232), .B2(n9494), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9495) );
  MUX2_X1 U11927 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9495), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9496) );
  NAND2_X1 U11928 ( .A1(n6592), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9497) );
  MUX2_X1 U11929 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9497), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n9498) );
  AOI21_X1 U11930 ( .B1(n13597), .B2(n9507), .A(n9833), .ZN(n10211) );
  INV_X1 U11931 ( .A(n13589), .ZN(n9838) );
  INV_X1 U11932 ( .A(n10210), .ZN(n10214) );
  INV_X1 U11933 ( .A(n10217), .ZN(n9499) );
  NAND4_X1 U11934 ( .A1(n14886), .A2(n9838), .A3(n10214), .A4(n13142), .ZN(
        n9500) );
  OAI211_X1 U11935 ( .C1(n8921), .C2(n9501), .A(n9500), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9504) );
  AOI21_X1 U11936 ( .B1(n6618), .B2(n10695), .A(n8922), .ZN(n9503) );
  INV_X4 U11937 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U11938 ( .A(n9507), .ZN(n9508) );
  NOR2_X1 U11939 ( .A1(n9833), .A2(n9508), .ZN(n9509) );
  NAND2_X1 U11940 ( .A1(n13597), .A2(n9509), .ZN(n9836) );
  XNOR2_X1 U11941 ( .A(n11264), .B(P3_B_REG_SCAN_IN), .ZN(n9510) );
  NAND2_X1 U11942 ( .A1(n9510), .A2(n11368), .ZN(n9511) );
  INV_X1 U11943 ( .A(n9512), .ZN(n11499) );
  NAND2_X1 U11944 ( .A1(n11499), .A2(n11264), .ZN(n9513) );
  NAND2_X1 U11945 ( .A1(n12948), .A2(n6507), .ZN(n9517) );
  NAND2_X1 U11946 ( .A1(n10614), .A2(n12550), .ZN(n9515) );
  NAND2_X1 U11947 ( .A1(n9515), .A2(n10563), .ZN(n9516) );
  NAND3_X1 U11948 ( .A1(n12463), .A2(n12296), .A3(n10945), .ZN(n9521) );
  NAND2_X1 U11949 ( .A1(n10737), .A2(n10870), .ZN(n10927) );
  NAND2_X1 U11950 ( .A1(n10927), .A2(n12296), .ZN(n9522) );
  NAND2_X1 U11951 ( .A1(n9523), .A2(n9522), .ZN(n9524) );
  XNOR2_X1 U11952 ( .A(n11040), .B(n12296), .ZN(n9526) );
  NAND2_X1 U11953 ( .A1(n9526), .A2(n11041), .ZN(n9527) );
  NAND2_X1 U11954 ( .A1(n9528), .A2(n9527), .ZN(n10953) );
  XNOR2_X1 U11955 ( .A(n9531), .B(n15186), .ZN(n10952) );
  INV_X1 U11956 ( .A(n9531), .ZN(n9532) );
  NAND2_X1 U11957 ( .A1(n9532), .A2(n12461), .ZN(n9533) );
  XNOR2_X1 U11958 ( .A(n9534), .B(n12296), .ZN(n9535) );
  XNOR2_X1 U11959 ( .A(n9535), .B(n12460), .ZN(n11217) );
  NAND2_X1 U11960 ( .A1(n9535), .A2(n15164), .ZN(n9536) );
  XNOR2_X1 U11961 ( .A(n15171), .B(n12296), .ZN(n9537) );
  XNOR2_X1 U11962 ( .A(n9537), .B(n12212), .ZN(n11307) );
  INV_X1 U11963 ( .A(n9537), .ZN(n9538) );
  NAND2_X1 U11964 ( .A1(n9538), .A2(n12212), .ZN(n9539) );
  NAND2_X1 U11965 ( .A1(n9540), .A2(n9539), .ZN(n12418) );
  XNOR2_X1 U11966 ( .A(n15149), .B(n12328), .ZN(n9541) );
  XNOR2_X1 U11967 ( .A(n9541), .B(n15163), .ZN(n12419) );
  INV_X1 U11968 ( .A(n9541), .ZN(n9542) );
  NAND2_X1 U11969 ( .A1(n12458), .A2(n9542), .ZN(n9543) );
  XNOR2_X1 U11970 ( .A(n15125), .B(n12296), .ZN(n11501) );
  NAND2_X1 U11971 ( .A1(n7045), .A2(n15143), .ZN(n9544) );
  XNOR2_X1 U11972 ( .A(n12225), .B(n12328), .ZN(n9545) );
  XNOR2_X1 U11973 ( .A(n9545), .B(n12457), .ZN(n11562) );
  INV_X1 U11974 ( .A(n9545), .ZN(n9546) );
  NAND2_X1 U11975 ( .A1(n9546), .A2(n12457), .ZN(n9547) );
  XNOR2_X1 U11976 ( .A(n15241), .B(n12328), .ZN(n9548) );
  XNOR2_X1 U11977 ( .A(n9548), .B(n15112), .ZN(n12375) );
  XNOR2_X1 U11978 ( .A(n14964), .B(n12296), .ZN(n9550) );
  XNOR2_X1 U11979 ( .A(n9550), .B(n14495), .ZN(n14961) );
  NAND2_X1 U11980 ( .A1(n9548), .A2(n15112), .ZN(n14957) );
  AND2_X1 U11981 ( .A1(n14961), .A2(n14957), .ZN(n9549) );
  NAND2_X1 U11982 ( .A1(n9550), .A2(n12456), .ZN(n9551) );
  XNOR2_X1 U11983 ( .A(n14497), .B(n12296), .ZN(n9553) );
  INV_X1 U11984 ( .A(n9552), .ZN(n9555) );
  INV_X1 U11985 ( .A(n9553), .ZN(n9554) );
  NAND2_X1 U11986 ( .A1(n9555), .A2(n9554), .ZN(n9597) );
  NAND2_X1 U11987 ( .A1(n9596), .A2(n9597), .ZN(n9556) );
  XNOR2_X1 U11988 ( .A(n9556), .B(n12797), .ZN(n9575) );
  OR2_X1 U11989 ( .A1(n9766), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9558) );
  NAND2_X1 U11990 ( .A1(n11499), .A2(n11368), .ZN(n9557) );
  AND2_X1 U11991 ( .A1(n9558), .A2(n9557), .ZN(n12946) );
  INV_X1 U11992 ( .A(n12946), .ZN(n10861) );
  AND2_X1 U11993 ( .A1(n10862), .A2(n10861), .ZN(n10630) );
  NOR2_X1 U11994 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n9562) );
  NOR4_X1 U11995 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9561) );
  NOR4_X1 U11996 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n9560) );
  NOR4_X1 U11997 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9559) );
  NAND4_X1 U11998 ( .A1(n9562), .A2(n9561), .A3(n9560), .A4(n9559), .ZN(n9568)
         );
  NOR4_X1 U11999 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9566) );
  NOR4_X1 U12000 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n9565) );
  NOR4_X1 U12001 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9564) );
  NOR4_X1 U12002 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9563) );
  NAND4_X1 U12003 ( .A1(n9566), .A2(n9565), .A3(n9564), .A4(n9563), .ZN(n9567)
         );
  NOR2_X1 U12004 ( .A1(n9568), .A2(n9567), .ZN(n9569) );
  AND2_X1 U12005 ( .A1(n10730), .A2(n12550), .ZN(n10928) );
  NAND2_X1 U12006 ( .A1(n10928), .A2(n6507), .ZN(n10605) );
  NAND2_X1 U12007 ( .A1(n10614), .A2(n10563), .ZN(n9570) );
  XNOR2_X1 U12008 ( .A(n10730), .B(n9570), .ZN(n9572) );
  NAND2_X1 U12009 ( .A1(n10614), .A2(n12523), .ZN(n9571) );
  AND2_X1 U12010 ( .A1(n9572), .A2(n9571), .ZN(n10610) );
  INV_X1 U12011 ( .A(n10610), .ZN(n10939) );
  NAND3_X1 U12012 ( .A1(n10608), .A2(n10939), .A3(n15219), .ZN(n9573) );
  OAI21_X1 U12013 ( .B1(n10611), .B2(n10605), .A(n9573), .ZN(n9574) );
  NOR2_X1 U12014 ( .A1(n9575), .A2(n12433), .ZN(n9595) );
  INV_X1 U12015 ( .A(n10608), .ZN(n9576) );
  NAND2_X1 U12016 ( .A1(n9576), .A2(n10946), .ZN(n9578) );
  AND2_X1 U12017 ( .A1(n10866), .A2(n15242), .ZN(n9577) );
  AND2_X1 U12018 ( .A1(n14965), .A2(n12229), .ZN(n9594) );
  INV_X1 U12019 ( .A(n10937), .ZN(n10635) );
  NAND2_X1 U12020 ( .A1(n9650), .A2(n10635), .ZN(n10631) );
  AND3_X1 U12021 ( .A1(n10631), .A2(n9607), .A3(n9649), .ZN(n9581) );
  INV_X1 U12022 ( .A(n10605), .ZN(n9579) );
  NAND2_X1 U12023 ( .A1(n10611), .A2(n9579), .ZN(n9580) );
  OAI211_X1 U12024 ( .C1(n10608), .C2(n10610), .A(n9581), .B(n9580), .ZN(n9582) );
  NAND2_X1 U12025 ( .A1(n9582), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9585) );
  NAND2_X1 U12026 ( .A1(n9650), .A2(n10937), .ZN(n10606) );
  INV_X1 U12027 ( .A(n10606), .ZN(n9583) );
  NAND3_X1 U12028 ( .A1(n10611), .A2(n10866), .A3(n9583), .ZN(n9584) );
  INV_X1 U12029 ( .A(n14498), .ZN(n9586) );
  NOR2_X1 U12030 ( .A1(n14971), .A2(n9586), .ZN(n9593) );
  NAND2_X1 U12031 ( .A1(n9657), .A2(n6722), .ZN(n9587) );
  NAND2_X1 U12032 ( .A1(n10866), .A2(n10937), .ZN(n9588) );
  NOR2_X1 U12033 ( .A1(n15185), .A2(n14968), .ZN(n12422) );
  INV_X1 U12034 ( .A(n12422), .ZN(n12440) );
  INV_X1 U12035 ( .A(n12414), .ZN(n12437) );
  NAND2_X1 U12036 ( .A1(n12456), .A2(n12437), .ZN(n9591) );
  INV_X1 U12037 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n9589) );
  NOR2_X1 U12038 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9589), .ZN(n11207) );
  INV_X1 U12039 ( .A(n11207), .ZN(n9590) );
  OAI211_X1 U12040 ( .C1(n12440), .C2(n14496), .A(n9591), .B(n9590), .ZN(n9592) );
  NAND2_X1 U12041 ( .A1(n9596), .A2(n14956), .ZN(n9598) );
  NAND2_X1 U12042 ( .A1(n9598), .A2(n9597), .ZN(n12267) );
  XNOR2_X1 U12043 ( .A(n12232), .B(n12328), .ZN(n12268) );
  XNOR2_X1 U12044 ( .A(n12455), .B(n12268), .ZN(n9599) );
  XNOR2_X1 U12045 ( .A(n12267), .B(n9599), .ZN(n9600) );
  NOR2_X1 U12046 ( .A1(n9600), .A2(n12433), .ZN(n9606) );
  AND2_X1 U12047 ( .A1(n14965), .A2(n12232), .ZN(n9605) );
  INV_X1 U12048 ( .A(n9601), .ZN(n12800) );
  NOR2_X1 U12049 ( .A1(n14971), .A2(n12800), .ZN(n9604) );
  NAND2_X1 U12050 ( .A1(n14956), .A2(n12437), .ZN(n9602) );
  INV_X1 U12051 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n10360) );
  OR2_X1 U12052 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10360), .ZN(n11427) );
  OAI211_X1 U12053 ( .C1(n12440), .C2(n12798), .A(n9602), .B(n11427), .ZN(
        n9603) );
  INV_X1 U12054 ( .A(n9607), .ZN(n9608) );
  AOI22_X1 U12055 ( .A1(n12125), .A2(n13770), .B1(n12118), .B2(n10532), .ZN(
        n9609) );
  XNOR2_X1 U12056 ( .A(n9609), .B(n12132), .ZN(n10758) );
  INV_X2 U12057 ( .A(n11396), .ZN(n12125) );
  AOI22_X1 U12058 ( .A1(n12068), .A2(n13770), .B1(n12125), .B2(n10532), .ZN(
        n10759) );
  XNOR2_X1 U12059 ( .A(n10758), .B(n10759), .ZN(n9629) );
  NAND2_X1 U12060 ( .A1(n11344), .A2(n10135), .ZN(n9611) );
  OR2_X1 U12061 ( .A1(n9634), .A2(n9760), .ZN(n9610) );
  OAI211_X1 U12062 ( .C1(n12131), .C2(n10130), .A(n9611), .B(n9610), .ZN(
        n10075) );
  INV_X1 U12063 ( .A(n9634), .ZN(n9612) );
  AOI222_X1 U12064 ( .A1(n10135), .A2(n12068), .B1(n7679), .B2(n11344), .C1(
        P1_IR_REG_0__SCAN_IN), .C2(n9612), .ZN(n10076) );
  NAND2_X1 U12065 ( .A1(n10076), .A2(n10075), .ZN(n10074) );
  AOI22_X1 U12066 ( .A1(n12118), .A2(n11778), .B1(n11344), .B2(n13772), .ZN(
        n9613) );
  INV_X1 U12067 ( .A(n13772), .ZN(n9614) );
  XNOR2_X1 U12068 ( .A(n9616), .B(n9617), .ZN(n10034) );
  NOR2_X1 U12069 ( .A1(n9618), .A2(n9617), .ZN(n9619) );
  AOI21_X1 U12070 ( .B1(n10033), .B2(n10034), .A(n9619), .ZN(n10099) );
  INV_X1 U12071 ( .A(n13771), .ZN(n10136) );
  AOI22_X1 U12072 ( .A1(n11344), .A2(n13771), .B1(n12118), .B2(n10114), .ZN(
        n9621) );
  XNOR2_X1 U12073 ( .A(n9621), .B(n12132), .ZN(n9622) );
  XOR2_X1 U12074 ( .A(n9623), .B(n9622), .Z(n10100) );
  INV_X1 U12075 ( .A(n9624), .ZN(n10516) );
  NAND2_X1 U12076 ( .A1(n10516), .A2(n9643), .ZN(n9632) );
  INV_X1 U12077 ( .A(n9644), .ZN(n9625) );
  NOR2_X1 U12078 ( .A1(n9632), .A2(n9625), .ZN(n9638) );
  NOR2_X1 U12079 ( .A1(n14724), .A2(n9626), .ZN(n9627) );
  AOI211_X1 U12080 ( .C1(n9629), .C2(n9628), .A(n13740), .B(n10763), .ZN(n9648) );
  INV_X1 U12081 ( .A(n9630), .ZN(n9631) );
  OAI21_X1 U12082 ( .B1(n9632), .B2(n9631), .A(n9639), .ZN(n9636) );
  INV_X1 U12083 ( .A(n9756), .ZN(n9633) );
  NAND3_X1 U12084 ( .A1(n9634), .A2(n9642), .A3(n9633), .ZN(n11992) );
  INV_X1 U12085 ( .A(n11992), .ZN(n9635) );
  NAND2_X1 U12086 ( .A1(n9636), .A2(n9635), .ZN(n10035) );
  MUX2_X1 U12087 ( .A(n13734), .B(P1_U3086), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n9647) );
  INV_X1 U12088 ( .A(n14560), .ZN(n9637) );
  NAND2_X1 U12089 ( .A1(n9638), .A2(n9637), .ZN(n9641) );
  INV_X1 U12090 ( .A(n9639), .ZN(n9640) );
  INV_X1 U12091 ( .A(n6462), .ZN(n13713) );
  OAI22_X1 U12092 ( .A1(n11798), .A2(n13713), .B1(n10136), .B2(n13711), .ZN(
        n10534) );
  INV_X1 U12093 ( .A(n10534), .ZN(n9645) );
  INV_X1 U12094 ( .A(n14552), .ZN(n13736) );
  OAI22_X1 U12095 ( .A1(n13730), .A2(n14703), .B1(n9645), .B2(n13736), .ZN(
        n9646) );
  OR3_X1 U12096 ( .A1(n9648), .A2(n9647), .A3(n9646), .ZN(P1_U3218) );
  NAND2_X1 U12097 ( .A1(n9650), .A2(n9649), .ZN(n9651) );
  NAND2_X1 U12098 ( .A1(n6722), .A2(n9651), .ZN(n9663) );
  INV_X1 U12099 ( .A(n9663), .ZN(n9653) );
  INV_X1 U12100 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10644) );
  MUX2_X1 U12101 ( .A(n10867), .B(n10644), .S(n12516), .Z(n9661) );
  NOR2_X1 U12102 ( .A1(n15067), .A2(n9661), .ZN(n9656) );
  INV_X1 U12103 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n9655) );
  MUX2_X1 U12104 ( .A(n15056), .B(n9656), .S(n9655), .Z(n9670) );
  INV_X1 U12105 ( .A(n9657), .ZN(n9658) );
  INV_X1 U12106 ( .A(n14480), .ZN(n15061) );
  INV_X1 U12107 ( .A(n15058), .ZN(n14998) );
  NAND3_X1 U12108 ( .A1(n15061), .A2(n15067), .A3(n14998), .ZN(n9662) );
  AND2_X1 U12109 ( .A1(n9661), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10474) );
  NAND2_X1 U12110 ( .A1(n9662), .A2(n10474), .ZN(n9668) );
  AOI22_X1 U12111 ( .A1(n15025), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n9667) );
  NAND2_X1 U12112 ( .A1(n14480), .A2(n10429), .ZN(n9666) );
  NOR2_X1 U12113 ( .A1(n10644), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10438) );
  NAND2_X1 U12114 ( .A1(n15058), .A2(n10438), .ZN(n9665) );
  NAND4_X1 U12115 ( .A1(n9668), .A2(n9667), .A3(n9666), .A4(n9665), .ZN(n9669)
         );
  OR2_X1 U12116 ( .A1(n9670), .A2(n9669), .ZN(P3_U3182) );
  NAND2_X2 U12117 ( .A1(n9685), .A2(P2_U3088), .ZN(n13587) );
  NOR2_X1 U12118 ( .A1(n9857), .A2(P2_U3088), .ZN(n14774) );
  AOI21_X1 U12119 ( .B1(n13585), .B2(P1_DATAO_REG_1__SCAN_IN), .A(n14774), 
        .ZN(n9671) );
  OAI21_X1 U12120 ( .B1(n9692), .B2(n13587), .A(n9671), .ZN(P2_U3326) );
  INV_X1 U12121 ( .A(n9672), .ZN(n9679) );
  AND2_X1 U12122 ( .A1(n9863), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14797) );
  AOI21_X1 U12123 ( .B1(n13585), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n14797), 
        .ZN(n9673) );
  OAI21_X1 U12124 ( .B1(n9679), .B2(n13587), .A(n9673), .ZN(P2_U3324) );
  INV_X1 U12125 ( .A(n13585), .ZN(n13599) );
  INV_X1 U12126 ( .A(n14787), .ZN(n9674) );
  OAI222_X1 U12127 ( .A1(n13599), .A2(n9675), .B1(n13587), .B2(n9690), .C1(
        P2_U3088), .C2(n9674), .ZN(P2_U3325) );
  INV_X1 U12128 ( .A(n9676), .ZN(n9695) );
  INV_X1 U12129 ( .A(n9937), .ZN(n9945) );
  OAI222_X1 U12130 ( .A1(n13599), .A2(n9677), .B1(n13587), .B2(n9695), .C1(
        P2_U3088), .C2(n9945), .ZN(P2_U3323) );
  INV_X1 U12131 ( .A(n13809), .ZN(n9680) );
  INV_X2 U12132 ( .A(n14235), .ZN(n14262) );
  OAI222_X1 U12133 ( .A1(P1_U3086), .A2(n9680), .B1(n14262), .B2(n9679), .C1(
        n9678), .C2(n14258), .ZN(P1_U3352) );
  INV_X1 U12134 ( .A(n9681), .ZN(n9697) );
  INV_X1 U12135 ( .A(n14817), .ZN(n9682) );
  OAI222_X1 U12136 ( .A1(n13599), .A2(n9683), .B1(n13587), .B2(n9697), .C1(
        P2_U3088), .C2(n9682), .ZN(P2_U3322) );
  NAND2_X1 U12137 ( .A1(n9685), .A2(P3_U3151), .ZN(n12966) );
  INV_X1 U12138 ( .A(SI_1_), .ZN(n9687) );
  INV_X1 U12139 ( .A(n6737), .ZN(n9686) );
  OAI222_X1 U12140 ( .A1(n6460), .A2(n9688), .B1(n12966), .B2(n9687), .C1(
        P3_U3151), .C2(n9686), .ZN(P3_U3294) );
  INV_X1 U12141 ( .A(n14258), .ZN(n14259) );
  INV_X1 U12142 ( .A(n14259), .ZN(n11694) );
  INV_X1 U12143 ( .A(n13792), .ZN(n9689) );
  OAI222_X1 U12144 ( .A1(n11694), .A2(n9691), .B1(n14262), .B2(n9690), .C1(
        P1_U3086), .C2(n9689), .ZN(P1_U3353) );
  OAI222_X1 U12145 ( .A1(n11694), .A2(n9693), .B1(n14262), .B2(n9692), .C1(
        P1_U3086), .C2(n9796), .ZN(P1_U3354) );
  INV_X1 U12146 ( .A(n13820), .ZN(n9694) );
  OAI222_X1 U12147 ( .A1(n11694), .A2(n9696), .B1(n14262), .B2(n9695), .C1(
        P1_U3086), .C2(n9694), .ZN(P1_U3351) );
  INV_X1 U12148 ( .A(n9801), .ZN(n9823) );
  OAI222_X1 U12149 ( .A1(n11694), .A2(n9698), .B1(n14262), .B2(n9697), .C1(
        P1_U3086), .C2(n9823), .ZN(P1_U3350) );
  INV_X1 U12150 ( .A(n9699), .ZN(n9701) );
  INV_X1 U12151 ( .A(n9805), .ZN(n10017) );
  OAI222_X1 U12152 ( .A1(n11694), .A2(n9700), .B1(n14262), .B2(n9701), .C1(
        P1_U3086), .C2(n10017), .ZN(P1_U3349) );
  INV_X1 U12153 ( .A(n9884), .ZN(n9875) );
  OAI222_X1 U12154 ( .A1(n13599), .A2(n9702), .B1(n13587), .B2(n9701), .C1(
        P2_U3088), .C2(n9875), .ZN(P2_U3321) );
  INV_X1 U12155 ( .A(n6475), .ZN(n10470) );
  INV_X1 U12156 ( .A(n12966), .ZN(n12952) );
  AOI222_X1 U12157 ( .A1(n9703), .A2(n10884), .B1(n10470), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_2_), .C2(n12952), .ZN(n9704) );
  INV_X1 U12158 ( .A(n9704), .ZN(P3_U3293) );
  AOI222_X1 U12159 ( .A1(n9705), .A2(n10884), .B1(SI_7_), .B2(n12952), .C1(
        n11126), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9706) );
  INV_X1 U12160 ( .A(n9706), .ZN(P3_U3288) );
  AOI222_X1 U12161 ( .A1(n9707), .A2(n10884), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15057), .C1(SI_9_), .C2(n12952), .ZN(n9708) );
  INV_X1 U12162 ( .A(n9708), .ZN(P3_U3286) );
  AOI222_X1 U12163 ( .A1(n9709), .A2(n10884), .B1(n14987), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_5_), .C2(n12952), .ZN(n9710) );
  INV_X1 U12164 ( .A(n9710), .ZN(P3_U3290) );
  INV_X1 U12165 ( .A(SI_8_), .ZN(n9711) );
  OAI222_X1 U12166 ( .A1(n6460), .A2(n9712), .B1(n12966), .B2(n9711), .C1(
        P3_U3151), .C2(n11133), .ZN(P3_U3287) );
  AOI222_X1 U12167 ( .A1(n9713), .A2(n10884), .B1(n10502), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_3_), .C2(n12952), .ZN(n9714) );
  INV_X1 U12168 ( .A(n9714), .ZN(P3_U3292) );
  AOI222_X1 U12169 ( .A1(n9715), .A2(n10884), .B1(SI_10_), .B2(n12952), .C1(
        n11144), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9716) );
  INV_X1 U12170 ( .A(n9716), .ZN(P3_U3285) );
  INV_X1 U12171 ( .A(SI_4_), .ZN(n9717) );
  OAI222_X1 U12172 ( .A1(P3_U3151), .A2(n11088), .B1(n6460), .B2(n9718), .C1(
        n9717), .C2(n12966), .ZN(P3_U3291) );
  OAI222_X1 U12173 ( .A1(n11422), .A2(P3_U3151), .B1(n6460), .B2(n9720), .C1(
        n9719), .C2(n12966), .ZN(P3_U3284) );
  INV_X1 U12174 ( .A(SI_6_), .ZN(n9721) );
  OAI222_X1 U12175 ( .A1(n11120), .A2(P3_U3151), .B1(n6461), .B2(n9722), .C1(
        n9721), .C2(n12966), .ZN(P3_U3289) );
  INV_X1 U12176 ( .A(n9723), .ZN(n9725) );
  INV_X1 U12177 ( .A(n9808), .ZN(n13830) );
  OAI222_X1 U12178 ( .A1(n11694), .A2(n9724), .B1(n14262), .B2(n9725), .C1(
        P1_U3086), .C2(n13830), .ZN(P1_U3348) );
  INV_X1 U12179 ( .A(n9920), .ZN(n9932) );
  OAI222_X1 U12180 ( .A1(n13599), .A2(n9726), .B1(n13587), .B2(n9725), .C1(
        P2_U3088), .C2(n9932), .ZN(P2_U3320) );
  INV_X1 U12181 ( .A(n9727), .ZN(n9729) );
  OAI222_X1 U12182 ( .A1(n11589), .A2(P3_U3151), .B1(n6461), .B2(n9729), .C1(
        n9728), .C2(n12966), .ZN(P3_U3283) );
  INV_X1 U12183 ( .A(n9730), .ZN(n9733) );
  INV_X1 U12184 ( .A(n9985), .ZN(n9731) );
  OAI222_X1 U12185 ( .A1(n13599), .A2(n9732), .B1(n13587), .B2(n9733), .C1(
        P2_U3088), .C2(n9731), .ZN(P2_U3319) );
  INV_X1 U12186 ( .A(n9811), .ZN(n9950) );
  OAI222_X1 U12187 ( .A1(n11694), .A2(n9734), .B1(n14262), .B2(n9733), .C1(
        P1_U3086), .C2(n9950), .ZN(P1_U3347) );
  NAND2_X1 U12188 ( .A1(n9735), .A2(n9753), .ZN(n14694) );
  INV_X1 U12189 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9739) );
  INV_X1 U12190 ( .A(n9736), .ZN(n9737) );
  AOI22_X1 U12191 ( .A1(n14694), .A2(n9739), .B1(n9738), .B2(n9737), .ZN(
        P1_U3445) );
  INV_X1 U12192 ( .A(n9740), .ZN(n9742) );
  OAI222_X1 U12193 ( .A1(n13599), .A2(n9741), .B1(n13587), .B2(n9742), .C1(
        P2_U3088), .C2(n10064), .ZN(P2_U3318) );
  INV_X1 U12194 ( .A(n9900), .ZN(n9895) );
  OAI222_X1 U12195 ( .A1(n11694), .A2(n9743), .B1(n14262), .B2(n9742), .C1(
        P1_U3086), .C2(n9895), .ZN(P1_U3346) );
  OAI222_X1 U12196 ( .A1(P3_U3151), .A2(n12469), .B1(n12966), .B2(n9745), .C1(
        n6460), .C2(n9744), .ZN(P3_U3282) );
  INV_X1 U12197 ( .A(n14694), .ZN(n14693) );
  OAI22_X1 U12198 ( .A1(n14693), .A2(P1_D_REG_1__SCAN_IN), .B1(n9747), .B2(
        n9746), .ZN(n9748) );
  INV_X1 U12199 ( .A(n9748), .ZN(P1_U3446) );
  INV_X1 U12200 ( .A(n9749), .ZN(n9751) );
  INV_X1 U12201 ( .A(n9904), .ZN(n9975) );
  OAI222_X1 U12202 ( .A1(n11694), .A2(n9750), .B1(n14262), .B2(n9751), .C1(
        P1_U3086), .C2(n9975), .ZN(P1_U3345) );
  INV_X1 U12203 ( .A(n10050), .ZN(n9996) );
  OAI222_X1 U12204 ( .A1(n13599), .A2(n9752), .B1(n13587), .B2(n9751), .C1(
        P2_U3088), .C2(n9996), .ZN(P2_U3317) );
  INV_X1 U12205 ( .A(n9753), .ZN(n9754) );
  NAND2_X1 U12206 ( .A1(n9756), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11993) );
  NAND2_X1 U12207 ( .A1(n9754), .A2(n11993), .ZN(n9759) );
  OAI21_X1 U12208 ( .B1(n11941), .B2(n9756), .A(n9755), .ZN(n9757) );
  NAND2_X1 U12209 ( .A1(n9759), .A2(n9757), .ZN(n14640) );
  INV_X1 U12210 ( .A(n9757), .ZN(n9758) );
  NAND2_X1 U12211 ( .A1(n9759), .A2(n9758), .ZN(n9792) );
  INV_X1 U12212 ( .A(n9792), .ZN(n9763) );
  NAND3_X1 U12213 ( .A1(n14631), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9760), .ZN(
        n9765) );
  OAI21_X1 U12214 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n14247), .A(n9791), .ZN(
        n13786) );
  AOI21_X1 U12215 ( .B1(n14247), .B2(n9760), .A(n13786), .ZN(n9761) );
  MUX2_X1 U12216 ( .A(n13786), .B(n9761), .S(n13785), .Z(n9762) );
  AOI22_X1 U12217 ( .A1(n9763), .A2(n9762), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9764) );
  OAI211_X1 U12218 ( .C1(n14640), .C2(n6760), .A(n9765), .B(n9764), .ZN(
        P1_U3243) );
  INV_X1 U12219 ( .A(n14640), .ZN(n13877) );
  NOR2_X1 U12220 ( .A1(n13877), .A2(n13788), .ZN(P1_U3085) );
  AND2_X1 U12221 ( .A1(n9767), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12222 ( .A1(n9767), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12223 ( .A1(n9767), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12224 ( .A1(n9767), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12225 ( .A1(n9767), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12226 ( .A1(n9767), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U12227 ( .A1(n9767), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12228 ( .A1(n9767), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12229 ( .A1(n9767), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12230 ( .A1(n9767), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12231 ( .A1(n9767), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12232 ( .A1(n9767), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12233 ( .A1(n9767), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12234 ( .A1(n9767), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12235 ( .A1(n9767), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12236 ( .A1(n9767), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12237 ( .A1(n9767), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12238 ( .A1(n9767), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12239 ( .A1(n9767), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12240 ( .A1(n9767), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12241 ( .A1(n9767), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12242 ( .A1(n9767), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12243 ( .A1(n9767), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12244 ( .A1(n9767), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12245 ( .A1(n9767), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12246 ( .A1(n9767), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12247 ( .A1(n9767), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12248 ( .A1(n9767), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12249 ( .A1(n9767), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12250 ( .A1(n9767), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  INV_X1 U12251 ( .A(n9768), .ZN(n9770) );
  INV_X1 U12252 ( .A(n10148), .ZN(n9910) );
  OAI222_X1 U12253 ( .A1(n11694), .A2(n9769), .B1(n14262), .B2(n9770), .C1(
        P1_U3086), .C2(n9910), .ZN(P1_U3344) );
  INV_X1 U12254 ( .A(n10083), .ZN(n10048) );
  OAI222_X1 U12255 ( .A1(n13599), .A2(n10368), .B1(n13587), .B2(n9770), .C1(
        P2_U3088), .C2(n10048), .ZN(P2_U3316) );
  OAI222_X1 U12256 ( .A1(P3_U3151), .A2(n12494), .B1(n12966), .B2(n9772), .C1(
        n6460), .C2(n9771), .ZN(P3_U3281) );
  NAND2_X1 U12257 ( .A1(n13788), .A2(n10135), .ZN(n9773) );
  OAI21_X1 U12258 ( .B1(n13788), .B2(n8895), .A(n9773), .ZN(P1_U3560) );
  INV_X1 U12259 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9774) );
  MUX2_X1 U12260 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9774), .S(n13792), .Z(
        n13795) );
  MUX2_X1 U12261 ( .A(n9775), .B(P1_REG2_REG_1__SCAN_IN), .S(n9796), .Z(n13774) );
  AND2_X1 U12262 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9776) );
  NAND2_X1 U12263 ( .A1(n13774), .A2(n9776), .ZN(n13773) );
  NAND2_X1 U12264 ( .A1(n13778), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9777) );
  NAND2_X1 U12265 ( .A1(n13773), .A2(n9777), .ZN(n13793) );
  NAND2_X1 U12266 ( .A1(n13795), .A2(n13793), .ZN(n9779) );
  NAND2_X1 U12267 ( .A1(n13792), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9778) );
  NAND2_X1 U12268 ( .A1(n9779), .A2(n9778), .ZN(n13806) );
  MUX2_X1 U12269 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10536), .S(n13809), .Z(
        n13807) );
  NAND2_X1 U12270 ( .A1(n13806), .A2(n13807), .ZN(n13823) );
  NAND2_X1 U12271 ( .A1(n13809), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n13822) );
  NAND2_X1 U12272 ( .A1(n13823), .A2(n13822), .ZN(n9782) );
  MUX2_X1 U12273 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9780), .S(n13820), .Z(n9781) );
  NAND2_X1 U12274 ( .A1(n9782), .A2(n9781), .ZN(n13825) );
  NAND2_X1 U12275 ( .A1(n13820), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9826) );
  MUX2_X1 U12276 ( .A(n9783), .B(P1_REG2_REG_5__SCAN_IN), .S(n9801), .Z(n9825)
         );
  AOI21_X1 U12277 ( .B1(n13825), .B2(n9826), .A(n9825), .ZN(n10010) );
  NOR2_X1 U12278 ( .A1(n9823), .A2(n9783), .ZN(n10009) );
  MUX2_X1 U12279 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9784), .S(n9805), .Z(n10008) );
  OAI21_X1 U12280 ( .B1(n10010), .B2(n10009), .A(n10008), .ZN(n13839) );
  NAND2_X1 U12281 ( .A1(n9805), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n13838) );
  MUX2_X1 U12282 ( .A(n10587), .B(P1_REG2_REG_7__SCAN_IN), .S(n9808), .Z(
        n13837) );
  AOI21_X1 U12283 ( .B1(n13839), .B2(n13838), .A(n13837), .ZN(n13836) );
  NOR2_X1 U12284 ( .A1(n13830), .A2(n10587), .ZN(n9953) );
  MUX2_X1 U12285 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n9785), .S(n9811), .Z(n9952)
         );
  OAI21_X1 U12286 ( .B1(n13836), .B2(n9953), .A(n9952), .ZN(n9951) );
  NAND2_X1 U12287 ( .A1(n9811), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9788) );
  MUX2_X1 U12288 ( .A(n10983), .B(P1_REG2_REG_9__SCAN_IN), .S(n9900), .Z(n9787) );
  AOI21_X1 U12289 ( .B1(n9951), .B2(n9788), .A(n9787), .ZN(n9970) );
  NAND2_X1 U12290 ( .A1(n9791), .A2(n11990), .ZN(n9786) );
  INV_X1 U12291 ( .A(n14627), .ZN(n13879) );
  NAND3_X1 U12292 ( .A1(n9951), .A2(n9788), .A3(n9787), .ZN(n9789) );
  NAND2_X1 U12293 ( .A1(n13879), .A2(n9789), .ZN(n9818) );
  NOR2_X1 U12294 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9790), .ZN(n11404) );
  OR2_X1 U12295 ( .A1(n9792), .A2(n9791), .ZN(n14636) );
  NOR2_X1 U12296 ( .A1(n14636), .A2(n9895), .ZN(n9793) );
  AOI211_X1 U12297 ( .C1(n13877), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n11404), .B(
        n9793), .ZN(n9817) );
  MUX2_X1 U12298 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9794), .S(n9900), .Z(n9814)
         );
  XNOR2_X1 U12299 ( .A(n13792), .B(n9795), .ZN(n13799) );
  XNOR2_X1 U12300 ( .A(n9796), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n13777) );
  AND2_X1 U12301 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n13776) );
  NAND2_X1 U12302 ( .A1(n13777), .A2(n13776), .ZN(n13775) );
  NAND2_X1 U12303 ( .A1(n13778), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9797) );
  NAND2_X1 U12304 ( .A1(n13775), .A2(n9797), .ZN(n13798) );
  NAND2_X1 U12305 ( .A1(n13799), .A2(n13798), .ZN(n13797) );
  NAND2_X1 U12306 ( .A1(n13792), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9798) );
  NAND2_X1 U12307 ( .A1(n13797), .A2(n9798), .ZN(n13804) );
  INV_X1 U12308 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n14757) );
  MUX2_X1 U12309 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n14757), .S(n13809), .Z(
        n13805) );
  NAND2_X1 U12310 ( .A1(n13804), .A2(n13805), .ZN(n13803) );
  NAND2_X1 U12311 ( .A1(n13809), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9799) );
  NAND2_X1 U12312 ( .A1(n13803), .A2(n9799), .ZN(n13818) );
  MUX2_X1 U12313 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n7726), .S(n13820), .Z(
        n13819) );
  NAND2_X1 U12314 ( .A1(n13818), .A2(n13819), .ZN(n13817) );
  NAND2_X1 U12315 ( .A1(n13820), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9800) );
  NAND2_X1 U12316 ( .A1(n13817), .A2(n9800), .ZN(n9821) );
  XNOR2_X1 U12317 ( .A(n9801), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9822) );
  OR2_X1 U12318 ( .A1(n9821), .A2(n9822), .ZN(n9819) );
  NAND2_X1 U12319 ( .A1(n9823), .A2(n9802), .ZN(n9803) );
  NAND2_X1 U12320 ( .A1(n9819), .A2(n9803), .ZN(n10006) );
  MUX2_X1 U12321 ( .A(n9804), .B(P1_REG1_REG_6__SCAN_IN), .S(n9805), .Z(n10007) );
  OR2_X1 U12322 ( .A1(n10006), .A2(n10007), .ZN(n10004) );
  NAND2_X1 U12323 ( .A1(n9805), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9806) );
  NAND2_X1 U12324 ( .A1(n10004), .A2(n9806), .ZN(n13834) );
  INV_X1 U12325 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9807) );
  XNOR2_X1 U12326 ( .A(n9808), .B(n9807), .ZN(n13835) );
  NAND2_X1 U12327 ( .A1(n13834), .A2(n13835), .ZN(n13833) );
  NAND2_X1 U12328 ( .A1(n9808), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9809) );
  AND2_X1 U12329 ( .A1(n13833), .A2(n9809), .ZN(n9948) );
  MUX2_X1 U12330 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9810), .S(n9811), .Z(n9947)
         );
  NAND2_X1 U12331 ( .A1(n9948), .A2(n9947), .ZN(n9946) );
  OR2_X1 U12332 ( .A1(n9811), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9812) );
  NAND2_X1 U12333 ( .A1(n9946), .A2(n9812), .ZN(n9813) );
  NAND2_X1 U12334 ( .A1(n9813), .A2(n9814), .ZN(n9902) );
  OAI21_X1 U12335 ( .B1(n9814), .B2(n9813), .A(n9902), .ZN(n9815) );
  NAND2_X1 U12336 ( .A1(n9815), .A2(n14631), .ZN(n9816) );
  OAI211_X1 U12337 ( .C1(n9970), .C2(n9818), .A(n9817), .B(n9816), .ZN(
        P1_U3252) );
  INV_X1 U12338 ( .A(n9819), .ZN(n9820) );
  AOI21_X1 U12339 ( .B1(n9822), .B2(n9821), .A(n9820), .ZN(n9831) );
  AND2_X1 U12340 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10840) );
  NOR2_X1 U12341 ( .A1(n14636), .A2(n9823), .ZN(n9824) );
  AOI211_X1 U12342 ( .C1(n13877), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n10840), .B(
        n9824), .ZN(n9830) );
  INV_X1 U12343 ( .A(n10010), .ZN(n9828) );
  NAND3_X1 U12344 ( .A1(n13825), .A2(n9826), .A3(n9825), .ZN(n9827) );
  NAND3_X1 U12345 ( .A1(n13879), .A2(n9828), .A3(n9827), .ZN(n9829) );
  OAI211_X1 U12346 ( .C1(n9831), .C2(n13860), .A(n9830), .B(n9829), .ZN(
        P1_U3248) );
  INV_X1 U12347 ( .A(n10218), .ZN(n9834) );
  OAI21_X1 U12348 ( .B1(n9834), .B2(n9833), .A(n9832), .ZN(n9835) );
  AND2_X1 U12349 ( .A1(n9836), .A2(n9835), .ZN(n9837) );
  AND2_X1 U12350 ( .A1(n14798), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14818) );
  AND2_X1 U12351 ( .A1(n9837), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14781) );
  INV_X1 U12352 ( .A(n14781), .ZN(n14825) );
  NOR2_X1 U12353 ( .A1(n10217), .A2(P2_U3088), .ZN(n13584) );
  AND2_X1 U12354 ( .A1(n13584), .A2(n9838), .ZN(n9839) );
  INV_X1 U12355 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10833) );
  MUX2_X1 U12356 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10833), .S(n9863), .Z(
        n14806) );
  INV_X1 U12357 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10898) );
  XNOR2_X1 U12358 ( .A(n14787), .B(n10898), .ZN(n14788) );
  XNOR2_X1 U12359 ( .A(n9857), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n14777) );
  INV_X1 U12360 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n14870) );
  NOR2_X1 U12361 ( .A1(n9840), .A2(n14870), .ZN(n14776) );
  NAND2_X1 U12362 ( .A1(n14777), .A2(n14776), .ZN(n14775) );
  NAND2_X1 U12363 ( .A1(n9859), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9841) );
  NAND2_X1 U12364 ( .A1(n14775), .A2(n9841), .ZN(n14789) );
  NAND2_X1 U12365 ( .A1(n14788), .A2(n14789), .ZN(n9843) );
  NAND2_X1 U12366 ( .A1(n14787), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9842) );
  NAND2_X1 U12367 ( .A1(n9843), .A2(n9842), .ZN(n14807) );
  NAND2_X1 U12368 ( .A1(n14806), .A2(n14807), .ZN(n14805) );
  NAND2_X1 U12369 ( .A1(n9863), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9939) );
  NAND2_X1 U12370 ( .A1(n14805), .A2(n9939), .ZN(n9846) );
  INV_X1 U12371 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9844) );
  MUX2_X1 U12372 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9844), .S(n9937), .Z(n9845)
         );
  NAND2_X1 U12373 ( .A1(n9846), .A2(n9845), .ZN(n9941) );
  NAND2_X1 U12374 ( .A1(n9937), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9847) );
  NAND2_X1 U12375 ( .A1(n9941), .A2(n9847), .ZN(n14822) );
  INV_X1 U12376 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10807) );
  MUX2_X1 U12377 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10807), .S(n14817), .Z(
        n14821) );
  NAND2_X1 U12378 ( .A1(n14822), .A2(n14821), .ZN(n14819) );
  NAND2_X1 U12379 ( .A1(n14817), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9851) );
  NAND2_X1 U12380 ( .A1(n14819), .A2(n9851), .ZN(n9849) );
  INV_X1 U12381 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10816) );
  MUX2_X1 U12382 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10816), .S(n9884), .Z(n9848) );
  NAND2_X1 U12383 ( .A1(n9849), .A2(n9848), .ZN(n9923) );
  MUX2_X1 U12384 ( .A(n10816), .B(P2_REG2_REG_6__SCAN_IN), .S(n9884), .Z(n9850) );
  NAND3_X1 U12385 ( .A1(n14819), .A2(n9851), .A3(n9850), .ZN(n9852) );
  NAND3_X1 U12386 ( .A1(n14820), .A2(n9923), .A3(n9852), .ZN(n9853) );
  OAI21_X1 U12387 ( .B1(n14825), .B2(n7231), .A(n9853), .ZN(n9873) );
  AND2_X1 U12388 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n10753) );
  AND2_X1 U12389 ( .A1(n13584), .A2(n13589), .ZN(n9854) );
  INV_X1 U12390 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n14952) );
  MUX2_X1 U12391 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n14952), .S(n9884), .Z(n9870) );
  INV_X1 U12392 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9856) );
  XNOR2_X1 U12393 ( .A(n14787), .B(n9856), .ZN(n14784) );
  XNOR2_X1 U12394 ( .A(n9857), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n14768) );
  INV_X1 U12395 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n14943) );
  AND2_X1 U12396 ( .A1(n14767), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9858) );
  NAND2_X1 U12397 ( .A1(n14768), .A2(n9858), .ZN(n14769) );
  NAND2_X1 U12398 ( .A1(n9859), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9860) );
  NAND2_X1 U12399 ( .A1(n14769), .A2(n9860), .ZN(n14783) );
  NAND2_X1 U12400 ( .A1(n14784), .A2(n14783), .ZN(n14782) );
  NAND2_X1 U12401 ( .A1(n14787), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9861) );
  NAND2_X1 U12402 ( .A1(n14782), .A2(n9861), .ZN(n14795) );
  INV_X1 U12403 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9862) );
  XNOR2_X1 U12404 ( .A(n9863), .B(n9862), .ZN(n14796) );
  NAND2_X1 U12405 ( .A1(n14795), .A2(n14796), .ZN(n14794) );
  NAND2_X1 U12406 ( .A1(n9863), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9864) );
  NAND2_X1 U12407 ( .A1(n14794), .A2(n9864), .ZN(n9934) );
  INV_X1 U12408 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9865) );
  XNOR2_X1 U12409 ( .A(n9937), .B(n9865), .ZN(n9935) );
  NAND2_X1 U12410 ( .A1(n9934), .A2(n9935), .ZN(n9933) );
  NAND2_X1 U12411 ( .A1(n9937), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9866) );
  NAND2_X1 U12412 ( .A1(n9933), .A2(n9866), .ZN(n14812) );
  INV_X1 U12413 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9867) );
  XNOR2_X1 U12414 ( .A(n14817), .B(n9867), .ZN(n14813) );
  NAND2_X1 U12415 ( .A1(n14812), .A2(n14813), .ZN(n14810) );
  NAND2_X1 U12416 ( .A1(n14817), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9868) );
  NAND2_X1 U12417 ( .A1(n14810), .A2(n9868), .ZN(n9869) );
  NAND2_X1 U12418 ( .A1(n9869), .A2(n9870), .ZN(n9877) );
  OAI21_X1 U12419 ( .B1(n9870), .B2(n9869), .A(n9877), .ZN(n9871) );
  NOR2_X1 U12420 ( .A1(n14803), .A2(n9871), .ZN(n9872) );
  NOR3_X1 U12421 ( .A1(n9873), .A2(n10753), .A3(n9872), .ZN(n9874) );
  OAI21_X1 U12422 ( .B1(n9875), .B2(n11524), .A(n9874), .ZN(P2_U3220) );
  NAND2_X1 U12423 ( .A1(n9884), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9876) );
  NAND2_X1 U12424 ( .A1(n9877), .A2(n9876), .ZN(n9928) );
  INV_X1 U12425 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9878) );
  MUX2_X1 U12426 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9878), .S(n9920), .Z(n9929)
         );
  NAND2_X1 U12427 ( .A1(n9928), .A2(n9929), .ZN(n9927) );
  NAND2_X1 U12428 ( .A1(n9920), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9879) );
  NAND2_X1 U12429 ( .A1(n9927), .A2(n9879), .ZN(n9880) );
  INV_X1 U12430 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n11339) );
  MUX2_X1 U12431 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n11339), .S(n9985), .Z(n9881) );
  AND2_X1 U12432 ( .A1(n9880), .A2(n9881), .ZN(n9980) );
  OAI21_X1 U12433 ( .B1(n9881), .B2(n9880), .A(n14811), .ZN(n9894) );
  INV_X1 U12434 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n9882) );
  NAND2_X1 U12435 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n11066) );
  OAI21_X1 U12436 ( .B1(n14825), .B2(n9882), .A(n11066), .ZN(n9883) );
  AOI21_X1 U12437 ( .B1(n9985), .B2(n14818), .A(n9883), .ZN(n9893) );
  NAND2_X1 U12438 ( .A1(n9884), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9922) );
  NAND2_X1 U12439 ( .A1(n9923), .A2(n9922), .ZN(n9886) );
  INV_X1 U12440 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n14829) );
  MUX2_X1 U12441 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n14829), .S(n9920), .Z(n9885) );
  NAND2_X1 U12442 ( .A1(n9886), .A2(n9885), .ZN(n9925) );
  NAND2_X1 U12443 ( .A1(n9920), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9890) );
  NAND2_X1 U12444 ( .A1(n9925), .A2(n9890), .ZN(n9888) );
  INV_X1 U12445 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10778) );
  MUX2_X1 U12446 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10778), .S(n9985), .Z(n9887) );
  NAND2_X1 U12447 ( .A1(n9888), .A2(n9887), .ZN(n9987) );
  MUX2_X1 U12448 ( .A(n10778), .B(P2_REG2_REG_8__SCAN_IN), .S(n9985), .Z(n9889) );
  NAND3_X1 U12449 ( .A1(n9925), .A2(n9890), .A3(n9889), .ZN(n9891) );
  NAND3_X1 U12450 ( .A1(n14820), .A2(n9987), .A3(n9891), .ZN(n9892) );
  OAI211_X1 U12451 ( .C1(n9980), .C2(n9894), .A(n9893), .B(n9892), .ZN(
        P2_U3222) );
  NOR2_X1 U12452 ( .A1(n9895), .A2(n10983), .ZN(n9969) );
  MUX2_X1 U12453 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11000), .S(n9904), .Z(
        n9968) );
  OAI21_X1 U12454 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(n9967) );
  NAND2_X1 U12455 ( .A1(n9904), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9898) );
  INV_X1 U12456 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9896) );
  MUX2_X1 U12457 ( .A(n9896), .B(P1_REG2_REG_11__SCAN_IN), .S(n10148), .Z(
        n9897) );
  AOI21_X1 U12458 ( .B1(n9967), .B2(n9898), .A(n9897), .ZN(n10143) );
  NAND3_X1 U12459 ( .A1(n9967), .A2(n9898), .A3(n9897), .ZN(n9899) );
  NAND2_X1 U12460 ( .A1(n9899), .A2(n13879), .ZN(n9914) );
  OR2_X1 U12461 ( .A1(n9900), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9901) );
  NAND2_X1 U12462 ( .A1(n9902), .A2(n9901), .ZN(n9965) );
  INV_X1 U12463 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9903) );
  MUX2_X1 U12464 ( .A(n9903), .B(P1_REG1_REG_10__SCAN_IN), .S(n9904), .Z(n9966) );
  OR2_X1 U12465 ( .A1(n9965), .A2(n9966), .ZN(n9963) );
  NAND2_X1 U12466 ( .A1(n9904), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9905) );
  AND2_X1 U12467 ( .A1(n9963), .A2(n9905), .ZN(n9908) );
  MUX2_X1 U12468 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9906), .S(n10148), .Z(
        n9907) );
  NAND2_X1 U12469 ( .A1(n9908), .A2(n9907), .ZN(n10150) );
  OAI21_X1 U12470 ( .B1(n9908), .B2(n9907), .A(n10150), .ZN(n9909) );
  NAND2_X1 U12471 ( .A1(n9909), .A2(n14631), .ZN(n9913) );
  AND2_X1 U12472 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n11655) );
  NOR2_X1 U12473 ( .A1(n14636), .A2(n9910), .ZN(n9911) );
  AOI211_X1 U12474 ( .C1(n13877), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n11655), 
        .B(n9911), .ZN(n9912) );
  OAI211_X1 U12475 ( .C1(n10143), .C2(n9914), .A(n9913), .B(n9912), .ZN(
        P1_U3254) );
  INV_X1 U12476 ( .A(n10556), .ZN(n10092) );
  INV_X1 U12477 ( .A(n9915), .ZN(n9918) );
  OAI222_X1 U12478 ( .A1(P2_U3088), .A2(n10092), .B1(n13587), .B2(n9918), .C1(
        n9916), .C2(n13599), .ZN(P2_U3315) );
  INV_X1 U12479 ( .A(n13854), .ZN(n9917) );
  OAI222_X1 U12480 ( .A1(n11694), .A2(n9919), .B1(n14262), .B2(n9918), .C1(
        n9917), .C2(P1_U3086), .ZN(P1_U3343) );
  AND2_X1 U12481 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10854) );
  MUX2_X1 U12482 ( .A(n14829), .B(P2_REG2_REG_7__SCAN_IN), .S(n9920), .Z(n9921) );
  NAND3_X1 U12483 ( .A1(n9923), .A2(n9922), .A3(n9921), .ZN(n9924) );
  AND3_X1 U12484 ( .A1(n14820), .A2(n9925), .A3(n9924), .ZN(n9926) );
  AOI211_X1 U12485 ( .C1(n14781), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n10854), .B(
        n9926), .ZN(n9931) );
  OAI211_X1 U12486 ( .C1(n9929), .C2(n9928), .A(n14811), .B(n9927), .ZN(n9930)
         );
  OAI211_X1 U12487 ( .C1(n11524), .C2(n9932), .A(n9931), .B(n9930), .ZN(
        P2_U3221) );
  OAI21_X1 U12488 ( .B1(n9935), .B2(n9934), .A(n9933), .ZN(n9936) );
  NAND2_X1 U12489 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n10574) );
  OAI21_X1 U12490 ( .B1(n14803), .B2(n9936), .A(n10574), .ZN(n9943) );
  MUX2_X1 U12491 ( .A(n9844), .B(P2_REG2_REG_4__SCAN_IN), .S(n9937), .Z(n9938)
         );
  NAND3_X1 U12492 ( .A1(n14805), .A2(n9939), .A3(n9938), .ZN(n9940) );
  AND3_X1 U12493 ( .A1(n14820), .A2(n9941), .A3(n9940), .ZN(n9942) );
  AOI211_X1 U12494 ( .C1(n14781), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n9943), .B(
        n9942), .ZN(n9944) );
  OAI21_X1 U12495 ( .B1(n9945), .B2(n11524), .A(n9944), .ZN(P2_U3218) );
  OAI21_X1 U12496 ( .B1(n9948), .B2(n9947), .A(n9946), .ZN(n9958) );
  AND2_X1 U12497 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11356) );
  AOI21_X1 U12498 ( .B1(n13877), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n11356), .ZN(
        n9949) );
  OAI21_X1 U12499 ( .B1(n9950), .B2(n14636), .A(n9949), .ZN(n9957) );
  INV_X1 U12500 ( .A(n9951), .ZN(n9955) );
  NOR3_X1 U12501 ( .A1(n13836), .A2(n9953), .A3(n9952), .ZN(n9954) );
  NOR3_X1 U12502 ( .A1(n9955), .A2(n14627), .A3(n9954), .ZN(n9956) );
  AOI211_X1 U12503 ( .C1(n14631), .C2(n9958), .A(n9957), .B(n9956), .ZN(n9959)
         );
  INV_X1 U12504 ( .A(n9959), .ZN(P1_U3251) );
  INV_X1 U12505 ( .A(n9960), .ZN(n9962) );
  OAI222_X1 U12506 ( .A1(n12540), .A2(P3_U3151), .B1(n6460), .B2(n9962), .C1(
        n9961), .C2(n12966), .ZN(P3_U3280) );
  INV_X1 U12507 ( .A(n9963), .ZN(n9964) );
  AOI211_X1 U12508 ( .C1(n9966), .C2(n9965), .A(n13860), .B(n9964), .ZN(n9978)
         );
  INV_X1 U12509 ( .A(n9967), .ZN(n9972) );
  NOR3_X1 U12510 ( .A1(n9970), .A2(n9969), .A3(n9968), .ZN(n9971) );
  NOR3_X1 U12511 ( .A1(n9972), .A2(n9971), .A3(n14627), .ZN(n9977) );
  INV_X1 U12512 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9973) );
  NOR2_X1 U12513 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9973), .ZN(n11487) );
  AOI21_X1 U12514 ( .B1(n13877), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n11487), 
        .ZN(n9974) );
  OAI21_X1 U12515 ( .B1(n9975), .B2(n14636), .A(n9974), .ZN(n9976) );
  OR3_X1 U12516 ( .A1(n9978), .A2(n9977), .A3(n9976), .ZN(P1_U3253) );
  INV_X1 U12517 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9979) );
  MUX2_X1 U12518 ( .A(n9979), .B(P2_REG1_REG_10__SCAN_IN), .S(n10050), .Z(
        n9984) );
  INV_X1 U12519 ( .A(n10064), .ZN(n9982) );
  INV_X1 U12520 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9981) );
  MUX2_X1 U12521 ( .A(n9981), .B(P2_REG1_REG_9__SCAN_IN), .S(n10064), .Z(
        n10067) );
  NAND2_X1 U12522 ( .A1(n10068), .A2(n10067), .ZN(n10066) );
  OAI21_X1 U12523 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n9982), .A(n10066), .ZN(
        n9983) );
  NOR2_X1 U12524 ( .A1(n9983), .A2(n9984), .ZN(n10049) );
  AOI211_X1 U12525 ( .C1(n9984), .C2(n9983), .A(n14803), .B(n10049), .ZN(n9998) );
  NAND2_X1 U12526 ( .A1(n9985), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9986) );
  NAND2_X1 U12527 ( .A1(n9987), .A2(n9986), .ZN(n10063) );
  INV_X1 U12528 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9988) );
  MUX2_X1 U12529 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n9988), .S(n10064), .Z(
        n10062) );
  OR2_X1 U12530 ( .A1(n10063), .A2(n10062), .ZN(n10060) );
  NAND2_X1 U12531 ( .A1(n10064), .A2(n9988), .ZN(n9989) );
  AND2_X1 U12532 ( .A1(n10060), .A2(n9989), .ZN(n9992) );
  INV_X1 U12533 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9990) );
  MUX2_X1 U12534 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n9990), .S(n10050), .Z(
        n9991) );
  NAND2_X1 U12535 ( .A1(n9992), .A2(n9991), .ZN(n10040) );
  OAI211_X1 U12536 ( .C1(n9992), .C2(n9991), .A(n10040), .B(n14820), .ZN(n9995) );
  NOR2_X1 U12537 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11301), .ZN(n9993) );
  AOI21_X1 U12538 ( .B1(n14781), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n9993), .ZN(
        n9994) );
  OAI211_X1 U12539 ( .C1(n11524), .C2(n9996), .A(n9995), .B(n9994), .ZN(n9997)
         );
  OR2_X1 U12540 ( .A1(n9998), .A2(n9997), .ZN(P2_U3224) );
  AOI22_X1 U12541 ( .A1(n14811), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n14820), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n10001) );
  NOR2_X1 U12542 ( .A1(n14803), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9999) );
  AOI211_X1 U12543 ( .C1(n14820), .C2(n14870), .A(n9999), .B(n14818), .ZN(
        n10000) );
  MUX2_X1 U12544 ( .A(n10001), .B(n10000), .S(n14767), .Z(n10003) );
  AOI22_X1 U12545 ( .A1(n14781), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n10002) );
  NAND2_X1 U12546 ( .A1(n10003), .A2(n10002), .ZN(P2_U3214) );
  INV_X1 U12547 ( .A(n10004), .ZN(n10005) );
  AOI211_X1 U12548 ( .C1(n10007), .C2(n10006), .A(n10005), .B(n13860), .ZN(
        n10014) );
  INV_X1 U12549 ( .A(n13839), .ZN(n10012) );
  NOR3_X1 U12550 ( .A1(n10010), .A2(n10009), .A3(n10008), .ZN(n10011) );
  NOR3_X1 U12551 ( .A1(n14627), .A2(n10012), .A3(n10011), .ZN(n10013) );
  NOR2_X1 U12552 ( .A1(n10014), .A2(n10013), .ZN(n10016) );
  INV_X1 U12553 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n10356) );
  NOR2_X1 U12554 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10356), .ZN(n11165) );
  AOI21_X1 U12555 ( .B1(n13877), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n11165), .ZN(
        n10015) );
  OAI211_X1 U12556 ( .C1(n10017), .C2(n14636), .A(n10016), .B(n10015), .ZN(
        P1_U3249) );
  INV_X1 U12557 ( .A(n10018), .ZN(n10021) );
  INV_X1 U12558 ( .A(n10169), .ZN(n10158) );
  OAI222_X1 U12559 ( .A1(n11694), .A2(n10019), .B1(n14262), .B2(n10021), .C1(
        n10158), .C2(P1_U3086), .ZN(P1_U3342) );
  OAI222_X1 U12560 ( .A1(P2_U3088), .A2(n10656), .B1(n13587), .B2(n10021), 
        .C1(n10020), .C2(n13599), .ZN(P2_U3314) );
  INV_X1 U12561 ( .A(n10022), .ZN(n10024) );
  OAI222_X1 U12562 ( .A1(n12538), .A2(P3_U3151), .B1(n6461), .B2(n10024), .C1(
        n10023), .C2(n12966), .ZN(P3_U3279) );
  NAND2_X1 U12563 ( .A1(n10135), .A2(n10130), .ZN(n11767) );
  AND2_X1 U12564 ( .A1(n11773), .A2(n11767), .ZN(n11953) );
  INV_X1 U12565 ( .A(n11953), .ZN(n10027) );
  OAI21_X1 U12566 ( .B1(n14664), .B2(n14753), .A(n10027), .ZN(n10031) );
  NAND2_X1 U12567 ( .A1(n13772), .A2(n6462), .ZN(n10596) );
  NAND2_X1 U12568 ( .A1(n7679), .A2(n10028), .ZN(n10029) );
  AND2_X1 U12569 ( .A1(n10596), .A2(n10029), .ZN(n10030) );
  AND2_X1 U12570 ( .A1(n10031), .A2(n10030), .ZN(n14695) );
  NAND2_X1 U12571 ( .A1(n14764), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10032) );
  OAI21_X1 U12572 ( .B1(n14764), .B2(n14695), .A(n10032), .ZN(P1_U3528) );
  XOR2_X1 U12573 ( .A(n10033), .B(n10034), .Z(n10038) );
  NOR2_X1 U12574 ( .A1(n13736), .A2(n13711), .ZN(n11357) );
  AOI22_X1 U12575 ( .A1(n11357), .A2(n10135), .B1(n11778), .B2(n14554), .ZN(
        n10037) );
  NAND2_X1 U12576 ( .A1(n14552), .A2(n6462), .ZN(n11490) );
  INV_X1 U12577 ( .A(n11490), .ZN(n10073) );
  OR2_X1 U12578 ( .A1(n10035), .A2(P1_U3086), .ZN(n10102) );
  AOI22_X1 U12579 ( .A1(n10073), .A2(n13771), .B1(n10102), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n10036) );
  OAI211_X1 U12580 ( .C1(n10038), .C2(n13740), .A(n10037), .B(n10036), .ZN(
        P1_U3222) );
  NAND2_X1 U12581 ( .A1(n10050), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10039) );
  NAND2_X1 U12582 ( .A1(n10040), .A2(n10039), .ZN(n10043) );
  INV_X1 U12583 ( .A(n10043), .ZN(n10045) );
  INV_X1 U12584 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10041) );
  MUX2_X1 U12585 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10041), .S(n10083), .Z(
        n10044) );
  MUX2_X1 U12586 ( .A(n10041), .B(P2_REG2_REG_11__SCAN_IN), .S(n10083), .Z(
        n10042) );
  OR2_X1 U12587 ( .A1(n10043), .A2(n10042), .ZN(n10089) );
  OAI21_X1 U12588 ( .B1(n10045), .B2(n10044), .A(n10089), .ZN(n10056) );
  AND2_X1 U12589 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10046) );
  AOI21_X1 U12590 ( .B1(n14781), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n10046), 
        .ZN(n10047) );
  OAI21_X1 U12591 ( .B1(n11524), .B2(n10048), .A(n10047), .ZN(n10055) );
  INV_X1 U12592 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10051) );
  MUX2_X1 U12593 ( .A(n10051), .B(P2_REG1_REG_11__SCAN_IN), .S(n10083), .Z(
        n10052) );
  NOR2_X1 U12594 ( .A1(n10053), .A2(n10052), .ZN(n10079) );
  AOI211_X1 U12595 ( .C1(n10053), .C2(n10052), .A(n14803), .B(n10079), .ZN(
        n10054) );
  AOI211_X1 U12596 ( .C1(n14820), .C2(n10056), .A(n10055), .B(n10054), .ZN(
        n10057) );
  INV_X1 U12597 ( .A(n10057), .ZN(P2_U3225) );
  OAI222_X1 U12598 ( .A1(P3_U3151), .A2(n12543), .B1(n12966), .B2(n10059), 
        .C1(n6461), .C2(n10058), .ZN(P3_U3278) );
  INV_X1 U12599 ( .A(n10060), .ZN(n10061) );
  AOI21_X1 U12600 ( .B1(n10063), .B2(n10062), .A(n10061), .ZN(n10072) );
  INV_X1 U12601 ( .A(n14820), .ZN(n13195) );
  AND2_X1 U12602 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n11234) );
  NOR2_X1 U12603 ( .A1(n11524), .A2(n10064), .ZN(n10065) );
  AOI211_X1 U12604 ( .C1(n14781), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n11234), .B(
        n10065), .ZN(n10071) );
  OAI21_X1 U12605 ( .B1(n10068), .B2(n10067), .A(n10066), .ZN(n10069) );
  NAND2_X1 U12606 ( .A1(n10069), .A2(n14811), .ZN(n10070) );
  OAI211_X1 U12607 ( .C1(n10072), .C2(n13195), .A(n10071), .B(n10070), .ZN(
        P2_U3223) );
  AOI22_X1 U12608 ( .A1(n10073), .A2(n13772), .B1(n10102), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n10078) );
  OAI21_X1 U12609 ( .B1(n10076), .B2(n10075), .A(n10074), .ZN(n13783) );
  AOI22_X1 U12610 ( .A1(n14550), .A2(n13783), .B1(n14554), .B2(n7679), .ZN(
        n10077) );
  NAND2_X1 U12611 ( .A1(n10078), .A2(n10077), .ZN(P1_U3232) );
  INV_X1 U12612 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10080) );
  MUX2_X1 U12613 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n10080), .S(n10556), .Z(
        n10081) );
  NAND2_X1 U12614 ( .A1(n10082), .A2(n10081), .ZN(n10555) );
  OAI21_X1 U12615 ( .B1(n10082), .B2(n10081), .A(n10555), .ZN(n10095) );
  OR2_X1 U12616 ( .A1(n10083), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10087) );
  NAND2_X1 U12617 ( .A1(n10089), .A2(n10087), .ZN(n10085) );
  INV_X1 U12618 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10084) );
  MUX2_X1 U12619 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n10084), .S(n10556), .Z(
        n10086) );
  NAND2_X1 U12620 ( .A1(n10085), .A2(n10086), .ZN(n10551) );
  INV_X1 U12621 ( .A(n10086), .ZN(n10088) );
  NAND3_X1 U12622 ( .A1(n10089), .A2(n10088), .A3(n10087), .ZN(n10090) );
  AOI21_X1 U12623 ( .B1(n10551), .B2(n10090), .A(n13195), .ZN(n10094) );
  NAND2_X1 U12624 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n11530)
         );
  NAND2_X1 U12625 ( .A1(n14781), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n10091) );
  OAI211_X1 U12626 ( .C1(n11524), .C2(n10092), .A(n11530), .B(n10091), .ZN(
        n10093) );
  AOI211_X1 U12627 ( .C1(n10095), .C2(n14811), .A(n10094), .B(n10093), .ZN(
        n10096) );
  INV_X1 U12628 ( .A(n10096), .ZN(P2_U3226) );
  OAI222_X1 U12629 ( .A1(P3_U3151), .A2(n12546), .B1(n12966), .B2(n10098), 
        .C1(n6461), .C2(n10097), .ZN(P3_U3277) );
  XOR2_X1 U12630 ( .A(n10100), .B(n10099), .Z(n10104) );
  AOI22_X1 U12631 ( .A1(n13725), .A2(n13772), .B1(n13770), .B2(n6462), .ZN(
        n10117) );
  OAI22_X1 U12632 ( .A1(n13730), .A2(n14682), .B1(n10117), .B2(n13736), .ZN(
        n10101) );
  AOI21_X1 U12633 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n10102), .A(n10101), .ZN(
        n10103) );
  OAI21_X1 U12634 ( .B1(n10104), .B2(n13740), .A(n10103), .ZN(P1_U3237) );
  INV_X1 U12635 ( .A(n10239), .ZN(n10105) );
  INV_X1 U12636 ( .A(n11176), .ZN(n10665) );
  OAI222_X1 U12637 ( .A1(n13599), .A2(n10106), .B1(n13587), .B2(n10105), .C1(
        P2_U3088), .C2(n10665), .ZN(P2_U3313) );
  INV_X1 U12638 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n10108) );
  NAND2_X1 U12639 ( .A1(n10737), .A2(P3_U3897), .ZN(n10107) );
  OAI21_X1 U12640 ( .B1(P3_U3897), .B2(n10108), .A(n10107), .ZN(P3_U3491) );
  OAI222_X1 U12641 ( .A1(n6461), .A2(n10110), .B1(n12966), .B2(n10109), .C1(
        P3_U3151), .C2(n12523), .ZN(P3_U3276) );
  XNOR2_X1 U12642 ( .A(n10111), .B(n11956), .ZN(n14687) );
  INV_X1 U12643 ( .A(n14724), .ZN(n14749) );
  INV_X1 U12644 ( .A(n10133), .ZN(n10113) );
  INV_X1 U12645 ( .A(n10112), .ZN(n10530) );
  AOI211_X1 U12646 ( .C1(n10114), .C2(n10113), .A(n14674), .B(n10530), .ZN(
        n14685) );
  INV_X1 U12647 ( .A(n14685), .ZN(n10115) );
  OAI21_X1 U12648 ( .B1(n14682), .B2(n14749), .A(n10115), .ZN(n10121) );
  XNOR2_X1 U12649 ( .A(n10116), .B(n11956), .ZN(n10118) );
  OAI21_X1 U12650 ( .B1(n10118), .B2(n14728), .A(n10117), .ZN(n10119) );
  AOI21_X1 U12651 ( .B1(n14687), .B2(n14732), .A(n10119), .ZN(n14691) );
  INV_X1 U12652 ( .A(n14691), .ZN(n10120) );
  AOI211_X1 U12653 ( .C1(n14745), .C2(n14687), .A(n10121), .B(n10120), .ZN(
        n14698) );
  NAND2_X1 U12654 ( .A1(n14764), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n10122) );
  OAI21_X1 U12655 ( .B1(n14698), .B2(n14764), .A(n10122), .ZN(P1_U3530) );
  INV_X1 U12656 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n10388) );
  NAND2_X1 U12657 ( .A1(n14956), .A2(P3_U3897), .ZN(n10123) );
  OAI21_X1 U12658 ( .B1(P3_U3897), .B2(n10388), .A(n10123), .ZN(P3_U3502) );
  INV_X1 U12659 ( .A(n10124), .ZN(n10126) );
  INV_X1 U12660 ( .A(n10918), .ZN(n14635) );
  OAI222_X1 U12661 ( .A1(n11694), .A2(n10125), .B1(n14262), .B2(n10126), .C1(
        P1_U3086), .C2(n14635), .ZN(P1_U3340) );
  INV_X1 U12662 ( .A(n11285), .ZN(n11278) );
  OAI222_X1 U12663 ( .A1(n13599), .A2(n10127), .B1(n13587), .B2(n10126), .C1(
        P2_U3088), .C2(n11278), .ZN(P2_U3312) );
  XOR2_X1 U12664 ( .A(n11954), .B(n10128), .Z(n10549) );
  INV_X1 U12665 ( .A(n10549), .ZN(n10141) );
  AOI21_X1 U12666 ( .B1(n11954), .B2(n10135), .A(n14728), .ZN(n10129) );
  NOR2_X1 U12667 ( .A1(n10129), .A2(n13725), .ZN(n10545) );
  NOR2_X1 U12668 ( .A1(n10131), .A2(n10130), .ZN(n10132) );
  NOR2_X1 U12669 ( .A1(n10133), .A2(n10132), .ZN(n10134) );
  XNOR2_X1 U12670 ( .A(n10134), .B(n13772), .ZN(n10544) );
  NOR3_X1 U12671 ( .A1(n10545), .A2(n14728), .A3(n10544), .ZN(n10140) );
  NAND2_X1 U12672 ( .A1(n10134), .A2(n14655), .ZN(n10540) );
  INV_X1 U12673 ( .A(n10540), .ZN(n10137) );
  OAI22_X1 U12674 ( .A1(n10545), .A2(n7680), .B1(n10136), .B2(n13713), .ZN(
        n10543) );
  AOI211_X1 U12675 ( .C1(n11778), .C2(n14724), .A(n10137), .B(n10543), .ZN(
        n10138) );
  OAI21_X1 U12676 ( .B1(n10549), .B2(n14700), .A(n10138), .ZN(n10139) );
  AOI211_X1 U12677 ( .C1(n14745), .C2(n10141), .A(n10140), .B(n10139), .ZN(
        n14697) );
  NAND2_X1 U12678 ( .A1(n14764), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10142) );
  OAI21_X1 U12679 ( .B1(n14697), .B2(n14764), .A(n10142), .ZN(P1_U3529) );
  AOI21_X1 U12680 ( .B1(n10148), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10143), 
        .ZN(n13846) );
  INV_X1 U12681 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10144) );
  MUX2_X1 U12682 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n10144), .S(n13854), .Z(
        n13847) );
  NAND2_X1 U12683 ( .A1(n13846), .A2(n13847), .ZN(n13845) );
  OAI21_X1 U12684 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n13854), .A(n13845), 
        .ZN(n10146) );
  MUX2_X1 U12685 ( .A(n11321), .B(P1_REG2_REG_13__SCAN_IN), .S(n10169), .Z(
        n10145) );
  NOR2_X1 U12686 ( .A1(n10146), .A2(n10145), .ZN(n10163) );
  AOI211_X1 U12687 ( .C1(n10146), .C2(n10145), .A(n14627), .B(n10163), .ZN(
        n10161) );
  INV_X1 U12688 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10147) );
  MUX2_X1 U12689 ( .A(n10147), .B(P1_REG1_REG_13__SCAN_IN), .S(n10169), .Z(
        n10155) );
  OR2_X1 U12690 ( .A1(n10148), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10149) );
  NAND2_X1 U12691 ( .A1(n10150), .A2(n10149), .ZN(n13851) );
  MUX2_X1 U12692 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10151), .S(n13854), .Z(
        n13852) );
  NAND2_X1 U12693 ( .A1(n13851), .A2(n13852), .ZN(n13850) );
  OR2_X1 U12694 ( .A1(n13854), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10152) );
  NAND2_X1 U12695 ( .A1(n13850), .A2(n10152), .ZN(n10154) );
  OR2_X1 U12696 ( .A1(n10154), .A2(n10155), .ZN(n10171) );
  INV_X1 U12697 ( .A(n10171), .ZN(n10153) );
  AOI211_X1 U12698 ( .C1(n10155), .C2(n10154), .A(n13860), .B(n10153), .ZN(
        n10160) );
  NAND2_X1 U12699 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n11720)
         );
  INV_X1 U12700 ( .A(n11720), .ZN(n10156) );
  AOI21_X1 U12701 ( .B1(n13877), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10156), 
        .ZN(n10157) );
  OAI21_X1 U12702 ( .B1(n10158), .B2(n14636), .A(n10157), .ZN(n10159) );
  OR3_X1 U12703 ( .A1(n10161), .A2(n10160), .A3(n10159), .ZN(P1_U3256) );
  MUX2_X1 U12704 ( .A(n10905), .B(P1_REG2_REG_14__SCAN_IN), .S(n10915), .Z(
        n10164) );
  NAND2_X1 U12705 ( .A1(n10169), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10165) );
  NAND2_X1 U12706 ( .A1(n10164), .A2(n10165), .ZN(n10162) );
  OAI21_X1 U12707 ( .B1(n10163), .B2(n10162), .A(n13879), .ZN(n10178) );
  INV_X1 U12708 ( .A(n10163), .ZN(n10166) );
  AOI21_X1 U12709 ( .B1(n10166), .B2(n10165), .A(n10164), .ZN(n10903) );
  NAND2_X1 U12710 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14555)
         );
  INV_X1 U12711 ( .A(n14555), .ZN(n10168) );
  INV_X1 U12712 ( .A(n10915), .ZN(n10906) );
  NOR2_X1 U12713 ( .A1(n14636), .A2(n10906), .ZN(n10167) );
  AOI211_X1 U12714 ( .C1(n13877), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n10168), 
        .B(n10167), .ZN(n10177) );
  NAND2_X1 U12715 ( .A1(n10169), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10170) );
  AND2_X1 U12716 ( .A1(n10171), .A2(n10170), .ZN(n10174) );
  MUX2_X1 U12717 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10172), .S(n10915), .Z(
        n10173) );
  NAND2_X1 U12718 ( .A1(n10174), .A2(n10173), .ZN(n10917) );
  OAI21_X1 U12719 ( .B1(n10174), .B2(n10173), .A(n10917), .ZN(n10175) );
  NAND2_X1 U12720 ( .A1(n10175), .A2(n14631), .ZN(n10176) );
  OAI211_X1 U12721 ( .C1(n10178), .C2(n10903), .A(n10177), .B(n10176), .ZN(
        P1_U3257) );
  AND2_X1 U12722 ( .A1(n8921), .A2(n10774), .ZN(n10180) );
  INV_X1 U12723 ( .A(n12002), .ZN(n10667) );
  OR2_X2 U12724 ( .A1(n14859), .A2(n10695), .ZN(n10723) );
  NAND2_X1 U12725 ( .A1(n10667), .A2(n10723), .ZN(n12001) );
  OAI21_X1 U12726 ( .B1(n10181), .B2(n8919), .A(n12001), .ZN(n10185) );
  NAND2_X1 U12727 ( .A1(n13182), .A2(n10723), .ZN(n10182) );
  NAND2_X1 U12728 ( .A1(n10183), .A2(n10182), .ZN(n10223) );
  OAI21_X1 U12729 ( .B1(n10183), .B2(n10182), .A(n10223), .ZN(n10184) );
  AOI21_X1 U12730 ( .B1(n10185), .B2(n10184), .A(n10225), .ZN(n10222) );
  XNOR2_X1 U12731 ( .A(n13597), .B(n12174), .ZN(n10186) );
  NAND2_X1 U12732 ( .A1(n10186), .A2(n13595), .ZN(n10187) );
  INV_X1 U12733 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14884) );
  NAND2_X1 U12734 ( .A1(n14874), .A2(n14884), .ZN(n10189) );
  NAND2_X1 U12735 ( .A1(n13595), .A2(n13593), .ZN(n10188) );
  NAND2_X1 U12736 ( .A1(n10189), .A2(n10188), .ZN(n14885) );
  NOR4_X1 U12737 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n10198) );
  INV_X1 U12738 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n14875) );
  INV_X1 U12739 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n14877) );
  INV_X1 U12740 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n14876) );
  INV_X1 U12741 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n14878) );
  NAND4_X1 U12742 ( .A1(n14875), .A2(n14877), .A3(n14876), .A4(n14878), .ZN(
        n10195) );
  NOR4_X1 U12743 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n10193) );
  NOR4_X1 U12744 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n10192) );
  NOR4_X1 U12745 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n10191) );
  NOR4_X1 U12746 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n10190) );
  NAND4_X1 U12747 ( .A1(n10193), .A2(n10192), .A3(n10191), .A4(n10190), .ZN(
        n10194) );
  NOR4_X1 U12748 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n10195), .A4(n10194), .ZN(n10197) );
  NOR4_X1 U12749 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n10196) );
  NAND3_X1 U12750 ( .A1(n10198), .A2(n10197), .A3(n10196), .ZN(n10199) );
  AND2_X1 U12751 ( .A1(n14874), .A2(n10199), .ZN(n10703) );
  INV_X1 U12752 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14880) );
  NAND2_X1 U12753 ( .A1(n14874), .A2(n14880), .ZN(n10202) );
  NOR2_X1 U12754 ( .A1(n13597), .A2(n10200), .ZN(n14881) );
  INV_X1 U12755 ( .A(n14881), .ZN(n10201) );
  OR3_X1 U12756 ( .A1(n14885), .A2(n10703), .A3(n11337), .ZN(n10209) );
  OR2_X1 U12757 ( .A1(n14859), .A2(n13213), .ZN(n10203) );
  NOR2_X1 U12758 ( .A1(n14933), .A2(n10218), .ZN(n10204) );
  INV_X1 U12759 ( .A(n10205), .ZN(n10780) );
  NAND2_X1 U12760 ( .A1(n10215), .A2(n10780), .ZN(n10207) );
  INV_X1 U12761 ( .A(n14859), .ZN(n10206) );
  INV_X1 U12762 ( .A(n10208), .ZN(n10704) );
  NAND2_X1 U12763 ( .A1(n10209), .A2(n10704), .ZN(n10213) );
  NAND2_X1 U12764 ( .A1(n10218), .A2(n10210), .ZN(n10701) );
  AND2_X1 U12765 ( .A1(n10211), .A2(n10701), .ZN(n10212) );
  NAND2_X1 U12766 ( .A1(n10213), .A2(n10212), .ZN(n10411) );
  OR2_X1 U12767 ( .A1(n10411), .A2(P2_U3088), .ZN(n12005) );
  AOI22_X1 U12768 ( .A1(n13149), .A2(n10677), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n12005), .ZN(n10221) );
  NAND2_X1 U12769 ( .A1(n10218), .A2(n10217), .ZN(n13074) );
  INV_X1 U12770 ( .A(n13074), .ZN(n13144) );
  NAND2_X1 U12771 ( .A1(n13144), .A2(n13181), .ZN(n10219) );
  OAI21_X1 U12772 ( .B1(n10216), .B2(n13072), .A(n10219), .ZN(n10876) );
  NAND2_X1 U12773 ( .A1(n13097), .A2(n10876), .ZN(n10220) );
  OAI211_X1 U12774 ( .C1(n10222), .C2(n13151), .A(n10221), .B(n10220), .ZN(
        P2_U3194) );
  INV_X1 U12775 ( .A(n10223), .ZN(n10224) );
  XNOR2_X1 U12776 ( .A(n10181), .B(n14903), .ZN(n10227) );
  NAND2_X1 U12777 ( .A1(n13181), .A2(n12981), .ZN(n10226) );
  NAND2_X1 U12778 ( .A1(n10227), .A2(n10226), .ZN(n10408) );
  OAI21_X1 U12779 ( .B1(n10227), .B2(n10226), .A(n10408), .ZN(n10228) );
  AOI21_X1 U12780 ( .B1(n10229), .B2(n10228), .A(n10410), .ZN(n10234) );
  AOI22_X1 U12781 ( .A1(n13149), .A2(n10900), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n12005), .ZN(n10233) );
  NAND2_X1 U12782 ( .A1(n13144), .A2(n13180), .ZN(n10231) );
  NAND2_X1 U12783 ( .A1(n13182), .A2(n13142), .ZN(n10230) );
  AND2_X1 U12784 ( .A1(n10231), .A2(n10230), .ZN(n10895) );
  OR2_X1 U12785 ( .A1(n13147), .A2(n10895), .ZN(n10232) );
  OAI211_X1 U12786 ( .C1(n10234), .C2(n13151), .A(n10233), .B(n10232), .ZN(
        P2_U3209) );
  INV_X1 U12787 ( .A(n10235), .ZN(n10238) );
  INV_X1 U12788 ( .A(n11615), .ZN(n11628) );
  OAI222_X1 U12789 ( .A1(n14258), .A2(n10236), .B1(n14262), .B2(n10238), .C1(
        n11628), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U12790 ( .A(n11508), .ZN(n11515) );
  OAI222_X1 U12791 ( .A1(P2_U3088), .A2(n11515), .B1(n13587), .B2(n10238), 
        .C1(n10237), .C2(n13599), .ZN(P2_U3311) );
  AOI222_X1 U12792 ( .A1(n10239), .A2(n14235), .B1(P2_DATAO_REG_14__SCAN_IN), 
        .B2(n14259), .C1(P1_STATE_REG_SCAN_IN), .C2(n10915), .ZN(n10407) );
  INV_X1 U12793 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U12794 ( .A1(n7227), .A2(keyinput111), .B1(n10377), .B2(keyinput76), 
        .ZN(n10240) );
  OAI221_X1 U12795 ( .B1(n7227), .B2(keyinput111), .C1(n10377), .C2(keyinput76), .A(n10240), .ZN(n10248) );
  INV_X1 U12796 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n11177) );
  AOI22_X1 U12797 ( .A1(n9810), .A2(keyinput89), .B1(n11177), .B2(keyinput97), 
        .ZN(n10241) );
  OAI221_X1 U12798 ( .B1(n9810), .B2(keyinput89), .C1(n11177), .C2(keyinput97), 
        .A(n10241), .ZN(n10247) );
  XOR2_X1 U12799 ( .A(n6762), .B(keyinput94), .Z(n10245) );
  XOR2_X1 U12800 ( .A(n10356), .B(keyinput121), .Z(n10244) );
  XNOR2_X1 U12801 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput91), .ZN(n10243) );
  XNOR2_X1 U12802 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput72), .ZN(n10242)
         );
  NAND4_X1 U12803 ( .A1(n10245), .A2(n10244), .A3(n10243), .A4(n10242), .ZN(
        n10246) );
  NOR3_X1 U12804 ( .A1(n10248), .A2(n10247), .A3(n10246), .ZN(n10282) );
  AOI22_X1 U12805 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(keyinput79), .B1(n14878), 
        .B2(keyinput82), .ZN(n10249) );
  OAI221_X1 U12806 ( .B1(P3_IR_REG_16__SCAN_IN), .B2(keyinput79), .C1(n14878), 
        .C2(keyinput82), .A(n10249), .ZN(n10257) );
  AOI22_X1 U12807 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput114), .B1(
        P2_D_REG_3__SCAN_IN), .B2(keyinput69), .ZN(n10250) );
  OAI221_X1 U12808 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput114), .C1(
        P2_D_REG_3__SCAN_IN), .C2(keyinput69), .A(n10250), .ZN(n10256) );
  AOI22_X1 U12809 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput66), .B1(
        P2_D_REG_17__SCAN_IN), .B2(keyinput95), .ZN(n10251) );
  OAI221_X1 U12810 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput66), .C1(
        P2_D_REG_17__SCAN_IN), .C2(keyinput95), .A(n10251), .ZN(n10255) );
  XOR2_X1 U12811 ( .A(n8455), .B(keyinput92), .Z(n10253) );
  XNOR2_X1 U12812 ( .A(SI_8_), .B(keyinput120), .ZN(n10252) );
  NAND2_X1 U12813 ( .A1(n10253), .A2(n10252), .ZN(n10254) );
  NOR4_X1 U12814 ( .A1(n10257), .A2(n10256), .A3(n10255), .A4(n10254), .ZN(
        n10281) );
  AOI22_X1 U12815 ( .A1(n10260), .A2(keyinput104), .B1(keyinput102), .B2(
        n10259), .ZN(n10258) );
  OAI221_X1 U12816 ( .B1(n10260), .B2(keyinput104), .C1(n10259), .C2(
        keyinput102), .A(n10258), .ZN(n10268) );
  AOI22_X1 U12817 ( .A1(n8456), .A2(keyinput127), .B1(n13465), .B2(keyinput83), 
        .ZN(n10261) );
  OAI221_X1 U12818 ( .B1(n8456), .B2(keyinput127), .C1(n13465), .C2(keyinput83), .A(n10261), .ZN(n10267) );
  INV_X1 U12819 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15255) );
  AOI22_X1 U12820 ( .A1(n15255), .A2(keyinput70), .B1(n6716), .B2(keyinput65), 
        .ZN(n10262) );
  OAI221_X1 U12821 ( .B1(n15255), .B2(keyinput70), .C1(n6716), .C2(keyinput65), 
        .A(n10262), .ZN(n10266) );
  XNOR2_X1 U12822 ( .A(P1_REG3_REG_9__SCAN_IN), .B(keyinput119), .ZN(n10264)
         );
  XNOR2_X1 U12823 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput109), .ZN(n10263) );
  NAND2_X1 U12824 ( .A1(n10264), .A2(n10263), .ZN(n10265) );
  NOR4_X1 U12825 ( .A1(n10268), .A2(n10267), .A3(n10266), .A4(n10265), .ZN(
        n10280) );
  INV_X1 U12826 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n14692) );
  INV_X1 U12827 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14604) );
  AOI22_X1 U12828 ( .A1(n14692), .A2(keyinput75), .B1(keyinput90), .B2(n14604), 
        .ZN(n10269) );
  OAI221_X1 U12829 ( .B1(n14692), .B2(keyinput75), .C1(n14604), .C2(keyinput90), .A(n10269), .ZN(n10278) );
  INV_X1 U12830 ( .A(P3_B_REG_SCAN_IN), .ZN(n10271) );
  AOI22_X1 U12831 ( .A1(n10271), .A2(keyinput85), .B1(n13076), .B2(keyinput93), 
        .ZN(n10270) );
  OAI221_X1 U12832 ( .B1(n10271), .B2(keyinput85), .C1(n13076), .C2(keyinput93), .A(n10270), .ZN(n10277) );
  XNOR2_X1 U12833 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(keyinput122), .ZN(n10275)
         );
  XNOR2_X1 U12834 ( .A(P3_IR_REG_6__SCAN_IN), .B(keyinput100), .ZN(n10274) );
  XNOR2_X1 U12835 ( .A(P3_REG0_REG_31__SCAN_IN), .B(keyinput77), .ZN(n10273)
         );
  XNOR2_X1 U12836 ( .A(SI_1_), .B(keyinput68), .ZN(n10272) );
  NAND4_X1 U12837 ( .A1(n10275), .A2(n10274), .A3(n10273), .A4(n10272), .ZN(
        n10276) );
  NOR3_X1 U12838 ( .A1(n10278), .A2(n10277), .A3(n10276), .ZN(n10279) );
  AND4_X1 U12839 ( .A1(n10282), .A2(n10281), .A3(n10280), .A4(n10279), .ZN(
        n10405) );
  OAI22_X1 U12840 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(keyinput86), .B1(
        keyinput98), .B2(P1_REG0_REG_23__SCAN_IN), .ZN(n10283) );
  AOI221_X1 U12841 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(keyinput86), .C1(
        P1_REG0_REG_23__SCAN_IN), .C2(keyinput98), .A(n10283), .ZN(n10290) );
  OAI22_X1 U12842 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(keyinput67), .B1(
        keyinput73), .B2(P3_REG1_REG_0__SCAN_IN), .ZN(n10284) );
  AOI221_X1 U12843 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput67), .C1(
        P3_REG1_REG_0__SCAN_IN), .C2(keyinput73), .A(n10284), .ZN(n10289) );
  OAI22_X1 U12844 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(keyinput103), .B1(
        P3_REG0_REG_3__SCAN_IN), .B2(keyinput110), .ZN(n10285) );
  AOI221_X1 U12845 ( .B1(P2_IR_REG_17__SCAN_IN), .B2(keyinput103), .C1(
        keyinput110), .C2(P3_REG0_REG_3__SCAN_IN), .A(n10285), .ZN(n10288) );
  OAI22_X1 U12846 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(keyinput101), .B1(
        keyinput107), .B2(P3_REG0_REG_30__SCAN_IN), .ZN(n10286) );
  AOI221_X1 U12847 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(keyinput101), .C1(
        P3_REG0_REG_30__SCAN_IN), .C2(keyinput107), .A(n10286), .ZN(n10287) );
  NAND4_X1 U12848 ( .A1(n10290), .A2(n10289), .A3(n10288), .A4(n10287), .ZN(
        n10318) );
  OAI22_X1 U12849 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput88), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput78), .ZN(n10291) );
  AOI221_X1 U12850 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput88), .C1(
        keyinput78), .C2(P2_DATAO_REG_21__SCAN_IN), .A(n10291), .ZN(n10298) );
  OAI22_X1 U12851 ( .A1(P2_D_REG_19__SCAN_IN), .A2(keyinput117), .B1(
        keyinput99), .B2(P3_REG0_REG_27__SCAN_IN), .ZN(n10292) );
  AOI221_X1 U12852 ( .B1(P2_D_REG_19__SCAN_IN), .B2(keyinput117), .C1(
        P3_REG0_REG_27__SCAN_IN), .C2(keyinput99), .A(n10292), .ZN(n10297) );
  OAI22_X1 U12853 ( .A1(P3_REG1_REG_29__SCAN_IN), .A2(keyinput80), .B1(
        keyinput64), .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n10293) );
  AOI221_X1 U12854 ( .B1(P3_REG1_REG_29__SCAN_IN), .B2(keyinput80), .C1(
        P1_DATAO_REG_30__SCAN_IN), .C2(keyinput64), .A(n10293), .ZN(n10296) );
  OAI22_X1 U12855 ( .A1(P3_DATAO_REG_4__SCAN_IN), .A2(keyinput112), .B1(
        P3_DATAO_REG_11__SCAN_IN), .B2(keyinput84), .ZN(n10294) );
  AOI221_X1 U12856 ( .B1(P3_DATAO_REG_4__SCAN_IN), .B2(keyinput112), .C1(
        keyinput84), .C2(P3_DATAO_REG_11__SCAN_IN), .A(n10294), .ZN(n10295) );
  NAND4_X1 U12857 ( .A1(n10298), .A2(n10297), .A3(n10296), .A4(n10295), .ZN(
        n10317) );
  OAI22_X1 U12858 ( .A1(P2_REG0_REG_17__SCAN_IN), .A2(keyinput105), .B1(
        keyinput116), .B2(P1_REG3_REG_7__SCAN_IN), .ZN(n10299) );
  AOI221_X1 U12859 ( .B1(P2_REG0_REG_17__SCAN_IN), .B2(keyinput105), .C1(
        P1_REG3_REG_7__SCAN_IN), .C2(keyinput116), .A(n10299), .ZN(n10306) );
  OAI22_X1 U12860 ( .A1(P2_D_REG_0__SCAN_IN), .A2(keyinput115), .B1(
        keyinput123), .B2(SI_31_), .ZN(n10300) );
  AOI221_X1 U12861 ( .B1(P2_D_REG_0__SCAN_IN), .B2(keyinput115), .C1(SI_31_), 
        .C2(keyinput123), .A(n10300), .ZN(n10305) );
  OAI22_X1 U12862 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(keyinput124), .B1(
        P1_REG3_REG_18__SCAN_IN), .B2(keyinput81), .ZN(n10301) );
  AOI221_X1 U12863 ( .B1(P1_ADDR_REG_19__SCAN_IN), .B2(keyinput124), .C1(
        keyinput81), .C2(P1_REG3_REG_18__SCAN_IN), .A(n10301), .ZN(n10304) );
  OAI22_X1 U12864 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(keyinput74), .B1(
        P3_REG1_REG_22__SCAN_IN), .B2(keyinput113), .ZN(n10302) );
  AOI221_X1 U12865 ( .B1(P3_REG3_REG_17__SCAN_IN), .B2(keyinput74), .C1(
        keyinput113), .C2(P3_REG1_REG_22__SCAN_IN), .A(n10302), .ZN(n10303) );
  NAND4_X1 U12866 ( .A1(n10306), .A2(n10305), .A3(n10304), .A4(n10303), .ZN(
        n10316) );
  OAI22_X1 U12867 ( .A1(P1_REG2_REG_26__SCAN_IN), .A2(keyinput126), .B1(
        P1_REG0_REG_13__SCAN_IN), .B2(keyinput106), .ZN(n10307) );
  AOI221_X1 U12868 ( .B1(P1_REG2_REG_26__SCAN_IN), .B2(keyinput126), .C1(
        keyinput106), .C2(P1_REG0_REG_13__SCAN_IN), .A(n10307), .ZN(n10314) );
  OAI22_X1 U12869 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput125), .B1(
        keyinput71), .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10308) );
  AOI221_X1 U12870 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput125), .C1(
        P3_DATAO_REG_30__SCAN_IN), .C2(keyinput71), .A(n10308), .ZN(n10313) );
  OAI22_X1 U12871 ( .A1(P1_D_REG_29__SCAN_IN), .A2(keyinput108), .B1(
        P1_REG1_REG_10__SCAN_IN), .B2(keyinput118), .ZN(n10309) );
  AOI221_X1 U12872 ( .B1(P1_D_REG_29__SCAN_IN), .B2(keyinput108), .C1(
        keyinput118), .C2(P1_REG1_REG_10__SCAN_IN), .A(n10309), .ZN(n10312) );
  OAI22_X1 U12873 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(keyinput96), .B1(keyinput87), .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n10310) );
  AOI221_X1 U12874 ( .B1(P3_IR_REG_1__SCAN_IN), .B2(keyinput96), .C1(
        P3_DATAO_REG_0__SCAN_IN), .C2(keyinput87), .A(n10310), .ZN(n10311) );
  NAND4_X1 U12875 ( .A1(n10314), .A2(n10313), .A3(n10312), .A4(n10311), .ZN(
        n10315) );
  NOR4_X1 U12876 ( .A1(n10318), .A2(n10317), .A3(n10316), .A4(n10315), .ZN(
        n10404) );
  AOI22_X1 U12877 ( .A1(P2_REG1_REG_26__SCAN_IN), .A2(keyinput40), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(keyinput14), .ZN(n10319) );
  OAI221_X1 U12878 ( .B1(P2_REG1_REG_26__SCAN_IN), .B2(keyinput40), .C1(
        P2_DATAO_REG_21__SCAN_IN), .C2(keyinput14), .A(n10319), .ZN(n10326) );
  AOI22_X1 U12879 ( .A1(P3_REG0_REG_3__SCAN_IN), .A2(keyinput46), .B1(
        P2_REG3_REG_8__SCAN_IN), .B2(keyinput24), .ZN(n10320) );
  OAI221_X1 U12880 ( .B1(P3_REG0_REG_3__SCAN_IN), .B2(keyinput46), .C1(
        P2_REG3_REG_8__SCAN_IN), .C2(keyinput24), .A(n10320), .ZN(n10325) );
  AOI22_X1 U12881 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(keyinput10), .B1(
        P3_B_REG_SCAN_IN), .B2(keyinput21), .ZN(n10321) );
  OAI221_X1 U12882 ( .B1(P3_REG3_REG_17__SCAN_IN), .B2(keyinput10), .C1(
        P3_B_REG_SCAN_IN), .C2(keyinput21), .A(n10321), .ZN(n10324) );
  AOI22_X1 U12883 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput45), .B1(
        P2_D_REG_19__SCAN_IN), .B2(keyinput53), .ZN(n10322) );
  OAI221_X1 U12884 ( .B1(P1_IR_REG_8__SCAN_IN), .B2(keyinput45), .C1(
        P2_D_REG_19__SCAN_IN), .C2(keyinput53), .A(n10322), .ZN(n10323) );
  NOR4_X1 U12885 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(n10323), .ZN(
        n10354) );
  AOI22_X1 U12886 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(keyinput22), .B1(
        P1_ADDR_REG_19__SCAN_IN), .B2(keyinput60), .ZN(n10327) );
  OAI221_X1 U12887 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(keyinput22), .C1(
        P1_ADDR_REG_19__SCAN_IN), .C2(keyinput60), .A(n10327), .ZN(n10334) );
  AOI22_X1 U12888 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(keyinput9), .B1(
        P2_REG1_REG_25__SCAN_IN), .B2(keyinput19), .ZN(n10328) );
  OAI221_X1 U12889 ( .B1(P3_REG1_REG_0__SCAN_IN), .B2(keyinput9), .C1(
        P2_REG1_REG_25__SCAN_IN), .C2(keyinput19), .A(n10328), .ZN(n10333) );
  AOI22_X1 U12890 ( .A1(P3_REG0_REG_27__SCAN_IN), .A2(keyinput35), .B1(
        P2_REG0_REG_17__SCAN_IN), .B2(keyinput41), .ZN(n10329) );
  OAI221_X1 U12891 ( .B1(P3_REG0_REG_27__SCAN_IN), .B2(keyinput35), .C1(
        P2_REG0_REG_17__SCAN_IN), .C2(keyinput41), .A(n10329), .ZN(n10332) );
  AOI22_X1 U12892 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(keyinput47), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput61), .ZN(n10330) );
  OAI221_X1 U12893 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(keyinput47), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput61), .A(n10330), .ZN(n10331) );
  NOR4_X1 U12894 ( .A1(n10334), .A2(n10333), .A3(n10332), .A4(n10331), .ZN(
        n10353) );
  AOI22_X1 U12895 ( .A1(P1_REG2_REG_26__SCAN_IN), .A2(keyinput62), .B1(
        P3_D_REG_0__SCAN_IN), .B2(keyinput1), .ZN(n10335) );
  OAI221_X1 U12896 ( .B1(P1_REG2_REG_26__SCAN_IN), .B2(keyinput62), .C1(
        P3_D_REG_0__SCAN_IN), .C2(keyinput1), .A(n10335), .ZN(n10342) );
  AOI22_X1 U12897 ( .A1(P3_REG0_REG_12__SCAN_IN), .A2(keyinput63), .B1(
        P2_IR_REG_17__SCAN_IN), .B2(keyinput39), .ZN(n10336) );
  OAI221_X1 U12898 ( .B1(P3_REG0_REG_12__SCAN_IN), .B2(keyinput63), .C1(
        P2_IR_REG_17__SCAN_IN), .C2(keyinput39), .A(n10336), .ZN(n10341) );
  AOI22_X1 U12899 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(keyinput0), .B1(
        P2_D_REG_3__SCAN_IN), .B2(keyinput5), .ZN(n10337) );
  OAI221_X1 U12900 ( .B1(P1_DATAO_REG_30__SCAN_IN), .B2(keyinput0), .C1(
        P2_D_REG_3__SCAN_IN), .C2(keyinput5), .A(n10337), .ZN(n10340) );
  AOI22_X1 U12901 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(keyinput25), .B1(
        P3_REG1_REG_29__SCAN_IN), .B2(keyinput16), .ZN(n10338) );
  OAI221_X1 U12902 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(keyinput25), .C1(
        P3_REG1_REG_29__SCAN_IN), .C2(keyinput16), .A(n10338), .ZN(n10339) );
  NOR4_X1 U12903 ( .A1(n10342), .A2(n10341), .A3(n10340), .A4(n10339), .ZN(
        n10352) );
  AOI22_X1 U12904 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(keyinput52), .B1(
        P1_RD_REG_SCAN_IN), .B2(keyinput27), .ZN(n10343) );
  OAI221_X1 U12905 ( .B1(P1_REG3_REG_7__SCAN_IN), .B2(keyinput52), .C1(
        P1_RD_REG_SCAN_IN), .C2(keyinput27), .A(n10343), .ZN(n10350) );
  AOI22_X1 U12906 ( .A1(P3_DATAO_REG_4__SCAN_IN), .A2(keyinput48), .B1(
        P1_D_REG_29__SCAN_IN), .B2(keyinput44), .ZN(n10344) );
  OAI221_X1 U12907 ( .B1(P3_DATAO_REG_4__SCAN_IN), .B2(keyinput48), .C1(
        P1_D_REG_29__SCAN_IN), .C2(keyinput44), .A(n10344), .ZN(n10349) );
  AOI22_X1 U12908 ( .A1(P3_DATAO_REG_0__SCAN_IN), .A2(keyinput23), .B1(
        P3_IR_REG_16__SCAN_IN), .B2(keyinput15), .ZN(n10345) );
  OAI221_X1 U12909 ( .B1(P3_DATAO_REG_0__SCAN_IN), .B2(keyinput23), .C1(
        P3_IR_REG_16__SCAN_IN), .C2(keyinput15), .A(n10345), .ZN(n10348) );
  AOI22_X1 U12910 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(keyinput55), .B1(SI_31_), 
        .B2(keyinput59), .ZN(n10346) );
  OAI221_X1 U12911 ( .B1(P1_REG3_REG_9__SCAN_IN), .B2(keyinput55), .C1(SI_31_), 
        .C2(keyinput59), .A(n10346), .ZN(n10347) );
  NOR4_X1 U12912 ( .A1(n10350), .A2(n10349), .A3(n10348), .A4(n10347), .ZN(
        n10351) );
  NAND4_X1 U12913 ( .A1(n10354), .A2(n10353), .A3(n10352), .A4(n10351), .ZN(
        n10403) );
  INV_X1 U12914 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n13715) );
  AOI22_X1 U12915 ( .A1(n13715), .A2(keyinput17), .B1(keyinput57), .B2(n10356), 
        .ZN(n10355) );
  OAI221_X1 U12916 ( .B1(n13715), .B2(keyinput17), .C1(n10356), .C2(keyinput57), .A(n10355), .ZN(n10364) );
  AOI22_X1 U12917 ( .A1(n9903), .A2(keyinput54), .B1(n7876), .B2(keyinput42), 
        .ZN(n10357) );
  OAI221_X1 U12918 ( .B1(n9903), .B2(keyinput54), .C1(n7876), .C2(keyinput42), 
        .A(n10357), .ZN(n10363) );
  INV_X1 U12919 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12846) );
  AOI22_X1 U12920 ( .A1(n11177), .A2(keyinput33), .B1(keyinput49), .B2(n12846), 
        .ZN(n10358) );
  OAI221_X1 U12921 ( .B1(n11177), .B2(keyinput33), .C1(n12846), .C2(keyinput49), .A(n10358), .ZN(n10362) );
  AOI22_X1 U12922 ( .A1(n13106), .A2(keyinput50), .B1(keyinput2), .B2(n10360), 
        .ZN(n10359) );
  OAI221_X1 U12923 ( .B1(n13106), .B2(keyinput50), .C1(n10360), .C2(keyinput2), 
        .A(n10359), .ZN(n10361) );
  NOR4_X1 U12924 ( .A1(n10364), .A2(n10363), .A3(n10362), .A4(n10361), .ZN(
        n10401) );
  AOI22_X1 U12925 ( .A1(n6762), .A2(keyinput30), .B1(n8455), .B2(keyinput28), 
        .ZN(n10365) );
  OAI221_X1 U12926 ( .B1(n6762), .B2(keyinput30), .C1(n8455), .C2(keyinput28), 
        .A(n10365), .ZN(n10374) );
  AOI22_X1 U12927 ( .A1(n14604), .A2(keyinput26), .B1(n14876), .B2(keyinput31), 
        .ZN(n10366) );
  OAI221_X1 U12928 ( .B1(n14604), .B2(keyinput26), .C1(n14876), .C2(keyinput31), .A(n10366), .ZN(n10373) );
  AOI22_X1 U12929 ( .A1(n10368), .A2(keyinput58), .B1(n14880), .B2(keyinput51), 
        .ZN(n10367) );
  OAI221_X1 U12930 ( .B1(n10368), .B2(keyinput58), .C1(n14880), .C2(keyinput51), .A(n10367), .ZN(n10372) );
  XNOR2_X1 U12931 ( .A(P1_REG1_REG_21__SCAN_IN), .B(keyinput38), .ZN(n10370)
         );
  XNOR2_X1 U12932 ( .A(SI_8_), .B(keyinput56), .ZN(n10369) );
  NAND2_X1 U12933 ( .A1(n10370), .A2(n10369), .ZN(n10371) );
  NOR4_X1 U12934 ( .A1(n10374), .A2(n10373), .A3(n10372), .A4(n10371), .ZN(
        n10400) );
  AOI22_X1 U12935 ( .A1(n14878), .A2(keyinput18), .B1(keyinput3), .B2(n11695), 
        .ZN(n10375) );
  OAI221_X1 U12936 ( .B1(n14878), .B2(keyinput18), .C1(n11695), .C2(keyinput3), 
        .A(n10375), .ZN(n10385) );
  XNOR2_X1 U12937 ( .A(n10376), .B(keyinput36), .ZN(n10384) );
  XNOR2_X1 U12938 ( .A(keyinput12), .B(n10377), .ZN(n10383) );
  XNOR2_X1 U12939 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput37), .ZN(n10381) );
  XNOR2_X1 U12940 ( .A(SI_1_), .B(keyinput4), .ZN(n10380) );
  XNOR2_X1 U12941 ( .A(P3_IR_REG_1__SCAN_IN), .B(keyinput32), .ZN(n10379) );
  XNOR2_X1 U12942 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput8), .ZN(n10378) );
  NAND4_X1 U12943 ( .A1(n10381), .A2(n10380), .A3(n10379), .A4(n10378), .ZN(
        n10382) );
  NOR4_X1 U12944 ( .A1(n10385), .A2(n10384), .A3(n10383), .A4(n10382), .ZN(
        n10399) );
  AOI22_X1 U12945 ( .A1(n10388), .A2(keyinput20), .B1(n10387), .B2(keyinput43), 
        .ZN(n10386) );
  OAI221_X1 U12946 ( .B1(n10388), .B2(keyinput20), .C1(n10387), .C2(keyinput43), .A(n10386), .ZN(n10397) );
  INV_X1 U12947 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n10990) );
  AOI22_X1 U12948 ( .A1(n10990), .A2(keyinput7), .B1(n10390), .B2(keyinput34), 
        .ZN(n10389) );
  OAI221_X1 U12949 ( .B1(n10990), .B2(keyinput7), .C1(n10390), .C2(keyinput34), 
        .A(n10389), .ZN(n10396) );
  AOI22_X1 U12950 ( .A1(n10392), .A2(keyinput13), .B1(keyinput11), .B2(n14692), 
        .ZN(n10391) );
  OAI221_X1 U12951 ( .B1(n10392), .B2(keyinput13), .C1(n14692), .C2(keyinput11), .A(n10391), .ZN(n10395) );
  AOI22_X1 U12952 ( .A1(n15255), .A2(keyinput6), .B1(n13076), .B2(keyinput29), 
        .ZN(n10393) );
  OAI221_X1 U12953 ( .B1(n15255), .B2(keyinput6), .C1(n13076), .C2(keyinput29), 
        .A(n10393), .ZN(n10394) );
  NOR4_X1 U12954 ( .A1(n10397), .A2(n10396), .A3(n10395), .A4(n10394), .ZN(
        n10398) );
  NAND4_X1 U12955 ( .A1(n10401), .A2(n10400), .A3(n10399), .A4(n10398), .ZN(
        n10402) );
  AOI211_X1 U12956 ( .C1(n10405), .C2(n10404), .A(n10403), .B(n10402), .ZN(
        n10406) );
  XNOR2_X1 U12957 ( .A(n10407), .B(n10406), .ZN(P1_U3341) );
  INV_X1 U12958 ( .A(n10408), .ZN(n10409) );
  XNOR2_X1 U12959 ( .A(n10181), .B(n14909), .ZN(n10567) );
  NAND2_X1 U12960 ( .A1(n13180), .A2(n12981), .ZN(n10566) );
  XNOR2_X1 U12961 ( .A(n10567), .B(n10566), .ZN(n10569) );
  XNOR2_X1 U12962 ( .A(n10570), .B(n10569), .ZN(n10414) );
  INV_X1 U12963 ( .A(n13181), .ZN(n10682) );
  INV_X1 U12964 ( .A(n13179), .ZN(n10689) );
  OAI22_X1 U12965 ( .A1(n10682), .A2(n13072), .B1(n10689), .B2(n13074), .ZN(
        n10831) );
  AND2_X1 U12966 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n14799) );
  NAND2_X1 U12967 ( .A1(n10411), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13104) );
  OAI22_X1 U12968 ( .A1(n13137), .A2(n10827), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13104), .ZN(n10412) );
  AOI211_X1 U12969 ( .C1(n13097), .C2(n10831), .A(n14799), .B(n10412), .ZN(
        n10413) );
  OAI21_X1 U12970 ( .B1(n10414), .B2(n13151), .A(n10413), .ZN(P2_U3190) );
  AOI22_X1 U12971 ( .A1(n12422), .A2(n12463), .B1(n14965), .B2(n10870), .ZN(
        n10416) );
  NAND2_X1 U12972 ( .A1(n14971), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10795) );
  NAND2_X1 U12973 ( .A1(n10795), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10415) );
  OAI211_X1 U12974 ( .C1(n10602), .C2(n12433), .A(n10416), .B(n10415), .ZN(
        P3_U3172) );
  MUX2_X1 U12975 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12516), .Z(n11110) );
  INV_X1 U12976 ( .A(n11088), .ZN(n11111) );
  XNOR2_X1 U12977 ( .A(n11110), .B(n11111), .ZN(n11108) );
  MUX2_X1 U12978 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n12516), .Z(n10417) );
  XNOR2_X1 U12979 ( .A(n10417), .B(n6737), .ZN(n10473) );
  NAND2_X1 U12980 ( .A1(n10473), .A2(n10474), .ZN(n10420) );
  INV_X1 U12981 ( .A(n10417), .ZN(n10418) );
  NAND2_X1 U12982 ( .A1(n10418), .A2(n6737), .ZN(n10419) );
  NAND2_X1 U12983 ( .A1(n10420), .A2(n10419), .ZN(n10457) );
  MUX2_X1 U12984 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12516), .Z(n10421) );
  XNOR2_X1 U12985 ( .A(n10421), .B(n10470), .ZN(n10458) );
  NAND2_X1 U12986 ( .A1(n10457), .A2(n10458), .ZN(n10424) );
  INV_X1 U12987 ( .A(n10421), .ZN(n10422) );
  NAND2_X1 U12988 ( .A1(n10422), .A2(n10470), .ZN(n10423) );
  NAND2_X1 U12989 ( .A1(n10424), .A2(n10423), .ZN(n10489) );
  MUX2_X1 U12990 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12516), .Z(n10425) );
  XNOR2_X1 U12991 ( .A(n10425), .B(n10502), .ZN(n10490) );
  NAND2_X1 U12992 ( .A1(n10489), .A2(n10490), .ZN(n10428) );
  INV_X1 U12993 ( .A(n10425), .ZN(n10426) );
  NAND2_X1 U12994 ( .A1(n10426), .A2(n10502), .ZN(n10427) );
  NAND2_X1 U12995 ( .A1(n10428), .A2(n10427), .ZN(n11109) );
  XOR2_X1 U12996 ( .A(n11108), .B(n11109), .Z(n10456) );
  INV_X1 U12997 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15206) );
  INV_X1 U12998 ( .A(n10429), .ZN(n10430) );
  NAND2_X1 U12999 ( .A1(n10486), .A2(n10430), .ZN(n10431) );
  NAND2_X1 U13000 ( .A1(n10461), .A2(n10460), .ZN(n10459) );
  NAND2_X1 U13001 ( .A1(n6475), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10433) );
  INV_X1 U13002 ( .A(n10502), .ZN(n10445) );
  AOI22_X1 U13003 ( .A1(n11111), .A2(P3_REG2_REG_4__SCAN_IN), .B1(n11332), 
        .B2(n11088), .ZN(n10436) );
  AOI21_X1 U13004 ( .B1(n10437), .B2(n10436), .A(n11087), .ZN(n10453) );
  AND2_X1 U13005 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n11220) );
  AOI21_X1 U13006 ( .B1(n15025), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n11220), .ZN(
        n10452) );
  INV_X1 U13007 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15259) );
  AOI22_X1 U13008 ( .A1(n11111), .A2(n15259), .B1(P3_REG1_REG_4__SCAN_IN), 
        .B2(n11088), .ZN(n10449) );
  XNOR2_X1 U13009 ( .A(n6475), .B(n15255), .ZN(n10464) );
  INV_X1 U13010 ( .A(n10438), .ZN(n10439) );
  NAND2_X1 U13011 ( .A1(n6737), .A2(n10439), .ZN(n10440) );
  OR3_X1 U13012 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n10644), .ZN(n10441) );
  NAND2_X1 U13013 ( .A1(n10440), .A2(n10441), .ZN(n10478) );
  INV_X1 U13014 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10477) );
  NAND2_X1 U13015 ( .A1(n10480), .A2(n10441), .ZN(n10463) );
  NAND2_X1 U13016 ( .A1(n10464), .A2(n10463), .ZN(n10444) );
  NAND2_X1 U13017 ( .A1(n6475), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10443) );
  NAND2_X1 U13018 ( .A1(n10444), .A2(n10443), .ZN(n10446) );
  NAND2_X1 U13019 ( .A1(n10446), .A2(n10445), .ZN(n10447) );
  XNOR2_X1 U13020 ( .A(n10446), .B(n10502), .ZN(n10496) );
  NAND2_X1 U13021 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(n10496), .ZN(n10495) );
  NAND2_X1 U13022 ( .A1(n10447), .A2(n10495), .ZN(n10448) );
  NAND2_X1 U13023 ( .A1(n10449), .A2(n10448), .ZN(n11095) );
  OAI21_X1 U13024 ( .B1(n10449), .B2(n10448), .A(n11095), .ZN(n10450) );
  NAND2_X1 U13025 ( .A1(n15058), .A2(n10450), .ZN(n10451) );
  OAI211_X1 U13026 ( .C1(n15061), .C2(n10453), .A(n10452), .B(n10451), .ZN(
        n10454) );
  AOI21_X1 U13027 ( .B1(n11111), .B2(n15056), .A(n10454), .ZN(n10455) );
  OAI21_X1 U13028 ( .B1(n10456), .B2(n15067), .A(n10455), .ZN(P3_U3186) );
  XOR2_X1 U13029 ( .A(n10458), .B(n10457), .Z(n10472) );
  OAI21_X1 U13030 ( .B1(n10461), .B2(n10460), .A(n10459), .ZN(n10462) );
  NAND2_X1 U13031 ( .A1(n14480), .A2(n10462), .ZN(n10468) );
  XNOR2_X1 U13032 ( .A(n10464), .B(n10463), .ZN(n10465) );
  NAND2_X1 U13033 ( .A1(n15058), .A2(n10465), .ZN(n10467) );
  AOI22_X1 U13034 ( .A1(n15025), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10466) );
  NAND3_X1 U13035 ( .A1(n10468), .A2(n10467), .A3(n10466), .ZN(n10469) );
  AOI21_X1 U13036 ( .B1(n10470), .B2(n15056), .A(n10469), .ZN(n10471) );
  OAI21_X1 U13037 ( .B1(n10472), .B2(n15067), .A(n10471), .ZN(P3_U3184) );
  XOR2_X1 U13038 ( .A(n10474), .B(n10473), .Z(n10488) );
  OAI21_X1 U13039 ( .B1(n6602), .B2(P3_REG2_REG_1__SCAN_IN), .A(n10475), .ZN(
        n10476) );
  NAND2_X1 U13040 ( .A1(n14480), .A2(n10476), .ZN(n10484) );
  NAND2_X1 U13041 ( .A1(n10478), .A2(n10477), .ZN(n10479) );
  NAND2_X1 U13042 ( .A1(n10480), .A2(n10479), .ZN(n10481) );
  NAND2_X1 U13043 ( .A1(n15058), .A2(n10481), .ZN(n10483) );
  AOI22_X1 U13044 ( .A1(n15025), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10482) );
  NAND3_X1 U13045 ( .A1(n10484), .A2(n10483), .A3(n10482), .ZN(n10485) );
  AOI21_X1 U13046 ( .B1(n6737), .B2(n15056), .A(n10485), .ZN(n10487) );
  OAI21_X1 U13047 ( .B1(n15067), .B2(n10488), .A(n10487), .ZN(P3_U3183) );
  XOR2_X1 U13048 ( .A(n10490), .B(n10489), .Z(n10504) );
  AOI21_X1 U13049 ( .B1(n10492), .B2(n8313), .A(n10491), .ZN(n10493) );
  INV_X1 U13050 ( .A(n10493), .ZN(n10494) );
  NAND2_X1 U13051 ( .A1(n14480), .A2(n10494), .ZN(n10500) );
  OAI21_X1 U13052 ( .B1(n10496), .B2(P3_REG1_REG_3__SCAN_IN), .A(n10495), .ZN(
        n10497) );
  NAND2_X1 U13053 ( .A1(n15058), .A2(n10497), .ZN(n10499) );
  AOI22_X1 U13054 ( .A1(n15025), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n10498) );
  NAND3_X1 U13055 ( .A1(n10500), .A2(n10499), .A3(n10498), .ZN(n10501) );
  AOI21_X1 U13056 ( .B1(n10502), .B2(n15056), .A(n10501), .ZN(n10503) );
  OAI21_X1 U13057 ( .B1(n10504), .B2(n15067), .A(n10503), .ZN(P3_U3185) );
  INV_X1 U13058 ( .A(n10505), .ZN(n10507) );
  INV_X1 U13059 ( .A(n11623), .ZN(n13865) );
  OAI222_X1 U13060 ( .A1(n11694), .A2(n10506), .B1(n14262), .B2(n10507), .C1(
        n13865), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U13061 ( .A(n13188), .ZN(n13184) );
  OAI222_X1 U13062 ( .A1(n13599), .A2(n10508), .B1(n13587), .B2(n10507), .C1(
        n13184), .C2(P2_U3088), .ZN(P2_U3310) );
  XNOR2_X1 U13063 ( .A(n10509), .B(n10513), .ZN(n10617) );
  OR2_X1 U13064 ( .A1(n11798), .A2(n13711), .ZN(n10511) );
  NAND2_X1 U13065 ( .A1(n13767), .A2(n6462), .ZN(n10510) );
  NAND2_X1 U13066 ( .A1(n10511), .A2(n10510), .ZN(n10841) );
  XNOR2_X1 U13067 ( .A(n10512), .B(n10513), .ZN(n10514) );
  NOR2_X1 U13068 ( .A1(n10514), .A2(n14728), .ZN(n10515) );
  AOI211_X1 U13069 ( .C1(n14732), .C2(n10617), .A(n10841), .B(n10515), .ZN(
        n10619) );
  NAND2_X1 U13070 ( .A1(n10517), .A2(n10516), .ZN(n13903) );
  OR2_X1 U13071 ( .A1(n10518), .A2(n14564), .ZN(n11942) );
  INV_X1 U13072 ( .A(n13988), .ZN(n14688) );
  NOR2_X1 U13073 ( .A1(n14667), .A2(n10844), .ZN(n10519) );
  AOI21_X1 U13074 ( .B1(n6476), .B2(P1_REG2_REG_5__SCAN_IN), .A(n10519), .ZN(
        n10524) );
  INV_X1 U13075 ( .A(n13903), .ZN(n10520) );
  AOI21_X1 U13076 ( .B1(n14673), .B2(n11804), .A(n14674), .ZN(n10521) );
  NAND2_X1 U13077 ( .A1(n10521), .A2(n14653), .ZN(n10618) );
  INV_X1 U13078 ( .A(n10618), .ZN(n10522) );
  NAND2_X1 U13079 ( .A1(n14686), .A2(n10522), .ZN(n10523) );
  OAI211_X1 U13080 ( .C1(n14683), .C2(n6699), .A(n10524), .B(n10523), .ZN(
        n10525) );
  AOI21_X1 U13081 ( .B1(n14688), .B2(n10617), .A(n10525), .ZN(n10526) );
  OAI21_X1 U13082 ( .B1(n10619), .B2(n6476), .A(n10526), .ZN(P1_U3288) );
  XNOR2_X1 U13083 ( .A(n10528), .B(n11789), .ZN(n14699) );
  INV_X1 U13084 ( .A(n10529), .ZN(n14675) );
  OAI211_X1 U13085 ( .C1(n14703), .C2(n10530), .A(n14675), .B(n14655), .ZN(
        n14701) );
  OAI22_X1 U13086 ( .A1(n14090), .A2(n14701), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14667), .ZN(n10531) );
  AOI21_X1 U13087 ( .B1(n14398), .B2(n10532), .A(n10531), .ZN(n10538) );
  XNOR2_X1 U13088 ( .A(n10533), .B(n11789), .ZN(n10535) );
  AOI21_X1 U13089 ( .B1(n10535), .B2(n14664), .A(n10534), .ZN(n14702) );
  MUX2_X1 U13090 ( .A(n14702), .B(n10536), .S(n6476), .Z(n10537) );
  OAI211_X1 U13091 ( .C1(n14077), .C2(n14699), .A(n10538), .B(n10537), .ZN(
        P1_U3290) );
  NOR2_X1 U13092 ( .A1(n14389), .A2(n9775), .ZN(n10542) );
  OAI22_X1 U13093 ( .A1(n14090), .A2(n10540), .B1(n10539), .B2(n14667), .ZN(
        n10541) );
  AOI211_X1 U13094 ( .C1(n14389), .C2(n10543), .A(n10542), .B(n10541), .ZN(
        n10548) );
  NOR3_X1 U13095 ( .A1(n14050), .A2(n10545), .A3(n10544), .ZN(n10546) );
  AOI21_X1 U13096 ( .B1(n14398), .B2(n11778), .A(n10546), .ZN(n10547) );
  OAI211_X1 U13097 ( .C1(n14077), .C2(n10549), .A(n10548), .B(n10547), .ZN(
        P1_U3292) );
  INV_X1 U13098 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10657) );
  MUX2_X1 U13099 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n10657), .S(n10656), .Z(
        n10654) );
  OR2_X1 U13100 ( .A1(n10556), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n10550) );
  NAND2_X1 U13101 ( .A1(n10551), .A2(n10550), .ZN(n10653) );
  XOR2_X1 U13102 ( .A(n10654), .B(n10653), .Z(n10561) );
  NOR2_X1 U13103 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11706), .ZN(n10552) );
  AOI21_X1 U13104 ( .B1(n14781), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n10552), 
        .ZN(n10553) );
  OAI21_X1 U13105 ( .B1(n11524), .B2(n10656), .A(n10553), .ZN(n10560) );
  INV_X1 U13106 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10554) );
  MUX2_X1 U13107 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n10554), .S(n10656), .Z(
        n10558) );
  OAI21_X1 U13108 ( .B1(n10556), .B2(P2_REG1_REG_12__SCAN_IN), .A(n10555), 
        .ZN(n10557) );
  NOR2_X1 U13109 ( .A1(n10557), .A2(n10558), .ZN(n10647) );
  AOI211_X1 U13110 ( .C1(n10558), .C2(n10557), .A(n14803), .B(n10647), .ZN(
        n10559) );
  AOI211_X1 U13111 ( .C1(n14820), .C2(n10561), .A(n10560), .B(n10559), .ZN(
        n10562) );
  INV_X1 U13112 ( .A(n10562), .ZN(P2_U3227) );
  OAI222_X1 U13113 ( .A1(n6461), .A2(n10565), .B1(n12966), .B2(n10564), .C1(
        P3_U3151), .C2(n10563), .ZN(P3_U3275) );
  INV_X1 U13114 ( .A(n10566), .ZN(n10568) );
  INV_X2 U13115 ( .A(n14525), .ZN(n14849) );
  AND2_X1 U13116 ( .A1(n13179), .A2(n14849), .ZN(n10572) );
  XNOR2_X1 U13117 ( .A(n10181), .B(n14850), .ZN(n10571) );
  NOR2_X1 U13118 ( .A1(n10571), .A2(n10572), .ZN(n10744) );
  AOI21_X1 U13119 ( .B1(n10572), .B2(n10571), .A(n10744), .ZN(n10573) );
  OAI21_X1 U13120 ( .B1(n6601), .B2(n10573), .A(n10746), .ZN(n10577) );
  AOI22_X1 U13121 ( .A1(n13144), .A2(n13178), .B1(n13180), .B2(n13142), .ZN(
        n14841) );
  INV_X1 U13122 ( .A(n13104), .ZN(n13145) );
  AOI22_X1 U13123 ( .A1(n13149), .A2(n14850), .B1(n14845), .B2(n13145), .ZN(
        n10575) );
  OAI211_X1 U13124 ( .C1(n14841), .C2(n13147), .A(n10575), .B(n10574), .ZN(
        n10576) );
  AOI21_X1 U13125 ( .B1(n10577), .B2(n13129), .A(n10576), .ZN(n10578) );
  INV_X1 U13126 ( .A(n10578), .ZN(P2_U3202) );
  INV_X1 U13127 ( .A(n10579), .ZN(n10580) );
  AOI21_X1 U13128 ( .B1(n10582), .B2(n10581), .A(n10580), .ZN(n14729) );
  INV_X1 U13129 ( .A(n11008), .ZN(n10584) );
  AOI21_X1 U13130 ( .B1(n14654), .B2(n14725), .A(n14674), .ZN(n10583) );
  NAND2_X1 U13131 ( .A1(n10584), .A2(n10583), .ZN(n14726) );
  NOR2_X1 U13132 ( .A1(n14090), .A2(n14726), .ZN(n10591) );
  NAND2_X1 U13133 ( .A1(n13725), .A2(n13767), .ZN(n10586) );
  NAND2_X1 U13134 ( .A1(n13765), .A2(n6462), .ZN(n10585) );
  NAND2_X1 U13135 ( .A1(n10586), .A2(n10585), .ZN(n14723) );
  INV_X1 U13136 ( .A(n14723), .ZN(n10588) );
  MUX2_X1 U13137 ( .A(n10588), .B(n10587), .S(n6476), .Z(n10589) );
  OAI21_X1 U13138 ( .B1(n14667), .B2(n11274), .A(n10589), .ZN(n10590) );
  AOI211_X1 U13139 ( .C1(n14398), .C2(n14725), .A(n10591), .B(n10590), .ZN(
        n10594) );
  XNOR2_X1 U13140 ( .A(n10592), .B(n11960), .ZN(n14722) );
  INV_X1 U13141 ( .A(n14722), .ZN(n14733) );
  INV_X1 U13142 ( .A(n14077), .ZN(n14677) );
  NAND2_X1 U13143 ( .A1(n14733), .A2(n14677), .ZN(n10593) );
  OAI211_X1 U13144 ( .C1(n14729), .C2(n14050), .A(n10594), .B(n10593), .ZN(
        P1_U3286) );
  NOR2_X1 U13145 ( .A1(n14677), .A2(n14055), .ZN(n10600) );
  NOR2_X1 U13146 ( .A1(n14090), .A2(n14674), .ZN(n14025) );
  OAI21_X1 U13147 ( .B1(n14025), .B2(n14398), .A(n7679), .ZN(n10599) );
  OAI22_X1 U13148 ( .A1(n6476), .A2(n10596), .B1(n10595), .B2(n14667), .ZN(
        n10597) );
  AOI21_X1 U13149 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n6476), .A(n10597), .ZN(
        n10598) );
  OAI211_X1 U13150 ( .C1(n11953), .C2(n10600), .A(n10599), .B(n10598), .ZN(
        P1_U3293) );
  NAND2_X1 U13151 ( .A1(n10606), .A2(n15219), .ZN(n10601) );
  OR2_X1 U13152 ( .A1(n10602), .A2(n10601), .ZN(n10604) );
  NAND2_X1 U13153 ( .A1(n12463), .A2(n15142), .ZN(n10603) );
  AND2_X1 U13154 ( .A1(n10604), .A2(n10603), .ZN(n10868) );
  NAND2_X1 U13155 ( .A1(n10606), .A2(n10605), .ZN(n10607) );
  NAND2_X1 U13156 ( .A1(n10608), .A2(n10607), .ZN(n10609) );
  OAI21_X1 U13157 ( .B1(n10611), .B2(n10610), .A(n10609), .ZN(n10612) );
  AOI22_X1 U13158 ( .A1(n12910), .A2(n10870), .B1(n15252), .B2(
        P3_REG0_REG_0__SCAN_IN), .ZN(n10613) );
  OAI21_X1 U13159 ( .B1(n10868), .B2(n15252), .A(n10613), .ZN(P3_U3390) );
  INV_X1 U13160 ( .A(SI_21_), .ZN(n10615) );
  OAI222_X1 U13161 ( .A1(n6461), .A2(n10616), .B1(n12966), .B2(n10615), .C1(
        P3_U3151), .C2(n10614), .ZN(P3_U3274) );
  INV_X1 U13162 ( .A(n10617), .ZN(n10620) );
  OAI211_X1 U13163 ( .C1(n10620), .C2(n14721), .A(n10619), .B(n10618), .ZN(
        n10625) );
  NAND2_X1 U13164 ( .A1(n10625), .A2(n14766), .ZN(n10622) );
  INV_X1 U13165 ( .A(n14190), .ZN(n14162) );
  NAND2_X1 U13166 ( .A1(n14162), .A2(n11804), .ZN(n10621) );
  OAI211_X1 U13167 ( .C1(n14766), .C2(n9802), .A(n10622), .B(n10621), .ZN(
        P1_U3533) );
  INV_X1 U13168 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10623) );
  OAI22_X1 U13169 ( .A1(n14232), .A2(n6699), .B1(n14756), .B2(n10623), .ZN(
        n10624) );
  AOI21_X1 U13170 ( .B1(n10625), .B2(n14756), .A(n10624), .ZN(n10626) );
  INV_X1 U13171 ( .A(n10626), .ZN(P1_U3474) );
  INV_X1 U13172 ( .A(n13204), .ZN(n13197) );
  OAI222_X1 U13173 ( .A1(n13599), .A2(n10627), .B1(n13587), .B2(n10628), .C1(
        n13197), .C2(P2_U3088), .ZN(P2_U3309) );
  INV_X1 U13174 ( .A(n11629), .ZN(n13874) );
  OAI222_X1 U13175 ( .A1(n11694), .A2(n10629), .B1(n14262), .B2(n10628), .C1(
        n13874), .C2(P1_U3086), .ZN(P1_U3337) );
  INV_X1 U13176 ( .A(n10630), .ZN(n10633) );
  NAND4_X1 U13177 ( .A1(n10633), .A2(n10866), .A3(n10632), .A4(n10631), .ZN(
        n10859) );
  NAND2_X1 U13178 ( .A1(n10730), .A2(n12523), .ZN(n10634) );
  OAI21_X1 U13179 ( .B1(n15219), .B2(n10638), .A(n10634), .ZN(n10636) );
  NAND2_X1 U13180 ( .A1(n10636), .A2(n10635), .ZN(n10637) );
  NAND3_X1 U13181 ( .A1(n10637), .A2(n10861), .A3(n10640), .ZN(n10642) );
  AND2_X1 U13182 ( .A1(n10638), .A2(n12523), .ZN(n10639) );
  NAND2_X1 U13183 ( .A1(n10730), .A2(n10639), .ZN(n10940) );
  NAND2_X1 U13184 ( .A1(n10640), .A2(n10940), .ZN(n10860) );
  NAND2_X1 U13185 ( .A1(n10860), .A2(n10862), .ZN(n10641) );
  NAND2_X1 U13186 ( .A1(n15269), .A2(n15242), .ZN(n12884) );
  MUX2_X1 U13187 ( .A(n10868), .B(n10644), .S(n15270), .Z(n10645) );
  OAI21_X1 U13188 ( .B1(n10646), .B2(n12884), .A(n10645), .ZN(P3_U3459) );
  INV_X1 U13189 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10649) );
  MUX2_X1 U13190 ( .A(n10649), .B(P2_REG1_REG_14__SCAN_IN), .S(n11176), .Z(
        n10650) );
  NOR2_X1 U13191 ( .A1(n10651), .A2(n10650), .ZN(n11175) );
  AOI211_X1 U13192 ( .C1(n10651), .C2(n10650), .A(n11175), .B(n14803), .ZN(
        n10652) );
  INV_X1 U13193 ( .A(n10652), .ZN(n10664) );
  NAND2_X1 U13194 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n11730)
         );
  INV_X1 U13195 ( .A(n11730), .ZN(n10662) );
  OR2_X1 U13196 ( .A1(n10654), .A2(n10653), .ZN(n10655) );
  OAI21_X1 U13197 ( .B1(n10657), .B2(n10656), .A(n10655), .ZN(n11171) );
  INV_X1 U13198 ( .A(n11171), .ZN(n10658) );
  XNOR2_X1 U13199 ( .A(n11176), .B(n10658), .ZN(n10659) );
  NAND2_X1 U13200 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n10659), .ZN(n11172) );
  OAI211_X1 U13201 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n10659), .A(n14820), 
        .B(n11172), .ZN(n10660) );
  INV_X1 U13202 ( .A(n10660), .ZN(n10661) );
  AOI211_X1 U13203 ( .C1(P2_ADDR_REG_14__SCAN_IN), .C2(n14781), .A(n10662), 
        .B(n10661), .ZN(n10663) );
  OAI211_X1 U13204 ( .C1(n11524), .C2(n10665), .A(n10664), .B(n10663), .ZN(
        P2_U3228) );
  INV_X1 U13205 ( .A(n10681), .ZN(n10893) );
  NAND2_X1 U13206 ( .A1(n10682), .A2(n14903), .ZN(n10668) );
  INV_X1 U13207 ( .A(n13180), .ZN(n10686) );
  NAND2_X1 U13208 ( .A1(n10686), .A2(n10827), .ZN(n10669) );
  NAND2_X1 U13209 ( .A1(n10689), .A2(n14917), .ZN(n10670) );
  NOR2_X1 U13210 ( .A1(n13087), .A2(n13178), .ZN(n10672) );
  NAND2_X1 U13211 ( .A1(n13087), .A2(n13178), .ZN(n10673) );
  INV_X1 U13212 ( .A(n10694), .ZN(n10674) );
  OAI21_X1 U13213 ( .B1(n10675), .B2(n10674), .A(n10712), .ZN(n14836) );
  NAND2_X1 U13214 ( .A1(n10826), .A2(n10827), .ZN(n14851) );
  INV_X1 U13215 ( .A(n10817), .ZN(n10676) );
  INV_X1 U13216 ( .A(n14831), .ZN(n10708) );
  AOI211_X1 U13217 ( .C1(n14831), .C2(n10676), .A(n14849), .B(n10724), .ZN(
        n14826) );
  AND2_X1 U13218 ( .A1(n10216), .A2(n8919), .ZN(n10873) );
  NAND2_X1 U13219 ( .A1(n10874), .A2(n10873), .ZN(n10680) );
  INV_X1 U13220 ( .A(n13182), .ZN(n10678) );
  NAND2_X1 U13221 ( .A1(n10678), .A2(n10677), .ZN(n10679) );
  NAND2_X1 U13222 ( .A1(n10680), .A2(n10679), .ZN(n10894) );
  NAND2_X1 U13223 ( .A1(n10894), .A2(n10681), .ZN(n10684) );
  NAND2_X1 U13224 ( .A1(n10682), .A2(n10900), .ZN(n10683) );
  NAND2_X1 U13225 ( .A1(n10684), .A2(n10683), .ZN(n10830) );
  INV_X1 U13226 ( .A(n10685), .ZN(n10829) );
  NAND2_X1 U13227 ( .A1(n10830), .A2(n10829), .ZN(n10688) );
  NAND2_X1 U13228 ( .A1(n10686), .A2(n14909), .ZN(n10687) );
  INV_X1 U13229 ( .A(n14847), .ZN(n14839) );
  NAND2_X1 U13230 ( .A1(n14840), .A2(n14839), .ZN(n10691) );
  NAND2_X1 U13231 ( .A1(n10689), .A2(n14850), .ZN(n10690) );
  INV_X1 U13232 ( .A(n13178), .ZN(n10752) );
  AND2_X1 U13233 ( .A1(n10752), .A2(n13087), .ZN(n10692) );
  NAND2_X1 U13234 ( .A1(n7200), .A2(n13178), .ZN(n10693) );
  INV_X1 U13235 ( .A(n10813), .ZN(n10810) );
  INV_X1 U13236 ( .A(n13177), .ZN(n10698) );
  XNOR2_X1 U13237 ( .A(n10715), .B(n10694), .ZN(n10699) );
  OR2_X1 U13238 ( .A1(n9441), .A2(n13213), .ZN(n10697) );
  NAND2_X1 U13239 ( .A1(n9442), .A2(n10695), .ZN(n10696) );
  OAI22_X1 U13240 ( .A1(n10698), .A2(n13072), .B1(n10965), .B2(n13074), .ZN(
        n10855) );
  AOI21_X1 U13241 ( .B1(n10699), .B2(n14860), .A(n10855), .ZN(n14838) );
  INV_X1 U13242 ( .A(n14838), .ZN(n10700) );
  AOI211_X1 U13243 ( .C1(n14921), .C2(n14836), .A(n14826), .B(n10700), .ZN(
        n11412) );
  INV_X1 U13244 ( .A(n10701), .ZN(n10702) );
  OR3_X1 U13245 ( .A1(n10703), .A2(n10702), .A3(n14883), .ZN(n10770) );
  NAND2_X1 U13246 ( .A1(n14885), .A2(n10704), .ZN(n10705) );
  INV_X1 U13247 ( .A(n11337), .ZN(n10706) );
  NAND2_X1 U13248 ( .A1(n14942), .A2(n14933), .ZN(n13557) );
  INV_X1 U13249 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10707) );
  OAI22_X1 U13250 ( .A1(n13557), .A2(n10708), .B1(n14942), .B2(n10707), .ZN(
        n10709) );
  INV_X1 U13251 ( .A(n10709), .ZN(n10710) );
  OAI21_X1 U13252 ( .B1(n11412), .B2(n14940), .A(n10710), .ZN(P2_U3451) );
  OR2_X1 U13253 ( .A1(n14831), .A2(n13176), .ZN(n10711) );
  INV_X1 U13254 ( .A(n10713), .ZN(n10714) );
  OAI21_X1 U13255 ( .B1(n10714), .B2(n10718), .A(n10961), .ZN(n10786) );
  INV_X1 U13256 ( .A(n13176), .ZN(n10751) );
  OAI21_X1 U13257 ( .B1(n10715), .B2(n14831), .A(n10751), .ZN(n10717) );
  NAND2_X1 U13258 ( .A1(n10715), .A2(n14831), .ZN(n10716) );
  AOI21_X1 U13259 ( .B1(n10719), .B2(n10718), .A(n13368), .ZN(n10722) );
  NAND2_X1 U13260 ( .A1(n13144), .A2(n13174), .ZN(n10721) );
  NAND2_X1 U13261 ( .A1(n13176), .A2(n13142), .ZN(n10720) );
  NAND2_X1 U13262 ( .A1(n10721), .A2(n10720), .ZN(n11065) );
  AOI21_X1 U13263 ( .B1(n10722), .B2(n10967), .A(n11065), .ZN(n10777) );
  INV_X1 U13264 ( .A(n11060), .ZN(n11340) );
  OAI21_X1 U13265 ( .B1(n10724), .B2(n11340), .A(n13405), .ZN(n10725) );
  OR2_X1 U13266 ( .A1(n10962), .A2(n10725), .ZN(n10779) );
  OAI211_X1 U13267 ( .C1(n10786), .C2(n14938), .A(n10777), .B(n10779), .ZN(
        n11342) );
  INV_X1 U13268 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10726) );
  OAI22_X1 U13269 ( .A1(n13557), .A2(n11340), .B1(n14942), .B2(n10726), .ZN(
        n10727) );
  AOI21_X1 U13270 ( .B1(n11342), .B2(n14942), .A(n10727), .ZN(n10728) );
  INV_X1 U13271 ( .A(n10728), .ZN(P2_U3454) );
  INV_X1 U13272 ( .A(n10729), .ZN(n10732) );
  OAI22_X1 U13273 ( .A1(n10730), .A2(P3_U3151), .B1(SI_22_), .B2(n12966), .ZN(
        n10731) );
  AOI21_X1 U13274 ( .B1(n10732), .B2(n10884), .A(n10731), .ZN(P3_U3273) );
  INV_X1 U13275 ( .A(n10795), .ZN(n10743) );
  INV_X1 U13276 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10742) );
  NAND3_X1 U13277 ( .A1(n10733), .A2(n10936), .A3(n12328), .ZN(n10734) );
  OAI211_X1 U13278 ( .C1(n6599), .C2(n10927), .A(n10735), .B(n10734), .ZN(
        n10736) );
  NAND2_X1 U13279 ( .A1(n10736), .A2(n14960), .ZN(n10741) );
  NAND2_X1 U13280 ( .A1(n10737), .A2(n15145), .ZN(n10932) );
  INV_X1 U13281 ( .A(n14965), .ZN(n14425) );
  OAI22_X1 U13282 ( .A1(n10932), .A2(n14968), .B1(n14425), .B2(n10738), .ZN(
        n10739) );
  AOI21_X1 U13283 ( .B1(n12422), .B2(n6736), .A(n10739), .ZN(n10740) );
  OAI211_X1 U13284 ( .C1(n10743), .C2(n10742), .A(n10741), .B(n10740), .ZN(
        P3_U3162) );
  INV_X1 U13285 ( .A(n10744), .ZN(n10745) );
  AND2_X1 U13286 ( .A1(n13178), .A2(n14849), .ZN(n10748) );
  XNOR2_X1 U13287 ( .A(n6682), .B(n13087), .ZN(n10747) );
  NOR2_X1 U13288 ( .A1(n10747), .A2(n10748), .ZN(n10749) );
  AOI21_X1 U13289 ( .B1(n10748), .B2(n10747), .A(n10749), .ZN(n13083) );
  NAND2_X1 U13290 ( .A1(n13082), .A2(n13083), .ZN(n13081) );
  INV_X1 U13291 ( .A(n10749), .ZN(n10750) );
  XNOR2_X1 U13292 ( .A(n14934), .B(n6682), .ZN(n10848) );
  AND2_X1 U13293 ( .A1(n13177), .A2(n14849), .ZN(n10849) );
  XNOR2_X1 U13294 ( .A(n10848), .B(n10849), .ZN(n10852) );
  XNOR2_X1 U13295 ( .A(n10853), .B(n10852), .ZN(n10756) );
  OAI22_X1 U13296 ( .A1(n10752), .A2(n13072), .B1(n10751), .B2(n13074), .ZN(
        n10814) );
  AOI21_X1 U13297 ( .B1(n13097), .B2(n10814), .A(n10753), .ZN(n10755) );
  AOI22_X1 U13298 ( .A1(n13149), .A2(n14934), .B1(n10819), .B2(n13145), .ZN(
        n10754) );
  OAI211_X1 U13299 ( .C1(n10756), .C2(n13151), .A(n10755), .B(n10754), .ZN(
        P2_U3211) );
  INV_X1 U13300 ( .A(n11344), .ZN(n11717) );
  OAI22_X1 U13301 ( .A1(n11798), .A2(n11717), .B1(n12131), .B2(n14708), .ZN(
        n10757) );
  XOR2_X1 U13302 ( .A(n12132), .B(n10757), .Z(n10765) );
  OAI22_X1 U13303 ( .A1(n9620), .A2(n11798), .B1(n14708), .B2(n11717), .ZN(
        n10836) );
  INV_X1 U13304 ( .A(n10758), .ZN(n10761) );
  INV_X1 U13305 ( .A(n10759), .ZN(n10760) );
  AOI211_X1 U13306 ( .C1(n10765), .C2(n10764), .A(n13740), .B(n10837), .ZN(
        n10766) );
  INV_X1 U13307 ( .A(n10766), .ZN(n10769) );
  AOI22_X1 U13308 ( .A1(n13725), .A2(n13770), .B1(n13768), .B2(n6462), .ZN(
        n14662) );
  NAND2_X1 U13309 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n13814) );
  OAI21_X1 U13310 ( .B1(n13736), .B2(n14662), .A(n13814), .ZN(n10767) );
  AOI21_X1 U13311 ( .B1(n14676), .B2(n14554), .A(n10767), .ZN(n10768) );
  OAI211_X1 U13312 ( .C1(n14557), .C2(n14666), .A(n10769), .B(n10768), .ZN(
        P1_U3230) );
  INV_X1 U13313 ( .A(n10770), .ZN(n10772) );
  INV_X1 U13314 ( .A(n14885), .ZN(n10771) );
  NAND3_X1 U13315 ( .A1(n10772), .A2(n10771), .A3(n11337), .ZN(n10773) );
  NOR2_X1 U13316 ( .A1(n10774), .A2(n13213), .ZN(n10775) );
  NAND2_X1 U13317 ( .A1(n14871), .A2(n10775), .ZN(n14867) );
  INV_X1 U13318 ( .A(n14925), .ZN(n14861) );
  NAND2_X1 U13319 ( .A1(n14871), .A2(n14861), .ZN(n10776) );
  MUX2_X1 U13320 ( .A(n10778), .B(n10777), .S(n14871), .Z(n10785) );
  INV_X1 U13321 ( .A(n10779), .ZN(n10783) );
  INV_X1 U13322 ( .A(n10781), .ZN(n11068) );
  OAI22_X1 U13323 ( .A1(n13420), .A2(n11340), .B1(n14865), .B2(n11068), .ZN(
        n10782) );
  AOI21_X1 U13324 ( .B1(n14854), .B2(n10783), .A(n10782), .ZN(n10784) );
  OAI211_X1 U13325 ( .C1(n13425), .C2(n10786), .A(n10785), .B(n10784), .ZN(
        P2_U3257) );
  INV_X1 U13326 ( .A(n10787), .ZN(n10789) );
  OAI222_X1 U13327 ( .A1(n13599), .A2(n10788), .B1(n13587), .B2(n10789), .C1(
        P2_U3088), .C2(n13213), .ZN(P2_U3308) );
  OAI222_X1 U13328 ( .A1(n14258), .A2(n10790), .B1(n14262), .B2(n10789), .C1(
        n14564), .C2(P1_U3086), .ZN(P1_U3336) );
  XOR2_X1 U13329 ( .A(n10792), .B(n10791), .Z(n10797) );
  AOI22_X1 U13330 ( .A1(n12461), .A2(n12422), .B1(n14965), .B2(n15198), .ZN(
        n10793) );
  OAI21_X1 U13331 ( .B1(n15188), .B2(n12414), .A(n10793), .ZN(n10794) );
  AOI21_X1 U13332 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10795), .A(n10794), .ZN(
        n10796) );
  OAI21_X1 U13333 ( .B1(n10797), .B2(n12433), .A(n10796), .ZN(P3_U3177) );
  XNOR2_X1 U13334 ( .A(n10798), .B(n10802), .ZN(n14924) );
  OAI211_X1 U13335 ( .C1(n7201), .C2(n7200), .A(n13405), .B(n10818), .ZN(
        n14926) );
  INV_X1 U13336 ( .A(n14926), .ZN(n10801) );
  INV_X1 U13337 ( .A(n13086), .ZN(n10799) );
  OAI22_X1 U13338 ( .A1(n13420), .A2(n7200), .B1(n10799), .B2(n14865), .ZN(
        n10800) );
  AOI21_X1 U13339 ( .B1(n14854), .B2(n10801), .A(n10800), .ZN(n10809) );
  XNOR2_X1 U13340 ( .A(n10803), .B(n10802), .ZN(n10806) );
  NAND2_X1 U13341 ( .A1(n13144), .A2(n13177), .ZN(n10805) );
  NAND2_X1 U13342 ( .A1(n13179), .A2(n13142), .ZN(n10804) );
  NAND2_X1 U13343 ( .A1(n10805), .A2(n10804), .ZN(n13085) );
  AOI21_X1 U13344 ( .B1(n10806), .B2(n14860), .A(n13085), .ZN(n14927) );
  MUX2_X1 U13345 ( .A(n10807), .B(n14927), .S(n14871), .Z(n10808) );
  OAI211_X1 U13346 ( .C1(n13425), .C2(n14924), .A(n10809), .B(n10808), .ZN(
        P2_U3260) );
  XNOR2_X1 U13347 ( .A(n10811), .B(n10810), .ZN(n14937) );
  OAI21_X1 U13348 ( .B1(n6595), .B2(n10813), .A(n10812), .ZN(n10815) );
  AOI21_X1 U13349 ( .B1(n10815), .B2(n14860), .A(n10814), .ZN(n14936) );
  MUX2_X1 U13350 ( .A(n14936), .B(n10816), .S(n14873), .Z(n10824) );
  AOI211_X1 U13351 ( .C1(n14934), .C2(n10818), .A(n12981), .B(n10817), .ZN(
        n14932) );
  INV_X1 U13352 ( .A(n14934), .ZN(n10821) );
  INV_X1 U13353 ( .A(n10819), .ZN(n10820) );
  OAI22_X1 U13354 ( .A1(n13420), .A2(n10821), .B1(n10820), .B2(n14865), .ZN(
        n10822) );
  AOI21_X1 U13355 ( .B1(n14854), .B2(n14932), .A(n10822), .ZN(n10823) );
  OAI211_X1 U13356 ( .C1(n13425), .C2(n14937), .A(n10824), .B(n10823), .ZN(
        P2_U3259) );
  XNOR2_X1 U13357 ( .A(n10825), .B(n10829), .ZN(n14912) );
  INV_X1 U13358 ( .A(n10826), .ZN(n10890) );
  AOI211_X1 U13359 ( .C1(n14909), .C2(n10890), .A(n12981), .B(n7202), .ZN(
        n14908) );
  OAI22_X1 U13360 ( .A1(n13420), .A2(n10827), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14865), .ZN(n10828) );
  AOI21_X1 U13361 ( .B1(n14854), .B2(n14908), .A(n10828), .ZN(n10835) );
  XNOR2_X1 U13362 ( .A(n10830), .B(n10829), .ZN(n10832) );
  AOI21_X1 U13363 ( .B1(n10832), .B2(n14860), .A(n10831), .ZN(n14910) );
  MUX2_X1 U13364 ( .A(n10833), .B(n14910), .S(n14871), .Z(n10834) );
  OAI211_X1 U13365 ( .C1(n13425), .C2(n14912), .A(n10835), .B(n10834), .ZN(
        P2_U3262) );
  AOI22_X1 U13366 ( .A1(n11804), .A2(n12118), .B1(n12125), .B2(n13768), .ZN(
        n10838) );
  XNOR2_X1 U13367 ( .A(n10838), .B(n12132), .ZN(n11158) );
  AOI22_X1 U13368 ( .A1(n12068), .A2(n13768), .B1(n12125), .B2(n11804), .ZN(
        n11159) );
  XNOR2_X1 U13369 ( .A(n11158), .B(n7326), .ZN(n10839) );
  XNOR2_X1 U13370 ( .A(n6591), .B(n10839), .ZN(n10846) );
  NAND2_X1 U13371 ( .A1(n14554), .A2(n11804), .ZN(n10843) );
  AOI21_X1 U13372 ( .B1(n14552), .B2(n10841), .A(n10840), .ZN(n10842) );
  OAI211_X1 U13373 ( .C1(n14557), .C2(n10844), .A(n10843), .B(n10842), .ZN(
        n10845) );
  AOI21_X1 U13374 ( .B1(n10846), .B2(n14550), .A(n10845), .ZN(n10847) );
  INV_X1 U13375 ( .A(n10847), .ZN(P1_U3227) );
  INV_X1 U13376 ( .A(n10848), .ZN(n10851) );
  INV_X1 U13377 ( .A(n10849), .ZN(n10850) );
  XNOR2_X1 U13378 ( .A(n14831), .B(n6682), .ZN(n11056) );
  NAND2_X1 U13379 ( .A1(n13176), .A2(n14849), .ZN(n11055) );
  XNOR2_X1 U13380 ( .A(n11056), .B(n11055), .ZN(n11058) );
  XNOR2_X1 U13381 ( .A(n11059), .B(n11058), .ZN(n10858) );
  AOI21_X1 U13382 ( .B1(n13097), .B2(n10855), .A(n10854), .ZN(n10857) );
  AOI22_X1 U13383 ( .A1(n13149), .A2(n14831), .B1(n14827), .B2(n13145), .ZN(
        n10856) );
  OAI211_X1 U13384 ( .C1(n10858), .C2(n13151), .A(n10857), .B(n10856), .ZN(
        P2_U3185) );
  INV_X1 U13385 ( .A(n10859), .ZN(n10864) );
  MUX2_X1 U13386 ( .A(n10862), .B(n10861), .S(n10860), .Z(n10863) );
  NOR2_X1 U13387 ( .A1(n15219), .A2(n10946), .ZN(n10865) );
  MUX2_X1 U13388 ( .A(n10868), .B(n10867), .S(n15177), .Z(n10872) );
  AOI22_X1 U13389 ( .A1(n12695), .A2(n10870), .B1(n15203), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10871) );
  NAND2_X1 U13390 ( .A1(n10872), .A2(n10871), .ZN(P3_U3233) );
  XNOR2_X1 U13391 ( .A(n10874), .B(n12002), .ZN(n14893) );
  XNOR2_X1 U13392 ( .A(n10874), .B(n10873), .ZN(n10875) );
  NAND2_X1 U13393 ( .A1(n10875), .A2(n14860), .ZN(n10878) );
  INV_X1 U13394 ( .A(n10876), .ZN(n10877) );
  NAND2_X1 U13395 ( .A1(n10878), .A2(n10877), .ZN(n14896) );
  INV_X1 U13396 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10880) );
  INV_X1 U13397 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10879) );
  OAI22_X1 U13398 ( .A1(n14871), .A2(n10880), .B1(n10879), .B2(n14865), .ZN(
        n10882) );
  OAI211_X1 U13399 ( .C1(n14895), .C2(n14858), .A(n13405), .B(n10889), .ZN(
        n14894) );
  OAI22_X1 U13400 ( .A1(n14833), .A2(n14894), .B1(n14895), .B2(n13420), .ZN(
        n10881) );
  AOI211_X1 U13401 ( .C1(n14871), .C2(n14896), .A(n10882), .B(n10881), .ZN(
        n10883) );
  OAI21_X1 U13402 ( .B1(n13425), .B2(n14893), .A(n10883), .ZN(P2_U3264) );
  INV_X1 U13403 ( .A(SI_23_), .ZN(n10888) );
  NAND2_X1 U13404 ( .A1(n10885), .A2(n10884), .ZN(n10887) );
  OAI211_X1 U13405 ( .C1(n10888), .C2(n12966), .A(n10887), .B(n10886), .ZN(
        P3_U3272) );
  INV_X1 U13406 ( .A(n10889), .ZN(n10891) );
  OAI211_X1 U13407 ( .C1(n14903), .C2(n10891), .A(n10890), .B(n13405), .ZN(
        n14902) );
  XNOR2_X1 U13408 ( .A(n10892), .B(n10893), .ZN(n14900) );
  XNOR2_X1 U13409 ( .A(n10894), .B(n10893), .ZN(n10896) );
  OAI21_X1 U13410 ( .B1(n10896), .B2(n13368), .A(n10895), .ZN(n14905) );
  AOI22_X1 U13411 ( .A1(n14855), .A2(n14900), .B1(n14871), .B2(n14905), .ZN(
        n10902) );
  INV_X1 U13412 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10897) );
  OAI22_X1 U13413 ( .A1(n14871), .A2(n10898), .B1(n10897), .B2(n14865), .ZN(
        n10899) );
  AOI21_X1 U13414 ( .B1(n14846), .B2(n10900), .A(n10899), .ZN(n10901) );
  OAI211_X1 U13415 ( .C1(n14833), .C2(n14902), .A(n10902), .B(n10901), .ZN(
        P2_U3263) );
  INV_X1 U13416 ( .A(n10903), .ZN(n10904) );
  OAI21_X1 U13417 ( .B1(n10906), .B2(n10905), .A(n10904), .ZN(n10907) );
  NOR2_X1 U13418 ( .A1(n10918), .A2(n10907), .ZN(n10908) );
  XNOR2_X1 U13419 ( .A(n10918), .B(n10907), .ZN(n14626) );
  NOR2_X1 U13420 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14626), .ZN(n14625) );
  NOR2_X1 U13421 ( .A1(n10908), .A2(n14625), .ZN(n10911) );
  INV_X1 U13422 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11627) );
  NOR2_X1 U13423 ( .A1(n11628), .A2(n11627), .ZN(n10909) );
  AOI21_X1 U13424 ( .B1(n11627), .B2(n11628), .A(n10909), .ZN(n10910) );
  NAND2_X1 U13425 ( .A1(n10910), .A2(n10911), .ZN(n11626) );
  OAI211_X1 U13426 ( .C1(n10911), .C2(n10910), .A(n13879), .B(n11626), .ZN(
        n10926) );
  INV_X1 U13427 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10914) );
  NOR2_X1 U13428 ( .A1(n10912), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13657) );
  INV_X1 U13429 ( .A(n13657), .ZN(n10913) );
  OAI21_X1 U13430 ( .B1(n14640), .B2(n10914), .A(n10913), .ZN(n10924) );
  OR2_X1 U13431 ( .A1(n10915), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n10916) );
  XNOR2_X1 U13432 ( .A(n10919), .B(n14635), .ZN(n14630) );
  NAND2_X1 U13433 ( .A1(n14630), .A2(n7916), .ZN(n14629) );
  OAI21_X1 U13434 ( .B1(n10919), .B2(n10918), .A(n14629), .ZN(n10922) );
  INV_X1 U13435 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14576) );
  NOR2_X1 U13436 ( .A1(n11615), .A2(n14576), .ZN(n10920) );
  AOI21_X1 U13437 ( .B1(n11615), .B2(n14576), .A(n10920), .ZN(n10921) );
  NOR2_X1 U13438 ( .A1(n10921), .A2(n10922), .ZN(n11614) );
  AOI211_X1 U13439 ( .C1(n10922), .C2(n10921), .A(n11614), .B(n13860), .ZN(
        n10923) );
  AOI211_X1 U13440 ( .C1(n13855), .C2(n11615), .A(n10924), .B(n10923), .ZN(
        n10925) );
  NAND2_X1 U13441 ( .A1(n10926), .A2(n10925), .ZN(P1_U3259) );
  OAI21_X1 U13442 ( .B1(n10936), .B2(n10927), .A(n15179), .ZN(n10934) );
  INV_X1 U13443 ( .A(n10928), .ZN(n10930) );
  NAND2_X1 U13444 ( .A1(n6736), .A2(n15142), .ZN(n10931) );
  NAND2_X1 U13445 ( .A1(n10932), .A2(n10931), .ZN(n10933) );
  AOI21_X1 U13446 ( .B1(n10934), .B2(n15183), .A(n10933), .ZN(n10943) );
  XNOR2_X1 U13447 ( .A(n10936), .B(n10935), .ZN(n15207) );
  AND2_X1 U13448 ( .A1(n15219), .A2(n10937), .ZN(n10938) );
  NAND2_X1 U13449 ( .A1(n10939), .A2(n10938), .ZN(n10941) );
  OR2_X1 U13450 ( .A1(n15207), .A2(n15169), .ZN(n10942) );
  NAND2_X1 U13451 ( .A1(n10943), .A2(n10942), .ZN(n15208) );
  NAND2_X1 U13452 ( .A1(n10944), .A2(n15199), .ZN(n15200) );
  AND2_X1 U13453 ( .A1(n10945), .A2(n15242), .ZN(n15209) );
  AOI22_X1 U13454 ( .A1(n15209), .A2(n10946), .B1(n15203), .B2(
        P3_REG3_REG_1__SCAN_IN), .ZN(n10947) );
  OAI21_X1 U13455 ( .B1(n15207), .B2(n15200), .A(n10947), .ZN(n10948) );
  NOR2_X1 U13456 ( .A1(n15208), .A2(n10948), .ZN(n10950) );
  MUX2_X1 U13457 ( .A(n10950), .B(n10949), .S(n15177), .Z(n10951) );
  INV_X1 U13458 ( .A(n10951), .ZN(P3_U3232) );
  AOI21_X1 U13459 ( .B1(n10953), .B2(n10952), .A(n12433), .ZN(n10955) );
  NAND2_X1 U13460 ( .A1(n10955), .A2(n10954), .ZN(n10959) );
  OAI22_X1 U13461 ( .A1(n14425), .A2(n6719), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n8311), .ZN(n10957) );
  OAI22_X1 U13462 ( .A1(n12440), .A2(n15164), .B1(n11041), .B2(n12414), .ZN(
        n10956) );
  AOI211_X1 U13463 ( .C1(n8311), .C2(n14436), .A(n10957), .B(n10956), .ZN(
        n10958) );
  NAND2_X1 U13464 ( .A1(n10959), .A2(n10958), .ZN(P3_U3158) );
  NAND2_X1 U13465 ( .A1(n11060), .A2(n13175), .ZN(n10960) );
  INV_X1 U13466 ( .A(n11027), .ZN(n10968) );
  XNOR2_X1 U13467 ( .A(n11028), .B(n10968), .ZN(n11079) );
  INV_X1 U13468 ( .A(n10962), .ZN(n10964) );
  INV_X1 U13469 ( .A(n11413), .ZN(n11238) );
  INV_X1 U13470 ( .A(n11033), .ZN(n10963) );
  AOI211_X1 U13471 ( .C1(n11413), .C2(n10964), .A(n14849), .B(n10963), .ZN(
        n11073) );
  OR2_X1 U13472 ( .A1(n11060), .A2(n10965), .ZN(n10966) );
  OAI211_X1 U13473 ( .C1(n10969), .C2(n10968), .A(n11021), .B(n14860), .ZN(
        n10972) );
  NAND2_X1 U13474 ( .A1(n13144), .A2(n13173), .ZN(n10971) );
  NAND2_X1 U13475 ( .A1(n13175), .A2(n13142), .ZN(n10970) );
  AND2_X1 U13476 ( .A1(n10971), .A2(n10970), .ZN(n11232) );
  NAND2_X1 U13477 ( .A1(n10972), .A2(n11232), .ZN(n11076) );
  AOI211_X1 U13478 ( .C1(n14921), .C2(n11079), .A(n11073), .B(n11076), .ZN(
        n11415) );
  INV_X1 U13479 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10973) );
  OAI22_X1 U13480 ( .A1(n13557), .A2(n11238), .B1(n14942), .B2(n10973), .ZN(
        n10974) );
  INV_X1 U13481 ( .A(n10974), .ZN(n10975) );
  OAI21_X1 U13482 ( .B1(n11415), .B2(n14940), .A(n10975), .ZN(P2_U3457) );
  INV_X1 U13483 ( .A(n11964), .ZN(n10976) );
  XNOR2_X1 U13484 ( .A(n10977), .B(n10976), .ZN(n14740) );
  XNOR2_X1 U13485 ( .A(n10978), .B(n11964), .ZN(n10981) );
  NAND2_X1 U13486 ( .A1(n13725), .A2(n13765), .ZN(n10980) );
  NAND2_X1 U13487 ( .A1(n13763), .A2(n6462), .ZN(n10979) );
  NAND2_X1 U13488 ( .A1(n10980), .A2(n10979), .ZN(n11405) );
  AOI21_X1 U13489 ( .B1(n10981), .B2(n14664), .A(n11405), .ZN(n10982) );
  OAI21_X1 U13490 ( .B1(n14740), .B2(n14700), .A(n10982), .ZN(n14742) );
  NAND2_X1 U13491 ( .A1(n14742), .A2(n14389), .ZN(n10987) );
  OAI22_X1 U13492 ( .A1(n14389), .A2(n10983), .B1(n11407), .B2(n14667), .ZN(
        n10985) );
  OAI211_X1 U13493 ( .C1(n7107), .C2(n7106), .A(n14655), .B(n10995), .ZN(
        n14741) );
  NOR2_X1 U13494 ( .A1(n14741), .A2(n14090), .ZN(n10984) );
  AOI211_X1 U13495 ( .C1(n14398), .C2(n11829), .A(n10985), .B(n10984), .ZN(
        n10986) );
  OAI211_X1 U13496 ( .C1(n14740), .C2(n13988), .A(n10987), .B(n10986), .ZN(
        P1_U3284) );
  INV_X1 U13497 ( .A(n12259), .ZN(n10988) );
  NAND2_X1 U13498 ( .A1(n10988), .A2(P3_U3897), .ZN(n10989) );
  OAI21_X1 U13499 ( .B1(P3_U3897), .B2(n10990), .A(n10989), .ZN(P3_U3521) );
  XNOR2_X1 U13500 ( .A(n10991), .B(n11965), .ZN(n10993) );
  AND2_X1 U13501 ( .A1(n13725), .A2(n13764), .ZN(n11488) );
  INV_X1 U13502 ( .A(n11488), .ZN(n10992) );
  OAI21_X1 U13503 ( .B1(n10993), .B2(n14728), .A(n10992), .ZN(n14751) );
  INV_X1 U13504 ( .A(n14751), .ZN(n11005) );
  XNOR2_X1 U13505 ( .A(n10994), .B(n11965), .ZN(n14754) );
  NAND2_X1 U13506 ( .A1(n10995), .A2(n14747), .ZN(n10996) );
  NAND2_X1 U13507 ( .A1(n10996), .A2(n14655), .ZN(n10997) );
  OR2_X1 U13508 ( .A1(n10997), .A2(n11190), .ZN(n10999) );
  NAND2_X1 U13509 ( .A1(n13762), .A2(n6462), .ZN(n10998) );
  AND2_X1 U13510 ( .A1(n10999), .A2(n10998), .ZN(n14748) );
  OAI22_X1 U13511 ( .A1(n14389), .A2(n11000), .B1(n11491), .B2(n14667), .ZN(
        n11001) );
  AOI21_X1 U13512 ( .B1(n14398), .B2(n14747), .A(n11001), .ZN(n11002) );
  OAI21_X1 U13513 ( .B1(n14748), .B2(n14090), .A(n11002), .ZN(n11003) );
  AOI21_X1 U13514 ( .B1(n14754), .B2(n14677), .A(n11003), .ZN(n11004) );
  OAI21_X1 U13515 ( .B1(n11005), .B2(n6476), .A(n11004), .ZN(P1_U3283) );
  XNOR2_X1 U13516 ( .A(n6683), .B(n11963), .ZN(n14738) );
  OAI211_X1 U13517 ( .C1(n11008), .C2(n14735), .A(n11007), .B(n14655), .ZN(
        n14734) );
  INV_X1 U13518 ( .A(n14667), .ZN(n14680) );
  INV_X1 U13519 ( .A(n11009), .ZN(n11360) );
  AOI22_X1 U13520 ( .A1(n14398), .A2(n11820), .B1(n14680), .B2(n11360), .ZN(
        n11010) );
  OAI21_X1 U13521 ( .B1(n14090), .B2(n14734), .A(n11010), .ZN(n11017) );
  AOI21_X1 U13522 ( .B1(n11011), .B2(n11963), .A(n14728), .ZN(n11013) );
  NAND2_X1 U13523 ( .A1(n11013), .A2(n11012), .ZN(n11015) );
  AOI22_X1 U13524 ( .A1(n13725), .A2(n13766), .B1(n13764), .B2(n6462), .ZN(
        n11014) );
  NAND2_X1 U13525 ( .A1(n11015), .A2(n11014), .ZN(n14736) );
  MUX2_X1 U13526 ( .A(n14736), .B(P1_REG2_REG_8__SCAN_IN), .S(n6476), .Z(
        n11016) );
  AOI211_X1 U13527 ( .C1(n14677), .C2(n14738), .A(n11017), .B(n11016), .ZN(
        n11018) );
  INV_X1 U13528 ( .A(n11018), .ZN(P1_U3285) );
  OR2_X1 U13529 ( .A1(n11413), .A2(n11019), .ZN(n11020) );
  INV_X1 U13530 ( .A(n11250), .ZN(n11031) );
  OAI211_X1 U13531 ( .C1(n11022), .C2(n11031), .A(n11243), .B(n14860), .ZN(
        n11026) );
  NAND2_X1 U13532 ( .A1(n13144), .A2(n13172), .ZN(n11024) );
  NAND2_X1 U13533 ( .A1(n13174), .A2(n13142), .ZN(n11023) );
  NAND2_X1 U13534 ( .A1(n11024), .A2(n11023), .ZN(n11299) );
  INV_X1 U13535 ( .A(n11299), .ZN(n11025) );
  NAND2_X1 U13536 ( .A1(n11026), .A2(n11025), .ZN(n11081) );
  INV_X1 U13537 ( .A(n11081), .ZN(n11038) );
  NAND2_X1 U13538 ( .A1(n11413), .A2(n13174), .ZN(n11029) );
  NAND2_X1 U13539 ( .A1(n11030), .A2(n11029), .ZN(n11251) );
  XNOR2_X1 U13540 ( .A(n11251), .B(n11031), .ZN(n11083) );
  INV_X1 U13541 ( .A(n11254), .ZN(n11032) );
  AOI211_X1 U13542 ( .C1(n11445), .C2(n11033), .A(n14849), .B(n11032), .ZN(
        n11082) );
  NAND2_X1 U13543 ( .A1(n11082), .A2(n14854), .ZN(n11035) );
  INV_X1 U13544 ( .A(n14865), .ZN(n14844) );
  AOI22_X1 U13545 ( .A1(n14873), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11304), 
        .B2(n14844), .ZN(n11034) );
  OAI211_X1 U13546 ( .C1(n6664), .C2(n13420), .A(n11035), .B(n11034), .ZN(
        n11036) );
  AOI21_X1 U13547 ( .B1(n11083), .B2(n14855), .A(n11036), .ZN(n11037) );
  OAI21_X1 U13548 ( .B1(n11038), .B2(n14873), .A(n11037), .ZN(P2_U3255) );
  INV_X1 U13549 ( .A(n11046), .ZN(n11048) );
  XNOR2_X1 U13550 ( .A(n11039), .B(n11048), .ZN(n15218) );
  INV_X1 U13551 ( .A(n15200), .ZN(n15170) );
  NAND2_X1 U13552 ( .A1(n15204), .A2(n15170), .ZN(n12657) );
  AOI22_X1 U13553 ( .A1(n15145), .A2(n6736), .B1(n12460), .B2(n15142), .ZN(
        n11051) );
  NAND2_X1 U13554 ( .A1(n11041), .A2(n11040), .ZN(n11043) );
  AND2_X1 U13555 ( .A1(n15178), .A2(n11043), .ZN(n11042) );
  NAND2_X1 U13556 ( .A1(n15179), .A2(n11042), .ZN(n11045) );
  NAND2_X1 U13557 ( .A1(n11043), .A2(n15190), .ZN(n11044) );
  INV_X1 U13558 ( .A(n11047), .ZN(n11049) );
  OAI211_X1 U13559 ( .C1(n11049), .C2(n11048), .A(n15183), .B(n15155), .ZN(
        n11050) );
  OAI211_X1 U13560 ( .C1(n15218), .C2(n15169), .A(n11051), .B(n11050), .ZN(
        n15220) );
  NAND2_X1 U13561 ( .A1(n15220), .A2(n15204), .ZN(n11054) );
  OAI22_X1 U13562 ( .A1(n15204), .A2(n8313), .B1(n15104), .B2(
        P3_REG3_REG_3__SCAN_IN), .ZN(n11052) );
  AOI21_X1 U13563 ( .B1(n12695), .B2(n11327), .A(n11052), .ZN(n11053) );
  OAI211_X1 U13564 ( .C1(n15218), .C2(n12657), .A(n11054), .B(n11053), .ZN(
        P3_U3230) );
  INV_X1 U13565 ( .A(n11055), .ZN(n11057) );
  AND2_X1 U13566 ( .A1(n13175), .A2(n14849), .ZN(n11062) );
  XNOR2_X1 U13567 ( .A(n11060), .B(n6682), .ZN(n11061) );
  NOR2_X1 U13568 ( .A1(n11061), .A2(n11062), .ZN(n11226) );
  AOI21_X1 U13569 ( .B1(n11062), .B2(n11061), .A(n11226), .ZN(n11063) );
  NAND2_X1 U13570 ( .A1(n11064), .A2(n11063), .ZN(n11228) );
  OAI21_X1 U13571 ( .B1(n11064), .B2(n11063), .A(n11228), .ZN(n11071) );
  NOR2_X1 U13572 ( .A1(n13137), .A2(n11340), .ZN(n11070) );
  NAND2_X1 U13573 ( .A1(n13097), .A2(n11065), .ZN(n11067) );
  OAI211_X1 U13574 ( .C1(n13104), .C2(n11068), .A(n11067), .B(n11066), .ZN(
        n11069) );
  AOI211_X1 U13575 ( .C1(n11071), .C2(n13129), .A(n11070), .B(n11069), .ZN(
        n11072) );
  INV_X1 U13576 ( .A(n11072), .ZN(P2_U3193) );
  INV_X1 U13577 ( .A(n11073), .ZN(n11075) );
  AOI22_X1 U13578 ( .A1(n14846), .A2(n11413), .B1(n11235), .B2(n14844), .ZN(
        n11074) );
  OAI21_X1 U13579 ( .B1(n11075), .B2(n14833), .A(n11074), .ZN(n11078) );
  MUX2_X1 U13580 ( .A(n11076), .B(P2_REG2_REG_9__SCAN_IN), .S(n14873), .Z(
        n11077) );
  AOI211_X1 U13581 ( .C1(n14855), .C2(n11079), .A(n11078), .B(n11077), .ZN(
        n11080) );
  INV_X1 U13582 ( .A(n11080), .ZN(P2_U3256) );
  AOI211_X1 U13583 ( .C1(n14921), .C2(n11083), .A(n11082), .B(n11081), .ZN(
        n11447) );
  INV_X1 U13584 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11084) );
  OAI22_X1 U13585 ( .A1(n13557), .A2(n6664), .B1(n14942), .B2(n11084), .ZN(
        n11085) );
  INV_X1 U13586 ( .A(n11085), .ZN(n11086) );
  OAI21_X1 U13587 ( .B1(n11447), .B2(n14940), .A(n11086), .ZN(P2_U3460) );
  MUX2_X1 U13588 ( .A(n11118), .B(P3_REG2_REG_6__SCAN_IN), .S(n11120), .Z(
        n14992) );
  AOI22_X1 U13589 ( .A1(n15043), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n11131), 
        .B2(n11133), .ZN(n15038) );
  NAND2_X1 U13590 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n11202), .ZN(n11092) );
  OAI21_X1 U13591 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11202), .A(n11092), 
        .ZN(n11093) );
  AOI21_X1 U13592 ( .B1(n11094), .B2(n11093), .A(n11196), .ZN(n11157) );
  INV_X1 U13593 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15271) );
  AOI22_X1 U13594 ( .A1(n11144), .A2(n15271), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n11202), .ZN(n11104) );
  INV_X1 U13595 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15266) );
  AOI22_X1 U13596 ( .A1(n15043), .A2(n15266), .B1(P3_REG1_REG_8__SCAN_IN), 
        .B2(n11133), .ZN(n15042) );
  INV_X1 U13597 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15263) );
  NAND2_X1 U13598 ( .A1(n11115), .A2(n11096), .ZN(n11097) );
  NAND2_X1 U13599 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n14976), .ZN(n14975) );
  AND2_X1 U13600 ( .A1(n11097), .A2(n14975), .ZN(n14996) );
  MUX2_X1 U13601 ( .A(n15263), .B(P3_REG1_REG_6__SCAN_IN), .S(n11120), .Z(
        n14995) );
  INV_X1 U13602 ( .A(n14994), .ZN(n11098) );
  NAND2_X1 U13603 ( .A1(n15021), .A2(n11099), .ZN(n11100) );
  XNOR2_X1 U13604 ( .A(n11126), .B(n11099), .ZN(n15027) );
  NAND2_X1 U13605 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n15027), .ZN(n15026) );
  NAND2_X1 U13606 ( .A1(n11100), .A2(n15026), .ZN(n15041) );
  NAND2_X1 U13607 ( .A1(n15042), .A2(n15041), .ZN(n15040) );
  NAND2_X1 U13608 ( .A1(n11139), .A2(n11101), .ZN(n11102) );
  XNOR2_X1 U13609 ( .A(n15057), .B(n11101), .ZN(n15055) );
  NAND2_X1 U13610 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n15055), .ZN(n15054) );
  NAND2_X1 U13611 ( .A1(n11102), .A2(n15054), .ZN(n11103) );
  NAND2_X1 U13612 ( .A1(n11104), .A2(n11103), .ZN(n11203) );
  OAI21_X1 U13613 ( .B1(n11104), .B2(n11103), .A(n11203), .ZN(n11155) );
  INV_X1 U13614 ( .A(n15056), .ZN(n15020) );
  INV_X1 U13615 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11105) );
  NOR2_X1 U13616 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11105), .ZN(n11106) );
  AOI21_X1 U13617 ( .B1(n15025), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11106), 
        .ZN(n11107) );
  OAI21_X1 U13618 ( .B1(n15020), .B2(n11202), .A(n11107), .ZN(n11154) );
  NAND2_X1 U13619 ( .A1(n11109), .A2(n11108), .ZN(n11114) );
  INV_X1 U13620 ( .A(n11110), .ZN(n11112) );
  NAND2_X1 U13621 ( .A1(n11112), .A2(n11111), .ZN(n11113) );
  NAND2_X1 U13622 ( .A1(n11114), .A2(n11113), .ZN(n14980) );
  MUX2_X1 U13623 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12516), .Z(n11116) );
  NAND2_X1 U13624 ( .A1(n11116), .A2(n11115), .ZN(n14981) );
  NAND2_X1 U13625 ( .A1(n14980), .A2(n14981), .ZN(n15003) );
  INV_X1 U13626 ( .A(n11116), .ZN(n11117) );
  NAND2_X1 U13627 ( .A1(n11117), .A2(n14987), .ZN(n15002) );
  NAND2_X1 U13628 ( .A1(n15003), .A2(n15002), .ZN(n11123) );
  MUX2_X1 U13629 ( .A(n11118), .B(n15263), .S(n12516), .Z(n11119) );
  NAND2_X1 U13630 ( .A1(n11119), .A2(n15007), .ZN(n15014) );
  INV_X1 U13631 ( .A(n11119), .ZN(n11121) );
  NAND2_X1 U13632 ( .A1(n11121), .A2(n11120), .ZN(n11122) );
  AND2_X1 U13633 ( .A1(n15014), .A2(n11122), .ZN(n15000) );
  NAND2_X1 U13634 ( .A1(n11123), .A2(n15000), .ZN(n15018) );
  NAND2_X1 U13635 ( .A1(n15018), .A2(n15014), .ZN(n11130) );
  INV_X1 U13636 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11124) );
  MUX2_X1 U13637 ( .A(n11125), .B(n11124), .S(n12516), .Z(n11127) );
  NAND2_X1 U13638 ( .A1(n11127), .A2(n11126), .ZN(n15034) );
  INV_X1 U13639 ( .A(n11127), .ZN(n11128) );
  NAND2_X1 U13640 ( .A1(n11128), .A2(n15021), .ZN(n11129) );
  AND2_X1 U13641 ( .A1(n15034), .A2(n11129), .ZN(n15016) );
  NAND2_X1 U13642 ( .A1(n11130), .A2(n15016), .ZN(n15035) );
  NAND2_X1 U13643 ( .A1(n15035), .A2(n15034), .ZN(n11136) );
  MUX2_X1 U13644 ( .A(n11131), .B(n15266), .S(n12516), .Z(n11132) );
  NAND2_X1 U13645 ( .A1(n11132), .A2(n15043), .ZN(n15065) );
  INV_X1 U13646 ( .A(n11132), .ZN(n11134) );
  NAND2_X1 U13647 ( .A1(n11134), .A2(n11133), .ZN(n11135) );
  AND2_X1 U13648 ( .A1(n15065), .A2(n11135), .ZN(n15032) );
  NAND2_X1 U13649 ( .A1(n11136), .A2(n15032), .ZN(n15066) );
  NAND2_X1 U13650 ( .A1(n15066), .A2(n15065), .ZN(n11142) );
  INV_X1 U13651 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11137) );
  MUX2_X1 U13652 ( .A(n15098), .B(n11137), .S(n12516), .Z(n11138) );
  NAND2_X1 U13653 ( .A1(n11138), .A2(n15057), .ZN(n11151) );
  INV_X1 U13654 ( .A(n11138), .ZN(n11140) );
  NAND2_X1 U13655 ( .A1(n11140), .A2(n11139), .ZN(n11141) );
  AND2_X1 U13656 ( .A1(n11151), .A2(n11141), .ZN(n15063) );
  NAND2_X1 U13657 ( .A1(n11142), .A2(n15063), .ZN(n15069) );
  NAND2_X1 U13658 ( .A1(n15069), .A2(n11151), .ZN(n11148) );
  MUX2_X1 U13659 ( .A(n11143), .B(n15271), .S(n12516), .Z(n11145) );
  NAND2_X1 U13660 ( .A1(n11145), .A2(n11144), .ZN(n11198) );
  INV_X1 U13661 ( .A(n11145), .ZN(n11146) );
  NAND2_X1 U13662 ( .A1(n11146), .A2(n11202), .ZN(n11147) );
  AND2_X1 U13663 ( .A1(n11198), .A2(n11147), .ZN(n11149) );
  NAND2_X1 U13664 ( .A1(n11148), .A2(n11149), .ZN(n11199) );
  INV_X1 U13665 ( .A(n11149), .ZN(n11150) );
  NAND3_X1 U13666 ( .A1(n15069), .A2(n11151), .A3(n11150), .ZN(n11152) );
  AOI21_X1 U13667 ( .B1(n11199), .B2(n11152), .A(n15067), .ZN(n11153) );
  AOI211_X1 U13668 ( .C1(n15058), .C2(n11155), .A(n11154), .B(n11153), .ZN(
        n11156) );
  OAI21_X1 U13669 ( .B1(n11157), .B2(n15061), .A(n11156), .ZN(P3_U3192) );
  AOI22_X1 U13670 ( .A1(n14648), .A2(n12125), .B1(n12068), .B2(n13767), .ZN(
        n11266) );
  NAND2_X1 U13671 ( .A1(n14648), .A2(n12118), .ZN(n11161) );
  NAND2_X1 U13672 ( .A1(n12125), .A2(n13767), .ZN(n11160) );
  NAND2_X1 U13673 ( .A1(n11161), .A2(n11160), .ZN(n11162) );
  XNOR2_X1 U13674 ( .A(n11162), .B(n12132), .ZN(n11265) );
  XOR2_X1 U13675 ( .A(n11266), .B(n11265), .Z(n11267) );
  XOR2_X1 U13676 ( .A(n11268), .B(n11267), .Z(n11169) );
  NAND2_X1 U13677 ( .A1(n14554), .A2(n14648), .ZN(n11167) );
  NAND2_X1 U13678 ( .A1(n13725), .A2(n13768), .ZN(n11164) );
  NAND2_X1 U13679 ( .A1(n13766), .A2(n6462), .ZN(n11163) );
  NAND2_X1 U13680 ( .A1(n11164), .A2(n11163), .ZN(n14647) );
  AOI21_X1 U13681 ( .B1(n14552), .B2(n14647), .A(n11165), .ZN(n11166) );
  OAI211_X1 U13682 ( .C1(n14557), .C2(n14649), .A(n11167), .B(n11166), .ZN(
        n11168) );
  AOI21_X1 U13683 ( .B1(n11169), .B2(n14550), .A(n11168), .ZN(n11170) );
  INV_X1 U13684 ( .A(n11170), .ZN(P1_U3239) );
  NAND2_X1 U13685 ( .A1(n11176), .A2(n11171), .ZN(n11173) );
  NAND2_X1 U13686 ( .A1(n11173), .A2(n11172), .ZN(n11284) );
  XNOR2_X1 U13687 ( .A(n11284), .B(n11278), .ZN(n11174) );
  NAND2_X1 U13688 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n11174), .ZN(n11286) );
  OAI211_X1 U13689 ( .C1(n11174), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14820), 
        .B(n11286), .ZN(n11182) );
  AND2_X1 U13690 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n11180) );
  XNOR2_X1 U13691 ( .A(n11278), .B(n11279), .ZN(n11178) );
  NOR2_X1 U13692 ( .A1(n11177), .A2(n11178), .ZN(n11280) );
  AOI211_X1 U13693 ( .C1(n11178), .C2(n11177), .A(n11280), .B(n14803), .ZN(
        n11179) );
  AOI211_X1 U13694 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n14781), .A(n11180), 
        .B(n11179), .ZN(n11181) );
  OAI211_X1 U13695 ( .C1(n11524), .C2(n11278), .A(n11182), .B(n11181), .ZN(
        P2_U3229) );
  XNOR2_X1 U13696 ( .A(n11183), .B(n11966), .ZN(n11187) );
  OR2_X1 U13697 ( .A1(n11841), .A2(n13713), .ZN(n11185) );
  NAND2_X1 U13698 ( .A1(n13725), .A2(n13763), .ZN(n11184) );
  NAND2_X1 U13699 ( .A1(n11185), .A2(n11184), .ZN(n11656) );
  INV_X1 U13700 ( .A(n11656), .ZN(n11186) );
  OAI21_X1 U13701 ( .B1(n11187), .B2(n14728), .A(n11186), .ZN(n14594) );
  INV_X1 U13702 ( .A(n14594), .ZN(n11195) );
  XNOR2_X1 U13703 ( .A(n11188), .B(n7116), .ZN(n14596) );
  INV_X1 U13704 ( .A(n14402), .ZN(n11189) );
  OAI211_X1 U13705 ( .C1(n14593), .C2(n11190), .A(n11189), .B(n14655), .ZN(
        n14592) );
  OAI22_X1 U13706 ( .A1(n14389), .A2(n9896), .B1(n11653), .B2(n14667), .ZN(
        n11191) );
  AOI21_X1 U13707 ( .B1(n14398), .B2(n11837), .A(n11191), .ZN(n11192) );
  OAI21_X1 U13708 ( .B1(n14592), .B2(n14090), .A(n11192), .ZN(n11193) );
  AOI21_X1 U13709 ( .B1(n14596), .B2(n14677), .A(n11193), .ZN(n11194) );
  OAI21_X1 U13710 ( .B1(n11195), .B2(n6476), .A(n11194), .ZN(P1_U3282) );
  NOR2_X1 U13711 ( .A1(n8438), .A2(n11197), .ZN(n11417) );
  AOI21_X1 U13712 ( .B1(n8438), .B2(n11197), .A(n11417), .ZN(n11213) );
  NAND2_X1 U13713 ( .A1(n11199), .A2(n11198), .ZN(n11201) );
  MUX2_X1 U13714 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12516), .Z(n11429) );
  INV_X1 U13715 ( .A(n11422), .ZN(n11430) );
  XNOR2_X1 U13716 ( .A(n11429), .B(n11430), .ZN(n11200) );
  NAND2_X1 U13717 ( .A1(n11201), .A2(n11200), .ZN(n11435) );
  OAI21_X1 U13718 ( .B1(n11201), .B2(n11200), .A(n11435), .ZN(n11211) );
  INV_X1 U13719 ( .A(n15067), .ZN(n14478) );
  NAND2_X1 U13720 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11202), .ZN(n11204) );
  NAND2_X1 U13721 ( .A1(n11204), .A2(n11203), .ZN(n11421) );
  XNOR2_X1 U13722 ( .A(n11430), .B(n11421), .ZN(n11205) );
  NAND2_X1 U13723 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n11205), .ZN(n11423) );
  OAI21_X1 U13724 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n11205), .A(n11423), 
        .ZN(n11206) );
  NAND2_X1 U13725 ( .A1(n11206), .A2(n15058), .ZN(n11209) );
  AOI21_X1 U13726 ( .B1(n15025), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11207), 
        .ZN(n11208) );
  OAI211_X1 U13727 ( .C1(n15020), .C2(n11422), .A(n11209), .B(n11208), .ZN(
        n11210) );
  AOI21_X1 U13728 ( .B1(n11211), .B2(n14478), .A(n11210), .ZN(n11212) );
  OAI21_X1 U13729 ( .B1(n11213), .B2(n15061), .A(n11212), .ZN(P3_U3193) );
  INV_X1 U13730 ( .A(n11214), .ZN(n11239) );
  OAI222_X1 U13731 ( .A1(n13599), .A2(n7009), .B1(n13587), .B2(n11239), .C1(
        n8923), .C2(P2_U3088), .ZN(P2_U3307) );
  INV_X1 U13732 ( .A(n11333), .ZN(n11223) );
  OAI21_X1 U13733 ( .B1(n11217), .B2(n11216), .A(n11215), .ZN(n11218) );
  NAND2_X1 U13734 ( .A1(n11218), .A2(n14960), .ZN(n11222) );
  OAI22_X1 U13735 ( .A1(n12440), .A2(n12212), .B1(n15186), .B2(n12414), .ZN(
        n11219) );
  AOI211_X1 U13736 ( .C1(n14965), .C2(n15223), .A(n11220), .B(n11219), .ZN(
        n11221) );
  OAI211_X1 U13737 ( .C1(n11223), .C2(n14971), .A(n11222), .B(n11221), .ZN(
        P3_U3170) );
  AND2_X1 U13738 ( .A1(n13174), .A2(n14849), .ZN(n11225) );
  XNOR2_X1 U13739 ( .A(n11413), .B(n6682), .ZN(n11224) );
  NOR2_X1 U13740 ( .A1(n11224), .A2(n11225), .ZN(n11296) );
  AOI21_X1 U13741 ( .B1(n11225), .B2(n11224), .A(n11296), .ZN(n11230) );
  INV_X1 U13742 ( .A(n11226), .ZN(n11227) );
  OAI21_X1 U13743 ( .B1(n11230), .B2(n6684), .A(n11298), .ZN(n11231) );
  NAND2_X1 U13744 ( .A1(n11231), .A2(n13129), .ZN(n11237) );
  NOR2_X1 U13745 ( .A1(n13147), .A2(n11232), .ZN(n11233) );
  AOI211_X1 U13746 ( .C1(n13145), .C2(n11235), .A(n11234), .B(n11233), .ZN(
        n11236) );
  OAI211_X1 U13747 ( .C1(n11238), .C2(n13137), .A(n11237), .B(n11236), .ZN(
        P2_U3203) );
  OAI222_X1 U13748 ( .A1(n11694), .A2(n11240), .B1(P1_U3086), .B2(n11938), 
        .C1(n14262), .C2(n11239), .ZN(P1_U3335) );
  OR2_X1 U13749 ( .A1(n11445), .A2(n11241), .ZN(n11242) );
  INV_X1 U13750 ( .A(n11450), .ZN(n11244) );
  AOI21_X1 U13751 ( .B1(n11455), .B2(n11245), .A(n11244), .ZN(n11249) );
  NAND2_X1 U13752 ( .A1(n13144), .A2(n13171), .ZN(n11247) );
  NAND2_X1 U13753 ( .A1(n13173), .A2(n13142), .ZN(n11246) );
  NAND2_X1 U13754 ( .A1(n11247), .A2(n11246), .ZN(n11377) );
  INV_X1 U13755 ( .A(n11377), .ZN(n11248) );
  OAI21_X1 U13756 ( .B1(n11249), .B2(n13368), .A(n11248), .ZN(n11384) );
  INV_X1 U13757 ( .A(n11384), .ZN(n11260) );
  NAND2_X1 U13758 ( .A1(n11251), .A2(n11250), .ZN(n11253) );
  NAND2_X1 U13759 ( .A1(n11445), .A2(n13173), .ZN(n11252) );
  XNOR2_X1 U13760 ( .A(n11456), .B(n6825), .ZN(n11386) );
  INV_X1 U13761 ( .A(n11457), .ZN(n11257) );
  AOI211_X1 U13762 ( .C1(n11457), .C2(n6465), .A(n14849), .B(n14527), .ZN(
        n11385) );
  NAND2_X1 U13763 ( .A1(n11385), .A2(n14854), .ZN(n11256) );
  AOI22_X1 U13764 ( .A1(n14873), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11376), 
        .B2(n14844), .ZN(n11255) );
  OAI211_X1 U13765 ( .C1(n11257), .C2(n13420), .A(n11256), .B(n11255), .ZN(
        n11258) );
  AOI21_X1 U13766 ( .B1(n11386), .B2(n14855), .A(n11258), .ZN(n11259) );
  OAI21_X1 U13767 ( .B1(n11260), .B2(n14873), .A(n11259), .ZN(P2_U3254) );
  INV_X1 U13768 ( .A(n11261), .ZN(n11263) );
  INV_X1 U13769 ( .A(SI_24_), .ZN(n11262) );
  OAI222_X1 U13770 ( .A1(n11264), .A2(P3_U3151), .B1(n6461), .B2(n11263), .C1(
        n11262), .C2(n12966), .ZN(P3_U3271) );
  NOR2_X1 U13771 ( .A1(n9620), .A2(n11269), .ZN(n11270) );
  AOI21_X1 U13772 ( .B1(n14725), .B2(n12125), .A(n11270), .ZN(n11347) );
  AOI22_X1 U13773 ( .A1(n14725), .A2(n12118), .B1(n12125), .B2(n13766), .ZN(
        n11271) );
  XNOR2_X1 U13774 ( .A(n11271), .B(n12132), .ZN(n11348) );
  XOR2_X1 U13775 ( .A(n11347), .B(n11348), .Z(n11351) );
  XOR2_X1 U13776 ( .A(n11352), .B(n11351), .Z(n11276) );
  NAND2_X1 U13777 ( .A1(n14554), .A2(n14725), .ZN(n11273) );
  AND2_X1 U13778 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n13832) );
  AOI21_X1 U13779 ( .B1(n14552), .B2(n14723), .A(n13832), .ZN(n11272) );
  OAI211_X1 U13780 ( .C1(n14557), .C2(n11274), .A(n11273), .B(n11272), .ZN(
        n11275) );
  AOI21_X1 U13781 ( .B1(n11276), .B2(n14550), .A(n11275), .ZN(n11277) );
  INV_X1 U13782 ( .A(n11277), .ZN(P1_U3213) );
  NOR2_X1 U13783 ( .A1(n11279), .A2(n11278), .ZN(n11281) );
  XNOR2_X1 U13784 ( .A(n11508), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n11282) );
  NOR2_X1 U13785 ( .A1(n11283), .A2(n11282), .ZN(n11507) );
  AOI211_X1 U13786 ( .C1(n11283), .C2(n11282), .A(n11507), .B(n14803), .ZN(
        n11295) );
  NAND2_X1 U13787 ( .A1(n11285), .A2(n11284), .ZN(n11287) );
  NAND2_X1 U13788 ( .A1(n11287), .A2(n11286), .ZN(n11290) );
  NOR2_X1 U13789 ( .A1(n11508), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11288) );
  AOI21_X1 U13790 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n11508), .A(n11288), 
        .ZN(n11289) );
  NAND2_X1 U13791 ( .A1(n11289), .A2(n11290), .ZN(n11513) );
  OAI211_X1 U13792 ( .C1(n11290), .C2(n11289), .A(n14820), .B(n11513), .ZN(
        n11293) );
  NOR2_X1 U13793 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13076), .ZN(n11291) );
  AOI21_X1 U13794 ( .B1(n14781), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n11291), 
        .ZN(n11292) );
  OAI211_X1 U13795 ( .C1(n11524), .C2(n11515), .A(n11293), .B(n11292), .ZN(
        n11294) );
  OR2_X1 U13796 ( .A1(n11295), .A2(n11294), .ZN(P2_U3230) );
  INV_X1 U13797 ( .A(n11296), .ZN(n11297) );
  NAND2_X1 U13798 ( .A1(n13173), .A2(n12981), .ZN(n11370) );
  XOR2_X1 U13799 ( .A(n11370), .B(n11369), .Z(n11371) );
  XNOR2_X1 U13800 ( .A(n11372), .B(n11371), .ZN(n11306) );
  NAND2_X1 U13801 ( .A1(n13097), .A2(n11299), .ZN(n11300) );
  OAI21_X1 U13802 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n11301), .A(n11300), .ZN(
        n11303) );
  NOR2_X1 U13803 ( .A1(n13137), .A2(n6664), .ZN(n11302) );
  AOI211_X1 U13804 ( .C1(n13145), .C2(n11304), .A(n11303), .B(n11302), .ZN(
        n11305) );
  OAI21_X1 U13805 ( .B1(n11306), .B2(n13151), .A(n11305), .ZN(P2_U3189) );
  XOR2_X1 U13806 ( .A(n11308), .B(n11307), .Z(n11313) );
  OAI22_X1 U13807 ( .A1(n14425), .A2(n12211), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11309), .ZN(n11311) );
  OAI22_X1 U13808 ( .A1(n12440), .A2(n15163), .B1(n15164), .B2(n12414), .ZN(
        n11310) );
  AOI211_X1 U13809 ( .C1(n15172), .C2(n14436), .A(n11311), .B(n11310), .ZN(
        n11312) );
  OAI21_X1 U13810 ( .B1(n11313), .B2(n12433), .A(n11312), .ZN(P3_U3167) );
  XNOR2_X1 U13811 ( .A(n11315), .B(n11314), .ZN(n14589) );
  XNOR2_X1 U13812 ( .A(n11316), .B(n11970), .ZN(n14591) );
  NAND2_X1 U13813 ( .A1(n14591), .A2(n14055), .ZN(n11325) );
  OR2_X1 U13814 ( .A1(n12016), .A2(n13713), .ZN(n11318) );
  OR2_X1 U13815 ( .A1(n11841), .A2(n13711), .ZN(n11317) );
  NAND2_X1 U13816 ( .A1(n11318), .A2(n11317), .ZN(n14584) );
  INV_X1 U13817 ( .A(n11721), .ZN(n11319) );
  AOI22_X1 U13818 ( .A1(n14389), .A2(n14584), .B1(n11319), .B2(n14680), .ZN(
        n11320) );
  OAI21_X1 U13819 ( .B1(n11321), .B2(n14389), .A(n11320), .ZN(n11323) );
  OAI211_X1 U13820 ( .C1(n14400), .C2(n11839), .A(n14655), .B(n11573), .ZN(
        n14586) );
  NOR2_X1 U13821 ( .A1(n14586), .A2(n14090), .ZN(n11322) );
  AOI211_X1 U13822 ( .C1(n14398), .C2(n14585), .A(n11323), .B(n11322), .ZN(
        n11324) );
  OAI211_X1 U13823 ( .C1(n14589), .C2(n14077), .A(n11325), .B(n11324), .ZN(
        P1_U3280) );
  INV_X1 U13824 ( .A(n15224), .ZN(n11336) );
  INV_X1 U13825 ( .A(n15169), .ZN(n15194) );
  OAI22_X1 U13826 ( .A1(n15186), .A2(n15187), .B1(n12212), .B2(n15185), .ZN(
        n11331) );
  NAND2_X1 U13827 ( .A1(n12461), .A2(n11327), .ZN(n12216) );
  NAND2_X1 U13828 ( .A1(n15155), .A2(n12216), .ZN(n11328) );
  XNOR2_X1 U13829 ( .A(n11328), .B(n12213), .ZN(n11329) );
  NOR2_X1 U13830 ( .A1(n11329), .A2(n15130), .ZN(n11330) );
  AOI211_X1 U13831 ( .C1(n15194), .C2(n15224), .A(n11331), .B(n11330), .ZN(
        n15226) );
  MUX2_X1 U13832 ( .A(n11332), .B(n15226), .S(n15204), .Z(n11335) );
  AOI22_X1 U13833 ( .A1(n12695), .A2(n15223), .B1(n15203), .B2(n11333), .ZN(
        n11334) );
  OAI211_X1 U13834 ( .C1(n11336), .C2(n12657), .A(n11335), .B(n11334), .ZN(
        P3_U3229) );
  OAI22_X1 U13835 ( .A1(n13486), .A2(n11340), .B1(n14535), .B2(n11339), .ZN(
        n11341) );
  AOI21_X1 U13836 ( .B1(n11342), .B2(n14535), .A(n11341), .ZN(n11343) );
  INV_X1 U13837 ( .A(n11343), .ZN(P2_U3507) );
  OAI22_X1 U13838 ( .A1(n14735), .A2(n11717), .B1(n11345), .B2(n9615), .ZN(
        n11393) );
  OAI22_X1 U13839 ( .A1(n14735), .A2(n12131), .B1(n11345), .B2(n11717), .ZN(
        n11346) );
  XNOR2_X1 U13840 ( .A(n11346), .B(n12132), .ZN(n11392) );
  XOR2_X1 U13841 ( .A(n11393), .B(n11392), .Z(n11354) );
  INV_X1 U13842 ( .A(n11347), .ZN(n11350) );
  INV_X1 U13843 ( .A(n11348), .ZN(n11349) );
  OAI21_X1 U13844 ( .B1(n11354), .B2(n11353), .A(n11401), .ZN(n11355) );
  NAND2_X1 U13845 ( .A1(n11355), .A2(n14550), .ZN(n11362) );
  AOI21_X1 U13846 ( .B1(n11357), .B2(n13766), .A(n11356), .ZN(n11358) );
  OAI21_X1 U13847 ( .B1(n11398), .B2(n11490), .A(n11358), .ZN(n11359) );
  AOI21_X1 U13848 ( .B1(n11360), .B2(n13734), .A(n11359), .ZN(n11361) );
  OAI211_X1 U13849 ( .C1(n14735), .C2(n13730), .A(n11362), .B(n11361), .ZN(
        P1_U3221) );
  INV_X1 U13850 ( .A(n11363), .ZN(n11390) );
  OAI222_X1 U13851 ( .A1(n13599), .A2(n11365), .B1(n13587), .B2(n11390), .C1(
        n6618), .C2(P2_U3088), .ZN(P2_U3306) );
  INV_X1 U13852 ( .A(n11366), .ZN(n11367) );
  OAI222_X1 U13853 ( .A1(P3_U3151), .A2(n11368), .B1(n6460), .B2(n11367), .C1(
        n7451), .C2(n12966), .ZN(P3_U3270) );
  INV_X1 U13854 ( .A(n6682), .ZN(n13006) );
  XNOR2_X1 U13855 ( .A(n11457), .B(n13006), .ZN(n11374) );
  NAND2_X1 U13856 ( .A1(n13172), .A2(n12981), .ZN(n11373) );
  NOR2_X1 U13857 ( .A1(n11374), .A2(n11373), .ZN(n11525) );
  NOR2_X1 U13858 ( .A1(n11525), .A2(n6593), .ZN(n11375) );
  XNOR2_X1 U13859 ( .A(n11526), .B(n11375), .ZN(n11383) );
  NAND2_X1 U13860 ( .A1(n13145), .A2(n11376), .ZN(n11379) );
  NAND2_X1 U13861 ( .A1(n13097), .A2(n11377), .ZN(n11378) );
  OAI211_X1 U13862 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n11380), .A(n11379), .B(
        n11378), .ZN(n11381) );
  AOI21_X1 U13863 ( .B1(n11457), .B2(n13149), .A(n11381), .ZN(n11382) );
  OAI21_X1 U13864 ( .B1(n11383), .B2(n13151), .A(n11382), .ZN(P2_U3208) );
  AOI211_X1 U13865 ( .C1(n14921), .C2(n11386), .A(n11385), .B(n11384), .ZN(
        n11444) );
  INV_X1 U13866 ( .A(n13557), .ZN(n13563) );
  INV_X1 U13867 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11387) );
  NOR2_X1 U13868 ( .A1(n14942), .A2(n11387), .ZN(n11388) );
  AOI21_X1 U13869 ( .B1(n13563), .B2(n11457), .A(n11388), .ZN(n11389) );
  OAI21_X1 U13870 ( .B1(n11444), .B2(n14940), .A(n11389), .ZN(P2_U3463) );
  OAI222_X1 U13871 ( .A1(n11694), .A2(n11391), .B1(P1_U3086), .B2(n11756), 
        .C1(n14262), .C2(n11390), .ZN(P1_U3334) );
  INV_X1 U13872 ( .A(n11392), .ZN(n11395) );
  INV_X1 U13873 ( .A(n11393), .ZN(n11394) );
  NAND2_X1 U13874 ( .A1(n11395), .A2(n11394), .ZN(n11400) );
  AND2_X1 U13875 ( .A1(n11401), .A2(n11400), .ZN(n11403) );
  OAI22_X1 U13876 ( .A1(n7106), .A2(n12131), .B1(n11398), .B2(n11396), .ZN(
        n11397) );
  XNOR2_X1 U13877 ( .A(n11397), .B(n12132), .ZN(n11480) );
  NOR2_X1 U13878 ( .A1(n9615), .A2(n11398), .ZN(n11399) );
  AOI21_X1 U13879 ( .B1(n11829), .B2(n12125), .A(n11399), .ZN(n11483) );
  XNOR2_X1 U13880 ( .A(n11480), .B(n11483), .ZN(n11402) );
  NAND3_X1 U13881 ( .A1(n11401), .A2(n11402), .A3(n11400), .ZN(n11481) );
  OAI211_X1 U13882 ( .C1(n11403), .C2(n11402), .A(n14550), .B(n11481), .ZN(
        n11410) );
  AOI21_X1 U13883 ( .B1(n14552), .B2(n11405), .A(n11404), .ZN(n11406) );
  OAI21_X1 U13884 ( .B1(n14557), .B2(n11407), .A(n11406), .ZN(n11408) );
  INV_X1 U13885 ( .A(n11408), .ZN(n11409) );
  OAI211_X1 U13886 ( .C1(n7106), .C2(n13730), .A(n11410), .B(n11409), .ZN(
        P1_U3231) );
  AOI22_X1 U13887 ( .A1(n13497), .A2(n14831), .B1(n14951), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n11411) );
  OAI21_X1 U13888 ( .B1(n11412), .B2(n14951), .A(n11411), .ZN(P2_U3506) );
  AOI22_X1 U13889 ( .A1(n13497), .A2(n11413), .B1(n14951), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11414) );
  OAI21_X1 U13890 ( .B1(n11415), .B2(n14951), .A(n11414), .ZN(P2_U3508) );
  NOR2_X1 U13891 ( .A1(n11430), .A2(n11416), .ZN(n11418) );
  AOI22_X1 U13892 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n11587), .B1(n11589), 
        .B2(n8455), .ZN(n11419) );
  NOR2_X1 U13893 ( .A1(n11420), .A2(n11419), .ZN(n11584) );
  AOI21_X1 U13894 ( .B1(n11420), .B2(n11419), .A(n11584), .ZN(n11442) );
  INV_X1 U13895 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14509) );
  AOI22_X1 U13896 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n11589), .B1(n11587), 
        .B2(n14509), .ZN(n11426) );
  NAND2_X1 U13897 ( .A1(n11422), .A2(n11421), .ZN(n11424) );
  NAND2_X1 U13898 ( .A1(n11424), .A2(n11423), .ZN(n11425) );
  NAND2_X1 U13899 ( .A1(n11426), .A2(n11425), .ZN(n11586) );
  OAI21_X1 U13900 ( .B1(n11426), .B2(n11425), .A(n11586), .ZN(n11440) );
  INV_X1 U13901 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14287) );
  NAND2_X1 U13902 ( .A1(n15056), .A2(n11587), .ZN(n11428) );
  OAI211_X1 U13903 ( .C1(n14287), .C2(n15074), .A(n11428), .B(n11427), .ZN(
        n11439) );
  MUX2_X1 U13904 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12516), .Z(n11590) );
  XNOR2_X1 U13905 ( .A(n11590), .B(n11587), .ZN(n11433) );
  INV_X1 U13906 ( .A(n11429), .ZN(n11431) );
  NAND2_X1 U13907 ( .A1(n11431), .A2(n11430), .ZN(n11434) );
  AND2_X1 U13908 ( .A1(n11433), .A2(n11434), .ZN(n11432) );
  NAND2_X1 U13909 ( .A1(n11435), .A2(n11432), .ZN(n11595) );
  INV_X1 U13910 ( .A(n11595), .ZN(n11437) );
  AOI21_X1 U13911 ( .B1(n11435), .B2(n11434), .A(n11433), .ZN(n11436) );
  NOR3_X1 U13912 ( .A1(n11437), .A2(n11436), .A3(n15067), .ZN(n11438) );
  AOI211_X1 U13913 ( .C1(n15058), .C2(n11440), .A(n11439), .B(n11438), .ZN(
        n11441) );
  OAI21_X1 U13914 ( .B1(n11442), .B2(n15061), .A(n11441), .ZN(P3_U3194) );
  AOI22_X1 U13915 ( .A1(n13497), .A2(n11457), .B1(n14951), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11443) );
  OAI21_X1 U13916 ( .B1(n11444), .B2(n14951), .A(n11443), .ZN(P2_U3510) );
  AOI22_X1 U13917 ( .A1(n13497), .A2(n11445), .B1(n14951), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n11446) );
  OAI21_X1 U13918 ( .B1(n11447), .B2(n14951), .A(n11446), .ZN(P2_U3509) );
  NAND2_X1 U13919 ( .A1(n11457), .A2(n11448), .ZN(n11449) );
  INV_X1 U13920 ( .A(n13171), .ZN(n11451) );
  NAND2_X1 U13921 ( .A1(n11452), .A2(n14537), .ZN(n11453) );
  XNOR2_X1 U13922 ( .A(n11535), .B(n11534), .ZN(n11454) );
  AOI22_X1 U13923 ( .A1(n13144), .A2(n13169), .B1(n13171), .B2(n13142), .ZN(
        n11707) );
  OAI21_X1 U13924 ( .B1(n11454), .B2(n13368), .A(n11707), .ZN(n11550) );
  INV_X1 U13925 ( .A(n11550), .ZN(n11466) );
  AND2_X1 U13926 ( .A1(n14522), .A2(n13171), .ZN(n11458) );
  OR2_X1 U13927 ( .A1(n14522), .A2(n13171), .ZN(n11459) );
  INV_X1 U13928 ( .A(n11534), .ZN(n11460) );
  XNOR2_X1 U13929 ( .A(n11541), .B(n11460), .ZN(n11552) );
  INV_X1 U13930 ( .A(n11461), .ZN(n14526) );
  AOI211_X1 U13931 ( .C1(n11696), .C2(n14526), .A(n14849), .B(n11544), .ZN(
        n11551) );
  NAND2_X1 U13932 ( .A1(n11551), .A2(n14854), .ZN(n11463) );
  AOI22_X1 U13933 ( .A1(n14873), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11709), 
        .B2(n14844), .ZN(n11462) );
  OAI211_X1 U13934 ( .C1(n11712), .C2(n13420), .A(n11463), .B(n11462), .ZN(
        n11464) );
  AOI21_X1 U13935 ( .B1(n11552), .B2(n14855), .A(n11464), .ZN(n11465) );
  OAI21_X1 U13936 ( .B1(n11466), .B2(n14873), .A(n11465), .ZN(P2_U3252) );
  XNOR2_X1 U13937 ( .A(n11468), .B(n11467), .ZN(n14580) );
  OAI21_X1 U13938 ( .B1(n6586), .B2(n11969), .A(n11469), .ZN(n14583) );
  INV_X1 U13939 ( .A(n11470), .ZN(n11572) );
  INV_X1 U13940 ( .A(n13738), .ZN(n14579) );
  OAI211_X1 U13941 ( .C1(n11572), .C2(n14579), .A(n14655), .B(n11604), .ZN(
        n14578) );
  OR2_X1 U13942 ( .A1(n12016), .A2(n13711), .ZN(n11472) );
  NAND2_X1 U13943 ( .A1(n13757), .A2(n6462), .ZN(n11471) );
  AND2_X1 U13944 ( .A1(n11472), .A2(n11471), .ZN(n14577) );
  INV_X1 U13945 ( .A(n14577), .ZN(n11473) );
  AOI22_X1 U13946 ( .A1(n14389), .A2(n11473), .B1(n13733), .B2(n14680), .ZN(
        n11474) );
  OAI21_X1 U13947 ( .B1(n11475), .B2(n14389), .A(n11474), .ZN(n11476) );
  AOI21_X1 U13948 ( .B1(n13738), .B2(n14398), .A(n11476), .ZN(n11477) );
  OAI21_X1 U13949 ( .B1(n14578), .B2(n14090), .A(n11477), .ZN(n11478) );
  AOI21_X1 U13950 ( .B1(n14583), .B2(n14677), .A(n11478), .ZN(n11479) );
  OAI21_X1 U13951 ( .B1(n14580), .B2(n14050), .A(n11479), .ZN(P1_U3278) );
  INV_X1 U13952 ( .A(n11480), .ZN(n11482) );
  NOR2_X1 U13953 ( .A1(n9620), .A2(n11484), .ZN(n11485) );
  AOI21_X1 U13954 ( .B1(n14747), .B2(n12125), .A(n11485), .ZN(n11644) );
  AOI22_X1 U13955 ( .A1(n14747), .A2(n12118), .B1(n12125), .B2(n13763), .ZN(
        n11486) );
  XNOR2_X1 U13956 ( .A(n11486), .B(n12132), .ZN(n11643) );
  XOR2_X1 U13957 ( .A(n11644), .B(n11643), .Z(n11648) );
  XNOR2_X1 U13958 ( .A(n11649), .B(n11648), .ZN(n11495) );
  AOI21_X1 U13959 ( .B1(n14552), .B2(n11488), .A(n11487), .ZN(n11489) );
  OAI21_X1 U13960 ( .B1(n11490), .B2(n11641), .A(n11489), .ZN(n11493) );
  NOR2_X1 U13961 ( .A1(n14557), .A2(n11491), .ZN(n11492) );
  AOI211_X1 U13962 ( .C1(n14747), .C2(n14554), .A(n11493), .B(n11492), .ZN(
        n11494) );
  OAI21_X1 U13963 ( .B1(n11495), .B2(n13740), .A(n11494), .ZN(P1_U3217) );
  INV_X1 U13964 ( .A(n11496), .ZN(n11498) );
  INV_X1 U13965 ( .A(SI_26_), .ZN(n11497) );
  OAI222_X1 U13966 ( .A1(n11499), .A2(P3_U3151), .B1(n6460), .B2(n11498), .C1(
        n11497), .C2(n12966), .ZN(P3_U3269) );
  OAI211_X1 U13967 ( .C1(n11502), .C2(n11501), .A(n11500), .B(n14960), .ZN(
        n11506) );
  INV_X1 U13968 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n15013) );
  OAI22_X1 U13969 ( .A1(n14425), .A2(n15132), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15013), .ZN(n11504) );
  OAI22_X1 U13970 ( .A1(n12440), .A2(n15127), .B1(n15163), .B2(n12414), .ZN(
        n11503) );
  AOI211_X1 U13971 ( .C1(n15133), .C2(n14436), .A(n11504), .B(n11503), .ZN(
        n11505) );
  NAND2_X1 U13972 ( .A1(n11506), .A2(n11505), .ZN(P3_U3153) );
  AOI21_X1 U13973 ( .B1(n11508), .B2(P2_REG1_REG_16__SCAN_IN), .A(n11507), 
        .ZN(n11510) );
  XNOR2_X1 U13974 ( .A(n13188), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n11509) );
  NOR2_X1 U13975 ( .A1(n11510), .A2(n11509), .ZN(n13187) );
  AOI211_X1 U13976 ( .C1(n11510), .C2(n11509), .A(n13187), .B(n14803), .ZN(
        n11522) );
  INV_X1 U13977 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n11519) );
  OR2_X1 U13978 ( .A1(n13188), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11512) );
  NAND2_X1 U13979 ( .A1(n13188), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11511) );
  AND2_X1 U13980 ( .A1(n11512), .A2(n11511), .ZN(n11517) );
  INV_X1 U13981 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11514) );
  OAI21_X1 U13982 ( .B1(n11515), .B2(n11514), .A(n11513), .ZN(n11516) );
  NAND2_X1 U13983 ( .A1(n11517), .A2(n11516), .ZN(n13183) );
  OAI211_X1 U13984 ( .C1(n11517), .C2(n11516), .A(n14820), .B(n13183), .ZN(
        n11518) );
  OAI21_X1 U13985 ( .B1(n14825), .B2(n11519), .A(n11518), .ZN(n11521) );
  AND2_X1 U13986 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n11520) );
  NOR3_X1 U13987 ( .A1(n11522), .A2(n11521), .A3(n11520), .ZN(n11523) );
  OAI21_X1 U13988 ( .B1(n13184), .B2(n11524), .A(n11523), .ZN(P2_U3231) );
  XNOR2_X1 U13989 ( .A(n14522), .B(n6682), .ZN(n11701) );
  NAND2_X1 U13990 ( .A1(n13171), .A2(n12981), .ZN(n11699) );
  XNOR2_X1 U13991 ( .A(n11701), .B(n11699), .ZN(n11527) );
  NAND2_X1 U13992 ( .A1(n11528), .A2(n11527), .ZN(n11700) );
  OAI21_X1 U13993 ( .B1(n11528), .B2(n11527), .A(n11700), .ZN(n11529) );
  NAND2_X1 U13994 ( .A1(n11529), .A2(n13129), .ZN(n11533) );
  AOI22_X1 U13995 ( .A1(n13144), .A2(n13170), .B1(n13172), .B2(n13142), .ZN(
        n14518) );
  OAI21_X1 U13996 ( .B1(n13147), .B2(n14518), .A(n11530), .ZN(n11531) );
  AOI21_X1 U13997 ( .B1(n14521), .B2(n13145), .A(n11531), .ZN(n11532) );
  OAI211_X1 U13998 ( .C1(n14537), .C2(n13137), .A(n11533), .B(n11532), .ZN(
        P2_U3196) );
  NAND2_X1 U13999 ( .A1(n11535), .A2(n11534), .ZN(n11538) );
  OR2_X1 U14000 ( .A1(n11696), .A2(n11536), .ZN(n11537) );
  NAND2_X1 U14001 ( .A1(n11538), .A2(n11537), .ZN(n11659) );
  XNOR2_X1 U14002 ( .A(n11659), .B(n11543), .ZN(n11539) );
  AOI22_X1 U14003 ( .A1(n13144), .A2(n13168), .B1(n13170), .B2(n13142), .ZN(
        n11731) );
  OAI21_X1 U14004 ( .B1(n11539), .B2(n13368), .A(n11731), .ZN(n14532) );
  INV_X1 U14005 ( .A(n14532), .ZN(n11549) );
  NOR2_X1 U14006 ( .A1(n11696), .A2(n13170), .ZN(n11540) );
  NAND2_X1 U14007 ( .A1(n11696), .A2(n13170), .ZN(n11542) );
  XNOR2_X1 U14008 ( .A(n11667), .B(n11543), .ZN(n14534) );
  OAI211_X1 U14009 ( .C1(n6663), .C2(n11544), .A(n13405), .B(n11663), .ZN(
        n14531) );
  AOI22_X1 U14010 ( .A1(n14873), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11733), 
        .B2(n14844), .ZN(n11546) );
  NAND2_X1 U14011 ( .A1(n11727), .A2(n14846), .ZN(n11545) );
  OAI211_X1 U14012 ( .C1(n14531), .C2(n14833), .A(n11546), .B(n11545), .ZN(
        n11547) );
  AOI21_X1 U14013 ( .B1(n14534), .B2(n14855), .A(n11547), .ZN(n11548) );
  OAI21_X1 U14014 ( .B1(n11549), .B2(n14873), .A(n11548), .ZN(P2_U3251) );
  AOI211_X1 U14015 ( .C1(n11552), .C2(n14921), .A(n11551), .B(n11550), .ZN(
        n11557) );
  AOI22_X1 U14016 ( .A1(n11696), .A2(n13497), .B1(n14951), .B2(
        P2_REG1_REG_13__SCAN_IN), .ZN(n11553) );
  OAI21_X1 U14017 ( .B1(n11557), .B2(n14951), .A(n11553), .ZN(P2_U3512) );
  INV_X1 U14018 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11554) );
  OAI22_X1 U14019 ( .A1(n11712), .A2(n13557), .B1(n14942), .B2(n11554), .ZN(
        n11555) );
  INV_X1 U14020 ( .A(n11555), .ZN(n11556) );
  OAI21_X1 U14021 ( .B1(n11557), .B2(n14940), .A(n11556), .ZN(P2_U3469) );
  INV_X1 U14022 ( .A(n11558), .ZN(n11560) );
  OAI222_X1 U14023 ( .A1(n6461), .A2(n11560), .B1(n12966), .B2(n11559), .C1(
        P3_U3151), .C2(n9654), .ZN(P3_U3268) );
  OAI211_X1 U14024 ( .C1(n11563), .C2(n11562), .A(n11561), .B(n14960), .ZN(
        n11568) );
  OAI22_X1 U14025 ( .A1(n14425), .A2(n15116), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11564), .ZN(n11566) );
  OAI22_X1 U14026 ( .A1(n12440), .A2(n15112), .B1(n15111), .B2(n12414), .ZN(
        n11565) );
  AOI211_X1 U14027 ( .C1(n15117), .C2(n14436), .A(n11566), .B(n11565), .ZN(
        n11567) );
  NAND2_X1 U14028 ( .A1(n11568), .A2(n11567), .ZN(P3_U3161) );
  NAND2_X1 U14029 ( .A1(n11569), .A2(n11968), .ZN(n11570) );
  AOI211_X1 U14030 ( .C1(n14558), .C2(n11573), .A(n14674), .B(n11572), .ZN(
        n14565) );
  OAI211_X1 U14031 ( .C1(n11575), .C2(n11968), .A(n11574), .B(n14664), .ZN(
        n11579) );
  OR2_X1 U14032 ( .A1(n12024), .A2(n13713), .ZN(n11577) );
  OR2_X1 U14033 ( .A1(n11840), .A2(n13711), .ZN(n11576) );
  NAND2_X1 U14034 ( .A1(n11577), .A2(n11576), .ZN(n14553) );
  INV_X1 U14035 ( .A(n14553), .ZN(n11578) );
  NAND2_X1 U14036 ( .A1(n11579), .A2(n11578), .ZN(n14562) );
  AOI211_X1 U14037 ( .C1(n14566), .C2(n14753), .A(n14565), .B(n14562), .ZN(
        n11583) );
  INV_X1 U14038 ( .A(n14232), .ZN(n14221) );
  NOR2_X1 U14039 ( .A1(n14756), .A2(n7895), .ZN(n11580) );
  AOI21_X1 U14040 ( .B1(n14558), .B2(n14221), .A(n11580), .ZN(n11581) );
  OAI21_X1 U14041 ( .B1(n11583), .B2(n14755), .A(n11581), .ZN(P1_U3501) );
  AOI22_X1 U14042 ( .A1(n14558), .A2(n14162), .B1(n14764), .B2(
        P1_REG1_REG_14__SCAN_IN), .ZN(n11582) );
  OAI21_X1 U14043 ( .B1(n11583), .B2(n14764), .A(n11582), .ZN(P1_U3542) );
  AOI21_X1 U14044 ( .B1(n8480), .B2(n11585), .A(n12465), .ZN(n11602) );
  XNOR2_X1 U14045 ( .A(n12468), .B(n12480), .ZN(n11588) );
  NAND2_X1 U14046 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n11588), .ZN(n12470) );
  OAI21_X1 U14047 ( .B1(n11588), .B2(P3_REG1_REG_13__SCAN_IN), .A(n12470), 
        .ZN(n11600) );
  NAND2_X1 U14048 ( .A1(n11590), .A2(n11589), .ZN(n11592) );
  MUX2_X1 U14049 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12516), .Z(n12479) );
  XNOR2_X1 U14050 ( .A(n12479), .B(n12480), .ZN(n11593) );
  AOI21_X1 U14051 ( .B1(n11595), .B2(n11592), .A(n11593), .ZN(n11591) );
  INV_X1 U14052 ( .A(n11591), .ZN(n11596) );
  AND2_X1 U14053 ( .A1(n11593), .A2(n11592), .ZN(n11594) );
  NAND2_X1 U14054 ( .A1(n11595), .A2(n11594), .ZN(n12487) );
  AOI21_X1 U14055 ( .B1(n11596), .B2(n12487), .A(n15067), .ZN(n11599) );
  NAND2_X1 U14056 ( .A1(n15056), .A2(n12480), .ZN(n11597) );
  NAND2_X1 U14057 ( .A1(P3_REG3_REG_13__SCAN_IN), .A2(P3_U3151), .ZN(n12394)
         );
  OAI211_X1 U14058 ( .C1(n14291), .C2(n15074), .A(n11597), .B(n12394), .ZN(
        n11598) );
  AOI211_X1 U14059 ( .C1(n11600), .C2(n15058), .A(n11599), .B(n11598), .ZN(
        n11601) );
  OAI21_X1 U14060 ( .B1(n11602), .B2(n15061), .A(n11601), .ZN(P3_U3195) );
  XNOR2_X1 U14061 ( .A(n11603), .B(n11972), .ZN(n14573) );
  OAI22_X1 U14062 ( .A1(n14389), .A2(n11627), .B1(n13655), .B2(n14667), .ZN(
        n11609) );
  AOI211_X1 U14063 ( .C1(n14571), .C2(n11604), .A(n14674), .B(n14082), .ZN(
        n14569) );
  NAND2_X1 U14064 ( .A1(n13756), .A2(n6462), .ZN(n11606) );
  OR2_X1 U14065 ( .A1(n12024), .A2(n13711), .ZN(n11605) );
  NAND2_X1 U14066 ( .A1(n11606), .A2(n11605), .ZN(n14570) );
  AOI21_X1 U14067 ( .B1(n14569), .B2(n14564), .A(n14570), .ZN(n11607) );
  NOR2_X1 U14068 ( .A1(n11607), .A2(n6476), .ZN(n11608) );
  AOI211_X1 U14069 ( .C1(n14398), .C2(n14571), .A(n11609), .B(n11608), .ZN(
        n11613) );
  XNOR2_X1 U14070 ( .A(n11611), .B(n11610), .ZN(n14575) );
  NAND2_X1 U14071 ( .A1(n14575), .A2(n14055), .ZN(n11612) );
  OAI211_X1 U14072 ( .C1(n14573), .C2(n14077), .A(n11613), .B(n11612), .ZN(
        P1_U3277) );
  INV_X1 U14073 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n11619) );
  AOI21_X1 U14074 ( .B1(n11615), .B2(P1_REG1_REG_16__SCAN_IN), .A(n11614), 
        .ZN(n13863) );
  INV_X1 U14075 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n11616) );
  OR2_X1 U14076 ( .A1(n11623), .A2(n11616), .ZN(n11618) );
  NAND2_X1 U14077 ( .A1(n11623), .A2(n11616), .ZN(n11617) );
  AND2_X1 U14078 ( .A1(n11618), .A2(n11617), .ZN(n13862) );
  NOR2_X1 U14079 ( .A1(n13863), .A2(n13862), .ZN(n13861) );
  AOI21_X1 U14080 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n11623), .A(n13861), 
        .ZN(n11620) );
  XNOR2_X1 U14081 ( .A(n13874), .B(n11620), .ZN(n13881) );
  NOR2_X1 U14082 ( .A1(n11619), .A2(n13881), .ZN(n13882) );
  NOR2_X1 U14083 ( .A1(n11620), .A2(n13874), .ZN(n11621) );
  NOR2_X1 U14084 ( .A1(n13882), .A2(n11621), .ZN(n11622) );
  XOR2_X1 U14085 ( .A(n11622), .B(n14176), .Z(n11636) );
  INV_X1 U14086 ( .A(n11636), .ZN(n11634) );
  INV_X1 U14087 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14086) );
  OR2_X1 U14088 ( .A1(n11623), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11625) );
  NAND2_X1 U14089 ( .A1(n11623), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n11624) );
  AND2_X1 U14090 ( .A1(n11625), .A2(n11624), .ZN(n13870) );
  OAI21_X1 U14091 ( .B1(n11628), .B2(n11627), .A(n11626), .ZN(n13869) );
  NAND2_X1 U14092 ( .A1(n13870), .A2(n13869), .ZN(n13868) );
  OAI21_X1 U14093 ( .B1(n14086), .B2(n13865), .A(n13868), .ZN(n11630) );
  NAND2_X1 U14094 ( .A1(n11629), .A2(n11630), .ZN(n11631) );
  XNOR2_X1 U14095 ( .A(n13874), .B(n11630), .ZN(n13880) );
  NAND2_X1 U14096 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n13880), .ZN(n13878) );
  NAND2_X1 U14097 ( .A1(n11631), .A2(n13878), .ZN(n11632) );
  XOR2_X1 U14098 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n11632), .Z(n11635) );
  OAI21_X1 U14099 ( .B1(n11635), .B2(n14627), .A(n14636), .ZN(n11633) );
  AOI21_X1 U14100 ( .B1(n11634), .B2(n14631), .A(n11633), .ZN(n11638) );
  AOI22_X1 U14101 ( .A1(n11636), .A2(n14631), .B1(n13879), .B2(n11635), .ZN(
        n11637) );
  MUX2_X1 U14102 ( .A(n11638), .B(n11637), .S(n14564), .Z(n11640) );
  AND2_X1 U14103 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13629) );
  INV_X1 U14104 ( .A(n13629), .ZN(n11639) );
  OAI211_X1 U14105 ( .C1(n7418), .C2(n14640), .A(n11640), .B(n11639), .ZN(
        P1_U3262) );
  OAI22_X1 U14106 ( .A1(n14593), .A2(n11717), .B1(n11641), .B2(n9620), .ZN(
        n11679) );
  OAI22_X1 U14107 ( .A1(n14593), .A2(n12131), .B1(n11641), .B2(n11717), .ZN(
        n11642) );
  XNOR2_X1 U14108 ( .A(n11642), .B(n12132), .ZN(n11678) );
  XOR2_X1 U14109 ( .A(n11679), .B(n11678), .Z(n11651) );
  INV_X1 U14110 ( .A(n11643), .ZN(n11646) );
  INV_X1 U14111 ( .A(n11644), .ZN(n11645) );
  OAI21_X1 U14112 ( .B1(n11651), .B2(n11650), .A(n11684), .ZN(n11652) );
  NAND2_X1 U14113 ( .A1(n11652), .A2(n14550), .ZN(n11658) );
  NOR2_X1 U14114 ( .A1(n14557), .A2(n11653), .ZN(n11654) );
  AOI211_X1 U14115 ( .C1(n14552), .C2(n11656), .A(n11655), .B(n11654), .ZN(
        n11657) );
  OAI211_X1 U14116 ( .C1(n14593), .C2(n13730), .A(n11658), .B(n11657), .ZN(
        P1_U3236) );
  INV_X1 U14117 ( .A(n13169), .ZN(n11660) );
  XOR2_X1 U14118 ( .A(n12146), .B(n12183), .Z(n11661) );
  INV_X1 U14119 ( .A(n13167), .ZN(n12148) );
  OAI22_X1 U14120 ( .A1(n11660), .A2(n13072), .B1(n12148), .B2(n13074), .ZN(
        n11744) );
  AOI21_X1 U14121 ( .B1(n11661), .B2(n14860), .A(n11744), .ZN(n13527) );
  INV_X1 U14122 ( .A(n13417), .ZN(n11662) );
  AOI211_X1 U14123 ( .C1(n13525), .C2(n11663), .A(n14849), .B(n11662), .ZN(
        n13524) );
  INV_X1 U14124 ( .A(n13525), .ZN(n11665) );
  AOI22_X1 U14125 ( .A1(n14873), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n11743), 
        .B2(n14844), .ZN(n11664) );
  OAI21_X1 U14126 ( .B1(n11665), .B2(n13420), .A(n11664), .ZN(n11670) );
  AND2_X1 U14127 ( .A1(n11727), .A2(n13169), .ZN(n11666) );
  OAI22_X1 U14128 ( .A1(n11667), .A2(n11666), .B1(n11727), .B2(n13169), .ZN(
        n12184) );
  INV_X1 U14129 ( .A(n12183), .ZN(n11668) );
  XNOR2_X1 U14130 ( .A(n12184), .B(n11668), .ZN(n13528) );
  NOR2_X1 U14131 ( .A1(n13528), .A2(n13425), .ZN(n11669) );
  AOI211_X1 U14132 ( .C1(n13524), .C2(n14854), .A(n11670), .B(n11669), .ZN(
        n11671) );
  OAI21_X1 U14133 ( .B1(n14873), .B2(n13527), .A(n11671), .ZN(P2_U3250) );
  INV_X1 U14134 ( .A(n11692), .ZN(n11674) );
  AOI21_X1 U14135 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n13585), .A(n11672), 
        .ZN(n11673) );
  OAI21_X1 U14136 ( .B1(n11674), .B2(n13587), .A(n11673), .ZN(P2_U3304) );
  INV_X1 U14137 ( .A(n11675), .ZN(n11676) );
  OAI222_X1 U14138 ( .A1(n13599), .A2(n11677), .B1(P2_U3088), .B2(n9441), .C1(
        n13587), .C2(n11676), .ZN(P2_U3305) );
  INV_X1 U14139 ( .A(n11678), .ZN(n11681) );
  INV_X1 U14140 ( .A(n11679), .ZN(n11680) );
  NAND2_X1 U14141 ( .A1(n11681), .A2(n11680), .ZN(n11683) );
  AND2_X1 U14142 ( .A1(n11684), .A2(n11683), .ZN(n11686) );
  OAI22_X1 U14143 ( .A1(n14407), .A2(n12131), .B1(n11841), .B2(n11717), .ZN(
        n11682) );
  XNOR2_X1 U14144 ( .A(n11682), .B(n12121), .ZN(n11713) );
  OAI22_X1 U14145 ( .A1(n14407), .A2(n11717), .B1(n11841), .B2(n9615), .ZN(
        n11714) );
  XNOR2_X1 U14146 ( .A(n11713), .B(n11714), .ZN(n11685) );
  OAI211_X1 U14147 ( .C1(n11686), .C2(n11685), .A(n14550), .B(n11716), .ZN(
        n11691) );
  OR2_X1 U14148 ( .A1(n11840), .A2(n13713), .ZN(n11688) );
  NAND2_X1 U14149 ( .A1(n13725), .A2(n13762), .ZN(n11687) );
  NAND2_X1 U14150 ( .A1(n11688), .A2(n11687), .ZN(n14395) );
  AND2_X1 U14151 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n13849) );
  NOR2_X1 U14152 ( .A1(n14557), .A2(n14396), .ZN(n11689) );
  AOI211_X1 U14153 ( .C1(n14552), .C2(n14395), .A(n13849), .B(n11689), .ZN(
        n11690) );
  OAI211_X1 U14154 ( .C1(n14407), .C2(n13730), .A(n11691), .B(n11690), .ZN(
        P1_U3224) );
  NAND2_X1 U14155 ( .A1(n11692), .A2(n14235), .ZN(n11693) );
  OAI211_X1 U14156 ( .C1(n11695), .C2(n11694), .A(n11693), .B(n11993), .ZN(
        P1_U3332) );
  XNOR2_X1 U14157 ( .A(n11696), .B(n6682), .ZN(n11698) );
  AND2_X1 U14158 ( .A1(n13170), .A2(n14849), .ZN(n11697) );
  NAND2_X1 U14159 ( .A1(n11698), .A2(n11697), .ZN(n11725) );
  OAI21_X1 U14160 ( .B1(n11698), .B2(n11697), .A(n11725), .ZN(n11704) );
  INV_X1 U14161 ( .A(n11699), .ZN(n11702) );
  AOI211_X1 U14162 ( .C1(n11704), .C2(n11703), .A(n13151), .B(n11726), .ZN(
        n11705) );
  INV_X1 U14163 ( .A(n11705), .ZN(n11711) );
  OAI22_X1 U14164 ( .A1(n13147), .A2(n11707), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11706), .ZN(n11708) );
  AOI21_X1 U14165 ( .B1(n11709), .B2(n13145), .A(n11708), .ZN(n11710) );
  OAI211_X1 U14166 ( .C1(n11712), .C2(n13137), .A(n11711), .B(n11710), .ZN(
        P2_U3206) );
  INV_X1 U14167 ( .A(n11713), .ZN(n11715) );
  OAI22_X1 U14168 ( .A1(n11839), .A2(n11717), .B1(n11840), .B2(n9620), .ZN(
        n12010) );
  OAI22_X1 U14169 ( .A1(n11839), .A2(n12131), .B1(n11840), .B2(n11717), .ZN(
        n11718) );
  XNOR2_X1 U14170 ( .A(n11718), .B(n12132), .ZN(n12011) );
  XOR2_X1 U14171 ( .A(n12010), .B(n12011), .Z(n12008) );
  XNOR2_X1 U14172 ( .A(n12009), .B(n12008), .ZN(n11724) );
  NAND2_X1 U14173 ( .A1(n14552), .A2(n14584), .ZN(n11719) );
  OAI211_X1 U14174 ( .C1(n14557), .C2(n11721), .A(n11720), .B(n11719), .ZN(
        n11722) );
  AOI21_X1 U14175 ( .B1(n14585), .B2(n14554), .A(n11722), .ZN(n11723) );
  OAI21_X1 U14176 ( .B1(n11724), .B2(n13740), .A(n11723), .ZN(P1_U3234) );
  XNOR2_X1 U14177 ( .A(n11727), .B(n6682), .ZN(n11739) );
  NAND2_X1 U14178 ( .A1(n13169), .A2(n12981), .ZN(n11737) );
  XNOR2_X1 U14179 ( .A(n11739), .B(n11737), .ZN(n11728) );
  OAI21_X1 U14180 ( .B1(n6590), .B2(n11728), .A(n11736), .ZN(n11729) );
  NAND2_X1 U14181 ( .A1(n11729), .A2(n13129), .ZN(n11735) );
  OAI21_X1 U14182 ( .B1(n13147), .B2(n11731), .A(n11730), .ZN(n11732) );
  AOI21_X1 U14183 ( .B1(n11733), .B2(n13145), .A(n11732), .ZN(n11734) );
  OAI211_X1 U14184 ( .C1(n6663), .C2(n13137), .A(n11735), .B(n11734), .ZN(
        P2_U3187) );
  INV_X1 U14185 ( .A(n11736), .ZN(n11740) );
  INV_X1 U14186 ( .A(n11737), .ZN(n11738) );
  NOR2_X1 U14187 ( .A1(n11739), .A2(n11738), .ZN(n12968) );
  NOR2_X1 U14188 ( .A1(n11740), .A2(n12968), .ZN(n11742) );
  XNOR2_X1 U14189 ( .A(n13525), .B(n13006), .ZN(n12970) );
  NAND2_X1 U14190 ( .A1(n13168), .A2(n14849), .ZN(n12969) );
  INV_X1 U14191 ( .A(n12969), .ZN(n12972) );
  XNOR2_X1 U14192 ( .A(n12970), .B(n12972), .ZN(n11741) );
  XNOR2_X1 U14193 ( .A(n11742), .B(n11741), .ZN(n11749) );
  INV_X1 U14194 ( .A(n11743), .ZN(n11746) );
  AOI22_X1 U14195 ( .A1(n13097), .A2(n11744), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11745) );
  OAI21_X1 U14196 ( .B1(n11746), .B2(n13104), .A(n11745), .ZN(n11747) );
  AOI21_X1 U14197 ( .B1(n13525), .B2(n13149), .A(n11747), .ZN(n11748) );
  OAI21_X1 U14198 ( .B1(n11749), .B2(n13151), .A(n11748), .ZN(P2_U3213) );
  NAND2_X1 U14199 ( .A1(n11998), .A2(n7923), .ZN(n11752) );
  OR2_X1 U14200 ( .A1(n11750), .A2(n11999), .ZN(n11751) );
  NAND2_X1 U14201 ( .A1(n11755), .A2(n8069), .ZN(n11758) );
  INV_X1 U14202 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14192) );
  NAND2_X1 U14203 ( .A1(n11759), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n11762) );
  NAND2_X1 U14204 ( .A1(n11760), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n11761) );
  OAI211_X1 U14205 ( .C1(n7673), .C2(n14192), .A(n11762), .B(n11761), .ZN(
        n13742) );
  INV_X1 U14206 ( .A(n11763), .ZN(n11764) );
  AOI21_X1 U14207 ( .B1(n11946), .B2(n13742), .A(n11764), .ZN(n11765) );
  OAI22_X1 U14208 ( .A1(n14197), .A2(n11946), .B1(n11927), .B2(n11765), .ZN(
        n11932) );
  INV_X1 U14209 ( .A(n11932), .ZN(n11933) );
  MUX2_X1 U14210 ( .A(n12138), .B(n14108), .S(n11946), .Z(n11924) );
  INV_X1 U14211 ( .A(n11924), .ZN(n11926) );
  MUX2_X1 U14212 ( .A(n13748), .B(n13972), .S(n11946), .Z(n11908) );
  NAND2_X1 U14213 ( .A1(n11767), .A2(n11766), .ZN(n11768) );
  NAND2_X1 U14214 ( .A1(n11768), .A2(n11773), .ZN(n11770) );
  NAND2_X1 U14215 ( .A1(n11774), .A2(n11773), .ZN(n11775) );
  MUX2_X1 U14216 ( .A(n11778), .B(n13772), .S(n11929), .Z(n11780) );
  NAND2_X1 U14217 ( .A1(n13772), .A2(n11778), .ZN(n11779) );
  AOI21_X1 U14218 ( .B1(n11780), .B2(n11779), .A(n11956), .ZN(n11781) );
  NAND2_X1 U14219 ( .A1(n11782), .A2(n11781), .ZN(n11790) );
  INV_X1 U14220 ( .A(n11783), .ZN(n11786) );
  INV_X1 U14221 ( .A(n11784), .ZN(n11785) );
  MUX2_X1 U14222 ( .A(n11786), .B(n11785), .S(n11929), .Z(n11787) );
  INV_X1 U14223 ( .A(n11787), .ZN(n11788) );
  NAND3_X1 U14224 ( .A1(n11790), .A2(n11789), .A3(n11788), .ZN(n11797) );
  INV_X1 U14225 ( .A(n11791), .ZN(n11794) );
  INV_X1 U14226 ( .A(n11792), .ZN(n11793) );
  INV_X1 U14227 ( .A(n11795), .ZN(n11796) );
  NAND2_X1 U14228 ( .A1(n11797), .A2(n11796), .ZN(n11801) );
  MUX2_X1 U14229 ( .A(n11798), .B(n14708), .S(n11929), .Z(n11800) );
  MUX2_X1 U14230 ( .A(n14676), .B(n13769), .S(n11929), .Z(n11799) );
  OAI21_X1 U14231 ( .B1(n11801), .B2(n11800), .A(n11799), .ZN(n11803) );
  NAND2_X1 U14232 ( .A1(n11801), .A2(n11800), .ZN(n11802) );
  NAND2_X1 U14233 ( .A1(n11803), .A2(n11802), .ZN(n11807) );
  MUX2_X1 U14234 ( .A(n11804), .B(n13768), .S(n11929), .Z(n11806) );
  MUX2_X1 U14235 ( .A(n13767), .B(n14648), .S(n11946), .Z(n11811) );
  MUX2_X1 U14236 ( .A(n13767), .B(n14648), .S(n11771), .Z(n11808) );
  NAND2_X1 U14237 ( .A1(n11809), .A2(n11808), .ZN(n11815) );
  INV_X1 U14238 ( .A(n11810), .ZN(n11813) );
  INV_X1 U14239 ( .A(n11811), .ZN(n11812) );
  NAND2_X1 U14240 ( .A1(n11813), .A2(n11812), .ZN(n11814) );
  NAND2_X1 U14241 ( .A1(n11815), .A2(n11814), .ZN(n11817) );
  MUX2_X1 U14242 ( .A(n13766), .B(n14725), .S(n11771), .Z(n11818) );
  MUX2_X1 U14243 ( .A(n13766), .B(n14725), .S(n11946), .Z(n11816) );
  INV_X1 U14244 ( .A(n11818), .ZN(n11819) );
  MUX2_X1 U14245 ( .A(n13765), .B(n11820), .S(n11946), .Z(n11824) );
  MUX2_X1 U14246 ( .A(n13765), .B(n11820), .S(n11771), .Z(n11821) );
  NAND2_X1 U14247 ( .A1(n11822), .A2(n11821), .ZN(n11828) );
  INV_X1 U14248 ( .A(n11823), .ZN(n11826) );
  INV_X1 U14249 ( .A(n11824), .ZN(n11825) );
  NAND2_X1 U14250 ( .A1(n11828), .A2(n11827), .ZN(n11831) );
  MUX2_X1 U14251 ( .A(n13764), .B(n11829), .S(n11771), .Z(n11832) );
  MUX2_X1 U14252 ( .A(n13764), .B(n11829), .S(n11946), .Z(n11830) );
  INV_X1 U14253 ( .A(n11832), .ZN(n11833) );
  MUX2_X1 U14254 ( .A(n13763), .B(n14747), .S(n11946), .Z(n11836) );
  MUX2_X1 U14255 ( .A(n13763), .B(n14747), .S(n11771), .Z(n11834) );
  MUX2_X1 U14256 ( .A(n13762), .B(n11837), .S(n11771), .Z(n11843) );
  MUX2_X1 U14257 ( .A(n13762), .B(n11837), .S(n11946), .Z(n11838) );
  MUX2_X1 U14258 ( .A(n11840), .B(n11839), .S(n11771), .Z(n11849) );
  MUX2_X1 U14259 ( .A(n13760), .B(n14585), .S(n11946), .Z(n11850) );
  MUX2_X1 U14260 ( .A(n11841), .B(n14407), .S(n11771), .Z(n11846) );
  MUX2_X1 U14261 ( .A(n13761), .B(n14399), .S(n11946), .Z(n11845) );
  AOI22_X1 U14262 ( .A1(n11849), .A2(n11850), .B1(n11846), .B2(n11845), .ZN(
        n11842) );
  INV_X1 U14263 ( .A(n11845), .ZN(n11848) );
  INV_X1 U14264 ( .A(n11846), .ZN(n11847) );
  INV_X1 U14265 ( .A(n11849), .ZN(n11852) );
  INV_X1 U14266 ( .A(n11850), .ZN(n11851) );
  OAI21_X1 U14267 ( .B1(n11853), .B2(n11852), .A(n11851), .ZN(n11855) );
  NAND2_X1 U14268 ( .A1(n11853), .A2(n11852), .ZN(n11854) );
  AND2_X1 U14269 ( .A1(n11863), .A2(n11857), .ZN(n11860) );
  AND2_X1 U14270 ( .A1(n11862), .A2(n11858), .ZN(n11859) );
  MUX2_X1 U14271 ( .A(n11860), .B(n11859), .S(n11771), .Z(n11861) );
  MUX2_X1 U14272 ( .A(n11863), .B(n11862), .S(n11946), .Z(n11864) );
  NAND2_X1 U14273 ( .A1(n11865), .A2(n11864), .ZN(n11867) );
  MUX2_X1 U14274 ( .A(n13757), .B(n14571), .S(n11771), .Z(n11868) );
  MUX2_X1 U14275 ( .A(n13757), .B(n14571), .S(n11946), .Z(n11866) );
  INV_X1 U14276 ( .A(n11868), .ZN(n11869) );
  MUX2_X1 U14277 ( .A(n13712), .B(n14233), .S(n11946), .Z(n11871) );
  MUX2_X1 U14278 ( .A(n13668), .B(n14074), .S(n11946), .Z(n11872) );
  NAND2_X1 U14279 ( .A1(n11875), .A2(n11874), .ZN(n11876) );
  NAND3_X1 U14280 ( .A1(n11877), .A2(n11876), .A3(n14051), .ZN(n11881) );
  MUX2_X1 U14281 ( .A(n11879), .B(n11878), .S(n11771), .Z(n11880) );
  NAND2_X1 U14282 ( .A1(n11881), .A2(n11880), .ZN(n11885) );
  MUX2_X1 U14283 ( .A(n14043), .B(n13753), .S(n11946), .Z(n11882) );
  INV_X1 U14284 ( .A(n11882), .ZN(n11884) );
  MUX2_X1 U14285 ( .A(n13753), .B(n14043), .S(n11946), .Z(n11883) );
  NAND2_X1 U14286 ( .A1(n11885), .A2(n11884), .ZN(n11886) );
  MUX2_X1 U14287 ( .A(n13752), .B(n14220), .S(n11946), .Z(n11889) );
  MUX2_X1 U14288 ( .A(n14220), .B(n13752), .S(n11946), .Z(n11888) );
  MUX2_X1 U14289 ( .A(n14217), .B(n13635), .S(n11946), .Z(n11893) );
  MUX2_X1 U14290 ( .A(n13635), .B(n14217), .S(n11946), .Z(n11890) );
  INV_X1 U14291 ( .A(n11890), .ZN(n11891) );
  MUX2_X1 U14292 ( .A(n13750), .B(n14212), .S(n11946), .Z(n11897) );
  MUX2_X1 U14293 ( .A(n14212), .B(n13750), .S(n11946), .Z(n11894) );
  NAND2_X1 U14294 ( .A1(n11895), .A2(n11894), .ZN(n11901) );
  INV_X1 U14295 ( .A(n11896), .ZN(n11899) );
  INV_X1 U14296 ( .A(n11897), .ZN(n11898) );
  MUX2_X1 U14297 ( .A(n13749), .B(n14132), .S(n11946), .Z(n11902) );
  NAND2_X1 U14298 ( .A1(n11907), .A2(n11908), .ZN(n11905) );
  MUX2_X1 U14299 ( .A(n13972), .B(n13748), .S(n11946), .Z(n11904) );
  NAND2_X1 U14300 ( .A1(n11905), .A2(n11904), .ZN(n11906) );
  MUX2_X1 U14301 ( .A(n14120), .B(n13747), .S(n11946), .Z(n11911) );
  MUX2_X1 U14302 ( .A(n14120), .B(n13747), .S(n11771), .Z(n11909) );
  MUX2_X1 U14303 ( .A(n13746), .B(n13939), .S(n11946), .Z(n11914) );
  MUX2_X1 U14304 ( .A(n13746), .B(n13939), .S(n11771), .Z(n11912) );
  NAND2_X1 U14305 ( .A1(n11913), .A2(n11912), .ZN(n11916) );
  INV_X1 U14306 ( .A(n11914), .ZN(n11915) );
  MUX2_X1 U14307 ( .A(n13745), .B(n13915), .S(n11771), .Z(n11917) );
  NAND2_X1 U14308 ( .A1(n11918), .A2(n11917), .ZN(n11921) );
  MUX2_X1 U14309 ( .A(n13745), .B(n13915), .S(n11946), .Z(n11920) );
  MUX2_X1 U14310 ( .A(n11922), .B(n13744), .S(n11946), .Z(n11923) );
  INV_X1 U14311 ( .A(n11927), .ZN(n13743) );
  OAI21_X1 U14312 ( .B1(n13742), .B2(n11928), .A(n13743), .ZN(n11930) );
  MUX2_X1 U14313 ( .A(n11930), .B(n14197), .S(n11946), .Z(n11931) );
  NAND2_X1 U14314 ( .A1(n14236), .A2(n7923), .ZN(n11937) );
  NAND2_X1 U14315 ( .A1(n11935), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n11936) );
  XNOR2_X1 U14316 ( .A(n11945), .B(n13742), .ZN(n11982) );
  NAND2_X1 U14317 ( .A1(n11939), .A2(n11938), .ZN(n11940) );
  NAND2_X1 U14318 ( .A1(n11941), .A2(n11940), .ZN(n11943) );
  NAND2_X1 U14319 ( .A1(n11943), .A2(n11942), .ZN(n11949) );
  INV_X1 U14320 ( .A(n11949), .ZN(n11944) );
  NOR2_X1 U14321 ( .A1(n11944), .A2(n11984), .ZN(n11985) );
  INV_X1 U14322 ( .A(n11985), .ZN(n11951) );
  INV_X1 U14323 ( .A(n13742), .ZN(n13889) );
  NOR2_X1 U14324 ( .A1(n11945), .A2(n13889), .ZN(n11948) );
  NOR2_X1 U14325 ( .A1(n14193), .A2(n13742), .ZN(n11947) );
  MUX2_X1 U14326 ( .A(n11948), .B(n11947), .S(n11946), .Z(n11986) );
  NOR2_X1 U14327 ( .A1(n11986), .A2(n11949), .ZN(n11950) );
  NAND2_X1 U14328 ( .A1(n11954), .A2(n11953), .ZN(n11955) );
  NOR4_X1 U14329 ( .A1(n14671), .A2(n11957), .A3(n11956), .A4(n11955), .ZN(
        n11961) );
  NAND4_X1 U14330 ( .A1(n11961), .A2(n11960), .A3(n11959), .A4(n11958), .ZN(
        n11962) );
  NOR4_X1 U14331 ( .A1(n11965), .A2(n11964), .A3(n11963), .A4(n11962), .ZN(
        n11967) );
  NAND4_X1 U14332 ( .A1(n11968), .A2(n11967), .A3(n11966), .A4(n14391), .ZN(
        n11971) );
  NOR4_X1 U14333 ( .A1(n14091), .A2(n11971), .A3(n11970), .A4(n11969), .ZN(
        n11973) );
  NAND4_X1 U14334 ( .A1(n14051), .A2(n11973), .A3(n14076), .A4(n11972), .ZN(
        n11974) );
  NOR4_X1 U14335 ( .A1(n14009), .A2(n14021), .A3(n11975), .A4(n11974), .ZN(
        n11976) );
  NAND4_X1 U14336 ( .A1(n13953), .A2(n11976), .A3(n13995), .A4(n13980), .ZN(
        n11977) );
  NOR4_X1 U14337 ( .A1(n13922), .A2(n11978), .A3(n13968), .A4(n11977), .ZN(
        n11981) );
  XNOR2_X1 U14338 ( .A(n13894), .B(n13743), .ZN(n11979) );
  NAND4_X1 U14339 ( .A1(n11982), .A2(n11981), .A3(n11980), .A4(n11979), .ZN(
        n11983) );
  XOR2_X1 U14340 ( .A(n14564), .B(n11983), .Z(n11989) );
  INV_X1 U14341 ( .A(n11984), .ZN(n11988) );
  AOI21_X1 U14342 ( .B1(n11986), .B2(n11985), .A(n11993), .ZN(n11987) );
  OAI21_X1 U14343 ( .B1(n11989), .B2(n11988), .A(n11987), .ZN(n11996) );
  NAND2_X1 U14344 ( .A1(n11990), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11991) );
  NOR3_X1 U14345 ( .A1(n11992), .A2(n13711), .A3(n11991), .ZN(n11995) );
  OAI21_X1 U14346 ( .B1(n11993), .B2(n14264), .A(P1_B_REG_SCAN_IN), .ZN(n11994) );
  OAI22_X1 U14347 ( .A1(n11997), .A2(n11996), .B1(n11995), .B2(n11994), .ZN(
        P1_U3242) );
  INV_X1 U14348 ( .A(n11998), .ZN(n13579) );
  OAI222_X1 U14349 ( .A1(n14262), .A2(n13579), .B1(P1_U3086), .B2(n12000), 
        .C1(n11999), .C2(n14258), .ZN(P1_U3325) );
  AOI21_X1 U14350 ( .B1(n13129), .B2(n12001), .A(n13149), .ZN(n12007) );
  NAND2_X1 U14351 ( .A1(n13144), .A2(n13182), .ZN(n14862) );
  NAND4_X1 U14352 ( .A1(n13129), .A2(n9472), .A3(n12002), .A4(n14849), .ZN(
        n12003) );
  OAI21_X1 U14353 ( .B1(n13147), .B2(n14862), .A(n12003), .ZN(n12004) );
  AOI21_X1 U14354 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n12005), .A(n12004), .ZN(
        n12006) );
  OAI21_X1 U14355 ( .B1(n12007), .B2(n14858), .A(n12006), .ZN(P2_U3204) );
  NAND2_X1 U14356 ( .A1(n12011), .A2(n12010), .ZN(n12012) );
  NAND2_X1 U14357 ( .A1(n14558), .A2(n12118), .ZN(n12014) );
  OR2_X1 U14358 ( .A1(n12016), .A2(n11717), .ZN(n12013) );
  NAND2_X1 U14359 ( .A1(n12014), .A2(n12013), .ZN(n12015) );
  XNOR2_X1 U14360 ( .A(n12015), .B(n12121), .ZN(n12019) );
  NOR2_X1 U14361 ( .A1(n9615), .A2(n12016), .ZN(n12017) );
  AOI21_X1 U14362 ( .B1(n14558), .B2(n12125), .A(n12017), .ZN(n12018) );
  NAND2_X1 U14363 ( .A1(n12019), .A2(n12018), .ZN(n12020) );
  OAI21_X1 U14364 ( .B1(n12019), .B2(n12018), .A(n12020), .ZN(n14546) );
  NAND2_X1 U14365 ( .A1(n13738), .A2(n12118), .ZN(n12022) );
  OR2_X1 U14366 ( .A1(n12024), .A2(n11717), .ZN(n12021) );
  NAND2_X1 U14367 ( .A1(n12022), .A2(n12021), .ZN(n12023) );
  XNOR2_X1 U14368 ( .A(n12023), .B(n12132), .ZN(n12025) );
  OAI22_X1 U14369 ( .A1(n14579), .A2(n11717), .B1(n12024), .B2(n9615), .ZN(
        n13731) );
  INV_X1 U14370 ( .A(n12025), .ZN(n12026) );
  NOR2_X1 U14371 ( .A1(n12027), .A2(n12026), .ZN(n12028) );
  AOI21_X1 U14372 ( .B1(n13732), .B2(n13731), .A(n12028), .ZN(n13652) );
  NAND2_X1 U14373 ( .A1(n14571), .A2(n12118), .ZN(n12030) );
  NAND2_X1 U14374 ( .A1(n12125), .A2(n13757), .ZN(n12029) );
  NAND2_X1 U14375 ( .A1(n12030), .A2(n12029), .ZN(n12031) );
  XNOR2_X1 U14376 ( .A(n12031), .B(n12132), .ZN(n12035) );
  NAND2_X1 U14377 ( .A1(n14571), .A2(n12125), .ZN(n12033) );
  NAND2_X1 U14378 ( .A1(n12068), .A2(n13757), .ZN(n12032) );
  NAND2_X1 U14379 ( .A1(n12033), .A2(n12032), .ZN(n12034) );
  NOR2_X1 U14380 ( .A1(n12035), .A2(n12034), .ZN(n13663) );
  AOI21_X1 U14381 ( .B1(n12035), .B2(n12034), .A(n13663), .ZN(n13653) );
  NAND2_X1 U14382 ( .A1(n13652), .A2(n13653), .ZN(n13661) );
  INV_X1 U14383 ( .A(n13663), .ZN(n12036) );
  NAND2_X1 U14384 ( .A1(n13661), .A2(n12036), .ZN(n12046) );
  NAND2_X1 U14385 ( .A1(n14088), .A2(n12118), .ZN(n12038) );
  NAND2_X1 U14386 ( .A1(n13756), .A2(n12125), .ZN(n12037) );
  NAND2_X1 U14387 ( .A1(n12038), .A2(n12037), .ZN(n12039) );
  XNOR2_X1 U14388 ( .A(n12039), .B(n12121), .ZN(n12041) );
  AND2_X1 U14389 ( .A1(n13756), .A2(n12068), .ZN(n12040) );
  AOI21_X1 U14390 ( .B1(n14088), .B2(n12125), .A(n12040), .ZN(n12042) );
  NAND2_X1 U14391 ( .A1(n12041), .A2(n12042), .ZN(n12047) );
  INV_X1 U14392 ( .A(n12041), .ZN(n12044) );
  INV_X1 U14393 ( .A(n12042), .ZN(n12043) );
  NAND2_X1 U14394 ( .A1(n12044), .A2(n12043), .ZN(n12045) );
  AND2_X1 U14395 ( .A1(n12047), .A2(n12045), .ZN(n13662) );
  NAND2_X1 U14396 ( .A1(n12046), .A2(n13662), .ZN(n13665) );
  NAND2_X1 U14397 ( .A1(n13665), .A2(n12047), .ZN(n13708) );
  OAI22_X1 U14398 ( .A1(n14074), .A2(n11717), .B1(n13668), .B2(n9620), .ZN(
        n12052) );
  OAI22_X1 U14399 ( .A1(n14074), .A2(n12131), .B1(n13668), .B2(n11717), .ZN(
        n12048) );
  XNOR2_X1 U14400 ( .A(n12048), .B(n12132), .ZN(n12051) );
  XOR2_X1 U14401 ( .A(n12052), .B(n12051), .Z(n13709) );
  NAND2_X1 U14402 ( .A1(n13708), .A2(n13709), .ZN(n13707) );
  NOR2_X1 U14403 ( .A1(n13714), .A2(n9615), .ZN(n12049) );
  AOI21_X1 U14404 ( .B1(n13621), .B2(n12125), .A(n12049), .ZN(n12055) );
  AOI22_X1 U14405 ( .A1(n13621), .A2(n12118), .B1(n12125), .B2(n13754), .ZN(
        n12050) );
  XNOR2_X1 U14406 ( .A(n12050), .B(n12132), .ZN(n12056) );
  XOR2_X1 U14407 ( .A(n12055), .B(n12056), .Z(n13624) );
  INV_X1 U14408 ( .A(n12051), .ZN(n12054) );
  INV_X1 U14409 ( .A(n12052), .ZN(n12053) );
  NAND2_X1 U14410 ( .A1(n12054), .A2(n12053), .ZN(n13622) );
  NAND3_X1 U14411 ( .A1(n13707), .A2(n13624), .A3(n13622), .ZN(n13623) );
  OR2_X1 U14412 ( .A1(n12056), .A2(n12055), .ZN(n12057) );
  OAI22_X1 U14413 ( .A1(n14165), .A2(n11717), .B1(n12058), .B2(n9620), .ZN(
        n12062) );
  NAND2_X1 U14414 ( .A1(n14043), .A2(n12118), .ZN(n12060) );
  NAND2_X1 U14415 ( .A1(n13753), .A2(n12125), .ZN(n12059) );
  NAND2_X1 U14416 ( .A1(n12060), .A2(n12059), .ZN(n12061) );
  XNOR2_X1 U14417 ( .A(n12061), .B(n12132), .ZN(n12063) );
  XOR2_X1 U14418 ( .A(n12062), .B(n12063), .Z(n13688) );
  NAND2_X1 U14419 ( .A1(n12063), .A2(n12062), .ZN(n12064) );
  NAND2_X1 U14420 ( .A1(n14220), .A2(n12118), .ZN(n12066) );
  NAND2_X1 U14421 ( .A1(n13752), .A2(n12125), .ZN(n12065) );
  NAND2_X1 U14422 ( .A1(n12066), .A2(n12065), .ZN(n12067) );
  XNOR2_X1 U14423 ( .A(n12067), .B(n12121), .ZN(n12071) );
  AND2_X1 U14424 ( .A1(n13752), .A2(n12068), .ZN(n12069) );
  AOI21_X1 U14425 ( .B1(n14220), .B2(n12125), .A(n12069), .ZN(n12070) );
  NAND2_X1 U14426 ( .A1(n12071), .A2(n12070), .ZN(n13696) );
  OAI21_X1 U14427 ( .B1(n12071), .B2(n12070), .A(n13696), .ZN(n13633) );
  OAI22_X1 U14428 ( .A1(n14217), .A2(n12131), .B1(n13635), .B2(n11717), .ZN(
        n12072) );
  XNOR2_X1 U14429 ( .A(n12072), .B(n12121), .ZN(n12075) );
  INV_X1 U14430 ( .A(n14217), .ZN(n12074) );
  NOR2_X1 U14431 ( .A1(n13635), .A2(n9615), .ZN(n12073) );
  AOI21_X1 U14432 ( .B1(n12074), .B2(n12125), .A(n12073), .ZN(n12076) );
  NAND2_X1 U14433 ( .A1(n12075), .A2(n12076), .ZN(n13611) );
  INV_X1 U14434 ( .A(n12075), .ZN(n12078) );
  INV_X1 U14435 ( .A(n12076), .ZN(n12077) );
  NAND2_X1 U14436 ( .A1(n12078), .A2(n12077), .ZN(n12079) );
  AND2_X1 U14437 ( .A1(n13611), .A2(n12079), .ZN(n13697) );
  NAND2_X1 U14438 ( .A1(n14212), .A2(n12118), .ZN(n12081) );
  NAND2_X1 U14439 ( .A1(n12125), .A2(n13750), .ZN(n12080) );
  NAND2_X1 U14440 ( .A1(n12081), .A2(n12080), .ZN(n12082) );
  XNOR2_X1 U14441 ( .A(n12082), .B(n12121), .ZN(n12086) );
  NOR2_X1 U14442 ( .A1(n9620), .A2(n12083), .ZN(n12084) );
  AOI21_X1 U14443 ( .B1(n14212), .B2(n12125), .A(n12084), .ZN(n12085) );
  NAND2_X1 U14444 ( .A1(n12086), .A2(n12085), .ZN(n13675) );
  OR2_X1 U14445 ( .A1(n12086), .A2(n12085), .ZN(n12087) );
  AND2_X1 U14446 ( .A1(n13675), .A2(n12087), .ZN(n13612) );
  NAND2_X1 U14447 ( .A1(n13613), .A2(n13675), .ZN(n12096) );
  NAND2_X1 U14448 ( .A1(n14132), .A2(n12118), .ZN(n12089) );
  NAND2_X1 U14449 ( .A1(n12125), .A2(n13749), .ZN(n12088) );
  NAND2_X1 U14450 ( .A1(n12089), .A2(n12088), .ZN(n12090) );
  XNOR2_X1 U14451 ( .A(n12090), .B(n12121), .ZN(n12094) );
  NOR2_X1 U14452 ( .A1(n9620), .A2(n12091), .ZN(n12092) );
  AOI21_X1 U14453 ( .B1(n14132), .B2(n12125), .A(n12092), .ZN(n12093) );
  NAND2_X1 U14454 ( .A1(n12094), .A2(n12093), .ZN(n13646) );
  OR2_X1 U14455 ( .A1(n12094), .A2(n12093), .ZN(n12095) );
  AND2_X1 U14456 ( .A1(n13646), .A2(n12095), .ZN(n13676) );
  NAND2_X1 U14457 ( .A1(n13679), .A2(n13646), .ZN(n12105) );
  NAND2_X1 U14458 ( .A1(n13972), .A2(n12118), .ZN(n12098) );
  NAND2_X1 U14459 ( .A1(n12125), .A2(n13748), .ZN(n12097) );
  NAND2_X1 U14460 ( .A1(n12098), .A2(n12097), .ZN(n12099) );
  XNOR2_X1 U14461 ( .A(n12099), .B(n12121), .ZN(n12103) );
  NOR2_X1 U14462 ( .A1(n9620), .A2(n12100), .ZN(n12101) );
  AOI21_X1 U14463 ( .B1(n13972), .B2(n12125), .A(n12101), .ZN(n12102) );
  NAND2_X1 U14464 ( .A1(n12103), .A2(n12102), .ZN(n12106) );
  OR2_X1 U14465 ( .A1(n12103), .A2(n12102), .ZN(n12104) );
  AND2_X1 U14466 ( .A1(n12106), .A2(n12104), .ZN(n13644) );
  NAND2_X1 U14467 ( .A1(n12105), .A2(n13644), .ZN(n13648) );
  NAND2_X1 U14468 ( .A1(n13648), .A2(n12106), .ZN(n13721) );
  NAND2_X1 U14469 ( .A1(n14120), .A2(n12118), .ZN(n12108) );
  NAND2_X1 U14470 ( .A1(n12125), .A2(n13747), .ZN(n12107) );
  NAND2_X1 U14471 ( .A1(n12108), .A2(n12107), .ZN(n12109) );
  XNOR2_X1 U14472 ( .A(n12109), .B(n12121), .ZN(n12113) );
  INV_X1 U14473 ( .A(n12113), .ZN(n12115) );
  NOR2_X1 U14474 ( .A1(n9615), .A2(n12110), .ZN(n12111) );
  AOI21_X1 U14475 ( .B1(n14120), .B2(n12125), .A(n12111), .ZN(n12112) );
  INV_X1 U14476 ( .A(n12112), .ZN(n12114) );
  AND2_X1 U14477 ( .A1(n12113), .A2(n12112), .ZN(n12116) );
  AOI21_X1 U14478 ( .B1(n12115), .B2(n12114), .A(n12116), .ZN(n13722) );
  INV_X1 U14479 ( .A(n12116), .ZN(n12117) );
  NAND2_X1 U14480 ( .A1(n13939), .A2(n12118), .ZN(n12120) );
  NAND2_X1 U14481 ( .A1(n12125), .A2(n13746), .ZN(n12119) );
  NAND2_X1 U14482 ( .A1(n12120), .A2(n12119), .ZN(n12122) );
  XNOR2_X1 U14483 ( .A(n12122), .B(n12121), .ZN(n12127) );
  INV_X1 U14484 ( .A(n12127), .ZN(n12129) );
  NOR2_X1 U14485 ( .A1(n9615), .A2(n12123), .ZN(n12124) );
  AOI21_X1 U14486 ( .B1(n13939), .B2(n12125), .A(n12124), .ZN(n12126) );
  INV_X1 U14487 ( .A(n12126), .ZN(n12128) );
  AND2_X1 U14488 ( .A1(n12127), .A2(n12126), .ZN(n12130) );
  AOI21_X1 U14489 ( .B1(n12129), .B2(n12128), .A(n12130), .ZN(n13604) );
  OAI22_X1 U14490 ( .A1(n14199), .A2(n12131), .B1(n12134), .B2(n11717), .ZN(
        n12133) );
  XNOR2_X1 U14491 ( .A(n12133), .B(n12132), .ZN(n12136) );
  OAI22_X1 U14492 ( .A1(n14199), .A2(n11717), .B1(n12134), .B2(n9615), .ZN(
        n12135) );
  XNOR2_X1 U14493 ( .A(n12136), .B(n12135), .ZN(n12137) );
  OR2_X1 U14494 ( .A1(n12138), .A2(n13713), .ZN(n12140) );
  NAND2_X1 U14495 ( .A1(n13725), .A2(n13746), .ZN(n12139) );
  AND2_X1 U14496 ( .A1(n12140), .A2(n12139), .ZN(n14109) );
  INV_X1 U14497 ( .A(n14109), .ZN(n12141) );
  AOI22_X1 U14498 ( .A1(n14552), .A2(n12141), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12142) );
  OAI21_X1 U14499 ( .B1(n14557), .B2(n13918), .A(n12142), .ZN(n12143) );
  AOI21_X1 U14500 ( .B1(n13915), .B2(n14554), .A(n12143), .ZN(n12144) );
  OAI21_X1 U14501 ( .B1(n12145), .B2(n13740), .A(n12144), .ZN(P1_U3220) );
  INV_X1 U14502 ( .A(n13232), .ZN(n12171) );
  INV_X1 U14503 ( .A(n13283), .ZN(n12168) );
  OR2_X1 U14504 ( .A1(n13520), .A2(n12148), .ZN(n12147) );
  NAND2_X1 U14505 ( .A1(n13520), .A2(n12148), .ZN(n12149) );
  OR2_X1 U14506 ( .A1(n13409), .A2(n13075), .ZN(n12151) );
  INV_X1 U14507 ( .A(n13165), .ZN(n13030) );
  NOR2_X1 U14508 ( .A1(n13507), .A2(n13030), .ZN(n12152) );
  INV_X1 U14509 ( .A(n13507), .ZN(n13394) );
  INV_X1 U14510 ( .A(n13379), .ZN(n13369) );
  INV_X1 U14511 ( .A(n13164), .ZN(n12153) );
  OR2_X1 U14512 ( .A1(n13500), .A2(n12153), .ZN(n12154) );
  NAND2_X1 U14513 ( .A1(n13562), .A2(n13031), .ZN(n12155) );
  INV_X1 U14514 ( .A(n13162), .ZN(n12156) );
  AND2_X1 U14515 ( .A1(n13488), .A2(n12156), .ZN(n12157) );
  NAND2_X1 U14516 ( .A1(n13327), .A2(n13326), .ZN(n12160) );
  OR2_X1 U14517 ( .A1(n13331), .A2(n12158), .ZN(n12159) );
  INV_X1 U14518 ( .A(n13160), .ZN(n12162) );
  NOR2_X1 U14519 ( .A1(n13476), .A2(n12162), .ZN(n12161) );
  NAND2_X1 U14520 ( .A1(n13476), .A2(n12162), .ZN(n12163) );
  INV_X1 U14521 ( .A(n13159), .ZN(n13062) );
  NAND2_X1 U14522 ( .A1(n13470), .A2(n13062), .ZN(n12164) );
  NAND2_X1 U14523 ( .A1(n12165), .A2(n12164), .ZN(n13278) );
  AND2_X1 U14524 ( .A1(n13288), .A2(n12166), .ZN(n12167) );
  AOI21_X1 U14525 ( .B1(n12168), .B2(n13278), .A(n12167), .ZN(n13267) );
  INV_X1 U14526 ( .A(n13157), .ZN(n13063) );
  OR2_X1 U14527 ( .A1(n13543), .A2(n13063), .ZN(n12169) );
  NAND2_X1 U14528 ( .A1(n13448), .A2(n12170), .ZN(n13231) );
  NOR2_X1 U14529 ( .A1(n13589), .A2(n12174), .ZN(n12175) );
  NOR2_X1 U14530 ( .A1(n13074), .A2(n12175), .ZN(n13221) );
  NAND2_X1 U14531 ( .A1(n13221), .A2(n13153), .ZN(n12176) );
  AOI21_X2 U14532 ( .B1(n12178), .B2(n14860), .A(n12177), .ZN(n13440) );
  INV_X1 U14533 ( .A(n13476), .ZN(n13319) );
  INV_X1 U14534 ( .A(n13488), .ZN(n13346) );
  INV_X1 U14535 ( .A(n13409), .ZN(n13512) );
  NAND2_X1 U14536 ( .A1(n13319), .A2(n13330), .ZN(n13315) );
  INV_X1 U14537 ( .A(n13242), .ZN(n12179) );
  AOI22_X1 U14538 ( .A1(n12180), .A2(n14844), .B1(n14873), .B2(
        P2_REG2_REG_29__SCAN_IN), .ZN(n12181) );
  OAI21_X1 U14539 ( .B1(n12182), .B2(n13420), .A(n12181), .ZN(n12209) );
  NAND2_X1 U14540 ( .A1(n12184), .A2(n12183), .ZN(n12186) );
  OR2_X1 U14541 ( .A1(n13525), .A2(n13168), .ZN(n12185) );
  NAND2_X1 U14542 ( .A1(n13500), .A2(n13164), .ZN(n12190) );
  NAND2_X1 U14543 ( .A1(n13380), .A2(n12190), .ZN(n12192) );
  OR2_X1 U14544 ( .A1(n13500), .A2(n13164), .ZN(n12191) );
  NOR2_X1 U14545 ( .A1(n13562), .A2(n13163), .ZN(n12193) );
  NAND2_X1 U14546 ( .A1(n13562), .A2(n13163), .ZN(n12194) );
  INV_X1 U14547 ( .A(n12196), .ZN(n12197) );
  INV_X1 U14548 ( .A(n13326), .ZN(n13324) );
  NAND2_X1 U14549 ( .A1(n13331), .A2(n13161), .ZN(n12198) );
  INV_X1 U14550 ( .A(n12199), .ZN(n12200) );
  NAND2_X1 U14551 ( .A1(n13470), .A2(n13159), .ZN(n12202) );
  OR2_X1 U14552 ( .A1(n13288), .A2(n13158), .ZN(n12204) );
  NAND2_X1 U14553 ( .A1(n13543), .A2(n13157), .ZN(n12205) );
  NAND2_X1 U14554 ( .A1(n13448), .A2(n13156), .ZN(n12206) );
  NAND2_X1 U14555 ( .A1(n13232), .A2(n13230), .ZN(n13229) );
  OAI21_X1 U14556 ( .B1(n13440), .B2(n14873), .A(n12210), .ZN(P2_U3236) );
  INV_X1 U14557 ( .A(n12585), .ZN(n12445) );
  NAND2_X1 U14558 ( .A1(n12212), .A2(n12211), .ZN(n12214) );
  NAND2_X1 U14559 ( .A1(n12460), .A2(n15223), .ZN(n12215) );
  AND2_X1 U14560 ( .A1(n12216), .A2(n12215), .ZN(n15154) );
  NAND2_X1 U14561 ( .A1(n15143), .A2(n12218), .ZN(n12220) );
  INV_X1 U14562 ( .A(n12220), .ZN(n12219) );
  NOR2_X1 U14563 ( .A1(n12219), .A2(n15125), .ZN(n12222) );
  NAND2_X1 U14564 ( .A1(n12458), .A2(n15149), .ZN(n15124) );
  AND2_X1 U14565 ( .A1(n15124), .A2(n12220), .ZN(n12221) );
  OR2_X1 U14566 ( .A1(n12222), .A2(n12221), .ZN(n12223) );
  NAND2_X1 U14567 ( .A1(n12224), .A2(n12223), .ZN(n15108) );
  AND2_X1 U14568 ( .A1(n12457), .A2(n12225), .ZN(n12226) );
  NAND2_X1 U14569 ( .A1(n12456), .A2(n14964), .ZN(n12227) );
  NAND2_X1 U14570 ( .A1(n12797), .A2(n14497), .ZN(n12228) );
  NAND2_X1 U14571 ( .A1(n14492), .A2(n12228), .ZN(n12231) );
  NAND2_X1 U14572 ( .A1(n14956), .A2(n12229), .ZN(n12230) );
  NAND2_X1 U14573 ( .A1(n12795), .A2(n12794), .ZN(n12234) );
  NAND2_X1 U14574 ( .A1(n12455), .A2(n12232), .ZN(n12233) );
  NOR2_X1 U14575 ( .A1(n12785), .A2(n12798), .ZN(n12763) );
  INV_X1 U14576 ( .A(n12781), .ZN(n12274) );
  NAND2_X1 U14577 ( .A1(n12785), .A2(n12798), .ZN(n12764) );
  AND2_X1 U14578 ( .A1(n12773), .A2(n12764), .ZN(n12767) );
  NAND2_X1 U14579 ( .A1(n12875), .A2(n12769), .ZN(n12235) );
  NAND2_X1 U14580 ( .A1(n12738), .A2(n12737), .ZN(n12238) );
  NAND2_X1 U14581 ( .A1(n14434), .A2(n12751), .ZN(n12237) );
  NAND2_X1 U14582 ( .A1(n12238), .A2(n12237), .ZN(n12725) );
  NAND2_X1 U14583 ( .A1(n12725), .A2(n12729), .ZN(n12240) );
  NAND2_X1 U14584 ( .A1(n12867), .A2(n12739), .ZN(n12239) );
  NAND2_X1 U14585 ( .A1(n12240), .A2(n12239), .ZN(n12712) );
  INV_X1 U14586 ( .A(n12712), .ZN(n12241) );
  OR2_X1 U14587 ( .A1(n12407), .A2(n12726), .ZN(n12242) );
  INV_X1 U14588 ( .A(n12453), .ZN(n12716) );
  OR2_X1 U14589 ( .A1(n12931), .A2(n12716), .ZN(n12243) );
  NAND2_X1 U14590 ( .A1(n12694), .A2(n12452), .ZN(n12244) );
  INV_X1 U14591 ( .A(n12685), .ZN(n12451) );
  OR2_X1 U14592 ( .A1(n12677), .A2(n12451), .ZN(n12247) );
  NAND2_X1 U14593 ( .A1(n12664), .A2(n12450), .ZN(n12248) );
  OR2_X1 U14594 ( .A1(n12664), .A2(n12450), .ZN(n12249) );
  NAND2_X1 U14595 ( .A1(n12622), .A2(n12630), .ZN(n12621) );
  INV_X1 U14596 ( .A(n12364), .ZN(n12448) );
  NAND2_X1 U14597 ( .A1(n12909), .A2(n12448), .ZN(n12250) );
  NAND2_X1 U14598 ( .A1(n12621), .A2(n12250), .ZN(n12610) );
  NAND2_X1 U14599 ( .A1(n12610), .A2(n12609), .ZN(n12608) );
  NAND2_X1 U14600 ( .A1(n12829), .A2(n12447), .ZN(n12251) );
  OR2_X1 U14601 ( .A1(n12602), .A2(n12446), .ZN(n12252) );
  NAND2_X1 U14602 ( .A1(n12595), .A2(n12252), .ZN(n12254) );
  NAND2_X1 U14603 ( .A1(n12602), .A2(n12446), .ZN(n12253) );
  OR2_X1 U14604 ( .A1(n12589), .A2(n12571), .ZN(n12255) );
  XNOR2_X1 U14605 ( .A(n12256), .B(n12264), .ZN(n12261) );
  NAND2_X1 U14606 ( .A1(n12257), .A2(P3_B_REG_SCAN_IN), .ZN(n12258) );
  NAND2_X1 U14607 ( .A1(n15142), .A2(n12258), .ZN(n12559) );
  OAI22_X1 U14608 ( .A1(n12585), .A2(n15187), .B1(n12259), .B2(n12559), .ZN(
        n12260) );
  INV_X1 U14609 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12263) );
  NAND2_X1 U14610 ( .A1(n12262), .A2(n15203), .ZN(n12561) );
  OAI21_X1 U14611 ( .B1(n15204), .B2(n12263), .A(n12561), .ZN(n12265) );
  NAND2_X1 U14612 ( .A1(n15169), .A2(n15200), .ZN(n15148) );
  XNOR2_X1 U14613 ( .A(n12589), .B(n12328), .ZN(n12326) );
  XNOR2_X1 U14614 ( .A(n12326), .B(n12571), .ZN(n12327) );
  NAND2_X1 U14615 ( .A1(n12268), .A2(n14496), .ZN(n12266) );
  INV_X1 U14616 ( .A(n12268), .ZN(n12269) );
  NAND2_X1 U14617 ( .A1(n12455), .A2(n12269), .ZN(n12270) );
  XNOR2_X1 U14618 ( .A(n12785), .B(n12296), .ZN(n12272) );
  NAND2_X1 U14619 ( .A1(n12272), .A2(n12798), .ZN(n12390) );
  INV_X1 U14620 ( .A(n12272), .ZN(n12273) );
  NAND2_X1 U14621 ( .A1(n12273), .A2(n12454), .ZN(n12391) );
  XNOR2_X1 U14622 ( .A(n14424), .B(n12328), .ZN(n12275) );
  XNOR2_X1 U14623 ( .A(n12275), .B(n12274), .ZN(n14418) );
  NAND2_X1 U14624 ( .A1(n12275), .A2(n12781), .ZN(n12276) );
  XNOR2_X1 U14625 ( .A(n12875), .B(n12328), .ZN(n12277) );
  XNOR2_X1 U14626 ( .A(n12277), .B(n12769), .ZN(n12435) );
  NAND2_X1 U14627 ( .A1(n12436), .A2(n12435), .ZN(n12434) );
  INV_X1 U14628 ( .A(n12277), .ZN(n12278) );
  NAND2_X1 U14629 ( .A1(n12278), .A2(n12769), .ZN(n12279) );
  NAND2_X1 U14630 ( .A1(n12434), .A2(n12279), .ZN(n14430) );
  XNOR2_X1 U14631 ( .A(n14434), .B(n12328), .ZN(n12281) );
  XNOR2_X1 U14632 ( .A(n12281), .B(n12439), .ZN(n14429) );
  NAND2_X1 U14633 ( .A1(n12281), .A2(n12439), .ZN(n12282) );
  XNOR2_X1 U14634 ( .A(n12867), .B(n12328), .ZN(n12283) );
  XNOR2_X1 U14635 ( .A(n12283), .B(n12715), .ZN(n12354) );
  XNOR2_X1 U14636 ( .A(n12407), .B(n12328), .ZN(n12286) );
  XNOR2_X1 U14637 ( .A(n12286), .B(n12726), .ZN(n12411) );
  INV_X1 U14638 ( .A(n12411), .ZN(n12285) );
  INV_X1 U14639 ( .A(n12283), .ZN(n12284) );
  NAND2_X1 U14640 ( .A1(n12284), .A2(n12739), .ZN(n12408) );
  INV_X1 U14641 ( .A(n12286), .ZN(n12287) );
  NAND2_X1 U14642 ( .A1(n12287), .A2(n12726), .ZN(n12288) );
  XNOR2_X1 U14643 ( .A(n12931), .B(n12328), .ZN(n12289) );
  XNOR2_X1 U14644 ( .A(n12289), .B(n12716), .ZN(n12319) );
  NAND2_X1 U14645 ( .A1(n12320), .A2(n12319), .ZN(n12318) );
  NAND2_X1 U14646 ( .A1(n12289), .A2(n12453), .ZN(n12290) );
  NAND2_X1 U14647 ( .A1(n12318), .A2(n12290), .ZN(n12385) );
  XNOR2_X1 U14648 ( .A(n12694), .B(n12328), .ZN(n12291) );
  XNOR2_X1 U14649 ( .A(n12291), .B(n12452), .ZN(n12384) );
  INV_X1 U14650 ( .A(n12291), .ZN(n12292) );
  NAND2_X1 U14651 ( .A1(n12292), .A2(n12452), .ZN(n12293) );
  XNOR2_X1 U14652 ( .A(n12677), .B(n12328), .ZN(n12294) );
  XNOR2_X1 U14653 ( .A(n12294), .B(n12685), .ZN(n12340) );
  NAND2_X1 U14654 ( .A1(n12294), .A2(n12685), .ZN(n12295) );
  XNOR2_X1 U14655 ( .A(n12664), .B(n12296), .ZN(n12297) );
  INV_X1 U14656 ( .A(n12297), .ZN(n12298) );
  AND2_X1 U14657 ( .A1(n12299), .A2(n12298), .ZN(n12300) );
  AOI21_X2 U14658 ( .B1(n12400), .B2(n12676), .A(n12300), .ZN(n12362) );
  XNOR2_X1 U14659 ( .A(n12909), .B(n12328), .ZN(n12365) );
  XNOR2_X1 U14660 ( .A(n12654), .B(n12328), .ZN(n12302) );
  OAI22_X1 U14661 ( .A1(n12365), .A2(n12364), .B1(n12401), .B2(n12302), .ZN(
        n12305) );
  INV_X1 U14662 ( .A(n12302), .ZN(n12361) );
  OAI21_X1 U14663 ( .B1(n12361), .B2(n12449), .A(n12448), .ZN(n12301) );
  NAND2_X1 U14664 ( .A1(n12365), .A2(n12301), .ZN(n12304) );
  NAND3_X1 U14665 ( .A1(n12302), .A2(n12401), .A3(n12364), .ZN(n12303) );
  OAI211_X2 U14666 ( .C1(n12362), .C2(n12305), .A(n12304), .B(n12303), .ZN(
        n12346) );
  XNOR2_X1 U14667 ( .A(n12829), .B(n12328), .ZN(n12306) );
  XNOR2_X1 U14668 ( .A(n12306), .B(n12447), .ZN(n12347) );
  XNOR2_X1 U14669 ( .A(n12602), .B(n12328), .ZN(n12307) );
  XNOR2_X1 U14670 ( .A(n12307), .B(n12584), .ZN(n12428) );
  AOI22_X1 U14671 ( .A1(n12446), .A2(n12437), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12309) );
  NAND2_X1 U14672 ( .A1(n12590), .A2(n14436), .ZN(n12308) );
  OAI211_X1 U14673 ( .C1(n12585), .C2(n12440), .A(n12309), .B(n12308), .ZN(
        n12310) );
  AOI21_X1 U14674 ( .B1(n12589), .B2(n14965), .A(n12310), .ZN(n12311) );
  OAI21_X1 U14675 ( .B1(n12312), .B2(n12433), .A(n12311), .ZN(P3_U3154) );
  XNOR2_X1 U14676 ( .A(n12362), .B(n12361), .ZN(n12363) );
  XNOR2_X1 U14677 ( .A(n12363), .B(n12401), .ZN(n12317) );
  INV_X1 U14678 ( .A(n12313), .ZN(n12651) );
  OAI22_X1 U14679 ( .A1(n12364), .A2(n15185), .B1(n12676), .B2(n15187), .ZN(
        n12648) );
  AOI22_X1 U14680 ( .A1(n12648), .A2(n14420), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12314) );
  OAI21_X1 U14681 ( .B1(n12651), .B2(n14971), .A(n12314), .ZN(n12315) );
  AOI21_X1 U14682 ( .B1(n12654), .B2(n14965), .A(n12315), .ZN(n12316) );
  OAI21_X1 U14683 ( .B1(n12317), .B2(n12433), .A(n12316), .ZN(P3_U3156) );
  OAI211_X1 U14684 ( .C1(n12320), .C2(n12319), .A(n12318), .B(n14960), .ZN(
        n12325) );
  AND2_X1 U14685 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12551) );
  AOI21_X1 U14686 ( .B1(n12452), .B2(n12422), .A(n12551), .ZN(n12321) );
  OAI21_X1 U14687 ( .B1(n12322), .B2(n12414), .A(n12321), .ZN(n12323) );
  AOI21_X1 U14688 ( .B1(n12705), .B2(n14436), .A(n12323), .ZN(n12324) );
  OAI211_X1 U14689 ( .C1(n14425), .C2(n12931), .A(n12325), .B(n12324), .ZN(
        P3_U3159) );
  XOR2_X1 U14690 ( .A(n12328), .B(n12565), .Z(n12329) );
  NAND2_X1 U14691 ( .A1(n12330), .A2(n14960), .ZN(n12336) );
  INV_X1 U14692 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n12331) );
  OAI22_X1 U14693 ( .A1(n12598), .A2(n12414), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12331), .ZN(n12332) );
  INV_X1 U14694 ( .A(n12332), .ZN(n12335) );
  AOI22_X1 U14695 ( .A1(n12570), .A2(n12422), .B1(n12577), .B2(n14436), .ZN(
        n12334) );
  NAND2_X1 U14696 ( .A1(n6693), .A2(n14965), .ZN(n12333) );
  NAND4_X1 U14697 ( .A1(n12336), .A2(n12335), .A3(n12334), .A4(n12333), .ZN(
        P3_U3160) );
  INV_X1 U14698 ( .A(n12337), .ZN(n12338) );
  AOI21_X1 U14699 ( .B1(n12340), .B2(n12339), .A(n12338), .ZN(n12345) );
  AOI22_X1 U14700 ( .A1(n12422), .A2(n12450), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12342) );
  NAND2_X1 U14701 ( .A1(n14436), .A2(n12678), .ZN(n12341) );
  OAI211_X1 U14702 ( .C1(n12704), .C2(n12414), .A(n12342), .B(n12341), .ZN(
        n12343) );
  AOI21_X1 U14703 ( .B1(n12677), .B2(n14965), .A(n12343), .ZN(n12344) );
  OAI21_X1 U14704 ( .B1(n12345), .B2(n12433), .A(n12344), .ZN(P3_U3163) );
  XOR2_X1 U14705 ( .A(n12347), .B(n12346), .Z(n12353) );
  NAND2_X1 U14706 ( .A1(n12446), .A2(n15142), .ZN(n12349) );
  OR2_X1 U14707 ( .A1(n12364), .A2(n15187), .ZN(n12348) );
  AND2_X1 U14708 ( .A1(n12349), .A2(n12348), .ZN(n12611) );
  AOI22_X1 U14709 ( .A1(n12616), .A2(n14436), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12350) );
  OAI21_X1 U14710 ( .B1(n12611), .B2(n14968), .A(n12350), .ZN(n12351) );
  AOI21_X1 U14711 ( .B1(n12829), .B2(n14965), .A(n12351), .ZN(n12352) );
  OAI21_X1 U14712 ( .B1(n12353), .B2(n12433), .A(n12352), .ZN(P3_U3165) );
  AOI21_X1 U14713 ( .B1(n12355), .B2(n12354), .A(n12433), .ZN(n12356) );
  OR2_X1 U14714 ( .A1(n12355), .A2(n12354), .ZN(n12409) );
  NAND2_X1 U14715 ( .A1(n12356), .A2(n12409), .ZN(n12360) );
  AOI22_X1 U14716 ( .A1(n12726), .A2(n12422), .B1(P3_REG3_REG_17__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12357) );
  OAI21_X1 U14717 ( .B1(n12439), .B2(n12414), .A(n12357), .ZN(n12358) );
  AOI21_X1 U14718 ( .B1(n12732), .B2(n14436), .A(n12358), .ZN(n12359) );
  OAI211_X1 U14719 ( .C1(n12734), .C2(n14425), .A(n12360), .B(n12359), .ZN(
        P3_U3168) );
  OAI22_X1 U14720 ( .A1(n12363), .A2(n12449), .B1(n12362), .B2(n12361), .ZN(
        n12367) );
  XNOR2_X1 U14721 ( .A(n12365), .B(n12364), .ZN(n12366) );
  XNOR2_X1 U14722 ( .A(n12367), .B(n12366), .ZN(n12374) );
  INV_X1 U14723 ( .A(n12634), .ZN(n12371) );
  OR2_X1 U14724 ( .A1(n12597), .A2(n15185), .ZN(n12369) );
  NAND2_X1 U14725 ( .A1(n12449), .A2(n15145), .ZN(n12368) );
  NAND2_X1 U14726 ( .A1(n12369), .A2(n12368), .ZN(n12623) );
  AOI22_X1 U14727 ( .A1(n12623), .A2(n14420), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12370) );
  OAI21_X1 U14728 ( .B1(n12371), .B2(n14971), .A(n12370), .ZN(n12372) );
  AOI21_X1 U14729 ( .B1(n12909), .B2(n14965), .A(n12372), .ZN(n12373) );
  OAI21_X1 U14730 ( .B1(n12374), .B2(n12433), .A(n12373), .ZN(P3_U3169) );
  NAND2_X1 U14731 ( .A1(n12376), .A2(n12375), .ZN(n12377) );
  AOI21_X1 U14732 ( .B1(n14958), .B2(n12377), .A(n12433), .ZN(n12382) );
  AOI22_X1 U14733 ( .A1(n12456), .A2(n15142), .B1(n15145), .B2(n12457), .ZN(
        n15090) );
  AOI22_X1 U14734 ( .A1(n14965), .A2(n15241), .B1(P3_REG3_REG_9__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12380) );
  NAND2_X1 U14735 ( .A1(n14436), .A2(n12378), .ZN(n12379) );
  OAI211_X1 U14736 ( .C1(n15090), .C2(n14968), .A(n12380), .B(n12379), .ZN(
        n12381) );
  OR2_X1 U14737 ( .A1(n12382), .A2(n12381), .ZN(P3_U3171) );
  OAI211_X1 U14738 ( .C1(n12385), .C2(n12384), .A(n12383), .B(n14960), .ZN(
        n12389) );
  AOI22_X1 U14739 ( .A1(n12451), .A2(n12422), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12386) );
  OAI21_X1 U14740 ( .B1(n12716), .B2(n12414), .A(n12386), .ZN(n12387) );
  AOI21_X1 U14741 ( .B1(n12686), .B2(n14436), .A(n12387), .ZN(n12388) );
  OAI211_X1 U14742 ( .C1(n12927), .C2(n14425), .A(n12389), .B(n12388), .ZN(
        P3_U3173) );
  NAND2_X1 U14743 ( .A1(n12391), .A2(n12390), .ZN(n12393) );
  XOR2_X1 U14744 ( .A(n12393), .B(n12392), .Z(n12399) );
  NAND2_X1 U14745 ( .A1(n12422), .A2(n12781), .ZN(n12395) );
  OAI211_X1 U14746 ( .C1(n14496), .C2(n12414), .A(n12395), .B(n12394), .ZN(
        n12397) );
  NOR2_X1 U14747 ( .A1(n12785), .A2(n14425), .ZN(n12396) );
  AOI211_X1 U14748 ( .C1(n12786), .C2(n14436), .A(n12397), .B(n12396), .ZN(
        n12398) );
  OAI21_X1 U14749 ( .B1(n12399), .B2(n12433), .A(n12398), .ZN(P3_U3174) );
  XNOR2_X1 U14750 ( .A(n12400), .B(n12450), .ZN(n12406) );
  INV_X1 U14751 ( .A(n12665), .ZN(n12403) );
  OAI22_X1 U14752 ( .A1(n12401), .A2(n15185), .B1(n12685), .B2(n15187), .ZN(
        n12660) );
  AOI22_X1 U14753 ( .A1(n12660), .A2(n14420), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12402) );
  OAI21_X1 U14754 ( .B1(n12403), .B2(n14971), .A(n12402), .ZN(n12404) );
  AOI21_X1 U14755 ( .B1(n12664), .B2(n14965), .A(n12404), .ZN(n12405) );
  OAI21_X1 U14756 ( .B1(n12406), .B2(n12433), .A(n12405), .ZN(P3_U3175) );
  INV_X1 U14757 ( .A(n12407), .ZN(n12935) );
  NAND2_X1 U14758 ( .A1(n12409), .A2(n12408), .ZN(n12412) );
  OAI211_X1 U14759 ( .C1(n12412), .C2(n12411), .A(n12410), .B(n14960), .ZN(
        n12417) );
  AOI22_X1 U14760 ( .A1(n12422), .A2(n12453), .B1(P3_REG3_REG_18__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12413) );
  OAI21_X1 U14761 ( .B1(n12715), .B2(n12414), .A(n12413), .ZN(n12415) );
  AOI21_X1 U14762 ( .B1(n12719), .B2(n14436), .A(n12415), .ZN(n12416) );
  OAI211_X1 U14763 ( .C1(n12935), .C2(n14425), .A(n12417), .B(n12416), .ZN(
        P3_U3178) );
  AOI21_X1 U14764 ( .B1(n12418), .B2(n12419), .A(n12433), .ZN(n12421) );
  NAND2_X1 U14765 ( .A1(n12421), .A2(n12420), .ZN(n12426) );
  AOI22_X1 U14766 ( .A1(n14965), .A2(n15149), .B1(P3_REG3_REG_6__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12425) );
  AOI22_X1 U14767 ( .A1(n12437), .A2(n15144), .B1(n15143), .B2(n12422), .ZN(
        n12424) );
  NAND2_X1 U14768 ( .A1(n14436), .A2(n15150), .ZN(n12423) );
  NAND4_X1 U14769 ( .A1(n12426), .A2(n12425), .A3(n12424), .A4(n12423), .ZN(
        P3_U3179) );
  AOI22_X1 U14770 ( .A1(n12447), .A2(n12437), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12430) );
  NAND2_X1 U14771 ( .A1(n12603), .A2(n14436), .ZN(n12429) );
  OAI211_X1 U14772 ( .C1(n12598), .C2(n12440), .A(n12430), .B(n12429), .ZN(
        n12431) );
  AOI21_X1 U14773 ( .B1(n12602), .B2(n14965), .A(n12431), .ZN(n12432) );
  OAI211_X1 U14774 ( .C1(n12436), .C2(n12435), .A(n12434), .B(n14960), .ZN(
        n12443) );
  NAND2_X1 U14775 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(P3_U3151), .ZN(n12500)
         );
  NAND2_X1 U14776 ( .A1(n12437), .A2(n12781), .ZN(n12438) );
  OAI211_X1 U14777 ( .C1(n12440), .C2(n12439), .A(n12500), .B(n12438), .ZN(
        n12441) );
  AOI21_X1 U14778 ( .B1(n12758), .B2(n14436), .A(n12441), .ZN(n12442) );
  OAI211_X1 U14779 ( .C1(n12760), .C2(n14425), .A(n12443), .B(n12442), .ZN(
        P3_U3181) );
  MUX2_X1 U14780 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12444), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14781 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12570), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U14782 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12445), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14783 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12571), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14784 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12446), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14785 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12447), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14786 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12448), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14787 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12449), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14788 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12450), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14789 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12451), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14790 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12452), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14791 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12453), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14792 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12726), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14793 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12739), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14794 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12751), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14795 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12769), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14796 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12781), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14797 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12454), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14798 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12455), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14799 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12456), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14800 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n14955), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14801 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12457), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14802 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n15143), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14803 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12458), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14804 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n15144), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14805 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12460), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14806 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12461), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14807 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12462), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14808 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n12463), .S(P3_U3897), .Z(
        P3_U3492) );
  NOR2_X1 U14809 ( .A1(n12480), .A2(n12464), .ZN(n12466) );
  NAND2_X1 U14810 ( .A1(n12494), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12503) );
  OAI21_X1 U14811 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n12494), .A(n12503), 
        .ZN(n12467) );
  AOI21_X1 U14812 ( .B1(n6585), .B2(n12467), .A(n12493), .ZN(n12492) );
  NAND2_X1 U14813 ( .A1(n12469), .A2(n12468), .ZN(n12471) );
  NAND2_X1 U14814 ( .A1(n12494), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12502) );
  OR2_X1 U14815 ( .A1(n12494), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12472) );
  AND2_X1 U14816 ( .A1(n12502), .A2(n12472), .ZN(n12483) );
  NAND2_X1 U14817 ( .A1(n12483), .A2(n12473), .ZN(n12497) );
  OAI21_X1 U14818 ( .B1(n12473), .B2(n12483), .A(n12497), .ZN(n12478) );
  INV_X1 U14819 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n12474) );
  NOR2_X1 U14820 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12474), .ZN(n12475) );
  AOI21_X1 U14821 ( .B1(n15025), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12475), 
        .ZN(n12476) );
  OAI21_X1 U14822 ( .B1(n15020), .B2(n12494), .A(n12476), .ZN(n12477) );
  AOI21_X1 U14823 ( .B1(n12478), .B2(n15058), .A(n12477), .ZN(n12491) );
  INV_X1 U14824 ( .A(n12479), .ZN(n12481) );
  NAND2_X1 U14825 ( .A1(n12481), .A2(n12480), .ZN(n12485) );
  AND2_X1 U14826 ( .A1(n12487), .A2(n12485), .ZN(n12489) );
  OR2_X1 U14827 ( .A1(n12494), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12482) );
  AND2_X1 U14828 ( .A1(n12503), .A2(n12482), .ZN(n12484) );
  MUX2_X1 U14829 ( .A(n12484), .B(n12483), .S(n12516), .Z(n12488) );
  AND2_X1 U14830 ( .A1(n12485), .A2(n12488), .ZN(n12486) );
  NAND2_X1 U14831 ( .A1(n12487), .A2(n12486), .ZN(n12505) );
  OAI211_X1 U14832 ( .C1(n12489), .C2(n12488), .A(n14478), .B(n12505), .ZN(
        n12490) );
  OAI211_X1 U14833 ( .C1(n12492), .C2(n15061), .A(n12491), .B(n12490), .ZN(
        P3_U3196) );
  AOI21_X1 U14834 ( .B1(n12496), .B2(n12495), .A(n12529), .ZN(n12512) );
  INV_X1 U14835 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14349) );
  NAND2_X1 U14836 ( .A1(n12502), .A2(n12497), .ZN(n12539) );
  XNOR2_X1 U14837 ( .A(n12528), .B(n12539), .ZN(n12498) );
  NAND2_X1 U14838 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12498), .ZN(n12541) );
  OAI21_X1 U14839 ( .B1(n12498), .B2(P3_REG1_REG_15__SCAN_IN), .A(n12541), 
        .ZN(n12499) );
  NAND2_X1 U14840 ( .A1(n15058), .A2(n12499), .ZN(n12501) );
  OAI211_X1 U14841 ( .C1(n14349), .C2(n15074), .A(n12501), .B(n12500), .ZN(
        n12510) );
  MUX2_X1 U14842 ( .A(n12503), .B(n12502), .S(n12516), .Z(n12504) );
  NAND2_X1 U14843 ( .A1(n12505), .A2(n12504), .ZN(n12513) );
  XNOR2_X1 U14844 ( .A(n12513), .B(n12540), .ZN(n12507) );
  MUX2_X1 U14845 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12516), .Z(n12506) );
  OR2_X1 U14846 ( .A1(n12507), .A2(n12506), .ZN(n12515) );
  NAND2_X1 U14847 ( .A1(n12507), .A2(n12506), .ZN(n12508) );
  AOI21_X1 U14848 ( .B1(n12515), .B2(n12508), .A(n15067), .ZN(n12509) );
  AOI211_X1 U14849 ( .C1(n15056), .C2(n12528), .A(n12510), .B(n12509), .ZN(
        n12511) );
  OAI21_X1 U14850 ( .B1(n12512), .B2(n15061), .A(n12511), .ZN(P3_U3197) );
  OR2_X1 U14851 ( .A1(n12513), .A2(n12540), .ZN(n12514) );
  NAND2_X1 U14852 ( .A1(n12515), .A2(n12514), .ZN(n14445) );
  MUX2_X1 U14853 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12516), .Z(n12517) );
  NAND2_X1 U14854 ( .A1(n12517), .A2(n12538), .ZN(n14443) );
  NAND2_X1 U14855 ( .A1(n14445), .A2(n14443), .ZN(n12519) );
  INV_X1 U14856 ( .A(n12517), .ZN(n12518) );
  NAND2_X1 U14857 ( .A1(n12518), .A2(n14439), .ZN(n14444) );
  NAND2_X1 U14858 ( .A1(n12519), .A2(n14444), .ZN(n14460) );
  MUX2_X1 U14859 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12516), .Z(n12520) );
  XNOR2_X1 U14860 ( .A(n12520), .B(n12543), .ZN(n14459) );
  NAND2_X1 U14861 ( .A1(n12520), .A2(n12543), .ZN(n12521) );
  NAND2_X1 U14862 ( .A1(n14461), .A2(n12521), .ZN(n12522) );
  XNOR2_X1 U14863 ( .A(n12522), .B(n14470), .ZN(n14476) );
  INV_X1 U14864 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12865) );
  MUX2_X1 U14865 ( .A(n12534), .B(n12865), .S(n12516), .Z(n14475) );
  NAND2_X1 U14866 ( .A1(n14476), .A2(n14475), .ZN(n14474) );
  OAI21_X1 U14867 ( .B1(n12522), .B2(n12546), .A(n14474), .ZN(n12526) );
  XNOR2_X1 U14868 ( .A(n12523), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12535) );
  INV_X1 U14869 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12861) );
  XNOR2_X1 U14870 ( .A(n12523), .B(n12861), .ZN(n12548) );
  INV_X1 U14871 ( .A(n12548), .ZN(n12524) );
  MUX2_X1 U14872 ( .A(n12535), .B(n12524), .S(n9654), .Z(n12525) );
  XNOR2_X1 U14873 ( .A(n12526), .B(n12525), .ZN(n12557) );
  NOR2_X1 U14874 ( .A1(n12528), .A2(n12527), .ZN(n12530) );
  AOI22_X1 U14875 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n14439), .B1(n12538), 
        .B2(n12531), .ZN(n14449) );
  NOR2_X1 U14876 ( .A1(n14456), .A2(n12532), .ZN(n12533) );
  XNOR2_X1 U14877 ( .A(n12536), .B(n12535), .ZN(n12537) );
  AOI22_X1 U14878 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n12546), .B1(n14470), 
        .B2(n12865), .ZN(n14473) );
  INV_X1 U14879 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12873) );
  AOI22_X1 U14880 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12538), .B1(n14439), 
        .B2(n12873), .ZN(n14442) );
  NAND2_X1 U14881 ( .A1(n12540), .A2(n12539), .ZN(n12542) );
  NAND2_X1 U14882 ( .A1(n12542), .A2(n12541), .ZN(n14441) );
  NAND2_X1 U14883 ( .A1(n14442), .A2(n14441), .ZN(n14440) );
  NAND2_X1 U14884 ( .A1(n12543), .A2(n12544), .ZN(n12545) );
  XNOR2_X1 U14885 ( .A(n14456), .B(n12544), .ZN(n14458) );
  NAND2_X1 U14886 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14458), .ZN(n14457) );
  NAND2_X1 U14887 ( .A1(n12545), .A2(n14457), .ZN(n14472) );
  NAND2_X1 U14888 ( .A1(n14473), .A2(n14472), .ZN(n14471) );
  NAND2_X1 U14889 ( .A1(n12546), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12547) );
  NAND2_X1 U14890 ( .A1(n14471), .A2(n12547), .ZN(n12549) );
  XNOR2_X1 U14891 ( .A(n12549), .B(n12548), .ZN(n12555) );
  NAND2_X1 U14892 ( .A1(n15056), .A2(n12550), .ZN(n12553) );
  AOI21_X1 U14893 ( .B1(n15025), .B2(P3_ADDR_REG_19__SCAN_IN), .A(n12551), 
        .ZN(n12552) );
  NAND2_X1 U14894 ( .A1(n12553), .A2(n12552), .ZN(n12554) );
  AOI21_X1 U14895 ( .B1(n12555), .B2(n15058), .A(n12554), .ZN(n12556) );
  OR2_X1 U14896 ( .A1(n12560), .A2(n12559), .ZN(n12885) );
  OAI21_X1 U14897 ( .B1(n12885), .B2(n15177), .A(n12561), .ZN(n12563) );
  AOI21_X1 U14898 ( .B1(P3_REG2_REG_31__SCAN_IN), .B2(n15177), .A(n12563), 
        .ZN(n12562) );
  OAI21_X1 U14899 ( .B1(n12887), .B2(n15100), .A(n12562), .ZN(P3_U3202) );
  AOI21_X1 U14900 ( .B1(P3_REG2_REG_30__SCAN_IN), .B2(n15177), .A(n12563), 
        .ZN(n12564) );
  OAI21_X1 U14901 ( .B1(n12890), .B2(n15100), .A(n12564), .ZN(P3_U3203) );
  NAND2_X1 U14902 ( .A1(n12566), .A2(n12565), .ZN(n12567) );
  NAND2_X1 U14903 ( .A1(n12567), .A2(n15183), .ZN(n12568) );
  OR2_X1 U14904 ( .A1(n12569), .A2(n12568), .ZN(n12573) );
  AOI22_X1 U14905 ( .A1(n12571), .A2(n15145), .B1(n12570), .B2(n15142), .ZN(
        n12572) );
  NAND2_X1 U14906 ( .A1(n12573), .A2(n12572), .ZN(n12819) );
  INV_X1 U14907 ( .A(n12819), .ZN(n12581) );
  XNOR2_X1 U14908 ( .A(n12575), .B(n12574), .ZN(n12817) );
  AOI22_X1 U14909 ( .A1(n12577), .A2(n15203), .B1(n15177), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12578) );
  OAI21_X1 U14910 ( .B1(n12897), .B2(n15100), .A(n12578), .ZN(n12579) );
  AOI21_X1 U14911 ( .B1(n12817), .B2(n15086), .A(n12579), .ZN(n12580) );
  OAI21_X1 U14912 ( .B1(n12581), .B2(n15177), .A(n12580), .ZN(P3_U3205) );
  INV_X1 U14913 ( .A(n12821), .ZN(n12594) );
  OAI21_X1 U14914 ( .B1(n12588), .B2(n12587), .A(n12586), .ZN(n12822) );
  AOI22_X1 U14915 ( .A1(n12590), .A2(n15203), .B1(n15177), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12591) );
  OAI21_X1 U14916 ( .B1(n12901), .B2(n15100), .A(n12591), .ZN(n12592) );
  AOI21_X1 U14917 ( .B1(n12822), .B2(n15086), .A(n12592), .ZN(n12593) );
  OAI21_X1 U14918 ( .B1(n12594), .B2(n15177), .A(n12593), .ZN(P3_U3206) );
  XOR2_X1 U14919 ( .A(n12595), .B(n12600), .Z(n12596) );
  OAI222_X1 U14920 ( .A1(n15185), .A2(n12598), .B1(n15187), .B2(n12597), .C1(
        n12596), .C2(n15130), .ZN(n12825) );
  INV_X1 U14921 ( .A(n12825), .ZN(n12607) );
  NAND2_X1 U14922 ( .A1(n12613), .A2(n12599), .ZN(n12601) );
  XNOR2_X1 U14923 ( .A(n12601), .B(n12600), .ZN(n12826) );
  AOI22_X1 U14924 ( .A1(n12603), .A2(n15203), .B1(n15177), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12604) );
  OAI21_X1 U14925 ( .B1(n12905), .B2(n15100), .A(n12604), .ZN(n12605) );
  AOI21_X1 U14926 ( .B1(n12826), .B2(n15086), .A(n12605), .ZN(n12606) );
  OAI21_X1 U14927 ( .B1(n12607), .B2(n15177), .A(n12606), .ZN(P3_U3207) );
  OAI211_X1 U14928 ( .C1(n12610), .C2(n12609), .A(n12608), .B(n15183), .ZN(
        n12612) );
  OAI21_X1 U14929 ( .B1(n12615), .B2(n12614), .A(n12613), .ZN(n12830) );
  INV_X1 U14930 ( .A(n12829), .ZN(n12618) );
  AOI22_X1 U14931 ( .A1(n12616), .A2(n15203), .B1(n15177), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12617) );
  OAI21_X1 U14932 ( .B1(n12618), .B2(n15100), .A(n12617), .ZN(n12619) );
  AOI21_X1 U14933 ( .B1(n12830), .B2(n15086), .A(n12619), .ZN(n12620) );
  OAI21_X1 U14934 ( .B1(n12832), .B2(n15177), .A(n12620), .ZN(P3_U3208) );
  OAI211_X1 U14935 ( .C1(n12622), .C2(n12630), .A(n12621), .B(n15183), .ZN(
        n12625) );
  INV_X1 U14936 ( .A(n12623), .ZN(n12624) );
  AND2_X1 U14937 ( .A1(n12627), .A2(n12626), .ZN(n12646) );
  INV_X1 U14938 ( .A(n12628), .ZN(n12629) );
  NAND2_X1 U14939 ( .A1(n12646), .A2(n12629), .ZN(n12631) );
  NAND2_X1 U14940 ( .A1(n12631), .A2(n12630), .ZN(n12633) );
  NAND2_X1 U14941 ( .A1(n12633), .A2(n12632), .ZN(n12833) );
  INV_X1 U14942 ( .A(n12909), .ZN(n12636) );
  AOI22_X1 U14943 ( .A1(n15177), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n12634), 
        .B2(n15203), .ZN(n12635) );
  OAI21_X1 U14944 ( .B1(n12636), .B2(n15100), .A(n12635), .ZN(n12637) );
  AOI21_X1 U14945 ( .B1(n12833), .B2(n15086), .A(n12637), .ZN(n12638) );
  OAI21_X1 U14946 ( .B1(n12835), .B2(n15177), .A(n12638), .ZN(P3_U3209) );
  NAND2_X1 U14947 ( .A1(n12639), .A2(n12640), .ZN(n12642) );
  NAND2_X1 U14948 ( .A1(n12642), .A2(n12641), .ZN(n12644) );
  OR2_X1 U14949 ( .A1(n12644), .A2(n12643), .ZN(n12645) );
  NAND2_X1 U14950 ( .A1(n12646), .A2(n12645), .ZN(n12839) );
  OAI211_X1 U14951 ( .C1(n6551), .C2(n7401), .A(n12647), .B(n15183), .ZN(
        n12650) );
  INV_X1 U14952 ( .A(n12648), .ZN(n12649) );
  OAI211_X1 U14953 ( .C1(n15169), .C2(n12839), .A(n12650), .B(n12649), .ZN(
        n12840) );
  NAND2_X1 U14954 ( .A1(n12840), .A2(n15204), .ZN(n12656) );
  INV_X1 U14955 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12652) );
  OAI22_X1 U14956 ( .A1(n15204), .A2(n12652), .B1(n12651), .B2(n15104), .ZN(
        n12653) );
  AOI21_X1 U14957 ( .B1(n12654), .B2(n12695), .A(n12653), .ZN(n12655) );
  OAI211_X1 U14958 ( .C1(n12839), .C2(n12657), .A(n12656), .B(n12655), .ZN(
        P3_U3210) );
  XNOR2_X1 U14959 ( .A(n12659), .B(n12658), .ZN(n12662) );
  INV_X1 U14960 ( .A(n12660), .ZN(n12661) );
  OAI21_X1 U14961 ( .B1(n12662), .B2(n15130), .A(n12661), .ZN(n12844) );
  INV_X1 U14962 ( .A(n12844), .ZN(n12669) );
  XNOR2_X1 U14963 ( .A(n12639), .B(n12663), .ZN(n12845) );
  INV_X1 U14964 ( .A(n12664), .ZN(n12919) );
  AOI22_X1 U14965 ( .A1(n15177), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15203), 
        .B2(n12665), .ZN(n12666) );
  OAI21_X1 U14966 ( .B1(n12919), .B2(n15100), .A(n12666), .ZN(n12667) );
  AOI21_X1 U14967 ( .B1(n12845), .B2(n15086), .A(n12667), .ZN(n12668) );
  OAI21_X1 U14968 ( .B1(n12669), .B2(n15177), .A(n12668), .ZN(P3_U3211) );
  XOR2_X1 U14969 ( .A(n12674), .B(n12670), .Z(n12849) );
  INV_X1 U14970 ( .A(n12849), .ZN(n12682) );
  INV_X1 U14971 ( .A(n12671), .ZN(n12672) );
  AOI21_X1 U14972 ( .B1(n12674), .B2(n12673), .A(n12672), .ZN(n12675) );
  OAI222_X1 U14973 ( .A1(n15185), .A2(n12676), .B1(n15187), .B2(n12704), .C1(
        n15130), .C2(n12675), .ZN(n12848) );
  INV_X1 U14974 ( .A(n12677), .ZN(n12923) );
  AOI22_X1 U14975 ( .A1(n15177), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15203), 
        .B2(n12678), .ZN(n12679) );
  OAI21_X1 U14976 ( .B1(n12923), .B2(n15100), .A(n12679), .ZN(n12680) );
  AOI21_X1 U14977 ( .B1(n12848), .B2(n15204), .A(n12680), .ZN(n12681) );
  OAI21_X1 U14978 ( .B1(n12682), .B2(n12805), .A(n12681), .ZN(P3_U3212) );
  XNOR2_X1 U14979 ( .A(n12683), .B(n12689), .ZN(n12684) );
  OAI222_X1 U14980 ( .A1(n15185), .A2(n12685), .B1(n15187), .B2(n12716), .C1(
        n15130), .C2(n12684), .ZN(n12854) );
  INV_X1 U14981 ( .A(n12854), .ZN(n12697) );
  INV_X1 U14982 ( .A(n12686), .ZN(n12687) );
  OAI22_X1 U14983 ( .A1(n15204), .A2(n12688), .B1(n12687), .B2(n15104), .ZN(
        n12693) );
  INV_X1 U14984 ( .A(n12855), .ZN(n12691) );
  AND2_X1 U14985 ( .A1(n12690), .A2(n12689), .ZN(n12853) );
  NOR3_X1 U14986 ( .A1(n12691), .A2(n12853), .A3(n12805), .ZN(n12692) );
  AOI211_X1 U14987 ( .C1(n12695), .C2(n12694), .A(n12693), .B(n12692), .ZN(
        n12696) );
  OAI21_X1 U14988 ( .B1(n12697), .B2(n15177), .A(n12696), .ZN(P3_U3213) );
  XNOR2_X1 U14989 ( .A(n12698), .B(n12700), .ZN(n12860) );
  INV_X1 U14990 ( .A(n12860), .ZN(n12709) );
  OAI211_X1 U14991 ( .C1(n12701), .C2(n12700), .A(n12699), .B(n15183), .ZN(
        n12703) );
  NAND2_X1 U14992 ( .A1(n12726), .A2(n15145), .ZN(n12702) );
  OAI211_X1 U14993 ( .C1(n12704), .C2(n15185), .A(n12703), .B(n12702), .ZN(
        n12859) );
  AOI22_X1 U14994 ( .A1(n15177), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15203), 
        .B2(n12705), .ZN(n12706) );
  OAI21_X1 U14995 ( .B1(n12931), .B2(n15100), .A(n12706), .ZN(n12707) );
  AOI21_X1 U14996 ( .B1(n12859), .B2(n15204), .A(n12707), .ZN(n12708) );
  OAI21_X1 U14997 ( .B1(n12709), .B2(n12805), .A(n12708), .ZN(P3_U3214) );
  INV_X1 U14998 ( .A(n12710), .ZN(n12711) );
  AOI21_X1 U14999 ( .B1(n12713), .B2(n12712), .A(n12711), .ZN(n12714) );
  OAI222_X1 U15000 ( .A1(n15185), .A2(n12716), .B1(n15187), .B2(n12715), .C1(
        n15130), .C2(n12714), .ZN(n12863) );
  INV_X1 U15001 ( .A(n12863), .ZN(n12723) );
  AOI21_X1 U15002 ( .B1(n12718), .B2(n12717), .A(n6529), .ZN(n12864) );
  AOI22_X1 U15003 ( .A1(n15177), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15203), 
        .B2(n12719), .ZN(n12720) );
  OAI21_X1 U15004 ( .B1(n12935), .B2(n15100), .A(n12720), .ZN(n12721) );
  AOI21_X1 U15005 ( .B1(n12864), .B2(n15086), .A(n12721), .ZN(n12722) );
  OAI21_X1 U15006 ( .B1(n12723), .B2(n15177), .A(n12722), .ZN(P3_U3215) );
  XNOR2_X1 U15007 ( .A(n12725), .B(n12724), .ZN(n12727) );
  AOI222_X1 U15008 ( .A1(n15183), .A2(n12727), .B1(n12726), .B2(n15142), .C1(
        n12751), .C2(n15145), .ZN(n12870) );
  NAND3_X1 U15009 ( .A1(n12743), .A2(n12729), .A3(n12728), .ZN(n12730) );
  NAND2_X1 U15010 ( .A1(n12731), .A2(n12730), .ZN(n12868) );
  AOI22_X1 U15011 ( .A1(n15177), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15203), 
        .B2(n12732), .ZN(n12733) );
  OAI21_X1 U15012 ( .B1(n12734), .B2(n15100), .A(n12733), .ZN(n12735) );
  AOI21_X1 U15013 ( .B1(n12868), .B2(n15086), .A(n12735), .ZN(n12736) );
  OAI21_X1 U15014 ( .B1(n12870), .B2(n15177), .A(n12736), .ZN(P3_U3216) );
  XNOR2_X1 U15015 ( .A(n12738), .B(n12737), .ZN(n12742) );
  NAND2_X1 U15016 ( .A1(n12739), .A2(n15142), .ZN(n12741) );
  NAND2_X1 U15017 ( .A1(n12769), .A2(n15145), .ZN(n12740) );
  AND2_X1 U15018 ( .A1(n12741), .A2(n12740), .ZN(n14438) );
  OAI21_X1 U15019 ( .B1(n12742), .B2(n15130), .A(n14438), .ZN(n12871) );
  INV_X1 U15020 ( .A(n12871), .ZN(n12749) );
  OAI21_X1 U15021 ( .B1(n12745), .B2(n12744), .A(n12743), .ZN(n12872) );
  INV_X1 U15022 ( .A(n14434), .ZN(n12940) );
  AOI22_X1 U15023 ( .A1(n15177), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15203), 
        .B2(n14435), .ZN(n12746) );
  OAI21_X1 U15024 ( .B1(n12940), .B2(n15100), .A(n12746), .ZN(n12747) );
  AOI21_X1 U15025 ( .B1(n12872), .B2(n15086), .A(n12747), .ZN(n12748) );
  OAI21_X1 U15026 ( .B1(n12749), .B2(n15177), .A(n12748), .ZN(P3_U3217) );
  XNOR2_X1 U15027 ( .A(n12750), .B(n12754), .ZN(n12752) );
  AOI222_X1 U15028 ( .A1(n15183), .A2(n12752), .B1(n12751), .B2(n15142), .C1(
        n12781), .C2(n15145), .ZN(n12878) );
  NAND3_X1 U15029 ( .A1(n12753), .A2(n7087), .A3(n12755), .ZN(n12756) );
  NAND2_X1 U15030 ( .A1(n12757), .A2(n12756), .ZN(n12876) );
  AOI22_X1 U15031 ( .A1(n15177), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15203), 
        .B2(n12758), .ZN(n12759) );
  OAI21_X1 U15032 ( .B1(n12760), .B2(n15100), .A(n12759), .ZN(n12761) );
  AOI21_X1 U15033 ( .B1(n12876), .B2(n15086), .A(n12761), .ZN(n12762) );
  OAI21_X1 U15034 ( .B1(n12878), .B2(n15177), .A(n12762), .ZN(P3_U3218) );
  OR2_X1 U15035 ( .A1(n12780), .A2(n12763), .ZN(n12768) );
  NAND2_X1 U15036 ( .A1(n12768), .A2(n12764), .ZN(n12766) );
  AOI21_X1 U15037 ( .B1(n12766), .B2(n12765), .A(n15130), .ZN(n12772) );
  NAND2_X1 U15038 ( .A1(n12768), .A2(n12767), .ZN(n12771) );
  NAND2_X1 U15039 ( .A1(n12769), .A2(n15142), .ZN(n12770) );
  OAI21_X1 U15040 ( .B1(n12798), .B2(n15187), .A(n12770), .ZN(n14421) );
  AOI21_X1 U15041 ( .B1(n12772), .B2(n12771), .A(n14421), .ZN(n12881) );
  NAND2_X1 U15042 ( .A1(n12774), .A2(n12773), .ZN(n12775) );
  NAND2_X1 U15043 ( .A1(n12753), .A2(n12775), .ZN(n12879) );
  AOI22_X1 U15044 ( .A1(n15177), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15203), 
        .B2(n12776), .ZN(n12777) );
  OAI21_X1 U15045 ( .B1(n15100), .B2(n14424), .A(n12777), .ZN(n12778) );
  AOI21_X1 U15046 ( .B1(n12879), .B2(n15086), .A(n12778), .ZN(n12779) );
  OAI21_X1 U15047 ( .B1(n12881), .B2(n15177), .A(n12779), .ZN(P3_U3219) );
  XNOR2_X1 U15048 ( .A(n12780), .B(n7489), .ZN(n12784) );
  NAND2_X1 U15049 ( .A1(n12781), .A2(n15142), .ZN(n12782) );
  OAI21_X1 U15050 ( .B1(n14496), .B2(n15187), .A(n12782), .ZN(n12783) );
  AOI21_X1 U15051 ( .B1(n12784), .B2(n15183), .A(n12783), .ZN(n14504) );
  NOR2_X1 U15052 ( .A1(n12785), .A2(n15219), .ZN(n14501) );
  INV_X1 U15053 ( .A(n12786), .ZN(n12787) );
  OAI22_X1 U15054 ( .A1(n15204), .A2(n8480), .B1(n12787), .B2(n15104), .ZN(
        n12788) );
  AOI21_X1 U15055 ( .B1(n14501), .B2(n15173), .A(n12788), .ZN(n12791) );
  XNOR2_X1 U15056 ( .A(n12789), .B(n7489), .ZN(n14502) );
  NAND2_X1 U15057 ( .A1(n14502), .A2(n15086), .ZN(n12790) );
  OAI211_X1 U15058 ( .C1(n14504), .C2(n15177), .A(n12791), .B(n12790), .ZN(
        P3_U3220) );
  XNOR2_X1 U15059 ( .A(n12793), .B(n12792), .ZN(n14508) );
  INV_X1 U15060 ( .A(n14508), .ZN(n12804) );
  XNOR2_X1 U15061 ( .A(n12795), .B(n12794), .ZN(n12796) );
  OAI222_X1 U15062 ( .A1(n15185), .A2(n12798), .B1(n15187), .B2(n12797), .C1(
        n12796), .C2(n15130), .ZN(n14506) );
  NAND2_X1 U15063 ( .A1(n14506), .A2(n15204), .ZN(n12803) );
  NOR2_X1 U15064 ( .A1(n12799), .A2(n15219), .ZN(n14507) );
  OAI22_X1 U15065 ( .A1(n15204), .A2(n8455), .B1(n12800), .B2(n15104), .ZN(
        n12801) );
  AOI21_X1 U15066 ( .B1(n15173), .B2(n14507), .A(n12801), .ZN(n12802) );
  OAI211_X1 U15067 ( .C1(n12805), .C2(n12804), .A(n12803), .B(n12802), .ZN(
        P3_U3221) );
  NOR2_X1 U15068 ( .A1(n12885), .A2(n15270), .ZN(n12807) );
  AOI21_X1 U15069 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n15270), .A(n12807), 
        .ZN(n12806) );
  OAI21_X1 U15070 ( .B1(n12887), .B2(n12884), .A(n12806), .ZN(P3_U3490) );
  AOI21_X1 U15071 ( .B1(P3_REG1_REG_30__SCAN_IN), .B2(n15270), .A(n12807), 
        .ZN(n12808) );
  OAI21_X1 U15072 ( .B1(n12890), .B2(n12884), .A(n12808), .ZN(P3_U3489) );
  NAND2_X1 U15073 ( .A1(n12810), .A2(n15199), .ZN(n12838) );
  INV_X1 U15074 ( .A(n12891), .ZN(n12814) );
  INV_X1 U15075 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12820) );
  AND2_X1 U15076 ( .A1(n12817), .A2(n12811), .ZN(n12818) );
  NOR2_X1 U15077 ( .A1(n12819), .A2(n12818), .ZN(n12895) );
  INV_X1 U15078 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12823) );
  AOI21_X1 U15079 ( .B1(n12811), .B2(n12822), .A(n12821), .ZN(n12898) );
  MUX2_X1 U15080 ( .A(n12823), .B(n12898), .S(n15269), .Z(n12824) );
  OAI21_X1 U15081 ( .B1(n12901), .B2(n12884), .A(n12824), .ZN(P3_U3486) );
  INV_X1 U15082 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12827) );
  AOI21_X1 U15083 ( .B1(n12826), .B2(n12811), .A(n12825), .ZN(n12902) );
  MUX2_X1 U15084 ( .A(n12827), .B(n12902), .S(n15269), .Z(n12828) );
  OAI21_X1 U15085 ( .B1(n12905), .B2(n12884), .A(n12828), .ZN(P3_U3485) );
  AOI22_X1 U15086 ( .A1(n12830), .A2(n12811), .B1(n15242), .B2(n12829), .ZN(
        n12831) );
  NAND2_X1 U15087 ( .A1(n12832), .A2(n12831), .ZN(n12906) );
  MUX2_X1 U15088 ( .A(n12906), .B(P3_REG1_REG_25__SCAN_IN), .S(n15270), .Z(
        P3_U3484) );
  NAND2_X1 U15089 ( .A1(n12833), .A2(n12811), .ZN(n12834) );
  NAND2_X1 U15090 ( .A1(n12835), .A2(n12834), .ZN(n12907) );
  MUX2_X1 U15091 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n12907), .S(n15269), .Z(
        n12836) );
  AOI21_X1 U15092 ( .B1(n6692), .B2(n12909), .A(n12836), .ZN(n12837) );
  INV_X1 U15093 ( .A(n12837), .ZN(P3_U3483) );
  INV_X1 U15094 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12842) );
  INV_X1 U15095 ( .A(n12839), .ZN(n12841) );
  AOI21_X1 U15096 ( .B1(n15243), .B2(n12841), .A(n12840), .ZN(n12912) );
  MUX2_X1 U15097 ( .A(n12842), .B(n12912), .S(n15269), .Z(n12843) );
  OAI21_X1 U15098 ( .B1(n12915), .B2(n12884), .A(n12843), .ZN(P3_U3482) );
  AOI21_X1 U15099 ( .B1(n12811), .B2(n12845), .A(n12844), .ZN(n12916) );
  MUX2_X1 U15100 ( .A(n12846), .B(n12916), .S(n15269), .Z(n12847) );
  OAI21_X1 U15101 ( .B1(n12919), .B2(n12884), .A(n12847), .ZN(P3_U3481) );
  INV_X1 U15102 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12850) );
  AOI21_X1 U15103 ( .B1(n12811), .B2(n12849), .A(n12848), .ZN(n12920) );
  MUX2_X1 U15104 ( .A(n12850), .B(n12920), .S(n15269), .Z(n12851) );
  OAI21_X1 U15105 ( .B1(n12923), .B2(n12884), .A(n12851), .ZN(P3_U3480) );
  INV_X1 U15106 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12857) );
  NOR2_X1 U15107 ( .A1(n12853), .A2(n12852), .ZN(n12856) );
  AOI21_X1 U15108 ( .B1(n12856), .B2(n12855), .A(n12854), .ZN(n12924) );
  MUX2_X1 U15109 ( .A(n12857), .B(n12924), .S(n15269), .Z(n12858) );
  OAI21_X1 U15110 ( .B1(n12927), .B2(n12884), .A(n12858), .ZN(P3_U3479) );
  AOI21_X1 U15111 ( .B1(n12811), .B2(n12860), .A(n12859), .ZN(n12928) );
  MUX2_X1 U15112 ( .A(n12861), .B(n12928), .S(n15269), .Z(n12862) );
  OAI21_X1 U15113 ( .B1(n12884), .B2(n12931), .A(n12862), .ZN(P3_U3478) );
  AOI21_X1 U15114 ( .B1(n12864), .B2(n12811), .A(n12863), .ZN(n12932) );
  MUX2_X1 U15115 ( .A(n12865), .B(n12932), .S(n15269), .Z(n12866) );
  OAI21_X1 U15116 ( .B1(n12935), .B2(n12884), .A(n12866), .ZN(P3_U3477) );
  AOI22_X1 U15117 ( .A1(n12868), .A2(n12811), .B1(n15242), .B2(n12867), .ZN(
        n12869) );
  NAND2_X1 U15118 ( .A1(n12870), .A2(n12869), .ZN(n12936) );
  MUX2_X1 U15119 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12936), .S(n15269), .Z(
        P3_U3476) );
  AOI21_X1 U15120 ( .B1(n12811), .B2(n12872), .A(n12871), .ZN(n12937) );
  MUX2_X1 U15121 ( .A(n12873), .B(n12937), .S(n15269), .Z(n12874) );
  OAI21_X1 U15122 ( .B1(n12940), .B2(n12884), .A(n12874), .ZN(P3_U3475) );
  AOI22_X1 U15123 ( .A1(n12876), .A2(n12811), .B1(n15242), .B2(n12875), .ZN(
        n12877) );
  NAND2_X1 U15124 ( .A1(n12878), .A2(n12877), .ZN(n12941) );
  MUX2_X1 U15125 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n12941), .S(n15269), .Z(
        P3_U3474) );
  NAND2_X1 U15126 ( .A1(n12879), .A2(n12811), .ZN(n12880) );
  AND2_X1 U15127 ( .A1(n12881), .A2(n12880), .ZN(n12943) );
  INV_X1 U15128 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12882) );
  MUX2_X1 U15129 ( .A(n12943), .B(n12882), .S(n15270), .Z(n12883) );
  OAI21_X1 U15130 ( .B1(n12884), .B2(n14424), .A(n12883), .ZN(P3_U3473) );
  INV_X1 U15131 ( .A(n12910), .ZN(n12945) );
  NOR2_X1 U15132 ( .A1(n12885), .A2(n15252), .ZN(n12888) );
  AOI21_X1 U15133 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n15252), .A(n12888), 
        .ZN(n12886) );
  OAI21_X1 U15134 ( .B1(n12887), .B2(n12945), .A(n12886), .ZN(P3_U3458) );
  AOI21_X1 U15135 ( .B1(P3_REG0_REG_30__SCAN_IN), .B2(n15252), .A(n12888), 
        .ZN(n12889) );
  OAI21_X1 U15136 ( .B1(n12890), .B2(n12945), .A(n12889), .ZN(P3_U3457) );
  INV_X1 U15137 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n12892) );
  MUX2_X1 U15138 ( .A(n12899), .B(n12898), .S(n15253), .Z(n12900) );
  OAI21_X1 U15139 ( .B1(n12901), .B2(n12945), .A(n12900), .ZN(P3_U3454) );
  MUX2_X1 U15140 ( .A(n12903), .B(n12902), .S(n15253), .Z(n12904) );
  OAI21_X1 U15141 ( .B1(n12905), .B2(n12945), .A(n12904), .ZN(P3_U3453) );
  MUX2_X1 U15142 ( .A(n12906), .B(P3_REG0_REG_25__SCAN_IN), .S(n15252), .Z(
        P3_U3452) );
  MUX2_X1 U15143 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n12907), .S(n15253), .Z(
        n12908) );
  AOI21_X1 U15144 ( .B1(n12910), .B2(n12909), .A(n12908), .ZN(n12911) );
  INV_X1 U15145 ( .A(n12911), .ZN(P3_U3451) );
  MUX2_X1 U15146 ( .A(n12913), .B(n12912), .S(n15253), .Z(n12914) );
  OAI21_X1 U15147 ( .B1(n12915), .B2(n12945), .A(n12914), .ZN(P3_U3450) );
  INV_X1 U15148 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12917) );
  MUX2_X1 U15149 ( .A(n12917), .B(n12916), .S(n15253), .Z(n12918) );
  OAI21_X1 U15150 ( .B1(n12919), .B2(n12945), .A(n12918), .ZN(P3_U3449) );
  MUX2_X1 U15151 ( .A(n12921), .B(n12920), .S(n15253), .Z(n12922) );
  OAI21_X1 U15152 ( .B1(n12923), .B2(n12945), .A(n12922), .ZN(P3_U3448) );
  MUX2_X1 U15153 ( .A(n12925), .B(n12924), .S(n15253), .Z(n12926) );
  OAI21_X1 U15154 ( .B1(n12927), .B2(n12945), .A(n12926), .ZN(P3_U3447) );
  INV_X1 U15155 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12929) );
  MUX2_X1 U15156 ( .A(n12929), .B(n12928), .S(n15253), .Z(n12930) );
  OAI21_X1 U15157 ( .B1(n12945), .B2(n12931), .A(n12930), .ZN(P3_U3446) );
  MUX2_X1 U15158 ( .A(n12933), .B(n12932), .S(n15253), .Z(n12934) );
  OAI21_X1 U15159 ( .B1(n12935), .B2(n12945), .A(n12934), .ZN(P3_U3444) );
  MUX2_X1 U15160 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n12936), .S(n15253), .Z(
        P3_U3441) );
  MUX2_X1 U15161 ( .A(n12938), .B(n12937), .S(n15253), .Z(n12939) );
  OAI21_X1 U15162 ( .B1(n12940), .B2(n12945), .A(n12939), .ZN(P3_U3438) );
  MUX2_X1 U15163 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n12941), .S(n15253), .Z(
        P3_U3435) );
  INV_X1 U15164 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12942) );
  MUX2_X1 U15165 ( .A(n12943), .B(n12942), .S(n15252), .Z(n12944) );
  OAI21_X1 U15166 ( .B1(n12945), .B2(n14424), .A(n12944), .ZN(P3_U3432) );
  MUX2_X1 U15167 ( .A(P3_D_REG_1__SCAN_IN), .B(n12946), .S(n12947), .Z(
        P3_U3377) );
  MUX2_X1 U15168 ( .A(P3_D_REG_0__SCAN_IN), .B(n12948), .S(n12947), .Z(
        P3_U3376) );
  INV_X1 U15169 ( .A(n12949), .ZN(n12954) );
  NOR4_X1 U15170 ( .A1(n12950), .A2(P3_IR_REG_30__SCAN_IN), .A3(n6724), .A4(
        P3_U3151), .ZN(n12951) );
  AOI21_X1 U15171 ( .B1(n12952), .B2(SI_31_), .A(n12951), .ZN(n12953) );
  OAI21_X1 U15172 ( .B1(n12954), .B2(n6460), .A(n12953), .ZN(P3_U3264) );
  INV_X1 U15173 ( .A(SI_30_), .ZN(n12957) );
  INV_X1 U15174 ( .A(n12955), .ZN(n12956) );
  OAI222_X1 U15175 ( .A1(n12958), .A2(P3_U3151), .B1(n12966), .B2(n12957), 
        .C1(n6461), .C2(n12956), .ZN(P3_U3265) );
  OAI222_X1 U15176 ( .A1(P3_U3151), .A2(n12960), .B1(n6461), .B2(n6589), .C1(
        n12959), .C2(n12966), .ZN(P3_U3266) );
  INV_X1 U15177 ( .A(n12961), .ZN(n12963) );
  OAI222_X1 U15178 ( .A1(n12966), .A2(n12965), .B1(n6460), .B2(n12963), .C1(
        n12962), .C2(P3_U3151), .ZN(P3_U3267) );
  MUX2_X1 U15179 ( .A(n12967), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  XNOR2_X1 U15180 ( .A(n13288), .B(n10181), .ZN(n13004) );
  NAND2_X1 U15181 ( .A1(n13158), .A2(n12981), .ZN(n13005) );
  XNOR2_X1 U15182 ( .A(n13470), .B(n10181), .ZN(n13002) );
  NAND2_X1 U15183 ( .A1(n13159), .A2(n12981), .ZN(n13003) );
  XNOR2_X1 U15184 ( .A(n13409), .B(n6682), .ZN(n12978) );
  INV_X1 U15185 ( .A(n12978), .ZN(n12980) );
  NAND2_X1 U15186 ( .A1(n13166), .A2(n12981), .ZN(n12979) );
  AOI21_X1 U15187 ( .B1(n12970), .B2(n12969), .A(n12968), .ZN(n12973) );
  INV_X1 U15188 ( .A(n12970), .ZN(n12971) );
  XNOR2_X1 U15189 ( .A(n13520), .B(n6682), .ZN(n12975) );
  NAND2_X1 U15190 ( .A1(n13167), .A2(n14849), .ZN(n12976) );
  XNOR2_X1 U15191 ( .A(n12975), .B(n12976), .ZN(n13069) );
  INV_X1 U15192 ( .A(n12975), .ZN(n12977) );
  NAND2_X1 U15193 ( .A1(n12977), .A2(n12976), .ZN(n13091) );
  XOR2_X1 U15194 ( .A(n12979), .B(n12978), .Z(n13092) );
  XNOR2_X1 U15195 ( .A(n13507), .B(n10181), .ZN(n12982) );
  NAND2_X1 U15196 ( .A1(n13165), .A2(n12981), .ZN(n12983) );
  XNOR2_X1 U15197 ( .A(n12982), .B(n12983), .ZN(n13131) );
  XNOR2_X1 U15198 ( .A(n13500), .B(n13006), .ZN(n12987) );
  NAND2_X1 U15199 ( .A1(n13164), .A2(n14849), .ZN(n12986) );
  NAND2_X1 U15200 ( .A1(n12987), .A2(n12986), .ZN(n13025) );
  NOR2_X1 U15201 ( .A1(n12987), .A2(n12986), .ZN(n13027) );
  AND2_X1 U15202 ( .A1(n13163), .A2(n14849), .ZN(n12989) );
  XNOR2_X1 U15203 ( .A(n13562), .B(n10181), .ZN(n12988) );
  NOR2_X1 U15204 ( .A1(n12988), .A2(n12989), .ZN(n12990) );
  AOI21_X1 U15205 ( .B1(n12989), .B2(n12988), .A(n12990), .ZN(n13113) );
  INV_X1 U15206 ( .A(n12990), .ZN(n12991) );
  NAND2_X1 U15207 ( .A1(n13162), .A2(n14849), .ZN(n12992) );
  XNOR2_X1 U15208 ( .A(n13488), .B(n10181), .ZN(n12994) );
  XOR2_X1 U15209 ( .A(n12992), .B(n12994), .Z(n13052) );
  INV_X1 U15210 ( .A(n12992), .ZN(n12993) );
  NAND2_X1 U15211 ( .A1(n12994), .A2(n12993), .ZN(n12995) );
  XNOR2_X1 U15212 ( .A(n13331), .B(n10181), .ZN(n12997) );
  NAND2_X1 U15213 ( .A1(n13161), .A2(n10723), .ZN(n13122) );
  INV_X1 U15214 ( .A(n12996), .ZN(n12999) );
  INV_X1 U15215 ( .A(n12997), .ZN(n12998) );
  XNOR2_X1 U15216 ( .A(n13476), .B(n10181), .ZN(n13001) );
  NAND2_X1 U15217 ( .A1(n13160), .A2(n10723), .ZN(n13017) );
  XNOR2_X1 U15218 ( .A(n13002), .B(n13003), .ZN(n13102) );
  XNOR2_X1 U15219 ( .A(n13004), .B(n13005), .ZN(n13060) );
  XNOR2_X1 U15220 ( .A(n13543), .B(n13006), .ZN(n13008) );
  NAND2_X1 U15221 ( .A1(n13157), .A2(n10723), .ZN(n13007) );
  NAND2_X1 U15222 ( .A1(n13008), .A2(n13007), .ZN(n13009) );
  OAI21_X1 U15223 ( .B1(n13008), .B2(n13007), .A(n13009), .ZN(n13140) );
  XNOR2_X1 U15224 ( .A(n13010), .B(n10181), .ZN(n13037) );
  NAND2_X1 U15225 ( .A1(n13156), .A2(n10723), .ZN(n13036) );
  XNOR2_X1 U15226 ( .A(n13037), .B(n13036), .ZN(n13038) );
  XNOR2_X1 U15227 ( .A(n13039), .B(n13038), .ZN(n13016) );
  INV_X1 U15228 ( .A(n13256), .ZN(n13013) );
  OAI22_X1 U15229 ( .A1(n13011), .A2(n13074), .B1(n13063), .B2(n13072), .ZN(
        n13251) );
  AOI22_X1 U15230 ( .A1(n13251), .A2(n13097), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13012) );
  OAI21_X1 U15231 ( .B1(n13013), .B2(n13104), .A(n13012), .ZN(n13014) );
  AOI21_X1 U15232 ( .B1(n13448), .B2(n13149), .A(n13014), .ZN(n13015) );
  OAI21_X1 U15233 ( .B1(n13016), .B2(n13151), .A(n13015), .ZN(P2_U3186) );
  XNOR2_X1 U15234 ( .A(n13018), .B(n13017), .ZN(n13024) );
  NAND2_X1 U15235 ( .A1(n13159), .A2(n13144), .ZN(n13020) );
  NAND2_X1 U15236 ( .A1(n13161), .A2(n13142), .ZN(n13019) );
  NAND2_X1 U15237 ( .A1(n13020), .A2(n13019), .ZN(n13475) );
  AOI22_X1 U15238 ( .A1(n13475), .A2(n13097), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13021) );
  OAI21_X1 U15239 ( .B1(n13313), .B2(n13104), .A(n13021), .ZN(n13022) );
  AOI21_X1 U15240 ( .B1(n13476), .B2(n13149), .A(n13022), .ZN(n13023) );
  OAI21_X1 U15241 ( .B1(n13024), .B2(n13151), .A(n13023), .ZN(P2_U3188) );
  INV_X1 U15242 ( .A(n13025), .ZN(n13026) );
  NOR2_X1 U15243 ( .A1(n13027), .A2(n13026), .ZN(n13028) );
  XNOR2_X1 U15244 ( .A(n13029), .B(n13028), .ZN(n13035) );
  OAI22_X1 U15245 ( .A1(n13031), .A2(n13074), .B1(n13030), .B2(n13072), .ZN(
        n13371) );
  NAND2_X1 U15246 ( .A1(n13097), .A2(n13371), .ZN(n13032) );
  NAND2_X1 U15247 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13216)
         );
  OAI211_X1 U15248 ( .C1(n13104), .C2(n13376), .A(n13032), .B(n13216), .ZN(
        n13033) );
  AOI21_X1 U15249 ( .B1(n13500), .B2(n13149), .A(n13033), .ZN(n13034) );
  OAI21_X1 U15250 ( .B1(n13035), .B2(n13151), .A(n13034), .ZN(P2_U3191) );
  NAND2_X1 U15251 ( .A1(n13155), .A2(n10723), .ZN(n13040) );
  XNOR2_X1 U15252 ( .A(n13040), .B(n10181), .ZN(n13041) );
  XNOR2_X1 U15253 ( .A(n13540), .B(n13041), .ZN(n13042) );
  NAND2_X1 U15254 ( .A1(n13043), .A2(n13129), .ZN(n13051) );
  OR2_X1 U15255 ( .A1(n13044), .A2(n13074), .ZN(n13046) );
  NAND2_X1 U15256 ( .A1(n13156), .A2(n13142), .ZN(n13045) );
  NAND2_X1 U15257 ( .A1(n13046), .A2(n13045), .ZN(n13236) );
  OAI22_X1 U15258 ( .A1(n13239), .A2(n13104), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13047), .ZN(n13049) );
  NOR2_X1 U15259 ( .A1(n13540), .A2(n13137), .ZN(n13048) );
  AOI211_X1 U15260 ( .C1(n13097), .C2(n13236), .A(n13049), .B(n13048), .ZN(
        n13050) );
  NAND2_X1 U15261 ( .A1(n13051), .A2(n13050), .ZN(P2_U3192) );
  XNOR2_X1 U15262 ( .A(n13053), .B(n13052), .ZN(n13059) );
  NAND2_X1 U15263 ( .A1(n13161), .A2(n13144), .ZN(n13055) );
  NAND2_X1 U15264 ( .A1(n13163), .A2(n13142), .ZN(n13054) );
  NAND2_X1 U15265 ( .A1(n13055), .A2(n13054), .ZN(n13338) );
  AOI22_X1 U15266 ( .A1(n13097), .A2(n13338), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13056) );
  OAI21_X1 U15267 ( .B1(n13343), .B2(n13104), .A(n13056), .ZN(n13057) );
  AOI21_X1 U15268 ( .B1(n13488), .B2(n13149), .A(n13057), .ZN(n13058) );
  OAI21_X1 U15269 ( .B1(n13059), .B2(n13151), .A(n13058), .ZN(P2_U3195) );
  XNOR2_X1 U15270 ( .A(n13061), .B(n13060), .ZN(n13067) );
  OAI22_X1 U15271 ( .A1(n13063), .A2(n13074), .B1(n13062), .B2(n13072), .ZN(
        n13279) );
  AOI22_X1 U15272 ( .A1(n13279), .A2(n13097), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13064) );
  OAI21_X1 U15273 ( .B1(n13289), .B2(n13104), .A(n13064), .ZN(n13065) );
  AOI21_X1 U15274 ( .B1(n13288), .B2(n13149), .A(n13065), .ZN(n13066) );
  OAI21_X1 U15275 ( .B1(n13067), .B2(n13151), .A(n13066), .ZN(P2_U3197) );
  INV_X1 U15276 ( .A(n13520), .ZN(n13421) );
  OAI21_X1 U15277 ( .B1(n13070), .B2(n13069), .A(n13068), .ZN(n13071) );
  NAND2_X1 U15278 ( .A1(n13071), .A2(n13129), .ZN(n13080) );
  OAI22_X1 U15279 ( .A1(n13075), .A2(n13074), .B1(n13073), .B2(n13072), .ZN(
        n13414) );
  INV_X1 U15280 ( .A(n13414), .ZN(n13077) );
  OAI22_X1 U15281 ( .A1(n13147), .A2(n13077), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13076), .ZN(n13078) );
  AOI21_X1 U15282 ( .B1(n13418), .B2(n13145), .A(n13078), .ZN(n13079) );
  OAI211_X1 U15283 ( .C1(n13421), .C2(n13137), .A(n13080), .B(n13079), .ZN(
        P2_U3198) );
  OAI21_X1 U15284 ( .B1(n13083), .B2(n13082), .A(n13081), .ZN(n13084) );
  NAND2_X1 U15285 ( .A1(n13084), .A2(n13129), .ZN(n13090) );
  AND2_X1 U15286 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n14816) );
  AOI21_X1 U15287 ( .B1(n13097), .B2(n13085), .A(n14816), .ZN(n13089) );
  AOI22_X1 U15288 ( .A1(n13149), .A2(n13087), .B1(n13086), .B2(n13145), .ZN(
        n13088) );
  NAND3_X1 U15289 ( .A1(n13090), .A2(n13089), .A3(n13088), .ZN(P2_U3199) );
  AND3_X1 U15290 ( .A1(n13068), .A2(n13092), .A3(n13091), .ZN(n13093) );
  OAI21_X1 U15291 ( .B1(n13094), .B2(n13093), .A(n13129), .ZN(n13101) );
  NAND2_X1 U15292 ( .A1(n13165), .A2(n13144), .ZN(n13096) );
  NAND2_X1 U15293 ( .A1(n13167), .A2(n13142), .ZN(n13095) );
  NAND2_X1 U15294 ( .A1(n13096), .A2(n13095), .ZN(n13400) );
  AOI22_X1 U15295 ( .A1(n13097), .A2(n13400), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13098) );
  OAI21_X1 U15296 ( .B1(n13406), .B2(n13104), .A(n13098), .ZN(n13099) );
  AOI21_X1 U15297 ( .B1(n13409), .B2(n13149), .A(n13099), .ZN(n13100) );
  NAND2_X1 U15298 ( .A1(n13101), .A2(n13100), .ZN(P2_U3200) );
  XNOR2_X1 U15299 ( .A(n13103), .B(n13102), .ZN(n13110) );
  NOR2_X1 U15300 ( .A1(n13104), .A2(n13304), .ZN(n13108) );
  AND2_X1 U15301 ( .A1(n13160), .A2(n13142), .ZN(n13105) );
  AOI21_X1 U15302 ( .B1(n13158), .B2(n13144), .A(n13105), .ZN(n13467) );
  OAI22_X1 U15303 ( .A1(n13467), .A2(n13147), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13106), .ZN(n13107) );
  AOI211_X1 U15304 ( .C1(n13470), .C2(n13149), .A(n13108), .B(n13107), .ZN(
        n13109) );
  OAI21_X1 U15305 ( .B1(n13110), .B2(n13151), .A(n13109), .ZN(P2_U3201) );
  INV_X1 U15306 ( .A(n13562), .ZN(n13365) );
  OAI21_X1 U15307 ( .B1(n13113), .B2(n13112), .A(n13111), .ZN(n13114) );
  NAND2_X1 U15308 ( .A1(n13114), .A2(n13129), .ZN(n13121) );
  NAND2_X1 U15309 ( .A1(n13162), .A2(n13144), .ZN(n13116) );
  NAND2_X1 U15310 ( .A1(n13164), .A2(n13142), .ZN(n13115) );
  NAND2_X1 U15311 ( .A1(n13116), .A2(n13115), .ZN(n13355) );
  INV_X1 U15312 ( .A(n13355), .ZN(n13118) );
  OAI22_X1 U15313 ( .A1(n13147), .A2(n13118), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13117), .ZN(n13119) );
  AOI21_X1 U15314 ( .B1(n13362), .B2(n13145), .A(n13119), .ZN(n13120) );
  OAI211_X1 U15315 ( .C1(n13365), .C2(n13137), .A(n13121), .B(n13120), .ZN(
        P2_U3205) );
  XNOR2_X1 U15316 ( .A(n13123), .B(n13122), .ZN(n13128) );
  AOI22_X1 U15317 ( .A1(n13160), .A2(n13144), .B1(n13142), .B2(n13162), .ZN(
        n13328) );
  OAI22_X1 U15318 ( .A1(n13147), .A2(n13328), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13124), .ZN(n13125) );
  AOI21_X1 U15319 ( .B1(n13332), .B2(n13145), .A(n13125), .ZN(n13127) );
  NAND2_X1 U15320 ( .A1(n13331), .A2(n13149), .ZN(n13126) );
  OAI211_X1 U15321 ( .C1(n13128), .C2(n13151), .A(n13127), .B(n13126), .ZN(
        P2_U3207) );
  OAI211_X1 U15322 ( .C1(n6587), .C2(n13131), .A(n13130), .B(n13129), .ZN(
        n13136) );
  INV_X1 U15323 ( .A(n13390), .ZN(n13134) );
  AND2_X1 U15324 ( .A1(n13166), .A2(n13142), .ZN(n13132) );
  AOI21_X1 U15325 ( .B1(n13164), .B2(n13144), .A(n13132), .ZN(n13504) );
  NAND2_X1 U15326 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13186)
         );
  OAI21_X1 U15327 ( .B1(n13147), .B2(n13504), .A(n13186), .ZN(n13133) );
  AOI21_X1 U15328 ( .B1(n13134), .B2(n13145), .A(n13133), .ZN(n13135) );
  OAI211_X1 U15329 ( .C1(n13394), .C2(n13137), .A(n13136), .B(n13135), .ZN(
        P2_U3210) );
  INV_X1 U15330 ( .A(n13138), .ZN(n13139) );
  AOI21_X1 U15331 ( .B1(n13141), .B2(n13140), .A(n13139), .ZN(n13152) );
  AND2_X1 U15332 ( .A1(n13158), .A2(n13142), .ZN(n13143) );
  AOI21_X1 U15333 ( .B1(n13156), .B2(n13144), .A(n13143), .ZN(n13268) );
  AOI22_X1 U15334 ( .A1(n13272), .A2(n13145), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13146) );
  OAI21_X1 U15335 ( .B1(n13268), .B2(n13147), .A(n13146), .ZN(n13148) );
  AOI21_X1 U15336 ( .B1(n13543), .B2(n13149), .A(n13148), .ZN(n13150) );
  OAI21_X1 U15337 ( .B1(n13152), .B2(n13151), .A(n13150), .ZN(P2_U3212) );
  MUX2_X1 U15338 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13220), .S(n6477), .Z(
        P2_U3562) );
  MUX2_X1 U15339 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13153), .S(n6477), .Z(
        P2_U3561) );
  MUX2_X1 U15340 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13154), .S(n6477), .Z(
        P2_U3560) );
  MUX2_X1 U15341 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13155), .S(n6477), .Z(
        P2_U3559) );
  MUX2_X1 U15342 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13156), .S(n6477), .Z(
        P2_U3558) );
  MUX2_X1 U15343 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13157), .S(n6477), .Z(
        P2_U3557) );
  MUX2_X1 U15344 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13158), .S(n6477), .Z(
        P2_U3556) );
  MUX2_X1 U15345 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13159), .S(n6477), .Z(
        P2_U3555) );
  MUX2_X1 U15346 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13160), .S(n6477), .Z(
        P2_U3554) );
  MUX2_X1 U15347 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13161), .S(n6477), .Z(
        P2_U3553) );
  MUX2_X1 U15348 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13162), .S(n6477), .Z(
        P2_U3552) );
  MUX2_X1 U15349 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13163), .S(n6477), .Z(
        P2_U3551) );
  MUX2_X1 U15350 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13164), .S(n6477), .Z(
        P2_U3550) );
  MUX2_X1 U15351 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13165), .S(n6477), .Z(
        P2_U3549) );
  MUX2_X1 U15352 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13166), .S(n6477), .Z(
        P2_U3548) );
  MUX2_X1 U15353 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13167), .S(n6477), .Z(
        P2_U3547) );
  MUX2_X1 U15354 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13168), .S(n6477), .Z(
        P2_U3546) );
  MUX2_X1 U15355 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13169), .S(n6477), .Z(
        P2_U3545) );
  MUX2_X1 U15356 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13170), .S(n6477), .Z(
        P2_U3544) );
  MUX2_X1 U15357 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13171), .S(n6477), .Z(
        P2_U3543) );
  MUX2_X1 U15358 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13172), .S(n6477), .Z(
        P2_U3542) );
  MUX2_X1 U15359 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13173), .S(n6477), .Z(
        P2_U3541) );
  MUX2_X1 U15360 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13174), .S(n6477), .Z(
        P2_U3540) );
  MUX2_X1 U15361 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13175), .S(n6477), .Z(
        P2_U3539) );
  MUX2_X1 U15362 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13176), .S(n6477), .Z(
        P2_U3538) );
  MUX2_X1 U15363 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13177), .S(n6477), .Z(
        P2_U3537) );
  MUX2_X1 U15364 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13178), .S(n6477), .Z(
        P2_U3536) );
  MUX2_X1 U15365 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13179), .S(n6477), .Z(
        P2_U3535) );
  MUX2_X1 U15366 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13180), .S(n6477), .Z(
        P2_U3534) );
  MUX2_X1 U15367 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13181), .S(n6477), .Z(
        P2_U3533) );
  MUX2_X1 U15368 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n13182), .S(n6477), .Z(
        P2_U3532) );
  MUX2_X1 U15369 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n9472), .S(n6477), .Z(
        P2_U3531) );
  OAI21_X1 U15370 ( .B1(n13184), .B2(n13407), .A(n13183), .ZN(n13203) );
  XOR2_X1 U15371 ( .A(n13203), .B(n13197), .Z(n13185) );
  NOR2_X1 U15372 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13185), .ZN(n13205) );
  AOI21_X1 U15373 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13185), .A(n13205), 
        .ZN(n13196) );
  INV_X1 U15374 ( .A(n13186), .ZN(n13192) );
  XNOR2_X1 U15375 ( .A(n13197), .B(n13198), .ZN(n13190) );
  INV_X1 U15376 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13189) );
  NOR2_X1 U15377 ( .A1(n13189), .A2(n13190), .ZN(n13200) );
  AOI211_X1 U15378 ( .C1(n13190), .C2(n13189), .A(n13200), .B(n14803), .ZN(
        n13191) );
  AOI211_X1 U15379 ( .C1(n14781), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n13192), 
        .B(n13191), .ZN(n13194) );
  NAND2_X1 U15380 ( .A1(n14818), .A2(n13204), .ZN(n13193) );
  OAI211_X1 U15381 ( .C1(n13196), .C2(n13195), .A(n13194), .B(n13193), .ZN(
        P2_U3232) );
  NOR2_X1 U15382 ( .A1(n13198), .A2(n13197), .ZN(n13199) );
  NOR2_X1 U15383 ( .A1(n13200), .A2(n13199), .ZN(n13202) );
  INV_X1 U15384 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13201) );
  XOR2_X1 U15385 ( .A(n13202), .B(n13201), .Z(n13212) );
  NOR2_X1 U15386 ( .A1(n13204), .A2(n13203), .ZN(n13206) );
  NOR2_X1 U15387 ( .A1(n13206), .A2(n13205), .ZN(n13207) );
  XNOR2_X1 U15388 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13207), .ZN(n13210) );
  AOI21_X1 U15389 ( .B1(n13210), .B2(n14820), .A(n14818), .ZN(n13208) );
  OAI21_X1 U15390 ( .B1(n13212), .B2(n14803), .A(n13208), .ZN(n13209) );
  INV_X1 U15391 ( .A(n13209), .ZN(n13215) );
  INV_X1 U15392 ( .A(n13210), .ZN(n13211) );
  AOI22_X1 U15393 ( .A1(n13212), .A2(n14811), .B1(n14820), .B2(n13211), .ZN(
        n13214) );
  MUX2_X1 U15394 ( .A(n13215), .B(n13214), .S(n13213), .Z(n13217) );
  OAI211_X1 U15395 ( .C1(n13218), .C2(n14825), .A(n13217), .B(n13216), .ZN(
        P2_U3233) );
  NAND2_X1 U15396 ( .A1(n13536), .A2(n13225), .ZN(n13224) );
  XNOR2_X1 U15397 ( .A(n9430), .B(n13224), .ZN(n13219) );
  NAND2_X1 U15398 ( .A1(n13430), .A2(n14854), .ZN(n13223) );
  AND2_X1 U15399 ( .A1(n13221), .A2(n13220), .ZN(n13429) );
  INV_X1 U15400 ( .A(n13429), .ZN(n13433) );
  NOR2_X1 U15401 ( .A1(n14873), .A2(n13433), .ZN(n13227) );
  AOI21_X1 U15402 ( .B1(n14873), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13227), 
        .ZN(n13222) );
  OAI211_X1 U15403 ( .C1(n13532), .C2(n13420), .A(n13223), .B(n13222), .ZN(
        P2_U3234) );
  OAI211_X1 U15404 ( .C1(n13536), .C2(n13225), .A(n13405), .B(n13224), .ZN(
        n13434) );
  NOR2_X1 U15405 ( .A1(n13536), .A2(n13420), .ZN(n13226) );
  AOI211_X1 U15406 ( .C1(n14873), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13227), 
        .B(n13226), .ZN(n13228) );
  OAI21_X1 U15407 ( .B1(n14833), .B2(n13434), .A(n13228), .ZN(P2_U3235) );
  OAI21_X1 U15408 ( .B1(n13232), .B2(n13230), .A(n13229), .ZN(n13444) );
  NAND2_X1 U15409 ( .A1(n13250), .A2(n13231), .ZN(n13233) );
  NAND2_X1 U15410 ( .A1(n13233), .A2(n13232), .ZN(n13234) );
  NAND3_X1 U15411 ( .A1(n13235), .A2(n14860), .A3(n13234), .ZN(n13238) );
  INV_X1 U15412 ( .A(n13236), .ZN(n13237) );
  OAI21_X1 U15413 ( .B1(n13239), .B2(n14865), .A(n13443), .ZN(n13240) );
  NAND2_X1 U15414 ( .A1(n13240), .A2(n14871), .ZN(n13247) );
  OAI21_X1 U15415 ( .B1(n13540), .B2(n13254), .A(n13405), .ZN(n13241) );
  INV_X1 U15416 ( .A(n13442), .ZN(n13245) );
  INV_X1 U15417 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13243) );
  OAI22_X1 U15418 ( .A1(n13540), .A2(n13420), .B1(n14871), .B2(n13243), .ZN(
        n13244) );
  AOI21_X1 U15419 ( .B1(n13245), .B2(n14854), .A(n13244), .ZN(n13246) );
  OAI211_X1 U15420 ( .C1(n13425), .C2(n13444), .A(n13247), .B(n13246), .ZN(
        P2_U3237) );
  NAND2_X1 U15421 ( .A1(n13248), .A2(n13260), .ZN(n13249) );
  NAND2_X1 U15422 ( .A1(n13250), .A2(n13249), .ZN(n13252) );
  AOI21_X1 U15423 ( .B1(n13252), .B2(n14860), .A(n13251), .ZN(n13453) );
  NAND2_X1 U15424 ( .A1(n13448), .A2(n13270), .ZN(n13253) );
  NAND2_X1 U15425 ( .A1(n13253), .A2(n13405), .ZN(n13255) );
  OR2_X1 U15426 ( .A1(n13255), .A2(n13254), .ZN(n13449) );
  AOI22_X1 U15427 ( .A1(n13256), .A2(n14844), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14873), .ZN(n13258) );
  NAND2_X1 U15428 ( .A1(n13448), .A2(n14846), .ZN(n13257) );
  OAI211_X1 U15429 ( .C1(n13449), .C2(n14833), .A(n13258), .B(n13257), .ZN(
        n13259) );
  INV_X1 U15430 ( .A(n13259), .ZN(n13263) );
  OR2_X1 U15431 ( .A1(n13261), .A2(n13260), .ZN(n13446) );
  NAND3_X1 U15432 ( .A1(n13447), .A2(n13446), .A3(n14855), .ZN(n13262) );
  OAI211_X1 U15433 ( .C1(n13453), .C2(n14873), .A(n13263), .B(n13262), .ZN(
        P2_U3238) );
  XNOR2_X1 U15434 ( .A(n13266), .B(n13264), .ZN(n13458) );
  OAI211_X1 U15435 ( .C1(n13267), .C2(n13266), .A(n13265), .B(n14860), .ZN(
        n13269) );
  AND2_X1 U15436 ( .A1(n13269), .A2(n13268), .ZN(n13457) );
  INV_X1 U15437 ( .A(n13457), .ZN(n13276) );
  AOI21_X1 U15438 ( .B1(n13543), .B2(n13285), .A(n14849), .ZN(n13271) );
  NAND2_X1 U15439 ( .A1(n13271), .A2(n13270), .ZN(n13456) );
  AOI22_X1 U15440 ( .A1(n13272), .A2(n14844), .B1(n14873), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n13274) );
  NAND2_X1 U15441 ( .A1(n13543), .A2(n14846), .ZN(n13273) );
  OAI211_X1 U15442 ( .C1(n13456), .C2(n14833), .A(n13274), .B(n13273), .ZN(
        n13275) );
  AOI21_X1 U15443 ( .B1(n13276), .B2(n14871), .A(n13275), .ZN(n13277) );
  OAI21_X1 U15444 ( .B1(n13425), .B2(n13458), .A(n13277), .ZN(P2_U3239) );
  XNOR2_X1 U15445 ( .A(n13278), .B(n13283), .ZN(n13281) );
  INV_X1 U15446 ( .A(n13279), .ZN(n13280) );
  OAI21_X1 U15447 ( .B1(n13281), .B2(n13368), .A(n13280), .ZN(n13463) );
  INV_X1 U15448 ( .A(n13463), .ZN(n13295) );
  OAI21_X1 U15449 ( .B1(n13284), .B2(n13283), .A(n13282), .ZN(n13464) );
  INV_X1 U15450 ( .A(n13297), .ZN(n13287) );
  INV_X1 U15451 ( .A(n13285), .ZN(n13286) );
  AOI211_X1 U15452 ( .C1(n13288), .C2(n13287), .A(n12981), .B(n13286), .ZN(
        n13462) );
  NAND2_X1 U15453 ( .A1(n13462), .A2(n14854), .ZN(n13292) );
  INV_X1 U15454 ( .A(n13289), .ZN(n13290) );
  AOI22_X1 U15455 ( .A1(n14873), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n13290), 
        .B2(n14844), .ZN(n13291) );
  OAI211_X1 U15456 ( .C1(n13551), .C2(n13420), .A(n13292), .B(n13291), .ZN(
        n13293) );
  AOI21_X1 U15457 ( .B1(n14855), .B2(n13464), .A(n13293), .ZN(n13294) );
  OAI21_X1 U15458 ( .B1(n14873), .B2(n13295), .A(n13294), .ZN(P2_U3240) );
  XNOR2_X1 U15459 ( .A(n13301), .B(n13296), .ZN(n13473) );
  AOI211_X1 U15460 ( .C1(n13470), .C2(n6466), .A(n14849), .B(n13297), .ZN(
        n13468) );
  INV_X1 U15461 ( .A(n13470), .ZN(n13299) );
  INV_X1 U15462 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13298) );
  OAI22_X1 U15463 ( .A1(n13299), .A2(n13420), .B1(n14871), .B2(n13298), .ZN(
        n13300) );
  AOI21_X1 U15464 ( .B1(n13468), .B2(n14854), .A(n13300), .ZN(n13307) );
  XNOR2_X1 U15465 ( .A(n13302), .B(n13301), .ZN(n13303) );
  NAND2_X1 U15466 ( .A1(n13303), .A2(n14860), .ZN(n13471) );
  OAI211_X1 U15467 ( .C1(n14865), .C2(n13304), .A(n13471), .B(n13467), .ZN(
        n13305) );
  NAND2_X1 U15468 ( .A1(n13305), .A2(n14871), .ZN(n13306) );
  OAI211_X1 U15469 ( .C1(n13425), .C2(n13473), .A(n13307), .B(n13306), .ZN(
        P2_U3241) );
  XNOR2_X1 U15470 ( .A(n13308), .B(n13309), .ZN(n13479) );
  XNOR2_X1 U15471 ( .A(n13310), .B(n13309), .ZN(n13311) );
  NAND2_X1 U15472 ( .A1(n13311), .A2(n14860), .ZN(n13477) );
  INV_X1 U15473 ( .A(n13475), .ZN(n13312) );
  OAI211_X1 U15474 ( .C1(n14865), .C2(n13313), .A(n13477), .B(n13312), .ZN(
        n13314) );
  NAND2_X1 U15475 ( .A1(n13314), .A2(n14871), .ZN(n13322) );
  INV_X1 U15476 ( .A(n6467), .ZN(n13317) );
  INV_X1 U15477 ( .A(n13315), .ZN(n13316) );
  AOI211_X1 U15478 ( .C1(n13476), .C2(n13317), .A(n14849), .B(n13316), .ZN(
        n13474) );
  INV_X1 U15479 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13318) );
  OAI22_X1 U15480 ( .A1(n13319), .A2(n13420), .B1(n13318), .B2(n14871), .ZN(
        n13320) );
  AOI21_X1 U15481 ( .B1(n13474), .B2(n14854), .A(n13320), .ZN(n13321) );
  OAI211_X1 U15482 ( .C1(n13425), .C2(n13479), .A(n13322), .B(n13321), .ZN(
        P2_U3242) );
  OAI21_X1 U15483 ( .B1(n13325), .B2(n13324), .A(n13323), .ZN(n13480) );
  XNOR2_X1 U15484 ( .A(n13327), .B(n13326), .ZN(n13329) );
  OAI21_X1 U15485 ( .B1(n13329), .B2(n13368), .A(n13328), .ZN(n13481) );
  NAND2_X1 U15486 ( .A1(n13481), .A2(n14871), .ZN(n13336) );
  AOI211_X1 U15487 ( .C1(n13331), .C2(n13340), .A(n14849), .B(n6467), .ZN(
        n13482) );
  INV_X1 U15488 ( .A(n13331), .ZN(n13558) );
  AOI22_X1 U15489 ( .A1(n14873), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13332), 
        .B2(n14844), .ZN(n13333) );
  OAI21_X1 U15490 ( .B1(n13558), .B2(n13420), .A(n13333), .ZN(n13334) );
  AOI21_X1 U15491 ( .B1(n13482), .B2(n14854), .A(n13334), .ZN(n13335) );
  OAI211_X1 U15492 ( .C1(n13425), .C2(n13480), .A(n13336), .B(n13335), .ZN(
        P2_U3243) );
  XOR2_X1 U15493 ( .A(n13337), .B(n13347), .Z(n13339) );
  AOI21_X1 U15494 ( .B1(n13339), .B2(n14860), .A(n13338), .ZN(n13490) );
  INV_X1 U15495 ( .A(n13361), .ZN(n13342) );
  INV_X1 U15496 ( .A(n13340), .ZN(n13341) );
  AOI211_X1 U15497 ( .C1(n13488), .C2(n13342), .A(n14849), .B(n13341), .ZN(
        n13487) );
  INV_X1 U15498 ( .A(n13343), .ZN(n13344) );
  AOI22_X1 U15499 ( .A1(n14873), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13344), 
        .B2(n14844), .ZN(n13345) );
  OAI21_X1 U15500 ( .B1(n13346), .B2(n13420), .A(n13345), .ZN(n13350) );
  XNOR2_X1 U15501 ( .A(n13348), .B(n13347), .ZN(n13491) );
  NOR2_X1 U15502 ( .A1(n13491), .A2(n13425), .ZN(n13349) );
  AOI211_X1 U15503 ( .C1(n13487), .C2(n14854), .A(n13350), .B(n13349), .ZN(
        n13351) );
  OAI21_X1 U15504 ( .B1(n13490), .B2(n14873), .A(n13351), .ZN(P2_U3244) );
  NAND2_X1 U15505 ( .A1(n13352), .A2(n13357), .ZN(n13353) );
  NAND2_X1 U15506 ( .A1(n13354), .A2(n13353), .ZN(n13356) );
  AOI21_X1 U15507 ( .B1(n13356), .B2(n14860), .A(n13355), .ZN(n13495) );
  XNOR2_X1 U15508 ( .A(n13358), .B(n13357), .ZN(n13493) );
  NAND2_X1 U15509 ( .A1(n13562), .A2(n13374), .ZN(n13359) );
  NAND2_X1 U15510 ( .A1(n13359), .A2(n13405), .ZN(n13360) );
  NOR2_X1 U15511 ( .A1(n13361), .A2(n13360), .ZN(n13492) );
  NAND2_X1 U15512 ( .A1(n13492), .A2(n14854), .ZN(n13364) );
  AOI22_X1 U15513 ( .A1(n14873), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13362), 
        .B2(n14844), .ZN(n13363) );
  OAI211_X1 U15514 ( .C1(n13365), .C2(n13420), .A(n13364), .B(n13363), .ZN(
        n13366) );
  AOI21_X1 U15515 ( .B1(n13493), .B2(n14855), .A(n13366), .ZN(n13367) );
  OAI21_X1 U15516 ( .B1(n13495), .B2(n14873), .A(n13367), .ZN(P2_U3245) );
  AOI21_X1 U15517 ( .B1(n13370), .B2(n13369), .A(n13368), .ZN(n13373) );
  AOI21_X1 U15518 ( .B1(n13373), .B2(n13372), .A(n13371), .ZN(n13502) );
  INV_X1 U15519 ( .A(n13374), .ZN(n13375) );
  AOI211_X1 U15520 ( .C1(n13500), .C2(n13392), .A(n14849), .B(n13375), .ZN(
        n13499) );
  INV_X1 U15521 ( .A(n13376), .ZN(n13377) );
  AOI22_X1 U15522 ( .A1(n14873), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13377), 
        .B2(n14844), .ZN(n13378) );
  OAI21_X1 U15523 ( .B1(n7207), .B2(n13420), .A(n13378), .ZN(n13382) );
  XNOR2_X1 U15524 ( .A(n13380), .B(n13379), .ZN(n13503) );
  NOR2_X1 U15525 ( .A1(n13503), .A2(n13425), .ZN(n13381) );
  AOI211_X1 U15526 ( .C1(n13499), .C2(n14854), .A(n13382), .B(n13381), .ZN(
        n13383) );
  OAI21_X1 U15527 ( .B1(n14873), .B2(n13502), .A(n13383), .ZN(P2_U3246) );
  OAI21_X1 U15528 ( .B1(n13385), .B2(n13387), .A(n13384), .ZN(n13386) );
  INV_X1 U15529 ( .A(n13386), .ZN(n13510) );
  XNOR2_X1 U15530 ( .A(n13388), .B(n13387), .ZN(n13389) );
  NAND2_X1 U15531 ( .A1(n13389), .A2(n14860), .ZN(n13508) );
  OAI211_X1 U15532 ( .C1(n14865), .C2(n13390), .A(n13508), .B(n13504), .ZN(
        n13391) );
  NAND2_X1 U15533 ( .A1(n13391), .A2(n14871), .ZN(n13397) );
  AOI211_X1 U15534 ( .C1(n13507), .C2(n13404), .A(n14849), .B(n7208), .ZN(
        n13505) );
  INV_X1 U15535 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13393) );
  OAI22_X1 U15536 ( .A1(n13394), .A2(n13420), .B1(n14871), .B2(n13393), .ZN(
        n13395) );
  AOI21_X1 U15537 ( .B1(n13505), .B2(n14854), .A(n13395), .ZN(n13396) );
  OAI211_X1 U15538 ( .C1(n13425), .C2(n13510), .A(n13397), .B(n13396), .ZN(
        P2_U3247) );
  INV_X1 U15539 ( .A(n13402), .ZN(n13398) );
  XNOR2_X1 U15540 ( .A(n13399), .B(n13398), .ZN(n13401) );
  AOI21_X1 U15541 ( .B1(n13401), .B2(n14860), .A(n13400), .ZN(n13516) );
  XNOR2_X1 U15542 ( .A(n13403), .B(n13402), .ZN(n13514) );
  OAI211_X1 U15543 ( .C1(n13416), .C2(n13512), .A(n13405), .B(n13404), .ZN(
        n13511) );
  OAI22_X1 U15544 ( .A1(n14871), .A2(n13407), .B1(n13406), .B2(n14865), .ZN(
        n13408) );
  AOI21_X1 U15545 ( .B1(n13409), .B2(n14846), .A(n13408), .ZN(n13410) );
  OAI21_X1 U15546 ( .B1(n13511), .B2(n14833), .A(n13410), .ZN(n13411) );
  AOI21_X1 U15547 ( .B1(n13514), .B2(n14855), .A(n13411), .ZN(n13412) );
  OAI21_X1 U15548 ( .B1(n13516), .B2(n14873), .A(n13412), .ZN(P2_U3248) );
  XNOR2_X1 U15549 ( .A(n13413), .B(n13422), .ZN(n13415) );
  AOI21_X1 U15550 ( .B1(n13415), .B2(n14860), .A(n13414), .ZN(n13522) );
  AOI211_X1 U15551 ( .C1(n13520), .C2(n13417), .A(n14849), .B(n13416), .ZN(
        n13519) );
  AOI22_X1 U15552 ( .A1(n14873), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n13418), 
        .B2(n14844), .ZN(n13419) );
  OAI21_X1 U15553 ( .B1(n13421), .B2(n13420), .A(n13419), .ZN(n13427) );
  NAND2_X1 U15554 ( .A1(n13423), .A2(n13422), .ZN(n13424) );
  NAND2_X1 U15555 ( .A1(n6832), .A2(n13424), .ZN(n13523) );
  NOR2_X1 U15556 ( .A1(n13523), .A2(n13425), .ZN(n13426) );
  AOI211_X1 U15557 ( .C1(n13519), .C2(n14854), .A(n13427), .B(n13426), .ZN(
        n13428) );
  OAI21_X1 U15558 ( .B1(n14873), .B2(n13522), .A(n13428), .ZN(P2_U3249) );
  NOR2_X1 U15559 ( .A1(n13430), .A2(n13429), .ZN(n13529) );
  MUX2_X1 U15560 ( .A(n13431), .B(n13529), .S(n14535), .Z(n13432) );
  AND2_X1 U15561 ( .A1(n13434), .A2(n13433), .ZN(n13533) );
  MUX2_X1 U15562 ( .A(n13435), .B(n13533), .S(n14535), .Z(n13436) );
  OAI21_X1 U15563 ( .B1(n13536), .B2(n13486), .A(n13436), .ZN(P2_U3529) );
  MUX2_X1 U15564 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13537), .S(n14954), .Z(
        P2_U3528) );
  OAI211_X1 U15565 ( .C1(n14938), .C2(n13444), .A(n13443), .B(n13442), .ZN(
        n13538) );
  OAI21_X1 U15566 ( .B1(n13540), .B2(n13486), .A(n13445), .ZN(P2_U3527) );
  NAND3_X1 U15567 ( .A1(n13447), .A2(n13446), .A3(n14921), .ZN(n13451) );
  NAND2_X1 U15568 ( .A1(n13448), .A2(n14933), .ZN(n13450) );
  AND3_X1 U15569 ( .A1(n13451), .A2(n13450), .A3(n13449), .ZN(n13452) );
  AND2_X1 U15570 ( .A1(n13453), .A2(n13452), .ZN(n13541) );
  MUX2_X1 U15571 ( .A(n13541), .B(n13454), .S(n14951), .Z(n13455) );
  INV_X1 U15572 ( .A(n13455), .ZN(P2_U3526) );
  OAI211_X1 U15573 ( .C1(n14938), .C2(n13458), .A(n13457), .B(n13456), .ZN(
        n13544) );
  MUX2_X1 U15574 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13544), .S(n14535), .Z(
        n13459) );
  INV_X1 U15575 ( .A(n13459), .ZN(n13461) );
  NAND2_X1 U15576 ( .A1(n13543), .A2(n13497), .ZN(n13460) );
  NAND2_X1 U15577 ( .A1(n13461), .A2(n13460), .ZN(P2_U3525) );
  AOI211_X1 U15578 ( .C1(n14921), .C2(n13464), .A(n13463), .B(n13462), .ZN(
        n13548) );
  MUX2_X1 U15579 ( .A(n13465), .B(n13548), .S(n14535), .Z(n13466) );
  OAI21_X1 U15580 ( .B1(n13551), .B2(n13486), .A(n13466), .ZN(P2_U3524) );
  INV_X1 U15581 ( .A(n13467), .ZN(n13469) );
  AOI211_X1 U15582 ( .C1(n13470), .C2(n14933), .A(n13469), .B(n13468), .ZN(
        n13472) );
  OAI211_X1 U15583 ( .C1(n14938), .C2(n13473), .A(n13472), .B(n13471), .ZN(
        n13552) );
  MUX2_X1 U15584 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13552), .S(n14535), .Z(
        P2_U3523) );
  AOI211_X1 U15585 ( .C1(n13476), .C2(n14933), .A(n13475), .B(n13474), .ZN(
        n13478) );
  OAI211_X1 U15586 ( .C1(n14938), .C2(n13479), .A(n13478), .B(n13477), .ZN(
        n13553) );
  MUX2_X1 U15587 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13553), .S(n14954), .Z(
        P2_U3522) );
  INV_X1 U15588 ( .A(n13480), .ZN(n13483) );
  AOI211_X1 U15589 ( .C1(n13483), .C2(n14921), .A(n13482), .B(n13481), .ZN(
        n13554) );
  MUX2_X1 U15590 ( .A(n13484), .B(n13554), .S(n14535), .Z(n13485) );
  OAI21_X1 U15591 ( .B1(n13558), .B2(n13486), .A(n13485), .ZN(P2_U3521) );
  AOI21_X1 U15592 ( .B1(n13488), .B2(n14933), .A(n13487), .ZN(n13489) );
  OAI211_X1 U15593 ( .C1(n14938), .C2(n13491), .A(n13490), .B(n13489), .ZN(
        n13559) );
  MUX2_X1 U15594 ( .A(n13559), .B(P2_REG1_REG_21__SCAN_IN), .S(n14951), .Z(
        P2_U3520) );
  AOI21_X1 U15595 ( .B1(n13493), .B2(n14921), .A(n13492), .ZN(n13494) );
  NAND2_X1 U15596 ( .A1(n13495), .A2(n13494), .ZN(n13560) );
  MUX2_X1 U15597 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13560), .S(n14535), .Z(
        n13496) );
  AOI21_X1 U15598 ( .B1(n13497), .B2(n13562), .A(n13496), .ZN(n13498) );
  INV_X1 U15599 ( .A(n13498), .ZN(P2_U3519) );
  AOI21_X1 U15600 ( .B1(n13500), .B2(n14933), .A(n13499), .ZN(n13501) );
  OAI211_X1 U15601 ( .C1(n14938), .C2(n13503), .A(n13502), .B(n13501), .ZN(
        n13565) );
  MUX2_X1 U15602 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13565), .S(n14535), .Z(
        P2_U3518) );
  INV_X1 U15603 ( .A(n13504), .ZN(n13506) );
  AOI211_X1 U15604 ( .C1(n13507), .C2(n14933), .A(n13506), .B(n13505), .ZN(
        n13509) );
  OAI211_X1 U15605 ( .C1(n13510), .C2(n14938), .A(n13509), .B(n13508), .ZN(
        n13566) );
  MUX2_X1 U15606 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13566), .S(n14535), .Z(
        P2_U3517) );
  INV_X1 U15607 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13517) );
  INV_X1 U15608 ( .A(n14933), .ZN(n14928) );
  OAI21_X1 U15609 ( .B1(n13512), .B2(n14928), .A(n13511), .ZN(n13513) );
  AOI21_X1 U15610 ( .B1(n13514), .B2(n14921), .A(n13513), .ZN(n13515) );
  AND2_X1 U15611 ( .A1(n13516), .A2(n13515), .ZN(n13567) );
  MUX2_X1 U15612 ( .A(n13517), .B(n13567), .S(n14535), .Z(n13518) );
  INV_X1 U15613 ( .A(n13518), .ZN(P2_U3516) );
  AOI21_X1 U15614 ( .B1(n13520), .B2(n14933), .A(n13519), .ZN(n13521) );
  OAI211_X1 U15615 ( .C1(n14938), .C2(n13523), .A(n13522), .B(n13521), .ZN(
        n13570) );
  MUX2_X1 U15616 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13570), .S(n14535), .Z(
        P2_U3515) );
  AOI21_X1 U15617 ( .B1(n13525), .B2(n14933), .A(n13524), .ZN(n13526) );
  OAI211_X1 U15618 ( .C1(n14938), .C2(n13528), .A(n13527), .B(n13526), .ZN(
        n13571) );
  MUX2_X1 U15619 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13571), .S(n14535), .Z(
        P2_U3514) );
  INV_X1 U15620 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13530) );
  MUX2_X1 U15621 ( .A(n13530), .B(n13529), .S(n14942), .Z(n13531) );
  OAI21_X1 U15622 ( .B1(n13532), .B2(n13557), .A(n13531), .ZN(P2_U3498) );
  INV_X1 U15623 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13534) );
  MUX2_X1 U15624 ( .A(n13534), .B(n13533), .S(n14942), .Z(n13535) );
  OAI21_X1 U15625 ( .B1(n13536), .B2(n13557), .A(n13535), .ZN(P2_U3497) );
  OAI21_X1 U15626 ( .B1(n13540), .B2(n13557), .A(n13539), .ZN(P2_U3495) );
  INV_X1 U15627 ( .A(n13541), .ZN(n13542) );
  MUX2_X1 U15628 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13542), .S(n14942), .Z(
        P2_U3494) );
  INV_X1 U15629 ( .A(n13543), .ZN(n13547) );
  MUX2_X1 U15630 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13544), .S(n14942), .Z(
        n13545) );
  INV_X1 U15631 ( .A(n13545), .ZN(n13546) );
  OAI21_X1 U15632 ( .B1(n13547), .B2(n13557), .A(n13546), .ZN(P2_U3493) );
  INV_X1 U15633 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n13549) );
  MUX2_X1 U15634 ( .A(n13549), .B(n13548), .S(n14942), .Z(n13550) );
  OAI21_X1 U15635 ( .B1(n13551), .B2(n13557), .A(n13550), .ZN(P2_U3492) );
  MUX2_X1 U15636 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13552), .S(n14942), .Z(
        P2_U3491) );
  MUX2_X1 U15637 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13553), .S(n14942), .Z(
        P2_U3490) );
  INV_X1 U15638 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n13555) );
  MUX2_X1 U15639 ( .A(n13555), .B(n13554), .S(n14942), .Z(n13556) );
  OAI21_X1 U15640 ( .B1(n13558), .B2(n13557), .A(n13556), .ZN(P2_U3489) );
  MUX2_X1 U15641 ( .A(n13559), .B(P2_REG0_REG_21__SCAN_IN), .S(n14940), .Z(
        P2_U3488) );
  MUX2_X1 U15642 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13560), .S(n14942), .Z(
        n13561) );
  AOI21_X1 U15643 ( .B1(n13563), .B2(n13562), .A(n13561), .ZN(n13564) );
  INV_X1 U15644 ( .A(n13564), .ZN(P2_U3487) );
  MUX2_X1 U15645 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13565), .S(n14942), .Z(
        P2_U3486) );
  MUX2_X1 U15646 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13566), .S(n14942), .Z(
        P2_U3484) );
  INV_X1 U15647 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n13568) );
  MUX2_X1 U15648 ( .A(n13568), .B(n13567), .S(n14942), .Z(n13569) );
  INV_X1 U15649 ( .A(n13569), .ZN(P2_U3481) );
  MUX2_X1 U15650 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13570), .S(n14942), .Z(
        P2_U3478) );
  MUX2_X1 U15651 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13571), .S(n14942), .Z(
        P2_U3475) );
  INV_X1 U15652 ( .A(n14236), .ZN(n13576) );
  NOR4_X1 U15653 ( .A1(n8887), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13573), .A4(
        P2_U3088), .ZN(n13574) );
  AOI21_X1 U15654 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n13585), .A(n13574), 
        .ZN(n13575) );
  OAI21_X1 U15655 ( .B1(n13576), .B2(n13587), .A(n13575), .ZN(P2_U3296) );
  AOI22_X1 U15656 ( .A1(n13577), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n13585), .ZN(n13578) );
  OAI21_X1 U15657 ( .B1(n13579), .B2(n13587), .A(n13578), .ZN(P2_U3297) );
  INV_X1 U15658 ( .A(n13580), .ZN(n14241) );
  OAI222_X1 U15659 ( .A1(n13599), .A2(n13582), .B1(n13587), .B2(n14241), .C1(
        n13581), .C2(P2_U3088), .ZN(P2_U3298) );
  INV_X1 U15660 ( .A(n13583), .ZN(n14244) );
  AOI21_X1 U15661 ( .B1(n13585), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13584), 
        .ZN(n13586) );
  OAI21_X1 U15662 ( .B1(n14244), .B2(n13587), .A(n13586), .ZN(P2_U3299) );
  INV_X1 U15663 ( .A(n13588), .ZN(n14248) );
  OAI222_X1 U15664 ( .A1(n13599), .A2(n13590), .B1(n13587), .B2(n14248), .C1(
        P2_U3088), .C2(n13589), .ZN(P2_U3300) );
  INV_X1 U15665 ( .A(n13591), .ZN(n14252) );
  OAI222_X1 U15666 ( .A1(n13593), .A2(P2_U3088), .B1(n13587), .B2(n14252), 
        .C1(n13592), .C2(n13599), .ZN(P2_U3301) );
  INV_X1 U15667 ( .A(n13594), .ZN(n14256) );
  OAI222_X1 U15668 ( .A1(n13599), .A2(n13596), .B1(n13587), .B2(n14256), .C1(
        n13595), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U15669 ( .A(n13597), .ZN(n13601) );
  INV_X1 U15670 ( .A(n13598), .ZN(n14263) );
  OAI222_X1 U15671 ( .A1(n13601), .A2(P2_U3088), .B1(n13587), .B2(n14263), 
        .C1(n13600), .C2(n13599), .ZN(P2_U3303) );
  INV_X1 U15672 ( .A(n13602), .ZN(n13603) );
  MUX2_X1 U15673 ( .A(n13603), .B(n14767), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3327) );
  NAND2_X1 U15674 ( .A1(n13725), .A2(n13747), .ZN(n13606) );
  NAND2_X1 U15675 ( .A1(n13745), .A2(n6462), .ZN(n13605) );
  NAND2_X1 U15676 ( .A1(n13606), .A2(n13605), .ZN(n13934) );
  AOI22_X1 U15677 ( .A1(n14552), .A2(n13934), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13607) );
  OAI21_X1 U15678 ( .B1(n14557), .B2(n13940), .A(n13607), .ZN(n13608) );
  AOI21_X1 U15679 ( .B1(n13939), .B2(n14554), .A(n13608), .ZN(n13609) );
  OAI21_X1 U15680 ( .B1(n13610), .B2(n13740), .A(n13609), .ZN(P1_U3214) );
  NOR2_X1 U15681 ( .A1(n13612), .A2(n7332), .ZN(n13614) );
  INV_X1 U15682 ( .A(n13613), .ZN(n13678) );
  AOI21_X1 U15683 ( .B1(n13614), .B2(n13699), .A(n13678), .ZN(n13620) );
  OR2_X1 U15684 ( .A1(n13635), .A2(n13711), .ZN(n13616) );
  NAND2_X1 U15685 ( .A1(n13749), .A2(n6462), .ZN(n13615) );
  NAND2_X1 U15686 ( .A1(n13616), .A2(n13615), .ZN(n14137) );
  AOI22_X1 U15687 ( .A1(n14137), .A2(n14552), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13617) );
  OAI21_X1 U15688 ( .B1(n14001), .B2(n14557), .A(n13617), .ZN(n13618) );
  AOI21_X1 U15689 ( .B1(n14212), .B2(n14554), .A(n13618), .ZN(n13619) );
  OAI21_X1 U15690 ( .B1(n13620), .B2(n13740), .A(n13619), .ZN(P1_U3216) );
  AND2_X1 U15691 ( .A1(n13707), .A2(n13622), .ZN(n13625) );
  OAI211_X1 U15692 ( .C1(n13625), .C2(n13624), .A(n14550), .B(n13623), .ZN(
        n13631) );
  NAND2_X1 U15693 ( .A1(n13753), .A2(n6462), .ZN(n13627) );
  OR2_X1 U15694 ( .A1(n13668), .A2(n13711), .ZN(n13626) );
  NAND2_X1 U15695 ( .A1(n13627), .A2(n13626), .ZN(n14057) );
  NOR2_X1 U15696 ( .A1(n14557), .A2(n14059), .ZN(n13628) );
  AOI211_X1 U15697 ( .C1(n14552), .C2(n14057), .A(n13629), .B(n13628), .ZN(
        n13630) );
  OAI211_X1 U15698 ( .C1(n14227), .C2(n13730), .A(n13631), .B(n13630), .ZN(
        P1_U3219) );
  INV_X1 U15699 ( .A(n13632), .ZN(n13698) );
  AOI21_X1 U15700 ( .B1(n13634), .B2(n13633), .A(n13698), .ZN(n13641) );
  OR2_X1 U15701 ( .A1(n13635), .A2(n13713), .ZN(n13637) );
  NAND2_X1 U15702 ( .A1(n13753), .A2(n13725), .ZN(n13636) );
  NAND2_X1 U15703 ( .A1(n13637), .A2(n13636), .ZN(n14156) );
  AOI22_X1 U15704 ( .A1(n14156), .A2(n14552), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13638) );
  OAI21_X1 U15705 ( .B1(n14026), .B2(n14557), .A(n13638), .ZN(n13639) );
  AOI21_X1 U15706 ( .B1(n14220), .B2(n14554), .A(n13639), .ZN(n13640) );
  OAI21_X1 U15707 ( .B1(n13641), .B2(n13740), .A(n13640), .ZN(P1_U3223) );
  AOI22_X1 U15708 ( .A1(n13725), .A2(n13749), .B1(n13747), .B2(n6462), .ZN(
        n13969) );
  INV_X1 U15709 ( .A(n13969), .ZN(n13642) );
  AOI22_X1 U15710 ( .A1(n14552), .A2(n13642), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13643) );
  OAI21_X1 U15711 ( .B1(n14557), .B2(n13965), .A(n13643), .ZN(n13650) );
  INV_X1 U15712 ( .A(n13644), .ZN(n13645) );
  NAND3_X1 U15713 ( .A1(n13679), .A2(n13646), .A3(n13645), .ZN(n13647) );
  AOI21_X1 U15714 ( .B1(n13648), .B2(n13647), .A(n13740), .ZN(n13649) );
  AOI211_X1 U15715 ( .C1(n13972), .C2(n14554), .A(n13650), .B(n13649), .ZN(
        n13651) );
  INV_X1 U15716 ( .A(n13651), .ZN(P1_U3225) );
  INV_X1 U15717 ( .A(n14571), .ZN(n13660) );
  OAI21_X1 U15718 ( .B1(n13653), .B2(n13652), .A(n13661), .ZN(n13654) );
  NAND2_X1 U15719 ( .A1(n13654), .A2(n14550), .ZN(n13659) );
  NOR2_X1 U15720 ( .A1(n14557), .A2(n13655), .ZN(n13656) );
  AOI211_X1 U15721 ( .C1(n14552), .C2(n14570), .A(n13657), .B(n13656), .ZN(
        n13658) );
  OAI211_X1 U15722 ( .C1(n13660), .C2(n13730), .A(n13659), .B(n13658), .ZN(
        P1_U3226) );
  INV_X1 U15723 ( .A(n13661), .ZN(n13664) );
  NOR3_X1 U15724 ( .A1(n13664), .A2(n13663), .A3(n13662), .ZN(n13667) );
  INV_X1 U15725 ( .A(n13665), .ZN(n13666) );
  OAI21_X1 U15726 ( .B1(n13667), .B2(n13666), .A(n14550), .ZN(n13674) );
  OR2_X1 U15727 ( .A1(n13668), .A2(n13713), .ZN(n13670) );
  NAND2_X1 U15728 ( .A1(n13757), .A2(n13725), .ZN(n13669) );
  NAND2_X1 U15729 ( .A1(n13670), .A2(n13669), .ZN(n14095) );
  NOR2_X1 U15730 ( .A1(n13671), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13867) );
  NOR2_X1 U15731 ( .A1(n14557), .A2(n14085), .ZN(n13672) );
  AOI211_X1 U15732 ( .C1(n14552), .C2(n14095), .A(n13867), .B(n13672), .ZN(
        n13673) );
  OAI211_X1 U15733 ( .C1(n14233), .C2(n13730), .A(n13674), .B(n13673), .ZN(
        P1_U3228) );
  INV_X1 U15734 ( .A(n14132), .ZN(n13987) );
  INV_X1 U15735 ( .A(n13675), .ZN(n13677) );
  NOR3_X1 U15736 ( .A1(n13678), .A2(n13677), .A3(n13676), .ZN(n13681) );
  INV_X1 U15737 ( .A(n13679), .ZN(n13680) );
  OAI21_X1 U15738 ( .B1(n13681), .B2(n13680), .A(n14550), .ZN(n13687) );
  INV_X1 U15739 ( .A(n13682), .ZN(n13985) );
  AOI22_X1 U15740 ( .A1(n13725), .A2(n13750), .B1(n13748), .B2(n6462), .ZN(
        n13982) );
  INV_X1 U15741 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13684) );
  OAI22_X1 U15742 ( .A1(n13736), .A2(n13982), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13684), .ZN(n13685) );
  AOI21_X1 U15743 ( .B1(n13985), .B2(n13734), .A(n13685), .ZN(n13686) );
  OAI211_X1 U15744 ( .C1(n13987), .C2(n13730), .A(n13687), .B(n13686), .ZN(
        P1_U3229) );
  XNOR2_X1 U15745 ( .A(n13689), .B(n13688), .ZN(n13695) );
  NOR2_X1 U15746 ( .A1(n14557), .A2(n14044), .ZN(n13693) );
  NOR2_X1 U15747 ( .A1(n13714), .A2(n13711), .ZN(n13690) );
  AOI21_X1 U15748 ( .B1(n13752), .B2(n6462), .A(n13690), .ZN(n14164) );
  OAI22_X1 U15749 ( .A1(n14164), .A2(n13736), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13691), .ZN(n13692) );
  AOI211_X1 U15750 ( .C1(n14043), .C2(n14554), .A(n13693), .B(n13692), .ZN(
        n13694) );
  OAI21_X1 U15751 ( .B1(n13695), .B2(n13740), .A(n13694), .ZN(P1_U3233) );
  NOR3_X1 U15752 ( .A1(n13698), .A2(n7333), .A3(n13697), .ZN(n13701) );
  INV_X1 U15753 ( .A(n13699), .ZN(n13700) );
  OAI21_X1 U15754 ( .B1(n13701), .B2(n13700), .A(n14550), .ZN(n13706) );
  AND2_X1 U15755 ( .A1(n13750), .A2(n6462), .ZN(n13702) );
  AOI21_X1 U15756 ( .B1(n13752), .B2(n13725), .A(n13702), .ZN(n14146) );
  INV_X1 U15757 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13703) );
  OAI22_X1 U15758 ( .A1(n14146), .A2(n13736), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13703), .ZN(n13704) );
  AOI21_X1 U15759 ( .B1(n14012), .B2(n13734), .A(n13704), .ZN(n13705) );
  OAI211_X1 U15760 ( .C1(n13730), .C2(n14217), .A(n13706), .B(n13705), .ZN(
        P1_U3235) );
  OAI21_X1 U15761 ( .B1(n13709), .B2(n13708), .A(n13707), .ZN(n13710) );
  NAND2_X1 U15762 ( .A1(n13710), .A2(n14550), .ZN(n13719) );
  OAI22_X1 U15763 ( .A1(n13714), .A2(n13713), .B1(n13712), .B2(n13711), .ZN(
        n14067) );
  NOR2_X1 U15764 ( .A1(n13715), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13876) );
  INV_X1 U15765 ( .A(n14072), .ZN(n13716) );
  NOR2_X1 U15766 ( .A1(n14557), .A2(n13716), .ZN(n13717) );
  AOI211_X1 U15767 ( .C1(n14552), .C2(n14067), .A(n13876), .B(n13717), .ZN(
        n13718) );
  OAI211_X1 U15768 ( .C1(n14074), .C2(n13730), .A(n13719), .B(n13718), .ZN(
        P1_U3238) );
  OAI21_X1 U15769 ( .B1(n13722), .B2(n13721), .A(n13720), .ZN(n13723) );
  NAND2_X1 U15770 ( .A1(n13723), .A2(n14550), .ZN(n13729) );
  INV_X1 U15771 ( .A(n13724), .ZN(n13948) );
  AOI22_X1 U15772 ( .A1(n13725), .A2(n13748), .B1(n13746), .B2(n6462), .ZN(
        n13954) );
  OAI22_X1 U15773 ( .A1(n13736), .A2(n13954), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13726), .ZN(n13727) );
  AOI21_X1 U15774 ( .B1(n13948), .B2(n13734), .A(n13727), .ZN(n13728) );
  OAI211_X1 U15775 ( .C1(n13950), .C2(n13730), .A(n13729), .B(n13728), .ZN(
        P1_U3240) );
  XNOR2_X1 U15776 ( .A(n13732), .B(n13731), .ZN(n13741) );
  NAND2_X1 U15777 ( .A1(n13734), .A2(n13733), .ZN(n13735) );
  NAND2_X1 U15778 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14638)
         );
  OAI211_X1 U15779 ( .C1(n14577), .C2(n13736), .A(n13735), .B(n14638), .ZN(
        n13737) );
  AOI21_X1 U15780 ( .B1(n13738), .B2(n14554), .A(n13737), .ZN(n13739) );
  OAI21_X1 U15781 ( .B1(n13741), .B2(n13740), .A(n13739), .ZN(P1_U3241) );
  MUX2_X1 U15782 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13742), .S(n13788), .Z(
        P1_U3591) );
  MUX2_X1 U15783 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13743), .S(n13788), .Z(
        P1_U3590) );
  MUX2_X1 U15784 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13744), .S(n13788), .Z(
        P1_U3589) );
  MUX2_X1 U15785 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13745), .S(n13788), .Z(
        P1_U3588) );
  MUX2_X1 U15786 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13746), .S(n13788), .Z(
        P1_U3587) );
  MUX2_X1 U15787 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13747), .S(n13788), .Z(
        P1_U3586) );
  MUX2_X1 U15788 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13748), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15789 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13749), .S(n13788), .Z(
        P1_U3584) );
  MUX2_X1 U15790 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13750), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15791 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13751), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15792 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13752), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15793 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13753), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15794 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13754), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15795 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13755), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15796 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13756), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15797 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13757), .S(n13788), .Z(
        P1_U3576) );
  MUX2_X1 U15798 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13758), .S(n13788), .Z(
        P1_U3575) );
  MUX2_X1 U15799 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13759), .S(n13788), .Z(
        P1_U3574) );
  MUX2_X1 U15800 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13760), .S(n13788), .Z(
        P1_U3573) );
  MUX2_X1 U15801 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13761), .S(n13788), .Z(
        P1_U3572) );
  MUX2_X1 U15802 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13762), .S(n13788), .Z(
        P1_U3571) );
  MUX2_X1 U15803 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13763), .S(n13788), .Z(
        P1_U3570) );
  MUX2_X1 U15804 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13764), .S(n13788), .Z(
        P1_U3569) );
  MUX2_X1 U15805 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13765), .S(n13788), .Z(
        P1_U3568) );
  MUX2_X1 U15806 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13766), .S(n13788), .Z(
        P1_U3567) );
  MUX2_X1 U15807 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13767), .S(n13788), .Z(
        P1_U3566) );
  MUX2_X1 U15808 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13768), .S(n13788), .Z(
        P1_U3565) );
  MUX2_X1 U15809 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13769), .S(n13788), .Z(
        P1_U3564) );
  MUX2_X1 U15810 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13770), .S(n13788), .Z(
        P1_U3563) );
  MUX2_X1 U15811 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13771), .S(n13788), .Z(
        P1_U3562) );
  MUX2_X1 U15812 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13772), .S(n13788), .Z(
        P1_U3561) );
  NAND2_X1 U15813 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13784) );
  OAI211_X1 U15814 ( .C1(n9776), .C2(n13774), .A(n13879), .B(n13773), .ZN(
        n13782) );
  OAI211_X1 U15815 ( .C1(n13777), .C2(n13776), .A(n14631), .B(n13775), .ZN(
        n13781) );
  AOI22_X1 U15816 ( .A1(n13877), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13780) );
  NAND2_X1 U15817 ( .A1(n13855), .A2(n13778), .ZN(n13779) );
  NAND4_X1 U15818 ( .A1(n13782), .A2(n13781), .A3(n13780), .A4(n13779), .ZN(
        P1_U3244) );
  MUX2_X1 U15819 ( .A(n13784), .B(n13783), .S(n14247), .Z(n13789) );
  NAND2_X1 U15820 ( .A1(n13786), .A2(n13785), .ZN(n13787) );
  OAI211_X1 U15821 ( .C1(n13789), .C2(n14245), .A(n13788), .B(n13787), .ZN(
        n13829) );
  OAI22_X1 U15822 ( .A1(n14640), .A2(n14269), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13790), .ZN(n13791) );
  AOI21_X1 U15823 ( .B1(n13792), .B2(n13855), .A(n13791), .ZN(n13802) );
  INV_X1 U15824 ( .A(n13793), .ZN(n13794) );
  XNOR2_X1 U15825 ( .A(n13795), .B(n13794), .ZN(n13796) );
  NAND2_X1 U15826 ( .A1(n13879), .A2(n13796), .ZN(n13801) );
  OAI211_X1 U15827 ( .C1(n13799), .C2(n13798), .A(n14631), .B(n13797), .ZN(
        n13800) );
  NAND4_X1 U15828 ( .A1(n13829), .A2(n13802), .A3(n13801), .A4(n13800), .ZN(
        P1_U3245) );
  OAI211_X1 U15829 ( .C1(n13805), .C2(n13804), .A(n14631), .B(n13803), .ZN(
        n13813) );
  OAI211_X1 U15830 ( .C1(n13807), .C2(n13806), .A(n13879), .B(n13823), .ZN(
        n13812) );
  AND2_X1 U15831 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n13808) );
  AOI21_X1 U15832 ( .B1(n13877), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n13808), .ZN(
        n13811) );
  NAND2_X1 U15833 ( .A1(n13855), .A2(n13809), .ZN(n13810) );
  NAND4_X1 U15834 ( .A1(n13813), .A2(n13812), .A3(n13811), .A4(n13810), .ZN(
        P1_U3246) );
  INV_X1 U15835 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n13815) );
  OAI21_X1 U15836 ( .B1(n14640), .B2(n13815), .A(n13814), .ZN(n13816) );
  AOI21_X1 U15837 ( .B1(n13820), .B2(n13855), .A(n13816), .ZN(n13828) );
  OAI211_X1 U15838 ( .C1(n13819), .C2(n13818), .A(n14631), .B(n13817), .ZN(
        n13827) );
  MUX2_X1 U15839 ( .A(n9780), .B(P1_REG2_REG_4__SCAN_IN), .S(n13820), .Z(
        n13821) );
  NAND3_X1 U15840 ( .A1(n13823), .A2(n13822), .A3(n13821), .ZN(n13824) );
  NAND3_X1 U15841 ( .A1(n13879), .A2(n13825), .A3(n13824), .ZN(n13826) );
  NAND4_X1 U15842 ( .A1(n13829), .A2(n13828), .A3(n13827), .A4(n13826), .ZN(
        P1_U3247) );
  NOR2_X1 U15843 ( .A1(n14636), .A2(n13830), .ZN(n13831) );
  AOI211_X1 U15844 ( .C1(n13877), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n13832), .B(
        n13831), .ZN(n13844) );
  OAI211_X1 U15845 ( .C1(n13835), .C2(n13834), .A(n14631), .B(n13833), .ZN(
        n13843) );
  INV_X1 U15846 ( .A(n13836), .ZN(n13841) );
  NAND3_X1 U15847 ( .A1(n13839), .A2(n13838), .A3(n13837), .ZN(n13840) );
  NAND3_X1 U15848 ( .A1(n13879), .A2(n13841), .A3(n13840), .ZN(n13842) );
  NAND3_X1 U15849 ( .A1(n13844), .A2(n13843), .A3(n13842), .ZN(P1_U3250) );
  OAI21_X1 U15850 ( .B1(n13847), .B2(n13846), .A(n13845), .ZN(n13848) );
  NAND2_X1 U15851 ( .A1(n13848), .A2(n13879), .ZN(n13859) );
  AOI21_X1 U15852 ( .B1(n13877), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n13849), 
        .ZN(n13858) );
  OAI21_X1 U15853 ( .B1(n13852), .B2(n13851), .A(n13850), .ZN(n13853) );
  NAND2_X1 U15854 ( .A1(n13853), .A2(n14631), .ZN(n13857) );
  NAND2_X1 U15855 ( .A1(n13855), .A2(n13854), .ZN(n13856) );
  NAND4_X1 U15856 ( .A1(n13859), .A2(n13858), .A3(n13857), .A4(n13856), .ZN(
        P1_U3255) );
  AOI211_X1 U15857 ( .C1(n13863), .C2(n13862), .A(n13861), .B(n13860), .ZN(
        n13864) );
  INV_X1 U15858 ( .A(n13864), .ZN(n13873) );
  NOR2_X1 U15859 ( .A1(n14636), .A2(n13865), .ZN(n13866) );
  AOI211_X1 U15860 ( .C1(n13877), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n13867), 
        .B(n13866), .ZN(n13872) );
  OAI211_X1 U15861 ( .C1(n13870), .C2(n13869), .A(n13879), .B(n13868), .ZN(
        n13871) );
  NAND3_X1 U15862 ( .A1(n13873), .A2(n13872), .A3(n13871), .ZN(P1_U3260) );
  NOR2_X1 U15863 ( .A1(n14636), .A2(n13874), .ZN(n13875) );
  AOI211_X1 U15864 ( .C1(n13877), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n13876), 
        .B(n13875), .ZN(n13887) );
  OAI211_X1 U15865 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n13880), .A(n13879), 
        .B(n13878), .ZN(n13886) );
  INV_X1 U15866 ( .A(n13881), .ZN(n13884) );
  INV_X1 U15867 ( .A(n13882), .ZN(n13883) );
  OAI211_X1 U15868 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n13884), .A(n14631), 
        .B(n13883), .ZN(n13885) );
  NAND3_X1 U15869 ( .A1(n13887), .A2(n13886), .A3(n13885), .ZN(P1_U3261) );
  NOR2_X1 U15870 ( .A1(n13888), .A2(n14674), .ZN(n14100) );
  NAND2_X1 U15871 ( .A1(n14100), .A2(n14686), .ZN(n13892) );
  OR2_X1 U15872 ( .A1(n13890), .A2(n13889), .ZN(n14099) );
  NOR2_X1 U15873 ( .A1(n6476), .A2(n14099), .ZN(n13897) );
  AOI21_X1 U15874 ( .B1(n6476), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13897), .ZN(
        n13891) );
  OAI211_X1 U15875 ( .C1(n14193), .C2(n14683), .A(n13892), .B(n13891), .ZN(
        P1_U3263) );
  AOI211_X1 U15876 ( .C1(n13895), .C2(n13894), .A(n14674), .B(n13893), .ZN(
        n14104) );
  NAND2_X1 U15877 ( .A1(n14104), .A2(n14686), .ZN(n13899) );
  AND2_X1 U15878 ( .A1(n6476), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n13896) );
  NOR2_X1 U15879 ( .A1(n13897), .A2(n13896), .ZN(n13898) );
  OAI211_X1 U15880 ( .C1(n14197), .C2(n14683), .A(n13899), .B(n13898), .ZN(
        P1_U3264) );
  INV_X1 U15881 ( .A(n13900), .ZN(n13913) );
  OAI22_X1 U15882 ( .A1(n13903), .A2(n13902), .B1(n13901), .B2(n14667), .ZN(
        n13906) );
  NOR2_X1 U15883 ( .A1(n6476), .A2(n13904), .ZN(n13905) );
  AOI211_X1 U15884 ( .C1(n6476), .C2(P1_REG2_REG_29__SCAN_IN), .A(n13906), .B(
        n13905), .ZN(n13907) );
  OAI21_X1 U15885 ( .B1(n14108), .B2(n14683), .A(n13907), .ZN(n13910) );
  NOR2_X1 U15886 ( .A1(n13908), .A2(n14090), .ZN(n13909) );
  AOI211_X1 U15887 ( .C1(n14055), .C2(n13911), .A(n13910), .B(n13909), .ZN(
        n13912) );
  OAI21_X1 U15888 ( .B1(n13913), .B2(n14077), .A(n13912), .ZN(P1_U3356) );
  XNOR2_X1 U15889 ( .A(n13914), .B(n13922), .ZN(n14111) );
  AOI21_X1 U15890 ( .B1(n13915), .B2(n13936), .A(n14674), .ZN(n13917) );
  NAND2_X1 U15891 ( .A1(n13917), .A2(n13916), .ZN(n14110) );
  INV_X1 U15892 ( .A(n14110), .ZN(n13926) );
  OAI22_X1 U15893 ( .A1(n6476), .A2(n14109), .B1(n13918), .B2(n14667), .ZN(
        n13919) );
  AOI21_X1 U15894 ( .B1(P1_REG2_REG_28__SCAN_IN), .B2(n6476), .A(n13919), .ZN(
        n13920) );
  OAI21_X1 U15895 ( .B1(n14199), .B2(n14683), .A(n13920), .ZN(n13925) );
  NOR2_X1 U15896 ( .A1(n14113), .A2(n14077), .ZN(n13924) );
  AOI211_X1 U15897 ( .C1(n14686), .C2(n13926), .A(n13925), .B(n13924), .ZN(
        n13927) );
  OAI21_X1 U15898 ( .B1(n14111), .B2(n14050), .A(n13927), .ZN(P1_U3265) );
  INV_X1 U15899 ( .A(n13928), .ZN(n13929) );
  OAI21_X1 U15900 ( .B1(n13933), .B2(n13932), .A(n13931), .ZN(n13935) );
  NAND2_X1 U15901 ( .A1(n14115), .A2(n14389), .ZN(n13945) );
  INV_X1 U15902 ( .A(n13947), .ZN(n13938) );
  INV_X1 U15903 ( .A(n13936), .ZN(n13937) );
  AOI211_X1 U15904 ( .C1(n13939), .C2(n13938), .A(n14674), .B(n13937), .ZN(
        n14116) );
  NOR2_X1 U15905 ( .A1(n14203), .A2(n14683), .ZN(n13943) );
  OAI22_X1 U15906 ( .A1(n14389), .A2(n13941), .B1(n13940), .B2(n14667), .ZN(
        n13942) );
  AOI211_X1 U15907 ( .C1(n14116), .C2(n14686), .A(n13943), .B(n13942), .ZN(
        n13944) );
  OAI211_X1 U15908 ( .C1(n14114), .C2(n13988), .A(n13945), .B(n13944), .ZN(
        P1_U3266) );
  XNOR2_X1 U15909 ( .A(n13946), .B(n13953), .ZN(n14124) );
  AOI21_X1 U15910 ( .B1(n14120), .B2(n13962), .A(n13947), .ZN(n14121) );
  AOI22_X1 U15911 ( .A1(n6476), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n13948), 
        .B2(n14680), .ZN(n13949) );
  OAI21_X1 U15912 ( .B1(n13950), .B2(n14683), .A(n13949), .ZN(n13958) );
  OAI21_X1 U15913 ( .B1(n13953), .B2(n13952), .A(n13951), .ZN(n13956) );
  INV_X1 U15914 ( .A(n13954), .ZN(n13955) );
  AOI21_X1 U15915 ( .B1(n13956), .B2(n14664), .A(n13955), .ZN(n14123) );
  NOR2_X1 U15916 ( .A1(n14123), .A2(n6476), .ZN(n13957) );
  AOI211_X1 U15917 ( .C1(n14121), .C2(n14025), .A(n13958), .B(n13957), .ZN(
        n13959) );
  OAI21_X1 U15918 ( .B1(n14077), .B2(n14124), .A(n13959), .ZN(P1_U3267) );
  OAI21_X1 U15919 ( .B1(n13968), .B2(n13961), .A(n13960), .ZN(n14125) );
  INV_X1 U15920 ( .A(n13984), .ZN(n13964) );
  INV_X1 U15921 ( .A(n13962), .ZN(n13963) );
  AOI211_X1 U15922 ( .C1(n13972), .C2(n13964), .A(n14674), .B(n13963), .ZN(
        n14127) );
  INV_X1 U15923 ( .A(n14127), .ZN(n13966) );
  OAI22_X1 U15924 ( .A1(n13966), .A2(n14058), .B1(n14667), .B2(n13965), .ZN(
        n13971) );
  AOI21_X1 U15925 ( .B1(n13968), .B2(n13967), .A(n6537), .ZN(n13970) );
  OAI21_X1 U15926 ( .B1(n13970), .B2(n14728), .A(n13969), .ZN(n14126) );
  OAI21_X1 U15927 ( .B1(n13971), .B2(n14126), .A(n14389), .ZN(n13974) );
  AOI22_X1 U15928 ( .A1(n13972), .A2(n14398), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n6476), .ZN(n13973) );
  OAI211_X1 U15929 ( .C1(n14125), .C2(n14077), .A(n13974), .B(n13973), .ZN(
        P1_U3268) );
  INV_X1 U15930 ( .A(n13975), .ZN(n13976) );
  AOI21_X1 U15931 ( .B1(n13980), .B2(n13977), .A(n13976), .ZN(n14135) );
  OAI211_X1 U15932 ( .C1(n13980), .C2(n13979), .A(n13978), .B(n14664), .ZN(
        n13981) );
  OAI211_X1 U15933 ( .C1(n14135), .C2(n14700), .A(n13982), .B(n13981), .ZN(
        n13983) );
  INV_X1 U15934 ( .A(n13983), .ZN(n14134) );
  AOI211_X1 U15935 ( .C1(n14132), .C2(n13997), .A(n14674), .B(n13984), .ZN(
        n14131) );
  AOI22_X1 U15936 ( .A1(n6476), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n13985), 
        .B2(n14680), .ZN(n13986) );
  OAI21_X1 U15937 ( .B1(n13987), .B2(n14683), .A(n13986), .ZN(n13990) );
  NOR2_X1 U15938 ( .A1(n14135), .A2(n13988), .ZN(n13989) );
  AOI211_X1 U15939 ( .C1(n14131), .C2(n14686), .A(n13990), .B(n13989), .ZN(
        n13991) );
  OAI21_X1 U15940 ( .B1(n6476), .B2(n14134), .A(n13991), .ZN(P1_U3269) );
  XNOR2_X1 U15941 ( .A(n13992), .B(n13995), .ZN(n14136) );
  OAI21_X1 U15942 ( .B1(n13995), .B2(n13994), .A(n13993), .ZN(n14140) );
  AOI21_X1 U15943 ( .B1(n14212), .B2(n13996), .A(n14674), .ZN(n13998) );
  NAND2_X1 U15944 ( .A1(n13998), .A2(n13997), .ZN(n14139) );
  NAND2_X1 U15945 ( .A1(n14137), .A2(n14389), .ZN(n14000) );
  NAND2_X1 U15946 ( .A1(n6476), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n13999) );
  OAI211_X1 U15947 ( .C1(n14667), .C2(n14001), .A(n14000), .B(n13999), .ZN(
        n14002) );
  AOI21_X1 U15948 ( .B1(n14212), .B2(n14398), .A(n14002), .ZN(n14003) );
  OAI21_X1 U15949 ( .B1(n14139), .B2(n14090), .A(n14003), .ZN(n14004) );
  AOI21_X1 U15950 ( .B1(n14140), .B2(n14055), .A(n14004), .ZN(n14005) );
  OAI21_X1 U15951 ( .B1(n14077), .B2(n14136), .A(n14005), .ZN(P1_U3270) );
  XNOR2_X1 U15952 ( .A(n14009), .B(n14006), .ZN(n14150) );
  INV_X1 U15953 ( .A(n14150), .ZN(n14019) );
  OAI21_X1 U15954 ( .B1(n14009), .B2(n14008), .A(n14007), .ZN(n14149) );
  INV_X1 U15955 ( .A(n14024), .ZN(n14010) );
  XNOR2_X1 U15956 ( .A(n14217), .B(n14010), .ZN(n14011) );
  NAND2_X1 U15957 ( .A1(n14011), .A2(n14655), .ZN(n14147) );
  INV_X1 U15958 ( .A(n14012), .ZN(n14013) );
  OAI22_X1 U15959 ( .A1(n14146), .A2(n6476), .B1(n14013), .B2(n14667), .ZN(
        n14015) );
  NOR2_X1 U15960 ( .A1(n14217), .A2(n14683), .ZN(n14014) );
  AOI211_X1 U15961 ( .C1(n6476), .C2(P1_REG2_REG_22__SCAN_IN), .A(n14015), .B(
        n14014), .ZN(n14016) );
  OAI21_X1 U15962 ( .B1(n14090), .B2(n14147), .A(n14016), .ZN(n14017) );
  AOI21_X1 U15963 ( .B1(n14677), .B2(n14149), .A(n14017), .ZN(n14018) );
  OAI21_X1 U15964 ( .B1(n14019), .B2(n14050), .A(n14018), .ZN(P1_U3271) );
  XNOR2_X1 U15965 ( .A(n14020), .B(n14021), .ZN(n14160) );
  XNOR2_X1 U15966 ( .A(n14022), .B(n14021), .ZN(n14155) );
  INV_X1 U15967 ( .A(n14220), .ZN(n14031) );
  AND2_X1 U15968 ( .A1(n14220), .A2(n14040), .ZN(n14023) );
  NOR2_X1 U15969 ( .A1(n14024), .A2(n14023), .ZN(n14157) );
  NAND2_X1 U15970 ( .A1(n14157), .A2(n14025), .ZN(n14030) );
  INV_X1 U15971 ( .A(n14156), .ZN(n14027) );
  OAI22_X1 U15972 ( .A1(n14027), .A2(n6476), .B1(n14026), .B2(n14667), .ZN(
        n14028) );
  AOI21_X1 U15973 ( .B1(P1_REG2_REG_21__SCAN_IN), .B2(n6476), .A(n14028), .ZN(
        n14029) );
  OAI211_X1 U15974 ( .C1(n14031), .C2(n14683), .A(n14030), .B(n14029), .ZN(
        n14032) );
  AOI21_X1 U15975 ( .B1(n14155), .B2(n14055), .A(n14032), .ZN(n14033) );
  OAI21_X1 U15976 ( .B1(n14160), .B2(n14077), .A(n14033), .ZN(P1_U3272) );
  OAI21_X1 U15977 ( .B1(n14035), .B2(n14039), .A(n14034), .ZN(n14170) );
  INV_X1 U15978 ( .A(n14036), .ZN(n14037) );
  AOI21_X1 U15979 ( .B1(n14039), .B2(n14038), .A(n14037), .ZN(n14168) );
  INV_X1 U15980 ( .A(n14040), .ZN(n14041) );
  AOI211_X1 U15981 ( .C1(n14043), .C2(n14042), .A(n14674), .B(n14041), .ZN(
        n14167) );
  NAND2_X1 U15982 ( .A1(n14167), .A2(n14686), .ZN(n14047) );
  OAI22_X1 U15983 ( .A1(n14164), .A2(n6476), .B1(n14044), .B2(n14667), .ZN(
        n14045) );
  AOI21_X1 U15984 ( .B1(P1_REG2_REG_20__SCAN_IN), .B2(n6476), .A(n14045), .ZN(
        n14046) );
  OAI211_X1 U15985 ( .C1(n14165), .C2(n14683), .A(n14047), .B(n14046), .ZN(
        n14048) );
  AOI21_X1 U15986 ( .B1(n14677), .B2(n14168), .A(n14048), .ZN(n14049) );
  OAI21_X1 U15987 ( .B1(n14050), .B2(n14170), .A(n14049), .ZN(P1_U3273) );
  XNOR2_X1 U15988 ( .A(n14052), .B(n14051), .ZN(n14173) );
  XNOR2_X1 U15989 ( .A(n14054), .B(n14053), .ZN(n14175) );
  NAND2_X1 U15990 ( .A1(n14175), .A2(n14055), .ZN(n14065) );
  XNOR2_X1 U15991 ( .A(n14227), .B(n14069), .ZN(n14056) );
  NAND2_X1 U15992 ( .A1(n14056), .A2(n14655), .ZN(n14171) );
  INV_X1 U15993 ( .A(n14057), .ZN(n14172) );
  OAI21_X1 U15994 ( .B1(n14171), .B2(n14058), .A(n14172), .ZN(n14063) );
  INV_X1 U15995 ( .A(n14059), .ZN(n14060) );
  AOI22_X1 U15996 ( .A1(n6476), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14060), 
        .B2(n14680), .ZN(n14061) );
  OAI21_X1 U15997 ( .B1(n14227), .B2(n14683), .A(n14061), .ZN(n14062) );
  AOI21_X1 U15998 ( .B1(n14063), .B2(n14389), .A(n14062), .ZN(n14064) );
  OAI211_X1 U15999 ( .C1(n14173), .C2(n14077), .A(n14065), .B(n14064), .ZN(
        P1_U3274) );
  XOR2_X1 U16000 ( .A(n14066), .B(n14076), .Z(n14068) );
  AOI21_X1 U16001 ( .B1(n14068), .B2(n14664), .A(n14067), .ZN(n14181) );
  INV_X1 U16002 ( .A(n14084), .ZN(n14071) );
  INV_X1 U16003 ( .A(n14069), .ZN(n14070) );
  AOI211_X1 U16004 ( .C1(n14179), .C2(n14071), .A(n14674), .B(n14070), .ZN(
        n14178) );
  AOI22_X1 U16005 ( .A1(n6476), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14072), 
        .B2(n14680), .ZN(n14073) );
  OAI21_X1 U16006 ( .B1(n14074), .B2(n14683), .A(n14073), .ZN(n14079) );
  XOR2_X1 U16007 ( .A(n14076), .B(n14075), .Z(n14182) );
  NOR2_X1 U16008 ( .A1(n14182), .A2(n14077), .ZN(n14078) );
  AOI211_X1 U16009 ( .C1(n14178), .C2(n14686), .A(n14079), .B(n14078), .ZN(
        n14080) );
  OAI21_X1 U16010 ( .B1(n6476), .B2(n14181), .A(n14080), .ZN(P1_U3275) );
  XNOR2_X1 U16011 ( .A(n14081), .B(n14091), .ZN(n14183) );
  OAI21_X1 U16012 ( .B1(n14082), .B2(n14233), .A(n14655), .ZN(n14083) );
  OR2_X1 U16013 ( .A1(n14084), .A2(n14083), .ZN(n14185) );
  OAI22_X1 U16014 ( .A1(n14389), .A2(n14086), .B1(n14085), .B2(n14667), .ZN(
        n14087) );
  AOI21_X1 U16015 ( .B1(n14088), .B2(n14398), .A(n14087), .ZN(n14089) );
  OAI21_X1 U16016 ( .B1(n14185), .B2(n14090), .A(n14089), .ZN(n14097) );
  AOI21_X1 U16017 ( .B1(n14092), .B2(n14091), .A(n14728), .ZN(n14094) );
  NAND2_X1 U16018 ( .A1(n14094), .A2(n14093), .ZN(n14186) );
  INV_X1 U16019 ( .A(n14095), .ZN(n14184) );
  AOI21_X1 U16020 ( .B1(n14186), .B2(n14184), .A(n6476), .ZN(n14096) );
  AOI211_X1 U16021 ( .C1(n14183), .C2(n14677), .A(n14097), .B(n14096), .ZN(
        n14098) );
  INV_X1 U16022 ( .A(n14098), .ZN(P1_U3276) );
  INV_X1 U16023 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14101) );
  INV_X1 U16024 ( .A(n14099), .ZN(n14103) );
  NOR2_X1 U16025 ( .A1(n14100), .A2(n14103), .ZN(n14191) );
  NOR2_X1 U16026 ( .A1(n14104), .A2(n14103), .ZN(n14194) );
  MUX2_X1 U16027 ( .A(n14105), .B(n14194), .S(n14766), .Z(n14106) );
  OAI21_X1 U16028 ( .B1(n14197), .B2(n14190), .A(n14106), .ZN(P1_U3558) );
  AND2_X1 U16029 ( .A1(n14110), .A2(n14109), .ZN(n14112) );
  INV_X1 U16030 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n14118) );
  INV_X1 U16031 ( .A(n14114), .ZN(n14117) );
  OAI21_X1 U16032 ( .B1(n14203), .B2(n14190), .A(n14119), .ZN(P1_U3555) );
  AOI22_X1 U16033 ( .A1(n14121), .A2(n14655), .B1(n14120), .B2(n14724), .ZN(
        n14122) );
  OAI211_X1 U16034 ( .C1(n14588), .C2(n14124), .A(n14123), .B(n14122), .ZN(
        n14204) );
  MUX2_X1 U16035 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14204), .S(n14766), .Z(
        P1_U3554) );
  INV_X1 U16036 ( .A(n14125), .ZN(n14128) );
  AOI211_X1 U16037 ( .C1(n14128), .C2(n14753), .A(n14127), .B(n14126), .ZN(
        n14205) );
  MUX2_X1 U16038 ( .A(n14129), .B(n14205), .S(n14766), .Z(n14130) );
  OAI21_X1 U16039 ( .B1(n14208), .B2(n14190), .A(n14130), .ZN(P1_U3553) );
  AOI21_X1 U16040 ( .B1(n14132), .B2(n14724), .A(n14131), .ZN(n14133) );
  OAI211_X1 U16041 ( .C1(n14135), .C2(n14721), .A(n14134), .B(n14133), .ZN(
        n14209) );
  MUX2_X1 U16042 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14209), .S(n14766), .Z(
        P1_U3552) );
  OR2_X1 U16043 ( .A1(n14136), .A2(n14588), .ZN(n14143) );
  INV_X1 U16044 ( .A(n14137), .ZN(n14138) );
  AND2_X1 U16045 ( .A1(n14139), .A2(n14138), .ZN(n14142) );
  NAND2_X1 U16046 ( .A1(n14140), .A2(n14664), .ZN(n14141) );
  NAND3_X1 U16047 ( .A1(n14143), .A2(n14142), .A3(n14141), .ZN(n14210) );
  MUX2_X1 U16048 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14210), .S(n14766), .Z(
        n14144) );
  AOI21_X1 U16049 ( .B1(n14162), .B2(n14212), .A(n14144), .ZN(n14145) );
  INV_X1 U16050 ( .A(n14145), .ZN(P1_U3551) );
  INV_X1 U16051 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n14153) );
  NAND2_X1 U16052 ( .A1(n14147), .A2(n14146), .ZN(n14148) );
  AOI21_X1 U16053 ( .B1(n14149), .B2(n14753), .A(n14148), .ZN(n14152) );
  NAND2_X1 U16054 ( .A1(n14150), .A2(n14664), .ZN(n14151) );
  AND2_X1 U16055 ( .A1(n14152), .A2(n14151), .ZN(n14214) );
  MUX2_X1 U16056 ( .A(n14153), .B(n14214), .S(n14766), .Z(n14154) );
  OAI21_X1 U16057 ( .B1(n14190), .B2(n14217), .A(n14154), .ZN(P1_U3550) );
  NAND2_X1 U16058 ( .A1(n14155), .A2(n14664), .ZN(n14159) );
  AOI21_X1 U16059 ( .B1(n14157), .B2(n14655), .A(n14156), .ZN(n14158) );
  OAI211_X1 U16060 ( .C1(n14160), .C2(n14588), .A(n14159), .B(n14158), .ZN(
        n14218) );
  MUX2_X1 U16061 ( .A(n14218), .B(P1_REG1_REG_21__SCAN_IN), .S(n14764), .Z(
        n14161) );
  AOI21_X1 U16062 ( .B1(n14162), .B2(n14220), .A(n14161), .ZN(n14163) );
  INV_X1 U16063 ( .A(n14163), .ZN(P1_U3549) );
  OAI21_X1 U16064 ( .B1(n14165), .B2(n14749), .A(n14164), .ZN(n14166) );
  AOI211_X1 U16065 ( .C1(n14168), .C2(n14753), .A(n14167), .B(n14166), .ZN(
        n14169) );
  OAI21_X1 U16066 ( .B1(n14728), .B2(n14170), .A(n14169), .ZN(n14223) );
  MUX2_X1 U16067 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14223), .S(n14766), .Z(
        P1_U3548) );
  OAI211_X1 U16068 ( .C1(n14173), .C2(n14588), .A(n14172), .B(n14171), .ZN(
        n14174) );
  AOI21_X1 U16069 ( .B1(n14664), .B2(n14175), .A(n14174), .ZN(n14224) );
  MUX2_X1 U16070 ( .A(n14176), .B(n14224), .S(n14766), .Z(n14177) );
  OAI21_X1 U16071 ( .B1(n14227), .B2(n14190), .A(n14177), .ZN(P1_U3547) );
  AOI21_X1 U16072 ( .B1(n14179), .B2(n14724), .A(n14178), .ZN(n14180) );
  OAI211_X1 U16073 ( .C1(n14588), .C2(n14182), .A(n14181), .B(n14180), .ZN(
        n14228) );
  MUX2_X1 U16074 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14228), .S(n14766), .Z(
        P1_U3546) );
  NAND2_X1 U16075 ( .A1(n14183), .A2(n14753), .ZN(n14188) );
  AND2_X1 U16076 ( .A1(n14185), .A2(n14184), .ZN(n14187) );
  MUX2_X1 U16077 ( .A(n11616), .B(n14230), .S(n14766), .Z(n14189) );
  OAI21_X1 U16078 ( .B1(n14233), .B2(n14190), .A(n14189), .ZN(P1_U3545) );
  MUX2_X1 U16079 ( .A(n14195), .B(n14194), .S(n14756), .Z(n14196) );
  OAI21_X1 U16080 ( .B1(n14197), .B2(n14232), .A(n14196), .ZN(P1_U3526) );
  MUX2_X1 U16081 ( .A(n14201), .B(n14200), .S(n14756), .Z(n14202) );
  OAI21_X1 U16082 ( .B1(n14203), .B2(n14232), .A(n14202), .ZN(P1_U3523) );
  MUX2_X1 U16083 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14204), .S(n14756), .Z(
        P1_U3522) );
  INV_X1 U16084 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n14206) );
  MUX2_X1 U16085 ( .A(n14206), .B(n14205), .S(n14756), .Z(n14207) );
  OAI21_X1 U16086 ( .B1(n14208), .B2(n14232), .A(n14207), .ZN(P1_U3521) );
  MUX2_X1 U16087 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14209), .S(n14756), .Z(
        P1_U3520) );
  MUX2_X1 U16088 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14210), .S(n14756), .Z(
        n14211) );
  AOI21_X1 U16089 ( .B1(n14221), .B2(n14212), .A(n14211), .ZN(n14213) );
  INV_X1 U16090 ( .A(n14213), .ZN(P1_U3519) );
  MUX2_X1 U16091 ( .A(n14215), .B(n14214), .S(n14756), .Z(n14216) );
  OAI21_X1 U16092 ( .B1(n14232), .B2(n14217), .A(n14216), .ZN(P1_U3518) );
  MUX2_X1 U16093 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14218), .S(n14756), .Z(
        n14219) );
  AOI21_X1 U16094 ( .B1(n14221), .B2(n14220), .A(n14219), .ZN(n14222) );
  INV_X1 U16095 ( .A(n14222), .ZN(P1_U3517) );
  MUX2_X1 U16096 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14223), .S(n14756), .Z(
        P1_U3516) );
  INV_X1 U16097 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n14225) );
  MUX2_X1 U16098 ( .A(n14225), .B(n14224), .S(n14756), .Z(n14226) );
  OAI21_X1 U16099 ( .B1(n14227), .B2(n14232), .A(n14226), .ZN(P1_U3515) );
  MUX2_X1 U16100 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14228), .S(n14756), .Z(
        P1_U3513) );
  INV_X1 U16101 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14229) );
  MUX2_X1 U16102 ( .A(n14230), .B(n14229), .S(n14755), .Z(n14231) );
  OAI21_X1 U16103 ( .B1(n14233), .B2(n14232), .A(n14231), .ZN(P1_U3510) );
  NAND3_X1 U16104 ( .A1(n14234), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n14239) );
  NAND2_X1 U16105 ( .A1(n14236), .A2(n14235), .ZN(n14238) );
  NAND2_X1 U16106 ( .A1(n14259), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n14237) );
  OAI211_X1 U16107 ( .C1(n14240), .C2(n14239), .A(n14238), .B(n14237), .ZN(
        P1_U3324) );
  OAI222_X1 U16108 ( .A1(n14258), .A2(n14243), .B1(P1_U3086), .B2(n14242), 
        .C1(n14262), .C2(n14241), .ZN(P1_U3326) );
  OAI222_X1 U16109 ( .A1(n14258), .A2(n14249), .B1(n14262), .B2(n14248), .C1(
        n14247), .C2(P1_U3086), .ZN(P1_U3328) );
  INV_X1 U16110 ( .A(n14250), .ZN(n14253) );
  OAI222_X1 U16111 ( .A1(P1_U3086), .A2(n14253), .B1(n14262), .B2(n14252), 
        .C1(n14251), .C2(n14258), .ZN(P1_U3329) );
  INV_X1 U16112 ( .A(n14254), .ZN(n14255) );
  OAI222_X1 U16113 ( .A1(n14258), .A2(n14257), .B1(n14262), .B2(n14256), .C1(
        P1_U3086), .C2(n14255), .ZN(P1_U3330) );
  AOI22_X1 U16114 ( .A1(n14260), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n14259), .ZN(n14261) );
  OAI21_X1 U16115 ( .B1(n14263), .B2(n14262), .A(n14261), .ZN(P1_U3331) );
  MUX2_X1 U16116 ( .A(n14265), .B(n14264), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U16117 ( .A(n14266), .ZN(n14267) );
  MUX2_X1 U16118 ( .A(n14267), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XOR2_X1 U16119 ( .A(n14343), .B(P1_ADDR_REG_14__SCAN_IN), .Z(n14290) );
  INV_X1 U16120 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14289) );
  XOR2_X1 U16121 ( .A(n14287), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n14340) );
  INV_X1 U16122 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14285) );
  INV_X1 U16123 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15075) );
  XOR2_X1 U16124 ( .A(n15075), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n14331) );
  INV_X1 U16125 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15051) );
  INV_X1 U16126 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14305) );
  XOR2_X1 U16127 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), .Z(
        n14301) );
  NOR2_X1 U16128 ( .A1(n14270), .A2(n7232), .ZN(n14272) );
  NOR2_X1 U16129 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(n14311), .ZN(n14271) );
  NOR2_X1 U16130 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n14315), .ZN(n14274) );
  AND2_X1 U16131 ( .A1(n15010), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n14276) );
  NOR2_X1 U16132 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14277), .ZN(n14279) );
  XNOR2_X1 U16133 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n14277), .ZN(n14323) );
  NOR2_X1 U16134 ( .A1(n14323), .A2(n14324), .ZN(n14278) );
  XOR2_X1 U16135 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), .Z(
        n14296) );
  NOR2_X1 U16136 ( .A1(n14297), .A2(n14296), .ZN(n14280) );
  NAND2_X1 U16137 ( .A1(n14331), .A2(n14330), .ZN(n14281) );
  XNOR2_X1 U16138 ( .A(n14283), .B(P1_ADDR_REG_10__SCAN_IN), .ZN(n14294) );
  NOR2_X1 U16139 ( .A1(n14295), .A2(n14294), .ZN(n14282) );
  XOR2_X1 U16140 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n14335) );
  NOR2_X1 U16141 ( .A1(n14336), .A2(n14335), .ZN(n14284) );
  NAND2_X1 U16142 ( .A1(n14340), .A2(n14339), .ZN(n14286) );
  NAND2_X1 U16143 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14291), .ZN(n14288) );
  XOR2_X1 U16144 ( .A(n14290), .B(n14345), .Z(n14617) );
  XOR2_X1 U16145 ( .A(n14291), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n14293) );
  XNOR2_X1 U16146 ( .A(n14293), .B(n14292), .ZN(n14611) );
  XOR2_X1 U16147 ( .A(n14295), .B(n14294), .Z(n14387) );
  XOR2_X1 U16148 ( .A(n14297), .B(n14296), .Z(n14327) );
  XNOR2_X1 U16149 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n14298), .ZN(n14299) );
  NAND2_X1 U16150 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14299), .ZN(n14314) );
  INV_X1 U16151 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14380) );
  XNOR2_X1 U16152 ( .A(n14301), .B(n14300), .ZN(n14310) );
  XNOR2_X1 U16153 ( .A(n14303), .B(n14302), .ZN(n14306) );
  NAND2_X1 U16154 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14306), .ZN(n14308) );
  AOI21_X1 U16155 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14305), .A(n14304), .ZN(
        n15278) );
  INV_X1 U16156 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15277) );
  NOR2_X1 U16157 ( .A1(n15278), .A2(n15277), .ZN(n15287) );
  XOR2_X1 U16158 ( .A(n14306), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n15286) );
  NAND2_X1 U16159 ( .A1(n15287), .A2(n15286), .ZN(n14307) );
  NAND2_X1 U16160 ( .A1(n14308), .A2(n14307), .ZN(n14309) );
  NAND2_X1 U16161 ( .A1(n14310), .A2(n14309), .ZN(n14377) );
  NOR2_X1 U16162 ( .A1(n14310), .A2(n14309), .ZN(n14378) );
  AOI21_X1 U16163 ( .B1(n14380), .B2(n14377), .A(n14378), .ZN(n15282) );
  XNOR2_X1 U16164 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14311), .ZN(n15283) );
  NOR2_X1 U16165 ( .A1(n15282), .A2(n15283), .ZN(n14312) );
  INV_X1 U16166 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15284) );
  NAND2_X1 U16167 ( .A1(n15282), .A2(n15283), .ZN(n15281) );
  OAI21_X1 U16168 ( .B1(n14312), .B2(n15284), .A(n15281), .ZN(n15273) );
  NAND2_X1 U16169 ( .A1(n15274), .A2(n15273), .ZN(n14313) );
  NAND2_X1 U16170 ( .A1(n14314), .A2(n14313), .ZN(n14317) );
  XNOR2_X1 U16171 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n14315), .ZN(n14316) );
  XNOR2_X1 U16172 ( .A(n14317), .B(n14316), .ZN(n15275) );
  NAND2_X1 U16173 ( .A1(n14318), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14321) );
  XOR2_X1 U16174 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n15010), .Z(n14320) );
  XOR2_X1 U16175 ( .A(n14320), .B(n14319), .Z(n14381) );
  NAND2_X1 U16176 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14322), .ZN(n14325) );
  XOR2_X1 U16177 ( .A(n14324), .B(n14323), .Z(n15279) );
  NOR2_X1 U16178 ( .A1(n14327), .A2(n14326), .ZN(n14329) );
  NOR2_X1 U16179 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n14383), .ZN(n14328) );
  XNOR2_X1 U16180 ( .A(n14331), .B(n14330), .ZN(n14333) );
  NAND2_X1 U16181 ( .A1(n14332), .A2(n14333), .ZN(n14334) );
  XOR2_X1 U16182 ( .A(n14336), .B(n14335), .Z(n14337) );
  NOR2_X1 U16183 ( .A1(n14338), .A2(n14337), .ZN(n14602) );
  XNOR2_X1 U16184 ( .A(n14340), .B(n14339), .ZN(n14607) );
  INV_X1 U16185 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14608) );
  INV_X1 U16186 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14613) );
  AND2_X1 U16187 ( .A1(n14617), .A2(n14616), .ZN(n14342) );
  NOR2_X1 U16188 ( .A1(n14617), .A2(n14616), .ZN(n14615) );
  INV_X1 U16189 ( .A(n14615), .ZN(n14341) );
  XOR2_X1 U16190 ( .A(n14641), .B(P3_ADDR_REG_15__SCAN_IN), .Z(n14346) );
  OR2_X1 U16191 ( .A1(n14343), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n14344) );
  AOI22_X1 U16192 ( .A1(n14345), .A2(n14344), .B1(P1_ADDR_REG_14__SCAN_IN), 
        .B2(n14343), .ZN(n14351) );
  XOR2_X1 U16193 ( .A(n14346), .B(n14351), .Z(n14348) );
  INV_X1 U16194 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14356) );
  XOR2_X1 U16195 ( .A(n14356), .B(P1_ADDR_REG_16__SCAN_IN), .Z(n14352) );
  NAND2_X1 U16196 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14349), .ZN(n14350) );
  AOI22_X1 U16197 ( .A1(n14351), .A2(n14350), .B1(P3_ADDR_REG_15__SCAN_IN), 
        .B2(n14641), .ZN(n14358) );
  XOR2_X1 U16198 ( .A(n14352), .B(n14358), .Z(n14353) );
  NOR2_X1 U16199 ( .A1(n14354), .A2(n14353), .ZN(n14623) );
  NOR2_X1 U16200 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n14622), .ZN(n14355) );
  INV_X1 U16201 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14360) );
  OR2_X1 U16202 ( .A1(n14356), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n14357) );
  AOI22_X1 U16203 ( .A1(n14358), .A2(n14357), .B1(P1_ADDR_REG_16__SCAN_IN), 
        .B2(n14356), .ZN(n14361) );
  XOR2_X1 U16204 ( .A(n14360), .B(n14361), .Z(n14362) );
  XNOR2_X1 U16205 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14362), .ZN(n14414) );
  NAND2_X1 U16206 ( .A1(n14415), .A2(n14414), .ZN(n14359) );
  NOR2_X1 U16207 ( .A1(n14415), .A2(n14414), .ZN(n14413) );
  NAND2_X1 U16208 ( .A1(n14361), .A2(n14360), .ZN(n14364) );
  NAND2_X1 U16209 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14362), .ZN(n14363) );
  NAND2_X1 U16210 ( .A1(n14364), .A2(n14363), .ZN(n14367) );
  INV_X1 U16211 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14370) );
  XOR2_X1 U16212 ( .A(n14370), .B(P1_ADDR_REG_18__SCAN_IN), .Z(n14368) );
  XNOR2_X1 U16213 ( .A(n14367), .B(n14368), .ZN(n14366) );
  NAND2_X1 U16214 ( .A1(n14368), .A2(n14367), .ZN(n14369) );
  OAI21_X1 U16215 ( .B1(n14370), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n14369), 
        .ZN(n14373) );
  XNOR2_X1 U16216 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n14371) );
  XNOR2_X1 U16217 ( .A(n14371), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n14372) );
  XNOR2_X1 U16218 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14374), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16219 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14375) );
  OAI21_X1 U16220 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14375), 
        .ZN(U28) );
  AOI21_X1 U16221 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14376) );
  OAI21_X1 U16222 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14376), 
        .ZN(U29) );
  INV_X1 U16223 ( .A(n14377), .ZN(n14379) );
  AOI222_X1 U16224 ( .A1(n14380), .A2(n14379), .B1(n14380), .B2(n14378), .C1(
        n15282), .C2(n14377), .ZN(SUB_1596_U61) );
  XOR2_X1 U16225 ( .A(n14382), .B(n14381), .Z(SUB_1596_U57) );
  XNOR2_X1 U16226 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14383), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U16227 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14384), .Z(SUB_1596_U54) );
  AOI21_X1 U16228 ( .B1(n14387), .B2(n14386), .A(n14385), .ZN(n14388) );
  XOR2_X1 U16229 ( .A(n14388), .B(P2_ADDR_REG_10__SCAN_IN), .Z(SUB_1596_U70)
         );
  XNOR2_X1 U16230 ( .A(n14390), .B(n7110), .ZN(n14411) );
  XNOR2_X1 U16231 ( .A(n14392), .B(n14391), .ZN(n14393) );
  NOR2_X1 U16232 ( .A1(n14393), .A2(n14728), .ZN(n14394) );
  AOI211_X1 U16233 ( .C1(n14732), .C2(n14411), .A(n14395), .B(n14394), .ZN(
        n14408) );
  INV_X1 U16234 ( .A(n14396), .ZN(n14397) );
  AOI222_X1 U16235 ( .A1(n14399), .A2(n14398), .B1(n14397), .B2(n14680), .C1(
        P1_REG2_REG_12__SCAN_IN), .C2(n6476), .ZN(n14405) );
  INV_X1 U16236 ( .A(n14400), .ZN(n14401) );
  OAI211_X1 U16237 ( .C1(n14407), .C2(n14402), .A(n14401), .B(n14655), .ZN(
        n14406) );
  INV_X1 U16238 ( .A(n14406), .ZN(n14403) );
  AOI22_X1 U16239 ( .A1(n14411), .A2(n14688), .B1(n14686), .B2(n14403), .ZN(
        n14404) );
  OAI211_X1 U16240 ( .C1(n6476), .C2(n14408), .A(n14405), .B(n14404), .ZN(
        P1_U3281) );
  OAI21_X1 U16241 ( .B1(n14407), .B2(n14749), .A(n14406), .ZN(n14410) );
  INV_X1 U16242 ( .A(n14408), .ZN(n14409) );
  AOI211_X1 U16243 ( .C1(n14745), .C2(n14411), .A(n14410), .B(n14409), .ZN(
        n14412) );
  AOI22_X1 U16244 ( .A1(n14756), .A2(n14412), .B1(n7855), .B2(n14755), .ZN(
        P1_U3495) );
  AOI22_X1 U16245 ( .A1(n14766), .A2(n14412), .B1(n10151), .B2(n14764), .ZN(
        P1_U3540) );
  AOI21_X1 U16246 ( .B1(n14415), .B2(n14414), .A(n14413), .ZN(n14416) );
  XOR2_X1 U16247 ( .A(n14416), .B(P2_ADDR_REG_17__SCAN_IN), .Z(SUB_1596_U63)
         );
  OAI211_X1 U16248 ( .C1(n14419), .C2(n14418), .A(n14417), .B(n14960), .ZN(
        n14423) );
  AOI22_X1 U16249 ( .A1(n14421), .A2(n14420), .B1(P3_REG3_REG_14__SCAN_IN), 
        .B2(P3_U3151), .ZN(n14422) );
  OAI211_X1 U16250 ( .C1(n14425), .C2(n14424), .A(n14423), .B(n14422), .ZN(
        n14426) );
  INV_X1 U16251 ( .A(n14426), .ZN(n14427) );
  OAI21_X1 U16252 ( .B1(n14428), .B2(n14971), .A(n14427), .ZN(P3_U3155) );
  NAND2_X1 U16253 ( .A1(n14430), .A2(n14429), .ZN(n14431) );
  NAND2_X1 U16254 ( .A1(n14432), .A2(n14431), .ZN(n14433) );
  AOI222_X1 U16255 ( .A1(n14436), .A2(n14435), .B1(n14434), .B2(n14965), .C1(
        n14433), .C2(n14960), .ZN(n14437) );
  NAND2_X1 U16256 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(P3_U3151), .ZN(n14453)
         );
  OAI211_X1 U16257 ( .C1(n14438), .C2(n14968), .A(n14437), .B(n14453), .ZN(
        P3_U3166) );
  AOI22_X1 U16258 ( .A1(n15056), .A2(n14439), .B1(n15025), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n14455) );
  OAI21_X1 U16259 ( .B1(n14442), .B2(n14441), .A(n14440), .ZN(n14448) );
  NAND2_X1 U16260 ( .A1(n14444), .A2(n14443), .ZN(n14446) );
  XOR2_X1 U16261 ( .A(n14446), .B(n14445), .Z(n14447) );
  AOI22_X1 U16262 ( .A1(n14448), .A2(n15058), .B1(n14478), .B2(n14447), .ZN(
        n14454) );
  OAI221_X1 U16263 ( .B1(n14451), .B2(n14450), .C1(n14451), .C2(n14449), .A(
        n14480), .ZN(n14452) );
  NAND4_X1 U16264 ( .A1(n14455), .A2(n14454), .A3(n14453), .A4(n14452), .ZN(
        P3_U3198) );
  AOI22_X1 U16265 ( .A1(n15056), .A2(n14456), .B1(n15025), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14469) );
  OAI21_X1 U16266 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n14458), .A(n14457), 
        .ZN(n14463) );
  AOI21_X1 U16267 ( .B1(n14460), .B2(n14459), .A(n15067), .ZN(n14462) );
  AOI22_X1 U16268 ( .A1(n14463), .A2(n15058), .B1(n14462), .B2(n14461), .ZN(
        n14468) );
  NAND2_X1 U16269 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_U3151), .ZN(n14467)
         );
  OAI221_X1 U16270 ( .B1(n14465), .B2(n8547), .C1(n14465), .C2(n14464), .A(
        n14480), .ZN(n14466) );
  NAND4_X1 U16271 ( .A1(n14469), .A2(n14468), .A3(n14467), .A4(n14466), .ZN(
        P3_U3199) );
  AOI22_X1 U16272 ( .A1(n15056), .A2(n14470), .B1(n15025), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n14487) );
  OAI21_X1 U16273 ( .B1(n14473), .B2(n14472), .A(n14471), .ZN(n14479) );
  OAI21_X1 U16274 ( .B1(n14476), .B2(n14475), .A(n14474), .ZN(n14477) );
  AOI22_X1 U16275 ( .A1(n14479), .A2(n15058), .B1(n14478), .B2(n14477), .ZN(
        n14486) );
  NAND2_X1 U16276 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(P3_U3151), .ZN(n14485)
         );
  OAI221_X1 U16277 ( .B1(n14483), .B2(n14482), .C1(n14483), .C2(n14481), .A(
        n14480), .ZN(n14484) );
  NAND4_X1 U16278 ( .A1(n14487), .A2(n14486), .A3(n14485), .A4(n14484), .ZN(
        P3_U3200) );
  INV_X1 U16279 ( .A(n14488), .ZN(n15082) );
  NOR2_X1 U16280 ( .A1(n15082), .A2(n14489), .ZN(n14491) );
  OAI21_X1 U16281 ( .B1(n14491), .B2(n14493), .A(n14490), .ZN(n14512) );
  XOR2_X1 U16282 ( .A(n14493), .B(n14492), .Z(n14494) );
  OAI222_X1 U16283 ( .A1(n15185), .A2(n14496), .B1(n15187), .B2(n14495), .C1(
        n14494), .C2(n15130), .ZN(n14510) );
  AOI21_X1 U16284 ( .B1(n15148), .B2(n14512), .A(n14510), .ZN(n14500) );
  NOR2_X1 U16285 ( .A1(n14497), .A2(n15219), .ZN(n14511) );
  AOI22_X1 U16286 ( .A1(n15173), .A2(n14511), .B1(n15203), .B2(n14498), .ZN(
        n14499) );
  OAI221_X1 U16287 ( .B1(n15177), .B2(n14500), .C1(n15204), .C2(n8438), .A(
        n14499), .ZN(P3_U3222) );
  INV_X2 U16288 ( .A(n15270), .ZN(n15269) );
  AOI21_X1 U16289 ( .B1(n14502), .B2(n12811), .A(n14501), .ZN(n14503) );
  AND2_X1 U16290 ( .A1(n14504), .A2(n14503), .ZN(n14514) );
  INV_X1 U16291 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14505) );
  AOI22_X1 U16292 ( .A1(n15269), .A2(n14514), .B1(n14505), .B2(n15270), .ZN(
        P3_U3472) );
  AOI211_X1 U16293 ( .C1(n14508), .C2(n12811), .A(n14507), .B(n14506), .ZN(
        n14515) );
  AOI22_X1 U16294 ( .A1(n15269), .A2(n14515), .B1(n14509), .B2(n15270), .ZN(
        P3_U3471) );
  AOI211_X1 U16295 ( .C1(n12811), .C2(n14512), .A(n14511), .B(n14510), .ZN(
        n14516) );
  INV_X1 U16296 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14513) );
  AOI22_X1 U16297 ( .A1(n15269), .A2(n14516), .B1(n14513), .B2(n15270), .ZN(
        P3_U3470) );
  AOI22_X1 U16298 ( .A1(n15253), .A2(n14514), .B1(n8481), .B2(n15252), .ZN(
        P3_U3429) );
  AOI22_X1 U16299 ( .A1(n15253), .A2(n14515), .B1(n8456), .B2(n15252), .ZN(
        P3_U3426) );
  AOI22_X1 U16300 ( .A1(n15253), .A2(n14516), .B1(n8439), .B2(n15252), .ZN(
        P3_U3423) );
  XNOR2_X1 U16301 ( .A(n14517), .B(n14523), .ZN(n14520) );
  INV_X1 U16302 ( .A(n14518), .ZN(n14519) );
  AOI21_X1 U16303 ( .B1(n14520), .B2(n14860), .A(n14519), .ZN(n14538) );
  AOI222_X1 U16304 ( .A1(n14522), .A2(n14846), .B1(P2_REG2_REG_12__SCAN_IN), 
        .B2(n14873), .C1(n14844), .C2(n14521), .ZN(n14530) );
  XNOR2_X1 U16305 ( .A(n14524), .B(n14523), .ZN(n14541) );
  OAI211_X1 U16306 ( .C1(n14537), .C2(n14527), .A(n14526), .B(n14525), .ZN(
        n14536) );
  INV_X1 U16307 ( .A(n14536), .ZN(n14528) );
  AOI22_X1 U16308 ( .A1(n14541), .A2(n14855), .B1(n14528), .B2(n14854), .ZN(
        n14529) );
  OAI211_X1 U16309 ( .C1(n14873), .C2(n14538), .A(n14530), .B(n14529), .ZN(
        P2_U3253) );
  OAI21_X1 U16310 ( .B1(n6663), .B2(n14928), .A(n14531), .ZN(n14533) );
  AOI211_X1 U16311 ( .C1(n14921), .C2(n14534), .A(n14533), .B(n14532), .ZN(
        n14543) );
  AOI22_X1 U16312 ( .A1(n14535), .A2(n14543), .B1(n10649), .B2(n14951), .ZN(
        P2_U3513) );
  OAI21_X1 U16313 ( .B1(n14537), .B2(n14928), .A(n14536), .ZN(n14540) );
  INV_X1 U16314 ( .A(n14538), .ZN(n14539) );
  AOI211_X1 U16315 ( .C1(n14921), .C2(n14541), .A(n14540), .B(n14539), .ZN(
        n14545) );
  AOI22_X1 U16316 ( .A1(n14954), .A2(n14545), .B1(n10080), .B2(n14951), .ZN(
        P2_U3511) );
  INV_X1 U16317 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14542) );
  AOI22_X1 U16318 ( .A1(n14942), .A2(n14543), .B1(n14542), .B2(n14940), .ZN(
        P2_U3472) );
  INV_X1 U16319 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14544) );
  AOI22_X1 U16320 ( .A1(n14942), .A2(n14545), .B1(n14544), .B2(n14940), .ZN(
        P2_U3466) );
  NAND2_X1 U16321 ( .A1(n14547), .A2(n14546), .ZN(n14548) );
  NAND2_X1 U16322 ( .A1(n14549), .A2(n14548), .ZN(n14551) );
  AOI222_X1 U16323 ( .A1(n14554), .A2(n14558), .B1(n14553), .B2(n14552), .C1(
        n14551), .C2(n14550), .ZN(n14556) );
  OAI211_X1 U16324 ( .C1(n14557), .C2(n14559), .A(n14556), .B(n14555), .ZN(
        P1_U3215) );
  INV_X1 U16325 ( .A(n14558), .ZN(n14561) );
  OAI22_X1 U16326 ( .A1(n14561), .A2(n14560), .B1(n14559), .B2(n14667), .ZN(
        n14563) );
  AOI211_X1 U16327 ( .C1(n14565), .C2(n14564), .A(n14563), .B(n14562), .ZN(
        n14568) );
  AOI22_X1 U16328 ( .A1(n14566), .A2(n14677), .B1(P1_REG2_REG_14__SCAN_IN), 
        .B2(n6476), .ZN(n14567) );
  OAI21_X1 U16329 ( .B1(n6476), .B2(n14568), .A(n14567), .ZN(P1_U3279) );
  AOI211_X1 U16330 ( .C1(n14571), .C2(n14724), .A(n14570), .B(n14569), .ZN(
        n14572) );
  OAI21_X1 U16331 ( .B1(n14573), .B2(n14588), .A(n14572), .ZN(n14574) );
  AOI21_X1 U16332 ( .B1(n14575), .B2(n14664), .A(n14574), .ZN(n14597) );
  AOI22_X1 U16333 ( .A1(n14766), .A2(n14597), .B1(n14576), .B2(n14764), .ZN(
        P1_U3544) );
  OAI211_X1 U16334 ( .C1(n14579), .C2(n14749), .A(n14578), .B(n14577), .ZN(
        n14582) );
  NOR2_X1 U16335 ( .A1(n14580), .A2(n14728), .ZN(n14581) );
  AOI211_X1 U16336 ( .C1(n14753), .C2(n14583), .A(n14582), .B(n14581), .ZN(
        n14598) );
  AOI22_X1 U16337 ( .A1(n14766), .A2(n14598), .B1(n7916), .B2(n14764), .ZN(
        P1_U3543) );
  AOI21_X1 U16338 ( .B1(n14585), .B2(n14724), .A(n14584), .ZN(n14587) );
  OAI211_X1 U16339 ( .C1(n14589), .C2(n14588), .A(n14587), .B(n14586), .ZN(
        n14590) );
  AOI21_X1 U16340 ( .B1(n14591), .B2(n14664), .A(n14590), .ZN(n14599) );
  AOI22_X1 U16341 ( .A1(n14766), .A2(n14599), .B1(n10147), .B2(n14764), .ZN(
        P1_U3541) );
  OAI21_X1 U16342 ( .B1(n14593), .B2(n14749), .A(n14592), .ZN(n14595) );
  AOI211_X1 U16343 ( .C1(n14596), .C2(n14753), .A(n14595), .B(n14594), .ZN(
        n14600) );
  AOI22_X1 U16344 ( .A1(n14766), .A2(n14600), .B1(n9906), .B2(n14764), .ZN(
        P1_U3539) );
  AOI22_X1 U16345 ( .A1(n14756), .A2(n14597), .B1(n7930), .B2(n14755), .ZN(
        P1_U3507) );
  AOI22_X1 U16346 ( .A1(n14756), .A2(n14598), .B1(n7915), .B2(n14755), .ZN(
        P1_U3504) );
  AOI22_X1 U16347 ( .A1(n14756), .A2(n14599), .B1(n7876), .B2(n14755), .ZN(
        P1_U3498) );
  AOI22_X1 U16348 ( .A1(n14756), .A2(n14600), .B1(n7843), .B2(n14755), .ZN(
        P1_U3492) );
  NOR2_X1 U16349 ( .A1(n14602), .A2(n14601), .ZN(n14603) );
  XNOR2_X1 U16350 ( .A(n14604), .B(n14603), .ZN(SUB_1596_U69) );
  OAI21_X1 U16351 ( .B1(n14607), .B2(n14606), .A(n14605), .ZN(n14609) );
  XOR2_X1 U16352 ( .A(n14609), .B(n14608), .Z(SUB_1596_U68) );
  OAI21_X1 U16353 ( .B1(n14612), .B2(n14611), .A(n14610), .ZN(n14614) );
  XOR2_X1 U16354 ( .A(n14614), .B(n14613), .Z(SUB_1596_U67) );
  AOI21_X1 U16355 ( .B1(n14617), .B2(n14616), .A(n14615), .ZN(n14618) );
  XOR2_X1 U16356 ( .A(n14618), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  NOR2_X1 U16357 ( .A1(n14620), .A2(n14619), .ZN(n14621) );
  XNOR2_X1 U16358 ( .A(n7227), .B(n14621), .ZN(SUB_1596_U65) );
  NOR2_X1 U16359 ( .A1(n14623), .A2(n14622), .ZN(n14624) );
  XOR2_X1 U16360 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14624), .Z(SUB_1596_U64)
         );
  AOI21_X1 U16361 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14626), .A(n14625), 
        .ZN(n14628) );
  OR2_X1 U16362 ( .A1(n14628), .A2(n14627), .ZN(n14634) );
  OAI21_X1 U16363 ( .B1(n14630), .B2(n7916), .A(n14629), .ZN(n14632) );
  NAND2_X1 U16364 ( .A1(n14632), .A2(n14631), .ZN(n14633) );
  OAI211_X1 U16365 ( .C1(n14636), .C2(n14635), .A(n14634), .B(n14633), .ZN(
        n14637) );
  INV_X1 U16366 ( .A(n14637), .ZN(n14639) );
  OAI211_X1 U16367 ( .C1(n14641), .C2(n14640), .A(n14639), .B(n14638), .ZN(
        P1_U3258) );
  XNOR2_X1 U16368 ( .A(n14642), .B(n14643), .ZN(n14719) );
  XNOR2_X1 U16369 ( .A(n14644), .B(n14643), .ZN(n14645) );
  NOR2_X1 U16370 ( .A1(n14645), .A2(n14728), .ZN(n14646) );
  AOI211_X1 U16371 ( .C1(n14732), .C2(n14719), .A(n14647), .B(n14646), .ZN(
        n14716) );
  INV_X1 U16372 ( .A(n14648), .ZN(n14715) );
  NOR2_X1 U16373 ( .A1(n14667), .A2(n14649), .ZN(n14650) );
  AOI21_X1 U16374 ( .B1(n6476), .B2(P1_REG2_REG_6__SCAN_IN), .A(n14650), .ZN(
        n14651) );
  OAI21_X1 U16375 ( .B1(n14683), .B2(n14715), .A(n14651), .ZN(n14652) );
  INV_X1 U16376 ( .A(n14652), .ZN(n14659) );
  INV_X1 U16377 ( .A(n14653), .ZN(n14656) );
  OAI211_X1 U16378 ( .C1(n14656), .C2(n14715), .A(n14655), .B(n14654), .ZN(
        n14714) );
  INV_X1 U16379 ( .A(n14714), .ZN(n14657) );
  AOI22_X1 U16380 ( .A1(n14719), .A2(n14688), .B1(n14686), .B2(n14657), .ZN(
        n14658) );
  OAI211_X1 U16381 ( .C1(n6476), .C2(n14716), .A(n14659), .B(n14658), .ZN(
        P1_U3287) );
  XNOR2_X1 U16382 ( .A(n14660), .B(n14661), .ZN(n14665) );
  INV_X1 U16383 ( .A(n14662), .ZN(n14663) );
  AOI21_X1 U16384 ( .B1(n14665), .B2(n14664), .A(n14663), .ZN(n14709) );
  NOR2_X1 U16385 ( .A1(n14667), .A2(n14666), .ZN(n14668) );
  AOI21_X1 U16386 ( .B1(n6476), .B2(P1_REG2_REG_4__SCAN_IN), .A(n14668), .ZN(
        n14669) );
  OAI21_X1 U16387 ( .B1(n14683), .B2(n14708), .A(n14669), .ZN(n14670) );
  INV_X1 U16388 ( .A(n14670), .ZN(n14679) );
  XNOR2_X1 U16389 ( .A(n14672), .B(n14671), .ZN(n14712) );
  AOI211_X1 U16390 ( .C1(n14676), .C2(n14675), .A(n14674), .B(n6700), .ZN(
        n14706) );
  AOI22_X1 U16391 ( .A1(n14677), .A2(n14712), .B1(n14686), .B2(n14706), .ZN(
        n14678) );
  OAI211_X1 U16392 ( .C1(n6476), .C2(n14709), .A(n14679), .B(n14678), .ZN(
        P1_U3289) );
  AOI22_X1 U16393 ( .A1(n6476), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n14680), .ZN(n14681) );
  OAI21_X1 U16394 ( .B1(n14683), .B2(n14682), .A(n14681), .ZN(n14684) );
  INV_X1 U16395 ( .A(n14684), .ZN(n14690) );
  AOI22_X1 U16396 ( .A1(n14688), .A2(n14687), .B1(n14686), .B2(n14685), .ZN(
        n14689) );
  OAI211_X1 U16397 ( .C1(n6476), .C2(n14691), .A(n14690), .B(n14689), .ZN(
        P1_U3291) );
  AND2_X1 U16398 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14694), .ZN(P1_U3294) );
  AND2_X1 U16399 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14694), .ZN(P1_U3295) );
  AND2_X1 U16400 ( .A1(n14694), .A2(P1_D_REG_29__SCAN_IN), .ZN(P1_U3296) );
  AND2_X1 U16401 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14694), .ZN(P1_U3297) );
  AND2_X1 U16402 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14694), .ZN(P1_U3298) );
  AND2_X1 U16403 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14694), .ZN(P1_U3299) );
  AND2_X1 U16404 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14694), .ZN(P1_U3300) );
  AND2_X1 U16405 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14694), .ZN(P1_U3301) );
  AND2_X1 U16406 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14694), .ZN(P1_U3302) );
  AND2_X1 U16407 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14694), .ZN(P1_U3303) );
  AND2_X1 U16408 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14694), .ZN(P1_U3304) );
  AND2_X1 U16409 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14694), .ZN(P1_U3305) );
  AND2_X1 U16410 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14694), .ZN(P1_U3306) );
  AND2_X1 U16411 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14694), .ZN(P1_U3307) );
  AND2_X1 U16412 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14694), .ZN(P1_U3308) );
  NOR2_X1 U16413 ( .A1(n14693), .A2(n14692), .ZN(P1_U3309) );
  AND2_X1 U16414 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14694), .ZN(P1_U3310) );
  AND2_X1 U16415 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14694), .ZN(P1_U3311) );
  AND2_X1 U16416 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14694), .ZN(P1_U3312) );
  AND2_X1 U16417 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14694), .ZN(P1_U3313) );
  AND2_X1 U16418 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14694), .ZN(P1_U3314) );
  AND2_X1 U16419 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14694), .ZN(P1_U3315) );
  AND2_X1 U16420 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14694), .ZN(P1_U3316) );
  AND2_X1 U16421 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14694), .ZN(P1_U3317) );
  AND2_X1 U16422 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14694), .ZN(P1_U3318) );
  AND2_X1 U16423 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14694), .ZN(P1_U3319) );
  AND2_X1 U16424 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14694), .ZN(P1_U3320) );
  AND2_X1 U16425 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14694), .ZN(P1_U3321) );
  AND2_X1 U16426 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14694), .ZN(P1_U3322) );
  AND2_X1 U16427 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14694), .ZN(P1_U3323) );
  AOI22_X1 U16428 ( .A1(n14756), .A2(n14695), .B1(n7672), .B2(n14755), .ZN(
        P1_U3459) );
  INV_X1 U16429 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14696) );
  AOI22_X1 U16430 ( .A1(n14756), .A2(n14697), .B1(n14696), .B2(n14755), .ZN(
        P1_U3462) );
  AOI22_X1 U16431 ( .A1(n14756), .A2(n14698), .B1(n7706), .B2(n14755), .ZN(
        P1_U3465) );
  AOI21_X1 U16432 ( .B1(n14700), .B2(n14721), .A(n14699), .ZN(n14705) );
  OAI211_X1 U16433 ( .C1(n14703), .C2(n14749), .A(n14702), .B(n14701), .ZN(
        n14704) );
  NOR2_X1 U16434 ( .A1(n14705), .A2(n14704), .ZN(n14758) );
  AOI22_X1 U16435 ( .A1(n14756), .A2(n14758), .B1(n7720), .B2(n14755), .ZN(
        P1_U3468) );
  INV_X1 U16436 ( .A(n14706), .ZN(n14707) );
  OAI21_X1 U16437 ( .B1(n14708), .B2(n14749), .A(n14707), .ZN(n14711) );
  INV_X1 U16438 ( .A(n14709), .ZN(n14710) );
  AOI211_X1 U16439 ( .C1(n14712), .C2(n14753), .A(n14711), .B(n14710), .ZN(
        n14759) );
  INV_X1 U16440 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14713) );
  AOI22_X1 U16441 ( .A1(n14756), .A2(n14759), .B1(n14713), .B2(n14755), .ZN(
        P1_U3471) );
  OAI21_X1 U16442 ( .B1(n14715), .B2(n14749), .A(n14714), .ZN(n14718) );
  INV_X1 U16443 ( .A(n14716), .ZN(n14717) );
  AOI211_X1 U16444 ( .C1(n14745), .C2(n14719), .A(n14718), .B(n14717), .ZN(
        n14760) );
  INV_X1 U16445 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14720) );
  AOI22_X1 U16446 ( .A1(n14756), .A2(n14760), .B1(n14720), .B2(n14755), .ZN(
        P1_U3477) );
  NOR2_X1 U16447 ( .A1(n14722), .A2(n14721), .ZN(n14731) );
  AOI21_X1 U16448 ( .B1(n14725), .B2(n14724), .A(n14723), .ZN(n14727) );
  OAI211_X1 U16449 ( .C1(n14729), .C2(n14728), .A(n14727), .B(n14726), .ZN(
        n14730) );
  AOI211_X1 U16450 ( .C1(n14733), .C2(n14732), .A(n14731), .B(n14730), .ZN(
        n14761) );
  AOI22_X1 U16451 ( .A1(n14756), .A2(n14761), .B1(n7780), .B2(n14755), .ZN(
        P1_U3480) );
  OAI21_X1 U16452 ( .B1(n14735), .B2(n14749), .A(n14734), .ZN(n14737) );
  AOI211_X1 U16453 ( .C1(n14738), .C2(n14753), .A(n14737), .B(n14736), .ZN(
        n14762) );
  INV_X1 U16454 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14739) );
  AOI22_X1 U16455 ( .A1(n14756), .A2(n14762), .B1(n14739), .B2(n14755), .ZN(
        P1_U3483) );
  INV_X1 U16456 ( .A(n14740), .ZN(n14744) );
  OAI21_X1 U16457 ( .B1(n7106), .B2(n14749), .A(n14741), .ZN(n14743) );
  AOI211_X1 U16458 ( .C1(n14745), .C2(n14744), .A(n14743), .B(n14742), .ZN(
        n14763) );
  INV_X1 U16459 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14746) );
  AOI22_X1 U16460 ( .A1(n14756), .A2(n14763), .B1(n14746), .B2(n14755), .ZN(
        P1_U3486) );
  INV_X1 U16461 ( .A(n14747), .ZN(n14750) );
  OAI21_X1 U16462 ( .B1(n14750), .B2(n14749), .A(n14748), .ZN(n14752) );
  AOI211_X1 U16463 ( .C1(n14754), .C2(n14753), .A(n14752), .B(n14751), .ZN(
        n14765) );
  AOI22_X1 U16464 ( .A1(n14756), .A2(n14765), .B1(n7826), .B2(n14755), .ZN(
        P1_U3489) );
  AOI22_X1 U16465 ( .A1(n14766), .A2(n14758), .B1(n14757), .B2(n14764), .ZN(
        P1_U3531) );
  AOI22_X1 U16466 ( .A1(n14766), .A2(n14759), .B1(n7726), .B2(n14764), .ZN(
        P1_U3532) );
  AOI22_X1 U16467 ( .A1(n14766), .A2(n14760), .B1(n9804), .B2(n14764), .ZN(
        P1_U3534) );
  AOI22_X1 U16468 ( .A1(n14766), .A2(n14761), .B1(n9807), .B2(n14764), .ZN(
        P1_U3535) );
  AOI22_X1 U16469 ( .A1(n14766), .A2(n14762), .B1(n9810), .B2(n14764), .ZN(
        P1_U3536) );
  AOI22_X1 U16470 ( .A1(n14766), .A2(n14763), .B1(n9794), .B2(n14764), .ZN(
        P1_U3537) );
  AOI22_X1 U16471 ( .A1(n14766), .A2(n14765), .B1(n9903), .B2(n14764), .ZN(
        P1_U3538) );
  NOR2_X1 U16472 ( .A1(n14781), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16473 ( .A1(n14781), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n14780) );
  NAND2_X1 U16474 ( .A1(n14767), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n14772) );
  INV_X1 U16475 ( .A(n14768), .ZN(n14771) );
  INV_X1 U16476 ( .A(n14769), .ZN(n14770) );
  AOI211_X1 U16477 ( .C1(n14772), .C2(n14771), .A(n14770), .B(n14803), .ZN(
        n14773) );
  AOI21_X1 U16478 ( .B1(n14798), .B2(n14774), .A(n14773), .ZN(n14779) );
  OAI211_X1 U16479 ( .C1(n14777), .C2(n14776), .A(n14820), .B(n14775), .ZN(
        n14778) );
  NAND3_X1 U16480 ( .A1(n14780), .A2(n14779), .A3(n14778), .ZN(P2_U3215) );
  AOI22_X1 U16481 ( .A1(n14781), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14793) );
  OAI211_X1 U16482 ( .C1(n14784), .C2(n14783), .A(n14811), .B(n14782), .ZN(
        n14785) );
  INV_X1 U16483 ( .A(n14785), .ZN(n14786) );
  AOI21_X1 U16484 ( .B1(n14818), .B2(n14787), .A(n14786), .ZN(n14792) );
  XOR2_X1 U16485 ( .A(n14789), .B(n14788), .Z(n14790) );
  NAND2_X1 U16486 ( .A1(n14820), .A2(n14790), .ZN(n14791) );
  NAND3_X1 U16487 ( .A1(n14793), .A2(n14792), .A3(n14791), .ZN(P2_U3216) );
  OAI21_X1 U16488 ( .B1(n14796), .B2(n14795), .A(n14794), .ZN(n14802) );
  NAND2_X1 U16489 ( .A1(n14798), .A2(n14797), .ZN(n14801) );
  INV_X1 U16490 ( .A(n14799), .ZN(n14800) );
  OAI211_X1 U16491 ( .C1(n14803), .C2(n14802), .A(n14801), .B(n14800), .ZN(
        n14804) );
  INV_X1 U16492 ( .A(n14804), .ZN(n14809) );
  OAI211_X1 U16493 ( .C1(n14807), .C2(n14806), .A(n14820), .B(n14805), .ZN(
        n14808) );
  OAI211_X1 U16494 ( .C1(n14825), .C2(n15284), .A(n14809), .B(n14808), .ZN(
        P2_U3217) );
  INV_X1 U16495 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15276) );
  OAI211_X1 U16496 ( .C1(n14813), .C2(n14812), .A(n14811), .B(n14810), .ZN(
        n14814) );
  INV_X1 U16497 ( .A(n14814), .ZN(n14815) );
  AOI211_X1 U16498 ( .C1(n14818), .C2(n14817), .A(n14816), .B(n14815), .ZN(
        n14824) );
  OAI211_X1 U16499 ( .C1(n14822), .C2(n14821), .A(n14820), .B(n14819), .ZN(
        n14823) );
  OAI211_X1 U16500 ( .C1(n14825), .C2(n15276), .A(n14824), .B(n14823), .ZN(
        P2_U3219) );
  INV_X1 U16501 ( .A(n14826), .ZN(n14834) );
  INV_X1 U16502 ( .A(n14827), .ZN(n14828) );
  OAI22_X1 U16503 ( .A1(n14871), .A2(n14829), .B1(n14828), .B2(n14865), .ZN(
        n14830) );
  AOI21_X1 U16504 ( .B1(n14846), .B2(n14831), .A(n14830), .ZN(n14832) );
  OAI21_X1 U16505 ( .B1(n14834), .B2(n14833), .A(n14832), .ZN(n14835) );
  AOI21_X1 U16506 ( .B1(n14855), .B2(n14836), .A(n14835), .ZN(n14837) );
  OAI21_X1 U16507 ( .B1(n14873), .B2(n14838), .A(n14837), .ZN(P2_U3258) );
  XNOR2_X1 U16508 ( .A(n14840), .B(n14839), .ZN(n14843) );
  INV_X1 U16509 ( .A(n14841), .ZN(n14842) );
  AOI21_X1 U16510 ( .B1(n14843), .B2(n14860), .A(n14842), .ZN(n14918) );
  XNOR2_X1 U16511 ( .A(n14848), .B(n14847), .ZN(n14922) );
  AOI21_X1 U16512 ( .B1(n14851), .B2(n14850), .A(n14849), .ZN(n14853) );
  AND2_X1 U16513 ( .A1(n14853), .A2(n14852), .ZN(n14915) );
  AOI22_X1 U16514 ( .A1(n14855), .A2(n14922), .B1(n14915), .B2(n14854), .ZN(
        n14856) );
  OAI211_X1 U16515 ( .C1(n14873), .C2(n14918), .A(n14857), .B(n14856), .ZN(
        P2_U3261) );
  NOR2_X1 U16516 ( .A1(n14859), .A2(n14858), .ZN(n14889) );
  NOR2_X1 U16517 ( .A1(n14861), .A2(n14860), .ZN(n14863) );
  OAI21_X1 U16518 ( .B1(n14863), .B2(n14887), .A(n14862), .ZN(n14888) );
  AOI21_X1 U16519 ( .B1(n14889), .B2(n14864), .A(n14888), .ZN(n14872) );
  INV_X1 U16520 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n14866) );
  OAI22_X1 U16521 ( .A1(n14867), .A2(n14887), .B1(n14866), .B2(n14865), .ZN(
        n14868) );
  INV_X1 U16522 ( .A(n14868), .ZN(n14869) );
  OAI221_X1 U16523 ( .B1(n14873), .B2(n14872), .C1(n14871), .C2(n14870), .A(
        n14869), .ZN(P2_U3265) );
  AND2_X1 U16524 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14879), .ZN(P2_U3266) );
  AND2_X1 U16525 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14879), .ZN(P2_U3267) );
  AND2_X1 U16526 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14879), .ZN(P2_U3268) );
  AND2_X1 U16527 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14879), .ZN(P2_U3269) );
  AND2_X1 U16528 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14879), .ZN(P2_U3270) );
  AND2_X1 U16529 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14879), .ZN(P2_U3271) );
  AND2_X1 U16530 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14879), .ZN(P2_U3272) );
  AND2_X1 U16531 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14879), .ZN(P2_U3273) );
  AND2_X1 U16532 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14879), .ZN(P2_U3274) );
  AND2_X1 U16533 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14879), .ZN(P2_U3275) );
  AND2_X1 U16534 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14879), .ZN(P2_U3276) );
  AND2_X1 U16535 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14879), .ZN(P2_U3277) );
  NOR2_X1 U16536 ( .A1(n14882), .A2(n14875), .ZN(P2_U3278) );
  AND2_X1 U16537 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14879), .ZN(P2_U3279) );
  NOR2_X1 U16538 ( .A1(n14882), .A2(n14876), .ZN(P2_U3280) );
  AND2_X1 U16539 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14879), .ZN(P2_U3281) );
  AND2_X1 U16540 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14879), .ZN(P2_U3282) );
  AND2_X1 U16541 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14879), .ZN(P2_U3283) );
  AND2_X1 U16542 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14879), .ZN(P2_U3284) );
  AND2_X1 U16543 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14879), .ZN(P2_U3285) );
  AND2_X1 U16544 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14879), .ZN(P2_U3286) );
  AND2_X1 U16545 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14879), .ZN(P2_U3287) );
  AND2_X1 U16546 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14879), .ZN(P2_U3288) );
  AND2_X1 U16547 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14879), .ZN(P2_U3289) );
  AND2_X1 U16548 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14879), .ZN(P2_U3290) );
  AND2_X1 U16549 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14879), .ZN(P2_U3291) );
  AND2_X1 U16550 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14879), .ZN(P2_U3292) );
  AND2_X1 U16551 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14879), .ZN(P2_U3293) );
  NOR2_X1 U16552 ( .A1(n14882), .A2(n14877), .ZN(P2_U3294) );
  NOR2_X1 U16553 ( .A1(n14882), .A2(n14878), .ZN(P2_U3295) );
  AOI22_X1 U16554 ( .A1(n14882), .A2(n14881), .B1(n14880), .B2(n14879), .ZN(
        P2_U3416) );
  AOI22_X1 U16555 ( .A1(n14886), .A2(n14885), .B1(n14884), .B2(n14883), .ZN(
        P2_U3417) );
  INV_X1 U16556 ( .A(n14887), .ZN(n14891) );
  INV_X1 U16557 ( .A(n10666), .ZN(n14890) );
  AOI211_X1 U16558 ( .C1(n14891), .C2(n14890), .A(n14889), .B(n14888), .ZN(
        n14944) );
  INV_X1 U16559 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14892) );
  AOI22_X1 U16560 ( .A1(n14942), .A2(n14944), .B1(n14892), .B2(n14940), .ZN(
        P2_U3430) );
  INV_X1 U16561 ( .A(n14893), .ZN(n14898) );
  OAI21_X1 U16562 ( .B1(n14928), .B2(n14895), .A(n14894), .ZN(n14897) );
  AOI211_X1 U16563 ( .C1(n14898), .C2(n14921), .A(n14897), .B(n14896), .ZN(
        n14946) );
  INV_X1 U16564 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n14899) );
  AOI22_X1 U16565 ( .A1(n14942), .A2(n14946), .B1(n14899), .B2(n14940), .ZN(
        P2_U3433) );
  INV_X1 U16566 ( .A(n14900), .ZN(n14901) );
  AOI21_X1 U16567 ( .B1(n10666), .B2(n14925), .A(n14901), .ZN(n14906) );
  OAI21_X1 U16568 ( .B1(n14903), .B2(n14928), .A(n14902), .ZN(n14904) );
  NOR3_X1 U16569 ( .A1(n14906), .A2(n14905), .A3(n14904), .ZN(n14947) );
  INV_X1 U16570 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14907) );
  AOI22_X1 U16571 ( .A1(n14942), .A2(n14947), .B1(n14907), .B2(n14940), .ZN(
        P2_U3436) );
  AOI21_X1 U16572 ( .B1(n14909), .B2(n14933), .A(n14908), .ZN(n14911) );
  OAI211_X1 U16573 ( .C1(n14938), .C2(n14912), .A(n14911), .B(n14910), .ZN(
        n14913) );
  INV_X1 U16574 ( .A(n14913), .ZN(n14948) );
  INV_X1 U16575 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14914) );
  AOI22_X1 U16576 ( .A1(n14942), .A2(n14948), .B1(n14914), .B2(n14940), .ZN(
        P2_U3439) );
  INV_X1 U16577 ( .A(n14915), .ZN(n14916) );
  OAI21_X1 U16578 ( .B1(n14917), .B2(n14928), .A(n14916), .ZN(n14920) );
  INV_X1 U16579 ( .A(n14918), .ZN(n14919) );
  AOI211_X1 U16580 ( .C1(n14922), .C2(n14921), .A(n14920), .B(n14919), .ZN(
        n14949) );
  INV_X1 U16581 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14923) );
  AOI22_X1 U16582 ( .A1(n14942), .A2(n14949), .B1(n14923), .B2(n14940), .ZN(
        P2_U3442) );
  AOI21_X1 U16583 ( .B1(n10666), .B2(n14925), .A(n14924), .ZN(n14930) );
  OAI211_X1 U16584 ( .C1(n7200), .C2(n14928), .A(n14927), .B(n14926), .ZN(
        n14929) );
  NOR2_X1 U16585 ( .A1(n14930), .A2(n14929), .ZN(n14950) );
  INV_X1 U16586 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14931) );
  AOI22_X1 U16587 ( .A1(n14942), .A2(n14950), .B1(n14931), .B2(n14940), .ZN(
        P2_U3445) );
  AOI21_X1 U16588 ( .B1(n14934), .B2(n14933), .A(n14932), .ZN(n14935) );
  OAI211_X1 U16589 ( .C1(n14938), .C2(n14937), .A(n14936), .B(n14935), .ZN(
        n14939) );
  INV_X1 U16590 ( .A(n14939), .ZN(n14953) );
  INV_X1 U16591 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n14941) );
  AOI22_X1 U16592 ( .A1(n14942), .A2(n14953), .B1(n14941), .B2(n14940), .ZN(
        P2_U3448) );
  AOI22_X1 U16593 ( .A1(n14954), .A2(n14944), .B1(n14943), .B2(n14951), .ZN(
        P2_U3499) );
  INV_X1 U16594 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n14945) );
  AOI22_X1 U16595 ( .A1(n14954), .A2(n14946), .B1(n14945), .B2(n14951), .ZN(
        P2_U3500) );
  AOI22_X1 U16596 ( .A1(n14954), .A2(n14947), .B1(n9856), .B2(n14951), .ZN(
        P2_U3501) );
  AOI22_X1 U16597 ( .A1(n14954), .A2(n14948), .B1(n9862), .B2(n14951), .ZN(
        P2_U3502) );
  AOI22_X1 U16598 ( .A1(n14954), .A2(n14949), .B1(n9865), .B2(n14951), .ZN(
        P2_U3503) );
  AOI22_X1 U16599 ( .A1(n14954), .A2(n14950), .B1(n9867), .B2(n14951), .ZN(
        P2_U3504) );
  AOI22_X1 U16600 ( .A1(n14954), .A2(n14953), .B1(n14952), .B2(n14951), .ZN(
        P2_U3505) );
  NOR2_X1 U16601 ( .A1(P3_U3897), .A2(n15025), .ZN(P3_U3150) );
  INV_X1 U16602 ( .A(n15081), .ZN(n14972) );
  AOI22_X1 U16603 ( .A1(n14956), .A2(n15142), .B1(n15145), .B2(n14955), .ZN(
        n15079) );
  AND2_X1 U16604 ( .A1(n14958), .A2(n14957), .ZN(n14962) );
  OAI211_X1 U16605 ( .C1(n14962), .C2(n14961), .A(n14959), .B(n14960), .ZN(
        n14967) );
  AOI22_X1 U16606 ( .A1(n14965), .A2(n14964), .B1(P3_REG3_REG_10__SCAN_IN), 
        .B2(P3_U3151), .ZN(n14966) );
  OAI211_X1 U16607 ( .C1(n15079), .C2(n14968), .A(n14967), .B(n14966), .ZN(
        n14969) );
  INV_X1 U16608 ( .A(n14969), .ZN(n14970) );
  OAI21_X1 U16609 ( .B1(n14972), .B2(n14971), .A(n14970), .ZN(P3_U3157) );
  AOI21_X1 U16610 ( .B1(n14974), .B2(n15175), .A(n14973), .ZN(n14979) );
  OAI21_X1 U16611 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n14976), .A(n14975), .ZN(
        n14977) );
  NAND2_X1 U16612 ( .A1(n15058), .A2(n14977), .ZN(n14978) );
  OAI21_X1 U16613 ( .B1(n15061), .B2(n14979), .A(n14978), .ZN(n14986) );
  INV_X1 U16614 ( .A(n15003), .ZN(n14983) );
  AOI21_X1 U16615 ( .B1(n14981), .B2(n15002), .A(n14980), .ZN(n14982) );
  AOI21_X1 U16616 ( .B1(n14983), .B2(n15002), .A(n14982), .ZN(n14984) );
  NOR2_X1 U16617 ( .A1(n14984), .A2(n15067), .ZN(n14985) );
  AOI211_X1 U16618 ( .C1(n15056), .C2(n14987), .A(n14986), .B(n14985), .ZN(
        n14989) );
  NAND2_X1 U16619 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(P3_U3151), .ZN(n14988) );
  OAI211_X1 U16620 ( .C1(n14990), .C2(n15074), .A(n14989), .B(n14988), .ZN(
        P3_U3187) );
  AOI21_X1 U16621 ( .B1(n14993), .B2(n14992), .A(n14991), .ZN(n14999) );
  AOI21_X1 U16622 ( .B1(n14996), .B2(n14995), .A(n14994), .ZN(n14997) );
  OAI22_X1 U16623 ( .A1(n14999), .A2(n15061), .B1(n14998), .B2(n14997), .ZN(
        n15006) );
  INV_X1 U16624 ( .A(n15000), .ZN(n15001) );
  NAND3_X1 U16625 ( .A1(n15003), .A2(n15002), .A3(n15001), .ZN(n15004) );
  AOI21_X1 U16626 ( .B1(n15018), .B2(n15004), .A(n15067), .ZN(n15005) );
  AOI211_X1 U16627 ( .C1(n15056), .C2(n15007), .A(n15006), .B(n15005), .ZN(
        n15009) );
  NAND2_X1 U16628 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n15008) );
  OAI211_X1 U16629 ( .C1(n15010), .C2(n15074), .A(n15009), .B(n15008), .ZN(
        P3_U3188) );
  AOI21_X1 U16630 ( .B1(n11125), .B2(n15012), .A(n15011), .ZN(n15031) );
  NOR2_X1 U16631 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15013), .ZN(n15024) );
  INV_X1 U16632 ( .A(n15014), .ZN(n15015) );
  NOR2_X1 U16633 ( .A1(n15016), .A2(n15015), .ZN(n15019) );
  INV_X1 U16634 ( .A(n15035), .ZN(n15017) );
  AOI21_X1 U16635 ( .B1(n15019), .B2(n15018), .A(n15017), .ZN(n15022) );
  OAI22_X1 U16636 ( .A1(n15022), .A2(n15067), .B1(n15021), .B2(n15020), .ZN(
        n15023) );
  AOI211_X1 U16637 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n15025), .A(n15024), .B(
        n15023), .ZN(n15030) );
  OAI21_X1 U16638 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n15027), .A(n15026), .ZN(
        n15028) );
  NAND2_X1 U16639 ( .A1(n15028), .A2(n15058), .ZN(n15029) );
  OAI211_X1 U16640 ( .C1(n15031), .C2(n15061), .A(n15030), .B(n15029), .ZN(
        P3_U3189) );
  INV_X1 U16641 ( .A(n15032), .ZN(n15033) );
  NAND3_X1 U16642 ( .A1(n15035), .A2(n15034), .A3(n15033), .ZN(n15036) );
  AOI21_X1 U16643 ( .B1(n15066), .B2(n15036), .A(n15067), .ZN(n15048) );
  AOI21_X1 U16644 ( .B1(n15039), .B2(n15038), .A(n15037), .ZN(n15046) );
  OAI21_X1 U16645 ( .B1(n15042), .B2(n15041), .A(n15040), .ZN(n15044) );
  AOI22_X1 U16646 ( .A1(n15044), .A2(n15058), .B1(n15043), .B2(n15056), .ZN(
        n15045) );
  OAI21_X1 U16647 ( .B1(n15046), .B2(n15061), .A(n15045), .ZN(n15047) );
  NOR2_X1 U16648 ( .A1(n15048), .A2(n15047), .ZN(n15050) );
  NAND2_X1 U16649 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n15049) );
  OAI211_X1 U16650 ( .C1(n15051), .C2(n15074), .A(n15050), .B(n15049), .ZN(
        P3_U3190) );
  AOI21_X1 U16651 ( .B1(n15053), .B2(n15098), .A(n15052), .ZN(n15062) );
  OAI21_X1 U16652 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n15055), .A(n15054), .ZN(
        n15059) );
  AOI22_X1 U16653 ( .A1(n15059), .A2(n15058), .B1(n15057), .B2(n15056), .ZN(
        n15060) );
  OAI21_X1 U16654 ( .B1(n15062), .B2(n15061), .A(n15060), .ZN(n15071) );
  INV_X1 U16655 ( .A(n15063), .ZN(n15064) );
  NAND3_X1 U16656 ( .A1(n15066), .A2(n15065), .A3(n15064), .ZN(n15068) );
  AOI21_X1 U16657 ( .B1(n15069), .B2(n15068), .A(n15067), .ZN(n15070) );
  NOR2_X1 U16658 ( .A1(n15071), .A2(n15070), .ZN(n15073) );
  NAND2_X1 U16659 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(P3_U3151), .ZN(n15072) );
  OAI211_X1 U16660 ( .C1(n15075), .C2(n15074), .A(n15073), .B(n15072), .ZN(
        P3_U3191) );
  NAND3_X1 U16661 ( .A1(n15091), .A2(n7384), .A3(n15076), .ZN(n15077) );
  NAND3_X1 U16662 ( .A1(n15078), .A2(n15183), .A3(n15077), .ZN(n15080) );
  AOI22_X1 U16663 ( .A1(n15177), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n15203), 
        .B2(n15081), .ZN(n15088) );
  AOI21_X1 U16664 ( .B1(n15084), .B2(n15083), .A(n15082), .ZN(n15251) );
  NOR2_X1 U16665 ( .A1(n15085), .A2(n15219), .ZN(n15250) );
  AOI22_X1 U16666 ( .A1(n15251), .A2(n15086), .B1(n15173), .B2(n15250), .ZN(
        n15087) );
  OAI211_X1 U16667 ( .C1(n15177), .C2(n15248), .A(n15088), .B(n15087), .ZN(
        P3_U3223) );
  XNOR2_X1 U16668 ( .A(n15089), .B(n15094), .ZN(n15244) );
  INV_X1 U16669 ( .A(n15244), .ZN(n15097) );
  INV_X1 U16670 ( .A(n15090), .ZN(n15096) );
  INV_X1 U16671 ( .A(n15091), .ZN(n15092) );
  AOI211_X1 U16672 ( .C1(n15094), .C2(n15093), .A(n15130), .B(n15092), .ZN(
        n15095) );
  AOI211_X1 U16673 ( .C1(n15194), .C2(n15244), .A(n15096), .B(n15095), .ZN(
        n15246) );
  OAI21_X1 U16674 ( .B1(n15097), .B2(n15200), .A(n15246), .ZN(n15102) );
  OAI22_X1 U16675 ( .A1(n15100), .A2(n15099), .B1(n15098), .B2(n15204), .ZN(
        n15101) );
  AOI21_X1 U16676 ( .B1(n15102), .B2(n15204), .A(n15101), .ZN(n15103) );
  OAI21_X1 U16677 ( .B1(n15105), .B2(n15104), .A(n15103), .ZN(P3_U3224) );
  OAI21_X1 U16678 ( .B1(n15107), .B2(n15110), .A(n15106), .ZN(n15239) );
  XOR2_X1 U16679 ( .A(n15110), .B(n15109), .Z(n15115) );
  OAI22_X1 U16680 ( .A1(n15112), .A2(n15185), .B1(n15111), .B2(n15187), .ZN(
        n15113) );
  AOI21_X1 U16681 ( .B1(n15239), .B2(n15194), .A(n15113), .ZN(n15114) );
  OAI21_X1 U16682 ( .B1(n15115), .B2(n15130), .A(n15114), .ZN(n15237) );
  AOI21_X1 U16683 ( .B1(n15170), .B2(n15239), .A(n15237), .ZN(n15119) );
  NOR2_X1 U16684 ( .A1(n15116), .A2(n15219), .ZN(n15238) );
  AOI22_X1 U16685 ( .A1(n15173), .A2(n15238), .B1(n15203), .B2(n15117), .ZN(
        n15118) );
  OAI221_X1 U16686 ( .B1(n15177), .B2(n15119), .C1(n15204), .C2(n11131), .A(
        n15118), .ZN(P3_U3225) );
  OAI21_X1 U16687 ( .B1(n15122), .B2(n15121), .A(n15120), .ZN(n15236) );
  NAND2_X1 U16688 ( .A1(n15123), .A2(n15159), .ZN(n15137) );
  OR2_X1 U16689 ( .A1(n15137), .A2(n15138), .ZN(n15139) );
  NAND2_X1 U16690 ( .A1(n15139), .A2(n15124), .ZN(n15126) );
  XNOR2_X1 U16691 ( .A(n15126), .B(n15125), .ZN(n15131) );
  OAI22_X1 U16692 ( .A1(n15127), .A2(n15185), .B1(n15163), .B2(n15187), .ZN(
        n15128) );
  AOI21_X1 U16693 ( .B1(n15236), .B2(n15194), .A(n15128), .ZN(n15129) );
  OAI21_X1 U16694 ( .B1(n15131), .B2(n15130), .A(n15129), .ZN(n15234) );
  AOI21_X1 U16695 ( .B1(n15170), .B2(n15236), .A(n15234), .ZN(n15135) );
  NOR2_X1 U16696 ( .A1(n15132), .A2(n15219), .ZN(n15235) );
  AOI22_X1 U16697 ( .A1(n15235), .A2(n15173), .B1(n15133), .B2(n15203), .ZN(
        n15134) );
  OAI221_X1 U16698 ( .B1(n15177), .B2(n15135), .C1(n15204), .C2(n11125), .A(
        n15134), .ZN(P3_U3226) );
  XNOR2_X1 U16699 ( .A(n15136), .B(n15138), .ZN(n15233) );
  INV_X1 U16700 ( .A(n15137), .ZN(n15141) );
  INV_X1 U16701 ( .A(n15138), .ZN(n15140) );
  OAI211_X1 U16702 ( .C1(n15141), .C2(n15140), .A(n15183), .B(n15139), .ZN(
        n15147) );
  AOI22_X1 U16703 ( .A1(n15145), .A2(n15144), .B1(n15143), .B2(n15142), .ZN(
        n15146) );
  NAND2_X1 U16704 ( .A1(n15147), .A2(n15146), .ZN(n15231) );
  AOI21_X1 U16705 ( .B1(n15233), .B2(n15148), .A(n15231), .ZN(n15152) );
  AND2_X1 U16706 ( .A1(n15149), .A2(n15242), .ZN(n15232) );
  AOI22_X1 U16707 ( .A1(n15173), .A2(n15232), .B1(n15203), .B2(n15150), .ZN(
        n15151) );
  OAI221_X1 U16708 ( .B1(n15177), .B2(n15152), .C1(n15204), .C2(n11118), .A(
        n15151), .ZN(P3_U3227) );
  XNOR2_X1 U16709 ( .A(n15153), .B(n15161), .ZN(n15168) );
  INV_X1 U16710 ( .A(n15168), .ZN(n15230) );
  NAND2_X1 U16711 ( .A1(n15155), .A2(n15154), .ZN(n15157) );
  NAND2_X1 U16712 ( .A1(n15157), .A2(n15156), .ZN(n15162) );
  AND2_X1 U16713 ( .A1(n15159), .A2(n15158), .ZN(n15160) );
  OAI21_X1 U16714 ( .B1(n15162), .B2(n15161), .A(n15160), .ZN(n15166) );
  OAI22_X1 U16715 ( .A1(n15164), .A2(n15187), .B1(n15163), .B2(n15185), .ZN(
        n15165) );
  AOI21_X1 U16716 ( .B1(n15166), .B2(n15183), .A(n15165), .ZN(n15167) );
  OAI21_X1 U16717 ( .B1(n15169), .B2(n15168), .A(n15167), .ZN(n15228) );
  AOI21_X1 U16718 ( .B1(n15170), .B2(n15230), .A(n15228), .ZN(n15176) );
  AND2_X1 U16719 ( .A1(n15171), .A2(n15242), .ZN(n15229) );
  AOI22_X1 U16720 ( .A1(n15173), .A2(n15229), .B1(n15203), .B2(n15172), .ZN(
        n15174) );
  OAI221_X1 U16721 ( .B1(n15177), .B2(n15176), .C1(n15204), .C2(n15175), .A(
        n15174), .ZN(P3_U3228) );
  NAND2_X1 U16722 ( .A1(n15179), .A2(n15178), .ZN(n15182) );
  NAND2_X1 U16723 ( .A1(n15182), .A2(n15181), .ZN(n15180) );
  OAI21_X1 U16724 ( .B1(n15182), .B2(n15181), .A(n15180), .ZN(n15184) );
  NAND2_X1 U16725 ( .A1(n15184), .A2(n15183), .ZN(n15197) );
  OAI22_X1 U16726 ( .A1(n15188), .A2(n15187), .B1(n15186), .B2(n15185), .ZN(
        n15189) );
  INV_X1 U16727 ( .A(n15189), .ZN(n15196) );
  OR2_X1 U16728 ( .A1(n15191), .A2(n15190), .ZN(n15192) );
  NAND2_X1 U16729 ( .A1(n15193), .A2(n15192), .ZN(n15211) );
  NAND2_X1 U16730 ( .A1(n15211), .A2(n15194), .ZN(n15195) );
  NAND3_X1 U16731 ( .A1(n15197), .A2(n15196), .A3(n15195), .ZN(n15215) );
  INV_X1 U16732 ( .A(n15211), .ZN(n15201) );
  NAND2_X1 U16733 ( .A1(n15198), .A2(n15242), .ZN(n15212) );
  OAI22_X1 U16734 ( .A1(n15201), .A2(n15200), .B1(n15199), .B2(n15212), .ZN(
        n15202) );
  AOI211_X1 U16735 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15203), .A(n15215), .B(
        n15202), .ZN(n15205) );
  AOI22_X1 U16736 ( .A1(n15177), .A2(n15206), .B1(n15205), .B2(n15204), .ZN(
        P3_U3231) );
  INV_X1 U16737 ( .A(n15207), .ZN(n15210) );
  AOI211_X1 U16738 ( .C1(n15243), .C2(n15210), .A(n15209), .B(n15208), .ZN(
        n15254) );
  AOI22_X1 U16739 ( .A1(n15253), .A2(n15254), .B1(n8292), .B2(n15252), .ZN(
        P3_U3393) );
  NAND2_X1 U16740 ( .A1(n15211), .A2(n15243), .ZN(n15213) );
  NAND2_X1 U16741 ( .A1(n15213), .A2(n15212), .ZN(n15214) );
  NOR2_X1 U16742 ( .A1(n15215), .A2(n15214), .ZN(n15256) );
  INV_X1 U16743 ( .A(n15256), .ZN(n15216) );
  OAI22_X1 U16744 ( .A1(n15252), .A2(n15216), .B1(P3_REG0_REG_2__SCAN_IN), 
        .B2(n15253), .ZN(n15217) );
  INV_X1 U16745 ( .A(n15217), .ZN(P3_U3396) );
  INV_X1 U16746 ( .A(n15218), .ZN(n15222) );
  NOR2_X1 U16747 ( .A1(n6719), .A2(n15219), .ZN(n15221) );
  AOI211_X1 U16748 ( .C1(n15222), .C2(n15243), .A(n15221), .B(n15220), .ZN(
        n15258) );
  AOI22_X1 U16749 ( .A1(n15253), .A2(n15258), .B1(n8312), .B2(n15252), .ZN(
        P3_U3399) );
  AOI22_X1 U16750 ( .A1(n15224), .A2(n15243), .B1(n15242), .B2(n15223), .ZN(
        n15225) );
  AND2_X1 U16751 ( .A1(n15226), .A2(n15225), .ZN(n15260) );
  INV_X1 U16752 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15227) );
  AOI22_X1 U16753 ( .A1(n15253), .A2(n15260), .B1(n15227), .B2(n15252), .ZN(
        P3_U3402) );
  AOI211_X1 U16754 ( .C1(n15230), .C2(n15243), .A(n15229), .B(n15228), .ZN(
        n15262) );
  AOI22_X1 U16755 ( .A1(n15253), .A2(n15262), .B1(n8345), .B2(n15252), .ZN(
        P3_U3405) );
  AOI211_X1 U16756 ( .C1(n15233), .C2(n12811), .A(n15232), .B(n15231), .ZN(
        n15264) );
  AOI22_X1 U16757 ( .A1(n15253), .A2(n15264), .B1(n8364), .B2(n15252), .ZN(
        P3_U3408) );
  AOI211_X1 U16758 ( .C1(n15243), .C2(n15236), .A(n15235), .B(n15234), .ZN(
        n15265) );
  AOI22_X1 U16759 ( .A1(n15253), .A2(n15265), .B1(n8378), .B2(n15252), .ZN(
        P3_U3411) );
  AOI211_X1 U16760 ( .C1(n15243), .C2(n15239), .A(n15238), .B(n15237), .ZN(
        n15267) );
  INV_X1 U16761 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15240) );
  AOI22_X1 U16762 ( .A1(n15253), .A2(n15267), .B1(n15240), .B2(n15252), .ZN(
        P3_U3414) );
  AOI22_X1 U16763 ( .A1(n15244), .A2(n15243), .B1(n15242), .B2(n15241), .ZN(
        n15245) );
  AND2_X1 U16764 ( .A1(n15246), .A2(n15245), .ZN(n15268) );
  INV_X1 U16765 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15247) );
  AOI22_X1 U16766 ( .A1(n15253), .A2(n15268), .B1(n15247), .B2(n15252), .ZN(
        P3_U3417) );
  INV_X1 U16767 ( .A(n15248), .ZN(n15249) );
  AOI211_X1 U16768 ( .C1(n15251), .C2(n12811), .A(n15250), .B(n15249), .ZN(
        n15272) );
  AOI22_X1 U16769 ( .A1(n15253), .A2(n15272), .B1(n8422), .B2(n15252), .ZN(
        P3_U3420) );
  AOI22_X1 U16770 ( .A1(n15269), .A2(n15254), .B1(n10477), .B2(n15270), .ZN(
        P3_U3460) );
  AOI22_X1 U16771 ( .A1(n15269), .A2(n15256), .B1(n15255), .B2(n15270), .ZN(
        P3_U3461) );
  INV_X1 U16772 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15257) );
  AOI22_X1 U16773 ( .A1(n15269), .A2(n15258), .B1(n15257), .B2(n15270), .ZN(
        P3_U3462) );
  AOI22_X1 U16774 ( .A1(n15269), .A2(n15260), .B1(n15259), .B2(n15270), .ZN(
        P3_U3463) );
  INV_X1 U16775 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15261) );
  AOI22_X1 U16776 ( .A1(n15269), .A2(n15262), .B1(n15261), .B2(n15270), .ZN(
        P3_U3464) );
  AOI22_X1 U16777 ( .A1(n15269), .A2(n15264), .B1(n15263), .B2(n15270), .ZN(
        P3_U3465) );
  AOI22_X1 U16778 ( .A1(n15269), .A2(n15265), .B1(n11124), .B2(n15270), .ZN(
        P3_U3466) );
  AOI22_X1 U16779 ( .A1(n15269), .A2(n15267), .B1(n15266), .B2(n15270), .ZN(
        P3_U3467) );
  AOI22_X1 U16780 ( .A1(n15269), .A2(n15268), .B1(n11137), .B2(n15270), .ZN(
        P3_U3468) );
  AOI22_X1 U16781 ( .A1(n15269), .A2(n15272), .B1(n15271), .B2(n15270), .ZN(
        P3_U3469) );
  XOR2_X1 U16782 ( .A(n15274), .B(n15273), .Z(SUB_1596_U59) );
  XOR2_X1 U16783 ( .A(n15276), .B(n15275), .Z(SUB_1596_U58) );
  AOI21_X1 U16784 ( .B1(n15278), .B2(n15277), .A(n15287), .ZN(SUB_1596_U53) );
  XOR2_X1 U16785 ( .A(n15280), .B(n15279), .Z(SUB_1596_U56) );
  OAI21_X1 U16786 ( .B1(n15283), .B2(n15282), .A(n15281), .ZN(n15285) );
  XOR2_X1 U16787 ( .A(n15285), .B(n15284), .Z(SUB_1596_U60) );
  XOR2_X1 U16788 ( .A(n15287), .B(n15286), .Z(SUB_1596_U5) );
  INV_X2 U7378 ( .A(n8049), .ZN(n7992) );
  CLKBUF_X2 U7230 ( .A(n9652), .Z(n6722) );
  INV_X1 U7266 ( .A(n12463), .ZN(n15188) );
  CLKBUF_X1 U7272 ( .A(n8678), .Z(n6473) );
  NAND2_X1 U7296 ( .A1(n10217), .A2(n13589), .ZN(n9832) );
  OAI211_X1 U7301 ( .C1(n9231), .C2(n9690), .A(n8949), .B(n8948), .ZN(n10900)
         );
  CLKBUF_X1 U7369 ( .A(n8529), .Z(n6469) );
endmodule

