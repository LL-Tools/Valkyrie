

module b20_C_SARLock_k_64_3 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10145;

  BUF_X1 U4774 ( .A(n6209), .Z(n4267) );
  AND2_X1 U4775 ( .A1(n5467), .A2(n5466), .ZN(n8573) );
  OR2_X1 U4776 ( .A1(n7508), .A2(n7853), .ZN(n7615) );
  INV_X1 U4777 ( .A(n5888), .ZN(n6500) );
  INV_X1 U4778 ( .A(n5693), .ZN(n6173) );
  INV_X1 U4779 ( .A(n5380), .ZN(n8367) );
  BUF_X1 U4780 ( .A(n7278), .Z(n4269) );
  NAND4_X1 U4781 ( .A1(n4952), .A2(n4951), .A3(n4950), .A4(n4949), .ZN(n6985)
         );
  INV_X1 U4782 ( .A(n6509), .ZN(n6161) );
  NAND2_X1 U4783 ( .A1(n5706), .A2(n5705), .ZN(n8975) );
  INV_X1 U4784 ( .A(n5718), .ZN(n5781) );
  AND2_X1 U4786 ( .A1(n8414), .A2(n4358), .ZN(n4485) );
  AOI21_X1 U4787 ( .B1(n4485), .B2(n8430), .A(n4484), .ZN(n4483) );
  NAND2_X1 U4788 ( .A1(n6984), .A2(n7931), .ZN(n5527) );
  BUF_X1 U4789 ( .A(n5726), .Z(n4274) );
  INV_X1 U4790 ( .A(n6755), .ZN(n6087) );
  OR2_X1 U4791 ( .A1(n9551), .A2(n9120), .ZN(n6591) );
  XNOR2_X1 U4792 ( .A(n7367), .B(n7220), .ZN(n7365) );
  INV_X2 U4793 ( .A(n8355), .ZN(n4275) );
  NAND2_X1 U4794 ( .A1(n5324), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5326) );
  AND2_X1 U4795 ( .A1(n5487), .A2(n5486), .ZN(n8564) );
  XNOR2_X1 U4796 ( .A(n4924), .B(P2_IR_REG_30__SCAN_IN), .ZN(n4929) );
  OAI211_X1 U4798 ( .C1(n5888), .C2(n6748), .A(n5792), .B(n5791), .ZN(n9932)
         );
  CLKBUF_X2 U4799 ( .A(n6505), .Z(n4268) );
  NAND2_X1 U4800 ( .A1(n5988), .A2(n5987), .ZN(n9817) );
  BUF_X1 U4801 ( .A(n4313), .Z(n4314) );
  AOI211_X1 U4802 ( .C1(n9933), .C2(n9521), .A(n9520), .B(n9519), .ZN(n9522)
         );
  XNOR2_X1 U4803 ( .A(n5112), .B(n5111), .ZN(n6757) );
  INV_X1 U4804 ( .A(n9671), .ZN(n9896) );
  NAND4_X2 U4805 ( .A1(n4912), .A2(n4790), .A3(n4886), .A4(n4885), .ZN(n4995)
         );
  INV_X2 U4806 ( .A(n5672), .ZN(n5674) );
  XNOR2_X2 U4807 ( .A(n5762), .B(n5745), .ZN(n6789) );
  OR2_X2 U4808 ( .A1(n5725), .A2(n5892), .ZN(n5762) );
  XNOR2_X1 U4809 ( .A(n5665), .B(n5633), .ZN(n6209) );
  OR2_X2 U4810 ( .A1(n5158), .A2(n4395), .ZN(n5523) );
  XNOR2_X2 U4811 ( .A(n8971), .B(n4270), .ZN(n7284) );
  NAND2_X4 U4812 ( .A1(n4938), .A2(n4937), .ZN(n5000) );
  NOR2_X2 U4813 ( .A1(n5271), .A2(n5270), .ZN(n5274) );
  NAND2_X1 U4814 ( .A1(n5672), .A2(n7920), .ZN(n6505) );
  NAND2_X2 U4815 ( .A1(n5917), .A2(n5916), .ZN(n7853) );
  INV_X2 U4816 ( .A(n6985), .ZN(n6984) );
  OAI22_X2 U4817 ( .A1(n7237), .A2(n7238), .B1(n6329), .B2(n7247), .ZN(n7351)
         );
  NOR2_X2 U4818 ( .A1(n7387), .A2(n4905), .ZN(n7370) );
  NOR2_X2 U4819 ( .A1(n7386), .A2(n7388), .ZN(n7387) );
  XNOR2_X1 U4820 ( .A(n7365), .B(n8459), .ZN(n7366) );
  NOR4_X2 U4821 ( .A1(n8674), .A2(n4353), .A3(n8399), .A4(n8398), .ZN(n8400)
         );
  AOI21_X2 U4822 ( .B1(n7132), .B2(n5531), .A(n4891), .ZN(n7205) );
  NAND2_X1 U4823 ( .A1(n5528), .A2(n7078), .ZN(n7132) );
  AOI21_X2 U4824 ( .B1(n9464), .B2(n9465), .A(n6679), .ZN(n9446) );
  OAI21_X2 U4825 ( .B1(n9474), .B2(n6678), .A(n6594), .ZN(n9464) );
  OAI21_X2 U4826 ( .B1(n7202), .B2(n7201), .A(n7199), .ZN(n7438) );
  NAND2_X1 U4827 ( .A1(n5028), .A2(n8233), .ZN(n7202) );
  NOR4_X2 U4828 ( .A1(n8404), .A2(n8615), .A3(n4701), .A4(n8403), .ZN(n8405)
         );
  CLKBUF_X1 U4829 ( .A(n9919), .Z(n4270) );
  AOI21_X2 U4830 ( .B1(n7124), .B2(n7125), .A(n6989), .ZN(n6997) );
  OAI22_X2 U4831 ( .A1(n7117), .A2(n7116), .B1(n6985), .B2(n6987), .ZN(n7124)
         );
  NOR4_X2 U4832 ( .A1(n8407), .A2(n8561), .A3(n8571), .A4(n8406), .ZN(n8409)
         );
  INV_X2 U4833 ( .A(n5234), .ZN(n7894) );
  OAI22_X2 U4834 ( .A1(n7743), .A2(n4705), .B1(n8099), .B2(n4704), .ZN(n5234)
         );
  OAI22_X2 U4835 ( .A1(n7515), .A2(n4531), .B1(n4314), .B2(n8973), .ZN(n9885)
         );
  XNOR2_X2 U4836 ( .A(n6449), .B(n4313), .ZN(n4531) );
  INV_X2 U4837 ( .A(n7363), .ZN(n7367) );
  NAND2_X2 U4838 ( .A1(n5636), .A2(n5635), .ZN(n9551) );
  BUF_X2 U4839 ( .A(n5718), .Z(n4272) );
  AND2_X1 U4841 ( .A1(n5672), .A2(n5675), .ZN(n5718) );
  NAND2_X4 U4842 ( .A1(n6039), .A2(n5693), .ZN(n5769) );
  AOI21_X1 U4843 ( .B1(n8865), .B2(n6715), .A(n6403), .ZN(n6718) );
  OR2_X1 U4844 ( .A1(n9188), .A2(n9159), .ZN(n4646) );
  AND2_X1 U4845 ( .A1(n8526), .A2(n8525), .ZN(n8529) );
  INV_X1 U4846 ( .A(n8711), .ZN(n8760) );
  OR2_X1 U4847 ( .A1(n6953), .A2(n5888), .ZN(n6028) );
  NAND2_X2 U4848 ( .A1(n8253), .A2(n8263), .ZN(n8391) );
  NAND2_X1 U4849 ( .A1(n5699), .A2(n6897), .ZN(n6862) );
  INV_X1 U4850 ( .A(n8245), .ZN(n8234) );
  INV_X1 U4851 ( .A(n7299), .ZN(n9925) );
  INV_X2 U4852 ( .A(n9932), .ZN(n7311) );
  INV_X2 U4853 ( .A(n6983), .ZN(n7931) );
  CLKBUF_X2 U4854 ( .A(n5693), .Z(n6394) );
  AND2_X1 U4856 ( .A1(n4684), .A2(n4929), .ZN(n5084) );
  INV_X1 U4857 ( .A(n6412), .ZN(n5682) );
  NAND2_X2 U4859 ( .A1(n6707), .A2(n6209), .ZN(n6755) );
  INV_X2 U4860 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4885) );
  OAI21_X1 U4861 ( .B1(n6701), .B2(n4291), .A(n4290), .ZN(n4289) );
  NAND2_X1 U4862 ( .A1(n8553), .A2(n7972), .ZN(n7973) );
  AOI21_X1 U4863 ( .B1(n7970), .B2(n8657), .A(n7969), .ZN(n8553) );
  OR2_X1 U4864 ( .A1(n8559), .A2(n10081), .ZN(n7972) );
  AND2_X1 U4865 ( .A1(n4690), .A2(n4324), .ZN(n8562) );
  OR2_X1 U4866 ( .A1(n6718), .A2(n6443), .ZN(n6444) );
  NOR2_X1 U4867 ( .A1(n4329), .A2(n4375), .ZN(n4557) );
  AND2_X1 U4868 ( .A1(n4831), .A2(n4832), .ZN(n9175) );
  MUX2_X1 U4869 ( .A(n6838), .B(n6633), .S(n9105), .Z(n6634) );
  NOR2_X1 U4870 ( .A1(n4300), .A2(n9137), .ZN(n9187) );
  OAI21_X1 U4871 ( .B1(n6630), .B2(n9163), .A(n6629), .ZN(n6633) );
  AND2_X1 U4872 ( .A1(n6702), .A2(n6703), .ZN(n4291) );
  AND2_X1 U4873 ( .A1(n8014), .A2(n8013), .ZN(n8074) );
  INV_X1 U4874 ( .A(n6713), .ZN(n4290) );
  NAND2_X1 U4875 ( .A1(n8602), .A2(n5387), .ZN(n8594) );
  NAND2_X1 U4876 ( .A1(n4693), .A2(n4691), .ZN(n8614) );
  NAND2_X1 U4877 ( .A1(n4276), .A2(n6608), .ZN(n6612) );
  NAND2_X1 U4878 ( .A1(n4280), .A2(n4279), .ZN(n4278) );
  NAND2_X1 U4879 ( .A1(n7936), .A2(n7937), .ZN(n7940) );
  NAND2_X1 U4880 ( .A1(n6603), .A2(n6838), .ZN(n4277) );
  NAND2_X1 U4881 ( .A1(n4281), .A2(n9150), .ZN(n4280) );
  AND2_X1 U4882 ( .A1(n6606), .A2(n4340), .ZN(n6609) );
  AND2_X1 U4883 ( .A1(n8760), .A2(n8573), .ZN(n8344) );
  OAI21_X1 U4884 ( .B1(n4655), .B2(n9151), .A(n9152), .ZN(n4654) );
  NAND2_X1 U4885 ( .A1(n4874), .A2(n4872), .ZN(n8198) );
  AND2_X1 U4886 ( .A1(n8081), .A2(n4862), .ZN(n4306) );
  NOR2_X1 U4887 ( .A1(n6604), .A2(n6838), .ZN(n4279) );
  NAND2_X1 U4888 ( .A1(n4442), .A2(n6022), .ZN(n4440) );
  NAND2_X1 U4889 ( .A1(n6366), .A2(n6365), .ZN(n9525) );
  OR2_X1 U4890 ( .A1(n8672), .A2(n5543), .ZN(n7935) );
  AND2_X1 U4891 ( .A1(n5460), .A2(n5459), .ZN(n8711) );
  NAND2_X1 U4892 ( .A1(n4719), .A2(n4718), .ZN(n6023) );
  NAND2_X1 U4893 ( .A1(n6160), .A2(n6159), .ZN(n9536) );
  AND2_X1 U4894 ( .A1(n8666), .A2(n5544), .ZN(n8665) );
  INV_X1 U4895 ( .A(n6588), .ZN(n4546) );
  NAND2_X1 U4896 ( .A1(n6126), .A2(n6125), .ZN(n9546) );
  NAND2_X1 U4897 ( .A1(n8402), .A2(n8299), .ZN(n8668) );
  NAND2_X1 U4898 ( .A1(n4907), .A2(n5540), .ZN(n7658) );
  AND2_X1 U4899 ( .A1(n5539), .A2(n8277), .ZN(n4907) );
  OAI21_X1 U4900 ( .B1(n5435), .B2(n5434), .A(n5433), .ZN(n5453) );
  NAND2_X1 U4901 ( .A1(n5371), .A2(n5370), .ZN(n5435) );
  NAND2_X1 U4902 ( .A1(n4296), .A2(n6576), .ZN(n6578) );
  NAND2_X1 U4903 ( .A1(n5311), .A2(n5310), .ZN(n8662) );
  OR2_X1 U4904 ( .A1(n7683), .A2(n7785), .ZN(n9810) );
  AND2_X1 U4905 ( .A1(n6675), .A2(n6672), .ZN(n6583) );
  OAI21_X1 U4906 ( .B1(n7856), .B2(n4792), .A(n4791), .ZN(n8465) );
  INV_X1 U4907 ( .A(n8289), .ZN(n8397) );
  NAND2_X1 U4908 ( .A1(n5329), .A2(n5328), .ZN(n8735) );
  NAND2_X1 U4909 ( .A1(n6089), .A2(n6088), .ZN(n9561) );
  NAND2_X1 U4910 ( .A1(n4587), .A2(n4585), .ZN(n7546) );
  NAND2_X1 U4911 ( .A1(n6028), .A2(n6027), .ZN(n9668) );
  OR2_X1 U4912 ( .A1(n7790), .A2(n9108), .ZN(n6669) );
  AOI21_X1 U4913 ( .B1(n4856), .B2(n4854), .A(n4371), .ZN(n4853) );
  NAND2_X1 U4914 ( .A1(n6010), .A2(n6009), .ZN(n7790) );
  AOI21_X1 U4915 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9758), .A(n9766), .ZN(
        n9047) );
  AND2_X1 U4916 ( .A1(n7165), .A2(n4723), .ZN(n4721) );
  NAND2_X1 U4917 ( .A1(n5265), .A2(n5264), .ZN(n5287) );
  NOR2_X1 U4918 ( .A1(n4857), .A2(n7595), .ZN(n4856) );
  NAND2_X1 U4919 ( .A1(n4294), .A2(n6552), .ZN(n4293) );
  AOI21_X1 U4920 ( .B1(n4882), .B2(n4904), .A(n4335), .ZN(n4875) );
  NAND2_X1 U4921 ( .A1(n5207), .A2(n5206), .ZN(n5214) );
  OR2_X1 U4922 ( .A1(n7853), .A2(n7611), .ZN(n6566) );
  NAND2_X1 U4923 ( .A1(n5201), .A2(n5178), .ZN(n6823) );
  OAI21_X1 U4924 ( .B1(n9859), .B2(n4676), .A(n4673), .ZN(n9843) );
  AND2_X1 U4925 ( .A1(n4434), .A2(n5776), .ZN(n4433) );
  NAND2_X1 U4926 ( .A1(n5201), .A2(n5200), .ZN(n5207) );
  NAND2_X1 U4927 ( .A1(n5867), .A2(n5866), .ZN(n7680) );
  NAND2_X1 U4928 ( .A1(n6547), .A2(n6550), .ZN(n7294) );
  OR2_X1 U4929 ( .A1(n5177), .A2(n5176), .ZN(n5201) );
  NAND2_X1 U4930 ( .A1(n9859), .A2(n6649), .ZN(n6547) );
  OAI22_X1 U4931 ( .A1(n5174), .A2(n5173), .B1(SI_11_), .B2(n5172), .ZN(n5177)
         );
  NAND2_X1 U4932 ( .A1(n7274), .A2(n6452), .ZN(n9859) );
  INV_X2 U4933 ( .A(n7363), .ZN(n8037) );
  AOI21_X1 U4934 ( .B1(n9874), .B2(n6451), .A(n6643), .ZN(n7275) );
  AOI21_X1 U4935 ( .B1(n6322), .B2(n6972), .A(n6955), .ZN(n7059) );
  NAND2_X1 U4936 ( .A1(n5064), .A2(n5063), .ZN(n5075) );
  AND2_X1 U4937 ( .A1(n7516), .A2(n6450), .ZN(n9874) );
  AOI21_X1 U4938 ( .B1(n6208), .B2(n9667), .A(n9847), .ZN(n8951) );
  INV_X1 U4939 ( .A(n7364), .ZN(n8457) );
  INV_X1 U4940 ( .A(n8462), .ZN(n4987) );
  BUF_X1 U4941 ( .A(n6449), .Z(n8973) );
  INV_X2 U4942 ( .A(n6039), .ZN(n6421) );
  AND2_X1 U4943 ( .A1(n4968), .A2(n4967), .ZN(n6983) );
  NAND4_X1 U4944 ( .A1(n5788), .A2(n5787), .A3(n5786), .A4(n5785), .ZN(n8969)
         );
  AOI21_X1 U4945 ( .B1(n6320), .B2(n7049), .A(n7033), .ZN(n6910) );
  AND2_X2 U4946 ( .A1(n5591), .A2(n6826), .ZN(n6977) );
  AND4_X1 U4947 ( .A1(n4933), .A2(n4932), .A3(n4931), .A4(n4930), .ZN(n7924)
         );
  NAND2_X1 U4948 ( .A1(n7494), .A2(n4427), .ZN(n6039) );
  NAND4_X1 U4949 ( .A1(n5744), .A2(n5743), .A3(n5742), .A4(n5741), .ZN(n8971)
         );
  NAND4_X1 U4950 ( .A1(n5724), .A2(n5723), .A3(n5722), .A4(n5721), .ZN(n8972)
         );
  NAND2_X1 U4951 ( .A1(n5589), .A2(n5588), .ZN(n5591) );
  CLKBUF_X3 U4952 ( .A(n5084), .Z(n5312) );
  INV_X2 U4953 ( .A(n4997), .ZN(n5509) );
  INV_X2 U4954 ( .A(n5039), .ZN(n8209) );
  OAI211_X1 U4955 ( .C1(n6755), .C2(n6790), .A(n5691), .B(n4299), .ZN(n4313)
         );
  NAND2_X1 U4956 ( .A1(n5309), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5323) );
  INV_X2 U4957 ( .A(n4274), .ZN(n6364) );
  AND2_X2 U4958 ( .A1(n8823), .A2(n4684), .ZN(n4971) );
  INV_X1 U4959 ( .A(n8827), .ZN(n4684) );
  OR2_X1 U4960 ( .A1(n5726), .A2(n6733), .ZN(n4299) );
  INV_X2 U4961 ( .A(n6316), .ZN(n8434) );
  INV_X1 U4962 ( .A(n7916), .ZN(n7795) );
  CLKBUF_X1 U4963 ( .A(n5604), .Z(n4310) );
  INV_X1 U4964 ( .A(n4929), .ZN(n8823) );
  NAND2_X1 U4965 ( .A1(n4927), .A2(n4926), .ZN(n8827) );
  AND2_X1 U4966 ( .A1(n5586), .A2(n5585), .ZN(n7916) );
  MUX2_X1 U4967 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4944), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n4947) );
  MUX2_X1 U4968 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4925), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n4927) );
  XNOR2_X1 U4969 ( .A(n5522), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8383) );
  OR2_X1 U4970 ( .A1(n5584), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U4971 ( .A1(n4926), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4924) );
  OR2_X1 U4972 ( .A1(n5668), .A2(n5892), .ZN(n5665) );
  AND2_X1 U4973 ( .A1(n4887), .A2(n4498), .ZN(n4621) );
  NAND2_X1 U4974 ( .A1(n4339), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5583) );
  AND2_X1 U4975 ( .A1(n4283), .A2(n4288), .ZN(n5668) );
  XNOR2_X1 U4976 ( .A(n5108), .B(SI_8_), .ZN(n5111) );
  OR2_X1 U4977 ( .A1(n5653), .A2(n5892), .ZN(n5634) );
  NAND2_X1 U4978 ( .A1(n5639), .A2(n5638), .ZN(n6046) );
  NAND2_X2 U4979 ( .A1(n4425), .A2(P1_U3086), .ZN(n9590) );
  BUF_X1 U4980 ( .A(n6735), .Z(n4425) );
  NOR2_X1 U4981 ( .A1(n4960), .A2(n4959), .ZN(n4962) );
  INV_X1 U4982 ( .A(n6024), .ZN(n5639) );
  AND2_X1 U4983 ( .A1(n4889), .A2(n4919), .ZN(n4887) );
  AND4_X1 U4984 ( .A1(n10145), .A2(n4286), .A3(n5630), .A4(n4285), .ZN(n4283)
         );
  NAND2_X2 U4985 ( .A1(n6736), .A2(P2_U3151), .ZN(n8822) );
  INV_X4 U4986 ( .A(n6736), .ZN(n6735) );
  INV_X1 U4987 ( .A(n4319), .ZN(n4286) );
  AND4_X1 U4988 ( .A1(n5629), .A2(n5628), .A3(n5627), .A4(n4454), .ZN(n5630)
         );
  NAND2_X1 U4990 ( .A1(n4282), .A2(n4287), .ZN(n4319) );
  INV_X1 U4991 ( .A(n4819), .ZN(n4282) );
  NOR2_X1 U4992 ( .A1(n4726), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n4288) );
  AND3_X1 U4993 ( .A1(n4915), .A2(n4914), .A3(n4913), .ZN(n4465) );
  AND2_X1 U4994 ( .A1(n5747), .A2(n5745), .ZN(n5760) );
  INV_X1 U4995 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4935) );
  INV_X4 U4996 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U4997 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5269) );
  INV_X4 U4998 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U4999 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5725) );
  NOR2_X1 U5000 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4916) );
  INV_X1 U5001 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6067) );
  INV_X1 U5002 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5146) );
  INV_X1 U5003 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4790) );
  NOR2_X1 U5004 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4804) );
  INV_X1 U5005 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4287) );
  NOR2_X1 U5006 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5632) );
  INV_X1 U5007 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5273) );
  INV_X1 U5008 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5267) );
  INV_X1 U5009 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4917) );
  NOR2_X1 U5010 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n4686) );
  INV_X1 U5011 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4285) );
  NAND3_X1 U5012 ( .A1(n4278), .A2(n4277), .A3(n6609), .ZN(n4276) );
  NAND4_X1 U5013 ( .A1(n6592), .A2(n6591), .A3(n6597), .A4(n6590), .ZN(n4281)
         );
  NAND3_X1 U5014 ( .A1(n4288), .A2(n5630), .A3(n10145), .ZN(n6200) );
  NAND3_X1 U5015 ( .A1(n6714), .A2(n6712), .A3(n4289), .ZN(P1_U3242) );
  NAND2_X1 U5016 ( .A1(n4292), .A2(n4572), .ZN(n4571) );
  NAND2_X1 U5017 ( .A1(n4293), .A2(n7318), .ZN(n4292) );
  NAND2_X1 U5018 ( .A1(n6551), .A2(n4295), .ZN(n4294) );
  AND2_X1 U5019 ( .A1(n6550), .A2(n6650), .ZN(n4295) );
  NAND2_X1 U5020 ( .A1(n7275), .A2(n7284), .ZN(n7274) );
  NAND3_X1 U5021 ( .A1(n4298), .A2(n4297), .A3(n7684), .ZN(n4296) );
  NAND3_X1 U5022 ( .A1(n6562), .A2(n6664), .A3(n6838), .ZN(n4297) );
  NAND3_X1 U5023 ( .A1(n6571), .A2(n6703), .A3(n6570), .ZN(n4298) );
  AND2_X1 U5024 ( .A1(n6669), .A2(n9660), .ZN(n6536) );
  NOR2_X2 U5025 ( .A1(n9490), .A2(n6470), .ZN(n9474) );
  AND2_X1 U5026 ( .A1(n4835), .A2(n4828), .ZN(n4300) );
  CLKBUF_X1 U5027 ( .A(n9851), .Z(n4301) );
  NAND4_X1 U5028 ( .A1(n5760), .A2(n4804), .A3(n5622), .A4(n5725), .ZN(n4302)
         );
  OR2_X1 U5030 ( .A1(n5243), .A2(n5242), .ZN(n5244) );
  OAI21_X1 U5031 ( .B1(n5287), .B2(n4776), .A(n4774), .ZN(n5337) );
  OAI21_X1 U5032 ( .B1(n5559), .B2(n4483), .A(n4479), .ZN(n4478) );
  OR2_X2 U5033 ( .A1(n5378), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5396) );
  OR2_X2 U5034 ( .A1(n5228), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5251) );
  OR2_X2 U5035 ( .A1(n5461), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U5036 ( .A1(n4809), .A2(n4812), .ZN(n7505) );
  NAND2_X1 U5037 ( .A1(n7479), .A2(n7478), .ZN(n9824) );
  NAND2_X2 U5038 ( .A1(n9232), .A2(n9131), .ZN(n9219) );
  NAND2_X1 U5039 ( .A1(n8080), .A2(n4306), .ZN(n4303) );
  AND2_X2 U5040 ( .A1(n4303), .A2(n4304), .ZN(n4860) );
  OR2_X1 U5041 ( .A1(n4305), .A2(n8002), .ZN(n4304) );
  INV_X1 U5042 ( .A(n4862), .ZN(n4305) );
  INV_X1 U5043 ( .A(n4859), .ZN(n4307) );
  NAND2_X1 U5044 ( .A1(n4308), .A2(n4860), .ZN(n8016) );
  NOR2_X1 U5045 ( .A1(n8009), .A2(n4307), .ZN(n4308) );
  CLKBUF_X1 U5046 ( .A(n7904), .Z(n4309) );
  XNOR2_X1 U5047 ( .A(n7901), .B(n7581), .ZN(n7904) );
  NAND2_X2 U5048 ( .A1(n7536), .A2(n7535), .ZN(n7597) );
  XNOR2_X1 U5049 ( .A(n5579), .B(n5578), .ZN(n5604) );
  NAND2_X1 U5050 ( .A1(n6755), .A2(n6735), .ZN(n4311) );
  NAND2_X1 U5051 ( .A1(n6755), .A2(n6735), .ZN(n4312) );
  NAND2_X1 U5052 ( .A1(n6755), .A2(n6735), .ZN(n5888) );
  OR2_X2 U5053 ( .A1(n5523), .A2(n4495), .ZN(n4339) );
  AND2_X1 U5054 ( .A1(n4464), .A2(n4465), .ZN(n4852) );
  AOI21_X2 U5055 ( .B1(n9472), .B2(n9475), .A(n4902), .ZN(n9458) );
  OAI21_X2 U5056 ( .B1(n9502), .B2(n9112), .A(n9493), .ZN(n9472) );
  NAND2_X2 U5057 ( .A1(n5587), .A2(n7916), .ZN(n5592) );
  NAND2_X2 U5058 ( .A1(n8198), .A2(n7991), .ZN(n8111) );
  OAI21_X2 U5059 ( .B1(n7366), .B2(n4876), .A(n4875), .ZN(n7386) );
  NAND2_X1 U5060 ( .A1(n4878), .A2(n7065), .ZN(n4876) );
  AOI21_X2 U5061 ( .B1(n7904), .B2(n7903), .A(n7902), .ZN(n7905) );
  NAND2_X2 U5062 ( .A1(n8433), .A2(n8412), .ZN(n6973) );
  NOR2_X2 U5063 ( .A1(n4995), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5037) );
  NOR2_X1 U5064 ( .A1(n5111), .A2(n4757), .ZN(n4756) );
  INV_X1 U5065 ( .A(n5080), .ZN(n4757) );
  OR2_X1 U5066 ( .A1(n8624), .A2(n8632), .ZN(n8332) );
  OR2_X1 U5067 ( .A1(n8748), .A2(n8678), .ZN(n8295) );
  INV_X1 U5068 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4919) );
  NAND2_X1 U5069 ( .A1(n8432), .A2(n4897), .ZN(n4484) );
  AND2_X1 U5070 ( .A1(n4916), .A2(n5146), .ZN(n4464) );
  XNOR2_X1 U5071 ( .A(n6269), .B(n7087), .ZN(n10019) );
  AOI21_X1 U5072 ( .B1(n4552), .B2(n4555), .A(n4551), .ZN(n4550) );
  INV_X1 U5073 ( .A(n4553), .ZN(n4552) );
  OAI21_X1 U5074 ( .B1(n4555), .B2(n6611), .A(n4554), .ZN(n4553) );
  AOI21_X1 U5075 ( .B1(n6976), .B2(n6975), .A(n6974), .ZN(n6978) );
  NAND2_X1 U5076 ( .A1(n8347), .A2(n8374), .ZN(n4509) );
  OR2_X1 U5077 ( .A1(n6277), .A2(n6922), .ZN(n6278) );
  AOI21_X1 U5078 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n6824), .A(n7886), .ZN(
        n6293) );
  NOR2_X1 U5079 ( .A1(n8556), .A2(n8564), .ZN(n8349) );
  AND2_X1 U5080 ( .A1(n5532), .A2(n8382), .ZN(n8240) );
  INV_X1 U5081 ( .A(n8349), .ZN(n4613) );
  OR2_X1 U5082 ( .A1(n8774), .A2(n8446), .ZN(n5426) );
  OR2_X1 U5083 ( .A1(n8774), .A2(n8596), .ZN(n8337) );
  OR2_X1 U5084 ( .A1(n8731), .A2(n8645), .ZN(n8320) );
  AND2_X1 U5085 ( .A1(n8208), .A2(n8678), .ZN(n5257) );
  INV_X1 U5086 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5608) );
  INV_X1 U5087 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4749) );
  INV_X1 U5088 ( .A(n4428), .ZN(n4427) );
  OAI21_X1 U5089 ( .B1(n6834), .B2(n6704), .A(n6731), .ZN(n4428) );
  INV_X1 U5090 ( .A(n4894), .ZN(n4716) );
  INV_X1 U5091 ( .A(n5738), .ZN(n4435) );
  AND2_X1 U5092 ( .A1(n4651), .A2(n9260), .ZN(n4649) );
  NAND2_X1 U5093 ( .A1(n4652), .A2(n4654), .ZN(n4651) );
  NOR2_X1 U5094 ( .A1(n7612), .A2(n4848), .ZN(n4847) );
  OR2_X1 U5095 ( .A1(n9510), .A2(n6510), .ZN(n6627) );
  NOR2_X1 U5096 ( .A1(n9510), .A2(n9515), .ZN(n4566) );
  INV_X1 U5097 ( .A(n7533), .ZN(n6644) );
  NAND2_X1 U5098 ( .A1(n5508), .A2(n5507), .ZN(n6493) );
  AND2_X1 U5099 ( .A1(n5491), .A2(n5476), .ZN(n5489) );
  OR2_X1 U5100 ( .A1(n6200), .A2(n4819), .ZN(n5651) );
  NAND2_X1 U5101 ( .A1(n4349), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5658) );
  OR2_X1 U5102 ( .A1(n5337), .A2(n5338), .ZN(n5342) );
  NAND2_X1 U5103 ( .A1(n5183), .A2(n5182), .ZN(n5194) );
  NOR2_X1 U5104 ( .A1(n6258), .A2(n7348), .ZN(n6259) );
  OR2_X1 U5105 ( .A1(n8465), .A2(n4411), .ZN(n4630) );
  NAND2_X1 U5106 ( .A1(n8465), .A2(n4632), .ZN(n4629) );
  AOI21_X1 U5107 ( .B1(n4701), .B2(n4345), .A(n4700), .ZN(n4699) );
  NOR2_X1 U5108 ( .A1(n5336), .A2(n8631), .ZN(n4700) );
  AND3_X1 U5109 ( .A1(n5364), .A2(n5363), .A3(n5362), .ZN(n8632) );
  NAND2_X1 U5110 ( .A1(n7992), .A2(n5298), .ZN(n5299) );
  OR2_X1 U5111 ( .A1(n7664), .A2(n8156), .ZN(n8281) );
  INV_X1 U5112 ( .A(n5132), .ZN(n4683) );
  XNOR2_X1 U5113 ( .A(n8358), .B(n8443), .ZN(n8408) );
  OR2_X1 U5114 ( .A1(n8735), .A2(n8631), .ZN(n8311) );
  INV_X1 U5115 ( .A(n8662), .ZN(n8742) );
  INV_X1 U5116 ( .A(n6242), .ZN(n5327) );
  NAND2_X1 U5117 ( .A1(n4590), .A2(n4594), .ZN(n5542) );
  INV_X1 U5118 ( .A(n4595), .ZN(n4594) );
  AND2_X1 U5119 ( .A1(n5520), .A2(n4344), .ZN(n8439) );
  INV_X1 U5120 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4912) );
  INV_X1 U5121 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4886) );
  NOR2_X1 U5122 ( .A1(n4462), .A2(n4365), .ZN(n4460) );
  AOI21_X1 U5123 ( .B1(n4341), .B2(n9159), .A(n4648), .ZN(n4647) );
  INV_X1 U5124 ( .A(n9160), .ZN(n4648) );
  NAND2_X1 U5125 ( .A1(n4821), .A2(n4824), .ZN(n9174) );
  AND2_X1 U5126 ( .A1(n4388), .A2(n4825), .ZN(n4824) );
  NAND2_X1 U5127 ( .A1(n4829), .A2(n4826), .ZN(n4825) );
  NAND2_X1 U5128 ( .A1(n4835), .A2(n4828), .ZN(n4833) );
  NAND2_X1 U5129 ( .A1(n5201), .A2(n4525), .ZN(n4527) );
  NOR2_X1 U5130 ( .A1(n5206), .A2(n4526), .ZN(n4525) );
  INV_X1 U5131 ( .A(n5200), .ZN(n4526) );
  INV_X1 U5132 ( .A(n9828), .ZN(n9876) );
  OR2_X1 U5133 ( .A1(n9171), .A2(n9828), .ZN(n4662) );
  AND2_X1 U5134 ( .A1(n4647), .A2(n4644), .ZN(n4643) );
  INV_X1 U5135 ( .A(n9181), .ZN(n4644) );
  NAND2_X1 U5136 ( .A1(n6627), .A2(n6628), .ZN(n9163) );
  NAND2_X1 U5137 ( .A1(n4450), .A2(n4449), .ZN(n5641) );
  AOI21_X1 U5138 ( .B1(n4452), .B2(n5892), .A(n5892), .ZN(n4449) );
  AND2_X1 U5139 ( .A1(n4751), .A2(n5074), .ZN(n4528) );
  NOR2_X1 U5140 ( .A1(n4755), .A2(n4752), .ZN(n4751) );
  OR3_X1 U5141 ( .A1(n7795), .A2(n5590), .A3(n5604), .ZN(n6999) );
  NAND2_X1 U5142 ( .A1(n4483), .A2(n4480), .ZN(n4479) );
  OR2_X1 U5143 ( .A1(n4485), .A2(n5559), .ZN(n4480) );
  OAI21_X1 U5144 ( .B1(n10019), .B2(n4639), .A(n4638), .ZN(n8523) );
  NAND2_X1 U5145 ( .A1(n4640), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4639) );
  OAI21_X1 U5146 ( .B1(n5572), .B2(n10037), .A(n5571), .ZN(n8544) );
  AOI21_X1 U5147 ( .B1(n5573), .B2(n7637), .A(n5570), .ZN(n5571) );
  INV_X1 U5148 ( .A(n5569), .ZN(n5570) );
  NAND2_X1 U5149 ( .A1(n8235), .A2(n8243), .ZN(n4491) );
  AND2_X1 U5150 ( .A1(n6553), .A2(n6838), .ZN(n4572) );
  INV_X1 U5151 ( .A(n8283), .ZN(n4470) );
  INV_X1 U5152 ( .A(n8293), .ZN(n4468) );
  NAND2_X1 U5153 ( .A1(n4489), .A2(n8355), .ZN(n4488) );
  INV_X1 U5154 ( .A(n8297), .ZN(n4489) );
  NOR2_X1 U5155 ( .A1(n6642), .A2(n4542), .ZN(n4541) );
  AND2_X1 U5156 ( .A1(n4391), .A2(n4533), .ZN(n4537) );
  NAND2_X1 U5157 ( .A1(n6605), .A2(n9270), .ZN(n6606) );
  AND2_X1 U5158 ( .A1(n7512), .A2(n6462), .ZN(n6563) );
  NAND2_X1 U5159 ( .A1(n4784), .A2(n4783), .ZN(n8417) );
  AND2_X1 U5160 ( .A1(n8442), .A2(n8211), .ZN(n4783) );
  OR2_X1 U5161 ( .A1(n5545), .A2(n8665), .ZN(n5547) );
  NAND2_X1 U5162 ( .A1(n4888), .A2(n4498), .ZN(n4497) );
  AND2_X1 U5163 ( .A1(n4919), .A2(n4920), .ZN(n4888) );
  INV_X1 U5164 ( .A(n8877), .ZN(n4712) );
  AOI21_X1 U5165 ( .B1(n4549), .B2(n6617), .A(n6616), .ZN(n4548) );
  INV_X1 U5166 ( .A(n4550), .ZN(n4549) );
  INV_X1 U5167 ( .A(n6563), .ZN(n6560) );
  INV_X1 U5168 ( .A(n5471), .ZN(n4764) );
  INV_X1 U5169 ( .A(n4763), .ZN(n4762) );
  OAI21_X1 U5170 ( .B1(n5469), .B2(n4764), .A(n5489), .ZN(n4763) );
  NAND2_X1 U5171 ( .A1(n5632), .A2(n4820), .ZN(n4819) );
  AND2_X1 U5172 ( .A1(n5430), .A2(n5429), .ZN(n5431) );
  NAND2_X1 U5173 ( .A1(n8357), .A2(n8362), .ZN(n4510) );
  NAND2_X1 U5174 ( .A1(n4355), .A2(n4322), .ZN(n4504) );
  NOR2_X1 U5175 ( .A1(n8356), .A2(n8350), .ZN(n4511) );
  OR2_X1 U5176 ( .A1(n5380), .A2(n4928), .ZN(n4931) );
  INV_X1 U5177 ( .A(n6964), .ZN(n4628) );
  NOR2_X1 U5178 ( .A1(n6966), .A2(n4356), .ZN(n6253) );
  AND2_X1 U5179 ( .A1(n8514), .A2(n6268), .ZN(n6269) );
  OR2_X1 U5180 ( .A1(n5618), .A2(n8046), .ZN(n8420) );
  NOR2_X1 U5181 ( .A1(n4703), .A2(n8641), .ZN(n4702) );
  INV_X1 U5182 ( .A(n5319), .ZN(n4703) );
  OR2_X1 U5183 ( .A1(n7900), .A2(n7661), .ZN(n8275) );
  OR2_X1 U5184 ( .A1(n10065), .A2(n7831), .ZN(n8260) );
  AND2_X1 U5185 ( .A1(n5606), .A2(n5605), .ZN(n6924) );
  AND2_X1 U5186 ( .A1(n8346), .A2(n8345), .ZN(n8374) );
  OR2_X1 U5187 ( .A1(n8786), .A2(n8620), .ZN(n8327) );
  AND2_X1 U5188 ( .A1(n8721), .A2(n8607), .ZN(n8377) );
  AOI21_X1 U5189 ( .B1(n4696), .B2(n4695), .A(n8616), .ZN(n4694) );
  INV_X1 U5190 ( .A(n4702), .ZN(n4695) );
  INV_X1 U5191 ( .A(n8311), .ZN(n4604) );
  OR2_X1 U5192 ( .A1(n8807), .A2(n8694), .ZN(n8305) );
  NOR2_X1 U5193 ( .A1(n8287), .A2(n4598), .ZN(n4597) );
  INV_X1 U5194 ( .A(n8281), .ZN(n4598) );
  XNOR2_X1 U5195 ( .A(n5970), .B(n6394), .ZN(n5972) );
  NOR2_X1 U5196 ( .A1(n8857), .A2(n4364), .ZN(n6137) );
  INV_X1 U5197 ( .A(n6357), .ZN(n4518) );
  NAND2_X1 U5198 ( .A1(n5682), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5687) );
  AND2_X1 U5199 ( .A1(n4834), .A2(n9138), .ZN(n4828) );
  NOR2_X1 U5200 ( .A1(n9668), .A2(n7790), .ZN(n4581) );
  NAND2_X1 U5201 ( .A1(n9977), .A2(n7784), .ZN(n4849) );
  INV_X1 U5202 ( .A(n4849), .ZN(n4841) );
  NAND2_X1 U5203 ( .A1(n7612), .A2(n6566), .ZN(n4672) );
  INV_X1 U5204 ( .A(n6566), .ZN(n4671) );
  OAI21_X1 U5205 ( .B1(n7501), .B2(n7506), .A(n6560), .ZN(n7486) );
  NOR2_X1 U5206 ( .A1(n4814), .A2(n4811), .ZN(n4810) );
  INV_X1 U5207 ( .A(n7567), .ZN(n4814) );
  INV_X1 U5208 ( .A(n9830), .ZN(n4811) );
  INV_X1 U5209 ( .A(n7481), .ZN(n4813) );
  INV_X1 U5210 ( .A(n6550), .ZN(n4678) );
  INV_X1 U5211 ( .A(n6653), .ZN(n4674) );
  INV_X1 U5212 ( .A(n4664), .ZN(n4663) );
  NAND2_X1 U5213 ( .A1(n5455), .A2(n5454), .ZN(n5470) );
  INV_X1 U5214 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5638) );
  INV_X1 U5215 ( .A(n4775), .ZN(n4774) );
  OAI21_X1 U5216 ( .B1(n4781), .B2(n4776), .A(n5320), .ZN(n4775) );
  INV_X1 U5217 ( .A(n4777), .ZN(n4776) );
  NOR2_X1 U5218 ( .A1(n5301), .A2(n4782), .ZN(n4781) );
  INV_X1 U5219 ( .A(n5286), .ZN(n4782) );
  AND2_X1 U5220 ( .A1(n5213), .A2(n5205), .ZN(n5206) );
  INV_X1 U5221 ( .A(n5136), .ZN(n4752) );
  XNOR2_X1 U5222 ( .A(n5134), .B(SI_9_), .ZN(n5136) );
  INV_X1 U5223 ( .A(n4756), .ZN(n4755) );
  AOI21_X1 U5224 ( .B1(n4754), .B2(n4756), .A(n4382), .ZN(n4753) );
  OAI21_X1 U5225 ( .B1(n6735), .B2(n4424), .A(n4423), .ZN(n5076) );
  NAND2_X1 U5226 ( .A1(n6735), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n4423) );
  NAND2_X1 U5227 ( .A1(n5001), .A2(SI_3_), .ZN(n5018) );
  OAI21_X1 U5228 ( .B1(n5000), .B2(n4523), .A(n4522), .ZN(n4521) );
  NAND3_X1 U5229 ( .A1(n4339), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_27__SCAN_IN), .ZN(n4943) );
  INV_X1 U5230 ( .A(n4903), .ZN(n4868) );
  INV_X1 U5231 ( .A(n8172), .ZN(n4867) );
  INV_X1 U5232 ( .A(n8456), .ZN(n7831) );
  AND2_X1 U5233 ( .A1(n8088), .A2(n4863), .ZN(n4862) );
  OR2_X1 U5234 ( .A1(n8144), .A2(n4864), .ZN(n4863) );
  INV_X1 U5235 ( .A(n8006), .ZN(n4864) );
  OR2_X1 U5236 ( .A1(n5165), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U5237 ( .A1(n4871), .A2(n4903), .ZN(n4870) );
  INV_X1 U5238 ( .A(n8111), .ZN(n4871) );
  AND2_X1 U5239 ( .A1(n8023), .A2(n8584), .ZN(n8183) );
  NAND2_X1 U5240 ( .A1(n8065), .A2(n8066), .ZN(n4874) );
  OAI21_X1 U5241 ( .B1(n6952), .B2(n4637), .A(n6245), .ZN(n6941) );
  AOI21_X1 U5242 ( .B1(n6959), .B2(n4741), .A(n4414), .ZN(n4740) );
  INV_X1 U5243 ( .A(n4797), .ZN(n4796) );
  NAND2_X1 U5244 ( .A1(n4748), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4745) );
  NAND2_X1 U5245 ( .A1(n6294), .A2(n4748), .ZN(n4744) );
  INV_X1 U5246 ( .A(n8475), .ZN(n4748) );
  OR2_X1 U5247 ( .A1(n7865), .A2(n7864), .ZN(n4747) );
  INV_X1 U5248 ( .A(n5562), .ZN(n6316) );
  NAND2_X1 U5249 ( .A1(n4633), .A2(n4342), .ZN(n4786) );
  NOR2_X1 U5250 ( .A1(n8344), .A2(n4615), .ZN(n4614) );
  INV_X1 U5251 ( .A(n8342), .ZN(n4615) );
  OAI22_X1 U5252 ( .A1(n8581), .A2(n4331), .B1(n4687), .B2(n4376), .ZN(n7966)
         );
  NAND2_X1 U5253 ( .A1(n4688), .A2(n4373), .ZN(n4687) );
  OR2_X1 U5254 ( .A1(n8349), .A2(n4368), .ZN(n8407) );
  NAND2_X1 U5255 ( .A1(n8443), .A2(n8653), .ZN(n7968) );
  OR2_X1 U5256 ( .A1(n5396), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U5257 ( .A1(n8652), .A2(n4702), .ZN(n4698) );
  OR2_X1 U5258 ( .A1(n5131), .A2(n5130), .ZN(n5132) );
  INV_X1 U5259 ( .A(n4586), .ZN(n4585) );
  NAND2_X1 U5260 ( .A1(n7458), .A2(n5536), .ZN(n4587) );
  OR2_X1 U5261 ( .A1(n5051), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5092) );
  OR2_X1 U5262 ( .A1(n8786), .A2(n8447), .ZN(n5387) );
  AOI21_X1 U5263 ( .B1(n4610), .B2(n4613), .A(n4368), .ZN(n4609) );
  NOR2_X1 U5264 ( .A1(n4614), .A2(n4611), .ZN(n4610) );
  NAND2_X1 U5265 ( .A1(n4607), .A2(n4606), .ZN(n4605) );
  NOR2_X1 U5266 ( .A1(n4612), .A2(n5555), .ZN(n4606) );
  NAND2_X1 U5267 ( .A1(n4613), .A2(n8345), .ZN(n4612) );
  AND2_X1 U5268 ( .A1(n5478), .A2(n5477), .ZN(n8026) );
  INV_X1 U5269 ( .A(n8374), .ZN(n8561) );
  NAND2_X1 U5270 ( .A1(n4607), .A2(n8341), .ZN(n4616) );
  AND2_X1 U5271 ( .A1(n8337), .A2(n5553), .ZN(n8582) );
  AND2_X1 U5272 ( .A1(n7080), .A2(n4275), .ZN(n8655) );
  INV_X1 U5273 ( .A(n10037), .ZN(n8657) );
  OAI21_X1 U5274 ( .B1(n8613), .B2(n5551), .A(n8332), .ZN(n8601) );
  NAND2_X1 U5275 ( .A1(n5549), .A2(n5548), .ZN(n8640) );
  NAND2_X1 U5276 ( .A1(n8640), .A2(n8641), .ZN(n8639) );
  NAND2_X1 U5277 ( .A1(n8680), .A2(n5285), .ZN(n7936) );
  INV_X1 U5278 ( .A(n8653), .ZN(n8695) );
  INV_X1 U5279 ( .A(n8291), .ZN(n4596) );
  INV_X1 U5280 ( .A(n8399), .ZN(n8690) );
  INV_X1 U5281 ( .A(n7839), .ZN(n10068) );
  AND2_X1 U5282 ( .A1(n5610), .A2(n8426), .ZN(n10037) );
  NAND2_X1 U5283 ( .A1(n4887), .A2(n4623), .ZN(n4617) );
  INV_X1 U5284 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5578) );
  INV_X1 U5285 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5575) );
  AND2_X1 U5286 ( .A1(n5912), .A2(n5911), .ZN(n7756) );
  NAND2_X1 U5287 ( .A1(n8916), .A2(n6086), .ZN(n4461) );
  NOR2_X1 U5288 ( .A1(n4330), .A2(n4362), .ZN(n4457) );
  INV_X1 U5289 ( .A(n6086), .ZN(n4458) );
  NAND2_X1 U5290 ( .A1(n6138), .A2(n4447), .ZN(n4446) );
  XNOR2_X1 U5291 ( .A(n5972), .B(n5973), .ZN(n7735) );
  XNOR2_X1 U5292 ( .A(n5731), .B(n6173), .ZN(n5735) );
  OR2_X1 U5293 ( .A1(n4518), .A2(n6183), .ZN(n4515) );
  INV_X1 U5294 ( .A(n4517), .ZN(n4516) );
  OAI21_X1 U5295 ( .B1(n6182), .B2(n4518), .A(n8866), .ZN(n4517) );
  NAND2_X1 U5296 ( .A1(n4444), .A2(n7471), .ZN(n6694) );
  NAND3_X1 U5297 ( .A1(n6188), .A2(n6184), .A3(n6185), .ZN(n6731) );
  NAND2_X1 U5298 ( .A1(n6522), .A2(n6521), .ZN(n9099) );
  OR2_X1 U5299 ( .A1(n9591), .A2(n5888), .ZN(n6522) );
  NAND2_X1 U5300 ( .A1(n9200), .A2(n9139), .ZN(n4832) );
  INV_X1 U5301 ( .A(n9158), .ZN(n9191) );
  OR2_X1 U5302 ( .A1(n9536), .A2(n9130), .ZN(n9131) );
  INV_X1 U5303 ( .A(n9283), .ZN(n4655) );
  CLKBUF_X1 U5304 ( .A(n9245), .Z(n9259) );
  OR2_X1 U5305 ( .A1(n9546), .A2(n9125), .ZN(n9126) );
  OR2_X1 U5306 ( .A1(n9278), .A2(n9124), .ZN(n4900) );
  NOR2_X1 U5307 ( .A1(n9284), .A2(n9283), .ZN(n9282) );
  OAI22_X2 U5308 ( .A1(n9806), .A2(n9808), .B1(n9817), .B2(n8960), .ZN(n9110)
         );
  AND2_X1 U5309 ( .A1(n6666), .A2(n9809), .ZN(n7684) );
  NOR2_X1 U5310 ( .A1(n4847), .A2(n4851), .ZN(n4838) );
  NAND2_X1 U5311 ( .A1(n6570), .A2(n6664), .ZN(n4837) );
  INV_X1 U5312 ( .A(n4837), .ZN(n7689) );
  OR2_X1 U5313 ( .A1(n7486), .A2(n7612), .ZN(n7488) );
  OAI22_X1 U5314 ( .A1(n9168), .A2(n9167), .B1(n9166), .B2(n9165), .ZN(n9169)
         );
  INV_X1 U5315 ( .A(n9105), .ZN(n9508) );
  NAND2_X1 U5316 ( .A1(n4568), .A2(n4567), .ZN(n9511) );
  NAND2_X1 U5317 ( .A1(n4564), .A2(n4563), .ZN(n4568) );
  OR2_X1 U5318 ( .A1(n9510), .A2(n9481), .ZN(n4563) );
  INV_X1 U5319 ( .A(n9481), .ZN(n9888) );
  NAND2_X1 U5320 ( .A1(n6072), .A2(n6071), .ZN(n9566) );
  OR2_X1 U5321 ( .A1(n7093), .A2(n5888), .ZN(n6072) );
  NAND2_X1 U5322 ( .A1(n6495), .A2(n6494), .ZN(n6516) );
  OR2_X1 U5323 ( .A1(n6493), .A2(n6492), .ZN(n6494) );
  OR2_X1 U5324 ( .A1(n6491), .A2(n6490), .ZN(n6495) );
  XNOR2_X1 U5325 ( .A(n6516), .B(n6515), .ZN(n8210) );
  NOR2_X1 U5326 ( .A1(n6200), .A2(n4319), .ZN(n5653) );
  XNOR2_X1 U5327 ( .A(n5415), .B(n5414), .ZN(n7722) );
  NAND2_X1 U5328 ( .A1(n5410), .A2(n5430), .ZN(n5415) );
  OR2_X1 U5329 ( .A1(n5435), .A2(n5428), .ZN(n5410) );
  XNOR2_X1 U5330 ( .A(n5393), .B(n5392), .ZN(n7699) );
  OAI21_X1 U5331 ( .B1(n5435), .B2(n5405), .A(n5407), .ZN(n5393) );
  NAND2_X1 U5332 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), 
        .ZN(n4729) );
  NOR2_X1 U5333 ( .A1(n5304), .A2(n4780), .ZN(n4777) );
  NAND2_X1 U5334 ( .A1(n4451), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U5335 ( .A1(n5639), .A2(n4323), .ZN(n4451) );
  INV_X1 U5336 ( .A(n4453), .ZN(n4452) );
  OAI21_X1 U5337 ( .B1(n4323), .B2(n5892), .A(n6067), .ZN(n4453) );
  NAND2_X1 U5338 ( .A1(n5259), .A2(n5258), .ZN(n5265) );
  NAND2_X1 U5339 ( .A1(n5243), .A2(n5242), .ZN(n5259) );
  NAND2_X1 U5340 ( .A1(n5985), .A2(n5637), .ZN(n6024) );
  AND2_X1 U5341 ( .A1(n5236), .A2(n5218), .ZN(n5219) );
  NAND3_X1 U5342 ( .A1(n4529), .A2(n5142), .A3(n4530), .ZN(n5157) );
  AND4_X1 U5343 ( .A1(n5318), .A2(n5317), .A3(n5316), .A4(n5315), .ZN(n8644)
         );
  AND3_X1 U5344 ( .A1(n5349), .A2(n5348), .A3(n5347), .ZN(n8645) );
  AND4_X1 U5345 ( .A1(n5199), .A2(n5198), .A3(n5197), .A4(n5196), .ZN(n8099)
         );
  AND4_X1 U5346 ( .A1(n5256), .A2(n5255), .A3(n5254), .A4(n5253), .ZN(n8678)
         );
  INV_X1 U5347 ( .A(n8607), .ZN(n8585) );
  AND2_X1 U5348 ( .A1(n5335), .A2(n5334), .ZN(n8631) );
  AND4_X1 U5349 ( .A1(n5189), .A2(n5188), .A3(n5187), .A4(n5186), .ZN(n8156)
         );
  NOR2_X1 U5350 ( .A1(n4374), .A2(n4422), .ZN(n4421) );
  INV_X1 U5351 ( .A(n8415), .ZN(n4422) );
  INV_X1 U5352 ( .A(n8440), .ZN(n4475) );
  NAND2_X1 U5353 ( .A1(n4483), .A2(n8433), .ZN(n4482) );
  INV_X1 U5354 ( .A(n8573), .ZN(n8445) );
  OR2_X1 U5355 ( .A1(n5380), .A2(n4948), .ZN(n4952) );
  NAND2_X1 U5356 ( .A1(n4798), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4797) );
  INV_X1 U5357 ( .A(n6259), .ZN(n4799) );
  NAND2_X1 U5358 ( .A1(n6259), .A2(n4636), .ZN(n4635) );
  INV_X1 U5359 ( .A(n7705), .ZN(n4636) );
  OR2_X1 U5360 ( .A1(P2_U3150), .A2(n6350), .ZN(n10010) );
  NOR2_X1 U5361 ( .A1(n8523), .A2(n6272), .ZN(n6273) );
  AND2_X1 U5362 ( .A1(P2_U3893), .A2(n5561), .ZN(n10031) );
  OR2_X1 U5363 ( .A1(n7093), .A2(n5039), .ZN(n5311) );
  NAND2_X1 U5364 ( .A1(n5212), .A2(n5211), .ZN(n9646) );
  INV_X1 U5365 ( .A(n8780), .ZN(n8721) );
  INV_X1 U5366 ( .A(n5618), .ZN(n8546) );
  NOR2_X1 U5367 ( .A1(n8544), .A2(n5574), .ZN(n6240) );
  NAND2_X1 U5368 ( .A1(n5494), .A2(n5493), .ZN(n8358) );
  INV_X1 U5369 ( .A(n8026), .ZN(n8556) );
  OR2_X1 U5370 ( .A1(n10087), .A2(n10079), .ZN(n8791) );
  INV_X1 U5371 ( .A(n8791), .ZN(n8806) );
  AND2_X1 U5372 ( .A1(n4887), .A2(n4619), .ZN(n4618) );
  AND2_X1 U5373 ( .A1(n4623), .A2(n4620), .ZN(n4619) );
  INV_X1 U5374 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4620) );
  AND2_X1 U5375 ( .A1(n4465), .A2(n4916), .ZN(n4466) );
  NAND2_X1 U5376 ( .A1(n6358), .A2(n4402), .ZN(n4429) );
  INV_X1 U5377 ( .A(n8921), .ZN(n8944) );
  INV_X1 U5378 ( .A(n8951), .ZN(n8934) );
  OR2_X1 U5379 ( .A1(n5781), .A2(n7340), .ZN(n5705) );
  AND2_X1 U5380 ( .A1(n5897), .A2(n5896), .ZN(n9602) );
  AND2_X1 U5381 ( .A1(n4662), .A2(n4582), .ZN(n4420) );
  INV_X1 U5382 ( .A(n4899), .ZN(n4582) );
  OR2_X1 U5383 ( .A1(n4643), .A2(n9162), .ZN(n4642) );
  OAI21_X1 U5384 ( .B1(n4659), .B2(n9990), .A(n4660), .ZN(n4657) );
  OR2_X1 U5385 ( .A1(n9991), .A2(n6426), .ZN(n4660) );
  AND2_X1 U5386 ( .A1(n6840), .A2(n6839), .ZN(n9828) );
  OR2_X1 U5388 ( .A1(n8384), .A2(n4357), .ZN(n4493) );
  NAND2_X1 U5389 ( .A1(n4569), .A2(n6559), .ZN(n6564) );
  NAND2_X1 U5390 ( .A1(n4469), .A2(n4467), .ZN(n8294) );
  NOR2_X1 U5391 ( .A1(n4360), .A2(n4468), .ZN(n4467) );
  NAND2_X1 U5392 ( .A1(n4486), .A2(n8300), .ZN(n8308) );
  NAND2_X1 U5393 ( .A1(n4490), .A2(n4487), .ZN(n4486) );
  AND2_X1 U5394 ( .A1(n8298), .A2(n4488), .ZN(n4487) );
  AND2_X1 U5395 ( .A1(n4546), .A2(n6577), .ZN(n4544) );
  NAND2_X1 U5396 ( .A1(n4546), .A2(n6585), .ZN(n4543) );
  NAND2_X1 U5397 ( .A1(n4546), .A2(n4534), .ZN(n4533) );
  NOR2_X1 U5398 ( .A1(n4538), .A2(n6589), .ZN(n4534) );
  INV_X1 U5399 ( .A(n4541), .ZN(n4538) );
  NOR2_X1 U5400 ( .A1(n6642), .A2(n4400), .ZN(n4540) );
  NAND2_X1 U5401 ( .A1(n9148), .A2(n6598), .ZN(n4545) );
  NAND2_X1 U5402 ( .A1(n6578), .A2(n4536), .ZN(n4535) );
  AND2_X1 U5403 ( .A1(n4546), .A2(n4392), .ZN(n4536) );
  INV_X1 U5404 ( .A(n6614), .ZN(n4555) );
  NAND2_X1 U5405 ( .A1(n6472), .A2(n9152), .ZN(n6604) );
  OR2_X1 U5406 ( .A1(n9539), .A2(n9128), .ZN(n6472) );
  NAND2_X1 U5407 ( .A1(n8462), .A2(n6979), .ZN(n8226) );
  INV_X1 U5408 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4934) );
  NOR2_X1 U5409 ( .A1(n9551), .A2(n9556), .ZN(n4575) );
  AND2_X1 U5410 ( .A1(n5367), .A2(n5354), .ZN(n4772) );
  INV_X1 U5411 ( .A(n7596), .ZN(n4854) );
  NOR2_X1 U5412 ( .A1(n6253), .A2(n7063), .ZN(n6254) );
  NOR2_X1 U5413 ( .A1(n7109), .A2(n4624), .ZN(n6256) );
  NOR2_X1 U5414 ( .A1(n6324), .A2(n6255), .ZN(n4624) );
  NOR2_X1 U5415 ( .A1(n7713), .A2(n6288), .ZN(n6289) );
  INV_X1 U5416 ( .A(n6287), .ZN(n6288) );
  INV_X1 U5417 ( .A(n8497), .ZN(n4632) );
  AND2_X1 U5418 ( .A1(n8500), .A2(n6299), .ZN(n6300) );
  NAND2_X1 U5419 ( .A1(n5558), .A2(n5557), .ZN(n8425) );
  NAND2_X1 U5420 ( .A1(n4605), .A2(n4328), .ZN(n5558) );
  NAND2_X1 U5421 ( .A1(n4325), .A2(n4689), .ZN(n4688) );
  OR2_X1 U5422 ( .A1(n5313), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5332) );
  NOR2_X1 U5423 ( .A1(n9646), .A2(n8452), .ZN(n4705) );
  INV_X1 U5424 ( .A(n9646), .ZN(n4704) );
  NAND2_X1 U5425 ( .A1(n7578), .A2(n4681), .ZN(n4680) );
  NAND2_X1 U5426 ( .A1(n7546), .A2(n8260), .ZN(n7635) );
  NAND2_X1 U5427 ( .A1(n5118), .A2(n5117), .ZN(n5150) );
  INV_X1 U5428 ( .A(n5119), .ZN(n5118) );
  INV_X1 U5429 ( .A(n8392), .ZN(n4588) );
  NAND2_X1 U5430 ( .A1(n5089), .A2(n5090), .ZN(n8253) );
  AND2_X1 U5431 ( .A1(n8248), .A2(n8247), .ZN(n8389) );
  NAND2_X1 U5432 ( .A1(n8227), .A2(n8226), .ZN(n8381) );
  OR2_X1 U5433 ( .A1(n7992), .A2(n8677), .ZN(n8663) );
  NOR2_X1 U5434 ( .A1(n4315), .A2(n4592), .ZN(n4591) );
  INV_X1 U5435 ( .A(n4597), .ZN(n4592) );
  OAI21_X1 U5436 ( .B1(n4320), .B2(n4315), .A(n8303), .ZN(n4595) );
  AND2_X1 U5437 ( .A1(n5607), .A2(n6235), .ZN(n7009) );
  NAND2_X1 U5438 ( .A1(n4496), .A2(n5608), .ZN(n4495) );
  INV_X1 U5439 ( .A(n4497), .ZN(n4496) );
  INV_X1 U5440 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5268) );
  OR2_X1 U5441 ( .A1(n5072), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U5442 ( .A1(n4327), .A2(n5913), .ZN(n4711) );
  NOR2_X1 U5443 ( .A1(n4712), .A2(n4439), .ZN(n4438) );
  INV_X1 U5444 ( .A(n8939), .ZN(n4439) );
  NOR2_X1 U5445 ( .A1(n4712), .A2(n6022), .ZN(n4437) );
  INV_X1 U5446 ( .A(n8833), .ZN(n4447) );
  INV_X1 U5447 ( .A(n4828), .ZN(n4826) );
  NOR2_X1 U5448 ( .A1(n4830), .A2(n4823), .ZN(n4822) );
  INV_X1 U5449 ( .A(n9135), .ZN(n4823) );
  NAND2_X1 U5450 ( .A1(n6368), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6408) );
  OR2_X1 U5451 ( .A1(n9536), .A2(n6478), .ZN(n9155) );
  NOR2_X1 U5452 ( .A1(n9546), .A2(n4574), .ZN(n4573) );
  INV_X1 U5453 ( .A(n4575), .ZN(n4574) );
  INV_X1 U5454 ( .A(n6128), .ZN(n6129) );
  NAND2_X1 U5455 ( .A1(n6129), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6142) );
  INV_X1 U5456 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9396) );
  OR3_X1 U5457 ( .A1(n6459), .A2(n6458), .A3(n7317), .ZN(n6526) );
  AND2_X1 U5458 ( .A1(n6565), .A2(n6560), .ZN(n6533) );
  NOR2_X1 U5459 ( .A1(n9853), .A2(n7324), .ZN(n7325) );
  NAND2_X1 U5460 ( .A1(n7279), .A2(n7287), .ZN(n7300) );
  NOR2_X1 U5461 ( .A1(n9887), .A2(n4269), .ZN(n7279) );
  NOR2_X1 U5462 ( .A1(n9515), .A2(n9481), .ZN(n4565) );
  NAND2_X1 U5463 ( .A1(n9449), .A2(n9092), .ZN(n9450) );
  INV_X1 U5464 ( .A(n6583), .ZN(n9662) );
  NOR2_X1 U5465 ( .A1(n7615), .A2(n6463), .ZN(n7693) );
  NAND2_X1 U5466 ( .A1(n4760), .A2(n4758), .ZN(n5505) );
  AOI21_X1 U5467 ( .B1(n4762), .B2(n4764), .A(n4759), .ZN(n4758) );
  INV_X1 U5468 ( .A(n5491), .ZN(n4759) );
  AND2_X1 U5469 ( .A1(n5471), .A2(n5458), .ZN(n5469) );
  OR2_X1 U5470 ( .A1(n5428), .A2(n5432), .ZN(n5434) );
  AND2_X1 U5471 ( .A1(n5454), .A2(n5439), .ZN(n5452) );
  OR2_X1 U5472 ( .A1(n5409), .A2(n5408), .ZN(n5430) );
  NAND2_X1 U5473 ( .A1(n5351), .A2(n5350), .ZN(n4773) );
  INV_X1 U5474 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5640) );
  NOR2_X1 U5475 ( .A1(n4767), .A2(n4771), .ZN(n4766) );
  INV_X1 U5476 ( .A(n5219), .ZN(n4771) );
  INV_X1 U5477 ( .A(n5206), .ZN(n4767) );
  INV_X1 U5478 ( .A(n5213), .ZN(n4770) );
  NAND2_X1 U5479 ( .A1(n5175), .A2(SI_12_), .ZN(n5200) );
  XNOR2_X1 U5480 ( .A(n5172), .B(SI_11_), .ZN(n5173) );
  CLKBUF_X1 U5481 ( .A(n4302), .Z(n5804) );
  AND2_X1 U5482 ( .A1(n8021), .A2(n8019), .ZN(n8132) );
  INV_X1 U5483 ( .A(n7598), .ZN(n4857) );
  NAND2_X1 U5484 ( .A1(n7597), .A2(n7596), .ZN(n4858) );
  INV_X1 U5485 ( .A(n7365), .ZN(n4881) );
  AND2_X1 U5486 ( .A1(n7015), .A2(n7204), .ZN(n8200) );
  NAND2_X1 U5487 ( .A1(n8348), .A2(n4321), .ZN(n4505) );
  MUX2_X1 U5488 ( .A(n8411), .B(n8421), .S(n8355), .Z(n8361) );
  NAND2_X1 U5489 ( .A1(n4507), .A2(n4508), .ZN(n8363) );
  AND2_X1 U5490 ( .A1(n4485), .A2(n5559), .ZN(n4481) );
  AND2_X1 U5491 ( .A1(n8373), .A2(n8372), .ZN(n8418) );
  AND4_X1 U5492 ( .A1(n5098), .A2(n5097), .A3(n5096), .A4(n5095), .ZN(n7364)
         );
  NOR2_X1 U5493 ( .A1(n6941), .A2(n6942), .ZN(n6940) );
  NAND2_X1 U5494 ( .A1(n7041), .A2(n7040), .ZN(n7039) );
  NOR2_X1 U5495 ( .A1(n7038), .A2(n7037), .ZN(n7036) );
  NAND2_X1 U5496 ( .A1(n4626), .A2(n4625), .ZN(n6966) );
  NAND2_X1 U5497 ( .A1(n6251), .A2(n4628), .ZN(n4625) );
  NAND2_X1 U5498 ( .A1(n6914), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6960) );
  AND2_X1 U5499 ( .A1(n4730), .A2(n7100), .ZN(n7054) );
  NAND2_X1 U5500 ( .A1(n7054), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7102) );
  AOI21_X1 U5501 ( .B1(n7107), .B2(n7105), .A(n7106), .ZN(n7109) );
  NAND2_X1 U5502 ( .A1(n7050), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7107) );
  XNOR2_X1 U5503 ( .A(n6256), .B(n7178), .ZN(n7176) );
  AOI21_X1 U5504 ( .B1(n7175), .B2(n4318), .A(n7240), .ZN(n7239) );
  NAND2_X1 U5505 ( .A1(n7176), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7175) );
  OR2_X1 U5506 ( .A1(n5103), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5113) );
  NOR2_X1 U5507 ( .A1(n7704), .A2(n6261), .ZN(n6262) );
  OAI21_X1 U5508 ( .B1(n7802), .B2(n4743), .A(n4742), .ZN(n7886) );
  NAND2_X1 U5509 ( .A1(n6292), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4743) );
  NAND2_X1 U5510 ( .A1(n6290), .A2(n6292), .ZN(n4742) );
  NOR2_X1 U5511 ( .A1(n7802), .A2(n9300), .ZN(n7801) );
  NAND2_X1 U5512 ( .A1(n4405), .A2(n4632), .ZN(n4631) );
  NAND2_X1 U5513 ( .A1(n4786), .A2(n4785), .ZN(n8514) );
  INV_X1 U5514 ( .A(n8511), .ZN(n4785) );
  AOI21_X1 U5515 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n6859), .A(n8474), .ZN(
        n6296) );
  OR2_X1 U5516 ( .A1(n5495), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U5517 ( .A1(n5479), .A2(n8028), .ZN(n5495) );
  INV_X1 U5518 ( .A(n5480), .ZN(n5479) );
  NAND2_X1 U5519 ( .A1(n5443), .A2(n5442), .ZN(n5461) );
  INV_X1 U5520 ( .A(n5444), .ZN(n5443) );
  NAND2_X1 U5521 ( .A1(n5359), .A2(n5358), .ZN(n5378) );
  INV_X1 U5522 ( .A(n5360), .ZN(n5359) );
  NAND2_X1 U5523 ( .A1(n5291), .A2(n10034), .ZN(n5313) );
  INV_X1 U5524 ( .A(n5292), .ZN(n5291) );
  NAND2_X1 U5525 ( .A1(n5250), .A2(n5249), .ZN(n5278) );
  NAND2_X1 U5526 ( .A1(n5193), .A2(n5192), .ZN(n5228) );
  INV_X1 U5527 ( .A(n5194), .ZN(n5193) );
  AND4_X1 U5528 ( .A1(n5170), .A2(n5169), .A3(n5168), .A4(n5167), .ZN(n7661)
         );
  NAND2_X1 U5529 ( .A1(n5082), .A2(n9405), .ZN(n5094) );
  INV_X1 U5530 ( .A(n5092), .ZN(n5082) );
  NAND2_X1 U5531 ( .A1(n5030), .A2(n5029), .ZN(n5051) );
  INV_X1 U5532 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5029) );
  INV_X1 U5533 ( .A(n5031), .ZN(n5030) );
  NAND2_X1 U5534 ( .A1(n7224), .A2(n5009), .ZN(n5031) );
  INV_X1 U5535 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5009) );
  NAND2_X1 U5536 ( .A1(n7144), .A2(n8224), .ZN(n7143) );
  AND2_X1 U5537 ( .A1(n6928), .A2(n5560), .ZN(n7637) );
  AND2_X1 U5538 ( .A1(n7002), .A2(n6230), .ZN(n6925) );
  AND2_X1 U5539 ( .A1(n7204), .A2(n4275), .ZN(n8653) );
  INV_X1 U5540 ( .A(n8325), .ZN(n8604) );
  AOI21_X1 U5541 ( .B1(n4694), .B2(n4697), .A(n4692), .ZN(n4691) );
  NAND2_X1 U5542 ( .A1(n8652), .A2(n4694), .ZN(n4693) );
  INV_X1 U5543 ( .A(n8615), .ZN(n4692) );
  AOI21_X1 U5544 ( .B1(n4603), .B2(n4701), .A(n4602), .ZN(n4601) );
  AND3_X1 U5545 ( .A1(n5070), .A2(n5069), .A3(n5068), .ZN(n10046) );
  OR2_X1 U5546 ( .A1(n6973), .A2(n8439), .ZN(n10069) );
  NAND2_X1 U5547 ( .A1(n7554), .A2(n10069), .ZN(n10049) );
  OR2_X1 U5548 ( .A1(n6228), .A2(n8355), .ZN(n7007) );
  AND2_X1 U5549 ( .A1(n7009), .A2(n8437), .ZN(n7013) );
  AND2_X1 U5550 ( .A1(n6999), .A2(n7118), .ZN(n8437) );
  NOR2_X1 U5551 ( .A1(n4923), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n4889) );
  NOR2_X1 U5552 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4623) );
  INV_X1 U5553 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4915) );
  INV_X1 U5554 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4914) );
  INV_X1 U5555 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5066) );
  INV_X1 U5556 ( .A(n6142), .ZN(n6143) );
  XNOR2_X1 U5557 ( .A(n5694), .B(n6173), .ZN(n5698) );
  NAND2_X1 U5558 ( .A1(n5692), .A2(n4426), .ZN(n5694) );
  NAND2_X1 U5559 ( .A1(n5769), .A2(n4314), .ZN(n4426) );
  NOR2_X1 U5560 ( .A1(n5798), .A2(n4725), .ZN(n4724) );
  INV_X1 U5561 ( .A(n5780), .ZN(n4725) );
  NAND2_X1 U5562 ( .A1(n8975), .A2(n6421), .ZN(n5710) );
  NOR2_X1 U5563 ( .A1(n6108), .A2(n9387), .ZN(n6110) );
  NAND2_X1 U5564 ( .A1(n6105), .A2(n4714), .ZN(n4713) );
  OR2_X1 U5565 ( .A1(n6104), .A2(n8847), .ZN(n4894) );
  NAND2_X1 U5566 ( .A1(n4461), .A2(n4460), .ZN(n6105) );
  NAND2_X1 U5567 ( .A1(n8904), .A2(n8905), .ZN(n8832) );
  NAND2_X1 U5568 ( .A1(n4433), .A2(n6901), .ZN(n4430) );
  INV_X1 U5569 ( .A(n6834), .ZN(n6708) );
  AND2_X1 U5570 ( .A1(n4561), .A2(n4444), .ZN(n4558) );
  AND2_X1 U5571 ( .A1(n6700), .A2(n6644), .ZN(n4561) );
  NOR2_X1 U5572 ( .A1(n4413), .A2(n4560), .ZN(n4559) );
  INV_X1 U5573 ( .A(n6637), .ZN(n4560) );
  OR2_X1 U5574 ( .A1(n6509), .A2(n5701), .ZN(n5702) );
  OR2_X1 U5575 ( .A1(n6412), .A2(n5700), .ZN(n5704) );
  AOI21_X1 U5576 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n6797), .A(n9702), .ZN(
        n9715) );
  AOI21_X1 U5577 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6803), .A(n9610), .ZN(
        n9627) );
  AOI21_X1 U5578 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9602), .A(n9597), .ZN(
        n9733) );
  AOI21_X1 U5579 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9754), .A(n9749), .ZN(
        n9764) );
  NOR2_X1 U5580 ( .A1(n9049), .A2(n9780), .ZN(n9052) );
  OR2_X1 U5581 ( .A1(n9796), .A2(n9797), .ZN(n9793) );
  NAND2_X1 U5582 ( .A1(n6448), .A2(n6447), .ZN(n9510) );
  NOR2_X1 U5583 ( .A1(n9530), .A2(n9237), .ZN(n9220) );
  AND2_X1 U5584 ( .A1(n9156), .A2(n4554), .ZN(n9226) );
  AND2_X1 U5585 ( .A1(n9155), .A2(n6613), .ZN(n9246) );
  NAND2_X1 U5586 ( .A1(n9236), .A2(n9239), .ZN(n9237) );
  INV_X1 U5587 ( .A(n9246), .ZN(n9233) );
  AND2_X1 U5588 ( .A1(n9539), .A2(n9129), .ZN(n4816) );
  NAND2_X1 U5589 ( .A1(n9258), .A2(n9128), .ZN(n4817) );
  NAND2_X1 U5590 ( .A1(n9449), .A2(n4573), .ZN(n9273) );
  OR2_X1 U5591 ( .A1(n9551), .A2(n9121), .ZN(n9122) );
  OR2_X1 U5592 ( .A1(n9293), .A2(n9120), .ZN(n4901) );
  NAND2_X1 U5593 ( .A1(n9818), .A2(n4577), .ZN(n9479) );
  NOR2_X1 U5594 ( .A1(n9566), .A2(n4579), .ZN(n4577) );
  AND2_X1 U5595 ( .A1(n6597), .A2(n6598), .ZN(n9465) );
  NAND2_X1 U5596 ( .A1(n6073), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6090) );
  AND2_X1 U5597 ( .A1(n6050), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6073) );
  NOR2_X1 U5598 ( .A1(n6030), .A2(n6029), .ZN(n6050) );
  NAND2_X1 U5599 ( .A1(n9818), .A2(n4581), .ZN(n9657) );
  NAND2_X1 U5600 ( .A1(n9818), .A2(n9689), .ZN(n9655) );
  OR2_X1 U5601 ( .A1(n6012), .A2(n6011), .ZN(n6030) );
  NAND2_X1 U5602 ( .A1(n9807), .A2(n6468), .ZN(n9661) );
  AND2_X1 U5603 ( .A1(n9820), .A2(n9984), .ZN(n9818) );
  AND2_X1 U5604 ( .A1(n7693), .A2(n9977), .ZN(n9820) );
  NAND2_X1 U5605 ( .A1(n9810), .A2(n6466), .ZN(n9807) );
  NAND2_X1 U5606 ( .A1(n4843), .A2(n4849), .ZN(n4839) );
  INV_X1 U5607 ( .A(n6575), .ZN(n9808) );
  NAND2_X1 U5608 ( .A1(n7689), .A2(n4672), .ZN(n4670) );
  AND2_X1 U5609 ( .A1(n4669), .A2(n6570), .ZN(n4668) );
  OR2_X1 U5610 ( .A1(n5870), .A2(n5670), .ZN(n5901) );
  INV_X1 U5611 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5900) );
  NOR2_X1 U5612 ( .A1(n5901), .A2(n5900), .ZN(n5918) );
  INV_X1 U5613 ( .A(n6533), .ZN(n7506) );
  AOI21_X1 U5614 ( .B1(n7567), .B2(n4813), .A(n4370), .ZN(n4812) );
  AND2_X1 U5615 ( .A1(n9838), .A2(n9946), .ZN(n7568) );
  OR2_X1 U5616 ( .A1(n6835), .A2(n6708), .ZN(n7268) );
  AND2_X1 U5617 ( .A1(n7325), .A2(n7477), .ZN(n9838) );
  OR2_X1 U5618 ( .A1(n5831), .A2(n7450), .ZN(n5870) );
  AOI21_X1 U5619 ( .B1(n4677), .B2(n4675), .A(n4674), .ZN(n4673) );
  INV_X1 U5620 ( .A(n4677), .ZN(n4676) );
  INV_X1 U5621 ( .A(n6649), .ZN(n4675) );
  AOI21_X1 U5622 ( .B1(n7309), .B2(n4807), .A(n4378), .ZN(n4805) );
  INV_X1 U5623 ( .A(n7292), .ZN(n4807) );
  NAND2_X1 U5624 ( .A1(n4562), .A2(n7311), .ZN(n9853) );
  INV_X1 U5625 ( .A(n9869), .ZN(n4562) );
  NOR2_X1 U5626 ( .A1(n5782), .A2(n7168), .ZN(n5809) );
  OR2_X1 U5627 ( .A1(n7300), .A2(n7299), .ZN(n9869) );
  NAND2_X1 U5628 ( .A1(n6731), .A2(n6729), .ZN(n7266) );
  NAND2_X1 U5629 ( .A1(n6385), .A2(n6384), .ZN(n9521) );
  INV_X1 U5630 ( .A(n9983), .ZN(n9933) );
  OAI21_X1 U5631 ( .B1(n7264), .B2(P1_D_REG_0__SCAN_IN), .A(n9584), .ZN(n7307)
         );
  AND2_X1 U5632 ( .A1(n7521), .A2(n9904), .ZN(n9937) );
  NAND2_X1 U5633 ( .A1(n9586), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5669) );
  XNOR2_X1 U5634 ( .A(n5490), .B(n5489), .ZN(n7827) );
  NAND2_X1 U5635 ( .A1(n4761), .A2(n5471), .ZN(n5490) );
  NAND2_X1 U5636 ( .A1(n5470), .A2(n5469), .ZN(n4761) );
  AND2_X1 U5637 ( .A1(n5655), .A2(n5654), .ZN(n6188) );
  XNOR2_X1 U5638 ( .A(n5470), .B(n5469), .ZN(n7793) );
  XNOR2_X1 U5639 ( .A(n5657), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6184) );
  AND2_X1 U5640 ( .A1(n5661), .A2(n5660), .ZN(n6185) );
  XNOR2_X1 U5641 ( .A(n5648), .B(n5644), .ZN(n6837) );
  NAND2_X1 U5642 ( .A1(n4727), .A2(n4347), .ZN(n5648) );
  NAND2_X1 U5643 ( .A1(n5287), .A2(n5286), .ZN(n5302) );
  AND2_X1 U5644 ( .A1(n5286), .A2(n5263), .ZN(n5264) );
  NAND2_X1 U5645 ( .A1(n4765), .A2(n4768), .ZN(n5243) );
  AOI21_X1 U5646 ( .B1(n5219), .B2(n4770), .A(n4769), .ZN(n4768) );
  NAND2_X1 U5647 ( .A1(n5207), .A2(n4766), .ZN(n4765) );
  INV_X1 U5648 ( .A(n5236), .ZN(n4769) );
  AND2_X1 U5649 ( .A1(n5258), .A2(n5241), .ZN(n5242) );
  AND2_X1 U5650 ( .A1(n5214), .A2(n4527), .ZN(n6828) );
  OAI21_X1 U5651 ( .B1(n5175), .B2(SI_12_), .A(n5200), .ZN(n5176) );
  AND2_X1 U5652 ( .A1(n5955), .A2(n5939), .ZN(n9045) );
  INV_X1 U5653 ( .A(n4750), .ZN(n4530) );
  OAI21_X1 U5654 ( .B1(n5100), .B2(n4755), .A(n4753), .ZN(n5137) );
  AND2_X1 U5655 ( .A1(n5080), .A2(n5079), .ZN(n5099) );
  NAND2_X1 U5656 ( .A1(n5100), .A2(n5099), .ZN(n5102) );
  AND2_X1 U5657 ( .A1(n5074), .A2(n5062), .ZN(n5063) );
  AND2_X1 U5658 ( .A1(n5057), .A2(n5045), .ZN(n5046) );
  NAND2_X1 U5659 ( .A1(n5024), .A2(n5023), .ZN(n5041) );
  AND2_X1 U5660 ( .A1(n5762), .A2(n5761), .ZN(n5764) );
  OR2_X1 U5661 ( .A1(n4521), .A2(SI_2_), .ZN(n4520) );
  AND4_X1 U5662 ( .A1(n5056), .A2(n5055), .A3(n5054), .A4(n5053), .ZN(n7378)
         );
  XNOR2_X1 U5663 ( .A(n8048), .B(n8444), .ZN(n8035) );
  AND2_X1 U5664 ( .A1(n5385), .A2(n5384), .ZN(n8620) );
  AOI21_X1 U5665 ( .B1(n4868), .B2(n4317), .A(n4867), .ZN(n4866) );
  NAND2_X1 U5666 ( .A1(n6981), .A2(n6980), .ZN(n6982) );
  NAND2_X1 U5667 ( .A1(n8143), .A2(n8144), .ZN(n4861) );
  AND2_X1 U5668 ( .A1(n5181), .A2(n5180), .ZN(n10080) );
  NAND2_X1 U5669 ( .A1(n8094), .A2(n8096), .ZN(n8095) );
  INV_X1 U5670 ( .A(n8460), .ZN(n7160) );
  INV_X1 U5671 ( .A(n4893), .ZN(n4869) );
  INV_X1 U5672 ( .A(n4876), .ZN(n7155) );
  AND2_X1 U5673 ( .A1(n7119), .A2(n8441), .ZN(n8031) );
  AND2_X1 U5674 ( .A1(n4858), .A2(n7594), .ZN(n7599) );
  NAND2_X1 U5675 ( .A1(n4858), .A2(n4856), .ZN(n7833) );
  NAND2_X1 U5676 ( .A1(n8095), .A2(n7983), .ZN(n8150) );
  NAND2_X1 U5677 ( .A1(n4860), .A2(n4859), .ZN(n8162) );
  AOI21_X1 U5678 ( .B1(n4862), .B2(n4864), .A(n4377), .ZN(n4859) );
  OAI21_X1 U5679 ( .B1(n8184), .B2(n8183), .A(n8182), .ZN(n8186) );
  INV_X1 U5680 ( .A(n8195), .ZN(n8185) );
  OR2_X1 U5681 ( .A1(n7014), .A2(n7204), .ZN(n8202) );
  NOR2_X1 U5682 ( .A1(n8196), .A2(n4873), .ZN(n4872) );
  INV_X1 U5683 ( .A(n7989), .ZN(n4873) );
  NAND2_X1 U5684 ( .A1(n4874), .A2(n7989), .ZN(n8197) );
  INV_X1 U5685 ( .A(n8031), .ZN(n8204) );
  INV_X1 U5686 ( .A(n8564), .ZN(n8444) );
  NAND2_X1 U5687 ( .A1(n5402), .A2(n5401), .ZN(n8607) );
  INV_X1 U5688 ( .A(n8620), .ZN(n8447) );
  INV_X1 U5689 ( .A(n8156), .ZN(n8453) );
  INV_X1 U5690 ( .A(n7378), .ZN(n8458) );
  INV_X1 U5691 ( .A(P2_U3893), .ZN(n8463) );
  AOI21_X1 U5692 ( .B1(n7243), .B2(n4735), .A(n4415), .ZN(n4733) );
  INV_X1 U5693 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n4735) );
  NAND2_X1 U5694 ( .A1(n4799), .A2(n4798), .ZN(n7344) );
  XNOR2_X1 U5695 ( .A(n6286), .B(n6769), .ZN(n7342) );
  XOR2_X1 U5696 ( .A(n6820), .B(n6262), .Z(n7800) );
  INV_X1 U5697 ( .A(n4794), .ZN(n7855) );
  INV_X1 U5698 ( .A(n4747), .ZN(n7863) );
  OR2_X1 U5699 ( .A1(n7856), .A2(n9650), .ZN(n4794) );
  INV_X1 U5700 ( .A(n6265), .ZN(n4793) );
  INV_X1 U5701 ( .A(n6294), .ZN(n4746) );
  NAND2_X1 U5702 ( .A1(n4795), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4792) );
  INV_X1 U5703 ( .A(n8466), .ZN(n4795) );
  OR2_X1 U5704 ( .A1(n8503), .A2(n8502), .ZN(n8500) );
  AOI21_X1 U5705 ( .B1(n10022), .B2(n10021), .A(n10020), .ZN(n10029) );
  INV_X1 U5706 ( .A(n10017), .ZN(n10022) );
  OAI21_X1 U5707 ( .B1(n8537), .B2(n10026), .A(n4802), .ZN(n4801) );
  NAND2_X1 U5708 ( .A1(n4608), .A2(n8345), .ZN(n7971) );
  NAND2_X1 U5709 ( .A1(n4616), .A2(n4614), .ZN(n4608) );
  NAND2_X1 U5710 ( .A1(n7968), .A2(n7967), .ZN(n7969) );
  XNOR2_X1 U5711 ( .A(n7966), .B(n8407), .ZN(n7970) );
  NAND2_X1 U5712 ( .A1(n8445), .A2(n8655), .ZN(n7967) );
  NAND2_X1 U5713 ( .A1(n5357), .A2(n5356), .ZN(n8624) );
  NAND2_X1 U5714 ( .A1(n4698), .A2(n4699), .ZN(n8628) );
  NAND2_X1 U5715 ( .A1(n5344), .A2(n5343), .ZN(n8731) );
  AOI21_X1 U5716 ( .B1(n8652), .B2(n5319), .A(n4345), .ZN(n8642) );
  NAND2_X1 U5717 ( .A1(n5248), .A2(n5247), .ZN(n8748) );
  AND2_X1 U5718 ( .A1(n5227), .A2(n5226), .ZN(n9640) );
  NAND2_X1 U5719 ( .A1(n4599), .A2(n8285), .ZN(n7897) );
  NAND2_X1 U5720 ( .A1(n7658), .A2(n8281), .ZN(n7748) );
  INV_X1 U5721 ( .A(n10080), .ZN(n7664) );
  OAI21_X1 U5722 ( .B1(n4683), .B2(n4679), .A(n4352), .ZN(n7579) );
  OR2_X1 U5723 ( .A1(n7458), .A2(n5534), .ZN(n4589) );
  NAND2_X1 U5724 ( .A1(n6927), .A2(n8437), .ZN(n8698) );
  INV_X1 U5725 ( .A(n8545), .ZN(n8702) );
  INV_X1 U5726 ( .A(n8698), .ZN(n8685) );
  INV_X1 U5727 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n4708) );
  OAI222_X1 U5728 ( .A1(n8695), .A2(n8564), .B1(n8693), .B2(n8584), .C1(n10037), .C2(n8563), .ZN(n8710) );
  OAI21_X1 U5729 ( .B1(n6737), .B2(n5039), .A(n4499), .ZN(n7225) );
  NOR2_X1 U5730 ( .A1(n4997), .A2(n9302), .ZN(n4501) );
  NAND2_X1 U5731 ( .A1(n4605), .A2(n4609), .ZN(n7951) );
  NAND2_X1 U5732 ( .A1(n4616), .A2(n8342), .ZN(n8560) );
  NAND2_X1 U5733 ( .A1(n5417), .A2(n5416), .ZN(n8774) );
  NAND2_X1 U5734 ( .A1(n5395), .A2(n5394), .ZN(n8780) );
  NAND2_X1 U5735 ( .A1(n5377), .A2(n5376), .ZN(n8786) );
  NAND2_X1 U5736 ( .A1(n8639), .A2(n8311), .ZN(n8627) );
  NAND2_X1 U5737 ( .A1(n5277), .A2(n5276), .ZN(n8807) );
  INV_X1 U5738 ( .A(n4593), .ZN(n8688) );
  AOI21_X1 U5739 ( .B1(n4599), .B2(n4320), .A(n4315), .ZN(n4593) );
  AND2_X1 U5740 ( .A1(n7012), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7118) );
  OR2_X1 U5741 ( .A1(n4945), .A2(n8816), .ZN(n4925) );
  NAND2_X1 U5742 ( .A1(n5577), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5579) );
  INV_X1 U5743 ( .A(n8479), .ZN(n6859) );
  INV_X1 U5744 ( .A(n6284), .ZN(n7247) );
  XNOR2_X1 U5745 ( .A(n5017), .B(n5016), .ZN(n6972) );
  OR2_X1 U5746 ( .A1(n4954), .A2(n4788), .ZN(n4787) );
  NAND2_X1 U5747 ( .A1(n8816), .A2(n4790), .ZN(n4789) );
  NAND2_X1 U5748 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4788) );
  NAND2_X1 U5749 ( .A1(n4956), .A2(n4955), .ZN(n6952) );
  MUX2_X1 U5750 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4953), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n4956) );
  AND2_X1 U5751 ( .A1(n4461), .A2(n4463), .ZN(n8850) );
  AOI21_X1 U5752 ( .B1(n6364), .B2(P2_DATAO_REG_19__SCAN_IN), .A(n4443), .ZN(
        n6088) );
  NOR2_X1 U5753 ( .A1(n6755), .A2(n7232), .ZN(n4443) );
  OR2_X1 U5754 ( .A1(n6442), .A2(n6441), .ZN(n6443) );
  NAND2_X1 U5755 ( .A1(n6436), .A2(n6435), .ZN(n6437) );
  AOI21_X1 U5756 ( .B1(n4457), .B2(n4459), .A(n4383), .ZN(n4455) );
  INV_X1 U5757 ( .A(n4460), .ZN(n4459) );
  NAND2_X1 U5758 ( .A1(n8876), .A2(n8877), .ZN(n8875) );
  NAND2_X1 U5759 ( .A1(n8938), .A2(n6023), .ZN(n8876) );
  INV_X1 U5760 ( .A(n4713), .ZN(n8897) );
  NAND2_X1 U5761 ( .A1(n7728), .A2(n4327), .ZN(n7732) );
  NAND2_X1 U5762 ( .A1(n4514), .A2(n4369), .ZN(n8925) );
  NAND2_X1 U5763 ( .A1(n4516), .A2(n4515), .ZN(n4513) );
  AND2_X1 U5764 ( .A1(n4440), .A2(n6023), .ZN(n8940) );
  INV_X1 U5765 ( .A(n8918), .ZN(n8948) );
  NAND2_X1 U5766 ( .A1(n8983), .A2(n8988), .ZN(n8982) );
  NAND2_X1 U5767 ( .A1(n9012), .A2(n9013), .ZN(n9011) );
  AOI21_X1 U5768 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9059), .A(n9057), .ZN(
        n9073) );
  NAND2_X1 U5769 ( .A1(n9095), .A2(n9888), .ZN(n9505) );
  NAND2_X1 U5770 ( .A1(n6502), .A2(n6501), .ZN(n9105) );
  XNOR2_X1 U5771 ( .A(n9141), .B(n9163), .ZN(n9513) );
  INV_X1 U5772 ( .A(n9511), .ZN(n9509) );
  NAND2_X1 U5773 ( .A1(n4645), .A2(n4647), .ZN(n9180) );
  NAND2_X1 U5774 ( .A1(n4833), .A2(n4829), .ZN(n4831) );
  NOR2_X1 U5775 ( .A1(n4827), .A2(n9134), .ZN(n9203) );
  INV_X1 U5776 ( .A(n4835), .ZN(n4827) );
  OAI21_X1 U5777 ( .B1(n9284), .B2(n4654), .A(n4652), .ZN(n9261) );
  NOR2_X1 U5778 ( .A1(n9282), .A2(n9151), .ZN(n9269) );
  OR2_X1 U5779 ( .A1(n6895), .A2(n5888), .ZN(n6010) );
  OR2_X1 U5780 ( .A1(n6858), .A2(n5888), .ZN(n5988) );
  NAND2_X1 U5781 ( .A1(n5958), .A2(n5957), .ZN(n7696) );
  NAND2_X1 U5782 ( .A1(n4524), .A2(n5214), .ZN(n5958) );
  AND2_X1 U5783 ( .A1(n4527), .A2(n6500), .ZN(n4524) );
  NAND2_X1 U5784 ( .A1(n4842), .A2(n4845), .ZN(n7786) );
  INV_X1 U5785 ( .A(n4844), .ZN(n4845) );
  NAND2_X1 U5786 ( .A1(n7613), .A2(n4846), .ZN(n4842) );
  NAND2_X1 U5787 ( .A1(n7488), .A2(n6566), .ZN(n7607) );
  AOI21_X1 U5788 ( .B1(n7613), .B2(n7612), .A(n4848), .ZN(n7690) );
  NAND2_X1 U5789 ( .A1(n5899), .A2(n5898), .ZN(n7512) );
  NAND2_X1 U5790 ( .A1(n9824), .A2(n9830), .ZN(n4815) );
  INV_X1 U5791 ( .A(n9879), .ZN(n9847) );
  OR2_X1 U5792 ( .A1(n9896), .A2(n7280), .ZN(n9883) );
  INV_X1 U5793 ( .A(n4531), .ZN(n4532) );
  INV_X1 U5794 ( .A(n9883), .ZN(n9835) );
  NAND2_X1 U5795 ( .A1(n7265), .A2(n7264), .ZN(n9901) );
  XNOR2_X1 U5796 ( .A(n6519), .B(n6518), .ZN(n9591) );
  INV_X1 U5797 ( .A(n6184), .ZN(n7727) );
  XNOR2_X1 U5798 ( .A(n5650), .B(n5649), .ZN(n7533) );
  OAI21_X1 U5799 ( .B1(n6046), .B2(n4728), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5650) );
  NAND2_X1 U5800 ( .A1(n4347), .A2(n5644), .ZN(n4728) );
  INV_X1 U5801 ( .A(n6837), .ZN(n7471) );
  NAND2_X1 U5802 ( .A1(n5306), .A2(n5321), .ZN(n7093) );
  NAND2_X1 U5803 ( .A1(n4778), .A2(n4777), .ZN(n5321) );
  NAND2_X1 U5804 ( .A1(n4448), .A2(n4452), .ZN(n6070) );
  OR2_X1 U5805 ( .A1(n5639), .A2(n5892), .ZN(n4448) );
  OAI21_X1 U5806 ( .B1(n5220), .B2(n5219), .A(n5237), .ZN(n6858) );
  NAND2_X1 U5807 ( .A1(n5220), .A2(n5219), .ZN(n5237) );
  NAND2_X1 U5808 ( .A1(n5214), .A2(n5213), .ZN(n5220) );
  INV_X1 U5809 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6771) );
  NOR2_X2 U5810 ( .A1(n6999), .A2(n7915), .ZN(P2_U3893) );
  NAND2_X1 U5811 ( .A1(n4478), .A2(n4421), .ZN(n4473) );
  AND2_X1 U5812 ( .A1(n4799), .A2(n4797), .ZN(n7706) );
  NAND2_X1 U5813 ( .A1(n4737), .A2(n7183), .ZN(n4736) );
  NAND2_X1 U5814 ( .A1(n4709), .A2(n4706), .ZN(P2_U3486) );
  AOI21_X1 U5815 ( .B1(n8556), .B2(n8744), .A(n4707), .ZN(n4706) );
  NAND2_X1 U5816 ( .A1(n7973), .A2(n10103), .ZN(n4709) );
  NOR2_X1 U5817 ( .A1(n10103), .A2(n4708), .ZN(n4707) );
  NOR2_X1 U5818 ( .A1(n5619), .A2(n5620), .ZN(n5621) );
  NAND2_X1 U5819 ( .A1(n7975), .A2(n7974), .ZN(n7976) );
  NAND2_X1 U5820 ( .A1(n10087), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7974) );
  NAND2_X1 U5821 ( .A1(n8865), .A2(n4429), .ZN(n8873) );
  MUX2_X1 U5822 ( .A(n9088), .B(n9089), .S(n7232), .Z(n9091) );
  NAND2_X1 U5823 ( .A1(n4418), .A2(n4406), .ZN(P1_U3551) );
  NAND2_X1 U5824 ( .A1(n4419), .A2(n10008), .ZN(n4418) );
  NAND2_X1 U5825 ( .A1(n4659), .A2(n4420), .ZN(n4419) );
  OAI211_X1 U5826 ( .C1(n9171), .C2(n4410), .A(n4658), .B(n4656), .ZN(P1_U3519) );
  NAND2_X1 U5827 ( .A1(n4899), .A2(n9991), .ZN(n4658) );
  INV_X1 U5828 ( .A(n4657), .ZN(n4656) );
  AND2_X1 U5829 ( .A1(n8292), .A2(n4596), .ZN(n4315) );
  AND2_X1 U5830 ( .A1(n4713), .A2(n6120), .ZN(n4316) );
  INV_X2 U5831 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5892) );
  NOR2_X1 U5832 ( .A1(n4893), .A2(n4389), .ZN(n4317) );
  OR2_X1 U5833 ( .A1(n6256), .A2(n6328), .ZN(n4318) );
  AND2_X1 U5834 ( .A1(n8292), .A2(n8285), .ZN(n4320) );
  AND2_X1 U5835 ( .A1(n4354), .A2(n4506), .ZN(n4321) );
  AND2_X1 U5836 ( .A1(n4511), .A2(n4506), .ZN(n4322) );
  AND2_X1 U5837 ( .A1(n5638), .A2(n4454), .ZN(n4323) );
  OR2_X1 U5838 ( .A1(n8767), .A2(n5451), .ZN(n4324) );
  AND2_X1 U5839 ( .A1(n4324), .A2(n5468), .ZN(n4325) );
  INV_X1 U5840 ( .A(n8319), .ZN(n4602) );
  INV_X1 U5841 ( .A(n8858), .ZN(n4717) );
  AND2_X1 U5842 ( .A1(n5548), .A2(n4603), .ZN(n4326) );
  AND2_X1 U5843 ( .A1(n7729), .A2(n7735), .ZN(n4327) );
  AND2_X1 U5844 ( .A1(n4384), .A2(n4609), .ZN(n4328) );
  AND2_X1 U5845 ( .A1(n6638), .A2(n7232), .ZN(n4329) );
  INV_X1 U5846 ( .A(n9566), .ZN(n9485) );
  OR2_X1 U5847 ( .A1(n8858), .A2(n4715), .ZN(n4330) );
  OR2_X1 U5848 ( .A1(n4687), .A2(n8582), .ZN(n4331) );
  OR2_X1 U5849 ( .A1(n4470), .A2(n4353), .ZN(n4332) );
  AND2_X1 U5850 ( .A1(n4348), .A2(n8524), .ZN(n4333) );
  NAND2_X1 U5851 ( .A1(n4850), .A2(n6464), .ZN(n4334) );
  AND2_X1 U5852 ( .A1(n4881), .A2(n4880), .ZN(n4335) );
  OR2_X1 U5853 ( .A1(n9515), .A2(n9168), .ZN(n9161) );
  NOR2_X1 U5854 ( .A1(n7705), .A2(n10094), .ZN(n4336) );
  AND2_X1 U5855 ( .A1(n4631), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4337) );
  AND2_X1 U5856 ( .A1(n4910), .A2(n7243), .ZN(n4338) );
  NAND2_X1 U5857 ( .A1(n9539), .A2(n9128), .ZN(n4340) );
  AND2_X1 U5858 ( .A1(n9191), .A2(n9192), .ZN(n4341) );
  OR2_X1 U5859 ( .A1(n8497), .A2(n6266), .ZN(n4342) );
  AND2_X1 U5860 ( .A1(n4698), .A2(n4696), .ZN(n4343) );
  OR2_X1 U5861 ( .A1(n5523), .A2(n4497), .ZN(n4344) );
  NAND2_X1 U5862 ( .A1(n4954), .A2(n4790), .ZN(n4975) );
  AND4_X1 U5863 ( .A1(n4993), .A2(n4992), .A3(n4991), .A4(n4990), .ZN(n7146)
         );
  AND2_X1 U5864 ( .A1(n8662), .A2(n8449), .ZN(n4345) );
  INV_X1 U5865 ( .A(n5769), .ZN(n5959) );
  AND2_X1 U5866 ( .A1(n4646), .A2(n4341), .ZN(n4346) );
  AND2_X1 U5867 ( .A1(n5643), .A2(n4729), .ZN(n4347) );
  NAND2_X1 U5868 ( .A1(n5541), .A2(n8692), .ZN(n8292) );
  NOR2_X1 U5869 ( .A1(n10017), .A2(n6270), .ZN(n4348) );
  OR2_X1 U5870 ( .A1(n6200), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4349) );
  NAND2_X1 U5871 ( .A1(n4622), .A2(n4618), .ZN(n4926) );
  OR2_X1 U5872 ( .A1(n7839), .A2(n8455), .ZN(n4350) );
  OR2_X1 U5873 ( .A1(n9146), .A2(n9983), .ZN(n4351) );
  NAND2_X1 U5874 ( .A1(n4512), .A2(n4516), .ZN(n8865) );
  OR2_X1 U5875 ( .A1(n10068), .A2(n7581), .ZN(n4352) );
  NAND2_X1 U5876 ( .A1(n9127), .A2(n9126), .ZN(n9253) );
  XOR2_X1 U5877 ( .A(n9646), .B(n8452), .Z(n4353) );
  AND2_X1 U5878 ( .A1(n4511), .A2(n8374), .ZN(n4354) );
  NAND2_X1 U5879 ( .A1(n8351), .A2(n4509), .ZN(n4355) );
  AND2_X1 U5880 ( .A1(n6972), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4356) );
  NAND2_X1 U5881 ( .A1(n6140), .A2(n6139), .ZN(n9539) );
  OR2_X1 U5882 ( .A1(n8244), .A2(n8245), .ZN(n4357) );
  XNOR2_X1 U5883 ( .A(n6137), .B(n4720), .ZN(n8904) );
  NAND2_X1 U5884 ( .A1(n6405), .A2(n6404), .ZN(n9515) );
  NOR2_X1 U5885 ( .A1(n5523), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U5886 ( .A1(n6360), .A2(n6359), .ZN(n9530) );
  NAND2_X1 U5887 ( .A1(n4519), .A2(n6182), .ZN(n6358) );
  OR2_X1 U5888 ( .A1(n8753), .A2(n8539), .ZN(n4358) );
  AND2_X1 U5889 ( .A1(n9176), .A2(n9093), .ZN(n4359) );
  AND2_X1 U5890 ( .A1(n8290), .A2(n4332), .ZN(n4360) );
  NAND2_X1 U5891 ( .A1(n5386), .A2(n8325), .ZN(n8602) );
  NAND2_X1 U5892 ( .A1(n5985), .A2(n5630), .ZN(n5645) );
  AND4_X1 U5893 ( .A1(n5088), .A2(n5087), .A3(n5086), .A4(n5085), .ZN(n7592)
         );
  INV_X1 U5894 ( .A(n7592), .ZN(n5090) );
  NOR2_X1 U5895 ( .A1(n4906), .A2(n8011), .ZN(n4361) );
  AND2_X1 U5896 ( .A1(n4460), .A2(n4458), .ZN(n4362) );
  AND2_X1 U5897 ( .A1(n4645), .A2(n4643), .ZN(n4363) );
  AND2_X1 U5898 ( .A1(n6124), .A2(n6123), .ZN(n4364) );
  INV_X1 U5899 ( .A(n9546), .ZN(n9278) );
  NOR2_X1 U5900 ( .A1(n8848), .A2(n6103), .ZN(n4365) );
  OR2_X1 U5901 ( .A1(n6463), .A2(n6464), .ZN(n6570) );
  AND2_X1 U5902 ( .A1(n8320), .A2(n8319), .ZN(n8629) );
  NAND2_X1 U5903 ( .A1(n10065), .A2(n8456), .ZN(n4366) );
  INV_X1 U5904 ( .A(n4697), .ZN(n4696) );
  NAND2_X1 U5905 ( .A1(n4699), .A2(n8404), .ZN(n4697) );
  INV_X1 U5906 ( .A(n4904), .ZN(n4877) );
  NOR2_X1 U5907 ( .A1(n5550), .A2(n4604), .ZN(n4603) );
  INV_X1 U5908 ( .A(n7790), .ZN(n9689) );
  NAND2_X1 U5909 ( .A1(n8663), .A2(n8402), .ZN(n4367) );
  AND2_X1 U5910 ( .A1(n8016), .A2(n8015), .ZN(n8133) );
  AND2_X1 U5911 ( .A1(n8556), .A2(n8564), .ZN(n4368) );
  AND2_X1 U5912 ( .A1(n4513), .A2(n6715), .ZN(n4369) );
  OR2_X1 U5913 ( .A1(n8767), .A2(n8584), .ZN(n8341) );
  AND2_X1 U5914 ( .A1(n8311), .A2(n8312), .ZN(n8641) );
  INV_X1 U5915 ( .A(n8641), .ZN(n4701) );
  INV_X1 U5916 ( .A(n9211), .ZN(n4554) );
  NOR2_X1 U5917 ( .A1(n7680), .A2(n8965), .ZN(n4370) );
  INV_X1 U5918 ( .A(n4830), .ZN(n4829) );
  NAND2_X1 U5919 ( .A1(n9158), .A2(n9136), .ZN(n4830) );
  NOR2_X1 U5920 ( .A1(n7832), .A2(n7831), .ZN(n4371) );
  AND3_X1 U5921 ( .A1(n4973), .A2(n4974), .A3(n4583), .ZN(n4372) );
  NAND2_X1 U5922 ( .A1(n8445), .A2(n8760), .ZN(n4373) );
  OR2_X1 U5923 ( .A1(n4481), .A2(n4475), .ZN(n4374) );
  INV_X1 U5924 ( .A(n6615), .ZN(n4551) );
  NOR2_X1 U5925 ( .A1(n4559), .A2(n7232), .ZN(n4375) );
  INV_X1 U5926 ( .A(n4851), .ZN(n4848) );
  NAND2_X1 U5927 ( .A1(n9964), .A2(n7611), .ZN(n4851) );
  AND2_X1 U5928 ( .A1(n4325), .A2(n5426), .ZN(n4376) );
  AND2_X1 U5929 ( .A1(n8008), .A2(n8632), .ZN(n4377) );
  AND2_X1 U5930 ( .A1(n7312), .A2(n7311), .ZN(n4378) );
  NAND2_X1 U5931 ( .A1(n5521), .A2(n4919), .ZN(n4379) );
  NAND2_X1 U5932 ( .A1(n4529), .A2(n4530), .ZN(n4380) );
  INV_X1 U5933 ( .A(n4579), .ZN(n4578) );
  NAND2_X1 U5934 ( .A1(n4581), .A2(n4580), .ZN(n4579) );
  INV_X1 U5935 ( .A(n4715), .ZN(n4714) );
  OR2_X1 U5936 ( .A1(n8898), .A2(n4716), .ZN(n4715) );
  INV_X1 U5937 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4920) );
  INV_X1 U5938 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5631) );
  AND2_X1 U5939 ( .A1(n4680), .A2(n5171), .ZN(n4381) );
  NAND2_X1 U5940 ( .A1(n5290), .A2(n5289), .ZN(n7992) );
  AND2_X1 U5941 ( .A1(n5110), .A2(n5109), .ZN(n4382) );
  AND2_X1 U5942 ( .A1(n4717), .A2(n6121), .ZN(n4383) );
  NAND2_X1 U5943 ( .A1(n8358), .A2(n5556), .ZN(n4384) );
  INV_X1 U5944 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8816) );
  NAND2_X1 U5945 ( .A1(n4861), .A2(n8006), .ZN(n8087) );
  OR2_X1 U5946 ( .A1(n8760), .A2(n8573), .ZN(n8345) );
  INV_X1 U5947 ( .A(n8345), .ZN(n4611) );
  AND2_X1 U5948 ( .A1(n4447), .A2(n8905), .ZN(n4385) );
  AND2_X1 U5949 ( .A1(n4482), .A2(n8440), .ZN(n4386) );
  AND2_X1 U5950 ( .A1(n7578), .A2(n4350), .ZN(n4387) );
  AND2_X1 U5951 ( .A1(n9181), .A2(n4832), .ZN(n4388) );
  AND2_X1 U5952 ( .A1(n7996), .A2(n8677), .ZN(n4389) );
  AND2_X1 U5953 ( .A1(n4573), .A2(n9258), .ZN(n4390) );
  NOR2_X1 U5954 ( .A1(n4540), .A2(n4545), .ZN(n4391) );
  NAND2_X1 U5955 ( .A1(n7790), .A2(n9108), .ZN(n9660) );
  INV_X1 U5956 ( .A(n9660), .ZN(n6580) );
  INV_X1 U5957 ( .A(n8767), .ZN(n8714) );
  NAND2_X1 U5958 ( .A1(n5441), .A2(n5440), .ZN(n8767) );
  AND2_X1 U5959 ( .A1(n4541), .A2(n6577), .ZN(n4392) );
  AND2_X1 U5960 ( .A1(n4341), .A2(n9161), .ZN(n4393) );
  INV_X1 U5961 ( .A(n4653), .ZN(n4652) );
  OAI21_X1 U5962 ( .B1(n4654), .B2(n9150), .A(n9153), .ZN(n4653) );
  AND2_X1 U5963 ( .A1(n7984), .A2(n7983), .ZN(n4394) );
  OR2_X1 U5964 ( .A1(n4685), .A2(n4918), .ZN(n4395) );
  AND2_X1 U5965 ( .A1(n4436), .A2(n6045), .ZN(n4396) );
  AND2_X1 U5966 ( .A1(n5826), .A2(n7447), .ZN(n4397) );
  INV_X1 U5967 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4498) );
  OR2_X1 U5968 ( .A1(n5135), .A2(SI_9_), .ZN(n4398) );
  INV_X1 U5969 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4454) );
  INV_X1 U5970 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5209) );
  INV_X1 U5971 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5159) );
  NAND2_X2 U5972 ( .A1(n8823), .A2(n8827), .ZN(n5380) );
  INV_X1 U5973 ( .A(n5011), .ZN(n5565) );
  NAND2_X1 U5974 ( .A1(n7658), .A2(n4597), .ZN(n4599) );
  NAND2_X1 U5975 ( .A1(n7753), .A2(n5914), .ZN(n7728) );
  NAND2_X1 U5976 ( .A1(n9818), .A2(n4578), .ZN(n4399) );
  INV_X1 U5977 ( .A(n8571), .ZN(n4689) );
  XNOR2_X1 U5978 ( .A(n6289), .B(n7812), .ZN(n7802) );
  NOR2_X1 U5979 ( .A1(n4302), .A2(n4726), .ZN(n5985) );
  INV_X1 U5980 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4523) );
  NAND2_X1 U5981 ( .A1(n4870), .A2(n4317), .ZN(n8171) );
  NAND2_X1 U5982 ( .A1(n5511), .A2(n5510), .ZN(n5618) );
  OR2_X1 U5983 ( .A1(n7232), .A2(n6704), .ZN(n6838) );
  AND2_X1 U5984 ( .A1(n6594), .A2(n6593), .ZN(n4400) );
  AND2_X1 U5985 ( .A1(n4870), .A2(n4869), .ZN(n8122) );
  NAND2_X1 U5986 ( .A1(n6105), .A2(n4894), .ZN(n8896) );
  NAND2_X1 U5987 ( .A1(n4456), .A2(n4455), .ZN(n8857) );
  OR2_X1 U5988 ( .A1(n9502), .A2(n6471), .ZN(n9473) );
  INV_X1 U5989 ( .A(n9473), .ZN(n4542) );
  NOR2_X1 U5990 ( .A1(n7801), .A2(n6290), .ZN(n4401) );
  NAND2_X1 U5991 ( .A1(n9449), .A2(n4575), .ZN(n4576) );
  AND2_X1 U5992 ( .A1(n8867), .A2(n6357), .ZN(n4402) );
  AND2_X1 U5993 ( .A1(n4794), .A2(n4793), .ZN(n4403) );
  AND2_X1 U5994 ( .A1(n4747), .A2(n4746), .ZN(n4404) );
  INV_X1 U5995 ( .A(n9134), .ZN(n4834) );
  AND2_X1 U5996 ( .A1(n9449), .A2(n4390), .ZN(n9236) );
  INV_X1 U5997 ( .A(n4780), .ZN(n4779) );
  NOR2_X1 U5998 ( .A1(n5300), .A2(SI_17_), .ZN(n4780) );
  INV_X1 U5999 ( .A(n4463), .ZN(n4462) );
  NAND2_X1 U6000 ( .A1(n6085), .A2(n6084), .ZN(n4463) );
  OAI21_X2 U6001 ( .B1(n6823), .B2(n5888), .A(n5940), .ZN(n6463) );
  INV_X1 U6002 ( .A(n6463), .ZN(n4850) );
  AND2_X1 U6003 ( .A1(n6208), .A2(n6202), .ZN(n8941) );
  AND2_X1 U6004 ( .A1(n6859), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4405) );
  NAND2_X1 U6005 ( .A1(n6049), .A2(n6048), .ZN(n9502) );
  INV_X1 U6006 ( .A(n9502), .ZN(n4580) );
  OR2_X1 U6007 ( .A1(n10008), .A2(n6425), .ZN(n4406) );
  NAND2_X1 U6008 ( .A1(n8439), .A2(n8383), .ZN(n8355) );
  OAI21_X1 U6009 ( .B1(n7635), .B2(n8259), .A(n8272), .ZN(n7577) );
  AND2_X1 U6010 ( .A1(n4876), .A2(n4877), .ZN(n4407) );
  NAND2_X1 U6011 ( .A1(n5133), .A2(n5132), .ZN(n4408) );
  NAND2_X1 U6012 ( .A1(n4808), .A2(n7292), .ZN(n7310) );
  NAND2_X1 U6013 ( .A1(n4815), .A2(n7481), .ZN(n7566) );
  AND2_X1 U6014 ( .A1(n4722), .A2(n5826), .ZN(n7446) );
  INV_X1 U6015 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4820) );
  NAND2_X1 U6016 ( .A1(n6107), .A2(n6106), .ZN(n9556) );
  INV_X1 U6017 ( .A(n9556), .ZN(n9092) );
  NAND2_X1 U6018 ( .A1(n6901), .A2(n5738), .ZN(n8840) );
  AND2_X1 U6019 ( .A1(n4796), .A2(n4799), .ZN(n4409) );
  OR2_X1 U6020 ( .A1(n9990), .A2(n9828), .ZN(n4410) );
  OR2_X1 U6021 ( .A1(n4405), .A2(n4632), .ZN(n4411) );
  AND2_X1 U6022 ( .A1(n4589), .A2(n5536), .ZN(n4412) );
  INV_X1 U6023 ( .A(n8459), .ZN(n4880) );
  NAND2_X1 U6024 ( .A1(n4338), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7182) );
  AND2_X1 U6025 ( .A1(n6644), .A2(n7587), .ZN(n4413) );
  INV_X1 U6026 ( .A(n4739), .ZN(n6914) );
  NAND2_X1 U6027 ( .A1(n6278), .A2(n6959), .ZN(n4739) );
  XOR2_X1 U6028 ( .A(n6972), .B(n7194), .Z(n4414) );
  XOR2_X1 U6029 ( .A(n6284), .B(P2_REG2_REG_8__SCAN_IN), .Z(n4415) );
  INV_X1 U6030 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n4741) );
  INV_X1 U6031 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n4584) );
  INV_X1 U6032 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n4424) );
  XNOR2_X1 U6033 ( .A(n6264), .B(n7869), .ZN(n7856) );
  XNOR2_X1 U6034 ( .A(n6300), .B(n7087), .ZN(n10024) );
  INV_X1 U6035 ( .A(n9892), .ZN(n9499) );
  NAND2_X1 U6036 ( .A1(n4962), .A2(n4963), .ZN(n4977) );
  NAND2_X1 U6037 ( .A1(n4981), .A2(n4980), .ZN(n4999) );
  NOR2_X2 U6038 ( .A1(n9225), .A2(n9157), .ZN(n9188) );
  INV_X1 U6039 ( .A(n6536), .ZN(n9109) );
  NAND2_X1 U6040 ( .A1(n4665), .A2(n4663), .ZN(n9664) );
  OAI21_X1 U6041 ( .B1(n4650), .B2(n4653), .A(n4649), .ZN(n9245) );
  NAND2_X1 U6042 ( .A1(n4773), .A2(n5354), .ZN(n5365) );
  NAND2_X1 U6043 ( .A1(n5128), .A2(n4898), .ZN(n7548) );
  NAND2_X1 U6044 ( .A1(n5091), .A2(n5107), .ZN(n5128) );
  NAND2_X2 U6045 ( .A1(n4416), .A2(n5081), .ZN(n10060) );
  NAND2_X1 U6046 ( .A1(n6757), .A2(n8209), .ZN(n4416) );
  NAND2_X1 U6047 ( .A1(n5102), .A2(n5080), .ZN(n5112) );
  NAND2_X1 U6048 ( .A1(n8570), .A2(n8571), .ZN(n4690) );
  NOR2_X1 U6049 ( .A1(n10024), .A2(n10025), .ZN(n10023) );
  NAND2_X1 U6050 ( .A1(n4417), .A2(n4740), .ZN(n6962) );
  NAND2_X1 U6051 ( .A1(n4738), .A2(n6959), .ZN(n4417) );
  NAND2_X1 U6052 ( .A1(n6281), .A2(n7099), .ZN(n7104) );
  NOR2_X1 U6053 ( .A1(n8522), .A2(n8521), .ZN(n8520) );
  XNOR2_X1 U6054 ( .A(n6303), .B(n6344), .ZN(n4737) );
  AOI22_X2 U6055 ( .A1(n9659), .A2(n9662), .B1(n9111), .B2(n9668), .ZN(n9495)
         );
  AOI21_X2 U6056 ( .B1(n9458), .B2(n9117), .A(n9116), .ZN(n9442) );
  AOI21_X2 U6057 ( .B1(n4818), .B2(n4817), .A(n4816), .ZN(n9234) );
  NAND2_X1 U6058 ( .A1(n4837), .A2(n4838), .ZN(n4836) );
  NOR2_X2 U6059 ( .A1(n4661), .A2(n9169), .ZN(n4659) );
  NOR2_X2 U6060 ( .A1(n4346), .A2(n9193), .ZN(n9195) );
  NOR2_X2 U6061 ( .A1(n9444), .A2(n9149), .ZN(n9284) );
  INV_X1 U6062 ( .A(n6466), .ZN(n4667) );
  NAND2_X1 U6063 ( .A1(n9810), .A2(n4666), .ZN(n4665) );
  OR2_X1 U6064 ( .A1(n8413), .A2(n8412), .ZN(n8414) );
  NAND2_X1 U6065 ( .A1(n9234), .A2(n9233), .ZN(n9232) );
  INV_X1 U6066 ( .A(n9253), .ZN(n4818) );
  OAI21_X1 U6067 ( .B1(n4844), .B2(n4846), .A(n7785), .ZN(n4843) );
  NOR2_X1 U6068 ( .A1(n9513), .A2(n9937), .ZN(n4661) );
  INV_X1 U6069 ( .A(n4801), .ZN(n4800) );
  NAND2_X1 U6070 ( .A1(n4622), .A2(n4621), .ZN(n4890) );
  INV_X1 U6071 ( .A(n8536), .ZN(n4802) );
  AOI21_X2 U6072 ( .B1(n6323), .B2(n6749), .A(n7058), .ZN(n7097) );
  INV_X1 U6073 ( .A(n5099), .ZN(n4754) );
  OAI21_X1 U6074 ( .B1(n4753), .B2(n4752), .A(n4398), .ZN(n4750) );
  OAI21_X1 U6075 ( .B1(n8592), .B2(n8377), .A(n8375), .ZN(n8580) );
  NAND2_X1 U6076 ( .A1(n4778), .A2(n4779), .ZN(n5305) );
  NAND3_X1 U6077 ( .A1(n4430), .A2(n4431), .A3(n5780), .ZN(n5799) );
  NAND2_X1 U6078 ( .A1(n8841), .A2(n4435), .ZN(n4434) );
  OAI21_X1 U6079 ( .B1(n6901), .B2(n4432), .A(n4433), .ZN(n7026) );
  NAND3_X1 U6080 ( .A1(n4434), .A2(n5776), .A3(n4432), .ZN(n4431) );
  INV_X1 U6081 ( .A(n8841), .ZN(n4432) );
  NAND2_X1 U6082 ( .A1(n8840), .A2(n8841), .ZN(n7024) );
  NAND2_X1 U6083 ( .A1(n4719), .A2(n4437), .ZN(n4436) );
  NAND3_X1 U6084 ( .A1(n4440), .A2(n8939), .A3(n6023), .ZN(n8938) );
  NAND3_X1 U6085 ( .A1(n4440), .A2(n4438), .A3(n6023), .ZN(n4441) );
  NAND2_X1 U6086 ( .A1(n4441), .A2(n4396), .ZN(n8885) );
  INV_X1 U6087 ( .A(n4719), .ZN(n4442) );
  INV_X1 U6088 ( .A(n5647), .ZN(n4444) );
  NOR2_X2 U6089 ( .A1(n9896), .A2(n4444), .ZN(n9892) );
  NAND2_X1 U6090 ( .A1(n8904), .A2(n4385), .ZN(n4445) );
  NAND2_X1 U6091 ( .A1(n4445), .A2(n4446), .ZN(n6181) );
  NAND3_X1 U6092 ( .A1(n4445), .A2(n4446), .A3(n6158), .ZN(n4519) );
  NAND2_X1 U6093 ( .A1(n5639), .A2(n4452), .ZN(n4450) );
  NAND2_X1 U6094 ( .A1(n8916), .A2(n4457), .ZN(n4456) );
  AND2_X1 U6095 ( .A1(n5037), .A2(n4466), .ZN(n5145) );
  NAND4_X1 U6096 ( .A1(n4472), .A2(n4471), .A3(n8290), .A4(n5540), .ZN(n4469)
         );
  NAND2_X1 U6097 ( .A1(n8279), .A2(n4275), .ZN(n4471) );
  NAND2_X1 U6098 ( .A1(n8280), .A2(n8355), .ZN(n4472) );
  OAI211_X1 U6099 ( .C1(n8415), .C2(n4474), .A(n4473), .B(n4477), .ZN(n4476)
         );
  NAND2_X1 U6100 ( .A1(n4478), .A2(n4386), .ZN(n4474) );
  INV_X1 U6101 ( .A(n4476), .ZN(P2_U3296) );
  NAND2_X1 U6102 ( .A1(n8440), .A2(n8441), .ZN(n4477) );
  NAND3_X1 U6103 ( .A1(n8296), .A2(n8297), .A3(n4275), .ZN(n4490) );
  NOR2_X1 U6104 ( .A1(n8384), .A2(n4491), .ZN(n4492) );
  NAND2_X1 U6105 ( .A1(n8236), .A2(n4492), .ZN(n4494) );
  NAND3_X1 U6106 ( .A1(n4494), .A2(n8247), .A3(n4493), .ZN(n8250) );
  NAND2_X1 U6107 ( .A1(n8236), .A2(n8235), .ZN(n8246) );
  NOR2_X1 U6108 ( .A1(n4501), .A2(n4500), .ZN(n4499) );
  NOR2_X1 U6109 ( .A1(n6242), .A2(n6922), .ZN(n4500) );
  NAND2_X2 U6110 ( .A1(n6242), .A2(n6735), .ZN(n4997) );
  NAND2_X2 U6111 ( .A1(n6242), .A2(n6736), .ZN(n5039) );
  NAND2_X4 U6112 ( .A1(n5562), .A2(n5561), .ZN(n6242) );
  NAND2_X1 U6113 ( .A1(n4355), .A2(n4511), .ZN(n4508) );
  NAND2_X1 U6114 ( .A1(n8348), .A2(n4354), .ZN(n4507) );
  NAND2_X1 U6115 ( .A1(n4505), .A2(n4502), .ZN(n8360) );
  INV_X1 U6116 ( .A(n4503), .ZN(n4502) );
  OAI21_X1 U6117 ( .B1(n8359), .B2(n4510), .A(n4504), .ZN(n4503) );
  INV_X1 U6118 ( .A(n8359), .ZN(n4506) );
  OR2_X1 U6119 ( .A1(n6181), .A2(n4515), .ZN(n4512) );
  NAND2_X1 U6120 ( .A1(n6181), .A2(n4516), .ZN(n4514) );
  NAND2_X1 U6121 ( .A1(n4998), .A2(n4520), .ZN(n4982) );
  NAND2_X1 U6122 ( .A1(n4521), .A2(SI_2_), .ZN(n4998) );
  NAND2_X1 U6123 ( .A1(n5000), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4522) );
  NAND2_X1 U6124 ( .A1(n4528), .A2(n5075), .ZN(n4529) );
  NAND2_X1 U6125 ( .A1(n5075), .A2(n5074), .ZN(n5100) );
  NAND2_X1 U6126 ( .A1(n7271), .A2(n4531), .ZN(n6529) );
  OAI21_X1 U6127 ( .B1(n7517), .B2(n4531), .A(n7516), .ZN(n7518) );
  NAND2_X1 U6128 ( .A1(n7517), .A2(n4531), .ZN(n7516) );
  XNOR2_X1 U6129 ( .A(n7515), .B(n4532), .ZN(n9905) );
  NAND2_X1 U6130 ( .A1(n4537), .A2(n4535), .ZN(n6602) );
  NAND2_X1 U6131 ( .A1(n6578), .A2(n4544), .ZN(n4539) );
  NAND2_X1 U6132 ( .A1(n4539), .A2(n4543), .ZN(n6595) );
  AND2_X1 U6133 ( .A1(n4547), .A2(n4548), .ZN(n6619) );
  NAND3_X1 U6134 ( .A1(n6612), .A2(n6617), .A3(n4552), .ZN(n4547) );
  AOI21_X1 U6135 ( .B1(n6612), .B2(n6611), .A(n4555), .ZN(n6620) );
  NAND2_X1 U6136 ( .A1(n4556), .A2(n4557), .ZN(n6639) );
  NAND3_X1 U6137 ( .A1(n6636), .A2(n6635), .A3(n4558), .ZN(n4556) );
  AND3_X1 U6138 ( .A1(n6636), .A2(n6700), .A3(n6635), .ZN(n6701) );
  NAND2_X1 U6139 ( .A1(n9176), .A2(n4566), .ZN(n4567) );
  INV_X1 U6140 ( .A(n4567), .ZN(n9142) );
  NAND2_X1 U6141 ( .A1(n9176), .A2(n4565), .ZN(n4564) );
  NAND3_X1 U6142 ( .A1(n4571), .A2(n6556), .A3(n4570), .ZN(n4569) );
  NAND4_X1 U6143 ( .A1(n6549), .A2(n7473), .A3(n7318), .A4(n6703), .ZN(n4570)
         );
  INV_X1 U6144 ( .A(n4576), .ZN(n9288) );
  NAND2_X1 U6145 ( .A1(n4372), .A2(n4972), .ZN(n8462) );
  OR2_X1 U6146 ( .A1(n5380), .A2(n4584), .ZN(n4583) );
  OAI21_X1 U6147 ( .B1(n5538), .B2(n5537), .A(n4588), .ZN(n4586) );
  NAND2_X1 U6148 ( .A1(n7658), .A2(n4591), .ZN(n4590) );
  NAND2_X1 U6149 ( .A1(n5549), .A2(n4326), .ZN(n4600) );
  NAND2_X1 U6150 ( .A1(n4600), .A2(n4601), .ZN(n8613) );
  INV_X1 U6151 ( .A(n8569), .ZN(n4607) );
  NOR2_X1 U6152 ( .A1(n5523), .A2(n4617), .ZN(n4945) );
  INV_X1 U6153 ( .A(n5523), .ZN(n4622) );
  NAND2_X1 U6154 ( .A1(n6913), .A2(n4627), .ZN(n4626) );
  NAND2_X1 U6155 ( .A1(n6913), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6912) );
  AND2_X1 U6156 ( .A1(n4628), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4627) );
  NOR2_X1 U6157 ( .A1(n8465), .A2(n4405), .ZN(n6266) );
  NAND3_X1 U6158 ( .A1(n4630), .A2(n4631), .A3(n4629), .ZN(n8493) );
  NAND3_X1 U6159 ( .A1(n4630), .A2(n4337), .A3(n4629), .ZN(n4633) );
  INV_X1 U6160 ( .A(n4633), .ZN(n8492) );
  NAND2_X1 U6161 ( .A1(n4798), .A2(n4336), .ZN(n4634) );
  NAND2_X1 U6162 ( .A1(n4635), .A2(n4634), .ZN(n7704) );
  INV_X1 U6163 ( .A(n6952), .ZN(n6317) );
  NOR2_X1 U6164 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(n6244), .ZN(n4637) );
  NOR2_X1 U6165 ( .A1(n10019), .A2(n10018), .ZN(n10017) );
  NAND2_X1 U6166 ( .A1(n6270), .A2(n4640), .ZN(n4638) );
  INV_X1 U6167 ( .A(n8524), .ZN(n4640) );
  OR2_X1 U6168 ( .A1(n4311), .A2(n6740), .ZN(n5691) );
  XNOR2_X2 U6169 ( .A(n5634), .B(n4285), .ZN(n6707) );
  NAND2_X1 U6170 ( .A1(n4641), .A2(n4642), .ZN(n9164) );
  NAND2_X1 U6171 ( .A1(n9188), .A2(n4393), .ZN(n4641) );
  NAND2_X1 U6172 ( .A1(n9188), .A2(n4341), .ZN(n4645) );
  INV_X1 U6173 ( .A(n9284), .ZN(n4650) );
  NAND2_X1 U6174 ( .A1(n4662), .A2(n9170), .ZN(n9512) );
  OAI21_X1 U6175 ( .B1(n6468), .B2(n6580), .A(n6583), .ZN(n4664) );
  NOR2_X1 U6176 ( .A1(n4667), .A2(n6580), .ZN(n4666) );
  OAI21_X1 U6177 ( .B1(n7486), .B2(n4670), .A(n4668), .ZN(n7683) );
  NAND3_X1 U6178 ( .A1(n7689), .A2(n4671), .A3(n4672), .ZN(n4669) );
  NOR2_X1 U6179 ( .A1(n7309), .A2(n4678), .ZN(n4677) );
  NAND2_X1 U6180 ( .A1(n9244), .A2(n9155), .ZN(n9225) );
  OAI211_X1 U6181 ( .C1(n8425), .C2(n8424), .A(n8423), .B(n8422), .ZN(n8427)
         );
  NOR2_X1 U6182 ( .A1(n10098), .A2(n7800), .ZN(n7799) );
  NOR2_X1 U6183 ( .A1(n6251), .A2(n6250), .ZN(n6913) );
  AOI21_X1 U6184 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7247), .A(n7239), .ZN(
        n6258) );
  AOI21_X1 U6185 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n6824), .A(n7877), .ZN(
        n6264) );
  NOR2_X1 U6186 ( .A1(n6263), .A2(n7799), .ZN(n7879) );
  NAND2_X1 U6187 ( .A1(n6265), .A2(n4795), .ZN(n4791) );
  INV_X1 U6188 ( .A(n8381), .ZN(n8224) );
  NAND2_X1 U6189 ( .A1(n6983), .A2(n6985), .ZN(n8222) );
  NOR2_X1 U6190 ( .A1(n9446), .A2(n9445), .ZN(n9444) );
  XNOR2_X1 U6191 ( .A(n5669), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5673) );
  OAI211_X1 U6192 ( .C1(n6356), .C2(n10020), .A(n6355), .B(n4736), .ZN(
        P2_U3201) );
  OAI21_X2 U6193 ( .B1(n4682), .B2(n4683), .A(n4381), .ZN(n7659) );
  NAND2_X1 U6194 ( .A1(n5133), .A2(n4350), .ZN(n4679) );
  INV_X1 U6195 ( .A(n4352), .ZN(n4681) );
  NAND2_X1 U6196 ( .A1(n5133), .A2(n4387), .ZN(n4682) );
  NAND4_X1 U6197 ( .A1(n4686), .A2(n4917), .A3(n5209), .A4(n5273), .ZN(n4685)
         );
  OAI21_X1 U6198 ( .B1(n8581), .B2(n8582), .A(n5426), .ZN(n8570) );
  INV_X1 U6199 ( .A(n5887), .ZN(n7753) );
  NAND3_X1 U6200 ( .A1(n4710), .A2(n4711), .A3(n5979), .ZN(n6004) );
  NAND2_X1 U6201 ( .A1(n5887), .A2(n4327), .ZN(n4710) );
  NAND2_X1 U6202 ( .A1(n8885), .A2(n8886), .ZN(n8884) );
  INV_X1 U6203 ( .A(n6022), .ZN(n4718) );
  NAND2_X1 U6204 ( .A1(n7817), .A2(n7816), .ZN(n4719) );
  NOR2_X1 U6205 ( .A1(n6137), .A2(n6136), .ZN(n6138) );
  INV_X1 U6206 ( .A(n6136), .ZN(n4720) );
  NAND2_X1 U6207 ( .A1(n4722), .A2(n4397), .ZN(n5846) );
  NAND2_X1 U6208 ( .A1(n5800), .A2(n4721), .ZN(n4722) );
  NAND2_X1 U6209 ( .A1(n5800), .A2(n7165), .ZN(n7254) );
  INV_X1 U6210 ( .A(n4722), .ZN(n7255) );
  INV_X1 U6211 ( .A(n7256), .ZN(n4723) );
  NAND2_X1 U6212 ( .A1(n7026), .A2(n4724), .ZN(n7164) );
  NAND4_X1 U6213 ( .A1(n5623), .A2(n5624), .A3(n5625), .A4(n5626), .ZN(n4726)
         );
  NAND3_X1 U6214 ( .A1(n6644), .A2(n6731), .A3(n7471), .ZN(n5688) );
  NAND2_X1 U6215 ( .A1(n6046), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4727) );
  NOR2_X1 U6216 ( .A1(n8482), .A2(n6297), .ZN(n8503) );
  NAND2_X1 U6217 ( .A1(n6280), .A2(n6749), .ZN(n7100) );
  NAND2_X1 U6218 ( .A1(n4731), .A2(n7063), .ZN(n4730) );
  INV_X1 U6219 ( .A(n6280), .ZN(n4731) );
  INV_X1 U6220 ( .A(n4910), .ZN(n4732) );
  NAND2_X1 U6221 ( .A1(n4732), .A2(n7243), .ZN(n4734) );
  NAND2_X1 U6222 ( .A1(n4734), .A2(n4733), .ZN(n7245) );
  INV_X1 U6223 ( .A(n6278), .ZN(n4738) );
  XNOR2_X1 U6224 ( .A(n6293), .B(n7869), .ZN(n7865) );
  OAI21_X1 U6225 ( .B1(n4745), .B2(n7865), .A(n4744), .ZN(n8474) );
  NAND3_X1 U6226 ( .A1(n4749), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4937) );
  NAND2_X1 U6227 ( .A1(n5470), .A2(n4762), .ZN(n4760) );
  NAND2_X1 U6228 ( .A1(n4773), .A2(n4772), .ZN(n5371) );
  NAND2_X1 U6229 ( .A1(n5287), .A2(n4781), .ZN(n4778) );
  NAND2_X1 U6230 ( .A1(n8210), .A2(n8209), .ZN(n4784) );
  NAND2_X1 U6231 ( .A1(n4784), .A2(n8211), .ZN(n8754) );
  INV_X1 U6232 ( .A(n4786), .ZN(n8512) );
  NAND3_X1 U6233 ( .A1(n4975), .A2(n4789), .A3(n4787), .ZN(n7049) );
  NAND2_X1 U6234 ( .A1(n6258), .A2(n7348), .ZN(n4798) );
  NAND2_X1 U6235 ( .A1(n4803), .A2(n4800), .ZN(P2_U3200) );
  OAI21_X1 U6236 ( .B1(n8523), .B2(n4333), .A(n7180), .ZN(n4803) );
  NAND3_X1 U6237 ( .A1(n5760), .A2(n5725), .A3(n4804), .ZN(n5801) );
  NAND3_X1 U6238 ( .A1(n9867), .A2(n9868), .A3(n7309), .ZN(n4806) );
  NAND2_X1 U6239 ( .A1(n9867), .A2(n9868), .ZN(n4808) );
  NAND2_X1 U6240 ( .A1(n4806), .A2(n4805), .ZN(n9851) );
  NAND2_X1 U6241 ( .A1(n9824), .A2(n4810), .ZN(n4809) );
  NAND2_X1 U6242 ( .A1(n9219), .A2(n9135), .ZN(n4835) );
  NAND2_X1 U6243 ( .A1(n9219), .A2(n4822), .ZN(n4821) );
  NAND2_X1 U6244 ( .A1(n4836), .A2(n4334), .ZN(n4844) );
  NOR2_X1 U6245 ( .A1(n7689), .A2(n4847), .ZN(n4846) );
  OAI21_X2 U6246 ( .B1(n4840), .B2(n7613), .A(n4839), .ZN(n9806) );
  OR2_X1 U6247 ( .A1(n4844), .A2(n4841), .ZN(n4840) );
  NAND2_X1 U6248 ( .A1(n5037), .A2(n4852), .ZN(n5158) );
  OAI21_X2 U6249 ( .B1(n7597), .B2(n4855), .A(n4853), .ZN(n7901) );
  INV_X1 U6250 ( .A(n4856), .ZN(n4855) );
  NAND2_X1 U6251 ( .A1(n8111), .A2(n4317), .ZN(n4865) );
  NAND2_X1 U6252 ( .A1(n4865), .A2(n4866), .ZN(n7999) );
  INV_X1 U6253 ( .A(n7366), .ZN(n4882) );
  NAND2_X1 U6254 ( .A1(n7065), .A2(n4883), .ZN(n7067) );
  NOR2_X1 U6255 ( .A1(n4879), .A2(n7068), .ZN(n4878) );
  INV_X1 U6256 ( .A(n4883), .ZN(n4879) );
  NAND2_X1 U6257 ( .A1(n4884), .A2(n8461), .ZN(n4883) );
  INV_X1 U6258 ( .A(n7066), .ZN(n4884) );
  NAND2_X1 U6259 ( .A1(n8095), .A2(n4394), .ZN(n8151) );
  NOR2_X2 U6260 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4954) );
  NAND2_X1 U6261 ( .A1(n4890), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4944) );
  AND2_X1 U6262 ( .A1(n6249), .A2(n6248), .ZN(n6250) );
  NAND2_X2 U6263 ( .A1(n7940), .A2(n5299), .ZN(n8652) );
  XNOR2_X1 U6264 ( .A(n6493), .B(n6492), .ZN(n6491) );
  INV_X1 U6265 ( .A(n5673), .ZN(n7920) );
  OAI21_X1 U6266 ( .B1(n6516), .B2(n6515), .A(n6514), .ZN(n6519) );
  NAND2_X2 U6267 ( .A1(n5527), .A2(n8222), .ZN(n8380) );
  OAI21_X1 U6268 ( .B1(n8380), .B2(n8217), .A(n5527), .ZN(n7144) );
  INV_X1 U6269 ( .A(n5005), .ZN(n5002) );
  XNOR2_X1 U6270 ( .A(n5505), .B(n5504), .ZN(n7874) );
  AOI22_X2 U6271 ( .A1(n8594), .A2(n5403), .B1(n8585), .B2(n8721), .ZN(n8581)
         );
  XNOR2_X1 U6272 ( .A(n5453), .B(n5452), .ZN(n7725) );
  NAND2_X1 U6273 ( .A1(n8074), .A2(n8585), .ZN(n8073) );
  NAND2_X1 U6274 ( .A1(n8180), .A2(n8024), .ZN(n8187) );
  XNOR2_X1 U6275 ( .A(n6491), .B(SI_29_), .ZN(n6446) );
  NAND2_X1 U6276 ( .A1(n8104), .A2(n8105), .ZN(n8180) );
  AND2_X1 U6277 ( .A1(n6988), .A2(n4987), .ZN(n6989) );
  OAI21_X1 U6278 ( .B1(n5000), .B2(n6741), .A(n4961), .ZN(n4963) );
  NAND2_X1 U6279 ( .A1(n5000), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4961) );
  NAND2_X1 U6280 ( .A1(n5000), .A2(n5707), .ZN(n4958) );
  AOI21_X2 U6281 ( .B1(n7659), .B2(n5191), .A(n5190), .ZN(n7743) );
  NAND2_X1 U6282 ( .A1(n5698), .A2(n5697), .ZN(n6897) );
  AOI22_X1 U6283 ( .A1(n9110), .A2(n9109), .B1(n9689), .B2(n9108), .ZN(n9659)
         );
  NOR2_X1 U6284 ( .A1(n5530), .A2(n7136), .ZN(n4891) );
  AND2_X1 U6285 ( .A1(n4896), .A2(n6239), .ZN(n4892) );
  NOR2_X1 U6286 ( .A1(n7994), .A2(n8120), .ZN(n4893) );
  NOR2_X1 U6287 ( .A1(n8556), .A2(n8444), .ZN(n4895) );
  OR2_X1 U6288 ( .A1(n8546), .A2(n8727), .ZN(n4896) );
  OR2_X1 U6289 ( .A1(n8431), .A2(n8430), .ZN(n4897) );
  NAND2_X1 U6290 ( .A1(n7626), .A2(n5107), .ZN(n4898) );
  NAND2_X1 U6291 ( .A1(n9511), .A2(n4351), .ZN(n4899) );
  AND2_X1 U6292 ( .A1(n9485), .A2(n9113), .ZN(n4902) );
  NOR2_X1 U6293 ( .A1(n8113), .A2(n7994), .ZN(n4903) );
  AND2_X1 U6294 ( .A1(n7154), .A2(n7160), .ZN(n4904) );
  AND2_X1 U6295 ( .A1(n7369), .A2(n8458), .ZN(n4905) );
  INV_X1 U6296 ( .A(n8433), .ZN(n5559) );
  XOR2_X1 U6297 ( .A(n8780), .B(n8037), .Z(n4906) );
  AND2_X1 U6298 ( .A1(n5450), .A2(n5449), .ZN(n8584) );
  INV_X1 U6299 ( .A(n8584), .ZN(n5451) );
  INV_X1 U6300 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5325) );
  INV_X1 U6301 ( .A(n8955), .ZN(n9168) );
  NOR2_X1 U6302 ( .A1(n8546), .A2(n8791), .ZN(n5619) );
  OR2_X1 U6303 ( .A1(n7306), .A2(n7307), .ZN(n10006) );
  INV_X1 U6304 ( .A(n10006), .ZN(n10008) );
  AND4_X1 U6305 ( .A1(n5297), .A2(n5296), .A3(n5295), .A4(n5294), .ZN(n8677)
         );
  INV_X1 U6306 ( .A(n8677), .ZN(n5298) );
  AND4_X1 U6307 ( .A1(n5283), .A2(n5282), .A3(n5281), .A4(n5280), .ZN(n8694)
         );
  INV_X1 U6308 ( .A(n8807), .ZN(n8115) );
  NAND2_X1 U6309 ( .A1(n7770), .A2(n7769), .ZN(n4908) );
  AND2_X1 U6310 ( .A1(n6698), .A2(n6697), .ZN(n4909) );
  INV_X1 U6311 ( .A(n9515), .ZN(n9093) );
  OR2_X1 U6312 ( .A1(n6283), .A2(n7178), .ZN(n4910) );
  OR2_X1 U6313 ( .A1(n8026), .A2(n8564), .ZN(n4911) );
  AND2_X2 U6314 ( .A1(n6925), .A2(n6238), .ZN(n10103) );
  AND2_X1 U6315 ( .A1(n5617), .A2(n5616), .ZN(n10087) );
  INV_X1 U6316 ( .A(n6607), .ZN(n6608) );
  AND2_X1 U6317 ( .A1(n9246), .A2(n6610), .ZN(n6611) );
  AND2_X1 U6318 ( .A1(n7460), .A2(n5127), .ZN(n5126) );
  INV_X1 U6319 ( .A(n5332), .ZN(n5331) );
  INV_X1 U6320 ( .A(n8694), .ZN(n5284) );
  NAND2_X1 U6321 ( .A1(n5008), .A2(n5007), .ZN(n7135) );
  INV_X1 U6322 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5622) );
  INV_X1 U6323 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5117) );
  NOR2_X1 U6324 ( .A1(n8530), .A2(n8660), .ZN(n6302) );
  NAND2_X1 U6325 ( .A1(n5331), .A2(n5330), .ZN(n5345) );
  AOI21_X1 U6326 ( .B1(n7966), .B2(n4911), .A(n4895), .ZN(n5488) );
  INV_X1 U6327 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4913) );
  OR2_X1 U6328 ( .A1(n5953), .A2(n5952), .ZN(n5954) );
  INV_X1 U6329 ( .A(n5688), .ZN(n6100) );
  INV_X1 U6330 ( .A(n6694), .ZN(n6695) );
  AND2_X1 U6331 ( .A1(n9246), .A2(n4340), .ZN(n9154) );
  NOR2_X1 U6332 ( .A1(n5961), .A2(n5960), .ZN(n5990) );
  INV_X1 U6333 ( .A(n7587), .ZN(n6704) );
  OR2_X1 U6334 ( .A1(n5405), .A2(n5409), .ZN(n5428) );
  NOR2_X1 U6335 ( .A1(n8012), .A2(n4361), .ZN(n8013) );
  INV_X1 U6336 ( .A(n5184), .ZN(n5183) );
  INV_X1 U6337 ( .A(n5419), .ZN(n5418) );
  INV_X1 U6338 ( .A(n7578), .ZN(n8396) );
  INV_X1 U6339 ( .A(n5251), .ZN(n5250) );
  INV_X1 U6340 ( .A(n6260), .ZN(n6261) );
  INV_X1 U6341 ( .A(n10060), .ZN(n5089) );
  OR2_X1 U6342 ( .A1(n5592), .A2(n5603), .ZN(n6229) );
  AOI21_X1 U6343 ( .B1(n8689), .B2(n8399), .A(n5257), .ZN(n8673) );
  OR2_X1 U6344 ( .A1(n5583), .A2(n5575), .ZN(n5576) );
  INV_X1 U6345 ( .A(n8866), .ZN(n8867) );
  NAND2_X1 U6346 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n6143), .ZN(n6164) );
  AND2_X1 U6347 ( .A1(n9561), .A2(n9115), .ZN(n9116) );
  OR2_X1 U6348 ( .A1(n6090), .A2(n8852), .ZN(n6108) );
  OR2_X1 U6349 ( .A1(n5942), .A2(n6881), .ZN(n5961) );
  NAND2_X1 U6350 ( .A1(n6755), .A2(n6736), .ZN(n5726) );
  NAND2_X1 U6351 ( .A1(n9092), .A2(n6475), .ZN(n9119) );
  NAND2_X1 U6352 ( .A1(n6644), .A2(n6837), .ZN(n6840) );
  OR2_X1 U6353 ( .A1(n5432), .A2(n5431), .ZN(n5433) );
  AND2_X1 U6354 ( .A1(n5895), .A2(n5894), .ZN(n5937) );
  NAND2_X1 U6355 ( .A1(n5076), .A2(SI_7_), .ZN(n5080) );
  OR2_X1 U6356 ( .A1(n7534), .A2(n8457), .ZN(n7535) );
  NAND2_X1 U6357 ( .A1(n5418), .A2(n8138), .ZN(n5444) );
  INV_X1 U6358 ( .A(n7594), .ZN(n7595) );
  NAND2_X1 U6359 ( .A1(n10019), .A2(n10018), .ZN(n10021) );
  AOI21_X1 U6360 ( .B1(n6354), .B2(n10031), .A(n6353), .ZN(n6355) );
  INV_X1 U6361 ( .A(n8284), .ZN(n5540) );
  NAND2_X1 U6362 ( .A1(n8341), .A2(n8342), .ZN(n8571) );
  INV_X1 U6363 ( .A(n8655), .ZN(n8693) );
  INV_X1 U6364 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7450) );
  NAND2_X1 U6365 ( .A1(n6004), .A2(n6003), .ZN(n7816) );
  INV_X1 U6366 ( .A(n5975), .ZN(n7766) );
  INV_X1 U6367 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7168) );
  INV_X1 U6368 ( .A(n9099), .ZN(n9094) );
  INV_X1 U6369 ( .A(n9176), .ZN(n9196) );
  NOR2_X1 U6370 ( .A1(n9530), .A2(n9132), .ZN(n9134) );
  INV_X1 U6371 ( .A(n9236), .ZN(n9254) );
  INV_X1 U6372 ( .A(n9449), .ZN(n9459) );
  AND2_X1 U6373 ( .A1(n6752), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6729) );
  INV_X1 U6374 ( .A(n7684), .ZN(n7785) );
  INV_X1 U6375 ( .A(n7271), .ZN(n9886) );
  INV_X1 U6376 ( .A(n5143), .ZN(n5142) );
  INV_X1 U6377 ( .A(n5024), .ZN(n5021) );
  AOI211_X1 U6378 ( .C1(n8444), .C2(n8039), .A(n8195), .B(n8047), .ZN(n8040)
         );
  NAND2_X1 U6379 ( .A1(n7017), .A2(n8698), .ZN(n8176) );
  AND2_X1 U6380 ( .A1(n5425), .A2(n5424), .ZN(n8596) );
  INV_X1 U6381 ( .A(n10010), .ZN(n7807) );
  NOR2_X1 U6382 ( .A1(n7342), .A2(n9303), .ZN(n7341) );
  INV_X1 U6383 ( .A(n10012), .ZN(n8528) );
  XNOR2_X1 U6384 ( .A(n8425), .B(n8356), .ZN(n5573) );
  INV_X1 U6385 ( .A(n8701), .ZN(n8699) );
  AND2_X1 U6386 ( .A1(n7007), .A2(n10079), .ZN(n6928) );
  INV_X1 U6387 ( .A(n8727), .ZN(n8744) );
  AND2_X1 U6388 ( .A1(n8539), .A2(n8538), .ZN(n8751) );
  INV_X1 U6389 ( .A(n10079), .ZN(n10066) );
  AND2_X1 U6390 ( .A1(n5225), .A2(n5245), .ZN(n8479) );
  OAI21_X1 U6391 ( .B1(n9200), .B2(n8951), .A(n6725), .ZN(n6726) );
  OAI211_X1 U6392 ( .C1(n6731), .C2(n6762), .A(n5710), .B(n5709), .ZN(n6852)
         );
  OR2_X1 U6393 ( .A1(n6412), .A2(n6720), .ZN(n6389) );
  AND2_X1 U6394 ( .A1(n6809), .A2(n6707), .ZN(n9763) );
  XNOR2_X1 U6395 ( .A(n9102), .B(n9094), .ZN(n9095) );
  OR2_X1 U6396 ( .A1(n7332), .A2(n6837), .ZN(n9481) );
  INV_X1 U6397 ( .A(n7309), .ZN(n7293) );
  INV_X1 U6398 ( .A(n9488), .ZN(n9893) );
  OR2_X1 U6399 ( .A1(n7332), .A2(n6708), .ZN(n9983) );
  INV_X1 U6400 ( .A(n9937), .ZN(n9979) );
  NAND2_X1 U6401 ( .A1(n6187), .A2(n6188), .ZN(n7264) );
  AND2_X1 U6402 ( .A1(n5850), .A2(n5864), .ZN(n6806) );
  INV_X1 U6403 ( .A(n7118), .ZN(n7915) );
  INV_X1 U6404 ( .A(n8200), .ZN(n8191) );
  AND2_X1 U6405 ( .A1(n6995), .A2(n6994), .ZN(n8195) );
  INV_X1 U6406 ( .A(n8418), .ZN(n8539) );
  INV_X1 U6407 ( .A(n8596), .ZN(n8446) );
  INV_X1 U6408 ( .A(n8099), .ZN(n8452) );
  INV_X1 U6409 ( .A(n8701), .ZN(n8682) );
  INV_X1 U6410 ( .A(n5573), .ZN(n8552) );
  NAND2_X1 U6411 ( .A1(n8699), .A2(n7191), .ZN(n8705) );
  AND2_X1 U6412 ( .A1(n6929), .A2(n8698), .ZN(n8701) );
  INV_X1 U6413 ( .A(n10103), .ZN(n10100) );
  XOR2_X1 U6414 ( .A(n8408), .B(n7951), .Z(n7965) );
  OR2_X1 U6415 ( .A1(n10087), .A2(n10081), .ZN(n8814) );
  INV_X2 U6416 ( .A(n10087), .ZN(n10085) );
  AND2_X1 U6417 ( .A1(n8437), .A2(n5592), .ZN(n6825) );
  INV_X1 U6418 ( .A(n6825), .ZN(n7919) );
  INV_X1 U6419 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6768) );
  NAND2_X1 U6420 ( .A1(n6225), .A2(n6224), .ZN(n6226) );
  INV_X1 U6421 ( .A(n7696), .ZN(n9977) );
  INV_X1 U6422 ( .A(n8941), .ZN(n8923) );
  OR2_X1 U6423 ( .A1(n6761), .A2(n6756), .ZN(n9805) );
  OR3_X1 U6424 ( .A1(n7266), .A2(n7232), .A3(n9481), .ZN(n9879) );
  AND2_X1 U6425 ( .A1(n7270), .A2(n9879), .ZN(n9881) );
  OR2_X1 U6426 ( .A1(n9881), .A2(n9670), .ZN(n9488) );
  INV_X1 U6427 ( .A(n10006), .ZN(n9569) );
  INV_X1 U6428 ( .A(n9991), .ZN(n9990) );
  AND2_X2 U6429 ( .A1(n7308), .A2(n7307), .ZN(n9991) );
  INV_X1 U6430 ( .A(n6185), .ZN(n7724) );
  OR2_X1 U6431 ( .A1(n6227), .A2(n6226), .ZN(P1_U3229) );
  NAND4_X1 U6432 ( .A1(n5269), .A2(n5267), .A3(n5159), .A4(n5325), .ZN(n4918)
         );
  NAND2_X1 U6433 ( .A1(n5575), .A2(n5578), .ZN(n5581) );
  INV_X1 U6434 ( .A(n5581), .ZN(n4922) );
  NOR2_X1 U6435 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4921) );
  NAND3_X1 U6436 ( .A1(n4922), .A2(n4921), .A3(n5608), .ZN(n4923) );
  NAND2_X1 U6437 ( .A1(n4971), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4933) );
  NAND2_X1 U6438 ( .A1(n5084), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n4932) );
  INV_X1 U6439 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n4928) );
  AND2_X2 U6440 ( .A1(n4929), .A2(n8827), .ZN(n5011) );
  NAND2_X1 U6441 ( .A1(n5011), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4930) );
  INV_X1 U6442 ( .A(n7924), .ZN(n8464) );
  INV_X1 U6443 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4936) );
  NAND3_X1 U6444 ( .A1(n4936), .A2(n4935), .A3(n4934), .ZN(n4938) );
  INV_X2 U6445 ( .A(n5000), .ZN(n6736) );
  NAND2_X1 U6446 ( .A1(n6736), .A2(SI_0_), .ZN(n4939) );
  XNOR2_X1 U6447 ( .A(n4939), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8828) );
  NAND2_X1 U6448 ( .A1(n9396), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4941) );
  XNOR2_X1 U6449 ( .A(P2_IR_REG_31__SCAN_IN), .B(P2_IR_REG_27__SCAN_IN), .ZN(
        n4940) );
  OAI21_X1 U6450 ( .B1(n5581), .B2(n4941), .A(n4940), .ZN(n4942) );
  NAND3_X2 U6451 ( .A1(n4890), .A2(n4943), .A3(n4942), .ZN(n5562) );
  INV_X1 U6452 ( .A(n4945), .ZN(n4946) );
  NAND2_X2 U6453 ( .A1(n4947), .A2(n4946), .ZN(n5561) );
  MUX2_X1 U6454 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8828), .S(n6242), .Z(n10040)
         );
  NAND2_X1 U6455 ( .A1(n8464), .A2(n10040), .ZN(n7922) );
  INV_X1 U6456 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n4948) );
  NAND2_X1 U6457 ( .A1(n5011), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4951) );
  NAND2_X1 U6458 ( .A1(n5084), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n4950) );
  NAND2_X1 U6459 ( .A1(n4971), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4949) );
  INV_X1 U6460 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6741) );
  NAND2_X1 U6461 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4953) );
  INV_X1 U6462 ( .A(n4954), .ZN(n4955) );
  OAI22_X1 U6463 ( .A1(n4997), .A2(n6741), .B1(n6242), .B2(n6952), .ZN(n4957)
         );
  INV_X1 U6464 ( .A(n4957), .ZN(n4968) );
  INV_X1 U6465 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5707) );
  OAI21_X1 U6466 ( .B1(n5000), .B2(P1_DATAO_REG_0__SCAN_IN), .A(n4958), .ZN(
        n4960) );
  INV_X1 U6467 ( .A(SI_0_), .ZN(n4959) );
  INV_X1 U6468 ( .A(n4962), .ZN(n4965) );
  INV_X1 U6469 ( .A(n4963), .ZN(n4964) );
  NAND2_X1 U6470 ( .A1(n4965), .A2(n4964), .ZN(n4978) );
  NAND2_X1 U6471 ( .A1(n4977), .A2(n4978), .ZN(n4966) );
  INV_X1 U6472 ( .A(SI_1_), .ZN(n4976) );
  XNOR2_X1 U6473 ( .A(n4966), .B(n4976), .ZN(n6740) );
  OR2_X1 U6474 ( .A1(n5039), .A2(n6740), .ZN(n4967) );
  NAND2_X1 U6475 ( .A1(n7922), .A2(n8380), .ZN(n4970) );
  NAND2_X1 U6476 ( .A1(n6984), .A2(n6983), .ZN(n4969) );
  NAND2_X1 U6477 ( .A1(n4970), .A2(n4969), .ZN(n7145) );
  NAND2_X1 U6478 ( .A1(n5084), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n4974) );
  NAND2_X1 U6479 ( .A1(n4971), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4973) );
  NAND2_X1 U6480 ( .A1(n5011), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4972) );
  OR2_X1 U6481 ( .A1(n4997), .A2(n4523), .ZN(n4986) );
  NAND2_X1 U6482 ( .A1(n4977), .A2(n4976), .ZN(n4979) );
  NAND2_X1 U6483 ( .A1(n4979), .A2(n4978), .ZN(n4983) );
  INV_X1 U6484 ( .A(n4983), .ZN(n4981) );
  INV_X1 U6485 ( .A(n4982), .ZN(n4980) );
  NAND2_X1 U6486 ( .A1(n4983), .A2(n4982), .ZN(n4984) );
  NAND2_X1 U6487 ( .A1(n4999), .A2(n4984), .ZN(n6746) );
  OR2_X1 U6488 ( .A1(n5039), .A2(n6746), .ZN(n4985) );
  OAI211_X1 U6489 ( .C1(n6242), .C2(n7049), .A(n4986), .B(n4985), .ZN(n7126)
         );
  NAND2_X1 U6490 ( .A1(n4987), .A2(n7126), .ZN(n8227) );
  INV_X1 U6491 ( .A(n7126), .ZN(n6979) );
  NAND2_X1 U6492 ( .A1(n7145), .A2(n8381), .ZN(n4989) );
  NAND2_X1 U6493 ( .A1(n4987), .A2(n6979), .ZN(n4988) );
  NAND2_X1 U6494 ( .A1(n4989), .A2(n4988), .ZN(n7077) );
  INV_X2 U6495 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7224) );
  NAND2_X1 U6496 ( .A1(n5312), .A2(n7224), .ZN(n4993) );
  NAND2_X1 U6497 ( .A1(n4971), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4992) );
  NAND2_X1 U6498 ( .A1(n8367), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n4991) );
  NAND2_X1 U6499 ( .A1(n5011), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4990) );
  NAND2_X1 U6500 ( .A1(n4975), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4994) );
  MUX2_X1 U6501 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4994), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n4996) );
  NAND2_X1 U6502 ( .A1(n4996), .A2(n4995), .ZN(n6922) );
  INV_X1 U6503 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9302) );
  NAND2_X1 U6504 ( .A1(n4999), .A2(n4998), .ZN(n5005) );
  MUX2_X1 U6505 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5000), .Z(n5001) );
  OAI21_X1 U6506 ( .B1(n5001), .B2(SI_3_), .A(n5018), .ZN(n5003) );
  NAND2_X1 U6507 ( .A1(n5002), .A2(n5003), .ZN(n5006) );
  INV_X1 U6508 ( .A(n5003), .ZN(n5004) );
  NAND2_X1 U6509 ( .A1(n5005), .A2(n5004), .ZN(n5019) );
  NAND2_X1 U6510 ( .A1(n5006), .A2(n5019), .ZN(n6737) );
  NAND2_X1 U6511 ( .A1(n7146), .A2(n7225), .ZN(n8243) );
  INV_X1 U6512 ( .A(n7146), .ZN(n8461) );
  INV_X1 U6513 ( .A(n7225), .ZN(n7082) );
  NAND2_X1 U6514 ( .A1(n8461), .A2(n7082), .ZN(n8237) );
  NAND2_X1 U6515 ( .A1(n8243), .A2(n8237), .ZN(n8379) );
  NAND2_X1 U6516 ( .A1(n7077), .A2(n8379), .ZN(n5008) );
  NAND2_X1 U6517 ( .A1(n7146), .A2(n7082), .ZN(n5007) );
  NAND2_X1 U6518 ( .A1(n4971), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5015) );
  NAND2_X1 U6519 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5010) );
  NAND2_X1 U6520 ( .A1(n5031), .A2(n5010), .ZN(n7195) );
  NAND2_X1 U6521 ( .A1(n5084), .A2(n7195), .ZN(n5014) );
  INV_X2 U6522 ( .A(n5565), .ZN(n8368) );
  NAND2_X1 U6523 ( .A1(n8368), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5013) );
  NAND2_X1 U6524 ( .A1(n8367), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5012) );
  NAND4_X1 U6525 ( .A1(n5015), .A2(n5014), .A3(n5013), .A4(n5012), .ZN(n8460)
         );
  NAND2_X1 U6526 ( .A1(n4995), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5017) );
  INV_X1 U6527 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5016) );
  INV_X1 U6528 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6739) );
  OR2_X1 U6529 ( .A1(n4997), .A2(n6739), .ZN(n5027) );
  NAND2_X1 U6530 ( .A1(n5019), .A2(n5018), .ZN(n5024) );
  MUX2_X1 U6531 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n6735), .Z(n5020) );
  NAND2_X1 U6532 ( .A1(n5020), .A2(SI_4_), .ZN(n5040) );
  OAI21_X1 U6533 ( .B1(n5020), .B2(SI_4_), .A(n5040), .ZN(n5022) );
  NAND2_X1 U6534 ( .A1(n5021), .A2(n5022), .ZN(n5025) );
  INV_X1 U6535 ( .A(n5022), .ZN(n5023) );
  NAND2_X1 U6536 ( .A1(n5025), .A2(n5041), .ZN(n6738) );
  OR2_X1 U6537 ( .A1(n5039), .A2(n6738), .ZN(n5026) );
  OAI211_X1 U6538 ( .C1(n6242), .C2(n6972), .A(n5027), .B(n5026), .ZN(n8245)
         );
  NAND2_X1 U6539 ( .A1(n8460), .A2(n8245), .ZN(n5529) );
  NAND2_X1 U6540 ( .A1(n7135), .A2(n5529), .ZN(n5028) );
  NAND2_X1 U6541 ( .A1(n7160), .A2(n8234), .ZN(n8233) );
  NAND2_X1 U6542 ( .A1(n4971), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5036) );
  NAND2_X1 U6543 ( .A1(n5031), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5032) );
  NAND2_X1 U6544 ( .A1(n5051), .A2(n5032), .ZN(n7207) );
  NAND2_X1 U6545 ( .A1(n5312), .A2(n7207), .ZN(n5035) );
  NAND2_X1 U6546 ( .A1(n8368), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5034) );
  NAND2_X1 U6547 ( .A1(n8367), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5033) );
  NAND4_X1 U6548 ( .A1(n5036), .A2(n5035), .A3(n5034), .A4(n5033), .ZN(n8459)
         );
  OR2_X1 U6549 ( .A1(n5037), .A2(n8816), .ZN(n5038) );
  XNOR2_X1 U6550 ( .A(n5038), .B(n5066), .ZN(n6749) );
  NAND2_X1 U6551 ( .A1(n5041), .A2(n5040), .ZN(n5047) );
  MUX2_X1 U6552 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6735), .Z(n5042) );
  NAND2_X1 U6553 ( .A1(n5042), .A2(SI_5_), .ZN(n5057) );
  INV_X1 U6554 ( .A(n5042), .ZN(n5044) );
  INV_X1 U6555 ( .A(SI_5_), .ZN(n5043) );
  NAND2_X1 U6556 ( .A1(n5044), .A2(n5043), .ZN(n5045) );
  NAND2_X1 U6557 ( .A1(n5047), .A2(n5046), .ZN(n5058) );
  OR2_X1 U6558 ( .A1(n5047), .A2(n5046), .ZN(n5048) );
  NAND2_X1 U6559 ( .A1(n5058), .A2(n5048), .ZN(n6748) );
  OR2_X1 U6560 ( .A1(n5039), .A2(n6748), .ZN(n5050) );
  INV_X1 U6561 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6747) );
  OR2_X1 U6562 ( .A1(n4997), .A2(n6747), .ZN(n5049) );
  OAI211_X1 U6563 ( .C1(n6242), .C2(n6749), .A(n5050), .B(n5049), .ZN(n7220)
         );
  NOR2_X1 U6564 ( .A1(n8459), .A2(n7220), .ZN(n7201) );
  NAND2_X1 U6565 ( .A1(n8459), .A2(n7220), .ZN(n7199) );
  NAND2_X1 U6566 ( .A1(n4971), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5056) );
  NAND2_X1 U6567 ( .A1(n5051), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5052) );
  NAND2_X1 U6568 ( .A1(n5092), .A2(n5052), .ZN(n7442) );
  NAND2_X1 U6569 ( .A1(n5312), .A2(n7442), .ZN(n5055) );
  NAND2_X1 U6570 ( .A1(n5011), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5054) );
  NAND2_X1 U6571 ( .A1(n8367), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U6572 ( .A1(n5058), .A2(n5057), .ZN(n5064) );
  MUX2_X1 U6573 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6735), .Z(n5059) );
  NAND2_X1 U6574 ( .A1(n5059), .A2(SI_6_), .ZN(n5074) );
  INV_X1 U6575 ( .A(n5059), .ZN(n5061) );
  INV_X1 U6576 ( .A(SI_6_), .ZN(n5060) );
  NAND2_X1 U6577 ( .A1(n5061), .A2(n5060), .ZN(n5062) );
  OR2_X1 U6578 ( .A1(n5064), .A2(n5063), .ZN(n5065) );
  NAND2_X1 U6579 ( .A1(n5075), .A2(n5065), .ZN(n6744) );
  OR2_X1 U6580 ( .A1(n6744), .A2(n5039), .ZN(n5070) );
  INV_X1 U6581 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6743) );
  OR2_X1 U6582 ( .A1(n4997), .A2(n6743), .ZN(n5069) );
  NAND2_X1 U6583 ( .A1(n5037), .A2(n5066), .ZN(n5072) );
  NAND2_X1 U6584 ( .A1(n5072), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5067) );
  XNOR2_X1 U6585 ( .A(n5067), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6324) );
  NAND2_X1 U6586 ( .A1(n5327), .A2(n6324), .ZN(n5068) );
  NAND2_X1 U6587 ( .A1(n7378), .A2(n10046), .ZN(n5071) );
  NAND2_X1 U6588 ( .A1(n7438), .A2(n5071), .ZN(n7461) );
  INV_X1 U6589 ( .A(n10046), .ZN(n7443) );
  NAND2_X1 U6590 ( .A1(n8458), .A2(n7443), .ZN(n7460) );
  NAND2_X1 U6591 ( .A1(n5113), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5073) );
  XNOR2_X1 U6592 ( .A(n5073), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6284) );
  AOI22_X1 U6593 ( .A1(n5509), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5327), .B2(
        n6284), .ZN(n5081) );
  INV_X1 U6594 ( .A(n5076), .ZN(n5078) );
  INV_X1 U6595 ( .A(SI_7_), .ZN(n5077) );
  NAND2_X1 U6596 ( .A1(n5078), .A2(n5077), .ZN(n5079) );
  MUX2_X1 U6597 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n6735), .Z(n5108) );
  NAND2_X1 U6598 ( .A1(n4971), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5088) );
  OR2_X2 U6599 ( .A1(n5094), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5119) );
  NAND2_X1 U6600 ( .A1(n5094), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5083) );
  NAND2_X1 U6601 ( .A1(n5119), .A2(n5083), .ZN(n7631) );
  NAND2_X1 U6602 ( .A1(n5084), .A2(n7631), .ZN(n5087) );
  NAND2_X1 U6603 ( .A1(n8368), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U6604 ( .A1(n8367), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5085) );
  NAND2_X1 U6605 ( .A1(n10060), .A2(n5090), .ZN(n5107) );
  NAND2_X1 U6606 ( .A1(n10060), .A2(n7592), .ZN(n8263) );
  INV_X1 U6607 ( .A(n8391), .ZN(n5091) );
  NAND2_X1 U6608 ( .A1(n4971), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5098) );
  NAND2_X1 U6609 ( .A1(n5092), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5093) );
  NAND2_X1 U6610 ( .A1(n5094), .A2(n5093), .ZN(n7465) );
  NAND2_X1 U6611 ( .A1(n5312), .A2(n7465), .ZN(n5097) );
  NAND2_X1 U6612 ( .A1(n8368), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5096) );
  NAND2_X1 U6613 ( .A1(n8367), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5095) );
  OR2_X1 U6614 ( .A1(n5100), .A2(n5099), .ZN(n5101) );
  NAND2_X1 U6615 ( .A1(n5102), .A2(n5101), .ZN(n6750) );
  OR2_X1 U6616 ( .A1(n6750), .A2(n5039), .ZN(n5106) );
  NAND2_X1 U6617 ( .A1(n5103), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5104) );
  XNOR2_X1 U6618 ( .A(n5104), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6328) );
  AOI22_X1 U6619 ( .A1(n5509), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5327), .B2(
        n6328), .ZN(n5105) );
  NAND2_X1 U6620 ( .A1(n5106), .A2(n5105), .ZN(n7375) );
  NAND2_X1 U6621 ( .A1(n8457), .A2(n7375), .ZN(n7626) );
  INV_X1 U6622 ( .A(n5108), .ZN(n5110) );
  INV_X1 U6623 ( .A(SI_8_), .ZN(n5109) );
  MUX2_X1 U6624 ( .A(n6768), .B(n6771), .S(n6735), .Z(n5134) );
  XNOR2_X1 U6625 ( .A(n5137), .B(n5136), .ZN(n6767) );
  NAND2_X1 U6626 ( .A1(n6767), .A2(n8209), .ZN(n5116) );
  OAI21_X1 U6627 ( .B1(n5113), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5114) );
  XNOR2_X1 U6628 ( .A(n5114), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7348) );
  AOI22_X1 U6629 ( .A1(n5509), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5327), .B2(
        n7348), .ZN(n5115) );
  NAND2_X1 U6630 ( .A1(n5116), .A2(n5115), .ZN(n10065) );
  NAND2_X1 U6631 ( .A1(n5513), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5124) );
  NAND2_X1 U6632 ( .A1(n5119), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5120) );
  NAND2_X1 U6633 ( .A1(n5150), .A2(n5120), .ZN(n7555) );
  NAND2_X1 U6634 ( .A1(n5312), .A2(n7555), .ZN(n5123) );
  NAND2_X1 U6635 ( .A1(n8368), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U6636 ( .A1(n8367), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5121) );
  NAND4_X1 U6637 ( .A1(n5124), .A2(n5123), .A3(n5122), .A4(n5121), .ZN(n8456)
         );
  NAND2_X1 U6638 ( .A1(n7548), .A2(n4366), .ZN(n5125) );
  OR2_X1 U6639 ( .A1(n10065), .A2(n8456), .ZN(n5129) );
  NAND2_X1 U6640 ( .A1(n5125), .A2(n5129), .ZN(n5127) );
  NAND2_X1 U6641 ( .A1(n7461), .A2(n5126), .ZN(n5133) );
  INV_X1 U6642 ( .A(n5127), .ZN(n5131) );
  NAND2_X1 U6643 ( .A1(n7364), .A2(n7375), .ZN(n8262) );
  INV_X1 U6644 ( .A(n7375), .ZN(n10051) );
  NAND2_X1 U6645 ( .A1(n8457), .A2(n10051), .ZN(n7622) );
  NAND2_X1 U6646 ( .A1(n8262), .A2(n7622), .ZN(n8256) );
  AND2_X1 U6647 ( .A1(n8256), .A2(n5128), .ZN(n7547) );
  AND2_X1 U6648 ( .A1(n7547), .A2(n5129), .ZN(n5130) );
  INV_X1 U6649 ( .A(n5134), .ZN(n5135) );
  MUX2_X1 U6650 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6735), .Z(n5138) );
  NAND2_X1 U6651 ( .A1(n5138), .A2(SI_10_), .ZN(n5156) );
  INV_X1 U6652 ( .A(n5138), .ZN(n5140) );
  INV_X1 U6653 ( .A(SI_10_), .ZN(n5139) );
  NAND2_X1 U6654 ( .A1(n5140), .A2(n5139), .ZN(n5141) );
  NAND2_X1 U6655 ( .A1(n5156), .A2(n5141), .ZN(n5143) );
  NAND2_X1 U6656 ( .A1(n4380), .A2(n5143), .ZN(n5144) );
  NAND2_X1 U6657 ( .A1(n5157), .A2(n5144), .ZN(n6774) );
  OR2_X1 U6658 ( .A1(n6774), .A2(n5039), .ZN(n5149) );
  OR2_X1 U6659 ( .A1(n5145), .A2(n8816), .ZN(n5147) );
  XNOR2_X1 U6660 ( .A(n5147), .B(n5146), .ZN(n6775) );
  INV_X1 U6661 ( .A(n6775), .ZN(n7719) );
  AOI22_X1 U6662 ( .A1(n5509), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5327), .B2(
        n7719), .ZN(n5148) );
  NAND2_X1 U6663 ( .A1(n5149), .A2(n5148), .ZN(n7839) );
  NAND2_X1 U6664 ( .A1(n5513), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5155) );
  OR2_X2 U6665 ( .A1(n5150), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U6666 ( .A1(n5150), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5151) );
  NAND2_X1 U6667 ( .A1(n5165), .A2(n5151), .ZN(n7641) );
  NAND2_X1 U6668 ( .A1(n5312), .A2(n7641), .ZN(n5154) );
  NAND2_X1 U6669 ( .A1(n8368), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5153) );
  NAND2_X1 U6670 ( .A1(n8367), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5152) );
  NAND4_X1 U6671 ( .A1(n5155), .A2(n5154), .A3(n5153), .A4(n5152), .ZN(n8455)
         );
  INV_X1 U6672 ( .A(n8455), .ZN(n7581) );
  NAND2_X1 U6673 ( .A1(n5157), .A2(n5156), .ZN(n5174) );
  MUX2_X1 U6674 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6735), .Z(n5172) );
  XNOR2_X1 U6675 ( .A(n5174), .B(n5173), .ZN(n6816) );
  NAND2_X1 U6676 ( .A1(n6816), .A2(n8209), .ZN(n5164) );
  INV_X1 U6677 ( .A(n5158), .ZN(n5160) );
  NAND2_X1 U6678 ( .A1(n5160), .A2(n5159), .ZN(n5208) );
  NAND2_X1 U6679 ( .A1(n5158), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5161) );
  MUX2_X1 U6680 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5161), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n5162) );
  AND2_X1 U6681 ( .A1(n5208), .A2(n5162), .ZN(n7812) );
  AOI22_X1 U6682 ( .A1(n5509), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5327), .B2(
        n7812), .ZN(n5163) );
  NAND2_X1 U6683 ( .A1(n5164), .A2(n5163), .ZN(n7900) );
  NAND2_X1 U6684 ( .A1(n5513), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6685 ( .A1(n5165), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6686 ( .A1(n5184), .A2(n5166), .ZN(n7910) );
  NAND2_X1 U6687 ( .A1(n5312), .A2(n7910), .ZN(n5169) );
  NAND2_X1 U6688 ( .A1(n8368), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U6689 ( .A1(n8367), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6690 ( .A1(n7900), .A2(n7661), .ZN(n8277) );
  NAND2_X1 U6691 ( .A1(n8275), .A2(n8277), .ZN(n7578) );
  INV_X1 U6692 ( .A(n7661), .ZN(n8454) );
  NAND2_X1 U6693 ( .A1(n7900), .A2(n8454), .ZN(n5171) );
  MUX2_X1 U6694 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6735), .Z(n5175) );
  NAND2_X1 U6695 ( .A1(n5177), .A2(n5176), .ZN(n5178) );
  OR2_X1 U6696 ( .A1(n6823), .A2(n5039), .ZN(n5181) );
  NAND2_X1 U6697 ( .A1(n5208), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5179) );
  XNOR2_X1 U6698 ( .A(n5179), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7891) );
  AOI22_X1 U6699 ( .A1(n5509), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5327), .B2(
        n7891), .ZN(n5180) );
  NAND2_X1 U6700 ( .A1(n8368), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5189) );
  NAND2_X1 U6701 ( .A1(n5513), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5188) );
  INV_X1 U6702 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U6703 ( .A1(n5184), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6704 ( .A1(n5194), .A2(n5185), .ZN(n8101) );
  NAND2_X1 U6705 ( .A1(n5312), .A2(n8101), .ZN(n5187) );
  NAND2_X1 U6706 ( .A1(n8367), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6707 ( .A1(n10080), .A2(n8156), .ZN(n5191) );
  AND2_X1 U6708 ( .A1(n7664), .A2(n8453), .ZN(n5190) );
  INV_X1 U6709 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6710 ( .A1(n5194), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5195) );
  NAND2_X1 U6711 ( .A1(n5228), .A2(n5195), .ZN(n8158) );
  NAND2_X1 U6712 ( .A1(n5312), .A2(n8158), .ZN(n5199) );
  NAND2_X1 U6713 ( .A1(n5513), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6714 ( .A1(n8367), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6715 ( .A1(n8368), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5196) );
  MUX2_X1 U6716 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6735), .Z(n5202) );
  NAND2_X1 U6717 ( .A1(n5202), .A2(SI_13_), .ZN(n5213) );
  INV_X1 U6718 ( .A(n5202), .ZN(n5204) );
  INV_X1 U6719 ( .A(SI_13_), .ZN(n5203) );
  NAND2_X1 U6720 ( .A1(n5204), .A2(n5203), .ZN(n5205) );
  NAND2_X1 U6721 ( .A1(n6828), .A2(n8209), .ZN(n5212) );
  INV_X1 U6722 ( .A(n5208), .ZN(n5210) );
  NAND2_X1 U6723 ( .A1(n5210), .A2(n5209), .ZN(n5271) );
  NAND2_X1 U6724 ( .A1(n5271), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5221) );
  XNOR2_X1 U6725 ( .A(n5221), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7869) );
  AOI22_X1 U6726 ( .A1(n5509), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5327), .B2(
        n7869), .ZN(n5211) );
  MUX2_X1 U6727 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6735), .Z(n5215) );
  NAND2_X1 U6728 ( .A1(n5215), .A2(SI_14_), .ZN(n5236) );
  INV_X1 U6729 ( .A(n5215), .ZN(n5217) );
  INV_X1 U6730 ( .A(SI_14_), .ZN(n5216) );
  NAND2_X1 U6731 ( .A1(n5217), .A2(n5216), .ZN(n5218) );
  OR2_X1 U6732 ( .A1(n6858), .A2(n5039), .ZN(n5227) );
  NAND2_X1 U6733 ( .A1(n5221), .A2(n5268), .ZN(n5222) );
  NAND2_X1 U6734 ( .A1(n5222), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5224) );
  INV_X1 U6735 ( .A(n5224), .ZN(n5223) );
  NAND2_X1 U6736 ( .A1(n5223), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6737 ( .A1(n5224), .A2(n5269), .ZN(n5245) );
  AOI22_X1 U6738 ( .A1(n5509), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5327), .B2(
        n8479), .ZN(n5226) );
  NOR2_X1 U6739 ( .A1(n7894), .A2(n9640), .ZN(n5235) );
  NAND2_X1 U6740 ( .A1(n5513), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U6741 ( .A1(n5228), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5229) );
  NAND2_X1 U6742 ( .A1(n5251), .A2(n5229), .ZN(n8070) );
  NAND2_X1 U6743 ( .A1(n5312), .A2(n8070), .ZN(n5232) );
  NAND2_X1 U6744 ( .A1(n8368), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5231) );
  NAND2_X1 U6745 ( .A1(n8367), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5230) );
  NAND4_X1 U6746 ( .A1(n5233), .A2(n5232), .A3(n5231), .A4(n5230), .ZN(n8451)
         );
  INV_X1 U6747 ( .A(n9640), .ZN(n5541) );
  OAI22_X1 U6748 ( .A1(n5235), .A2(n8451), .B1(n5541), .B2(n5234), .ZN(n8689)
         );
  MUX2_X1 U6749 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n5000), .Z(n5238) );
  NAND2_X1 U6750 ( .A1(n5238), .A2(SI_15_), .ZN(n5258) );
  INV_X1 U6751 ( .A(n5238), .ZN(n5240) );
  INV_X1 U6752 ( .A(SI_15_), .ZN(n5239) );
  NAND2_X1 U6753 ( .A1(n5240), .A2(n5239), .ZN(n5241) );
  NAND2_X1 U6754 ( .A1(n5259), .A2(n5244), .ZN(n6895) );
  OR2_X1 U6755 ( .A1(n6895), .A2(n5039), .ZN(n5248) );
  NAND2_X1 U6756 ( .A1(n5245), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5246) );
  XNOR2_X1 U6757 ( .A(n5246), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8497) );
  AOI22_X1 U6758 ( .A1(n5509), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5327), .B2(
        n8497), .ZN(n5247) );
  NAND2_X1 U6759 ( .A1(n5513), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U6760 ( .A1(n8368), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5255) );
  INV_X1 U6761 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6762 ( .A1(n5251), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6763 ( .A1(n5278), .A2(n5252), .ZN(n8696) );
  NAND2_X1 U6764 ( .A1(n5312), .A2(n8696), .ZN(n5254) );
  NAND2_X1 U6765 ( .A1(n8367), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5253) );
  NAND2_X1 U6766 ( .A1(n8748), .A2(n8678), .ZN(n8303) );
  NAND2_X1 U6767 ( .A1(n8295), .A2(n8303), .ZN(n8399) );
  INV_X1 U6768 ( .A(n8748), .ZN(n8208) );
  MUX2_X1 U6769 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n5000), .Z(n5260) );
  NAND2_X1 U6770 ( .A1(n5260), .A2(SI_16_), .ZN(n5286) );
  INV_X1 U6771 ( .A(n5260), .ZN(n5262) );
  INV_X1 U6772 ( .A(SI_16_), .ZN(n5261) );
  NAND2_X1 U6773 ( .A1(n5262), .A2(n5261), .ZN(n5263) );
  OR2_X1 U6774 ( .A1(n5265), .A2(n5264), .ZN(n5266) );
  NAND2_X1 U6775 ( .A1(n5287), .A2(n5266), .ZN(n6953) );
  OR2_X1 U6776 ( .A1(n6953), .A2(n5039), .ZN(n5277) );
  NAND3_X1 U6777 ( .A1(n5269), .A2(n5268), .A3(n5267), .ZN(n5270) );
  NOR2_X1 U6778 ( .A1(n5274), .A2(n8816), .ZN(n5272) );
  MUX2_X1 U6779 ( .A(n8816), .B(n5272), .S(P2_IR_REG_16__SCAN_IN), .Z(n5275)
         );
  NAND2_X1 U6780 ( .A1(n5274), .A2(n5273), .ZN(n5307) );
  NOR2_X1 U6781 ( .A1(n5275), .A2(n5308), .ZN(n8517) );
  AOI22_X1 U6782 ( .A1(n5509), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5327), .B2(
        n8517), .ZN(n5276) );
  NAND2_X1 U6783 ( .A1(n8368), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5283) );
  NAND2_X1 U6784 ( .A1(n5513), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5282) );
  OR2_X2 U6785 ( .A1(n5278), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5292) );
  NAND2_X1 U6786 ( .A1(n5278), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5279) );
  NAND2_X1 U6787 ( .A1(n5292), .A2(n5279), .ZN(n8684) );
  NAND2_X1 U6788 ( .A1(n5312), .A2(n8684), .ZN(n5281) );
  NAND2_X1 U6789 ( .A1(n8367), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U6790 ( .A1(n8807), .A2(n8694), .ZN(n8297) );
  NAND2_X1 U6791 ( .A1(n8305), .A2(n8297), .ZN(n8674) );
  NAND2_X1 U6792 ( .A1(n8673), .A2(n8674), .ZN(n8680) );
  NAND2_X1 U6793 ( .A1(n8807), .A2(n5284), .ZN(n5285) );
  MUX2_X1 U6794 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n4425), .Z(n5300) );
  XNOR2_X1 U6795 ( .A(n5300), .B(SI_17_), .ZN(n5301) );
  XNOR2_X1 U6796 ( .A(n5302), .B(n5301), .ZN(n7088) );
  NAND2_X1 U6797 ( .A1(n7088), .A2(n8209), .ZN(n5290) );
  NAND2_X1 U6798 ( .A1(n5307), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5288) );
  XNOR2_X1 U6799 ( .A(n5288), .B(P2_IR_REG_17__SCAN_IN), .ZN(n7087) );
  AOI22_X1 U6800 ( .A1(n5509), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5327), .B2(
        n7087), .ZN(n5289) );
  NAND2_X1 U6801 ( .A1(n5513), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5297) );
  INV_X1 U6802 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10034) );
  NAND2_X1 U6803 ( .A1(n5292), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6804 ( .A1(n5313), .A2(n5293), .ZN(n8128) );
  NAND2_X1 U6805 ( .A1(n5312), .A2(n8128), .ZN(n5296) );
  NAND2_X1 U6806 ( .A1(n8368), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5295) );
  NAND2_X1 U6807 ( .A1(n8367), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U6808 ( .A1(n7992), .A2(n8677), .ZN(n8666) );
  NAND2_X1 U6809 ( .A1(n8663), .A2(n8666), .ZN(n7937) );
  INV_X1 U6810 ( .A(n7992), .ZN(n8131) );
  MUX2_X1 U6811 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5000), .Z(n5303) );
  NAND2_X1 U6812 ( .A1(n5303), .A2(SI_18_), .ZN(n5320) );
  OAI21_X1 U6813 ( .B1(n5303), .B2(SI_18_), .A(n5320), .ZN(n5304) );
  NAND2_X1 U6814 ( .A1(n5305), .A2(n5304), .ZN(n5306) );
  INV_X1 U6815 ( .A(n5307), .ZN(n5308) );
  NAND2_X1 U6816 ( .A1(n5308), .A2(n4917), .ZN(n5309) );
  XNOR2_X1 U6817 ( .A(n5323), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8530) );
  AOI22_X1 U6818 ( .A1(n5509), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5327), .B2(
        n8530), .ZN(n5310) );
  NAND2_X1 U6819 ( .A1(n5513), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5318) );
  NAND2_X1 U6820 ( .A1(n8367), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6821 ( .A1(n5313), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5314) );
  NAND2_X1 U6822 ( .A1(n5332), .A2(n5314), .ZN(n8658) );
  NAND2_X1 U6823 ( .A1(n5312), .A2(n8658), .ZN(n5316) );
  NAND2_X1 U6824 ( .A1(n8368), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5315) );
  NAND2_X1 U6825 ( .A1(n8742), .A2(n8644), .ZN(n5319) );
  INV_X1 U6826 ( .A(n8644), .ZN(n8449) );
  MUX2_X1 U6827 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n4425), .Z(n5339) );
  XNOR2_X1 U6828 ( .A(n5339), .B(SI_19_), .ZN(n5338) );
  XNOR2_X1 U6829 ( .A(n5337), .B(n5338), .ZN(n7231) );
  NAND2_X1 U6830 ( .A1(n7231), .A2(n8209), .ZN(n5329) );
  INV_X1 U6831 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6832 ( .A1(n5323), .A2(n5322), .ZN(n5324) );
  XNOR2_X2 U6833 ( .A(n5326), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8433) );
  AOI22_X1 U6834 ( .A1(n5509), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8433), .B2(
        n5327), .ZN(n5328) );
  INV_X1 U6835 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5330) );
  NAND2_X1 U6836 ( .A1(n5332), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6837 ( .A1(n5345), .A2(n5333), .ZN(n8646) );
  AOI22_X1 U6838 ( .A1(n8646), .A2(n5312), .B1(n5011), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n5335) );
  AOI22_X1 U6839 ( .A1(n5513), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n8367), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6840 ( .A1(n8735), .A2(n8631), .ZN(n8312) );
  INV_X1 U6841 ( .A(n8735), .ZN(n5336) );
  INV_X1 U6842 ( .A(n5339), .ZN(n5340) );
  INV_X1 U6843 ( .A(SI_19_), .ZN(n9323) );
  NAND2_X1 U6844 ( .A1(n5340), .A2(n9323), .ZN(n5341) );
  NAND2_X1 U6845 ( .A1(n5342), .A2(n5341), .ZN(n5351) );
  INV_X1 U6846 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7436) );
  INV_X1 U6847 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7472) );
  MUX2_X1 U6848 ( .A(n7436), .B(n7472), .S(n4425), .Z(n5353) );
  XNOR2_X1 U6849 ( .A(n5353), .B(SI_20_), .ZN(n5350) );
  XNOR2_X1 U6850 ( .A(n5351), .B(n5350), .ZN(n7435) );
  NAND2_X1 U6851 ( .A1(n7435), .A2(n8209), .ZN(n5344) );
  NAND2_X1 U6852 ( .A1(n5509), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5343) );
  OR2_X2 U6853 ( .A1(n5345), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U6854 ( .A1(n5345), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6855 ( .A1(n5360), .A2(n5346), .ZN(n8633) );
  NAND2_X1 U6856 ( .A1(n8633), .A2(n5312), .ZN(n5349) );
  AOI22_X1 U6857 ( .A1(n5513), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n5011), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U6858 ( .A1(n8367), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U6859 ( .A1(n8731), .A2(n8645), .ZN(n8319) );
  INV_X1 U6860 ( .A(n8645), .ZN(n8448) );
  NOR2_X1 U6861 ( .A1(n8731), .A2(n8448), .ZN(n8616) );
  INV_X1 U6862 ( .A(SI_20_), .ZN(n5352) );
  NAND2_X1 U6863 ( .A1(n5353), .A2(n5352), .ZN(n5354) );
  INV_X1 U6864 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7530) );
  INV_X1 U6865 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7531) );
  MUX2_X1 U6866 ( .A(n7530), .B(n7531), .S(n4425), .Z(n5368) );
  XNOR2_X1 U6867 ( .A(n5368), .B(SI_21_), .ZN(n5355) );
  XNOR2_X1 U6868 ( .A(n5365), .B(n5355), .ZN(n7529) );
  NAND2_X1 U6869 ( .A1(n7529), .A2(n8209), .ZN(n5357) );
  NAND2_X1 U6870 ( .A1(n5509), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5356) );
  INV_X1 U6871 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U6872 ( .A1(n5360), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6873 ( .A1(n5378), .A2(n5361), .ZN(n8623) );
  NAND2_X1 U6874 ( .A1(n8623), .A2(n5312), .ZN(n5364) );
  AOI22_X1 U6875 ( .A1(n5513), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n5011), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n5363) );
  NAND2_X1 U6876 ( .A1(n8367), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6877 ( .A1(n8624), .A2(n8632), .ZN(n8326) );
  NAND2_X1 U6878 ( .A1(n8332), .A2(n8326), .ZN(n8615) );
  INV_X1 U6879 ( .A(n8624), .ZN(n8792) );
  NAND2_X1 U6880 ( .A1(n8792), .A2(n8632), .ZN(n8603) );
  NAND2_X1 U6881 ( .A1(n8614), .A2(n8603), .ZN(n5386) );
  INV_X1 U6882 ( .A(SI_21_), .ZN(n5366) );
  NAND2_X1 U6883 ( .A1(n5368), .A2(n5366), .ZN(n5367) );
  INV_X1 U6884 ( .A(n5368), .ZN(n5369) );
  NAND2_X1 U6885 ( .A1(n5369), .A2(SI_21_), .ZN(n5370) );
  INV_X1 U6886 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7588) );
  INV_X1 U6887 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9413) );
  MUX2_X1 U6888 ( .A(n7588), .B(n9413), .S(n4425), .Z(n5373) );
  INV_X1 U6889 ( .A(SI_22_), .ZN(n5372) );
  NAND2_X1 U6890 ( .A1(n5373), .A2(n5372), .ZN(n5407) );
  INV_X1 U6891 ( .A(n5373), .ZN(n5374) );
  NAND2_X1 U6892 ( .A1(n5374), .A2(SI_22_), .ZN(n5375) );
  NAND2_X1 U6893 ( .A1(n5407), .A2(n5375), .ZN(n5405) );
  XNOR2_X1 U6894 ( .A(n5435), .B(n5405), .ZN(n7586) );
  NAND2_X1 U6895 ( .A1(n7586), .A2(n8209), .ZN(n5377) );
  NAND2_X1 U6896 ( .A1(n5509), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6897 ( .A1(n5378), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6898 ( .A1(n5396), .A2(n5379), .ZN(n8610) );
  NAND2_X1 U6899 ( .A1(n8610), .A2(n5312), .ZN(n5385) );
  INV_X1 U6900 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8785) );
  NAND2_X1 U6901 ( .A1(n5513), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U6902 ( .A1(n8368), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5381) );
  OAI211_X1 U6903 ( .C1(n8785), .C2(n5380), .A(n5382), .B(n5381), .ZN(n5383)
         );
  INV_X1 U6904 ( .A(n5383), .ZN(n5384) );
  NAND2_X1 U6905 ( .A1(n8786), .A2(n8620), .ZN(n8334) );
  NAND2_X1 U6906 ( .A1(n8327), .A2(n8334), .ZN(n8325) );
  INV_X1 U6907 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5389) );
  INV_X1 U6908 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5388) );
  MUX2_X1 U6909 ( .A(n5389), .B(n5388), .S(n4425), .Z(n5390) );
  INV_X1 U6910 ( .A(SI_23_), .ZN(n9395) );
  NAND2_X1 U6911 ( .A1(n5390), .A2(n9395), .ZN(n5406) );
  INV_X1 U6912 ( .A(n5390), .ZN(n5391) );
  NAND2_X1 U6913 ( .A1(n5391), .A2(SI_23_), .ZN(n5404) );
  AND2_X1 U6914 ( .A1(n5406), .A2(n5404), .ZN(n5392) );
  NAND2_X1 U6915 ( .A1(n7699), .A2(n8209), .ZN(n5395) );
  NAND2_X1 U6916 ( .A1(n5509), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5394) );
  NAND2_X1 U6917 ( .A1(n5396), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6918 ( .A1(n5419), .A2(n5397), .ZN(n8598) );
  NAND2_X1 U6919 ( .A1(n8598), .A2(n5312), .ZN(n5402) );
  INV_X1 U6920 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8779) );
  NAND2_X1 U6921 ( .A1(n5513), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U6922 ( .A1(n8368), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5398) );
  OAI211_X1 U6923 ( .C1(n8779), .C2(n5380), .A(n5399), .B(n5398), .ZN(n5400)
         );
  INV_X1 U6924 ( .A(n5400), .ZN(n5401) );
  NAND2_X1 U6925 ( .A1(n8780), .A2(n8607), .ZN(n5403) );
  INV_X1 U6926 ( .A(n5404), .ZN(n5409) );
  AND2_X1 U6927 ( .A1(n5407), .A2(n5406), .ZN(n5408) );
  INV_X1 U6928 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8058) );
  INV_X1 U6929 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7723) );
  MUX2_X1 U6930 ( .A(n8058), .B(n7723), .S(n4425), .Z(n5412) );
  INV_X1 U6931 ( .A(SI_24_), .ZN(n5411) );
  NAND2_X1 U6932 ( .A1(n5412), .A2(n5411), .ZN(n5429) );
  INV_X1 U6933 ( .A(n5412), .ZN(n5413) );
  NAND2_X1 U6934 ( .A1(n5413), .A2(SI_24_), .ZN(n5427) );
  AND2_X1 U6935 ( .A1(n5429), .A2(n5427), .ZN(n5414) );
  NAND2_X1 U6936 ( .A1(n7722), .A2(n8209), .ZN(n5417) );
  NAND2_X1 U6937 ( .A1(n5509), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5416) );
  INV_X1 U6938 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8138) );
  NAND2_X1 U6939 ( .A1(n5419), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6940 ( .A1(n5444), .A2(n5420), .ZN(n8586) );
  NAND2_X1 U6941 ( .A1(n8586), .A2(n5312), .ZN(n5425) );
  INV_X1 U6942 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8773) );
  NAND2_X1 U6943 ( .A1(n5513), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U6944 ( .A1(n8368), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5421) );
  OAI211_X1 U6945 ( .C1(n8773), .C2(n5380), .A(n5422), .B(n5421), .ZN(n5423)
         );
  INV_X1 U6946 ( .A(n5423), .ZN(n5424) );
  NAND2_X1 U6947 ( .A1(n8774), .A2(n8596), .ZN(n5553) );
  INV_X1 U6948 ( .A(n5427), .ZN(n5432) );
  INV_X1 U6949 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7913) );
  INV_X1 U6950 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7726) );
  MUX2_X1 U6951 ( .A(n7913), .B(n7726), .S(n4425), .Z(n5437) );
  INV_X1 U6952 ( .A(SI_25_), .ZN(n5436) );
  NAND2_X1 U6953 ( .A1(n5437), .A2(n5436), .ZN(n5454) );
  INV_X1 U6954 ( .A(n5437), .ZN(n5438) );
  NAND2_X1 U6955 ( .A1(n5438), .A2(SI_25_), .ZN(n5439) );
  NAND2_X1 U6956 ( .A1(n7725), .A2(n8209), .ZN(n5441) );
  NAND2_X1 U6957 ( .A1(n5509), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5440) );
  INV_X1 U6958 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U6959 ( .A1(n5444), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U6960 ( .A1(n5461), .A2(n5445), .ZN(n8574) );
  NAND2_X1 U6961 ( .A1(n8574), .A2(n5312), .ZN(n5450) );
  INV_X1 U6962 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8766) );
  NAND2_X1 U6963 ( .A1(n5513), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6964 ( .A1(n5011), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5446) );
  OAI211_X1 U6965 ( .C1(n5380), .C2(n8766), .A(n5447), .B(n5446), .ZN(n5448)
         );
  INV_X1 U6966 ( .A(n5448), .ZN(n5449) );
  NAND2_X1 U6967 ( .A1(n8767), .A2(n8584), .ZN(n8342) );
  NAND2_X1 U6968 ( .A1(n5453), .A2(n5452), .ZN(n5455) );
  INV_X1 U6969 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7794) );
  INV_X1 U6970 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7796) );
  MUX2_X1 U6971 ( .A(n7794), .B(n7796), .S(n4425), .Z(n5456) );
  INV_X1 U6972 ( .A(SI_26_), .ZN(n9384) );
  NAND2_X1 U6973 ( .A1(n5456), .A2(n9384), .ZN(n5471) );
  INV_X1 U6974 ( .A(n5456), .ZN(n5457) );
  NAND2_X1 U6975 ( .A1(n5457), .A2(SI_26_), .ZN(n5458) );
  NAND2_X1 U6976 ( .A1(n7793), .A2(n8209), .ZN(n5460) );
  NAND2_X1 U6977 ( .A1(n5509), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U6978 ( .A1(n5461), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U6979 ( .A1(n5480), .A2(n5462), .ZN(n8566) );
  NAND2_X1 U6980 ( .A1(n8566), .A2(n5312), .ZN(n5467) );
  INV_X1 U6981 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8759) );
  NAND2_X1 U6982 ( .A1(n5513), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U6983 ( .A1(n5011), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5463) );
  OAI211_X1 U6984 ( .C1(n8759), .C2(n5380), .A(n5464), .B(n5463), .ZN(n5465)
         );
  INV_X1 U6985 ( .A(n5465), .ZN(n5466) );
  NAND2_X1 U6986 ( .A1(n8711), .A2(n8573), .ZN(n5468) );
  INV_X1 U6987 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5472) );
  INV_X1 U6988 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9408) );
  MUX2_X1 U6989 ( .A(n5472), .B(n9408), .S(n4425), .Z(n5474) );
  INV_X1 U6990 ( .A(SI_27_), .ZN(n5473) );
  NAND2_X1 U6991 ( .A1(n5474), .A2(n5473), .ZN(n5491) );
  INV_X1 U6992 ( .A(n5474), .ZN(n5475) );
  NAND2_X1 U6993 ( .A1(n5475), .A2(SI_27_), .ZN(n5476) );
  NAND2_X1 U6994 ( .A1(n7827), .A2(n8209), .ZN(n5478) );
  NAND2_X1 U6995 ( .A1(n5509), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5477) );
  INV_X1 U6996 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8028) );
  NAND2_X1 U6997 ( .A1(n5480), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5481) );
  NAND2_X1 U6998 ( .A1(n5495), .A2(n5481), .ZN(n8027) );
  NAND2_X1 U6999 ( .A1(n8027), .A2(n5312), .ZN(n5487) );
  INV_X1 U7000 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U7001 ( .A1(n5513), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U7002 ( .A1(n5011), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5482) );
  OAI211_X1 U7003 ( .C1(n5484), .C2(n5380), .A(n5483), .B(n5482), .ZN(n5485)
         );
  INV_X1 U7004 ( .A(n5485), .ZN(n5486) );
  INV_X1 U7005 ( .A(n5488), .ZN(n7952) );
  INV_X1 U7006 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5492) );
  INV_X1 U7007 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8057) );
  MUX2_X1 U7008 ( .A(n5492), .B(n8057), .S(n4425), .Z(n5506) );
  XNOR2_X1 U7009 ( .A(n5506), .B(SI_28_), .ZN(n5504) );
  NAND2_X1 U7010 ( .A1(n7874), .A2(n8209), .ZN(n5494) );
  NAND2_X1 U7011 ( .A1(n5509), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U7012 ( .A1(n5495), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U7013 ( .A1(n8540), .A2(n5496), .ZN(n8043) );
  NAND2_X1 U7014 ( .A1(n8043), .A2(n5312), .ZN(n5501) );
  INV_X1 U7015 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n7955) );
  NAND2_X1 U7016 ( .A1(n5513), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U7017 ( .A1(n5011), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5497) );
  OAI211_X1 U7018 ( .C1(n7955), .C2(n5380), .A(n5498), .B(n5497), .ZN(n5499)
         );
  INV_X1 U7019 ( .A(n5499), .ZN(n5500) );
  NAND2_X2 U7020 ( .A1(n5501), .A2(n5500), .ZN(n8443) );
  NOR2_X1 U7021 ( .A1(n8358), .A2(n8443), .ZN(n5503) );
  INV_X1 U7022 ( .A(n8358), .ZN(n5502) );
  INV_X1 U7023 ( .A(n8443), .ZN(n5556) );
  OAI22_X1 U7024 ( .A1(n7952), .A2(n5503), .B1(n5502), .B2(n5556), .ZN(n5518)
         );
  NAND2_X1 U7025 ( .A1(n5505), .A2(n5504), .ZN(n5508) );
  NAND2_X1 U7026 ( .A1(n5506), .A2(n9427), .ZN(n5507) );
  INV_X1 U7027 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8825) );
  INV_X1 U7028 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8063) );
  MUX2_X1 U7029 ( .A(n8825), .B(n8063), .S(n4425), .Z(n6492) );
  NAND2_X1 U7030 ( .A1(n6446), .A2(n8209), .ZN(n5511) );
  NAND2_X1 U7031 ( .A1(n5509), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5510) );
  INV_X1 U7032 ( .A(n8540), .ZN(n5512) );
  NAND2_X1 U7033 ( .A1(n5512), .A2(n5312), .ZN(n8373) );
  INV_X1 U7034 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9316) );
  NAND2_X1 U7035 ( .A1(n5513), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5515) );
  NAND2_X1 U7036 ( .A1(n5011), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5514) );
  OAI211_X1 U7037 ( .C1(n5380), .C2(n9316), .A(n5515), .B(n5514), .ZN(n5516)
         );
  INV_X1 U7038 ( .A(n5516), .ZN(n5517) );
  AND2_X2 U7039 ( .A1(n8373), .A2(n5517), .ZN(n8046) );
  NAND2_X1 U7040 ( .A1(n5618), .A2(n8046), .ZN(n8353) );
  NAND2_X2 U7041 ( .A1(n8420), .A2(n8353), .ZN(n8356) );
  XNOR2_X1 U7042 ( .A(n5518), .B(n8356), .ZN(n5572) );
  NAND2_X1 U7043 ( .A1(n4379), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5519) );
  MUX2_X1 U7044 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5519), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n5520) );
  NAND2_X1 U7045 ( .A1(n8433), .A2(n8439), .ZN(n5610) );
  INV_X1 U7046 ( .A(n5521), .ZN(n5525) );
  NAND2_X1 U7047 ( .A1(n5525), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7048 ( .A1(n5523), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5524) );
  MUX2_X1 U7049 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5524), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5526) );
  NAND2_X1 U7050 ( .A1(n5526), .A2(n5525), .ZN(n8412) );
  INV_X1 U7051 ( .A(n8412), .ZN(n8430) );
  NAND2_X1 U7052 ( .A1(n8383), .A2(n8430), .ZN(n8426) );
  NAND2_X1 U7053 ( .A1(n7924), .A2(n10040), .ZN(n8217) );
  NAND2_X1 U7054 ( .A1(n7143), .A2(n8227), .ZN(n5528) );
  INV_X1 U7055 ( .A(n8379), .ZN(n7078) );
  NAND2_X1 U7056 ( .A1(n7160), .A2(n8245), .ZN(n8238) );
  AND2_X1 U7057 ( .A1(n8243), .A2(n8238), .ZN(n5531) );
  INV_X1 U7058 ( .A(n8238), .ZN(n5530) );
  NAND2_X1 U7059 ( .A1(n8233), .A2(n5529), .ZN(n7136) );
  NAND2_X1 U7060 ( .A1(n8458), .A2(n10046), .ZN(n8248) );
  INV_X1 U7061 ( .A(n7220), .ZN(n7217) );
  NAND2_X1 U7062 ( .A1(n8459), .A2(n7217), .ZN(n8247) );
  NAND2_X1 U7063 ( .A1(n7205), .A2(n8389), .ZN(n5533) );
  NOR2_X1 U7064 ( .A1(n8459), .A2(n7217), .ZN(n8384) );
  NAND2_X1 U7065 ( .A1(n8389), .A2(n8384), .ZN(n5532) );
  NAND2_X1 U7066 ( .A1(n7378), .A2(n7443), .ZN(n8382) );
  NAND2_X1 U7067 ( .A1(n5533), .A2(n8240), .ZN(n7458) );
  INV_X1 U7068 ( .A(n8263), .ZN(n5535) );
  OR2_X1 U7069 ( .A1(n8256), .A2(n5535), .ZN(n5534) );
  INV_X1 U7070 ( .A(n5534), .ZN(n5538) );
  AND2_X1 U7071 ( .A1(n8253), .A2(n7622), .ZN(n8261) );
  OR2_X1 U7072 ( .A1(n5535), .A2(n8261), .ZN(n5536) );
  INV_X1 U7073 ( .A(n5536), .ZN(n5537) );
  NAND2_X1 U7074 ( .A1(n10065), .A2(n7831), .ZN(n8264) );
  NAND2_X1 U7075 ( .A1(n8260), .A2(n8264), .ZN(n8392) );
  AND2_X1 U7076 ( .A1(n10068), .A2(n8455), .ZN(n8259) );
  NAND2_X1 U7077 ( .A1(n7839), .A2(n7581), .ZN(n8272) );
  NAND2_X1 U7078 ( .A1(n7577), .A2(n8396), .ZN(n5539) );
  NAND2_X1 U7079 ( .A1(n7664), .A2(n8156), .ZN(n8282) );
  NAND2_X1 U7080 ( .A1(n8281), .A2(n8282), .ZN(n8284) );
  NOR2_X1 U7081 ( .A1(n9646), .A2(n8099), .ZN(n8287) );
  NAND2_X1 U7082 ( .A1(n9646), .A2(n8099), .ZN(n8285) );
  NAND2_X1 U7083 ( .A1(n9640), .A2(n8451), .ZN(n8291) );
  INV_X1 U7084 ( .A(n8451), .ZN(n8692) );
  NAND2_X1 U7085 ( .A1(n5542), .A2(n8295), .ZN(n8672) );
  INV_X1 U7086 ( .A(n8305), .ZN(n5543) );
  OR2_X2 U7087 ( .A1(n8662), .A2(n8644), .ZN(n8402) );
  INV_X1 U7088 ( .A(n8402), .ZN(n5545) );
  NAND2_X1 U7089 ( .A1(n8662), .A2(n8644), .ZN(n8299) );
  INV_X1 U7090 ( .A(n8668), .ZN(n5544) );
  AND2_X1 U7091 ( .A1(n8297), .A2(n5547), .ZN(n5546) );
  NAND2_X1 U7092 ( .A1(n7935), .A2(n5546), .ZN(n5549) );
  NAND2_X1 U7093 ( .A1(n5547), .A2(n4367), .ZN(n5548) );
  INV_X1 U7094 ( .A(n8320), .ZN(n5550) );
  INV_X1 U7095 ( .A(n8326), .ZN(n5551) );
  NAND2_X1 U7096 ( .A1(n8601), .A2(n8334), .ZN(n5552) );
  NAND2_X1 U7097 ( .A1(n5552), .A2(n8327), .ZN(n8592) );
  NAND2_X1 U7098 ( .A1(n8780), .A2(n8585), .ZN(n8375) );
  INV_X1 U7099 ( .A(n5553), .ZN(n5554) );
  OAI21_X1 U7100 ( .B1(n8580), .B2(n5554), .A(n8337), .ZN(n8569) );
  INV_X1 U7101 ( .A(n8341), .ZN(n5555) );
  OR2_X1 U7102 ( .A1(n8358), .A2(n5556), .ZN(n5557) );
  NAND2_X1 U7103 ( .A1(n5559), .A2(n8412), .ZN(n6228) );
  INV_X1 U7104 ( .A(n8439), .ZN(n7590) );
  NAND2_X1 U7105 ( .A1(n7590), .A2(n6975), .ZN(n10079) );
  NAND2_X1 U7106 ( .A1(n5559), .A2(n8439), .ZN(n6231) );
  NAND2_X1 U7107 ( .A1(n6228), .A2(n6231), .ZN(n5560) );
  XNOR2_X1 U7108 ( .A(n5561), .B(n8434), .ZN(n7204) );
  INV_X1 U7109 ( .A(n7204), .ZN(n7080) );
  INV_X1 U7110 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n9399) );
  NAND2_X1 U7111 ( .A1(n5513), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7112 ( .A1(n8367), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5563) );
  OAI211_X1 U7113 ( .C1(n5565), .C2(n9399), .A(n5564), .B(n5563), .ZN(n5566)
         );
  INV_X1 U7114 ( .A(n5566), .ZN(n5567) );
  NAND2_X1 U7115 ( .A1(n8373), .A2(n5567), .ZN(n8442) );
  NAND2_X1 U7116 ( .A1(n6242), .A2(P2_B_REG_SCAN_IN), .ZN(n5568) );
  AND2_X1 U7117 ( .A1(n8653), .A2(n5568), .ZN(n8538) );
  AOI22_X1 U7118 ( .A1(n8655), .A2(n8443), .B1(n8442), .B2(n8538), .ZN(n5569)
         );
  NOR2_X1 U7119 ( .A1(n8552), .A2(n10069), .ZN(n5574) );
  NAND2_X1 U7120 ( .A1(n5583), .A2(n5575), .ZN(n5577) );
  NAND2_X1 U7121 ( .A1(n5576), .A2(n5577), .ZN(n5590) );
  XNOR2_X1 U7122 ( .A(n5590), .B(P2_B_REG_SCAN_IN), .ZN(n5580) );
  NAND2_X1 U7123 ( .A1(n5580), .A2(n5604), .ZN(n5587) );
  NAND2_X1 U7124 ( .A1(n5581), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U7125 ( .A1(n5583), .A2(n5582), .ZN(n5584) );
  NAND2_X1 U7126 ( .A1(n5584), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n5585) );
  INV_X1 U7127 ( .A(n5592), .ZN(n5589) );
  INV_X1 U7128 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7129 ( .A1(n7795), .A2(n5590), .ZN(n6826) );
  NOR2_X1 U7130 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .ZN(
        n5596) );
  NOR4_X1 U7131 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n5595) );
  NOR4_X1 U7132 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5594) );
  NOR4_X1 U7133 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n5593) );
  NAND4_X1 U7134 ( .A1(n5596), .A2(n5595), .A3(n5594), .A4(n5593), .ZN(n5602)
         );
  NOR4_X1 U7135 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5600) );
  NOR4_X1 U7136 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5599) );
  NOR4_X1 U7137 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5598) );
  NOR4_X1 U7138 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5597) );
  NAND4_X1 U7139 ( .A1(n5600), .A2(n5599), .A3(n5598), .A4(n5597), .ZN(n5601)
         );
  NOR2_X1 U7140 ( .A1(n5602), .A2(n5601), .ZN(n5603) );
  INV_X1 U7141 ( .A(n6229), .ZN(n7001) );
  NOR2_X1 U7142 ( .A1(n6977), .A2(n7001), .ZN(n5607) );
  OR2_X1 U7143 ( .A1(n5592), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7144 ( .A1(n4310), .A2(n7795), .ZN(n5605) );
  INV_X1 U7145 ( .A(n6924), .ZN(n6235) );
  NAND2_X1 U7146 ( .A1(n4344), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5609) );
  XNOR2_X1 U7147 ( .A(n5609), .B(n5608), .ZN(n7012) );
  OR2_X1 U7148 ( .A1(n5610), .A2(n8412), .ZN(n5613) );
  NOR2_X1 U7149 ( .A1(n4275), .A2(n10066), .ZN(n5611) );
  NAND2_X1 U7150 ( .A1(n5613), .A2(n5611), .ZN(n6992) );
  NAND2_X1 U7151 ( .A1(n6973), .A2(n10066), .ZN(n8588) );
  NAND2_X1 U7152 ( .A1(n6992), .A2(n8588), .ZN(n7000) );
  NAND2_X1 U7153 ( .A1(n7013), .A2(n7000), .ZN(n5617) );
  NAND2_X1 U7154 ( .A1(n6977), .A2(n6924), .ZN(n7002) );
  NAND2_X1 U7155 ( .A1(n6229), .A2(n8437), .ZN(n5612) );
  NOR2_X1 U7156 ( .A1(n7002), .A2(n5612), .ZN(n7016) );
  INV_X1 U7157 ( .A(n5613), .ZN(n5614) );
  NAND2_X1 U7158 ( .A1(n5614), .A2(n6975), .ZN(n7005) );
  NAND2_X1 U7159 ( .A1(n7005), .A2(n7007), .ZN(n5615) );
  NAND2_X1 U7160 ( .A1(n7016), .A2(n5615), .ZN(n5616) );
  NOR2_X1 U7161 ( .A1(n10085), .A2(n9316), .ZN(n5620) );
  OAI21_X1 U7162 ( .B1(n6240), .B2(n10087), .A(n5621), .ZN(P2_U3456) );
  NOR2_X1 U7163 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5626) );
  NOR2_X1 U7164 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5625) );
  NOR2_X1 U7165 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5624) );
  NOR2_X1 U7166 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5623) );
  NAND2_X1 U7167 ( .A1(n6067), .A2(n5640), .ZN(n5642) );
  INV_X1 U7168 ( .A(n5642), .ZN(n5629) );
  NOR2_X1 U7169 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5628) );
  NOR2_X1 U7170 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5627) );
  INV_X1 U7171 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U7172 ( .A1(n7529), .A2(n6500), .ZN(n5636) );
  NAND2_X1 U7173 ( .A1(n6364), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5635) );
  INV_X1 U7174 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5637) );
  XNOR2_X1 U7175 ( .A(n5641), .B(n5640), .ZN(n5647) );
  NAND2_X1 U7176 ( .A1(n5642), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5643) );
  INV_X1 U7177 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U7178 ( .A1(n7232), .A2(n7471), .ZN(n6834) );
  NAND2_X1 U7179 ( .A1(n5645), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5646) );
  XNOR2_X1 U7180 ( .A(n5646), .B(n5631), .ZN(n7587) );
  INV_X1 U7181 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5649) );
  OR2_X1 U7182 ( .A1(n6694), .A2(n7533), .ZN(n7494) );
  NAND2_X1 U7183 ( .A1(n5651), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5652) );
  MUX2_X1 U7184 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5652), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n5655) );
  INV_X1 U7185 ( .A(n5653), .ZN(n5654) );
  INV_X1 U7186 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U7187 ( .A1(n5658), .A2(n5656), .ZN(n5660) );
  NAND2_X1 U7188 ( .A1(n5660), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5657) );
  INV_X1 U7189 ( .A(n5658), .ZN(n5659) );
  NAND2_X1 U7190 ( .A1(n5659), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7191 ( .A1(n7232), .A2(n6704), .ZN(n6832) );
  NAND2_X1 U7192 ( .A1(n7533), .A2(n6832), .ZN(n5662) );
  NAND2_X1 U7193 ( .A1(n6840), .A2(n5662), .ZN(n5663) );
  NAND2_X1 U7194 ( .A1(n5663), .A2(n6731), .ZN(n5693) );
  NAND2_X1 U7195 ( .A1(n9551), .A2(n5769), .ZN(n5680) );
  NAND2_X1 U7196 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5664) );
  NAND2_X1 U7197 ( .A1(n5665), .A2(n5664), .ZN(n5666) );
  XNOR2_X2 U7198 ( .A(n5666), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5672) );
  NOR2_X1 U7199 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n5667) );
  NAND2_X1 U7200 ( .A1(n5668), .A2(n5667), .ZN(n9586) );
  INV_X1 U7201 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U7202 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5782) );
  NAND2_X1 U7203 ( .A1(n5809), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5831) );
  NAND2_X1 U7204 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n5670) );
  NAND2_X1 U7205 ( .A1(n5918), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5942) );
  INV_X1 U7206 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6881) );
  INV_X1 U7207 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5960) );
  NAND2_X1 U7208 ( .A1(n5990), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6012) );
  INV_X1 U7209 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6011) );
  INV_X1 U7210 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6029) );
  INV_X1 U7211 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8852) );
  INV_X1 U7212 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9387) );
  OR2_X1 U7213 ( .A1(n6110), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U7214 ( .A1(n6110), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7215 ( .A1(n5671), .A2(n6128), .ZN(n9289) );
  NAND2_X4 U7216 ( .A1(n5674), .A2(n5675), .ZN(n6412) );
  OR2_X1 U7217 ( .A1(n9289), .A2(n6412), .ZN(n5677) );
  NAND2_X4 U7218 ( .A1(n5674), .A2(n7920), .ZN(n6509) );
  AOI22_X1 U7219 ( .A1(n6161), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n4272), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n5676) );
  OAI211_X1 U7220 ( .C1(n4268), .C2(n5678), .A(n5677), .B(n5676), .ZN(n9121)
         );
  NAND2_X1 U7221 ( .A1(n9121), .A2(n6422), .ZN(n5679) );
  NAND2_X1 U7222 ( .A1(n5680), .A2(n5679), .ZN(n5681) );
  XNOR2_X1 U7223 ( .A(n5681), .B(n6394), .ZN(n6122) );
  INV_X1 U7224 ( .A(n6122), .ZN(n6124) );
  INV_X2 U7225 ( .A(n5688), .ZN(n6422) );
  AOI22_X1 U7226 ( .A1(n9551), .A2(n6422), .B1(n6421), .B2(n9121), .ZN(n6123)
         );
  NAND2_X1 U7227 ( .A1(n6111), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5686) );
  INV_X1 U7228 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5683) );
  OR2_X1 U7229 ( .A1(n6509), .A2(n5683), .ZN(n5685) );
  NAND2_X1 U7230 ( .A1(n4273), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5684) );
  NAND4_X1 U7231 ( .A1(n5687), .A2(n5686), .A3(n5685), .A4(n5684), .ZN(n6449)
         );
  NAND2_X1 U7232 ( .A1(n6449), .A2(n6100), .ZN(n5692) );
  INV_X1 U7233 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5690) );
  NAND2_X1 U7234 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5689) );
  XNOR2_X1 U7235 ( .A(n5690), .B(n5689), .ZN(n6790) );
  INV_X1 U7236 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6733) );
  INV_X1 U7237 ( .A(n5698), .ZN(n5696) );
  AOI22_X1 U7238 ( .A1(n8973), .A2(n6421), .B1(n6100), .B2(n4314), .ZN(n5697)
         );
  INV_X1 U7239 ( .A(n5697), .ZN(n5695) );
  NAND2_X1 U7240 ( .A1(n5696), .A2(n5695), .ZN(n5699) );
  INV_X1 U7241 ( .A(n6862), .ZN(n5717) );
  INV_X1 U7242 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6762) );
  INV_X1 U7243 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7244 ( .A1(n6111), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5703) );
  INV_X1 U7245 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5701) );
  AND3_X1 U7246 ( .A1(n5704), .A2(n5703), .A3(n5702), .ZN(n5706) );
  INV_X1 U7247 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7340) );
  NAND2_X1 U7248 ( .A1(n6735), .A2(SI_0_), .ZN(n5708) );
  XNOR2_X1 U7249 ( .A(n5708), .B(n5707), .ZN(n9592) );
  MUX2_X1 U7250 ( .A(n6762), .B(n9592), .S(n6755), .Z(n7523) );
  INV_X1 U7251 ( .A(n7523), .ZN(n7330) );
  NAND2_X1 U7252 ( .A1(n7330), .A2(n6100), .ZN(n5709) );
  NAND2_X1 U7253 ( .A1(n8975), .A2(n6100), .ZN(n5713) );
  INV_X1 U7254 ( .A(n6731), .ZN(n5711) );
  NAND2_X1 U7255 ( .A1(n5711), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5712) );
  OAI211_X1 U7256 ( .C1(n5959), .C2(n7523), .A(n5713), .B(n5712), .ZN(n6853)
         );
  NAND2_X1 U7257 ( .A1(n6852), .A2(n6853), .ZN(n5715) );
  NAND2_X1 U7258 ( .A1(n7523), .A2(n6173), .ZN(n5714) );
  NAND2_X1 U7259 ( .A1(n5715), .A2(n5714), .ZN(n6861) );
  INV_X1 U7260 ( .A(n6861), .ZN(n5716) );
  NAND2_X1 U7261 ( .A1(n5717), .A2(n5716), .ZN(n6863) );
  NAND2_X1 U7262 ( .A1(n6863), .A2(n6897), .ZN(n5737) );
  NAND2_X1 U7263 ( .A1(n4272), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5724) );
  INV_X1 U7264 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9878) );
  OR2_X1 U7265 ( .A1(n6412), .A2(n9878), .ZN(n5723) );
  INV_X1 U7266 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5719) );
  OR2_X1 U7267 ( .A1(n6505), .A2(n5719), .ZN(n5722) );
  INV_X1 U7268 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5720) );
  OR2_X1 U7269 ( .A1(n6509), .A2(n5720), .ZN(n5721) );
  NAND2_X1 U7270 ( .A1(n8972), .A2(n6100), .ZN(n5730) );
  INV_X1 U7271 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5745) );
  OR2_X1 U7272 ( .A1(n4312), .A2(n6746), .ZN(n5728) );
  INV_X1 U7273 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6732) );
  OR2_X1 U7274 ( .A1(n4274), .A2(n6732), .ZN(n5727) );
  OAI211_X1 U7275 ( .C1(n6755), .C2(n6789), .A(n5728), .B(n5727), .ZN(n7278)
         );
  NAND2_X1 U7276 ( .A1(n4269), .A2(n5769), .ZN(n5729) );
  NAND2_X1 U7277 ( .A1(n5730), .A2(n5729), .ZN(n5731) );
  INV_X1 U7278 ( .A(n5735), .ZN(n5733) );
  AOI22_X1 U7279 ( .A1(n8972), .A2(n6421), .B1(n6100), .B2(n4269), .ZN(n5734)
         );
  INV_X1 U7280 ( .A(n5734), .ZN(n5732) );
  NAND2_X1 U7281 ( .A1(n5733), .A2(n5732), .ZN(n5736) );
  NAND2_X1 U7282 ( .A1(n5735), .A2(n5734), .ZN(n5738) );
  AND2_X1 U7283 ( .A1(n5736), .A2(n5738), .ZN(n6898) );
  NAND2_X1 U7284 ( .A1(n5737), .A2(n6898), .ZN(n6901) );
  NAND2_X1 U7285 ( .A1(n4272), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5744) );
  OR2_X1 U7286 ( .A1(n6412), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5743) );
  INV_X1 U7287 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5739) );
  OR2_X1 U7288 ( .A1(n4268), .A2(n5739), .ZN(n5742) );
  INV_X1 U7289 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5740) );
  OR2_X1 U7290 ( .A1(n6509), .A2(n5740), .ZN(n5741) );
  NAND2_X1 U7291 ( .A1(n8971), .A2(n6422), .ZN(n5752) );
  NAND2_X1 U7292 ( .A1(n5762), .A2(n5745), .ZN(n5746) );
  NAND2_X1 U7293 ( .A1(n5746), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5748) );
  INV_X1 U7294 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5747) );
  XNOR2_X1 U7295 ( .A(n5748), .B(n5747), .ZN(n6793) );
  OR2_X1 U7296 ( .A1(n5888), .A2(n6737), .ZN(n5750) );
  INV_X1 U7297 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6734) );
  OR2_X1 U7298 ( .A1(n4274), .A2(n6734), .ZN(n5749) );
  OAI211_X1 U7299 ( .C1(n6755), .C2(n6793), .A(n5750), .B(n5749), .ZN(n9919)
         );
  NAND2_X1 U7300 ( .A1(n4271), .A2(n5769), .ZN(n5751) );
  NAND2_X1 U7301 ( .A1(n5752), .A2(n5751), .ZN(n5753) );
  XNOR2_X1 U7302 ( .A(n5753), .B(n6394), .ZN(n5773) );
  AOI22_X1 U7303 ( .A1(n8971), .A2(n6421), .B1(n6422), .B2(n4271), .ZN(n5774)
         );
  XNOR2_X1 U7304 ( .A(n5773), .B(n5774), .ZN(n8841) );
  NAND2_X1 U7305 ( .A1(n6111), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5759) );
  INV_X1 U7306 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5754) );
  OR2_X1 U7307 ( .A1(n5781), .A2(n5754), .ZN(n5758) );
  OAI21_X1 U7308 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5782), .ZN(n9863) );
  OR2_X1 U7309 ( .A1(n6412), .A2(n9863), .ZN(n5757) );
  INV_X1 U7310 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5755) );
  OR2_X1 U7311 ( .A1(n6509), .A2(n5755), .ZN(n5756) );
  NAND4_X1 U7312 ( .A1(n5759), .A2(n5758), .A3(n5757), .A4(n5756), .ZN(n8970)
         );
  NAND2_X1 U7313 ( .A1(n8970), .A2(n6100), .ZN(n5771) );
  OR2_X1 U7314 ( .A1(n5760), .A2(n5892), .ZN(n5761) );
  INV_X1 U7315 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U7316 ( .A1(n5764), .A2(n5763), .ZN(n5789) );
  INV_X1 U7317 ( .A(n5764), .ZN(n5765) );
  NAND2_X1 U7318 ( .A1(n5765), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5766) );
  NAND2_X1 U7319 ( .A1(n5789), .A2(n5766), .ZN(n6795) );
  OR2_X1 U7320 ( .A1(n5888), .A2(n6738), .ZN(n5768) );
  INV_X1 U7321 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9416) );
  OR2_X1 U7322 ( .A1(n4274), .A2(n9416), .ZN(n5767) );
  OAI211_X1 U7323 ( .C1(n6755), .C2(n6795), .A(n5768), .B(n5767), .ZN(n7299)
         );
  NAND2_X1 U7324 ( .A1(n7299), .A2(n5769), .ZN(n5770) );
  NAND2_X1 U7325 ( .A1(n5771), .A2(n5770), .ZN(n5772) );
  XNOR2_X1 U7326 ( .A(n5772), .B(n6394), .ZN(n5779) );
  AOI22_X1 U7327 ( .A1(n8970), .A2(n6421), .B1(n6422), .B2(n7299), .ZN(n5777)
         );
  XNOR2_X1 U7328 ( .A(n5779), .B(n5777), .ZN(n7027) );
  INV_X1 U7329 ( .A(n5773), .ZN(n5775) );
  NAND2_X1 U7330 ( .A1(n5775), .A2(n5774), .ZN(n7025) );
  AND2_X1 U7331 ( .A1(n7027), .A2(n7025), .ZN(n5776) );
  INV_X1 U7332 ( .A(n5777), .ZN(n5778) );
  NAND2_X1 U7333 ( .A1(n5779), .A2(n5778), .ZN(n5780) );
  NAND2_X1 U7334 ( .A1(n6161), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5788) );
  INV_X1 U7335 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7298) );
  OR2_X1 U7336 ( .A1(n5781), .A2(n7298), .ZN(n5787) );
  AND2_X1 U7337 ( .A1(n5782), .A2(n7168), .ZN(n5783) );
  OR2_X1 U7338 ( .A1(n5783), .A2(n5809), .ZN(n7302) );
  OR2_X1 U7339 ( .A1(n6412), .A2(n7302), .ZN(n5786) );
  INV_X1 U7340 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5784) );
  OR2_X1 U7341 ( .A1(n4268), .A2(n5784), .ZN(n5785) );
  NAND2_X1 U7342 ( .A1(n8969), .A2(n6422), .ZN(n5794) );
  NAND2_X1 U7343 ( .A1(n6364), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U7344 ( .A1(n5789), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5790) );
  XNOR2_X1 U7345 ( .A(n5790), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6797) );
  NAND2_X1 U7346 ( .A1(n6087), .A2(n6797), .ZN(n5791) );
  NAND2_X1 U7347 ( .A1(n9932), .A2(n5769), .ZN(n5793) );
  NAND2_X1 U7348 ( .A1(n5794), .A2(n5793), .ZN(n5795) );
  XNOR2_X1 U7349 ( .A(n5795), .B(n6394), .ZN(n5798) );
  NAND2_X1 U7350 ( .A1(n8969), .A2(n6421), .ZN(n5797) );
  NAND2_X1 U7351 ( .A1(n9932), .A2(n6422), .ZN(n5796) );
  NAND2_X1 U7352 ( .A1(n5797), .A2(n5796), .ZN(n7167) );
  NAND2_X1 U7353 ( .A1(n7164), .A2(n7167), .ZN(n5800) );
  NAND2_X1 U7354 ( .A1(n5799), .A2(n5798), .ZN(n7165) );
  OR2_X1 U7355 ( .A1(n6744), .A2(n5888), .ZN(n5807) );
  NAND2_X1 U7356 ( .A1(n5801), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5802) );
  MUX2_X1 U7357 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5802), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5805) );
  AND2_X1 U7358 ( .A1(n5805), .A2(n5804), .ZN(n6801) );
  AOI22_X1 U7359 ( .A1(n6364), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6087), .B2(
        n6801), .ZN(n5806) );
  NAND2_X1 U7360 ( .A1(n5807), .A2(n5806), .ZN(n7324) );
  NAND2_X1 U7361 ( .A1(n7324), .A2(n5769), .ZN(n5817) );
  NAND2_X1 U7362 ( .A1(n6161), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5815) );
  INV_X1 U7363 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5808) );
  OR2_X1 U7364 ( .A1(n5781), .A2(n5808), .ZN(n5814) );
  OR2_X1 U7365 ( .A1(n5809), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U7366 ( .A1(n5831), .A2(n5810), .ZN(n7259) );
  OR2_X1 U7367 ( .A1(n6412), .A2(n7259), .ZN(n5813) );
  INV_X1 U7368 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5811) );
  OR2_X1 U7369 ( .A1(n4268), .A2(n5811), .ZN(n5812) );
  NAND4_X1 U7370 ( .A1(n5815), .A2(n5814), .A3(n5813), .A4(n5812), .ZN(n8968)
         );
  NAND2_X1 U7371 ( .A1(n8968), .A2(n6422), .ZN(n5816) );
  NAND2_X1 U7372 ( .A1(n5817), .A2(n5816), .ZN(n5818) );
  XNOR2_X1 U7373 ( .A(n5818), .B(n6173), .ZN(n5821) );
  NAND2_X1 U7374 ( .A1(n7324), .A2(n6422), .ZN(n5820) );
  NAND2_X1 U7375 ( .A1(n8968), .A2(n6421), .ZN(n5819) );
  AND2_X1 U7376 ( .A1(n5820), .A2(n5819), .ZN(n5822) );
  NAND2_X1 U7377 ( .A1(n5821), .A2(n5822), .ZN(n5826) );
  INV_X1 U7378 ( .A(n5821), .ZN(n5824) );
  INV_X1 U7379 ( .A(n5822), .ZN(n5823) );
  NAND2_X1 U7380 ( .A1(n5824), .A2(n5823), .ZN(n5825) );
  NAND2_X1 U7381 ( .A1(n5826), .A2(n5825), .ZN(n7256) );
  OR2_X1 U7382 ( .A1(n6750), .A2(n5888), .ZN(n5829) );
  NAND2_X1 U7383 ( .A1(n5804), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5827) );
  XNOR2_X1 U7384 ( .A(n5827), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6803) );
  AOI22_X1 U7385 ( .A1(n6364), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6087), .B2(
        n6803), .ZN(n5828) );
  NAND2_X1 U7386 ( .A1(n5829), .A2(n5828), .ZN(n7455) );
  NAND2_X1 U7387 ( .A1(n7455), .A2(n5769), .ZN(n5839) );
  NAND2_X1 U7388 ( .A1(n6161), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5837) );
  INV_X1 U7389 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5830) );
  OR2_X1 U7390 ( .A1(n5781), .A2(n5830), .ZN(n5836) );
  NAND2_X1 U7391 ( .A1(n5831), .A2(n7450), .ZN(n5832) );
  NAND2_X1 U7392 ( .A1(n5870), .A2(n5832), .ZN(n7452) );
  OR2_X1 U7393 ( .A1(n6412), .A2(n7452), .ZN(n5835) );
  INV_X1 U7394 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5833) );
  OR2_X1 U7395 ( .A1(n4268), .A2(n5833), .ZN(n5834) );
  NAND4_X1 U7396 ( .A1(n5837), .A2(n5836), .A3(n5835), .A4(n5834), .ZN(n8967)
         );
  NAND2_X1 U7397 ( .A1(n8967), .A2(n6100), .ZN(n5838) );
  NAND2_X1 U7398 ( .A1(n5839), .A2(n5838), .ZN(n5840) );
  XNOR2_X1 U7399 ( .A(n5840), .B(n6173), .ZN(n5842) );
  AND2_X1 U7400 ( .A1(n8967), .A2(n6421), .ZN(n5841) );
  AOI21_X1 U7401 ( .B1(n7455), .B2(n6422), .A(n5841), .ZN(n5843) );
  NAND2_X1 U7402 ( .A1(n5842), .A2(n5843), .ZN(n7447) );
  INV_X1 U7403 ( .A(n5842), .ZN(n5845) );
  INV_X1 U7404 ( .A(n5843), .ZN(n5844) );
  NAND2_X1 U7405 ( .A1(n5845), .A2(n5844), .ZN(n7448) );
  NAND2_X1 U7406 ( .A1(n5846), .A2(n7448), .ZN(n7646) );
  NAND2_X1 U7407 ( .A1(n6757), .A2(n6500), .ZN(n5852) );
  NOR2_X1 U7408 ( .A1(n5804), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5890) );
  OR2_X1 U7409 ( .A1(n5890), .A2(n5892), .ZN(n5849) );
  INV_X1 U7410 ( .A(n5849), .ZN(n5847) );
  NAND2_X1 U7411 ( .A1(n5847), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5850) );
  INV_X1 U7412 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5848) );
  NAND2_X1 U7413 ( .A1(n5849), .A2(n5848), .ZN(n5864) );
  AOI22_X1 U7414 ( .A1(n6364), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6087), .B2(
        n6806), .ZN(n5851) );
  NAND2_X1 U7415 ( .A1(n5852), .A2(n5851), .ZN(n9836) );
  NAND2_X1 U7416 ( .A1(n9836), .A2(n5769), .ZN(n5860) );
  NAND2_X1 U7417 ( .A1(n4273), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5858) );
  INV_X1 U7418 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5853) );
  OR2_X1 U7419 ( .A1(n6509), .A2(n5853), .ZN(n5857) );
  INV_X1 U7420 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7654) );
  XNOR2_X1 U7421 ( .A(n5870), .B(n7654), .ZN(n7651) );
  OR2_X1 U7422 ( .A1(n6412), .A2(n7651), .ZN(n5856) );
  INV_X1 U7423 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5854) );
  OR2_X1 U7424 ( .A1(n4268), .A2(n5854), .ZN(n5855) );
  NAND4_X1 U7425 ( .A1(n5858), .A2(n5857), .A3(n5856), .A4(n5855), .ZN(n8966)
         );
  NAND2_X1 U7426 ( .A1(n8966), .A2(n6100), .ZN(n5859) );
  NAND2_X1 U7427 ( .A1(n5860), .A2(n5859), .ZN(n5861) );
  XNOR2_X1 U7428 ( .A(n5861), .B(n6394), .ZN(n7668) );
  INV_X1 U7429 ( .A(n7668), .ZN(n7647) );
  NAND2_X1 U7430 ( .A1(n9836), .A2(n6100), .ZN(n5863) );
  NAND2_X1 U7431 ( .A1(n8966), .A2(n6421), .ZN(n5862) );
  NAND2_X1 U7432 ( .A1(n5863), .A2(n5862), .ZN(n5881) );
  INV_X1 U7433 ( .A(n5881), .ZN(n7649) );
  NAND2_X1 U7434 ( .A1(n6767), .A2(n6500), .ZN(n5867) );
  NAND2_X1 U7435 ( .A1(n5864), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5865) );
  XNOR2_X1 U7436 ( .A(n5865), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6876) );
  AOI22_X1 U7437 ( .A1(n6364), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6087), .B2(
        n6876), .ZN(n5866) );
  NAND2_X1 U7438 ( .A1(n7680), .A2(n5769), .ZN(n5877) );
  NAND2_X1 U7439 ( .A1(n6111), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5875) );
  INV_X1 U7440 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5868) );
  OR2_X1 U7441 ( .A1(n6509), .A2(n5868), .ZN(n5874) );
  INV_X1 U7442 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7571) );
  OR2_X1 U7443 ( .A1(n5781), .A2(n7571), .ZN(n5873) );
  INV_X1 U7444 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5869) );
  OAI21_X1 U7445 ( .B1(n5870), .B2(n7654), .A(n5869), .ZN(n5871) );
  NAND2_X1 U7446 ( .A1(n5871), .A2(n5901), .ZN(n7678) );
  OR2_X1 U7447 ( .A1(n6412), .A2(n7678), .ZN(n5872) );
  NAND4_X1 U7448 ( .A1(n5875), .A2(n5874), .A3(n5873), .A4(n5872), .ZN(n8965)
         );
  NAND2_X1 U7449 ( .A1(n8965), .A2(n6100), .ZN(n5876) );
  NAND2_X1 U7450 ( .A1(n5877), .A2(n5876), .ZN(n5878) );
  XNOR2_X1 U7451 ( .A(n5878), .B(n6173), .ZN(n5884) );
  INV_X1 U7452 ( .A(n5884), .ZN(n7671) );
  NAND2_X1 U7453 ( .A1(n7680), .A2(n6100), .ZN(n5880) );
  NAND2_X1 U7454 ( .A1(n8965), .A2(n6421), .ZN(n5879) );
  NAND2_X1 U7455 ( .A1(n5880), .A2(n5879), .ZN(n7670) );
  NAND2_X1 U7456 ( .A1(n7671), .A2(n7670), .ZN(n7669) );
  OAI21_X1 U7457 ( .B1(n7647), .B2(n7649), .A(n7669), .ZN(n5886) );
  OAI21_X1 U7458 ( .B1(n7668), .B2(n5881), .A(n7670), .ZN(n5883) );
  NOR2_X1 U7459 ( .A1(n7670), .A2(n5881), .ZN(n5882) );
  AOI22_X1 U7460 ( .A1(n5884), .A2(n5883), .B1(n5882), .B2(n7647), .ZN(n5885)
         );
  OAI21_X1 U7461 ( .B1(n7646), .B2(n5886), .A(n5885), .ZN(n5887) );
  OR2_X1 U7462 ( .A1(n6774), .A2(n5888), .ZN(n5899) );
  NOR2_X1 U7463 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5889) );
  AND2_X1 U7464 ( .A1(n5890), .A2(n5889), .ZN(n5895) );
  NOR2_X1 U7465 ( .A1(n5895), .A2(n5892), .ZN(n5891) );
  MUX2_X1 U7466 ( .A(n5892), .B(n5891), .S(P1_IR_REG_10__SCAN_IN), .Z(n5893)
         );
  INV_X1 U7467 ( .A(n5893), .ZN(n5897) );
  INV_X1 U7468 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5894) );
  INV_X1 U7469 ( .A(n5937), .ZN(n5896) );
  AOI22_X1 U7470 ( .A1(n6364), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6087), .B2(
        n9602), .ZN(n5898) );
  NAND2_X1 U7471 ( .A1(n7512), .A2(n5769), .ZN(n5909) );
  NAND2_X1 U7472 ( .A1(n6111), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5907) );
  INV_X1 U7473 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7507) );
  OR2_X1 U7474 ( .A1(n5781), .A2(n7507), .ZN(n5906) );
  INV_X1 U7475 ( .A(n5918), .ZN(n5903) );
  NAND2_X1 U7476 ( .A1(n5901), .A2(n5900), .ZN(n5902) );
  NAND2_X1 U7477 ( .A1(n5903), .A2(n5902), .ZN(n7758) );
  OR2_X1 U7478 ( .A1(n6412), .A2(n7758), .ZN(n5905) );
  INV_X1 U7479 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6874) );
  OR2_X1 U7480 ( .A1(n6509), .A2(n6874), .ZN(n5904) );
  NAND4_X1 U7481 ( .A1(n5907), .A2(n5906), .A3(n5905), .A4(n5904), .ZN(n8964)
         );
  NAND2_X1 U7482 ( .A1(n8964), .A2(n6100), .ZN(n5908) );
  NAND2_X1 U7483 ( .A1(n5909), .A2(n5908), .ZN(n5910) );
  XNOR2_X1 U7484 ( .A(n5910), .B(n6173), .ZN(n5933) );
  NAND2_X1 U7485 ( .A1(n7512), .A2(n6100), .ZN(n5912) );
  NAND2_X1 U7486 ( .A1(n8964), .A2(n6421), .ZN(n5911) );
  AND2_X1 U7487 ( .A1(n5933), .A2(n7756), .ZN(n5913) );
  INV_X1 U7488 ( .A(n5913), .ZN(n5914) );
  NAND2_X1 U7489 ( .A1(n6816), .A2(n6500), .ZN(n5917) );
  OR2_X1 U7490 ( .A1(n5937), .A2(n5892), .ZN(n5915) );
  XNOR2_X1 U7491 ( .A(n5915), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9728) );
  AOI22_X1 U7492 ( .A1(n6364), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6087), .B2(
        n9728), .ZN(n5916) );
  NAND2_X1 U7493 ( .A1(n7853), .A2(n5769), .ZN(n5925) );
  NAND2_X1 U7494 ( .A1(n6111), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5923) );
  INV_X1 U7495 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7496) );
  OR2_X1 U7496 ( .A1(n5781), .A2(n7496), .ZN(n5922) );
  INV_X1 U7497 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6877) );
  OR2_X1 U7498 ( .A1(n6509), .A2(n6877), .ZN(n5921) );
  OR2_X1 U7499 ( .A1(n5918), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U7500 ( .A1(n5942), .A2(n5919), .ZN(n7844) );
  OR2_X1 U7501 ( .A1(n6412), .A2(n7844), .ZN(n5920) );
  NAND4_X1 U7502 ( .A1(n5923), .A2(n5922), .A3(n5921), .A4(n5920), .ZN(n8963)
         );
  NAND2_X1 U7503 ( .A1(n8963), .A2(n6100), .ZN(n5924) );
  NAND2_X1 U7504 ( .A1(n5925), .A2(n5924), .ZN(n5926) );
  XNOR2_X1 U7505 ( .A(n5926), .B(n6173), .ZN(n5928) );
  AND2_X1 U7506 ( .A1(n8963), .A2(n6421), .ZN(n5927) );
  AOI21_X1 U7507 ( .B1(n7853), .B2(n6422), .A(n5927), .ZN(n5929) );
  NAND2_X1 U7508 ( .A1(n5928), .A2(n5929), .ZN(n7765) );
  INV_X1 U7509 ( .A(n5928), .ZN(n5931) );
  INV_X1 U7510 ( .A(n5929), .ZN(n5930) );
  NAND2_X1 U7511 ( .A1(n5931), .A2(n5930), .ZN(n5932) );
  NAND2_X1 U7512 ( .A1(n7765), .A2(n5932), .ZN(n7847) );
  INV_X1 U7513 ( .A(n5933), .ZN(n7754) );
  INV_X1 U7514 ( .A(n7756), .ZN(n5934) );
  AND2_X1 U7515 ( .A1(n7754), .A2(n5934), .ZN(n5935) );
  NOR2_X1 U7516 ( .A1(n7847), .A2(n5935), .ZN(n7764) );
  INV_X1 U7517 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U7518 ( .A1(n5937), .A2(n5936), .ZN(n5983) );
  NAND2_X1 U7519 ( .A1(n5983), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5938) );
  INV_X1 U7520 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7521 ( .A1(n5938), .A2(n5981), .ZN(n5955) );
  OR2_X1 U7522 ( .A1(n5938), .A2(n5981), .ZN(n5939) );
  AOI22_X1 U7523 ( .A1(n6364), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6087), .B2(
        n9045), .ZN(n5940) );
  NAND2_X1 U7524 ( .A1(n6463), .A2(n5769), .ZN(n5949) );
  NAND2_X1 U7525 ( .A1(n6111), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5947) );
  INV_X1 U7526 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5941) );
  OR2_X1 U7527 ( .A1(n6509), .A2(n5941), .ZN(n5946) );
  INV_X1 U7528 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7614) );
  OR2_X1 U7529 ( .A1(n5781), .A2(n7614), .ZN(n5945) );
  NAND2_X1 U7530 ( .A1(n5942), .A2(n6881), .ZN(n5943) );
  NAND2_X1 U7531 ( .A1(n5961), .A2(n5943), .ZN(n7772) );
  OR2_X1 U7532 ( .A1(n6412), .A2(n7772), .ZN(n5944) );
  NAND4_X1 U7533 ( .A1(n5947), .A2(n5946), .A3(n5945), .A4(n5944), .ZN(n8962)
         );
  NAND2_X1 U7534 ( .A1(n8962), .A2(n6422), .ZN(n5948) );
  NAND2_X1 U7535 ( .A1(n5949), .A2(n5948), .ZN(n5950) );
  XNOR2_X1 U7536 ( .A(n5950), .B(n6173), .ZN(n5953) );
  AND2_X1 U7537 ( .A1(n8962), .A2(n6421), .ZN(n5951) );
  AOI21_X1 U7538 ( .B1(n6463), .B2(n6422), .A(n5951), .ZN(n5952) );
  NAND2_X1 U7539 ( .A1(n5953), .A2(n5952), .ZN(n5976) );
  NAND2_X1 U7540 ( .A1(n5954), .A2(n5976), .ZN(n5975) );
  AND2_X1 U7541 ( .A1(n7764), .A2(n7766), .ZN(n7729) );
  NAND2_X1 U7542 ( .A1(n5955), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5956) );
  XNOR2_X1 U7543 ( .A(n5956), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9754) );
  AOI22_X1 U7544 ( .A1(n6364), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6087), .B2(
        n9754), .ZN(n5957) );
  NAND2_X1 U7545 ( .A1(n7696), .A2(n5769), .ZN(n5969) );
  NAND2_X1 U7546 ( .A1(n6111), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5967) );
  INV_X1 U7547 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7691) );
  OR2_X1 U7548 ( .A1(n5781), .A2(n7691), .ZN(n5966) );
  INV_X1 U7549 ( .A(n5990), .ZN(n5963) );
  NAND2_X1 U7550 ( .A1(n5961), .A2(n5960), .ZN(n5962) );
  NAND2_X1 U7551 ( .A1(n5963), .A2(n5962), .ZN(n7737) );
  OR2_X1 U7552 ( .A1(n6412), .A2(n7737), .ZN(n5965) );
  INV_X1 U7553 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9033) );
  OR2_X1 U7554 ( .A1(n6509), .A2(n9033), .ZN(n5964) );
  NAND4_X1 U7555 ( .A1(n5967), .A2(n5966), .A3(n5965), .A4(n5964), .ZN(n8961)
         );
  NAND2_X1 U7556 ( .A1(n8961), .A2(n6422), .ZN(n5968) );
  NAND2_X1 U7557 ( .A1(n5969), .A2(n5968), .ZN(n5970) );
  AND2_X1 U7558 ( .A1(n8961), .A2(n6421), .ZN(n5971) );
  AOI21_X1 U7559 ( .B1(n7696), .B2(n6422), .A(n5971), .ZN(n5973) );
  INV_X1 U7560 ( .A(n5972), .ZN(n5974) );
  NAND2_X1 U7561 ( .A1(n5974), .A2(n5973), .ZN(n5978) );
  INV_X1 U7562 ( .A(n7735), .ZN(n5977) );
  OR2_X1 U7563 ( .A1(n5975), .A2(n7765), .ZN(n7769) );
  AND2_X1 U7564 ( .A1(n7769), .A2(n5976), .ZN(n7730) );
  OR2_X1 U7565 ( .A1(n5977), .A2(n7730), .ZN(n7731) );
  AND2_X1 U7566 ( .A1(n5978), .A2(n7731), .ZN(n5979) );
  INV_X1 U7567 ( .A(n6004), .ZN(n6000) );
  INV_X1 U7568 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U7569 ( .A1(n5981), .A2(n5980), .ZN(n5982) );
  OAI21_X1 U7570 ( .B1(n5983), .B2(n5982), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5984) );
  MUX2_X1 U7571 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5984), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5986) );
  INV_X1 U7572 ( .A(n5985), .ZN(n6006) );
  AND2_X1 U7573 ( .A1(n5986), .A2(n6006), .ZN(n9758) );
  AOI22_X1 U7574 ( .A1(n6364), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6087), .B2(
        n9758), .ZN(n5987) );
  NAND2_X1 U7575 ( .A1(n9817), .A2(n5769), .ZN(n5997) );
  NAND2_X1 U7576 ( .A1(n4273), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5995) );
  INV_X1 U7577 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5989) );
  OR2_X1 U7578 ( .A1(n4268), .A2(n5989), .ZN(n5994) );
  OR2_X1 U7579 ( .A1(n5990), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7580 ( .A1(n6012), .A2(n5991), .ZN(n9815) );
  OR2_X1 U7581 ( .A1(n6412), .A2(n9815), .ZN(n5993) );
  INV_X1 U7582 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9035) );
  OR2_X1 U7583 ( .A1(n6509), .A2(n9035), .ZN(n5992) );
  NAND4_X1 U7584 ( .A1(n5995), .A2(n5994), .A3(n5993), .A4(n5992), .ZN(n8960)
         );
  NAND2_X1 U7585 ( .A1(n8960), .A2(n6100), .ZN(n5996) );
  NAND2_X1 U7586 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  XNOR2_X1 U7587 ( .A(n5998), .B(n6173), .ZN(n6003) );
  INV_X1 U7588 ( .A(n6003), .ZN(n5999) );
  NAND2_X1 U7589 ( .A1(n6000), .A2(n5999), .ZN(n7815) );
  NAND2_X1 U7590 ( .A1(n9817), .A2(n6422), .ZN(n6002) );
  NAND2_X1 U7591 ( .A1(n8960), .A2(n6421), .ZN(n6001) );
  NAND2_X1 U7592 ( .A1(n6002), .A2(n6001), .ZN(n7820) );
  INV_X1 U7593 ( .A(n7820), .ZN(n6005) );
  NAND3_X1 U7594 ( .A1(n7815), .A2(n6005), .A3(n7816), .ZN(n7817) );
  NAND2_X1 U7595 ( .A1(n6006), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6007) );
  MUX2_X1 U7596 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6007), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n6008) );
  NAND2_X1 U7597 ( .A1(n6008), .A2(n6024), .ZN(n9048) );
  INV_X1 U7598 ( .A(n9048), .ZN(n9784) );
  AOI22_X1 U7599 ( .A1(n6364), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6087), .B2(
        n9784), .ZN(n6009) );
  NAND2_X1 U7600 ( .A1(n7790), .A2(n5769), .ZN(n6020) );
  NAND2_X1 U7601 ( .A1(n6111), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7602 ( .A1(n6012), .A2(n6011), .ZN(n6013) );
  NAND2_X1 U7603 ( .A1(n6030), .A2(n6013), .ZN(n8943) );
  OR2_X1 U7604 ( .A1(n6412), .A2(n8943), .ZN(n6017) );
  INV_X1 U7605 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7787) );
  OR2_X1 U7606 ( .A1(n5781), .A2(n7787), .ZN(n6016) );
  INV_X1 U7607 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6014) );
  OR2_X1 U7608 ( .A1(n6509), .A2(n6014), .ZN(n6015) );
  NAND4_X1 U7609 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .ZN(n8959)
         );
  NAND2_X1 U7610 ( .A1(n8959), .A2(n6422), .ZN(n6019) );
  NAND2_X1 U7611 ( .A1(n6020), .A2(n6019), .ZN(n6021) );
  XNOR2_X1 U7612 ( .A(n6021), .B(n6394), .ZN(n6022) );
  AOI22_X1 U7613 ( .A1(n7790), .A2(n6422), .B1(n6421), .B2(n8959), .ZN(n8939)
         );
  NAND2_X1 U7614 ( .A1(n6024), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6025) );
  MUX2_X1 U7615 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6025), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n6026) );
  AND2_X1 U7616 ( .A1(n6026), .A2(n6046), .ZN(n9059) );
  AOI22_X1 U7617 ( .A1(n6364), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6087), .B2(
        n9059), .ZN(n6027) );
  INV_X1 U7618 ( .A(n9668), .ZN(n9683) );
  AND2_X1 U7619 ( .A1(n6030), .A2(n6029), .ZN(n6031) );
  OR2_X1 U7620 ( .A1(n6031), .A2(n6050), .ZN(n9675) );
  OR2_X1 U7621 ( .A1(n9675), .A2(n6412), .ZN(n6038) );
  INV_X1 U7622 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n6032) );
  OR2_X1 U7623 ( .A1(n5781), .A2(n6032), .ZN(n6037) );
  INV_X1 U7624 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n6033) );
  OR2_X1 U7625 ( .A1(n4268), .A2(n6033), .ZN(n6036) );
  INV_X1 U7626 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n6034) );
  OR2_X1 U7627 ( .A1(n6509), .A2(n6034), .ZN(n6035) );
  NAND4_X1 U7628 ( .A1(n6038), .A2(n6037), .A3(n6036), .A4(n6035), .ZN(n9111)
         );
  INV_X1 U7629 ( .A(n9111), .ZN(n6469) );
  OAI22_X1 U7630 ( .A1(n9683), .A2(n5688), .B1(n6469), .B2(n6039), .ZN(n6043)
         );
  NAND2_X1 U7631 ( .A1(n9668), .A2(n5769), .ZN(n6041) );
  NAND2_X1 U7632 ( .A1(n9111), .A2(n6100), .ZN(n6040) );
  NAND2_X1 U7633 ( .A1(n6041), .A2(n6040), .ZN(n6042) );
  XNOR2_X1 U7634 ( .A(n6042), .B(n6394), .ZN(n6044) );
  XOR2_X1 U7635 ( .A(n6043), .B(n6044), .Z(n8877) );
  OR2_X1 U7636 ( .A1(n6044), .A2(n6043), .ZN(n6045) );
  NAND2_X1 U7637 ( .A1(n7088), .A2(n6500), .ZN(n6049) );
  NAND2_X1 U7638 ( .A1(n6046), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6047) );
  XNOR2_X1 U7639 ( .A(n6047), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9079) );
  AOI22_X1 U7640 ( .A1(n6364), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6087), .B2(
        n9079), .ZN(n6048) );
  NAND2_X1 U7641 ( .A1(n9502), .A2(n5769), .ZN(n6059) );
  NOR2_X1 U7642 ( .A1(n6050), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6051) );
  OR2_X1 U7643 ( .A1(n6073), .A2(n6051), .ZN(n9496) );
  INV_X1 U7644 ( .A(n9496), .ZN(n6052) );
  NAND2_X1 U7645 ( .A1(n5682), .A2(n6052), .ZN(n6057) );
  INV_X1 U7646 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9497) );
  OR2_X1 U7647 ( .A1(n5781), .A2(n9497), .ZN(n6056) );
  INV_X1 U7648 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n6053) );
  OR2_X1 U7649 ( .A1(n4268), .A2(n6053), .ZN(n6055) );
  INV_X1 U7650 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9060) );
  OR2_X1 U7651 ( .A1(n6509), .A2(n9060), .ZN(n6054) );
  NAND4_X1 U7652 ( .A1(n6057), .A2(n6056), .A3(n6055), .A4(n6054), .ZN(n9112)
         );
  NAND2_X1 U7653 ( .A1(n9112), .A2(n6100), .ZN(n6058) );
  NAND2_X1 U7654 ( .A1(n6059), .A2(n6058), .ZN(n6060) );
  XNOR2_X1 U7655 ( .A(n6060), .B(n6394), .ZN(n6063) );
  NAND2_X1 U7656 ( .A1(n9502), .A2(n6100), .ZN(n6062) );
  NAND2_X1 U7657 ( .A1(n9112), .A2(n6421), .ZN(n6061) );
  NAND2_X1 U7658 ( .A1(n6062), .A2(n6061), .ZN(n6064) );
  NAND2_X1 U7659 ( .A1(n6063), .A2(n6064), .ZN(n8886) );
  INV_X1 U7660 ( .A(n6063), .ZN(n6066) );
  INV_X1 U7661 ( .A(n6064), .ZN(n6065) );
  NAND2_X1 U7662 ( .A1(n6066), .A2(n6065), .ZN(n8888) );
  NAND2_X1 U7663 ( .A1(n8884), .A2(n8888), .ZN(n8916) );
  OR2_X1 U7664 ( .A1(n6068), .A2(n6067), .ZN(n6069) );
  AND2_X1 U7665 ( .A1(n6070), .A2(n6069), .ZN(n9800) );
  AOI22_X1 U7666 ( .A1(n6364), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6087), .B2(
        n9800), .ZN(n6071) );
  NAND2_X1 U7667 ( .A1(n9566), .A2(n5769), .ZN(n6080) );
  OR2_X1 U7668 ( .A1(n6073), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6074) );
  AND2_X1 U7669 ( .A1(n6090), .A2(n6074), .ZN(n9482) );
  NAND2_X1 U7670 ( .A1(n9482), .A2(n5682), .ZN(n6078) );
  NAND2_X1 U7671 ( .A1(n4273), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7672 ( .A1(n6111), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7673 ( .A1(n6161), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6075) );
  NAND4_X1 U7674 ( .A1(n6078), .A2(n6077), .A3(n6076), .A4(n6075), .ZN(n8958)
         );
  NAND2_X1 U7675 ( .A1(n8958), .A2(n6100), .ZN(n6079) );
  NAND2_X1 U7676 ( .A1(n6080), .A2(n6079), .ZN(n6081) );
  XNOR2_X1 U7677 ( .A(n6081), .B(n6394), .ZN(n8914) );
  NAND2_X1 U7678 ( .A1(n9566), .A2(n6422), .ZN(n6083) );
  NAND2_X1 U7679 ( .A1(n8958), .A2(n6421), .ZN(n6082) );
  NAND2_X1 U7680 ( .A1(n6083), .A2(n6082), .ZN(n8913) );
  NAND2_X1 U7681 ( .A1(n8914), .A2(n8913), .ZN(n6086) );
  INV_X1 U7682 ( .A(n8914), .ZN(n6085) );
  INV_X1 U7683 ( .A(n8913), .ZN(n6084) );
  NAND2_X1 U7684 ( .A1(n7231), .A2(n6500), .ZN(n6089) );
  NAND2_X1 U7685 ( .A1(n9561), .A2(n5769), .ZN(n6098) );
  INV_X1 U7686 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U7687 ( .A1(n6090), .A2(n8852), .ZN(n6091) );
  NAND2_X1 U7688 ( .A1(n6108), .A2(n6091), .ZN(n9468) );
  OR2_X1 U7689 ( .A1(n9468), .A2(n6412), .ZN(n6095) );
  INV_X1 U7690 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9461) );
  OR2_X1 U7691 ( .A1(n5781), .A2(n9461), .ZN(n6093) );
  INV_X1 U7692 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9081) );
  OR2_X1 U7693 ( .A1(n6509), .A2(n9081), .ZN(n6092) );
  AND2_X1 U7694 ( .A1(n6093), .A2(n6092), .ZN(n6094) );
  OAI211_X1 U7695 ( .C1(n4268), .C2(n6096), .A(n6095), .B(n6094), .ZN(n9115)
         );
  NAND2_X1 U7696 ( .A1(n9115), .A2(n6422), .ZN(n6097) );
  NAND2_X1 U7697 ( .A1(n6098), .A2(n6097), .ZN(n6099) );
  XNOR2_X1 U7698 ( .A(n6099), .B(n6394), .ZN(n8848) );
  NAND2_X1 U7699 ( .A1(n9561), .A2(n6100), .ZN(n6102) );
  NAND2_X1 U7700 ( .A1(n9115), .A2(n6421), .ZN(n6101) );
  NAND2_X1 U7701 ( .A1(n6102), .A2(n6101), .ZN(n6103) );
  INV_X1 U7702 ( .A(n8848), .ZN(n6104) );
  INV_X1 U7703 ( .A(n6103), .ZN(n8847) );
  NAND2_X1 U7704 ( .A1(n7435), .A2(n6500), .ZN(n6107) );
  NAND2_X1 U7705 ( .A1(n6364), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U7706 ( .A1(n9556), .A2(n5769), .ZN(n6115) );
  AND2_X1 U7707 ( .A1(n6108), .A2(n9387), .ZN(n6109) );
  OR2_X1 U7708 ( .A1(n6110), .A2(n6109), .ZN(n9452) );
  AOI22_X1 U7709 ( .A1(n6161), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n4272), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7710 ( .A1(n6111), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6112) );
  OAI211_X1 U7711 ( .C1(n9452), .C2(n6412), .A(n6113), .B(n6112), .ZN(n9118)
         );
  NAND2_X1 U7712 ( .A1(n9118), .A2(n6422), .ZN(n6114) );
  NAND2_X1 U7713 ( .A1(n6115), .A2(n6114), .ZN(n6116) );
  XNOR2_X1 U7714 ( .A(n6116), .B(n6173), .ZN(n6119) );
  AND2_X1 U7715 ( .A1(n9118), .A2(n6421), .ZN(n6117) );
  AOI21_X1 U7716 ( .B1(n9556), .B2(n6422), .A(n6117), .ZN(n6118) );
  NAND2_X1 U7717 ( .A1(n6119), .A2(n6118), .ZN(n6120) );
  OAI21_X1 U7718 ( .B1(n6119), .B2(n6118), .A(n6120), .ZN(n8898) );
  INV_X1 U7719 ( .A(n6120), .ZN(n6121) );
  XOR2_X1 U7720 ( .A(n6123), .B(n6122), .Z(n8858) );
  NAND2_X1 U7721 ( .A1(n7586), .A2(n6500), .ZN(n6126) );
  OR2_X1 U7722 ( .A1(n4274), .A2(n9413), .ZN(n6125) );
  NAND2_X1 U7723 ( .A1(n4273), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6134) );
  INV_X1 U7724 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n6127) );
  OR2_X1 U7725 ( .A1(n4268), .A2(n6127), .ZN(n6133) );
  OAI21_X1 U7726 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n6129), .A(n6142), .ZN(
        n8907) );
  OR2_X1 U7727 ( .A1(n6412), .A2(n8907), .ZN(n6132) );
  INV_X1 U7728 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n6130) );
  OR2_X1 U7729 ( .A1(n6509), .A2(n6130), .ZN(n6131) );
  NAND4_X1 U7730 ( .A1(n6134), .A2(n6133), .A3(n6132), .A4(n6131), .ZN(n9125)
         );
  AOI22_X1 U7731 ( .A1(n9546), .A2(n5769), .B1(n6422), .B2(n9125), .ZN(n6135)
         );
  XOR2_X1 U7732 ( .A(n6394), .B(n6135), .Z(n6136) );
  AOI22_X1 U7733 ( .A1(n9546), .A2(n6422), .B1(n6421), .B2(n9125), .ZN(n8905)
         );
  INV_X1 U7734 ( .A(n6138), .ZN(n8834) );
  NAND2_X1 U7735 ( .A1(n7699), .A2(n6500), .ZN(n6140) );
  NAND2_X1 U7736 ( .A1(n6364), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7737 ( .A1(n9539), .A2(n5769), .ZN(n6150) );
  NAND2_X1 U7738 ( .A1(n6161), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6148) );
  INV_X1 U7739 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6141) );
  OR2_X1 U7740 ( .A1(n5781), .A2(n6141), .ZN(n6147) );
  OAI21_X1 U7741 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n6143), .A(n6164), .ZN(
        n9255) );
  OR2_X1 U7742 ( .A1(n6412), .A2(n9255), .ZN(n6146) );
  INV_X1 U7743 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n6144) );
  OR2_X1 U7744 ( .A1(n4268), .A2(n6144), .ZN(n6145) );
  NAND4_X1 U7745 ( .A1(n6148), .A2(n6147), .A3(n6146), .A4(n6145), .ZN(n9129)
         );
  NAND2_X1 U7746 ( .A1(n9129), .A2(n6422), .ZN(n6149) );
  NAND2_X1 U7747 ( .A1(n6150), .A2(n6149), .ZN(n6151) );
  XNOR2_X1 U7748 ( .A(n6151), .B(n6173), .ZN(n6153) );
  AND2_X1 U7749 ( .A1(n9129), .A2(n6421), .ZN(n6152) );
  AOI21_X1 U7750 ( .B1(n9539), .B2(n6422), .A(n6152), .ZN(n6154) );
  NAND2_X1 U7751 ( .A1(n6153), .A2(n6154), .ZN(n6158) );
  INV_X1 U7752 ( .A(n6153), .ZN(n6156) );
  INV_X1 U7753 ( .A(n6154), .ZN(n6155) );
  NAND2_X1 U7754 ( .A1(n6156), .A2(n6155), .ZN(n6157) );
  NAND2_X1 U7755 ( .A1(n6158), .A2(n6157), .ZN(n8833) );
  INV_X1 U7756 ( .A(n6158), .ZN(n6183) );
  NAND2_X1 U7757 ( .A1(n7722), .A2(n6500), .ZN(n6160) );
  NAND2_X1 U7758 ( .A1(n6364), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6159) );
  NAND2_X1 U7759 ( .A1(n9536), .A2(n5769), .ZN(n6172) );
  NAND2_X1 U7760 ( .A1(n6161), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6170) );
  INV_X1 U7761 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9241) );
  OR2_X1 U7762 ( .A1(n5781), .A2(n9241), .ZN(n6169) );
  INV_X1 U7763 ( .A(n6164), .ZN(n6162) );
  NAND2_X1 U7764 ( .A1(n6162), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6213) );
  INV_X1 U7765 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7766 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  NAND2_X1 U7767 ( .A1(n6213), .A2(n6165), .ZN(n9240) );
  OR2_X1 U7768 ( .A1(n6412), .A2(n9240), .ZN(n6168) );
  INV_X1 U7769 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n6166) );
  OR2_X1 U7770 ( .A1(n4268), .A2(n6166), .ZN(n6167) );
  NAND4_X1 U7771 ( .A1(n6170), .A2(n6169), .A3(n6168), .A4(n6167), .ZN(n9130)
         );
  NAND2_X1 U7772 ( .A1(n9130), .A2(n6422), .ZN(n6171) );
  NAND2_X1 U7773 ( .A1(n6172), .A2(n6171), .ZN(n6174) );
  XNOR2_X1 U7774 ( .A(n6174), .B(n6173), .ZN(n6176) );
  AND2_X1 U7775 ( .A1(n9130), .A2(n6421), .ZN(n6175) );
  AOI21_X1 U7776 ( .B1(n9536), .B2(n6422), .A(n6175), .ZN(n6177) );
  NAND2_X1 U7777 ( .A1(n6176), .A2(n6177), .ZN(n6357) );
  INV_X1 U7778 ( .A(n6176), .ZN(n6179) );
  INV_X1 U7779 ( .A(n6177), .ZN(n6178) );
  NAND2_X1 U7780 ( .A1(n6179), .A2(n6178), .ZN(n6180) );
  AND2_X1 U7781 ( .A1(n6357), .A2(n6180), .ZN(n6182) );
  OR3_X1 U7782 ( .A1(n6181), .A2(n6183), .A3(n6182), .ZN(n6203) );
  NAND2_X1 U7783 ( .A1(n7727), .A2(P1_B_REG_SCAN_IN), .ZN(n6186) );
  MUX2_X1 U7784 ( .A(P1_B_REG_SCAN_IN), .B(n6186), .S(n7724), .Z(n6187) );
  INV_X1 U7785 ( .A(n6188), .ZN(n7798) );
  NAND2_X1 U7786 ( .A1(n7798), .A2(n7724), .ZN(n9584) );
  NOR4_X1 U7787 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6192) );
  NOR4_X1 U7788 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6191) );
  NOR4_X1 U7789 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6190) );
  NOR4_X1 U7790 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6189) );
  NAND4_X1 U7791 ( .A1(n6192), .A2(n6191), .A3(n6190), .A4(n6189), .ZN(n6198)
         );
  NOR2_X1 U7792 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n6196) );
  NOR4_X1 U7793 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6195) );
  NOR4_X1 U7794 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6194) );
  NOR4_X1 U7795 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6193) );
  NAND4_X1 U7796 ( .A1(n6196), .A2(n6195), .A3(n6194), .A4(n6193), .ZN(n6197)
         );
  NOR2_X1 U7797 ( .A1(n6198), .A2(n6197), .ZN(n6843) );
  AND2_X1 U7798 ( .A1(n6843), .A2(P1_D_REG_1__SCAN_IN), .ZN(n7263) );
  NAND2_X1 U7799 ( .A1(n7798), .A2(n7727), .ZN(n9583) );
  OAI21_X1 U7800 ( .B1(n7264), .B2(n7263), .A(n9583), .ZN(n6199) );
  OR2_X1 U7801 ( .A1(n7307), .A2(n6199), .ZN(n6204) );
  NAND2_X1 U7802 ( .A1(n6200), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6201) );
  XNOR2_X1 U7803 ( .A(n6201), .B(n4820), .ZN(n6752) );
  NOR2_X1 U7804 ( .A1(n6204), .A2(n7266), .ZN(n6208) );
  NAND2_X1 U7805 ( .A1(n7533), .A2(n7587), .ZN(n7332) );
  NAND2_X1 U7806 ( .A1(n6644), .A2(n6704), .ZN(n6835) );
  AND2_X1 U7807 ( .A1(n9983), .A2(n6835), .ZN(n6202) );
  AOI21_X1 U7808 ( .B1(n6358), .B2(n6203), .A(n8923), .ZN(n6227) );
  NOR2_X1 U7809 ( .A1(n7332), .A2(n7471), .ZN(n9667) );
  NAND2_X1 U7810 ( .A1(n9536), .A2(n8934), .ZN(n6225) );
  OAI21_X1 U7811 ( .B1(n9667), .B2(n9983), .A(n6204), .ZN(n6205) );
  NAND3_X1 U7812 ( .A1(n6205), .A2(n6731), .A3(n7268), .ZN(n6206) );
  NAND2_X1 U7813 ( .A1(n6206), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6207) );
  OR2_X1 U7814 ( .A1(n6752), .A2(P1_U3086), .ZN(n7702) );
  NAND2_X1 U7815 ( .A1(n6207), .A2(n7702), .ZN(n8921) );
  NAND2_X1 U7816 ( .A1(n6208), .A2(n6708), .ZN(n8918) );
  INV_X1 U7817 ( .A(n6835), .ZN(n6523) );
  INV_X1 U7818 ( .A(n4267), .ZN(n8990) );
  AND2_X2 U7819 ( .A1(n6523), .A2(n8990), .ZN(n8928) );
  NAND2_X1 U7820 ( .A1(n9129), .A2(n8928), .ZN(n6221) );
  NAND2_X1 U7821 ( .A1(n4273), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6219) );
  INV_X1 U7822 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n6210) );
  OR2_X1 U7823 ( .A1(n4268), .A2(n6210), .ZN(n6218) );
  INV_X1 U7824 ( .A(n6213), .ZN(n6211) );
  NAND2_X1 U7825 ( .A1(n6211), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6370) );
  INV_X1 U7826 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7827 ( .A1(n6213), .A2(n6212), .ZN(n6214) );
  NAND2_X1 U7828 ( .A1(n6370), .A2(n6214), .ZN(n9221) );
  OR2_X1 U7829 ( .A1(n6412), .A2(n9221), .ZN(n6217) );
  INV_X1 U7830 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6215) );
  OR2_X1 U7831 ( .A1(n6509), .A2(n6215), .ZN(n6216) );
  NAND4_X1 U7832 ( .A1(n6219), .A2(n6218), .A3(n6217), .A4(n6216), .ZN(n9132)
         );
  NAND2_X1 U7833 ( .A1(n6523), .A2(n4267), .ZN(n7569) );
  INV_X2 U7834 ( .A(n7569), .ZN(n8929) );
  NAND2_X1 U7835 ( .A1(n9132), .A2(n8929), .ZN(n6220) );
  NAND2_X1 U7836 ( .A1(n6221), .A2(n6220), .ZN(n9247) );
  AOI22_X1 U7837 ( .A1(n8948), .A2(n9247), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n6222) );
  OAI21_X1 U7838 ( .B1(n8944), .B2(n9240), .A(n6222), .ZN(n6223) );
  INV_X1 U7839 ( .A(n6223), .ZN(n6224) );
  NAND2_X1 U7840 ( .A1(n6228), .A2(n4275), .ZN(n6998) );
  AND3_X1 U7841 ( .A1(n6229), .A2(n8437), .A3(n6998), .ZN(n6230) );
  INV_X1 U7842 ( .A(n6977), .ZN(n6233) );
  NOR2_X1 U7843 ( .A1(n10069), .A2(n8383), .ZN(n6927) );
  OR2_X1 U7844 ( .A1(n6231), .A2(n8412), .ZN(n6232) );
  AND2_X1 U7845 ( .A1(n6232), .A2(n8355), .ZN(n6923) );
  OAI21_X1 U7846 ( .B1(n6233), .B2(n6927), .A(n6923), .ZN(n6237) );
  INV_X1 U7847 ( .A(n6923), .ZN(n6234) );
  NAND2_X1 U7848 ( .A1(n6235), .A2(n6234), .ZN(n6236) );
  AND2_X1 U7849 ( .A1(n6237), .A2(n6236), .ZN(n6238) );
  NAND2_X1 U7850 ( .A1(n10103), .A2(n10066), .ZN(n8727) );
  NAND2_X1 U7851 ( .A1(n10100), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6239) );
  OAI21_X1 U7852 ( .B1(n6240), .B2(n10100), .A(n4892), .ZN(P2_U3488) );
  NAND2_X1 U7853 ( .A1(n6999), .A2(n8355), .ZN(n6241) );
  NAND2_X1 U7854 ( .A1(n6241), .A2(n7012), .ZN(n6347) );
  NAND2_X1 U7855 ( .A1(n6347), .A2(n6242), .ZN(n6243) );
  NAND2_X1 U7856 ( .A1(n6243), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  XNOR2_X1 U7857 ( .A(n5559), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n6343) );
  INV_X1 U7858 ( .A(n7891), .ZN(n6824) );
  INV_X1 U7859 ( .A(n6324), .ZN(n7115) );
  INV_X1 U7860 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U7861 ( .A1(n4954), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6245) );
  INV_X1 U7862 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6942) );
  INV_X1 U7863 ( .A(n6245), .ZN(n6246) );
  NOR2_X1 U7864 ( .A1(n6940), .A2(n6246), .ZN(n7038) );
  INV_X1 U7865 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6247) );
  MUX2_X1 U7866 ( .A(n6247), .B(P2_REG1_REG_2__SCAN_IN), .S(n7049), .Z(n7037)
         );
  AOI21_X1 U7867 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n7049), .A(n7036), .ZN(
        n6249) );
  INV_X1 U7868 ( .A(n6922), .ZN(n6248) );
  NOR2_X1 U7869 ( .A1(n6249), .A2(n6248), .ZN(n6251) );
  INV_X1 U7870 ( .A(n6251), .ZN(n6963) );
  INV_X1 U7871 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6252) );
  MUX2_X1 U7872 ( .A(n6252), .B(P2_REG1_REG_4__SCAN_IN), .S(n6972), .Z(n6964)
         );
  INV_X1 U7873 ( .A(n6749), .ZN(n7063) );
  AOI21_X1 U7874 ( .B1(n6253), .B2(n7063), .A(n6254), .ZN(n7050) );
  INV_X1 U7875 ( .A(n6254), .ZN(n7105) );
  INV_X1 U7876 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6255) );
  XNOR2_X1 U7877 ( .A(n6324), .B(n6255), .ZN(n7106) );
  INV_X1 U7878 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6257) );
  XNOR2_X1 U7879 ( .A(n6284), .B(n6257), .ZN(n7240) );
  INV_X1 U7880 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10094) );
  NAND2_X1 U7881 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n6775), .ZN(n6260) );
  OAI21_X1 U7882 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n6775), .A(n6260), .ZN(
        n7705) );
  NOR2_X1 U7883 ( .A1(n7812), .A2(n6262), .ZN(n6263) );
  INV_X1 U7884 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10098) );
  INV_X1 U7885 ( .A(n7812), .ZN(n6820) );
  INV_X1 U7886 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10101) );
  AOI22_X1 U7887 ( .A1(n7891), .A2(P2_REG1_REG_12__SCAN_IN), .B1(n10101), .B2(
        n6824), .ZN(n7878) );
  NOR2_X1 U7888 ( .A1(n7879), .A2(n7878), .ZN(n7877) );
  INV_X1 U7889 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9650) );
  NOR2_X1 U7890 ( .A1(n7869), .A2(n6264), .ZN(n6265) );
  INV_X1 U7891 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9644) );
  AOI22_X1 U7892 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8479), .B1(n6859), .B2(
        n9644), .ZN(n8466) );
  INV_X1 U7893 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9298) );
  INV_X1 U7894 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8743) );
  OR2_X1 U7895 ( .A1(n8517), .A2(n8743), .ZN(n6268) );
  NAND2_X1 U7896 ( .A1(n8517), .A2(n8743), .ZN(n6267) );
  NAND2_X1 U7897 ( .A1(n6268), .A2(n6267), .ZN(n8511) );
  INV_X1 U7898 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n10018) );
  NOR2_X1 U7899 ( .A1(n7087), .A2(n6269), .ZN(n6270) );
  INV_X1 U7900 ( .A(n8530), .ZN(n7091) );
  NAND2_X1 U7901 ( .A1(n7091), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6271) );
  OAI21_X1 U7902 ( .B1(n7091), .B2(P2_REG1_REG_18__SCAN_IN), .A(n6271), .ZN(
        n8524) );
  INV_X1 U7903 ( .A(n6271), .ZN(n6272) );
  XOR2_X1 U7904 ( .A(n6343), .B(n6273), .Z(n6356) );
  NOR2_X1 U7905 ( .A1(n5561), .A2(P2_U3151), .ZN(n7875) );
  AND2_X1 U7906 ( .A1(n6347), .A2(n7875), .ZN(n6890) );
  NAND2_X1 U7907 ( .A1(n6890), .A2(n8434), .ZN(n10020) );
  XNOR2_X1 U7908 ( .A(n5559), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n6344) );
  INV_X1 U7909 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8483) );
  INV_X1 U7910 ( .A(n7348), .ZN(n6769) );
  INV_X1 U7911 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9331) );
  MUX2_X1 U7912 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9331), .S(n7049), .Z(n7041)
         );
  AND2_X1 U7913 ( .A1(n4885), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U7914 ( .A1(n4954), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6275) );
  OAI21_X1 U7915 ( .B1(n6952), .B2(n6274), .A(n6275), .ZN(n6945) );
  INV_X1 U7916 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6946) );
  OR2_X1 U7917 ( .A1(n6945), .A2(n6946), .ZN(n6943) );
  NAND2_X1 U7918 ( .A1(n6943), .A2(n6275), .ZN(n7040) );
  NAND2_X1 U7919 ( .A1(n7049), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6276) );
  NAND2_X1 U7920 ( .A1(n7039), .A2(n6276), .ZN(n6277) );
  NAND2_X1 U7921 ( .A1(n6277), .A2(n6922), .ZN(n6959) );
  INV_X1 U7922 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7194) );
  NAND2_X1 U7923 ( .A1(n6972), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U7924 ( .A1(n6962), .A2(n6279), .ZN(n6280) );
  NAND2_X1 U7925 ( .A1(n7102), .A2(n7100), .ZN(n6281) );
  XNOR2_X1 U7926 ( .A(n6324), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n7099) );
  INV_X1 U7927 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7441) );
  OR2_X1 U7928 ( .A1(n6324), .A2(n7441), .ZN(n6282) );
  NAND2_X1 U7929 ( .A1(n7104), .A2(n6282), .ZN(n6283) );
  INV_X1 U7930 ( .A(n6328), .ZN(n7178) );
  NAND2_X1 U7931 ( .A1(n6283), .A2(n7178), .ZN(n7243) );
  NAND2_X1 U7932 ( .A1(n7247), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7933 ( .A1(n7245), .A2(n6285), .ZN(n6286) );
  INV_X1 U7934 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9303) );
  AOI21_X1 U7935 ( .B1(n6769), .B2(n6286), .A(n7341), .ZN(n7715) );
  NAND2_X1 U7936 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n6775), .ZN(n6287) );
  OAI21_X1 U7937 ( .B1(n6775), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6287), .ZN(
        n7714) );
  NOR2_X1 U7938 ( .A1(n7715), .A2(n7714), .ZN(n7713) );
  NOR2_X1 U7939 ( .A1(n7812), .A2(n6289), .ZN(n6290) );
  INV_X1 U7940 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9300) );
  INV_X1 U7941 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6291) );
  MUX2_X1 U7942 ( .A(n6291), .B(P2_REG2_REG_12__SCAN_IN), .S(n7891), .Z(n6292)
         );
  INV_X1 U7943 ( .A(n6292), .ZN(n7887) );
  NOR2_X1 U7944 ( .A1(n7869), .A2(n6293), .ZN(n6294) );
  INV_X1 U7945 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7864) );
  INV_X1 U7946 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6295) );
  AOI22_X1 U7947 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8479), .B1(n6859), .B2(
        n6295), .ZN(n8475) );
  XNOR2_X1 U7948 ( .A(n6296), .B(n8497), .ZN(n8484) );
  NOR2_X1 U7949 ( .A1(n8483), .A2(n8484), .ZN(n8482) );
  NOR2_X1 U7950 ( .A1(n8497), .A2(n6296), .ZN(n6297) );
  INV_X1 U7951 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8683) );
  OR2_X1 U7952 ( .A1(n8517), .A2(n8683), .ZN(n6299) );
  NAND2_X1 U7953 ( .A1(n8517), .A2(n8683), .ZN(n6298) );
  NAND2_X1 U7954 ( .A1(n6299), .A2(n6298), .ZN(n8502) );
  NOR2_X1 U7955 ( .A1(n7087), .A2(n6300), .ZN(n6301) );
  INV_X1 U7956 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n10025) );
  NOR2_X1 U7957 ( .A1(n6301), .A2(n10023), .ZN(n8522) );
  INV_X1 U7958 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8660) );
  MUX2_X1 U7959 ( .A(P2_REG2_REG_18__SCAN_IN), .B(n8660), .S(n8530), .Z(n8521)
         );
  NOR2_X1 U7960 ( .A1(n8520), .A2(n6302), .ZN(n6303) );
  NAND2_X1 U7961 ( .A1(n6890), .A2(n6316), .ZN(n10026) );
  MUX2_X1 U7962 ( .A(n10025), .B(n10018), .S(n8434), .Z(n6304) );
  NAND2_X1 U7963 ( .A1(n6304), .A2(n7087), .ZN(n6338) );
  XOR2_X1 U7964 ( .A(n7087), .B(n6304), .Z(n10016) );
  MUX2_X1 U7965 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8434), .Z(n6306) );
  INV_X1 U7966 ( .A(n6306), .ZN(n6305) );
  NAND2_X1 U7967 ( .A1(n8517), .A2(n6305), .ZN(n6337) );
  XNOR2_X1 U7968 ( .A(n6306), .B(n8517), .ZN(n8506) );
  MUX2_X1 U7969 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8434), .Z(n6308) );
  INV_X1 U7970 ( .A(n6308), .ZN(n6307) );
  NAND2_X1 U7971 ( .A1(n8497), .A2(n6307), .ZN(n6336) );
  XNOR2_X1 U7972 ( .A(n6308), .B(n8497), .ZN(n8487) );
  MUX2_X1 U7973 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8434), .Z(n6309) );
  OR2_X1 U7974 ( .A1(n6309), .A2(n6859), .ZN(n6335) );
  XNOR2_X1 U7975 ( .A(n6309), .B(n8479), .ZN(n8469) );
  MUX2_X1 U7976 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8434), .Z(n6311) );
  INV_X1 U7977 ( .A(n6311), .ZN(n6310) );
  NAND2_X1 U7978 ( .A1(n7869), .A2(n6310), .ZN(n6334) );
  XNOR2_X1 U7979 ( .A(n6311), .B(n7869), .ZN(n7858) );
  MUX2_X1 U7980 ( .A(n6291), .B(n10101), .S(n8434), .Z(n6312) );
  NAND2_X1 U7981 ( .A1(n6312), .A2(n7891), .ZN(n6333) );
  XNOR2_X1 U7982 ( .A(n6312), .B(n6824), .ZN(n7882) );
  MUX2_X1 U7983 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8434), .Z(n6313) );
  OR2_X1 U7984 ( .A1(n6313), .A2(n6820), .ZN(n6332) );
  XNOR2_X1 U7985 ( .A(n6313), .B(n7812), .ZN(n7805) );
  MUX2_X1 U7986 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8434), .Z(n6314) );
  OR2_X1 U7987 ( .A1(n6314), .A2(n6775), .ZN(n6331) );
  XNOR2_X1 U7988 ( .A(n6314), .B(n7719), .ZN(n7709) );
  MUX2_X1 U7989 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8434), .Z(n6315) );
  OR2_X1 U7990 ( .A1(n6315), .A2(n6769), .ZN(n6330) );
  XNOR2_X1 U7991 ( .A(n6315), .B(n7348), .ZN(n7350) );
  MUX2_X1 U7992 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8434), .Z(n6325) );
  MUX2_X1 U7993 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8434), .Z(n6323) );
  MUX2_X1 U7994 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8434), .Z(n6322) );
  MUX2_X1 U7995 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8434), .Z(n6321) );
  MUX2_X1 U7996 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n5562), .Z(n6320) );
  MUX2_X1 U7997 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n5562), .Z(n6319) );
  XNOR2_X1 U7998 ( .A(n6317), .B(n6319), .ZN(n6936) );
  INV_X1 U7999 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6318) );
  MUX2_X1 U8000 ( .A(n6318), .B(n6244), .S(n5562), .Z(n6888) );
  NAND2_X1 U8001 ( .A1(n6888), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6935) );
  AND2_X1 U8002 ( .A1(n6936), .A2(n6935), .ZN(n6938) );
  AOI21_X1 U8003 ( .B1(n6319), .B2(n6952), .A(n6938), .ZN(n7034) );
  XNOR2_X1 U8004 ( .A(n6320), .B(n7049), .ZN(n7035) );
  NOR2_X1 U8005 ( .A1(n7034), .A2(n7035), .ZN(n7033) );
  XOR2_X1 U8006 ( .A(n6922), .B(n6321), .Z(n6909) );
  NAND2_X1 U8007 ( .A1(n6910), .A2(n6909), .ZN(n6908) );
  OAI21_X1 U8008 ( .B1(n6321), .B2(n6922), .A(n6908), .ZN(n6956) );
  XNOR2_X1 U8009 ( .A(n6322), .B(n6972), .ZN(n6957) );
  NOR2_X1 U8010 ( .A1(n6956), .A2(n6957), .ZN(n6955) );
  XNOR2_X1 U8011 ( .A(n6323), .B(n6749), .ZN(n7060) );
  NOR2_X1 U8012 ( .A1(n7059), .A2(n7060), .ZN(n7058) );
  XNOR2_X1 U8013 ( .A(n6325), .B(n6324), .ZN(n7096) );
  NAND2_X1 U8014 ( .A1(n7097), .A2(n7096), .ZN(n7095) );
  OAI21_X1 U8015 ( .B1(n6325), .B2(n7115), .A(n7095), .ZN(n7173) );
  MUX2_X1 U8016 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8434), .Z(n6326) );
  XNOR2_X1 U8017 ( .A(n6326), .B(n6328), .ZN(n7174) );
  INV_X1 U8018 ( .A(n6326), .ZN(n6327) );
  AOI22_X1 U8019 ( .A1(n7173), .A2(n7174), .B1(n6328), .B2(n6327), .ZN(n7237)
         );
  MUX2_X1 U8020 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8434), .Z(n6329) );
  XNOR2_X1 U8021 ( .A(n6329), .B(n7247), .ZN(n7238) );
  NAND2_X1 U8022 ( .A1(n7350), .A2(n7351), .ZN(n7349) );
  NAND2_X1 U8023 ( .A1(n6330), .A2(n7349), .ZN(n7708) );
  NAND2_X1 U8024 ( .A1(n7709), .A2(n7708), .ZN(n7707) );
  NAND2_X1 U8025 ( .A1(n6331), .A2(n7707), .ZN(n7804) );
  NAND2_X1 U8026 ( .A1(n7805), .A2(n7804), .ZN(n7803) );
  NAND2_X1 U8027 ( .A1(n6332), .A2(n7803), .ZN(n7881) );
  NAND2_X1 U8028 ( .A1(n7882), .A2(n7881), .ZN(n7880) );
  NAND2_X1 U8029 ( .A1(n6333), .A2(n7880), .ZN(n7859) );
  NAND2_X1 U8030 ( .A1(n7858), .A2(n7859), .ZN(n7857) );
  NAND2_X1 U8031 ( .A1(n6334), .A2(n7857), .ZN(n8468) );
  NAND2_X1 U8032 ( .A1(n8469), .A2(n8468), .ZN(n8467) );
  NAND2_X1 U8033 ( .A1(n6335), .A2(n8467), .ZN(n8486) );
  NAND2_X1 U8034 ( .A1(n8487), .A2(n8486), .ZN(n8485) );
  NAND2_X1 U8035 ( .A1(n6336), .A2(n8485), .ZN(n8505) );
  NAND2_X1 U8036 ( .A1(n8506), .A2(n8505), .ZN(n8504) );
  NAND2_X1 U8037 ( .A1(n6337), .A2(n8504), .ZN(n10015) );
  NAND2_X1 U8038 ( .A1(n10016), .A2(n10015), .ZN(n10014) );
  NAND2_X1 U8039 ( .A1(n6338), .A2(n10014), .ZN(n6341) );
  INV_X1 U8040 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n6339) );
  MUX2_X1 U8041 ( .A(n8660), .B(n6339), .S(n8434), .Z(n6340) );
  NAND2_X1 U8042 ( .A1(n6341), .A2(n6340), .ZN(n8525) );
  NAND2_X1 U8043 ( .A1(n8525), .A2(n7091), .ZN(n6342) );
  OR2_X1 U8044 ( .A1(n6341), .A2(n6340), .ZN(n8526) );
  NAND2_X1 U8045 ( .A1(n6342), .A2(n8526), .ZN(n6346) );
  MUX2_X1 U8046 ( .A(n6344), .B(n6343), .S(n8434), .Z(n6345) );
  XNOR2_X1 U8047 ( .A(n6346), .B(n6345), .ZN(n6354) );
  NOR2_X1 U8048 ( .A1(n8434), .A2(P2_U3151), .ZN(n7828) );
  NAND2_X1 U8049 ( .A1(n6347), .A2(n7828), .ZN(n6348) );
  INV_X1 U8050 ( .A(n5561), .ZN(n8435) );
  MUX2_X1 U8051 ( .A(n6348), .B(n8463), .S(n8435), .Z(n10012) );
  INV_X1 U8052 ( .A(n7012), .ZN(n6349) );
  NOR2_X1 U8053 ( .A1(n6999), .A2(n6349), .ZN(n6350) );
  NAND2_X1 U8054 ( .A1(n7807), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n6352) );
  NAND2_X1 U8055 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3151), .ZN(n6351) );
  OAI211_X1 U8056 ( .C1(n10012), .C2(n5559), .A(n6352), .B(n6351), .ZN(n6353)
         );
  NAND2_X1 U8057 ( .A1(n7725), .A2(n6500), .ZN(n6360) );
  NAND2_X1 U8058 ( .A1(n6364), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6359) );
  NAND2_X1 U8059 ( .A1(n9530), .A2(n5769), .ZN(n6362) );
  NAND2_X1 U8060 ( .A1(n9132), .A2(n6422), .ZN(n6361) );
  NAND2_X1 U8061 ( .A1(n6362), .A2(n6361), .ZN(n6363) );
  XNOR2_X1 U8062 ( .A(n6363), .B(n6394), .ZN(n6381) );
  AOI22_X1 U8063 ( .A1(n9530), .A2(n6422), .B1(n6421), .B2(n9132), .ZN(n6382)
         );
  XNOR2_X1 U8064 ( .A(n6381), .B(n6382), .ZN(n8866) );
  NAND2_X1 U8065 ( .A1(n7793), .A2(n6500), .ZN(n6366) );
  NAND2_X1 U8066 ( .A1(n6364), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6365) );
  NAND2_X1 U8067 ( .A1(n9525), .A2(n5769), .ZN(n6378) );
  NAND2_X1 U8068 ( .A1(n4272), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6376) );
  INV_X1 U8069 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n6367) );
  OR2_X1 U8070 ( .A1(n4268), .A2(n6367), .ZN(n6375) );
  INV_X1 U8071 ( .A(n6370), .ZN(n6368) );
  INV_X1 U8072 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6369) );
  NAND2_X1 U8073 ( .A1(n6370), .A2(n6369), .ZN(n6371) );
  NAND2_X1 U8074 ( .A1(n6408), .A2(n6371), .ZN(n9207) );
  OR2_X1 U8075 ( .A1(n6412), .A2(n9207), .ZN(n6374) );
  INV_X1 U8076 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6372) );
  OR2_X1 U8077 ( .A1(n6509), .A2(n6372), .ZN(n6373) );
  NAND4_X1 U8078 ( .A1(n6376), .A2(n6375), .A3(n6374), .A4(n6373), .ZN(n8957)
         );
  NAND2_X1 U8079 ( .A1(n8957), .A2(n6422), .ZN(n6377) );
  NAND2_X1 U8080 ( .A1(n6378), .A2(n6377), .ZN(n6379) );
  XNOR2_X1 U8081 ( .A(n6379), .B(n6394), .ZN(n6402) );
  AND2_X1 U8082 ( .A1(n8957), .A2(n6421), .ZN(n6380) );
  AOI21_X1 U8083 ( .B1(n9525), .B2(n6422), .A(n6380), .ZN(n6400) );
  XNOR2_X1 U8084 ( .A(n6402), .B(n6400), .ZN(n8926) );
  INV_X1 U8085 ( .A(n6381), .ZN(n6383) );
  NAND2_X1 U8086 ( .A1(n6383), .A2(n6382), .ZN(n8927) );
  AND2_X1 U8087 ( .A1(n8926), .A2(n8927), .ZN(n6715) );
  NAND2_X1 U8088 ( .A1(n7827), .A2(n6500), .ZN(n6385) );
  OR2_X1 U8089 ( .A1(n4274), .A2(n9408), .ZN(n6384) );
  NAND2_X1 U8090 ( .A1(n9521), .A2(n5769), .ZN(n6393) );
  NAND2_X1 U8091 ( .A1(n4272), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6391) );
  INV_X1 U8092 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6386) );
  OR2_X1 U8093 ( .A1(n6509), .A2(n6386), .ZN(n6390) );
  INV_X1 U8094 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6723) );
  XNOR2_X1 U8095 ( .A(n6408), .B(n6723), .ZN(n6720) );
  INV_X1 U8096 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n6387) );
  OR2_X1 U8097 ( .A1(n4268), .A2(n6387), .ZN(n6388) );
  NAND4_X1 U8098 ( .A1(n6391), .A2(n6390), .A3(n6389), .A4(n6388), .ZN(n8956)
         );
  NAND2_X1 U8099 ( .A1(n8956), .A2(n6422), .ZN(n6392) );
  NAND2_X1 U8100 ( .A1(n6393), .A2(n6392), .ZN(n6395) );
  XNOR2_X1 U8101 ( .A(n6395), .B(n6394), .ZN(n6399) );
  NAND2_X1 U8102 ( .A1(n9521), .A2(n6422), .ZN(n6397) );
  NAND2_X1 U8103 ( .A1(n8956), .A2(n6421), .ZN(n6396) );
  NAND2_X1 U8104 ( .A1(n6397), .A2(n6396), .ZN(n6398) );
  NOR2_X1 U8105 ( .A1(n6399), .A2(n6398), .ZN(n6439) );
  AOI21_X1 U8106 ( .B1(n6399), .B2(n6398), .A(n6439), .ZN(n6716) );
  INV_X1 U8107 ( .A(n6400), .ZN(n6401) );
  NAND2_X1 U8108 ( .A1(n6402), .A2(n6401), .ZN(n6717) );
  NAND2_X1 U8109 ( .A1(n6716), .A2(n6717), .ZN(n6403) );
  NAND2_X1 U8110 ( .A1(n7874), .A2(n6500), .ZN(n6405) );
  OR2_X1 U8111 ( .A1(n4274), .A2(n8057), .ZN(n6404) );
  NAND2_X1 U8112 ( .A1(n9515), .A2(n5769), .ZN(n6419) );
  NAND2_X1 U8113 ( .A1(n4273), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6417) );
  INV_X1 U8114 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6406) );
  OR2_X1 U8115 ( .A1(n4268), .A2(n6406), .ZN(n6416) );
  INV_X1 U8116 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6407) );
  OAI21_X1 U8117 ( .B1(n6408), .B2(n6723), .A(n6407), .ZN(n6411) );
  INV_X1 U8118 ( .A(n6408), .ZN(n6410) );
  AND2_X1 U8119 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .ZN(n6409) );
  NAND2_X1 U8120 ( .A1(n6410), .A2(n6409), .ZN(n9143) );
  NAND2_X1 U8121 ( .A1(n6411), .A2(n9143), .ZN(n9177) );
  OR2_X1 U8122 ( .A1(n6412), .A2(n9177), .ZN(n6415) );
  INV_X1 U8123 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6413) );
  OR2_X1 U8124 ( .A1(n6509), .A2(n6413), .ZN(n6414) );
  NAND4_X1 U8125 ( .A1(n6417), .A2(n6416), .A3(n6415), .A4(n6414), .ZN(n8955)
         );
  NAND2_X1 U8126 ( .A1(n8955), .A2(n6422), .ZN(n6418) );
  NAND2_X1 U8127 ( .A1(n6419), .A2(n6418), .ZN(n6420) );
  XNOR2_X1 U8128 ( .A(n6420), .B(n6394), .ZN(n6424) );
  AOI22_X1 U8129 ( .A1(n9515), .A2(n6422), .B1(n6421), .B2(n8955), .ZN(n6423)
         );
  XNOR2_X1 U8130 ( .A(n6424), .B(n6423), .ZN(n6442) );
  AND2_X1 U8131 ( .A1(n6442), .A2(n8941), .ZN(n6438) );
  NAND3_X1 U8132 ( .A1(n6442), .A2(n8941), .A3(n6439), .ZN(n6436) );
  NAND2_X1 U8133 ( .A1(n4272), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6430) );
  INV_X1 U8134 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6425) );
  OR2_X1 U8135 ( .A1(n6509), .A2(n6425), .ZN(n6429) );
  OR2_X1 U8136 ( .A1(n6412), .A2(n9143), .ZN(n6428) );
  INV_X1 U8137 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6426) );
  OR2_X1 U8138 ( .A1(n4268), .A2(n6426), .ZN(n6427) );
  NAND4_X1 U8139 ( .A1(n6430), .A2(n6429), .A3(n6428), .A4(n6427), .ZN(n8954)
         );
  NAND2_X1 U8140 ( .A1(n8954), .A2(n8929), .ZN(n6432) );
  NAND2_X1 U8141 ( .A1(n8956), .A2(n8928), .ZN(n6431) );
  NAND2_X1 U8142 ( .A1(n6432), .A2(n6431), .ZN(n9182) );
  AOI22_X1 U8143 ( .A1(n8948), .A2(n9182), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6433) );
  OAI21_X1 U8144 ( .B1(n8944), .B2(n9177), .A(n6433), .ZN(n6434) );
  AOI21_X1 U8145 ( .B1(n9515), .B2(n8934), .A(n6434), .ZN(n6435) );
  AOI21_X1 U8146 ( .B1(n6718), .B2(n6438), .A(n6437), .ZN(n6445) );
  INV_X1 U8147 ( .A(n6439), .ZN(n6440) );
  NAND2_X1 U8148 ( .A1(n6440), .A2(n8941), .ZN(n6441) );
  NAND2_X1 U8149 ( .A1(n6445), .A2(n6444), .ZN(P1_U3220) );
  NAND2_X1 U8150 ( .A1(n6446), .A2(n6500), .ZN(n6448) );
  OR2_X1 U8151 ( .A1(n4274), .A2(n8063), .ZN(n6447) );
  INV_X1 U8152 ( .A(n8954), .ZN(n6510) );
  AND2_X1 U8153 ( .A1(n6627), .A2(n9161), .ZN(n6640) );
  NOR2_X1 U8154 ( .A1(n8975), .A2(n7523), .ZN(n7517) );
  INV_X1 U8155 ( .A(n8973), .ZN(n6904) );
  NAND2_X1 U8156 ( .A1(n6904), .A2(n4314), .ZN(n6450) );
  INV_X1 U8157 ( .A(n8972), .ZN(n7276) );
  NAND2_X1 U8158 ( .A1(n7276), .A2(n4269), .ZN(n6451) );
  INV_X1 U8159 ( .A(n4269), .ZN(n9913) );
  AND2_X1 U8160 ( .A1(n9913), .A2(n8972), .ZN(n6643) );
  INV_X1 U8161 ( .A(n8971), .ZN(n7288) );
  NAND2_X1 U8162 ( .A1(n7288), .A2(n4271), .ZN(n6452) );
  NAND2_X1 U8163 ( .A1(n8970), .A2(n9925), .ZN(n6649) );
  INV_X1 U8164 ( .A(n8970), .ZN(n7291) );
  NAND2_X1 U8165 ( .A1(n7291), .A2(n7299), .ZN(n6550) );
  INV_X1 U8166 ( .A(n8969), .ZN(n7312) );
  NAND2_X1 U8167 ( .A1(n7312), .A2(n9932), .ZN(n6650) );
  NAND2_X1 U8168 ( .A1(n7311), .A2(n8969), .ZN(n6653) );
  NAND2_X1 U8169 ( .A1(n6650), .A2(n6653), .ZN(n7309) );
  INV_X1 U8170 ( .A(n8965), .ZN(n6455) );
  NAND2_X1 U8171 ( .A1(n7680), .A2(n6455), .ZN(n7482) );
  INV_X1 U8172 ( .A(n8966), .ZN(n7563) );
  NAND2_X1 U8173 ( .A1(n9836), .A2(n7563), .ZN(n7480) );
  INV_X1 U8174 ( .A(n8967), .ZN(n7476) );
  NAND2_X1 U8175 ( .A1(n7455), .A2(n7476), .ZN(n7559) );
  AND2_X1 U8176 ( .A1(n7480), .A2(n7559), .ZN(n6554) );
  AND2_X1 U8177 ( .A1(n7482), .A2(n6554), .ZN(n6532) );
  INV_X1 U8178 ( .A(n6532), .ZN(n6456) );
  INV_X1 U8179 ( .A(n8968), .ZN(n7314) );
  NAND2_X1 U8180 ( .A1(n7314), .A2(n7324), .ZN(n7318) );
  INV_X1 U8181 ( .A(n7318), .ZN(n6453) );
  NOR2_X1 U8182 ( .A1(n6456), .A2(n6453), .ZN(n6454) );
  NAND2_X1 U8183 ( .A1(n9843), .A2(n6454), .ZN(n6461) );
  OR2_X1 U8184 ( .A1(n7680), .A2(n6455), .ZN(n7483) );
  OR2_X1 U8185 ( .A1(n9836), .A2(n7563), .ZN(n7561) );
  AND2_X1 U8186 ( .A1(n7483), .A2(n7561), .ZN(n6557) );
  INV_X1 U8187 ( .A(n6557), .ZN(n6459) );
  NAND2_X1 U8188 ( .A1(n6459), .A2(n7482), .ZN(n6457) );
  NAND2_X1 U8189 ( .A1(n6457), .A2(n6456), .ZN(n6659) );
  INV_X1 U8190 ( .A(n7455), .ZN(n7477) );
  NAND2_X1 U8191 ( .A1(n7477), .A2(n8967), .ZN(n6553) );
  INV_X1 U8192 ( .A(n6553), .ZN(n6458) );
  INV_X1 U8193 ( .A(n7324), .ZN(n9940) );
  NAND2_X1 U8194 ( .A1(n9940), .A2(n8968), .ZN(n7313) );
  INV_X1 U8195 ( .A(n7313), .ZN(n7317) );
  NAND2_X1 U8196 ( .A1(n6659), .A2(n6526), .ZN(n6460) );
  NAND2_X1 U8197 ( .A1(n6461), .A2(n6460), .ZN(n7501) );
  INV_X1 U8198 ( .A(n8964), .ZN(n6462) );
  OR2_X1 U8199 ( .A1(n7512), .A2(n6462), .ZN(n6565) );
  INV_X1 U8200 ( .A(n8963), .ZN(n7611) );
  NAND2_X1 U8201 ( .A1(n7853), .A2(n7611), .ZN(n6567) );
  NAND2_X1 U8202 ( .A1(n6566), .A2(n6567), .ZN(n7612) );
  INV_X1 U8203 ( .A(n8962), .ZN(n6464) );
  NAND2_X1 U8204 ( .A1(n6463), .A2(n6464), .ZN(n6664) );
  INV_X1 U8205 ( .A(n8961), .ZN(n7784) );
  OR2_X1 U8206 ( .A1(n7696), .A2(n7784), .ZN(n6666) );
  NAND2_X1 U8207 ( .A1(n7696), .A2(n7784), .ZN(n9809) );
  INV_X1 U8208 ( .A(n8960), .ZN(n6465) );
  OR2_X2 U8209 ( .A1(n9817), .A2(n6465), .ZN(n7778) );
  NAND2_X1 U8210 ( .A1(n9817), .A2(n6465), .ZN(n6584) );
  NAND2_X1 U8211 ( .A1(n7778), .A2(n6584), .ZN(n6575) );
  INV_X1 U8212 ( .A(n9809), .ZN(n6572) );
  NOR2_X1 U8213 ( .A1(n6575), .A2(n6572), .ZN(n6466) );
  INV_X1 U8214 ( .A(n8959), .ZN(n9108) );
  INV_X1 U8215 ( .A(n7778), .ZN(n6467) );
  NOR2_X1 U8216 ( .A1(n9109), .A2(n6467), .ZN(n6468) );
  OR2_X1 U8217 ( .A1(n9668), .A2(n6469), .ZN(n6675) );
  NAND2_X1 U8218 ( .A1(n9668), .A2(n6469), .ZN(n6672) );
  NAND2_X1 U8219 ( .A1(n9664), .A2(n6672), .ZN(n9490) );
  INV_X1 U8220 ( .A(n9112), .ZN(n6471) );
  NAND2_X1 U8221 ( .A1(n9502), .A2(n6471), .ZN(n6593) );
  INV_X1 U8222 ( .A(n6593), .ZN(n6470) );
  INV_X1 U8223 ( .A(n8958), .ZN(n9113) );
  OR2_X1 U8224 ( .A1(n9566), .A2(n9113), .ZN(n6596) );
  NAND2_X1 U8225 ( .A1(n6596), .A2(n9473), .ZN(n6678) );
  NAND2_X1 U8226 ( .A1(n9566), .A2(n9113), .ZN(n6594) );
  INV_X1 U8227 ( .A(n9115), .ZN(n9114) );
  OR2_X1 U8228 ( .A1(n9561), .A2(n9114), .ZN(n6597) );
  NAND2_X1 U8229 ( .A1(n9561), .A2(n9114), .ZN(n6598) );
  INV_X1 U8230 ( .A(n6598), .ZN(n6679) );
  INV_X1 U8231 ( .A(n8956), .ZN(n9139) );
  NOR2_X1 U8232 ( .A1(n9521), .A2(n9139), .ZN(n6616) );
  INV_X1 U8233 ( .A(n6616), .ZN(n6621) );
  INV_X1 U8234 ( .A(n8957), .ZN(n6481) );
  OR2_X1 U8235 ( .A1(n9525), .A2(n6481), .ZN(n9192) );
  INV_X1 U8236 ( .A(n9132), .ZN(n9133) );
  OR2_X1 U8237 ( .A1(n9530), .A2(n9133), .ZN(n9156) );
  AND2_X1 U8238 ( .A1(n9192), .A2(n9156), .ZN(n6615) );
  INV_X1 U8239 ( .A(n9129), .ZN(n9128) );
  INV_X1 U8240 ( .A(n9125), .ZN(n9124) );
  OR2_X1 U8241 ( .A1(n9124), .A2(n9546), .ZN(n9152) );
  INV_X1 U8242 ( .A(n9121), .ZN(n9120) );
  INV_X1 U8243 ( .A(n9118), .ZN(n6475) );
  OR2_X1 U8244 ( .A1(n9556), .A2(n6475), .ZN(n6590) );
  AND2_X1 U8245 ( .A1(n6591), .A2(n6590), .ZN(n6601) );
  INV_X1 U8246 ( .A(n6601), .ZN(n6473) );
  NOR2_X1 U8247 ( .A1(n6604), .A2(n6473), .ZN(n6474) );
  INV_X1 U8248 ( .A(n9130), .ZN(n6478) );
  NAND4_X1 U8249 ( .A1(n6621), .A2(n6615), .A3(n6474), .A4(n9155), .ZN(n6683)
         );
  NAND2_X1 U8250 ( .A1(n9515), .A2(n9168), .ZN(n6623) );
  NAND2_X1 U8251 ( .A1(n9521), .A2(n9139), .ZN(n9160) );
  NAND2_X1 U8252 ( .A1(n6623), .A2(n9160), .ZN(n6618) );
  NAND2_X1 U8253 ( .A1(n9546), .A2(n9124), .ZN(n9153) );
  NAND2_X1 U8254 ( .A1(n9551), .A2(n9120), .ZN(n6599) );
  NAND2_X1 U8255 ( .A1(n9556), .A2(n6475), .ZN(n9148) );
  NAND2_X1 U8256 ( .A1(n6599), .A2(n9148), .ZN(n6476) );
  NAND2_X1 U8257 ( .A1(n6476), .A2(n6591), .ZN(n9150) );
  AND2_X1 U8258 ( .A1(n9153), .A2(n9150), .ZN(n6477) );
  OAI21_X1 U8259 ( .B1(n6604), .B2(n6477), .A(n4340), .ZN(n6480) );
  NAND2_X1 U8260 ( .A1(n9536), .A2(n6478), .ZN(n6613) );
  INV_X1 U8261 ( .A(n6613), .ZN(n6479) );
  AOI21_X1 U8262 ( .B1(n9155), .B2(n6480), .A(n6479), .ZN(n6482) );
  NAND2_X1 U8263 ( .A1(n9525), .A2(n6481), .ZN(n6617) );
  AND2_X1 U8264 ( .A1(n9530), .A2(n9133), .ZN(n9211) );
  NAND2_X1 U8265 ( .A1(n6617), .A2(n4554), .ZN(n9159) );
  NAND2_X1 U8266 ( .A1(n9159), .A2(n9192), .ZN(n9189) );
  OAI21_X1 U8267 ( .B1(n4551), .B2(n6482), .A(n9189), .ZN(n6483) );
  AND2_X1 U8268 ( .A1(n6483), .A2(n6621), .ZN(n6484) );
  NOR2_X1 U8269 ( .A1(n6618), .A2(n6484), .ZN(n6641) );
  OAI21_X1 U8270 ( .B1(n9446), .B2(n6683), .A(n6641), .ZN(n6503) );
  NAND2_X1 U8271 ( .A1(n4272), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6489) );
  INV_X1 U8272 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6485) );
  OR2_X1 U8273 ( .A1(n6509), .A2(n6485), .ZN(n6488) );
  INV_X1 U8274 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6486) );
  OR2_X1 U8275 ( .A1(n4268), .A2(n6486), .ZN(n6487) );
  AND3_X1 U8276 ( .A1(n6489), .A2(n6488), .A3(n6487), .ZN(n9098) );
  INV_X1 U8277 ( .A(SI_29_), .ZN(n6490) );
  INV_X1 U8278 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8820) );
  INV_X1 U8279 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7921) );
  MUX2_X1 U8280 ( .A(n8820), .B(n7921), .S(n4425), .Z(n6497) );
  INV_X1 U8281 ( .A(SI_30_), .ZN(n6496) );
  NAND2_X1 U8282 ( .A1(n6497), .A2(n6496), .ZN(n6514) );
  INV_X1 U8283 ( .A(n6497), .ZN(n6498) );
  NAND2_X1 U8284 ( .A1(n6498), .A2(SI_30_), .ZN(n6499) );
  NAND2_X1 U8285 ( .A1(n6514), .A2(n6499), .ZN(n6515) );
  NAND2_X1 U8286 ( .A1(n8210), .A2(n6500), .ZN(n6502) );
  OR2_X1 U8287 ( .A1(n4274), .A2(n7921), .ZN(n6501) );
  AOI22_X1 U8288 ( .A1(n6640), .A2(n6503), .B1(n9098), .B2(n9105), .ZN(n6513)
         );
  INV_X1 U8289 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6508) );
  NAND2_X1 U8290 ( .A1(n4273), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6507) );
  INV_X1 U8291 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n6504) );
  OR2_X1 U8292 ( .A1(n4268), .A2(n6504), .ZN(n6506) );
  OAI211_X1 U8293 ( .C1(n6509), .C2(n6508), .A(n6507), .B(n6506), .ZN(n8953)
         );
  INV_X1 U8294 ( .A(n8953), .ZN(n9165) );
  NAND2_X1 U8295 ( .A1(n9105), .A2(n9165), .ZN(n6511) );
  NAND2_X1 U8296 ( .A1(n9510), .A2(n6510), .ZN(n6628) );
  AND2_X1 U8297 ( .A1(n6511), .A2(n6628), .ZN(n6688) );
  INV_X1 U8298 ( .A(n9098), .ZN(n8952) );
  NAND2_X1 U8299 ( .A1(n8952), .A2(n8953), .ZN(n6631) );
  INV_X1 U8300 ( .A(n6631), .ZN(n6512) );
  AOI22_X1 U8301 ( .A1(n6513), .A2(n6688), .B1(n9508), .B2(n6512), .ZN(n6525)
         );
  MUX2_X1 U8302 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n4425), .Z(n6517) );
  XNOR2_X1 U8303 ( .A(n6517), .B(SI_31_), .ZN(n6518) );
  INV_X1 U8304 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6520) );
  OR2_X1 U8305 ( .A1(n4274), .A2(n6520), .ZN(n6521) );
  OR2_X1 U8306 ( .A1(n9099), .A2(n9098), .ZN(n6706) );
  INV_X1 U8307 ( .A(n6706), .ZN(n6524) );
  NAND2_X1 U8308 ( .A1(n9099), .A2(n9098), .ZN(n6700) );
  OAI211_X1 U8309 ( .C1(n6525), .C2(n6524), .A(n6523), .B(n6700), .ZN(n6546)
         );
  NAND2_X1 U8310 ( .A1(n9161), .A2(n6623), .ZN(n9181) );
  NAND2_X1 U8311 ( .A1(n6621), .A2(n9160), .ZN(n9158) );
  OR2_X1 U8312 ( .A1(n9525), .A2(n8957), .ZN(n9138) );
  NAND2_X1 U8313 ( .A1(n9525), .A2(n8957), .ZN(n9136) );
  NAND2_X1 U8314 ( .A1(n9138), .A2(n9136), .ZN(n9213) );
  NAND2_X1 U8315 ( .A1(n9152), .A2(n9153), .ZN(n9270) );
  NAND2_X1 U8316 ( .A1(n6590), .A2(n9148), .ZN(n9445) );
  NAND2_X1 U8317 ( .A1(n6591), .A2(n6599), .ZN(n9283) );
  NAND2_X1 U8318 ( .A1(n6596), .A2(n6594), .ZN(n9475) );
  NAND2_X1 U8319 ( .A1(n9473), .A2(n6593), .ZN(n9494) );
  INV_X1 U8320 ( .A(n6526), .ZN(n6656) );
  AND2_X1 U8321 ( .A1(n6550), .A2(n6649), .ZN(n9860) );
  INV_X1 U8322 ( .A(n7517), .ZN(n6527) );
  NAND2_X1 U8323 ( .A1(n8975), .A2(n7523), .ZN(n6648) );
  AND2_X1 U8324 ( .A1(n6527), .A2(n6648), .ZN(n7331) );
  NAND4_X1 U8325 ( .A1(n7293), .A2(n9860), .A3(n7331), .A4(n7533), .ZN(n6530)
         );
  XNOR2_X1 U8326 ( .A(n8972), .B(n7278), .ZN(n7271) );
  NAND2_X1 U8327 ( .A1(n7284), .A2(n7318), .ZN(n6528) );
  NOR3_X1 U8328 ( .A1(n6530), .A2(n6529), .A3(n6528), .ZN(n6531) );
  NAND4_X1 U8329 ( .A1(n6533), .A2(n6656), .A3(n6532), .A4(n6531), .ZN(n6534)
         );
  NOR3_X1 U8330 ( .A1(n4837), .A2(n7612), .A3(n6534), .ZN(n6535) );
  NAND4_X1 U8331 ( .A1(n6536), .A2(n9808), .A3(n7684), .A4(n6535), .ZN(n6537)
         );
  NOR4_X1 U8332 ( .A1(n9475), .A2(n9494), .A3(n9662), .A4(n6537), .ZN(n6538)
         );
  NAND2_X1 U8333 ( .A1(n9465), .A2(n6538), .ZN(n6539) );
  OR4_X1 U8334 ( .A1(n9270), .A2(n9445), .A3(n9283), .A4(n6539), .ZN(n6540) );
  NOR2_X1 U8335 ( .A1(n9233), .A2(n6540), .ZN(n6541) );
  XNOR2_X1 U8336 ( .A(n9539), .B(n9129), .ZN(n9260) );
  NAND4_X1 U8337 ( .A1(n9213), .A2(n9226), .A3(n6541), .A4(n9260), .ZN(n6542)
         );
  OR3_X1 U8338 ( .A1(n9181), .A2(n9158), .A3(n6542), .ZN(n6543) );
  NOR2_X1 U8339 ( .A1(n9163), .A2(n6543), .ZN(n6545) );
  XNOR2_X1 U8340 ( .A(n9105), .B(n8953), .ZN(n6544) );
  NAND4_X1 U8341 ( .A1(n6706), .A2(n6700), .A3(n6545), .A4(n6544), .ZN(n6637)
         );
  AND2_X1 U8342 ( .A1(n6546), .A2(n6637), .ZN(n6638) );
  INV_X1 U8343 ( .A(n6838), .ZN(n6703) );
  MUX2_X1 U8344 ( .A(n6547), .B(n7294), .S(n6703), .Z(n6551) );
  INV_X1 U8345 ( .A(n6650), .ZN(n6548) );
  AND2_X1 U8346 ( .A1(n7313), .A2(n6653), .ZN(n6552) );
  OAI21_X1 U8347 ( .B1(n6551), .B2(n6548), .A(n6552), .ZN(n6549) );
  XNOR2_X1 U8348 ( .A(n7455), .B(n8967), .ZN(n7473) );
  AND2_X1 U8349 ( .A1(n7561), .A2(n6553), .ZN(n6555) );
  MUX2_X1 U8350 ( .A(n6555), .B(n6554), .S(n6838), .Z(n6556) );
  AND2_X1 U8351 ( .A1(n7482), .A2(n7480), .ZN(n6558) );
  MUX2_X1 U8352 ( .A(n6558), .B(n6557), .S(n6838), .Z(n6559) );
  INV_X1 U8353 ( .A(n6565), .ZN(n6658) );
  AOI21_X1 U8354 ( .B1(n6564), .B2(n7482), .A(n6658), .ZN(n6561) );
  NAND2_X1 U8355 ( .A1(n6567), .A2(n6560), .ZN(n6662) );
  AND2_X1 U8356 ( .A1(n6570), .A2(n6566), .ZN(n6661) );
  OAI21_X1 U8357 ( .B1(n6561), .B2(n6662), .A(n6661), .ZN(n6562) );
  AOI21_X1 U8358 ( .B1(n6564), .B2(n7483), .A(n6563), .ZN(n6569) );
  NAND2_X1 U8359 ( .A1(n6566), .A2(n6565), .ZN(n6568) );
  OAI211_X1 U8360 ( .C1(n6569), .C2(n6568), .A(n6567), .B(n6664), .ZN(n6571)
         );
  INV_X1 U8361 ( .A(n6666), .ZN(n6573) );
  MUX2_X1 U8362 ( .A(n6573), .B(n6572), .S(n6838), .Z(n6574) );
  NOR2_X1 U8363 ( .A1(n6575), .A2(n6574), .ZN(n6576) );
  NAND2_X1 U8364 ( .A1(n6669), .A2(n7778), .ZN(n6674) );
  NAND2_X1 U8365 ( .A1(n6674), .A2(n6838), .ZN(n6577) );
  INV_X1 U8366 ( .A(n6669), .ZN(n6579) );
  MUX2_X1 U8367 ( .A(n6580), .B(n6579), .S(n6703), .Z(n6581) );
  INV_X1 U8368 ( .A(n6581), .ZN(n6582) );
  NAND2_X1 U8369 ( .A1(n6583), .A2(n6582), .ZN(n6585) );
  INV_X1 U8370 ( .A(n6585), .ZN(n6589) );
  INV_X1 U8371 ( .A(n6675), .ZN(n6587) );
  AND2_X1 U8372 ( .A1(n9660), .A2(n6584), .ZN(n6668) );
  OAI211_X1 U8373 ( .C1(n6585), .C2(n6668), .A(n6593), .B(n6672), .ZN(n6586)
         );
  MUX2_X1 U8374 ( .A(n6587), .B(n6586), .S(n6703), .Z(n6588) );
  OAI211_X1 U8375 ( .C1(n6595), .C2(n6678), .A(n6598), .B(n6594), .ZN(n6592)
         );
  NAND2_X1 U8376 ( .A1(n6597), .A2(n6596), .ZN(n6642) );
  INV_X1 U8377 ( .A(n6599), .ZN(n6600) );
  AOI21_X1 U8378 ( .B1(n6602), .B2(n6601), .A(n6600), .ZN(n6603) );
  NAND2_X1 U8379 ( .A1(n6604), .A2(n6703), .ZN(n6605) );
  AOI21_X1 U8380 ( .B1(n4340), .B2(n9153), .A(n6703), .ZN(n6607) );
  INV_X1 U8381 ( .A(n9539), .ZN(n9258) );
  NAND3_X1 U8382 ( .A1(n9258), .A2(n9129), .A3(n6838), .ZN(n6610) );
  MUX2_X1 U8383 ( .A(n9155), .B(n6613), .S(n6838), .Z(n6614) );
  OAI21_X1 U8384 ( .B1(n6619), .B2(n6618), .A(n9161), .ZN(n6626) );
  OAI211_X1 U8385 ( .C1(n6620), .C2(n4551), .A(n9160), .B(n9189), .ZN(n6622)
         );
  NAND3_X1 U8386 ( .A1(n6622), .A2(n9161), .A3(n6621), .ZN(n6624) );
  NAND2_X1 U8387 ( .A1(n6624), .A2(n6623), .ZN(n6625) );
  MUX2_X1 U8388 ( .A(n6626), .B(n6625), .S(n6838), .Z(n6630) );
  MUX2_X1 U8389 ( .A(n6628), .B(n6627), .S(n6838), .Z(n6629) );
  MUX2_X1 U8390 ( .A(n6633), .B(n6703), .S(n9105), .Z(n6632) );
  NAND3_X1 U8391 ( .A1(n6632), .A2(n6706), .A3(n6631), .ZN(n6636) );
  NAND3_X1 U8392 ( .A1(n6634), .A2(n9099), .A3(n8953), .ZN(n6635) );
  NAND2_X1 U8393 ( .A1(n6639), .A2(n6837), .ZN(n6699) );
  INV_X1 U8394 ( .A(n6640), .ZN(n6687) );
  INV_X1 U8395 ( .A(n6641), .ZN(n6685) );
  INV_X1 U8396 ( .A(n6642), .ZN(n6681) );
  INV_X1 U8397 ( .A(n6643), .ZN(n6647) );
  INV_X1 U8398 ( .A(n4271), .ZN(n7287) );
  NAND2_X1 U8399 ( .A1(n8971), .A2(n7287), .ZN(n6646) );
  INV_X1 U8400 ( .A(n4314), .ZN(n9907) );
  NAND2_X1 U8401 ( .A1(n8973), .A2(n9907), .ZN(n6645) );
  NAND4_X1 U8402 ( .A1(n6647), .A2(n6646), .A3(n6645), .A4(n6644), .ZN(n6652)
         );
  NAND2_X1 U8403 ( .A1(n6649), .A2(n6648), .ZN(n6651) );
  OAI21_X1 U8404 ( .B1(n6652), .B2(n6651), .A(n6650), .ZN(n6654) );
  OAI21_X1 U8405 ( .B1(n7294), .B2(n6654), .A(n6653), .ZN(n6655) );
  NAND2_X1 U8406 ( .A1(n6655), .A2(n7318), .ZN(n6657) );
  NAND2_X1 U8407 ( .A1(n6657), .A2(n6656), .ZN(n6660) );
  AOI21_X1 U8408 ( .B1(n6660), .B2(n6659), .A(n6658), .ZN(n6663) );
  OAI21_X1 U8409 ( .B1(n6663), .B2(n6662), .A(n6661), .ZN(n6665) );
  NAND3_X1 U8410 ( .A1(n6665), .A2(n9809), .A3(n6664), .ZN(n6667) );
  NAND2_X1 U8411 ( .A1(n6667), .A2(n6666), .ZN(n6673) );
  INV_X1 U8412 ( .A(n6668), .ZN(n6670) );
  NAND2_X1 U8413 ( .A1(n6670), .A2(n6669), .ZN(n6671) );
  OAI211_X1 U8414 ( .C1(n6674), .C2(n6673), .A(n6672), .B(n6671), .ZN(n6676)
         );
  NAND2_X1 U8415 ( .A1(n6676), .A2(n6675), .ZN(n6677) );
  OAI21_X1 U8416 ( .B1(n6678), .B2(n6677), .A(n4400), .ZN(n6680) );
  AOI21_X1 U8417 ( .B1(n6681), .B2(n6680), .A(n6679), .ZN(n6682) );
  NOR2_X1 U8418 ( .A1(n6683), .A2(n6682), .ZN(n6684) );
  NOR2_X1 U8419 ( .A1(n6685), .A2(n6684), .ZN(n6686) );
  NOR2_X1 U8420 ( .A1(n6687), .A2(n6686), .ZN(n6690) );
  INV_X1 U8421 ( .A(n6688), .ZN(n6689) );
  OAI22_X1 U8422 ( .A1(n6690), .A2(n6689), .B1(n9165), .B2(n9105), .ZN(n6691)
         );
  NAND2_X1 U8423 ( .A1(n6691), .A2(n6706), .ZN(n6692) );
  NAND2_X1 U8424 ( .A1(n6692), .A2(n6700), .ZN(n6693) );
  AOI21_X1 U8425 ( .B1(n6693), .B2(n6708), .A(n7702), .ZN(n6698) );
  INV_X1 U8426 ( .A(n6693), .ZN(n6696) );
  NAND2_X1 U8427 ( .A1(n6696), .A2(n6695), .ZN(n6697) );
  NAND2_X1 U8428 ( .A1(n6699), .A2(n4909), .ZN(n6714) );
  INV_X1 U8429 ( .A(n6700), .ZN(n6702) );
  NOR2_X1 U8430 ( .A1(n7702), .A2(n6704), .ZN(n6709) );
  INV_X1 U8431 ( .A(n6840), .ZN(n6705) );
  OAI211_X1 U8432 ( .C1(n6706), .C2(n7232), .A(n6709), .B(n6705), .ZN(n6713)
         );
  INV_X1 U8433 ( .A(n7266), .ZN(n7265) );
  INV_X1 U8434 ( .A(n6707), .ZN(n8987) );
  NAND4_X1 U8435 ( .A1(n8928), .A2(n7265), .A3(n8987), .A4(n6708), .ZN(n6711)
         );
  INV_X1 U8436 ( .A(n6709), .ZN(n6710) );
  NAND3_X1 U8437 ( .A1(n6711), .A2(P1_B_REG_SCAN_IN), .A3(n6710), .ZN(n6712)
         );
  AOI21_X1 U8438 ( .B1(n8925), .B2(n6717), .A(n6716), .ZN(n6719) );
  OAI21_X1 U8439 ( .B1(n6719), .B2(n6718), .A(n8941), .ZN(n6728) );
  INV_X1 U8440 ( .A(n9521), .ZN(n9200) );
  INV_X1 U8441 ( .A(n6720), .ZN(n9197) );
  NAND2_X1 U8442 ( .A1(n8955), .A2(n8929), .ZN(n6722) );
  NAND2_X1 U8443 ( .A1(n8957), .A2(n8928), .ZN(n6721) );
  AND2_X1 U8444 ( .A1(n6722), .A2(n6721), .ZN(n9194) );
  OAI22_X1 U8445 ( .A1(n9194), .A2(n8918), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6723), .ZN(n6724) );
  AOI21_X1 U8446 ( .B1(n9197), .B2(n8921), .A(n6724), .ZN(n6725) );
  INV_X1 U8447 ( .A(n6726), .ZN(n6727) );
  NAND2_X1 U8448 ( .A1(n6728), .A2(n6727), .ZN(P1_U3214) );
  INV_X1 U8449 ( .A(n6729), .ZN(n6730) );
  OR2_X2 U8450 ( .A1(n6731), .A2(n6730), .ZN(n8974) );
  INV_X1 U8451 ( .A(n8974), .ZN(P1_U3973) );
  NOR2_X1 U8452 ( .A1(n4425), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9588) );
  INV_X1 U8453 ( .A(n9588), .ZN(n8064) );
  OAI222_X1 U8454 ( .A1(n8064), .A2(n6732), .B1(n9590), .B2(n6746), .C1(n6789), 
        .C2(P1_U3086), .ZN(P1_U3353) );
  OAI222_X1 U8455 ( .A1(P1_U3086), .A2(n6790), .B1(n8064), .B2(n6733), .C1(
        n9590), .C2(n6740), .ZN(P1_U3354) );
  OAI222_X1 U8456 ( .A1(n8064), .A2(n6734), .B1(n9590), .B2(n6737), .C1(n6793), 
        .C2(P1_U3086), .ZN(P1_U3352) );
  OAI222_X1 U8457 ( .A1(n8064), .A2(n9416), .B1(n9590), .B2(n6738), .C1(n6795), 
        .C2(P1_U3086), .ZN(P1_U3351) );
  AND2_X1 U8458 ( .A1(n4425), .A2(P2_U3151), .ZN(n8818) );
  INV_X1 U8459 ( .A(n8818), .ZN(n8824) );
  OAI222_X1 U8460 ( .A1(n8824), .A2(n9302), .B1(n8822), .B2(n6737), .C1(
        P2_U3151), .C2(n6922), .ZN(P2_U3292) );
  OAI222_X1 U8461 ( .A1(n8824), .A2(n6739), .B1(n8822), .B2(n6738), .C1(
        P2_U3151), .C2(n6972), .ZN(P2_U3291) );
  OAI222_X1 U8462 ( .A1(n6952), .A2(P2_U3151), .B1(n8824), .B2(n6741), .C1(
        n8822), .C2(n6740), .ZN(P2_U3294) );
  INV_X1 U8463 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6742) );
  INV_X1 U8464 ( .A(n6797), .ZN(n9706) );
  OAI222_X1 U8465 ( .A1(n8064), .A2(n6742), .B1(n9590), .B2(n6748), .C1(n9706), 
        .C2(P1_U3086), .ZN(P1_U3350) );
  OAI222_X1 U8466 ( .A1(P2_U3151), .A2(n7115), .B1(n8822), .B2(n6744), .C1(
        n6743), .C2(n8824), .ZN(P2_U3289) );
  INV_X1 U8467 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6745) );
  INV_X1 U8468 ( .A(n6801), .ZN(n9723) );
  OAI222_X1 U8469 ( .A1(n8064), .A2(n6745), .B1(n9590), .B2(n6744), .C1(n9723), 
        .C2(P1_U3086), .ZN(P1_U3349) );
  OAI222_X1 U8470 ( .A1(n8824), .A2(n4523), .B1(n8822), .B2(n6746), .C1(
        P2_U3151), .C2(n7049), .ZN(P2_U3293) );
  OAI222_X1 U8471 ( .A1(P2_U3151), .A2(n6749), .B1(n8822), .B2(n6748), .C1(
        n6747), .C2(n8824), .ZN(P2_U3290) );
  OAI222_X1 U8472 ( .A1(P2_U3151), .A2(n7178), .B1(n8822), .B2(n6750), .C1(
        n4424), .C2(n8824), .ZN(P2_U3288) );
  INV_X1 U8473 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6751) );
  INV_X1 U8474 ( .A(n6803), .ZN(n9618) );
  OAI222_X1 U8475 ( .A1(n8064), .A2(n6751), .B1(n9590), .B2(n6750), .C1(n9618), 
        .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U8476 ( .A(n6752), .ZN(n6753) );
  OR2_X1 U8477 ( .A1(n6835), .A2(n6753), .ZN(n6754) );
  AND2_X1 U8478 ( .A1(n6755), .A2(n6754), .ZN(n6761) );
  NAND2_X1 U8479 ( .A1(n7266), .A2(n7702), .ZN(n6760) );
  INV_X1 U8480 ( .A(n6760), .ZN(n6756) );
  INV_X1 U8481 ( .A(n9805), .ZN(n9064) );
  NOR2_X1 U8482 ( .A1(n9064), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8483 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9398) );
  INV_X1 U8484 ( .A(n6757), .ZN(n6759) );
  INV_X1 U8485 ( .A(n6806), .ZN(n9635) );
  OAI222_X1 U8486 ( .A1(n8064), .A2(n9398), .B1(n9590), .B2(n6759), .C1(
        P1_U3086), .C2(n9635), .ZN(P1_U3347) );
  INV_X1 U8487 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6758) );
  OAI222_X1 U8488 ( .A1(n7247), .A2(P2_U3151), .B1(n8822), .B2(n6759), .C1(
        n6758), .C2(n8824), .ZN(P2_U3287) );
  AND2_X1 U8489 ( .A1(n6761), .A2(n6760), .ZN(n6809) );
  INV_X1 U8490 ( .A(n6809), .ZN(n6766) );
  AOI21_X1 U8491 ( .B1(n8987), .B2(n7340), .A(n4267), .ZN(n8993) );
  OAI21_X1 U8492 ( .B1(n8987), .B2(P1_REG1_REG_0__SCAN_IN), .A(n8993), .ZN(
        n6763) );
  XNOR2_X1 U8493 ( .A(n6763), .B(n6762), .ZN(n6765) );
  AOI22_X1 U8494 ( .A1(n9064), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n6764) );
  OAI21_X1 U8495 ( .B1(n6766), .B2(n6765), .A(n6764), .ZN(P1_U3243) );
  INV_X1 U8496 ( .A(n6767), .ZN(n6770) );
  OAI222_X1 U8497 ( .A1(P2_U3151), .A2(n6769), .B1(n8822), .B2(n6770), .C1(
        n6768), .C2(n8824), .ZN(P2_U3286) );
  INV_X1 U8498 ( .A(n6876), .ZN(n6811) );
  OAI222_X1 U8499 ( .A1(n8064), .A2(n6771), .B1(n9590), .B2(n6770), .C1(n6811), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8500 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6772) );
  INV_X1 U8501 ( .A(n9602), .ZN(n6869) );
  OAI222_X1 U8502 ( .A1(n8064), .A2(n6772), .B1(n9590), .B2(n6774), .C1(n6869), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U8503 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6773) );
  OAI222_X1 U8504 ( .A1(P2_U3151), .A2(n6775), .B1(n8822), .B2(n6774), .C1(
        n6773), .C2(n8824), .ZN(P2_U3285) );
  INV_X1 U8505 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n9312) );
  NOR2_X1 U8506 ( .A1(n6825), .A2(n9312), .ZN(P2_U3242) );
  NOR2_X1 U8507 ( .A1(n6876), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6776) );
  AOI21_X1 U8508 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6876), .A(n6776), .ZN(
        n6785) );
  INV_X1 U8509 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6777) );
  MUX2_X1 U8510 ( .A(n6777), .B(P1_REG2_REG_2__SCAN_IN), .S(n6789), .Z(n8999)
         );
  INV_X1 U8511 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7522) );
  MUX2_X1 U8512 ( .A(n7522), .B(P1_REG2_REG_1__SCAN_IN), .S(n6790), .Z(n8983)
         );
  AND2_X1 U8513 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n8988) );
  INV_X1 U8514 ( .A(n6790), .ZN(n8978) );
  NAND2_X1 U8515 ( .A1(n8978), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U8516 ( .A1(n8982), .A2(n6778), .ZN(n8998) );
  NAND2_X1 U8517 ( .A1(n8999), .A2(n8998), .ZN(n8997) );
  INV_X1 U8518 ( .A(n6789), .ZN(n8996) );
  NAND2_X1 U8519 ( .A1(n8996), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6779) );
  NAND2_X1 U8520 ( .A1(n8997), .A2(n6779), .ZN(n9012) );
  INV_X1 U8521 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9431) );
  MUX2_X1 U8522 ( .A(n9431), .B(P1_REG2_REG_3__SCAN_IN), .S(n6793), .Z(n9013)
         );
  INV_X1 U8523 ( .A(n6793), .ZN(n9010) );
  NAND2_X1 U8524 ( .A1(n9010), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6780) );
  NAND2_X1 U8525 ( .A1(n9011), .A2(n6780), .ZN(n9027) );
  XNOR2_X1 U8526 ( .A(n6795), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U8527 ( .A1(n9027), .A2(n9028), .ZN(n9026) );
  INV_X1 U8528 ( .A(n6795), .ZN(n9022) );
  NAND2_X1 U8529 ( .A1(n9022), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6781) );
  NAND2_X1 U8530 ( .A1(n9026), .A2(n6781), .ZN(n9700) );
  MUX2_X1 U8531 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7298), .S(n6797), .Z(n9699)
         );
  AND2_X1 U8532 ( .A1(n9700), .A2(n9699), .ZN(n9702) );
  NAND2_X1 U8533 ( .A1(n6801), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6782) );
  OAI21_X1 U8534 ( .B1(n6801), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6782), .ZN(
        n9716) );
  NOR2_X1 U8535 ( .A1(n9715), .A2(n9716), .ZN(n9717) );
  AOI21_X1 U8536 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6801), .A(n9717), .ZN(
        n9612) );
  AOI22_X1 U8537 ( .A1(n6803), .A2(n5830), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n9618), .ZN(n9611) );
  NOR2_X1 U8538 ( .A1(n9612), .A2(n9611), .ZN(n9610) );
  NAND2_X1 U8539 ( .A1(n6806), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6783) );
  OAI21_X1 U8540 ( .B1(n6806), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6783), .ZN(
        n9628) );
  NOR2_X1 U8541 ( .A1(n9627), .A2(n9628), .ZN(n9629) );
  AOI21_X1 U8542 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6806), .A(n9629), .ZN(
        n6784) );
  NAND2_X1 U8543 ( .A1(n6785), .A2(n6784), .ZN(n6870) );
  OAI21_X1 U8544 ( .B1(n6785), .B2(n6784), .A(n6870), .ZN(n6787) );
  NOR2_X1 U8545 ( .A1(n4267), .A2(n6707), .ZN(n6786) );
  NAND2_X1 U8546 ( .A1(n6809), .A2(n6786), .ZN(n9795) );
  INV_X1 U8547 ( .A(n9795), .ZN(n9086) );
  NAND2_X1 U8548 ( .A1(n6787), .A2(n9086), .ZN(n6815) );
  NOR2_X1 U8549 ( .A1(n6876), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6788) );
  AOI21_X1 U8550 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n6876), .A(n6788), .ZN(
        n6808) );
  MUX2_X1 U8551 ( .A(n5720), .B(P1_REG1_REG_2__SCAN_IN), .S(n6789), .Z(n9003)
         );
  MUX2_X1 U8552 ( .A(n5683), .B(P1_REG1_REG_1__SCAN_IN), .S(n6790), .Z(n8981)
         );
  AND2_X1 U8553 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n8980) );
  NAND2_X1 U8554 ( .A1(n8981), .A2(n8980), .ZN(n8979) );
  NAND2_X1 U8555 ( .A1(n8978), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6791) );
  NAND2_X1 U8556 ( .A1(n8979), .A2(n6791), .ZN(n9002) );
  NAND2_X1 U8557 ( .A1(n9003), .A2(n9002), .ZN(n9001) );
  NAND2_X1 U8558 ( .A1(n8996), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6792) );
  NAND2_X1 U8559 ( .A1(n9001), .A2(n6792), .ZN(n9015) );
  MUX2_X1 U8560 ( .A(n5740), .B(P1_REG1_REG_3__SCAN_IN), .S(n6793), .Z(n9016)
         );
  NAND2_X1 U8561 ( .A1(n9015), .A2(n9016), .ZN(n9014) );
  NAND2_X1 U8562 ( .A1(n9010), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6794) );
  NAND2_X1 U8563 ( .A1(n9014), .A2(n6794), .ZN(n9024) );
  XNOR2_X1 U8564 ( .A(n6795), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9025) );
  NAND2_X1 U8565 ( .A1(n9024), .A2(n9025), .ZN(n9023) );
  NAND2_X1 U8566 ( .A1(n9022), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6796) );
  NAND2_X1 U8567 ( .A1(n9023), .A2(n6796), .ZN(n9697) );
  OR2_X1 U8568 ( .A1(n6797), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6798) );
  NAND2_X1 U8569 ( .A1(n6797), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6799) );
  AND2_X1 U8570 ( .A1(n6798), .A2(n6799), .ZN(n9698) );
  NAND2_X1 U8571 ( .A1(n9697), .A2(n9698), .ZN(n9696) );
  AND2_X1 U8572 ( .A1(n9696), .A2(n6799), .ZN(n9713) );
  NAND2_X1 U8573 ( .A1(n6801), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6800) );
  OAI21_X1 U8574 ( .B1(n6801), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6800), .ZN(
        n9712) );
  NOR2_X1 U8575 ( .A1(n9713), .A2(n9712), .ZN(n9711) );
  AOI21_X1 U8576 ( .B1(n6801), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9711), .ZN(
        n9607) );
  INV_X1 U8577 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6802) );
  MUX2_X1 U8578 ( .A(n6802), .B(P1_REG1_REG_7__SCAN_IN), .S(n6803), .Z(n9608)
         );
  NOR2_X1 U8579 ( .A1(n9607), .A2(n9608), .ZN(n9606) );
  AOI21_X1 U8580 ( .B1(n6803), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9606), .ZN(
        n9624) );
  OR2_X1 U8581 ( .A1(n6806), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6805) );
  NAND2_X1 U8582 ( .A1(n6806), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U8583 ( .A1(n6805), .A2(n6804), .ZN(n9625) );
  NOR2_X1 U8584 ( .A1(n9624), .A2(n9625), .ZN(n9623) );
  AOI21_X1 U8585 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6806), .A(n9623), .ZN(
        n6807) );
  NAND2_X1 U8586 ( .A1(n6808), .A2(n6807), .ZN(n6875) );
  OAI21_X1 U8587 ( .B1(n6808), .B2(n6807), .A(n6875), .ZN(n6813) );
  NAND2_X1 U8588 ( .A1(n6809), .A2(n4267), .ZN(n9773) );
  NAND2_X1 U8589 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7676) );
  NAND2_X1 U8590 ( .A1(n9064), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n6810) );
  OAI211_X1 U8591 ( .C1(n9773), .C2(n6811), .A(n7676), .B(n6810), .ZN(n6812)
         );
  AOI21_X1 U8592 ( .B1(n6813), .B2(n9763), .A(n6812), .ZN(n6814) );
  NAND2_X1 U8593 ( .A1(n6815), .A2(n6814), .ZN(P1_U3252) );
  INV_X1 U8594 ( .A(n6816), .ZN(n6819) );
  AOI22_X1 U8595 ( .A1(n9728), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9588), .ZN(n6817) );
  OAI21_X1 U8596 ( .B1(n6819), .B2(n9590), .A(n6817), .ZN(P1_U3344) );
  INV_X1 U8597 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6818) );
  OAI222_X1 U8598 ( .A1(n6820), .A2(P2_U3151), .B1(n8822), .B2(n6819), .C1(
        n6818), .C2(n8824), .ZN(P2_U3284) );
  AND2_X1 U8599 ( .A1(n7919), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8600 ( .A1(n7919), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8601 ( .A1(n7919), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8602 ( .A1(n7919), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8603 ( .A1(n7919), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8604 ( .A1(n7919), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8605 ( .A1(n7919), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8606 ( .A1(n7919), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8607 ( .A1(n7919), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8608 ( .A1(n7919), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8609 ( .A1(n7919), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8610 ( .A1(n7919), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  INV_X1 U8611 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6821) );
  INV_X1 U8612 ( .A(n9045), .ZN(n6884) );
  OAI222_X1 U8613 ( .A1(n8064), .A2(n6821), .B1(n9590), .B2(n6823), .C1(n6884), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8614 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6822) );
  OAI222_X1 U8615 ( .A1(P2_U3151), .A2(n6824), .B1(n8822), .B2(n6823), .C1(
        n6822), .C2(n8824), .ZN(P2_U3283) );
  INV_X1 U8616 ( .A(n6826), .ZN(n6827) );
  AOI22_X1 U8617 ( .A1(n7919), .A2(n5588), .B1(n7118), .B2(n6827), .ZN(
        P2_U3376) );
  AND2_X1 U8618 ( .A1(n7919), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8619 ( .A1(n7919), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8620 ( .A1(n7919), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8621 ( .A1(n7919), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8622 ( .A1(n7919), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8623 ( .A1(n7919), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8624 ( .A1(n7919), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8625 ( .A1(n7919), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8626 ( .A1(n7919), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8627 ( .A1(n7919), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8628 ( .A1(n7919), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8629 ( .A1(n7919), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8630 ( .A1(n7919), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8631 ( .A1(n7919), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8632 ( .A1(n7919), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8633 ( .A1(n7919), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8634 ( .A1(n7919), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  INV_X1 U8635 ( .A(n6828), .ZN(n6831) );
  AOI22_X1 U8636 ( .A1(n9754), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9588), .ZN(n6829) );
  OAI21_X1 U8637 ( .B1(n6831), .B2(n9590), .A(n6829), .ZN(P1_U3342) );
  AOI22_X1 U8638 ( .A1(n7869), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n8818), .ZN(n6830) );
  OAI21_X1 U8639 ( .B1(n6831), .B2(n8822), .A(n6830), .ZN(P2_U3282) );
  INV_X1 U8640 ( .A(n7332), .ZN(n6842) );
  NAND2_X1 U8641 ( .A1(n8973), .A2(n8929), .ZN(n7335) );
  INV_X1 U8642 ( .A(n7335), .ZN(n6854) );
  NAND2_X1 U8643 ( .A1(n6834), .A2(n6832), .ZN(n6833) );
  AND2_X1 U8644 ( .A1(n7332), .A2(n6833), .ZN(n6836) );
  OR2_X1 U8645 ( .A1(n6835), .A2(n6834), .ZN(n7333) );
  NAND2_X1 U8646 ( .A1(n6836), .A2(n7333), .ZN(n7521) );
  OR2_X1 U8647 ( .A1(n6838), .A2(n6837), .ZN(n9904) );
  OR2_X1 U8648 ( .A1(n7232), .A2(n7587), .ZN(n6839) );
  AOI21_X1 U8649 ( .B1(n9937), .B2(n9828), .A(n7331), .ZN(n6841) );
  AOI211_X1 U8650 ( .C1(n6842), .C2(n7330), .A(n6854), .B(n6841), .ZN(n9903)
         );
  AND2_X1 U8651 ( .A1(n7265), .A2(n7268), .ZN(n6849) );
  OAI21_X1 U8652 ( .B1(n7264), .B2(P1_D_REG_1__SCAN_IN), .A(n9583), .ZN(n6848)
         );
  INV_X1 U8653 ( .A(n7264), .ZN(n6845) );
  INV_X1 U8654 ( .A(n6843), .ZN(n6844) );
  NAND2_X1 U8655 ( .A1(n6845), .A2(n6844), .ZN(n6847) );
  OR2_X1 U8656 ( .A1(n9481), .A2(n7232), .ZN(n6846) );
  NAND4_X1 U8657 ( .A1(n6849), .A2(n6848), .A3(n6847), .A4(n6846), .ZN(n7306)
         );
  NAND2_X1 U8658 ( .A1(n10006), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6850) );
  OAI21_X1 U8659 ( .B1(n9903), .B2(n10006), .A(n6850), .ZN(P1_U3522) );
  AOI22_X1 U8660 ( .A1(n9758), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9588), .ZN(n6851) );
  OAI21_X1 U8661 ( .B1(n6858), .B2(n9590), .A(n6851), .ZN(P1_U3341) );
  XNOR2_X1 U8662 ( .A(n6853), .B(n6852), .ZN(n8989) );
  AOI22_X1 U8663 ( .A1(n8934), .A2(n7330), .B1(n8948), .B2(n6854), .ZN(n6856)
         );
  NOR2_X1 U8664 ( .A1(n8921), .A2(P1_U3086), .ZN(n6907) );
  INV_X1 U8665 ( .A(n6907), .ZN(n6865) );
  NAND2_X1 U8666 ( .A1(n6865), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6855) );
  OAI211_X1 U8667 ( .C1(n8989), .C2(n8923), .A(n6856), .B(n6855), .ZN(P1_U3232) );
  INV_X1 U8668 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6857) );
  OAI222_X1 U8669 ( .A1(P2_U3151), .A2(n6859), .B1(n8822), .B2(n6858), .C1(
        n6857), .C2(n8824), .ZN(P2_U3281) );
  AOI22_X1 U8670 ( .A1(n8497), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n8818), .ZN(n6860) );
  OAI21_X1 U8671 ( .B1(n6895), .B2(n8822), .A(n6860), .ZN(P2_U3280) );
  INV_X1 U8672 ( .A(n6863), .ZN(n6900) );
  AOI21_X1 U8673 ( .B1(n6861), .B2(n6862), .A(n6900), .ZN(n6867) );
  AOI22_X1 U8674 ( .A1(n8928), .A2(n8975), .B1(n8972), .B2(n8929), .ZN(n7520)
         );
  OAI22_X1 U8675 ( .A1(n9907), .A2(n8951), .B1(n7520), .B2(n8918), .ZN(n6864)
         );
  AOI21_X1 U8676 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6865), .A(n6864), .ZN(
        n6866) );
  OAI21_X1 U8677 ( .B1(n6867), .B2(n8923), .A(n6866), .ZN(P1_U3222) );
  NOR2_X1 U8678 ( .A1(n9045), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6868) );
  AOI21_X1 U8679 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9045), .A(n6868), .ZN(
        n6873) );
  AOI22_X1 U8680 ( .A1(n9602), .A2(n7507), .B1(P1_REG2_REG_10__SCAN_IN), .B2(
        n6869), .ZN(n9598) );
  OAI21_X1 U8681 ( .B1(n6876), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6870), .ZN(
        n9599) );
  NOR2_X1 U8682 ( .A1(n9598), .A2(n9599), .ZN(n9597) );
  NAND2_X1 U8683 ( .A1(n9728), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6871) );
  OAI21_X1 U8684 ( .B1(n9728), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6871), .ZN(
        n9734) );
  NOR2_X1 U8685 ( .A1(n9733), .A2(n9734), .ZN(n9735) );
  AOI21_X1 U8686 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9728), .A(n9735), .ZN(
        n6872) );
  NAND2_X1 U8687 ( .A1(n6873), .A2(n6872), .ZN(n9044) );
  OAI21_X1 U8688 ( .B1(n6873), .B2(n6872), .A(n9044), .ZN(n6886) );
  MUX2_X1 U8689 ( .A(n6874), .B(P1_REG1_REG_10__SCAN_IN), .S(n9602), .Z(n9595)
         );
  OAI21_X1 U8690 ( .B1(n6876), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6875), .ZN(
        n9596) );
  NOR2_X1 U8691 ( .A1(n9595), .A2(n9596), .ZN(n9594) );
  AOI21_X1 U8692 ( .B1(n9602), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9594), .ZN(
        n9730) );
  MUX2_X1 U8693 ( .A(n6877), .B(P1_REG1_REG_11__SCAN_IN), .S(n9728), .Z(n9731)
         );
  NOR2_X1 U8694 ( .A1(n9730), .A2(n9731), .ZN(n9729) );
  AOI21_X1 U8695 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9728), .A(n9729), .ZN(
        n6879) );
  AOI22_X1 U8696 ( .A1(n9045), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n5941), .B2(
        n6884), .ZN(n6878) );
  NAND2_X1 U8697 ( .A1(n6879), .A2(n6878), .ZN(n9034) );
  OAI21_X1 U8698 ( .B1(n6879), .B2(n6878), .A(n9034), .ZN(n6880) );
  NAND2_X1 U8699 ( .A1(n6880), .A2(n9763), .ZN(n6883) );
  NOR2_X1 U8700 ( .A1(n6881), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7774) );
  AOI21_X1 U8701 ( .B1(n9064), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n7774), .ZN(
        n6882) );
  OAI211_X1 U8702 ( .C1(n9773), .C2(n6884), .A(n6883), .B(n6882), .ZN(n6885)
         );
  AOI21_X1 U8703 ( .B1(n6886), .B2(n9086), .A(n6885), .ZN(n6887) );
  INV_X1 U8704 ( .A(n6887), .ZN(P1_U3255) );
  INV_X1 U8705 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6892) );
  OAI21_X1 U8706 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6888), .A(n6935), .ZN(n6889) );
  OAI21_X1 U8707 ( .B1(n10031), .B2(n6890), .A(n6889), .ZN(n6891) );
  OAI21_X1 U8708 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6892), .A(n6891), .ZN(n6893) );
  AOI21_X1 U8709 ( .B1(n7807), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n6893), .ZN(
        n6894) );
  OAI21_X1 U8710 ( .B1(n4885), .B2(n10012), .A(n6894), .ZN(P2_U3182) );
  INV_X1 U8711 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6896) );
  OAI222_X1 U8712 ( .A1(n8064), .A2(n6896), .B1(n9590), .B2(n6895), .C1(n9048), 
        .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U8713 ( .A(n6897), .ZN(n6899) );
  NOR3_X1 U8714 ( .A1(n6900), .A2(n6899), .A3(n6898), .ZN(n6903) );
  INV_X1 U8715 ( .A(n6901), .ZN(n6902) );
  OAI21_X1 U8716 ( .B1(n6903), .B2(n6902), .A(n8941), .ZN(n6906) );
  INV_X1 U8717 ( .A(n8928), .ZN(n9167) );
  OAI22_X1 U8718 ( .A1(n7288), .A2(n7569), .B1(n6904), .B2(n9167), .ZN(n9875)
         );
  AOI22_X1 U8719 ( .A1(n8934), .A2(n4269), .B1(n9875), .B2(n8948), .ZN(n6905)
         );
  OAI211_X1 U8720 ( .C1(n6907), .C2(n9878), .A(n6906), .B(n6905), .ZN(P1_U3237) );
  OAI21_X1 U8721 ( .B1(n6910), .B2(n6909), .A(n6908), .ZN(n6911) );
  NAND2_X1 U8722 ( .A1(n6911), .A2(n10031), .ZN(n6921) );
  INV_X1 U8723 ( .A(n10020), .ZN(n7180) );
  OAI21_X1 U8724 ( .B1(n6913), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6912), .ZN(
        n6919) );
  AND2_X1 U8725 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7018) );
  INV_X1 U8726 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6917) );
  INV_X1 U8727 ( .A(n6960), .ZN(n6915) );
  AOI21_X1 U8728 ( .B1(n4741), .B2(n4739), .A(n6915), .ZN(n6916) );
  OAI22_X1 U8729 ( .A1(n10010), .A2(n6917), .B1(n10026), .B2(n6916), .ZN(n6918) );
  AOI211_X1 U8730 ( .C1(n7180), .C2(n6919), .A(n7018), .B(n6918), .ZN(n6920)
         );
  OAI211_X1 U8731 ( .C1(n10012), .C2(n6922), .A(n6921), .B(n6920), .ZN(
        P2_U3185) );
  MUX2_X1 U8732 ( .A(n6977), .B(n6924), .S(n6923), .Z(n6926) );
  NAND2_X1 U8733 ( .A1(n6926), .A2(n6925), .ZN(n6929) );
  INV_X1 U8734 ( .A(n10040), .ZN(n6980) );
  AND2_X1 U8735 ( .A1(n8464), .A2(n6980), .ZN(n8218) );
  INV_X1 U8736 ( .A(n8218), .ZN(n8219) );
  NAND2_X1 U8737 ( .A1(n8219), .A2(n8217), .ZN(n10035) );
  NOR2_X1 U8738 ( .A1(n6984), .A2(n8695), .ZN(n10039) );
  AOI21_X1 U8739 ( .B1(n6928), .B2(n10035), .A(n10039), .ZN(n6933) );
  INV_X1 U8740 ( .A(n6929), .ZN(n6930) );
  INV_X1 U8741 ( .A(n8588), .ZN(n7747) );
  NAND2_X1 U8742 ( .A1(n6930), .A2(n7747), .ZN(n8545) );
  AOI22_X1 U8743 ( .A1(n8702), .A2(n10040), .B1(n8701), .B2(
        P2_REG2_REG_0__SCAN_IN), .ZN(n6932) );
  NAND2_X1 U8744 ( .A1(n8685), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6931) );
  OAI211_X1 U8745 ( .C1(n8701), .C2(n6933), .A(n6932), .B(n6931), .ZN(P2_U3233) );
  AOI22_X1 U8746 ( .A1(n8517), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n8818), .ZN(n6934) );
  OAI21_X1 U8747 ( .B1(n6953), .B2(n8822), .A(n6934), .ZN(P2_U3279) );
  OAI21_X1 U8748 ( .B1(n6936), .B2(n6935), .A(n10031), .ZN(n6939) );
  INV_X1 U8749 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6937) );
  OAI22_X1 U8750 ( .A1(n6939), .A2(n6938), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6937), .ZN(n6950) );
  AOI21_X1 U8751 ( .B1(n6942), .B2(n6941), .A(n6940), .ZN(n6948) );
  INV_X1 U8752 ( .A(n6943), .ZN(n6944) );
  AOI21_X1 U8753 ( .B1(n6946), .B2(n6945), .A(n6944), .ZN(n6947) );
  OAI22_X1 U8754 ( .A1(n6948), .A2(n10020), .B1(n10026), .B2(n6947), .ZN(n6949) );
  AOI211_X1 U8755 ( .C1(n7807), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n6950), .B(
        n6949), .ZN(n6951) );
  OAI21_X1 U8756 ( .B1(n6952), .B2(n10012), .A(n6951), .ZN(P2_U3183) );
  INV_X1 U8757 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6954) );
  INV_X1 U8758 ( .A(n9059), .ZN(n9042) );
  OAI222_X1 U8759 ( .A1(n8064), .A2(n6954), .B1(n9590), .B2(n6953), .C1(n9042), 
        .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U8760 ( .A(n10031), .ZN(n7252) );
  AOI211_X1 U8761 ( .C1(n6957), .C2(n6956), .A(n7252), .B(n6955), .ZN(n6958)
         );
  INV_X1 U8762 ( .A(n6958), .ZN(n6971) );
  NAND3_X1 U8763 ( .A1(n6960), .A2(n4414), .A3(n6959), .ZN(n6961) );
  AOI21_X1 U8764 ( .B1(n6962), .B2(n6961), .A(n10026), .ZN(n6969) );
  AND3_X1 U8765 ( .A1(n6912), .A2(n6964), .A3(n6963), .ZN(n6965) );
  OAI21_X1 U8766 ( .B1(n6966), .B2(n6965), .A(n7180), .ZN(n6967) );
  NAND2_X1 U8767 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7069) );
  NAND2_X1 U8768 ( .A1(n6967), .A2(n7069), .ZN(n6968) );
  AOI211_X1 U8769 ( .C1(n7807), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6969), .B(
        n6968), .ZN(n6970) );
  OAI211_X1 U8770 ( .C1(n10012), .C2(n6972), .A(n6971), .B(n6970), .ZN(
        P2_U3186) );
  INV_X1 U8771 ( .A(n6973), .ZN(n6976) );
  INV_X1 U8772 ( .A(n8383), .ZN(n6975) );
  INV_X1 U8773 ( .A(n8426), .ZN(n6974) );
  NAND2_X2 U8774 ( .A1(n6978), .A2(n6977), .ZN(n6990) );
  CLKBUF_X1 U8775 ( .A(n6990), .Z(n6981) );
  XNOR2_X1 U8776 ( .A(n6981), .B(n6979), .ZN(n6988) );
  XNOR2_X1 U8777 ( .A(n6988), .B(n8462), .ZN(n7125) );
  AND2_X1 U8778 ( .A1(n6982), .A2(n8217), .ZN(n7117) );
  XNOR2_X2 U8779 ( .A(n6990), .B(n6983), .ZN(n6986) );
  XNOR2_X2 U8780 ( .A(n6986), .B(n6984), .ZN(n7116) );
  INV_X1 U8781 ( .A(n6986), .ZN(n6987) );
  INV_X2 U8782 ( .A(n6990), .ZN(n7363) );
  XNOR2_X1 U8783 ( .A(n7082), .B(n7367), .ZN(n7066) );
  XNOR2_X1 U8784 ( .A(n7066), .B(n8461), .ZN(n6996) );
  NAND2_X1 U8785 ( .A1(n6997), .A2(n6996), .ZN(n7065) );
  INV_X1 U8786 ( .A(n7005), .ZN(n6991) );
  NAND2_X1 U8787 ( .A1(n7013), .A2(n6991), .ZN(n6995) );
  INV_X1 U8788 ( .A(n6992), .ZN(n6993) );
  NAND2_X1 U8789 ( .A1(n7016), .A2(n6993), .ZN(n6994) );
  OAI211_X1 U8790 ( .C1(n6997), .C2(n6996), .A(n7065), .B(n8185), .ZN(n7023)
         );
  AND2_X1 U8791 ( .A1(n6999), .A2(n6998), .ZN(n7004) );
  OAI21_X1 U8792 ( .B1(n7002), .B2(n7001), .A(n7000), .ZN(n7003) );
  OAI211_X1 U8793 ( .C1(n7009), .C2(n7005), .A(n7004), .B(n7003), .ZN(n7006)
         );
  NAND2_X1 U8794 ( .A1(n7006), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7011) );
  INV_X1 U8795 ( .A(n7007), .ZN(n8436) );
  NAND2_X1 U8796 ( .A1(n8437), .A2(n8436), .ZN(n7008) );
  OR2_X1 U8797 ( .A1(n7009), .A2(n7008), .ZN(n7010) );
  AND2_X1 U8798 ( .A1(n7011), .A2(n7010), .ZN(n7119) );
  OR2_X1 U8799 ( .A1(n7012), .A2(P2_U3151), .ZN(n8441) );
  NAND2_X1 U8800 ( .A1(n7013), .A2(n8436), .ZN(n7014) );
  INV_X1 U8801 ( .A(n7014), .ZN(n7015) );
  NAND2_X1 U8802 ( .A1(n8200), .A2(n8460), .ZN(n7020) );
  NAND2_X1 U8803 ( .A1(n7016), .A2(n10066), .ZN(n7017) );
  AOI21_X1 U8804 ( .B1(n8176), .B2(n7225), .A(n7018), .ZN(n7019) );
  OAI211_X1 U8805 ( .C1(n4987), .C2(n8202), .A(n7020), .B(n7019), .ZN(n7021)
         );
  AOI21_X1 U8806 ( .B1(n7224), .B2(n8204), .A(n7021), .ZN(n7022) );
  NAND2_X1 U8807 ( .A1(n7023), .A2(n7022), .ZN(P2_U3158) );
  AND2_X1 U8808 ( .A1(n7024), .A2(n7025), .ZN(n7028) );
  OAI211_X1 U8809 ( .C1(n7028), .C2(n7027), .A(n8941), .B(n7026), .ZN(n7032)
         );
  OAI22_X1 U8810 ( .A1(n7288), .A2(n9167), .B1(n7312), .B2(n7569), .ZN(n9861)
         );
  INV_X1 U8811 ( .A(n9861), .ZN(n7029) );
  INV_X1 U8812 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9309) );
  OAI22_X1 U8813 ( .A1(n7029), .A2(n8918), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9309), .ZN(n7030) );
  AOI21_X1 U8814 ( .B1(n7299), .B2(n8934), .A(n7030), .ZN(n7031) );
  OAI211_X1 U8815 ( .C1(n8944), .C2(n9863), .A(n7032), .B(n7031), .ZN(P1_U3230) );
  AOI211_X1 U8816 ( .C1(n7035), .C2(n7034), .A(n7252), .B(n7033), .ZN(n7047)
         );
  AOI21_X1 U8817 ( .B1(n7038), .B2(n7037), .A(n7036), .ZN(n7045) );
  INV_X1 U8818 ( .A(n10026), .ZN(n7183) );
  OAI21_X1 U8819 ( .B1(n7041), .B2(n7040), .A(n7039), .ZN(n7042) );
  AOI22_X1 U8820 ( .A1(n7807), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n7183), .B2(
        n7042), .ZN(n7044) );
  NAND2_X1 U8821 ( .A1(P2_U3151), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7043) );
  OAI211_X1 U8822 ( .C1(n7045), .C2(n10020), .A(n7044), .B(n7043), .ZN(n7046)
         );
  NOR2_X1 U8823 ( .A1(n7047), .A2(n7046), .ZN(n7048) );
  OAI21_X1 U8824 ( .B1(n7049), .B2(n10012), .A(n7048), .ZN(P2_U3184) );
  INV_X1 U8825 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7053) );
  INV_X1 U8826 ( .A(n7050), .ZN(n7052) );
  INV_X1 U8827 ( .A(n7107), .ZN(n7051) );
  AOI21_X1 U8828 ( .B1(n7053), .B2(n7052), .A(n7051), .ZN(n7057) );
  NAND2_X1 U8829 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7156) );
  OAI21_X1 U8830 ( .B1(n7054), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7102), .ZN(
        n7055) );
  AOI22_X1 U8831 ( .A1(n7807), .A2(P2_ADDR_REG_5__SCAN_IN), .B1(n7183), .B2(
        n7055), .ZN(n7056) );
  OAI211_X1 U8832 ( .C1(n7057), .C2(n10020), .A(n7156), .B(n7056), .ZN(n7062)
         );
  AOI211_X1 U8833 ( .C1(n7060), .C2(n7059), .A(n7252), .B(n7058), .ZN(n7061)
         );
  AOI211_X1 U8834 ( .C1(n8528), .C2(n7063), .A(n7062), .B(n7061), .ZN(n7064)
         );
  INV_X1 U8835 ( .A(n7064), .ZN(P2_U3187) );
  XNOR2_X1 U8836 ( .A(n7367), .B(n8234), .ZN(n7154) );
  XNOR2_X1 U8837 ( .A(n7154), .B(n7160), .ZN(n7068) );
  AOI21_X1 U8838 ( .B1(n7068), .B2(n7067), .A(n7155), .ZN(n7075) );
  NAND2_X1 U8839 ( .A1(n8200), .A2(n8459), .ZN(n7072) );
  INV_X1 U8840 ( .A(n7069), .ZN(n7070) );
  AOI21_X1 U8841 ( .B1(n8176), .B2(n8245), .A(n7070), .ZN(n7071) );
  OAI211_X1 U8842 ( .C1(n7146), .C2(n8202), .A(n7072), .B(n7071), .ZN(n7073)
         );
  AOI21_X1 U8843 ( .B1(n7195), .B2(n8204), .A(n7073), .ZN(n7074) );
  OAI21_X1 U8844 ( .B1(n7075), .B2(n8195), .A(n7074), .ZN(P2_U3170) );
  INV_X1 U8845 ( .A(n7637), .ZN(n7554) );
  NAND3_X1 U8846 ( .A1(n7143), .A2(n8227), .A3(n8379), .ZN(n7076) );
  NAND2_X1 U8847 ( .A1(n7132), .A2(n7076), .ZN(n7228) );
  NAND2_X1 U8848 ( .A1(n8460), .A2(n4275), .ZN(n8244) );
  XNOR2_X1 U8849 ( .A(n7077), .B(n7078), .ZN(n7079) );
  OAI222_X1 U8850 ( .A1(n8693), .A2(n4987), .B1(n8244), .B2(n7080), .C1(n10037), .C2(n7079), .ZN(n7223) );
  AOI21_X1 U8851 ( .B1(n10049), .B2(n7228), .A(n7223), .ZN(n7086) );
  INV_X1 U8852 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7081) );
  OAI22_X1 U8853 ( .A1(n7082), .A2(n8791), .B1(n10085), .B2(n7081), .ZN(n7083)
         );
  INV_X1 U8854 ( .A(n7083), .ZN(n7084) );
  OAI21_X1 U8855 ( .B1(n7086), .B2(n10087), .A(n7084), .ZN(P2_U3399) );
  AOI22_X1 U8856 ( .A1(n8744), .A2(n7225), .B1(n10100), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n7085) );
  OAI21_X1 U8857 ( .B1(n7086), .B2(n10100), .A(n7085), .ZN(P2_U3462) );
  INV_X1 U8858 ( .A(n7087), .ZN(n10011) );
  INV_X1 U8859 ( .A(n7088), .ZN(n7089) );
  INV_X1 U8860 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9310) );
  OAI222_X1 U8861 ( .A1(n10011), .A2(P2_U3151), .B1(n8822), .B2(n7089), .C1(
        n9310), .C2(n8824), .ZN(P2_U3278) );
  INV_X1 U8862 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7090) );
  INV_X1 U8863 ( .A(n9079), .ZN(n9067) );
  OAI222_X1 U8864 ( .A1(n8064), .A2(n7090), .B1(n9590), .B2(n7089), .C1(
        P1_U3086), .C2(n9067), .ZN(P1_U3338) );
  INV_X1 U8865 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7092) );
  OAI222_X1 U8866 ( .A1(n8824), .A2(n7092), .B1(n8822), .B2(n7093), .C1(
        P2_U3151), .C2(n7091), .ZN(P2_U3277) );
  INV_X1 U8867 ( .A(n9800), .ZN(n7094) );
  INV_X1 U8868 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9385) );
  OAI222_X1 U8869 ( .A1(P1_U3086), .A2(n7094), .B1(n9590), .B2(n7093), .C1(
        n9385), .C2(n8064), .ZN(P1_U3337) );
  OAI21_X1 U8870 ( .B1(n7097), .B2(n7096), .A(n7095), .ZN(n7098) );
  NAND2_X1 U8871 ( .A1(n7098), .A2(n10031), .ZN(n7114) );
  INV_X1 U8872 ( .A(n7099), .ZN(n7101) );
  NAND3_X1 U8873 ( .A1(n7102), .A2(n7101), .A3(n7100), .ZN(n7103) );
  AOI21_X1 U8874 ( .B1(n7104), .B2(n7103), .A(n10026), .ZN(n7112) );
  AND3_X1 U8875 ( .A1(n7107), .A2(n7106), .A3(n7105), .ZN(n7108) );
  OAI21_X1 U8876 ( .B1(n7109), .B2(n7108), .A(n7180), .ZN(n7110) );
  NAND2_X1 U8877 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7382) );
  NAND2_X1 U8878 ( .A1(n7110), .A2(n7382), .ZN(n7111) );
  AOI211_X1 U8879 ( .C1(n7807), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n7112), .B(
        n7111), .ZN(n7113) );
  OAI211_X1 U8880 ( .C1(n10012), .C2(n7115), .A(n7114), .B(n7113), .ZN(
        P2_U3188) );
  XOR2_X1 U8881 ( .A(n7117), .B(n7116), .Z(n7123) );
  NAND2_X1 U8882 ( .A1(n7119), .A2(n7118), .ZN(n8060) );
  INV_X1 U8883 ( .A(n8202), .ZN(n8189) );
  AOI22_X1 U8884 ( .A1(n8189), .A2(n8464), .B1(n7931), .B2(n8176), .ZN(n7120)
         );
  OAI21_X1 U8885 ( .B1(n4987), .B2(n8191), .A(n7120), .ZN(n7121) );
  AOI21_X1 U8886 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n8060), .A(n7121), .ZN(
        n7122) );
  OAI21_X1 U8887 ( .B1(n8195), .B2(n7123), .A(n7122), .ZN(P2_U3162) );
  XOR2_X1 U8888 ( .A(n7124), .B(n7125), .Z(n7130) );
  AOI22_X1 U8889 ( .A1(n8189), .A2(n6985), .B1(n7126), .B2(n8176), .ZN(n7127)
         );
  OAI21_X1 U8890 ( .B1(n7146), .B2(n8191), .A(n7127), .ZN(n7128) );
  AOI21_X1 U8891 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n8060), .A(n7128), .ZN(
        n7129) );
  OAI21_X1 U8892 ( .B1(n8195), .B2(n7130), .A(n7129), .ZN(P2_U3177) );
  NAND2_X1 U8893 ( .A1(n7132), .A2(n8243), .ZN(n7131) );
  NAND2_X1 U8894 ( .A1(n7131), .A2(n7136), .ZN(n7134) );
  INV_X1 U8895 ( .A(n7136), .ZN(n8386) );
  NAND3_X1 U8896 ( .A1(n7132), .A2(n8386), .A3(n8243), .ZN(n7133) );
  NAND2_X1 U8897 ( .A1(n7134), .A2(n7133), .ZN(n7188) );
  XNOR2_X1 U8898 ( .A(n7135), .B(n7136), .ZN(n7137) );
  OAI222_X1 U8899 ( .A1(n8695), .A2(n4880), .B1(n8693), .B2(n7146), .C1(n7137), 
        .C2(n10037), .ZN(n7192) );
  AOI21_X1 U8900 ( .B1(n10049), .B2(n7188), .A(n7192), .ZN(n7142) );
  AOI22_X1 U8901 ( .A1(n8744), .A2(n8245), .B1(n10100), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n7138) );
  OAI21_X1 U8902 ( .B1(n7142), .B2(n10100), .A(n7138), .ZN(P2_U3463) );
  INV_X1 U8903 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7139) );
  OAI22_X1 U8904 ( .A1(n8234), .A2(n8791), .B1(n10085), .B2(n7139), .ZN(n7140)
         );
  INV_X1 U8905 ( .A(n7140), .ZN(n7141) );
  OAI21_X1 U8906 ( .B1(n7142), .B2(n10087), .A(n7141), .ZN(P2_U3402) );
  OAI21_X1 U8907 ( .B1(n7144), .B2(n8224), .A(n7143), .ZN(n7148) );
  INV_X1 U8908 ( .A(n7148), .ZN(n10041) );
  NOR2_X1 U8909 ( .A1(n6973), .A2(n6975), .ZN(n7189) );
  NAND2_X1 U8910 ( .A1(n8699), .A2(n7189), .ZN(n8551) );
  NOR2_X1 U8911 ( .A1(n6979), .A2(n8588), .ZN(n7151) );
  XNOR2_X1 U8912 ( .A(n7145), .B(n8224), .ZN(n7150) );
  OAI22_X1 U8913 ( .A1(n6984), .A2(n8693), .B1(n7146), .B2(n8695), .ZN(n7147)
         );
  AOI21_X1 U8914 ( .B1(n7148), .B2(n7637), .A(n7147), .ZN(n7149) );
  OAI21_X1 U8915 ( .B1(n10037), .B2(n7150), .A(n7149), .ZN(n10043) );
  AOI211_X1 U8916 ( .C1(n8685), .C2(P2_REG3_REG_2__SCAN_IN), .A(n7151), .B(
        n10043), .ZN(n7152) );
  MUX2_X1 U8917 ( .A(n9331), .B(n7152), .S(n8682), .Z(n7153) );
  OAI21_X1 U8918 ( .B1(n10041), .B2(n8551), .A(n7153), .ZN(P2_U3231) );
  XOR2_X1 U8919 ( .A(n7366), .B(n4407), .Z(n7163) );
  NAND2_X1 U8920 ( .A1(n8200), .A2(n8458), .ZN(n7159) );
  INV_X1 U8921 ( .A(n7156), .ZN(n7157) );
  AOI21_X1 U8922 ( .B1(n8176), .B2(n7220), .A(n7157), .ZN(n7158) );
  OAI211_X1 U8923 ( .C1(n7160), .C2(n8202), .A(n7159), .B(n7158), .ZN(n7161)
         );
  AOI21_X1 U8924 ( .B1(n7207), .B2(n8204), .A(n7161), .ZN(n7162) );
  OAI21_X1 U8925 ( .B1(n7163), .B2(n8195), .A(n7162), .ZN(P2_U3167) );
  NAND2_X1 U8926 ( .A1(n7164), .A2(n7165), .ZN(n7166) );
  XOR2_X1 U8927 ( .A(n7167), .B(n7166), .Z(n7172) );
  NOR2_X1 U8928 ( .A1(n8944), .A2(n7302), .ZN(n7170) );
  AOI22_X1 U8929 ( .A1(n8928), .A2(n8970), .B1(n8968), .B2(n8929), .ZN(n7295)
         );
  OAI22_X1 U8930 ( .A1(n7295), .A2(n8918), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7168), .ZN(n7169) );
  AOI211_X1 U8931 ( .C1(n9932), .C2(n8934), .A(n7170), .B(n7169), .ZN(n7171)
         );
  OAI21_X1 U8932 ( .B1(n7172), .B2(n8923), .A(n7171), .ZN(P1_U3227) );
  XOR2_X1 U8933 ( .A(n7174), .B(n7173), .Z(n7187) );
  OAI21_X1 U8934 ( .B1(n7176), .B2(P2_REG1_REG_7__SCAN_IN), .A(n7175), .ZN(
        n7181) );
  NAND2_X1 U8935 ( .A1(n7807), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7177) );
  NAND2_X1 U8936 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7373) );
  OAI211_X1 U8937 ( .C1(n10012), .C2(n7178), .A(n7177), .B(n7373), .ZN(n7179)
         );
  AOI21_X1 U8938 ( .B1(n7181), .B2(n7180), .A(n7179), .ZN(n7186) );
  OAI21_X1 U8939 ( .B1(n4338), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7182), .ZN(
        n7184) );
  NAND2_X1 U8940 ( .A1(n7184), .A2(n7183), .ZN(n7185) );
  OAI211_X1 U8941 ( .C1(n7187), .C2(n7252), .A(n7186), .B(n7185), .ZN(P2_U3189) );
  INV_X1 U8942 ( .A(n7188), .ZN(n7198) );
  INV_X1 U8943 ( .A(n7189), .ZN(n7190) );
  NAND2_X1 U8944 ( .A1(n7554), .A2(n7190), .ZN(n7191) );
  INV_X1 U8945 ( .A(n7192), .ZN(n7193) );
  MUX2_X1 U8946 ( .A(n7194), .B(n7193), .S(n8682), .Z(n7197) );
  AOI22_X1 U8947 ( .A1(n8702), .A2(n8245), .B1(n8685), .B2(n7195), .ZN(n7196)
         );
  OAI211_X1 U8948 ( .C1(n7198), .C2(n8705), .A(n7197), .B(n7196), .ZN(P2_U3229) );
  INV_X1 U8949 ( .A(n7199), .ZN(n7200) );
  NOR2_X1 U8950 ( .A1(n7201), .A2(n7200), .ZN(n7206) );
  XOR2_X1 U8951 ( .A(n7206), .B(n7202), .Z(n7203) );
  OAI222_X1 U8952 ( .A1(n8244), .A2(n7204), .B1(n7203), .B2(n10037), .C1(n8695), .C2(n7378), .ZN(n7214) );
  INV_X1 U8953 ( .A(n7214), .ZN(n7213) );
  XOR2_X1 U8954 ( .A(n7206), .B(n7205), .Z(n7215) );
  INV_X1 U8955 ( .A(n8705), .ZN(n7211) );
  INV_X1 U8956 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7209) );
  AOI22_X1 U8957 ( .A1(n8702), .A2(n7220), .B1(n8685), .B2(n7207), .ZN(n7208)
         );
  OAI21_X1 U8958 ( .B1(n7209), .B2(n8682), .A(n7208), .ZN(n7210) );
  AOI21_X1 U8959 ( .B1(n7215), .B2(n7211), .A(n7210), .ZN(n7212) );
  OAI21_X1 U8960 ( .B1(n7213), .B2(n8701), .A(n7212), .ZN(P2_U3228) );
  AOI21_X1 U8961 ( .B1(n10049), .B2(n7215), .A(n7214), .ZN(n7222) );
  INV_X1 U8962 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7216) );
  OAI22_X1 U8963 ( .A1(n7217), .A2(n8791), .B1(n10085), .B2(n7216), .ZN(n7218)
         );
  INV_X1 U8964 ( .A(n7218), .ZN(n7219) );
  OAI21_X1 U8965 ( .B1(n7222), .B2(n10087), .A(n7219), .ZN(P2_U3405) );
  AOI22_X1 U8966 ( .A1(n8744), .A2(n7220), .B1(n10100), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n7221) );
  OAI21_X1 U8967 ( .B1(n7222), .B2(n10100), .A(n7221), .ZN(P2_U3464) );
  INV_X1 U8968 ( .A(n7223), .ZN(n7230) );
  AOI22_X1 U8969 ( .A1(n8702), .A2(n7225), .B1(n8685), .B2(n7224), .ZN(n7226)
         );
  OAI21_X1 U8970 ( .B1(n4741), .B2(n8682), .A(n7226), .ZN(n7227) );
  AOI21_X1 U8971 ( .B1(n7211), .B2(n7228), .A(n7227), .ZN(n7229) );
  OAI21_X1 U8972 ( .B1(n7230), .B2(n8701), .A(n7229), .ZN(P2_U3230) );
  INV_X1 U8973 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7233) );
  INV_X1 U8974 ( .A(n7231), .ZN(n7235) );
  OAI222_X1 U8975 ( .A1(n8064), .A2(n7233), .B1(n9590), .B2(n7235), .C1(
        P1_U3086), .C2(n7232), .ZN(P1_U3336) );
  INV_X1 U8976 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7234) );
  OAI222_X1 U8977 ( .A1(n5559), .A2(P2_U3151), .B1(n8822), .B2(n7235), .C1(
        n7234), .C2(n8824), .ZN(P2_U3276) );
  NAND2_X1 U8978 ( .A1(n8463), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7236) );
  OAI21_X1 U8979 ( .B1(n8046), .B2(n8463), .A(n7236), .ZN(P2_U3520) );
  XOR2_X1 U8980 ( .A(n7238), .B(n7237), .Z(n7253) );
  INV_X1 U8981 ( .A(n7239), .ZN(n7242) );
  NAND3_X1 U8982 ( .A1(n7175), .A2(n7240), .A3(n4318), .ZN(n7241) );
  AOI21_X1 U8983 ( .B1(n7242), .B2(n7241), .A(n10020), .ZN(n7250) );
  NAND3_X1 U8984 ( .A1(n7182), .A2(n4415), .A3(n7243), .ZN(n7244) );
  AOI21_X1 U8985 ( .B1(n7245), .B2(n7244), .A(n10026), .ZN(n7249) );
  NAND2_X1 U8986 ( .A1(n7807), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7246) );
  NAND2_X1 U8987 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7537) );
  OAI211_X1 U8988 ( .C1(n10012), .C2(n7247), .A(n7246), .B(n7537), .ZN(n7248)
         );
  NOR3_X1 U8989 ( .A1(n7250), .A2(n7249), .A3(n7248), .ZN(n7251) );
  OAI21_X1 U8990 ( .B1(n7253), .B2(n7252), .A(n7251), .ZN(P2_U3190) );
  AOI21_X1 U8991 ( .B1(n7256), .B2(n7254), .A(n7255), .ZN(n7262) );
  NAND2_X1 U8992 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9725) );
  INV_X1 U8993 ( .A(n9725), .ZN(n7258) );
  AOI22_X1 U8994 ( .A1(n8928), .A2(n8969), .B1(n8967), .B2(n8929), .ZN(n9844)
         );
  NOR2_X1 U8995 ( .A1(n9844), .A2(n8918), .ZN(n7257) );
  AOI211_X1 U8996 ( .C1(n7324), .C2(n8934), .A(n7258), .B(n7257), .ZN(n7261)
         );
  INV_X1 U8997 ( .A(n7259), .ZN(n9848) );
  NAND2_X1 U8998 ( .A1(n8921), .A2(n9848), .ZN(n7260) );
  OAI211_X1 U8999 ( .C1(n7262), .C2(n8923), .A(n7261), .B(n7260), .ZN(P1_U3239) );
  INV_X1 U9000 ( .A(n7263), .ZN(n7267) );
  OAI21_X1 U9001 ( .B1(n7267), .B2(n7266), .A(n9901), .ZN(n7269) );
  NAND4_X1 U9002 ( .A1(n7269), .A2(n7307), .A3(n9583), .A4(n7268), .ZN(n7270)
         );
  AND2_X1 U9003 ( .A1(n7521), .A2(n7494), .ZN(n9670) );
  AND2_X1 U9004 ( .A1(n8975), .A2(n7330), .ZN(n7515) );
  NAND2_X1 U9005 ( .A1(n9885), .A2(n9886), .ZN(n7273) );
  NAND2_X1 U9006 ( .A1(n7276), .A2(n9913), .ZN(n7272) );
  NAND2_X1 U9007 ( .A1(n7273), .A2(n7272), .ZN(n7286) );
  XNOR2_X1 U9008 ( .A(n7286), .B(n7284), .ZN(n9922) );
  OAI21_X1 U9009 ( .B1(n7275), .B2(n7284), .A(n7274), .ZN(n7277) );
  OAI22_X1 U9010 ( .A1(n7291), .A2(n7569), .B1(n7276), .B2(n9167), .ZN(n8843)
         );
  AOI21_X1 U9011 ( .B1(n7277), .B2(n9876), .A(n8843), .ZN(n9920) );
  INV_X2 U9012 ( .A(n9881), .ZN(n9671) );
  MUX2_X1 U9013 ( .A(n9431), .B(n9920), .S(n9671), .Z(n7283) );
  NAND2_X1 U9014 ( .A1(n9907), .A2(n7523), .ZN(n9887) );
  INV_X1 U9015 ( .A(n7279), .ZN(n9889) );
  INV_X1 U9016 ( .A(n7300), .ZN(n9870) );
  AOI211_X1 U9017 ( .C1(n4271), .C2(n9889), .A(n9481), .B(n9870), .ZN(n9918)
         );
  INV_X1 U9018 ( .A(n9667), .ZN(n7280) );
  OAI22_X1 U9019 ( .A1(n9883), .A2(n7287), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9879), .ZN(n7281) );
  AOI21_X1 U9020 ( .B1(n9918), .B2(n9892), .A(n7281), .ZN(n7282) );
  OAI211_X1 U9021 ( .C1(n9488), .C2(n9922), .A(n7283), .B(n7282), .ZN(P1_U3290) );
  INV_X1 U9022 ( .A(n7284), .ZN(n7285) );
  NAND2_X1 U9023 ( .A1(n7286), .A2(n7285), .ZN(n7290) );
  NAND2_X1 U9024 ( .A1(n7288), .A2(n7287), .ZN(n7289) );
  NAND2_X1 U9025 ( .A1(n7290), .A2(n7289), .ZN(n9867) );
  INV_X1 U9026 ( .A(n9860), .ZN(n9868) );
  NAND2_X1 U9027 ( .A1(n7291), .A2(n9925), .ZN(n7292) );
  XNOR2_X1 U9028 ( .A(n7310), .B(n7293), .ZN(n9936) );
  XNOR2_X1 U9029 ( .A(n7294), .B(n7293), .ZN(n7297) );
  INV_X1 U9030 ( .A(n7295), .ZN(n7296) );
  AOI21_X1 U9031 ( .B1(n7297), .B2(n9876), .A(n7296), .ZN(n9935) );
  MUX2_X1 U9032 ( .A(n7298), .B(n9935), .S(n9671), .Z(n7305) );
  AOI21_X1 U9033 ( .B1(n9869), .B2(n9932), .A(n9481), .ZN(n7301) );
  AND2_X1 U9034 ( .A1(n7301), .A2(n9853), .ZN(n9931) );
  OAI22_X1 U9035 ( .A1(n9883), .A2(n7311), .B1(n9879), .B2(n7302), .ZN(n7303)
         );
  AOI21_X1 U9036 ( .B1(n9931), .B2(n9892), .A(n7303), .ZN(n7304) );
  OAI211_X1 U9037 ( .C1(n9936), .C2(n9488), .A(n7305), .B(n7304), .ZN(P1_U3288) );
  INV_X1 U9038 ( .A(n7306), .ZN(n7308) );
  NAND2_X1 U9039 ( .A1(n7313), .A2(n7318), .ZN(n9852) );
  NAND2_X1 U9040 ( .A1(n9851), .A2(n9852), .ZN(n7316) );
  NAND2_X1 U9041 ( .A1(n9940), .A2(n7314), .ZN(n7315) );
  NAND2_X1 U9042 ( .A1(n7316), .A2(n7315), .ZN(n7475) );
  XNOR2_X1 U9043 ( .A(n7475), .B(n7473), .ZN(n7359) );
  AOI21_X1 U9044 ( .B1(n9843), .B2(n7318), .A(n7317), .ZN(n7319) );
  NAND2_X1 U9045 ( .A1(n7319), .A2(n7473), .ZN(n7560) );
  OAI21_X1 U9046 ( .B1(n7319), .B2(n7473), .A(n7560), .ZN(n7323) );
  NAND2_X1 U9047 ( .A1(n8968), .A2(n8928), .ZN(n7321) );
  NAND2_X1 U9048 ( .A1(n8966), .A2(n8929), .ZN(n7320) );
  AND2_X1 U9049 ( .A1(n7321), .A2(n7320), .ZN(n7451) );
  INV_X1 U9050 ( .A(n7451), .ZN(n7322) );
  AOI21_X1 U9051 ( .B1(n7323), .B2(n9876), .A(n7322), .ZN(n7362) );
  INV_X1 U9052 ( .A(n7325), .ZN(n9854) );
  AOI211_X1 U9053 ( .C1(n7455), .C2(n9854), .A(n9481), .B(n9838), .ZN(n7358)
         );
  AOI21_X1 U9054 ( .B1(n9933), .B2(n7455), .A(n7358), .ZN(n7326) );
  OAI211_X1 U9055 ( .C1(n9937), .C2(n7359), .A(n7362), .B(n7326), .ZN(n7328)
         );
  NAND2_X1 U9056 ( .A1(n7328), .A2(n9991), .ZN(n7327) );
  OAI21_X1 U9057 ( .B1(n9991), .B2(n5833), .A(n7327), .ZN(P1_U3474) );
  NAND2_X1 U9058 ( .A1(n7328), .A2(n9569), .ZN(n7329) );
  OAI21_X1 U9059 ( .B1(n9569), .B2(n6802), .A(n7329), .ZN(P1_U3529) );
  NOR2_X1 U9060 ( .A1(n9499), .A2(n9481), .ZN(n9266) );
  OAI21_X1 U9061 ( .B1(n9266), .B2(n9835), .A(n7330), .ZN(n7339) );
  INV_X1 U9062 ( .A(n7331), .ZN(n7334) );
  NAND3_X1 U9063 ( .A1(n7334), .A2(n7333), .A3(n7332), .ZN(n7336) );
  OAI211_X1 U9064 ( .C1(n5700), .C2(n9879), .A(n7336), .B(n7335), .ZN(n7337)
         );
  NAND2_X1 U9065 ( .A1(n7337), .A2(n9671), .ZN(n7338) );
  OAI211_X1 U9066 ( .C1(n9671), .C2(n7340), .A(n7339), .B(n7338), .ZN(P1_U3293) );
  AOI21_X1 U9067 ( .B1(n9303), .B2(n7342), .A(n7341), .ZN(n7355) );
  INV_X1 U9068 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7409) );
  AND2_X1 U9069 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7600) );
  INV_X1 U9070 ( .A(n7600), .ZN(n7343) );
  OAI21_X1 U9071 ( .B1(n10010), .B2(n7409), .A(n7343), .ZN(n7347) );
  AOI21_X1 U9072 ( .B1(n7344), .B2(n10094), .A(n4409), .ZN(n7345) );
  NOR2_X1 U9073 ( .A1(n7345), .A2(n10020), .ZN(n7346) );
  AOI211_X1 U9074 ( .C1(n8528), .C2(n7348), .A(n7347), .B(n7346), .ZN(n7354)
         );
  OAI21_X1 U9075 ( .B1(n7351), .B2(n7350), .A(n7349), .ZN(n7352) );
  NAND2_X1 U9076 ( .A1(n7352), .A2(n10031), .ZN(n7353) );
  OAI211_X1 U9077 ( .C1(n7355), .C2(n10026), .A(n7354), .B(n7353), .ZN(
        P2_U3191) );
  NOR2_X1 U9078 ( .A1(n7477), .A2(n9883), .ZN(n7357) );
  OAI22_X1 U9079 ( .A1(n9671), .A2(n5830), .B1(n7452), .B2(n9879), .ZN(n7356)
         );
  AOI211_X1 U9080 ( .C1(n7358), .C2(n9892), .A(n7357), .B(n7356), .ZN(n7361)
         );
  OR2_X1 U9081 ( .A1(n7359), .A2(n9488), .ZN(n7360) );
  OAI211_X1 U9082 ( .C1(n7362), .C2(n9896), .A(n7361), .B(n7360), .ZN(P1_U3286) );
  XNOR2_X1 U9083 ( .A(n8037), .B(n7375), .ZN(n7534) );
  XNOR2_X1 U9084 ( .A(n7534), .B(n7364), .ZN(n7371) );
  XNOR2_X1 U9085 ( .A(n7367), .B(n10046), .ZN(n7368) );
  XNOR2_X1 U9086 ( .A(n7368), .B(n7378), .ZN(n7388) );
  INV_X1 U9087 ( .A(n7368), .ZN(n7369) );
  NAND2_X1 U9088 ( .A1(n7370), .A2(n7371), .ZN(n7536) );
  OAI21_X1 U9089 ( .B1(n7371), .B2(n7370), .A(n7536), .ZN(n7372) );
  NAND2_X1 U9090 ( .A1(n7372), .A2(n8185), .ZN(n7381) );
  NAND2_X1 U9091 ( .A1(n8200), .A2(n5090), .ZN(n7377) );
  INV_X1 U9092 ( .A(n7373), .ZN(n7374) );
  AOI21_X1 U9093 ( .B1(n8176), .B2(n7375), .A(n7374), .ZN(n7376) );
  OAI211_X1 U9094 ( .C1(n7378), .C2(n8202), .A(n7377), .B(n7376), .ZN(n7379)
         );
  AOI21_X1 U9095 ( .B1(n7465), .B2(n8204), .A(n7379), .ZN(n7380) );
  NAND2_X1 U9096 ( .A1(n7381), .A2(n7380), .ZN(P2_U3153) );
  NAND2_X1 U9097 ( .A1(n8200), .A2(n8457), .ZN(n7385) );
  INV_X1 U9098 ( .A(n7382), .ZN(n7383) );
  AOI21_X1 U9099 ( .B1(n8176), .B2(n7443), .A(n7383), .ZN(n7384) );
  OAI211_X1 U9100 ( .C1(n4880), .C2(n8202), .A(n7385), .B(n7384), .ZN(n7390)
         );
  AOI211_X1 U9101 ( .C1(n7388), .C2(n7386), .A(n8195), .B(n7387), .ZN(n7389)
         );
  AOI211_X1 U9102 ( .C1(n7442), .C2(n8204), .A(n7390), .B(n7389), .ZN(n7391)
         );
  INV_X1 U9103 ( .A(n7391), .ZN(P2_U3179) );
  NOR2_X1 U9104 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7430) );
  NOR2_X1 U9105 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7428) );
  NOR2_X1 U9106 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n7426) );
  NOR2_X1 U9107 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7424) );
  NOR2_X1 U9108 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7422) );
  NOR2_X1 U9109 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(P2_ADDR_REG_12__SCAN_IN), 
        .ZN(n7420) );
  NOR2_X1 U9110 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7417) );
  NOR2_X1 U9111 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7414) );
  NOR2_X1 U9112 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7412) );
  NOR2_X1 U9113 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7408) );
  NOR2_X1 U9114 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7406) );
  NOR2_X1 U9115 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7404) );
  NOR2_X1 U9116 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7402) );
  NOR2_X1 U9117 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7400) );
  NAND2_X1 U9118 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7398) );
  INV_X1 U9119 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9008) );
  XNOR2_X1 U9120 ( .A(n9008), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n10139) );
  NAND2_X1 U9121 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7396) );
  AOI21_X1 U9122 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10105) );
  INV_X1 U9123 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7393) );
  NAND2_X1 U9124 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7392) );
  NOR2_X1 U9125 ( .A1(n7393), .A2(n7392), .ZN(n10104) );
  NOR2_X1 U9126 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10104), .ZN(n7394) );
  NOR2_X1 U9127 ( .A1(n10105), .A2(n7394), .ZN(n10137) );
  XOR2_X1 U9128 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10136) );
  NAND2_X1 U9129 ( .A1(n10137), .A2(n10136), .ZN(n7395) );
  NAND2_X1 U9130 ( .A1(n7396), .A2(n7395), .ZN(n10138) );
  NAND2_X1 U9131 ( .A1(n10139), .A2(n10138), .ZN(n7397) );
  NAND2_X1 U9132 ( .A1(n7398), .A2(n7397), .ZN(n10141) );
  XNOR2_X1 U9133 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10140) );
  NOR2_X1 U9134 ( .A1(n10141), .A2(n10140), .ZN(n7399) );
  NOR2_X1 U9135 ( .A1(n7400), .A2(n7399), .ZN(n10129) );
  INV_X1 U9136 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9710) );
  XOR2_X1 U9137 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n9710), .Z(n10128) );
  NOR2_X1 U9138 ( .A1(n10129), .A2(n10128), .ZN(n7401) );
  NOR2_X1 U9139 ( .A1(n7402), .A2(n7401), .ZN(n10127) );
  INV_X1 U9140 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9727) );
  XOR2_X1 U9141 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n9727), .Z(n10126) );
  NOR2_X1 U9142 ( .A1(n10127), .A2(n10126), .ZN(n7403) );
  NOR2_X1 U9143 ( .A1(n7404), .A2(n7403), .ZN(n10133) );
  INV_X1 U9144 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9622) );
  XOR2_X1 U9145 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n9622), .Z(n10132) );
  NOR2_X1 U9146 ( .A1(n10133), .A2(n10132), .ZN(n7405) );
  NOR2_X1 U9147 ( .A1(n7406), .A2(n7405), .ZN(n10135) );
  INV_X1 U9148 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9639) );
  XOR2_X1 U9149 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n9639), .Z(n10134) );
  NOR2_X1 U9150 ( .A1(n10135), .A2(n10134), .ZN(n7407) );
  NOR2_X1 U9151 ( .A1(n7408), .A2(n7407), .ZN(n10131) );
  INV_X1 U9152 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7410) );
  AOI22_X1 U9153 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7410), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n7409), .ZN(n10130) );
  NOR2_X1 U9154 ( .A1(n10131), .A2(n10130), .ZN(n7411) );
  NOR2_X1 U9155 ( .A1(n7412), .A2(n7411), .ZN(n10125) );
  INV_X1 U9156 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9605) );
  INV_X1 U9157 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7712) );
  AOI22_X1 U9158 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n9605), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n7712), .ZN(n10124) );
  NOR2_X1 U9159 ( .A1(n10125), .A2(n10124), .ZN(n7413) );
  NOR2_X1 U9160 ( .A1(n7414), .A2(n7413), .ZN(n10123) );
  INV_X1 U9161 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9745) );
  INV_X1 U9162 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7415) );
  AOI22_X1 U9163 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n9745), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n7415), .ZN(n10122) );
  NOR2_X1 U9164 ( .A1(n10123), .A2(n10122), .ZN(n7416) );
  NOR2_X1 U9165 ( .A1(n7417), .A2(n7416), .ZN(n10121) );
  INV_X1 U9166 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7885) );
  INV_X1 U9167 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7418) );
  AOI22_X1 U9168 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(n7885), .B1(
        P2_ADDR_REG_12__SCAN_IN), .B2(n7418), .ZN(n10120) );
  NOR2_X1 U9169 ( .A1(n10121), .A2(n10120), .ZN(n7419) );
  NOR2_X1 U9170 ( .A1(n7420), .A2(n7419), .ZN(n10119) );
  INV_X1 U9171 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9757) );
  XOR2_X1 U9172 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n9757), .Z(n10118) );
  NOR2_X1 U9173 ( .A1(n10119), .A2(n10118), .ZN(n7421) );
  NOR2_X1 U9174 ( .A1(n7422), .A2(n7421), .ZN(n10117) );
  INV_X1 U9175 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9777) );
  XOR2_X1 U9176 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n9777), .Z(n10116) );
  NOR2_X1 U9177 ( .A1(n10117), .A2(n10116), .ZN(n7423) );
  NOR2_X1 U9178 ( .A1(n7424), .A2(n7423), .ZN(n10115) );
  INV_X1 U9179 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8491) );
  INV_X1 U9180 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9787) );
  AOI22_X1 U9181 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n8491), .B1(
        P2_ADDR_REG_15__SCAN_IN), .B2(n9787), .ZN(n10114) );
  NOR2_X1 U9182 ( .A1(n10115), .A2(n10114), .ZN(n7425) );
  NOR2_X1 U9183 ( .A1(n7426), .A2(n7425), .ZN(n10113) );
  XNOR2_X1 U9184 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10112) );
  NOR2_X1 U9185 ( .A1(n10113), .A2(n10112), .ZN(n7427) );
  NOR2_X1 U9186 ( .A1(n7428), .A2(n7427), .ZN(n10111) );
  XNOR2_X1 U9187 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10110) );
  NOR2_X1 U9188 ( .A1(n10111), .A2(n10110), .ZN(n7429) );
  NOR2_X1 U9189 ( .A1(n7430), .A2(n7429), .ZN(n7431) );
  AND2_X1 U9190 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7431), .ZN(n10107) );
  NOR2_X1 U9191 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10107), .ZN(n7432) );
  NOR2_X1 U9192 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n7431), .ZN(n10108) );
  NOR2_X1 U9193 ( .A1(n7432), .A2(n10108), .ZN(n7434) );
  XNOR2_X1 U9194 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7433) );
  XNOR2_X1 U9195 ( .A(n7434), .B(n7433), .ZN(ADD_1068_U4) );
  INV_X1 U9196 ( .A(n7435), .ZN(n7470) );
  OAI222_X1 U9197 ( .A1(P2_U3151), .A2(n8412), .B1(n8822), .B2(n7470), .C1(
        n7436), .C2(n8824), .ZN(P2_U3275) );
  NAND2_X1 U9198 ( .A1(n8382), .A2(n8248), .ZN(n7439) );
  OAI21_X1 U9199 ( .B1(n7205), .B2(n8384), .A(n8247), .ZN(n7437) );
  XOR2_X1 U9200 ( .A(n7439), .B(n7437), .Z(n10044) );
  XOR2_X1 U9201 ( .A(n7439), .B(n7438), .Z(n7440) );
  AOI222_X1 U9202 ( .A1(n8657), .A2(n7440), .B1(n8457), .B2(n8653), .C1(n8459), 
        .C2(n8655), .ZN(n10045) );
  MUX2_X1 U9203 ( .A(n7441), .B(n10045), .S(n8682), .Z(n7445) );
  AOI22_X1 U9204 ( .A1(n8702), .A2(n7443), .B1(n8685), .B2(n7442), .ZN(n7444)
         );
  OAI211_X1 U9205 ( .C1(n10044), .C2(n8705), .A(n7445), .B(n7444), .ZN(
        P2_U3227) );
  NAND2_X1 U9206 ( .A1(n7448), .A2(n7447), .ZN(n7449) );
  XOR2_X1 U9207 ( .A(n7446), .B(n7449), .Z(n7457) );
  OAI22_X1 U9208 ( .A1(n7451), .A2(n8918), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7450), .ZN(n7454) );
  NOR2_X1 U9209 ( .A1(n8944), .A2(n7452), .ZN(n7453) );
  AOI211_X1 U9210 ( .C1(n7455), .C2(n8934), .A(n7454), .B(n7453), .ZN(n7456)
         );
  OAI21_X1 U9211 ( .B1(n7457), .B2(n8923), .A(n7456), .ZN(P1_U3213) );
  OR2_X1 U9212 ( .A1(n7458), .A2(n8256), .ZN(n7623) );
  NAND2_X1 U9213 ( .A1(n7458), .A2(n8256), .ZN(n7459) );
  NAND2_X1 U9214 ( .A1(n7623), .A2(n7459), .ZN(n10052) );
  NAND2_X1 U9215 ( .A1(n7461), .A2(n7460), .ZN(n7625) );
  INV_X1 U9216 ( .A(n8256), .ZN(n8388) );
  XNOR2_X1 U9217 ( .A(n7625), .B(n8388), .ZN(n7462) );
  NAND2_X1 U9218 ( .A1(n7462), .A2(n8657), .ZN(n7464) );
  AOI22_X1 U9219 ( .A1(n8655), .A2(n8458), .B1(n5090), .B2(n8653), .ZN(n7463)
         );
  OAI211_X1 U9220 ( .C1(n7554), .C2(n10052), .A(n7464), .B(n7463), .ZN(n10054)
         );
  NAND2_X1 U9221 ( .A1(n10054), .A2(n8699), .ZN(n7469) );
  INV_X1 U9222 ( .A(n7465), .ZN(n7466) );
  OAI22_X1 U9223 ( .A1(n8545), .A2(n10051), .B1(n7466), .B2(n8698), .ZN(n7467)
         );
  AOI21_X1 U9224 ( .B1(n8701), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7467), .ZN(
        n7468) );
  OAI211_X1 U9225 ( .C1(n10052), .C2(n8551), .A(n7469), .B(n7468), .ZN(
        P2_U3226) );
  OAI222_X1 U9226 ( .A1(n8064), .A2(n7472), .B1(P1_U3086), .B2(n7471), .C1(
        n9590), .C2(n7470), .ZN(P1_U3335) );
  INV_X1 U9227 ( .A(n7473), .ZN(n7474) );
  NAND2_X1 U9228 ( .A1(n7475), .A2(n7474), .ZN(n7479) );
  NAND2_X1 U9229 ( .A1(n7477), .A2(n7476), .ZN(n7478) );
  NAND2_X1 U9230 ( .A1(n7561), .A2(n7480), .ZN(n9830) );
  OR2_X1 U9231 ( .A1(n9836), .A2(n8966), .ZN(n7481) );
  NAND2_X1 U9232 ( .A1(n7483), .A2(n7482), .ZN(n7567) );
  NAND2_X1 U9233 ( .A1(n7505), .A2(n7506), .ZN(n7485) );
  OR2_X1 U9234 ( .A1(n7512), .A2(n8964), .ZN(n7484) );
  NAND2_X2 U9235 ( .A1(n7485), .A2(n7484), .ZN(n7613) );
  XNOR2_X1 U9236 ( .A(n7613), .B(n7612), .ZN(n9966) );
  INV_X1 U9237 ( .A(n7521), .ZN(n9833) );
  NAND2_X1 U9238 ( .A1(n7486), .A2(n7612), .ZN(n7487) );
  NAND3_X1 U9239 ( .A1(n7488), .A2(n9876), .A3(n7487), .ZN(n7492) );
  NAND2_X1 U9240 ( .A1(n8964), .A2(n8928), .ZN(n7490) );
  NAND2_X1 U9241 ( .A1(n8962), .A2(n8929), .ZN(n7489) );
  NAND2_X1 U9242 ( .A1(n7490), .A2(n7489), .ZN(n7842) );
  INV_X1 U9243 ( .A(n7842), .ZN(n7491) );
  NAND2_X1 U9244 ( .A1(n7492), .A2(n7491), .ZN(n7493) );
  AOI21_X1 U9245 ( .B1(n9966), .B2(n9833), .A(n7493), .ZN(n9968) );
  NOR2_X1 U9246 ( .A1(n9896), .A2(n7494), .ZN(n9840) );
  INV_X1 U9247 ( .A(n9836), .ZN(n9946) );
  INV_X1 U9248 ( .A(n7680), .ZN(n9952) );
  INV_X1 U9249 ( .A(n7512), .ZN(n9959) );
  NAND3_X1 U9250 ( .A1(n7568), .A2(n9952), .A3(n9959), .ZN(n7508) );
  AOI21_X1 U9251 ( .B1(n7508), .B2(n7853), .A(n9481), .ZN(n7495) );
  NAND2_X1 U9252 ( .A1(n7495), .A2(n7615), .ZN(n9963) );
  OAI22_X1 U9253 ( .A1(n9671), .A2(n7496), .B1(n7844), .B2(n9879), .ZN(n7497)
         );
  AOI21_X1 U9254 ( .B1(n7853), .B2(n9835), .A(n7497), .ZN(n7498) );
  OAI21_X1 U9255 ( .B1(n9963), .B2(n9499), .A(n7498), .ZN(n7499) );
  AOI21_X1 U9256 ( .B1(n9966), .B2(n9840), .A(n7499), .ZN(n7500) );
  OAI21_X1 U9257 ( .B1(n9968), .B2(n9881), .A(n7500), .ZN(P1_U3282) );
  XNOR2_X1 U9258 ( .A(n7501), .B(n7506), .ZN(n7504) );
  NAND2_X1 U9259 ( .A1(n8965), .A2(n8928), .ZN(n7503) );
  NAND2_X1 U9260 ( .A1(n8963), .A2(n8929), .ZN(n7502) );
  NAND2_X1 U9261 ( .A1(n7503), .A2(n7502), .ZN(n7761) );
  AOI21_X1 U9262 ( .B1(n7504), .B2(n9876), .A(n7761), .ZN(n9958) );
  XNOR2_X1 U9263 ( .A(n7505), .B(n7506), .ZN(n9961) );
  NAND2_X1 U9264 ( .A1(n9961), .A2(n9893), .ZN(n7514) );
  OAI22_X1 U9265 ( .A1(n9671), .A2(n7507), .B1(n7758), .B2(n9879), .ZN(n7511)
         );
  INV_X1 U9266 ( .A(n7568), .ZN(n9837) );
  OAI21_X1 U9267 ( .B1(n9837), .B2(n7680), .A(n7512), .ZN(n7509) );
  NAND3_X1 U9268 ( .A1(n7509), .A2(n9888), .A3(n7508), .ZN(n9957) );
  NOR2_X1 U9269 ( .A1(n9957), .A2(n9499), .ZN(n7510) );
  AOI211_X1 U9270 ( .C1(n9835), .C2(n7512), .A(n7511), .B(n7510), .ZN(n7513)
         );
  OAI211_X1 U9271 ( .C1(n9896), .C2(n9958), .A(n7514), .B(n7513), .ZN(P1_U3283) );
  INV_X1 U9272 ( .A(n9840), .ZN(n7528) );
  NAND2_X1 U9273 ( .A1(n7518), .A2(n9876), .ZN(n7519) );
  OAI211_X1 U9274 ( .C1(n9905), .C2(n7521), .A(n7520), .B(n7519), .ZN(n9908)
         );
  NAND2_X1 U9275 ( .A1(n9908), .A2(n9671), .ZN(n7527) );
  INV_X1 U9276 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n8976) );
  OAI22_X1 U9277 ( .A1(n9671), .A2(n7522), .B1(n8976), .B2(n9879), .ZN(n7525)
         );
  OAI211_X1 U9278 ( .C1(n9907), .C2(n7523), .A(n9888), .B(n9887), .ZN(n9906)
         );
  NOR2_X1 U9279 ( .A1(n9499), .A2(n9906), .ZN(n7524) );
  AOI211_X1 U9280 ( .C1(n9835), .C2(n4314), .A(n7525), .B(n7524), .ZN(n7526)
         );
  OAI211_X1 U9281 ( .C1(n9905), .C2(n7528), .A(n7527), .B(n7526), .ZN(P1_U3292) );
  INV_X1 U9282 ( .A(n7529), .ZN(n7532) );
  OAI222_X1 U9283 ( .A1(P2_U3151), .A2(n6975), .B1(n8822), .B2(n7532), .C1(
        n7530), .C2(n8824), .ZN(P2_U3274) );
  OAI222_X1 U9284 ( .A1(P1_U3086), .A2(n7533), .B1(n9590), .B2(n7532), .C1(
        n7531), .C2(n8064), .ZN(P1_U3334) );
  XNOR2_X1 U9285 ( .A(n10060), .B(n8037), .ZN(n7591) );
  XNOR2_X1 U9286 ( .A(n7591), .B(n7592), .ZN(n7596) );
  XOR2_X1 U9287 ( .A(n7596), .B(n7597), .Z(n7544) );
  INV_X1 U9288 ( .A(n7631), .ZN(n7541) );
  INV_X1 U9289 ( .A(n7537), .ZN(n7538) );
  AOI21_X1 U9290 ( .B1(n8189), .B2(n8457), .A(n7538), .ZN(n7540) );
  NAND2_X1 U9291 ( .A1(n8200), .A2(n8456), .ZN(n7539) );
  OAI211_X1 U9292 ( .C1(n8031), .C2(n7541), .A(n7540), .B(n7539), .ZN(n7542)
         );
  AOI21_X1 U9293 ( .B1(n10060), .B2(n8176), .A(n7542), .ZN(n7543) );
  OAI21_X1 U9294 ( .B1(n7544), .B2(n8195), .A(n7543), .ZN(P2_U3161) );
  NAND2_X1 U9295 ( .A1(n4412), .A2(n8392), .ZN(n7545) );
  NAND2_X1 U9296 ( .A1(n7546), .A2(n7545), .ZN(n10062) );
  NAND2_X1 U9297 ( .A1(n7625), .A2(n7547), .ZN(n7549) );
  NAND2_X1 U9298 ( .A1(n7549), .A2(n7548), .ZN(n7550) );
  XOR2_X1 U9299 ( .A(n8392), .B(n7550), .Z(n7551) );
  NAND2_X1 U9300 ( .A1(n7551), .A2(n8657), .ZN(n7553) );
  AOI22_X1 U9301 ( .A1(n5090), .A2(n8655), .B1(n8653), .B2(n8455), .ZN(n7552)
         );
  OAI211_X1 U9302 ( .C1(n7554), .C2(n10062), .A(n7553), .B(n7552), .ZN(n10063)
         );
  NAND2_X1 U9303 ( .A1(n10063), .A2(n8699), .ZN(n7558) );
  INV_X1 U9304 ( .A(n7555), .ZN(n7603) );
  OAI22_X1 U9305 ( .A1(n8682), .A2(n9303), .B1(n7603), .B2(n8698), .ZN(n7556)
         );
  AOI21_X1 U9306 ( .B1(n8702), .B2(n10065), .A(n7556), .ZN(n7557) );
  OAI211_X1 U9307 ( .C1(n10062), .C2(n8551), .A(n7558), .B(n7557), .ZN(
        P2_U3224) );
  NAND2_X1 U9308 ( .A1(n7560), .A2(n7559), .ZN(n9829) );
  OR2_X1 U9309 ( .A1(n9829), .A2(n9830), .ZN(n9826) );
  NAND2_X1 U9310 ( .A1(n9826), .A2(n7561), .ZN(n7562) );
  XOR2_X1 U9311 ( .A(n7567), .B(n7562), .Z(n7565) );
  NOR2_X1 U9312 ( .A1(n7563), .A2(n9167), .ZN(n7675) );
  INV_X1 U9313 ( .A(n7675), .ZN(n7564) );
  OAI21_X1 U9314 ( .B1(n7565), .B2(n9828), .A(n7564), .ZN(n9953) );
  INV_X1 U9315 ( .A(n9953), .ZN(n7576) );
  XNOR2_X1 U9316 ( .A(n7566), .B(n7567), .ZN(n9955) );
  XNOR2_X1 U9317 ( .A(n7568), .B(n7680), .ZN(n7570) );
  AND2_X1 U9318 ( .A1(n8964), .A2(n8929), .ZN(n7674) );
  AOI21_X1 U9319 ( .B1(n7570), .B2(n9888), .A(n7674), .ZN(n9951) );
  OAI22_X1 U9320 ( .A1(n9671), .A2(n7571), .B1(n7678), .B2(n9879), .ZN(n7572)
         );
  AOI21_X1 U9321 ( .B1(n7680), .B2(n9835), .A(n7572), .ZN(n7573) );
  OAI21_X1 U9322 ( .B1(n9951), .B2(n9499), .A(n7573), .ZN(n7574) );
  AOI21_X1 U9323 ( .B1(n9955), .B2(n9893), .A(n7574), .ZN(n7575) );
  OAI21_X1 U9324 ( .B1(n7576), .B2(n9881), .A(n7575), .ZN(P1_U3284) );
  XNOR2_X1 U9325 ( .A(n7577), .B(n7578), .ZN(n10075) );
  XNOR2_X1 U9326 ( .A(n7579), .B(n7578), .ZN(n7580) );
  OAI222_X1 U9327 ( .A1(n8695), .A2(n8156), .B1(n8693), .B2(n7581), .C1(n7580), 
        .C2(n10037), .ZN(n10077) );
  NAND2_X1 U9328 ( .A1(n10077), .A2(n8682), .ZN(n7585) );
  INV_X1 U9329 ( .A(n7910), .ZN(n7582) );
  OAI22_X1 U9330 ( .A1(n8699), .A2(n9300), .B1(n7582), .B2(n8698), .ZN(n7583)
         );
  AOI21_X1 U9331 ( .B1(n7900), .B2(n8702), .A(n7583), .ZN(n7584) );
  OAI211_X1 U9332 ( .C1(n8705), .C2(n10075), .A(n7585), .B(n7584), .ZN(
        P2_U3222) );
  INV_X1 U9333 ( .A(n7586), .ZN(n7589) );
  OAI222_X1 U9334 ( .A1(n8064), .A2(n9413), .B1(n9590), .B2(n7589), .C1(
        P1_U3086), .C2(n7587), .ZN(P1_U3333) );
  OAI222_X1 U9335 ( .A1(n7590), .A2(P2_U3151), .B1(n8822), .B2(n7589), .C1(
        n7588), .C2(n8824), .ZN(P2_U3273) );
  INV_X1 U9336 ( .A(n7591), .ZN(n7593) );
  NAND2_X1 U9337 ( .A1(n7593), .A2(n7592), .ZN(n7594) );
  XNOR2_X1 U9338 ( .A(n10065), .B(n8037), .ZN(n7830) );
  XNOR2_X1 U9339 ( .A(n7830), .B(n7831), .ZN(n7598) );
  OAI211_X1 U9340 ( .C1(n7599), .C2(n7598), .A(n7833), .B(n8185), .ZN(n7606)
         );
  AOI21_X1 U9341 ( .B1(n8189), .B2(n5090), .A(n7600), .ZN(n7602) );
  NAND2_X1 U9342 ( .A1(n8200), .A2(n8455), .ZN(n7601) );
  OAI211_X1 U9343 ( .C1(n8031), .C2(n7603), .A(n7602), .B(n7601), .ZN(n7604)
         );
  AOI21_X1 U9344 ( .B1(n10065), .B2(n8176), .A(n7604), .ZN(n7605) );
  NAND2_X1 U9345 ( .A1(n7606), .A2(n7605), .ZN(P2_U3171) );
  XNOR2_X1 U9346 ( .A(n7607), .B(n4837), .ZN(n7610) );
  NAND2_X1 U9347 ( .A1(n8963), .A2(n8928), .ZN(n7609) );
  NAND2_X1 U9348 ( .A1(n8961), .A2(n8929), .ZN(n7608) );
  NAND2_X1 U9349 ( .A1(n7609), .A2(n7608), .ZN(n7775) );
  AOI21_X1 U9350 ( .B1(n7610), .B2(n9876), .A(n7775), .ZN(n9971) );
  INV_X1 U9351 ( .A(n7853), .ZN(n9964) );
  XNOR2_X1 U9352 ( .A(n7690), .B(n7689), .ZN(n9973) );
  NAND2_X1 U9353 ( .A1(n9973), .A2(n9893), .ZN(n7621) );
  OAI22_X1 U9354 ( .A1(n9671), .A2(n7614), .B1(n7772), .B2(n9879), .ZN(n7619)
         );
  INV_X1 U9355 ( .A(n7615), .ZN(n7617) );
  INV_X1 U9356 ( .A(n7693), .ZN(n7616) );
  OAI211_X1 U9357 ( .C1(n4850), .C2(n7617), .A(n7616), .B(n9888), .ZN(n9970)
         );
  NOR2_X1 U9358 ( .A1(n9970), .A2(n9499), .ZN(n7618) );
  AOI211_X1 U9359 ( .C1(n9835), .C2(n6463), .A(n7619), .B(n7618), .ZN(n7620)
         );
  OAI211_X1 U9360 ( .C1(n9896), .C2(n9971), .A(n7621), .B(n7620), .ZN(P1_U3281) );
  NAND2_X1 U9361 ( .A1(n7623), .A2(n7622), .ZN(n7624) );
  XOR2_X1 U9362 ( .A(n8391), .B(n7624), .Z(n10056) );
  INV_X1 U9363 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7630) );
  NAND2_X1 U9364 ( .A1(n7625), .A2(n8256), .ZN(n7627) );
  NAND2_X1 U9365 ( .A1(n7627), .A2(n7626), .ZN(n7628) );
  XOR2_X1 U9366 ( .A(n8391), .B(n7628), .Z(n7629) );
  AOI222_X1 U9367 ( .A1(n8657), .A2(n7629), .B1(n8457), .B2(n8655), .C1(n8456), 
        .C2(n8653), .ZN(n10057) );
  MUX2_X1 U9368 ( .A(n7630), .B(n10057), .S(n8682), .Z(n7633) );
  AOI22_X1 U9369 ( .A1(n8702), .A2(n10060), .B1(n8685), .B2(n7631), .ZN(n7632)
         );
  OAI211_X1 U9370 ( .C1(n10056), .C2(n8705), .A(n7633), .B(n7632), .ZN(
        P2_U3225) );
  INV_X1 U9371 ( .A(n8272), .ZN(n7634) );
  OR2_X1 U9372 ( .A1(n8259), .A2(n7634), .ZN(n8393) );
  XNOR2_X1 U9373 ( .A(n7635), .B(n8393), .ZN(n7638) );
  INV_X1 U9374 ( .A(n7638), .ZN(n10070) );
  XOR2_X1 U9375 ( .A(n8393), .B(n4408), .Z(n7640) );
  OAI22_X1 U9376 ( .A1(n7831), .A2(n8693), .B1(n7661), .B2(n8695), .ZN(n7636)
         );
  AOI21_X1 U9377 ( .B1(n7638), .B2(n7637), .A(n7636), .ZN(n7639) );
  OAI21_X1 U9378 ( .B1(n7640), .B2(n10037), .A(n7639), .ZN(n10072) );
  NAND2_X1 U9379 ( .A1(n10072), .A2(n8699), .ZN(n7645) );
  INV_X1 U9380 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7642) );
  INV_X1 U9381 ( .A(n7641), .ZN(n7837) );
  OAI22_X1 U9382 ( .A1(n8682), .A2(n7642), .B1(n7837), .B2(n8698), .ZN(n7643)
         );
  AOI21_X1 U9383 ( .B1(n8702), .B2(n7839), .A(n7643), .ZN(n7644) );
  OAI211_X1 U9384 ( .C1(n10070), .C2(n8551), .A(n7645), .B(n7644), .ZN(
        P2_U3223) );
  XNOR2_X1 U9385 ( .A(n7646), .B(n7647), .ZN(n7648) );
  NAND2_X1 U9386 ( .A1(n7648), .A2(n7649), .ZN(n7667) );
  OAI21_X1 U9387 ( .B1(n7649), .B2(n7648), .A(n7667), .ZN(n7650) );
  NAND2_X1 U9388 ( .A1(n7650), .A2(n8941), .ZN(n7657) );
  INV_X1 U9389 ( .A(n7651), .ZN(n9834) );
  NAND2_X1 U9390 ( .A1(n8967), .A2(n8928), .ZN(n7653) );
  NAND2_X1 U9391 ( .A1(n8965), .A2(n8929), .ZN(n7652) );
  AND2_X1 U9392 ( .A1(n7653), .A2(n7652), .ZN(n9825) );
  OAI22_X1 U9393 ( .A1(n9825), .A2(n8918), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7654), .ZN(n7655) );
  AOI21_X1 U9394 ( .B1(n9834), .B2(n8921), .A(n7655), .ZN(n7656) );
  OAI211_X1 U9395 ( .C1(n9946), .C2(n8951), .A(n7657), .B(n7656), .ZN(P1_U3221) );
  OAI21_X1 U9396 ( .B1(n4907), .B2(n5540), .A(n7658), .ZN(n10082) );
  XNOR2_X1 U9397 ( .A(n7659), .B(n8284), .ZN(n7660) );
  OAI222_X1 U9398 ( .A1(n8693), .A2(n7661), .B1(n8695), .B2(n8099), .C1(n7660), 
        .C2(n10037), .ZN(n10084) );
  NAND2_X1 U9399 ( .A1(n10084), .A2(n8699), .ZN(n7666) );
  INV_X1 U9400 ( .A(n8101), .ZN(n7662) );
  OAI22_X1 U9401 ( .A1(n8699), .A2(n6291), .B1(n7662), .B2(n8698), .ZN(n7663)
         );
  AOI21_X1 U9402 ( .B1(n7664), .B2(n8702), .A(n7663), .ZN(n7665) );
  OAI211_X1 U9403 ( .C1(n8705), .C2(n10082), .A(n7666), .B(n7665), .ZN(
        P2_U3221) );
  OAI21_X1 U9404 ( .B1(n7668), .B2(n7646), .A(n7667), .ZN(n7673) );
  OAI21_X1 U9405 ( .B1(n7671), .B2(n7670), .A(n7669), .ZN(n7672) );
  XNOR2_X1 U9406 ( .A(n7673), .B(n7672), .ZN(n7682) );
  OAI21_X1 U9407 ( .B1(n7675), .B2(n7674), .A(n8948), .ZN(n7677) );
  OAI211_X1 U9408 ( .C1(n8944), .C2(n7678), .A(n7677), .B(n7676), .ZN(n7679)
         );
  AOI21_X1 U9409 ( .B1(n7680), .B2(n8934), .A(n7679), .ZN(n7681) );
  OAI21_X1 U9410 ( .B1(n7682), .B2(n8923), .A(n7681), .ZN(P1_U3231) );
  INV_X1 U9411 ( .A(n7683), .ZN(n7685) );
  OAI21_X1 U9412 ( .B1(n7685), .B2(n7684), .A(n9810), .ZN(n7688) );
  NAND2_X1 U9413 ( .A1(n8962), .A2(n8928), .ZN(n7687) );
  NAND2_X1 U9414 ( .A1(n8960), .A2(n8929), .ZN(n7686) );
  NAND2_X1 U9415 ( .A1(n7687), .A2(n7686), .ZN(n7740) );
  AOI21_X1 U9416 ( .B1(n7688), .B2(n9876), .A(n7740), .ZN(n9976) );
  XNOR2_X1 U9417 ( .A(n7786), .B(n7785), .ZN(n9980) );
  NAND2_X1 U9418 ( .A1(n9980), .A2(n9893), .ZN(n7698) );
  OAI22_X1 U9419 ( .A1(n9671), .A2(n7691), .B1(n7737), .B2(n9879), .ZN(n7695)
         );
  INV_X1 U9420 ( .A(n9820), .ZN(n7692) );
  OAI211_X1 U9421 ( .C1(n9977), .C2(n7693), .A(n7692), .B(n9888), .ZN(n9975)
         );
  NOR2_X1 U9422 ( .A1(n9975), .A2(n9499), .ZN(n7694) );
  AOI211_X1 U9423 ( .C1(n9835), .C2(n7696), .A(n7695), .B(n7694), .ZN(n7697)
         );
  OAI211_X1 U9424 ( .C1(n9896), .C2(n9976), .A(n7698), .B(n7697), .ZN(P1_U3280) );
  INV_X1 U9425 ( .A(n7699), .ZN(n7703) );
  NAND2_X1 U9426 ( .A1(n8818), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7700) );
  OAI211_X1 U9427 ( .C1(n7703), .C2(n8822), .A(n8441), .B(n7700), .ZN(P2_U3272) );
  NAND2_X1 U9428 ( .A1(n9588), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7701) );
  OAI211_X1 U9429 ( .C1(n7703), .C2(n9590), .A(n7702), .B(n7701), .ZN(P1_U3332) );
  AOI21_X1 U9430 ( .B1(n7706), .B2(n7705), .A(n7704), .ZN(n7721) );
  OAI21_X1 U9431 ( .B1(n7709), .B2(n7708), .A(n7707), .ZN(n7710) );
  AND2_X1 U9432 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7834) );
  AOI21_X1 U9433 ( .B1(n7710), .B2(n10031), .A(n7834), .ZN(n7711) );
  OAI21_X1 U9434 ( .B1(n7712), .B2(n10010), .A(n7711), .ZN(n7718) );
  AOI21_X1 U9435 ( .B1(n7715), .B2(n7714), .A(n7713), .ZN(n7716) );
  NOR2_X1 U9436 ( .A1(n7716), .A2(n10026), .ZN(n7717) );
  AOI211_X1 U9437 ( .C1(n8528), .C2(n7719), .A(n7718), .B(n7717), .ZN(n7720)
         );
  OAI21_X1 U9438 ( .B1(n7721), .B2(n10020), .A(n7720), .ZN(P2_U3192) );
  INV_X1 U9439 ( .A(n7722), .ZN(n8059) );
  OAI222_X1 U9440 ( .A1(n7724), .A2(P1_U3086), .B1(n9590), .B2(n8059), .C1(
        n7723), .C2(n8064), .ZN(P1_U3331) );
  INV_X1 U9441 ( .A(n7725), .ZN(n7914) );
  OAI222_X1 U9442 ( .A1(n7727), .A2(P1_U3086), .B1(n9590), .B2(n7914), .C1(
        n7726), .C2(n8064), .ZN(P1_U3330) );
  NAND2_X1 U9443 ( .A1(n7728), .A2(n7729), .ZN(n7770) );
  NAND2_X1 U9444 ( .A1(n7770), .A2(n7730), .ZN(n7734) );
  AND2_X1 U9445 ( .A1(n7732), .A2(n7731), .ZN(n7733) );
  OAI21_X1 U9446 ( .B1(n7735), .B2(n7734), .A(n7733), .ZN(n7736) );
  NAND2_X1 U9447 ( .A1(n7736), .A2(n8941), .ZN(n7742) );
  NAND2_X1 U9448 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9755) );
  INV_X1 U9449 ( .A(n9755), .ZN(n7739) );
  NOR2_X1 U9450 ( .A1(n8944), .A2(n7737), .ZN(n7738) );
  AOI211_X1 U9451 ( .C1(n8948), .C2(n7740), .A(n7739), .B(n7738), .ZN(n7741)
         );
  OAI211_X1 U9452 ( .C1(n9977), .C2(n8951), .A(n7742), .B(n7741), .ZN(P1_U3234) );
  XNOR2_X1 U9453 ( .A(n7743), .B(n4353), .ZN(n7744) );
  NAND2_X1 U9454 ( .A1(n7744), .A2(n8657), .ZN(n7746) );
  AOI22_X1 U9455 ( .A1(n8453), .A2(n8655), .B1(n8653), .B2(n8451), .ZN(n7745)
         );
  NAND2_X1 U9456 ( .A1(n7746), .A2(n7745), .ZN(n9649) );
  AOI21_X1 U9457 ( .B1(n7747), .B2(n9646), .A(n9649), .ZN(n7752) );
  XNOR2_X1 U9458 ( .A(n7748), .B(n4353), .ZN(n9645) );
  INV_X1 U9459 ( .A(n8158), .ZN(n7749) );
  OAI22_X1 U9460 ( .A1(n8682), .A2(n7864), .B1(n7749), .B2(n8698), .ZN(n7750)
         );
  AOI21_X1 U9461 ( .B1(n9645), .B2(n7211), .A(n7750), .ZN(n7751) );
  OAI21_X1 U9462 ( .B1(n7752), .B2(n8701), .A(n7751), .ZN(P2_U3220) );
  NOR2_X1 U9463 ( .A1(n7753), .A2(n7754), .ZN(n7845) );
  AOI21_X1 U9464 ( .B1(n7753), .B2(n7754), .A(n7845), .ZN(n7755) );
  NAND2_X1 U9465 ( .A1(n7755), .A2(n7756), .ZN(n7848) );
  OAI21_X1 U9466 ( .B1(n7756), .B2(n7755), .A(n7848), .ZN(n7757) );
  NAND2_X1 U9467 ( .A1(n7757), .A2(n8941), .ZN(n7763) );
  NAND2_X1 U9468 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9603) );
  INV_X1 U9469 ( .A(n9603), .ZN(n7760) );
  NOR2_X1 U9470 ( .A1(n8944), .A2(n7758), .ZN(n7759) );
  AOI211_X1 U9471 ( .C1(n8948), .C2(n7761), .A(n7760), .B(n7759), .ZN(n7762)
         );
  OAI211_X1 U9472 ( .C1(n9959), .C2(n8951), .A(n7763), .B(n7762), .ZN(P1_U3217) );
  NAND2_X1 U9473 ( .A1(n7728), .A2(n7764), .ZN(n7849) );
  INV_X1 U9474 ( .A(n7849), .ZN(n7768) );
  INV_X1 U9475 ( .A(n7765), .ZN(n7767) );
  NOR3_X1 U9476 ( .A1(n7768), .A2(n7767), .A3(n7766), .ZN(n7771) );
  OAI21_X1 U9477 ( .B1(n7771), .B2(n4908), .A(n8941), .ZN(n7777) );
  NOR2_X1 U9478 ( .A1(n8944), .A2(n7772), .ZN(n7773) );
  AOI211_X1 U9479 ( .C1(n8948), .C2(n7775), .A(n7774), .B(n7773), .ZN(n7776)
         );
  OAI211_X1 U9480 ( .C1(n4850), .C2(n8951), .A(n7777), .B(n7776), .ZN(P1_U3224) );
  NAND2_X1 U9481 ( .A1(n9807), .A2(n7778), .ZN(n7779) );
  NAND2_X1 U9482 ( .A1(n7779), .A2(n9109), .ZN(n7780) );
  NAND2_X1 U9483 ( .A1(n7780), .A2(n9661), .ZN(n7783) );
  NAND2_X1 U9484 ( .A1(n8960), .A2(n8928), .ZN(n7782) );
  NAND2_X1 U9485 ( .A1(n9111), .A2(n8929), .ZN(n7781) );
  NAND2_X1 U9486 ( .A1(n7782), .A2(n7781), .ZN(n8947) );
  AOI21_X1 U9487 ( .B1(n7783), .B2(n9876), .A(n8947), .ZN(n9688) );
  XNOR2_X1 U9488 ( .A(n9110), .B(n9109), .ZN(n9691) );
  NAND2_X1 U9489 ( .A1(n9691), .A2(n9893), .ZN(n7792) );
  OAI22_X1 U9490 ( .A1(n9671), .A2(n7787), .B1(n8943), .B2(n9879), .ZN(n7789)
         );
  INV_X1 U9491 ( .A(n9817), .ZN(n9984) );
  OAI211_X1 U9492 ( .C1(n9818), .C2(n9689), .A(n9888), .B(n9655), .ZN(n9687)
         );
  NOR2_X1 U9493 ( .A1(n9687), .A2(n9499), .ZN(n7788) );
  AOI211_X1 U9494 ( .C1(n9835), .C2(n7790), .A(n7789), .B(n7788), .ZN(n7791)
         );
  OAI211_X1 U9495 ( .C1(n9881), .C2(n9688), .A(n7792), .B(n7791), .ZN(P1_U3278) );
  INV_X1 U9496 ( .A(n7793), .ZN(n7797) );
  OAI222_X1 U9497 ( .A1(n7795), .A2(P2_U3151), .B1(n8822), .B2(n7797), .C1(
        n7794), .C2(n8824), .ZN(P2_U3269) );
  OAI222_X1 U9498 ( .A1(n7798), .A2(P1_U3086), .B1(n9590), .B2(n7797), .C1(
        n7796), .C2(n8064), .ZN(P1_U3329) );
  AOI21_X1 U9499 ( .B1(n10098), .B2(n7800), .A(n7799), .ZN(n7814) );
  AOI21_X1 U9500 ( .B1(n7802), .B2(n9300), .A(n7801), .ZN(n7810) );
  OAI21_X1 U9501 ( .B1(n7805), .B2(n7804), .A(n7803), .ZN(n7806) );
  AOI22_X1 U9502 ( .A1(n7807), .A2(P2_ADDR_REG_11__SCAN_IN), .B1(n10031), .B2(
        n7806), .ZN(n7809) );
  AND2_X1 U9503 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7907) );
  INV_X1 U9504 ( .A(n7907), .ZN(n7808) );
  OAI211_X1 U9505 ( .C1(n7810), .C2(n10026), .A(n7809), .B(n7808), .ZN(n7811)
         );
  AOI21_X1 U9506 ( .B1(n7812), .B2(n8528), .A(n7811), .ZN(n7813) );
  OAI21_X1 U9507 ( .B1(n7814), .B2(n10020), .A(n7813), .ZN(P2_U3193) );
  NAND2_X1 U9508 ( .A1(n7816), .A2(n7815), .ZN(n7819) );
  INV_X1 U9509 ( .A(n7817), .ZN(n7818) );
  AOI21_X1 U9510 ( .B1(n7820), .B2(n7819), .A(n7818), .ZN(n7826) );
  NAND2_X1 U9511 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U9512 ( .A1(n8961), .A2(n8928), .ZN(n7822) );
  NAND2_X1 U9513 ( .A1(n8959), .A2(n8929), .ZN(n7821) );
  NAND2_X1 U9514 ( .A1(n7822), .A2(n7821), .ZN(n9813) );
  NAND2_X1 U9515 ( .A1(n8948), .A2(n9813), .ZN(n7823) );
  OAI211_X1 U9516 ( .C1(n8944), .C2(n9815), .A(n9775), .B(n7823), .ZN(n7824)
         );
  AOI21_X1 U9517 ( .B1(n9817), .B2(n8934), .A(n7824), .ZN(n7825) );
  OAI21_X1 U9518 ( .B1(n7826), .B2(n8923), .A(n7825), .ZN(P1_U3215) );
  INV_X1 U9519 ( .A(n7827), .ZN(n7873) );
  AOI21_X1 U9520 ( .B1(n8818), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7828), .ZN(
        n7829) );
  OAI21_X1 U9521 ( .B1(n7873), .B2(n8822), .A(n7829), .ZN(P2_U3268) );
  INV_X1 U9522 ( .A(n7830), .ZN(n7832) );
  XNOR2_X1 U9523 ( .A(n10068), .B(n8037), .ZN(n7903) );
  XOR2_X1 U9524 ( .A(n4309), .B(n7903), .Z(n7841) );
  AOI21_X1 U9525 ( .B1(n8189), .B2(n8456), .A(n7834), .ZN(n7836) );
  NAND2_X1 U9526 ( .A1(n8200), .A2(n8454), .ZN(n7835) );
  OAI211_X1 U9527 ( .C1(n8031), .C2(n7837), .A(n7836), .B(n7835), .ZN(n7838)
         );
  AOI21_X1 U9528 ( .B1(n7839), .B2(n8176), .A(n7838), .ZN(n7840) );
  OAI21_X1 U9529 ( .B1(n7841), .B2(n8195), .A(n7840), .ZN(P2_U3157) );
  NAND2_X1 U9530 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9743) );
  NAND2_X1 U9531 ( .A1(n8948), .A2(n7842), .ZN(n7843) );
  OAI211_X1 U9532 ( .C1(n8944), .C2(n7844), .A(n9743), .B(n7843), .ZN(n7852)
         );
  INV_X1 U9533 ( .A(n7845), .ZN(n7846) );
  NAND3_X1 U9534 ( .A1(n7848), .A2(n7847), .A3(n7846), .ZN(n7850) );
  AOI21_X1 U9535 ( .B1(n7850), .B2(n7849), .A(n8923), .ZN(n7851) );
  AOI211_X1 U9536 ( .C1(n7853), .C2(n8934), .A(n7852), .B(n7851), .ZN(n7854)
         );
  INV_X1 U9537 ( .A(n7854), .ZN(P1_U3236) );
  AOI21_X1 U9538 ( .B1(n9650), .B2(n7856), .A(n7855), .ZN(n7872) );
  INV_X1 U9539 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7862) );
  OAI21_X1 U9540 ( .B1(n7859), .B2(n7858), .A(n7857), .ZN(n7860) );
  NAND2_X1 U9541 ( .A1(n7860), .A2(n10031), .ZN(n7861) );
  OAI21_X1 U9542 ( .B1(n10010), .B2(n7862), .A(n7861), .ZN(n7868) );
  AOI21_X1 U9543 ( .B1(n7865), .B2(n7864), .A(n7863), .ZN(n7866) );
  NAND2_X1 U9544 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8154) );
  OAI21_X1 U9545 ( .B1(n10026), .B2(n7866), .A(n8154), .ZN(n7867) );
  NOR2_X1 U9546 ( .A1(n7868), .A2(n7867), .ZN(n7871) );
  NAND2_X1 U9547 ( .A1(n8528), .A2(n7869), .ZN(n7870) );
  OAI211_X1 U9548 ( .C1(n7872), .C2(n10020), .A(n7871), .B(n7870), .ZN(
        P2_U3195) );
  OAI222_X1 U9549 ( .A1(n8064), .A2(n9408), .B1(P1_U3086), .B2(n6707), .C1(
        n9590), .C2(n7873), .ZN(P1_U3328) );
  INV_X1 U9550 ( .A(n7874), .ZN(n8056) );
  AOI21_X1 U9551 ( .B1(n8818), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n7875), .ZN(
        n7876) );
  OAI21_X1 U9552 ( .B1(n8056), .B2(n8822), .A(n7876), .ZN(P2_U3267) );
  AOI21_X1 U9553 ( .B1(n7879), .B2(n7878), .A(n7877), .ZN(n7893) );
  OAI21_X1 U9554 ( .B1(n7882), .B2(n7881), .A(n7880), .ZN(n7883) );
  AND2_X1 U9555 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8097) );
  AOI21_X1 U9556 ( .B1(n7883), .B2(n10031), .A(n8097), .ZN(n7884) );
  OAI21_X1 U9557 ( .B1(n7885), .B2(n10010), .A(n7884), .ZN(n7890) );
  AOI21_X1 U9558 ( .B1(n4401), .B2(n7887), .A(n7886), .ZN(n7888) );
  NOR2_X1 U9559 ( .A1(n7888), .A2(n10026), .ZN(n7889) );
  AOI211_X1 U9560 ( .C1(n8528), .C2(n7891), .A(n7890), .B(n7889), .ZN(n7892)
         );
  OAI21_X1 U9561 ( .B1(n7893), .B2(n10020), .A(n7892), .ZN(P2_U3194) );
  NOR2_X1 U9562 ( .A1(n9640), .A2(n8588), .ZN(n7896) );
  NAND2_X1 U9563 ( .A1(n8292), .A2(n8291), .ZN(n8289) );
  XNOR2_X1 U9564 ( .A(n7894), .B(n8397), .ZN(n7895) );
  OAI222_X1 U9565 ( .A1(n8693), .A2(n8099), .B1(n8695), .B2(n8678), .C1(n7895), 
        .C2(n10037), .ZN(n9641) );
  AOI211_X1 U9566 ( .C1(n8685), .C2(n8070), .A(n7896), .B(n9641), .ZN(n7899)
         );
  XNOR2_X1 U9567 ( .A(n7897), .B(n8397), .ZN(n9643) );
  AOI22_X1 U9568 ( .A1(n9643), .A2(n7211), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n8701), .ZN(n7898) );
  OAI21_X1 U9569 ( .B1(n7899), .B2(n8701), .A(n7898), .ZN(P2_U3219) );
  INV_X1 U9570 ( .A(n7900), .ZN(n10074) );
  INV_X1 U9571 ( .A(n8176), .ZN(n8207) );
  NOR2_X1 U9572 ( .A1(n7901), .A2(n8455), .ZN(n7902) );
  XNOR2_X1 U9573 ( .A(n8396), .B(n8037), .ZN(n7978) );
  INV_X1 U9574 ( .A(n7978), .ZN(n7906) );
  NAND2_X1 U9575 ( .A1(n7905), .A2(n7906), .ZN(n7980) );
  OAI211_X1 U9576 ( .C1(n7905), .C2(n7906), .A(n8185), .B(n7980), .ZN(n7912)
         );
  AOI21_X1 U9577 ( .B1(n8189), .B2(n8455), .A(n7907), .ZN(n7908) );
  OAI21_X1 U9578 ( .B1(n8191), .B2(n8156), .A(n7908), .ZN(n7909) );
  AOI21_X1 U9579 ( .B1(n7910), .B2(n8204), .A(n7909), .ZN(n7911) );
  OAI211_X1 U9580 ( .C1(n10074), .C2(n8207), .A(n7912), .B(n7911), .ZN(
        P2_U3176) );
  OAI222_X1 U9581 ( .A1(n4310), .A2(P2_U3151), .B1(n8822), .B2(n7914), .C1(
        n7913), .C2(n8824), .ZN(P2_U3270) );
  INV_X1 U9582 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n7918) );
  NOR2_X1 U9583 ( .A1(n7916), .A2(n7915), .ZN(n7917) );
  AOI22_X1 U9584 ( .A1(n7919), .A2(n7918), .B1(n7917), .B2(n4310), .ZN(
        P2_U3377) );
  INV_X1 U9585 ( .A(n8210), .ZN(n8821) );
  OAI222_X1 U9586 ( .A1(n8064), .A2(n7921), .B1(n9590), .B2(n8821), .C1(n7920), 
        .C2(P1_U3086), .ZN(P1_U3325) );
  XNOR2_X1 U9587 ( .A(n8380), .B(n8217), .ZN(n7928) );
  XOR2_X1 U9588 ( .A(n7922), .B(n8380), .Z(n7923) );
  OAI222_X1 U9589 ( .A1(n8695), .A2(n4987), .B1(n8693), .B2(n7924), .C1(n10037), .C2(n7923), .ZN(n7929) );
  AOI21_X1 U9590 ( .B1(n10049), .B2(n7928), .A(n7929), .ZN(n7927) );
  AOI22_X1 U9591 ( .A1(n8806), .A2(n7931), .B1(n10087), .B2(
        P2_REG0_REG_1__SCAN_IN), .ZN(n7925) );
  OAI21_X1 U9592 ( .B1(n7927), .B2(n10087), .A(n7925), .ZN(P2_U3393) );
  AOI22_X1 U9593 ( .A1(n8744), .A2(n7931), .B1(n10100), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n7926) );
  OAI21_X1 U9594 ( .B1(n7927), .B2(n10100), .A(n7926), .ZN(P2_U3460) );
  INV_X1 U9595 ( .A(n7928), .ZN(n7934) );
  INV_X1 U9596 ( .A(n7929), .ZN(n7930) );
  MUX2_X1 U9597 ( .A(n6946), .B(n7930), .S(n8682), .Z(n7933) );
  AOI22_X1 U9598 ( .A1(n8702), .A2(n7931), .B1(n8685), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7932) );
  OAI211_X1 U9599 ( .C1(n7934), .C2(n8705), .A(n7933), .B(n7932), .ZN(P2_U3232) );
  NAND2_X1 U9600 ( .A1(n7935), .A2(n8297), .ZN(n8664) );
  XNOR2_X1 U9601 ( .A(n8664), .B(n7937), .ZN(n7950) );
  INV_X1 U9602 ( .A(n10049), .ZN(n10081) );
  INV_X1 U9603 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n7942) );
  INV_X1 U9604 ( .A(n7936), .ZN(n7938) );
  INV_X1 U9605 ( .A(n7937), .ZN(n8298) );
  AOI21_X1 U9606 ( .B1(n7938), .B2(n8298), .A(n10037), .ZN(n7941) );
  OAI22_X1 U9607 ( .A1(n8694), .A2(n8693), .B1(n8644), .B2(n8695), .ZN(n7939)
         );
  AOI21_X1 U9608 ( .B1(n7941), .B2(n7940), .A(n7939), .ZN(n7947) );
  MUX2_X1 U9609 ( .A(n7942), .B(n7947), .S(n10085), .Z(n7944) );
  NAND2_X1 U9610 ( .A1(n7992), .A2(n8806), .ZN(n7943) );
  OAI211_X1 U9611 ( .C1(n7950), .C2(n8814), .A(n7944), .B(n7943), .ZN(P2_U3441) );
  NAND2_X1 U9612 ( .A1(n10103), .A2(n10049), .ZN(n8750) );
  MUX2_X1 U9613 ( .A(n10018), .B(n7947), .S(n10103), .Z(n7946) );
  NAND2_X1 U9614 ( .A1(n7992), .A2(n8744), .ZN(n7945) );
  OAI211_X1 U9615 ( .C1(n8750), .C2(n7950), .A(n7946), .B(n7945), .ZN(P2_U3476) );
  MUX2_X1 U9616 ( .A(n10025), .B(n7947), .S(n8682), .Z(n7949) );
  AOI22_X1 U9617 ( .A1(n7992), .A2(n8702), .B1(n8685), .B2(n8128), .ZN(n7948)
         );
  OAI211_X1 U9618 ( .C1(n7950), .C2(n8705), .A(n7949), .B(n7948), .ZN(P2_U3216) );
  XOR2_X1 U9619 ( .A(n8408), .B(n7952), .Z(n7954) );
  OAI22_X1 U9620 ( .A1(n8046), .A2(n8695), .B1(n8564), .B2(n8693), .ZN(n7953)
         );
  AOI21_X1 U9621 ( .B1(n7954), .B2(n8657), .A(n7953), .ZN(n7961) );
  MUX2_X1 U9622 ( .A(n7955), .B(n7961), .S(n10085), .Z(n7957) );
  NAND2_X1 U9623 ( .A1(n8358), .A2(n8806), .ZN(n7956) );
  OAI211_X1 U9624 ( .C1(n7965), .C2(n8814), .A(n7957), .B(n7956), .ZN(P2_U3455) );
  INV_X1 U9625 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n7958) );
  MUX2_X1 U9626 ( .A(n7958), .B(n7961), .S(n10103), .Z(n7960) );
  NAND2_X1 U9627 ( .A1(n8358), .A2(n8744), .ZN(n7959) );
  OAI211_X1 U9628 ( .C1(n7965), .C2(n8750), .A(n7960), .B(n7959), .ZN(P2_U3487) );
  INV_X1 U9629 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n7962) );
  MUX2_X1 U9630 ( .A(n7962), .B(n7961), .S(n8682), .Z(n7964) );
  AOI22_X1 U9631 ( .A1(n8358), .A2(n8702), .B1(n8685), .B2(n8043), .ZN(n7963)
         );
  OAI211_X1 U9632 ( .C1(n7965), .C2(n8705), .A(n7964), .B(n7963), .ZN(P2_U3205) );
  XOR2_X1 U9633 ( .A(n7971), .B(n8407), .Z(n8559) );
  NAND2_X1 U9634 ( .A1(n7973), .A2(n10085), .ZN(n7975) );
  AOI21_X1 U9635 ( .B1(n8806), .B2(n8556), .A(n7976), .ZN(n7977) );
  INV_X1 U9636 ( .A(n7977), .ZN(P2_U3454) );
  NAND2_X1 U9637 ( .A1(n7978), .A2(n8454), .ZN(n7979) );
  NAND2_X1 U9638 ( .A1(n7980), .A2(n7979), .ZN(n8094) );
  XNOR2_X1 U9639 ( .A(n10080), .B(n8037), .ZN(n7981) );
  XNOR2_X1 U9640 ( .A(n7981), .B(n8453), .ZN(n8096) );
  INV_X1 U9641 ( .A(n7981), .ZN(n7982) );
  NAND2_X1 U9642 ( .A1(n7982), .A2(n8453), .ZN(n7983) );
  XNOR2_X1 U9643 ( .A(n9646), .B(n8037), .ZN(n7985) );
  XNOR2_X1 U9644 ( .A(n7985), .B(n8452), .ZN(n8153) );
  INV_X1 U9645 ( .A(n8153), .ZN(n7984) );
  INV_X1 U9646 ( .A(n7985), .ZN(n7986) );
  NAND2_X1 U9647 ( .A1(n7986), .A2(n8099), .ZN(n7987) );
  NAND2_X1 U9648 ( .A1(n8151), .A2(n7987), .ZN(n8065) );
  XNOR2_X1 U9649 ( .A(n9640), .B(n8037), .ZN(n7988) );
  XNOR2_X1 U9650 ( .A(n7988), .B(n8451), .ZN(n8066) );
  NAND2_X1 U9651 ( .A1(n7988), .A2(n8692), .ZN(n7989) );
  XNOR2_X1 U9652 ( .A(n8748), .B(n8037), .ZN(n7990) );
  XOR2_X1 U9653 ( .A(n8678), .B(n7990), .Z(n8196) );
  INV_X1 U9654 ( .A(n8678), .ZN(n8450) );
  NAND2_X1 U9655 ( .A1(n7990), .A2(n8450), .ZN(n7991) );
  XNOR2_X1 U9656 ( .A(n8115), .B(n8037), .ZN(n7993) );
  XNOR2_X1 U9657 ( .A(n7993), .B(n8694), .ZN(n8113) );
  XNOR2_X1 U9658 ( .A(n7992), .B(n8037), .ZN(n7995) );
  XNOR2_X1 U9659 ( .A(n7995), .B(n8677), .ZN(n8124) );
  INV_X1 U9660 ( .A(n8124), .ZN(n7994) );
  NAND2_X1 U9661 ( .A1(n7993), .A2(n8694), .ZN(n8120) );
  INV_X1 U9662 ( .A(n7995), .ZN(n7996) );
  XNOR2_X1 U9663 ( .A(n8742), .B(n8037), .ZN(n7997) );
  XNOR2_X1 U9664 ( .A(n7997), .B(n8449), .ZN(n8172) );
  NAND2_X1 U9665 ( .A1(n7997), .A2(n8644), .ZN(n7998) );
  NAND2_X1 U9666 ( .A1(n7999), .A2(n7998), .ZN(n8080) );
  XNOR2_X1 U9667 ( .A(n8735), .B(n8037), .ZN(n8000) );
  XNOR2_X1 U9668 ( .A(n8000), .B(n8631), .ZN(n8081) );
  NAND2_X1 U9669 ( .A1(n8080), .A2(n8081), .ZN(n8003) );
  INV_X1 U9670 ( .A(n8000), .ZN(n8001) );
  NAND2_X1 U9671 ( .A1(n8001), .A2(n8631), .ZN(n8002) );
  NAND2_X1 U9672 ( .A1(n8003), .A2(n8002), .ZN(n8143) );
  XNOR2_X1 U9673 ( .A(n8731), .B(n8037), .ZN(n8004) );
  XNOR2_X1 U9674 ( .A(n8004), .B(n8645), .ZN(n8144) );
  INV_X1 U9675 ( .A(n8004), .ZN(n8005) );
  NAND2_X1 U9676 ( .A1(n8005), .A2(n8645), .ZN(n8006) );
  XNOR2_X1 U9677 ( .A(n8624), .B(n8037), .ZN(n8007) );
  XNOR2_X1 U9678 ( .A(n8007), .B(n8632), .ZN(n8088) );
  INV_X1 U9679 ( .A(n8007), .ZN(n8008) );
  XNOR2_X1 U9680 ( .A(n8786), .B(n8037), .ZN(n8163) );
  NOR2_X1 U9681 ( .A1(n8163), .A2(n8447), .ZN(n8009) );
  NAND2_X1 U9682 ( .A1(n8163), .A2(n8447), .ZN(n8011) );
  AND2_X1 U9683 ( .A1(n4906), .A2(n8011), .ZN(n8015) );
  NAND2_X1 U9684 ( .A1(n8016), .A2(n8015), .ZN(n8014) );
  OR2_X1 U9685 ( .A1(n8009), .A2(n4906), .ZN(n8010) );
  NOR2_X1 U9686 ( .A1(n8162), .A2(n8010), .ZN(n8012) );
  NAND2_X1 U9687 ( .A1(n8073), .A2(n8014), .ZN(n8020) );
  XNOR2_X1 U9688 ( .A(n8774), .B(n7363), .ZN(n8017) );
  NAND2_X1 U9689 ( .A1(n8017), .A2(n8596), .ZN(n8021) );
  INV_X1 U9690 ( .A(n8017), .ZN(n8018) );
  NAND2_X1 U9691 ( .A1(n8018), .A2(n8446), .ZN(n8019) );
  NAND2_X1 U9692 ( .A1(n8020), .A2(n8132), .ZN(n8135) );
  NAND2_X1 U9693 ( .A1(n8135), .A2(n8021), .ZN(n8104) );
  XNOR2_X1 U9694 ( .A(n8767), .B(n8037), .ZN(n8022) );
  XNOR2_X1 U9695 ( .A(n8022), .B(n8584), .ZN(n8105) );
  XNOR2_X1 U9696 ( .A(n8711), .B(n8037), .ZN(n8181) );
  INV_X1 U9697 ( .A(n8022), .ZN(n8023) );
  AOI21_X1 U9698 ( .B1(n8181), .B2(n8573), .A(n8183), .ZN(n8024) );
  INV_X1 U9699 ( .A(n8181), .ZN(n8025) );
  NAND2_X1 U9700 ( .A1(n8025), .A2(n8445), .ZN(n8179) );
  NAND2_X1 U9701 ( .A1(n8187), .A2(n8179), .ZN(n8036) );
  XNOR2_X1 U9702 ( .A(n8026), .B(n8037), .ZN(n8048) );
  XNOR2_X1 U9703 ( .A(n8036), .B(n8035), .ZN(n8034) );
  INV_X1 U9704 ( .A(n8027), .ZN(n8554) );
  OAI22_X1 U9705 ( .A1(n8573), .A2(n8202), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8028), .ZN(n8029) );
  AOI21_X1 U9706 ( .B1(n8443), .B2(n8200), .A(n8029), .ZN(n8030) );
  OAI21_X1 U9707 ( .B1(n8554), .B2(n8031), .A(n8030), .ZN(n8032) );
  AOI21_X1 U9708 ( .B1(n8556), .B2(n8176), .A(n8032), .ZN(n8033) );
  OAI21_X1 U9709 ( .B1(n8034), .B2(n8195), .A(n8033), .ZN(P2_U3154) );
  NAND2_X1 U9710 ( .A1(n8036), .A2(n8035), .ZN(n8055) );
  XNOR2_X1 U9711 ( .A(n8443), .B(n8037), .ZN(n8038) );
  XNOR2_X1 U9712 ( .A(n8358), .B(n8038), .ZN(n8047) );
  NAND2_X1 U9713 ( .A1(n8047), .A2(n8185), .ZN(n8054) );
  INV_X1 U9714 ( .A(n8048), .ZN(n8039) );
  NAND2_X1 U9715 ( .A1(n8055), .A2(n8040), .ZN(n8053) );
  INV_X1 U9716 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8041) );
  OAI22_X1 U9717 ( .A1(n8564), .A2(n8202), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8041), .ZN(n8042) );
  INV_X1 U9718 ( .A(n8042), .ZN(n8045) );
  NAND2_X1 U9719 ( .A1(n8043), .A2(n8204), .ZN(n8044) );
  OAI211_X1 U9720 ( .C1(n8046), .C2(n8191), .A(n8045), .B(n8044), .ZN(n8051)
         );
  INV_X1 U9721 ( .A(n8047), .ZN(n8049) );
  NOR4_X1 U9722 ( .A1(n8049), .A2(n8048), .A3(n8564), .A4(n8195), .ZN(n8050)
         );
  AOI211_X1 U9723 ( .C1(n8358), .C2(n8176), .A(n8051), .B(n8050), .ZN(n8052)
         );
  OAI211_X1 U9724 ( .C1(n8055), .C2(n8054), .A(n8053), .B(n8052), .ZN(P2_U3160) );
  OAI222_X1 U9725 ( .A1(n8064), .A2(n8057), .B1(P1_U3086), .B2(n4267), .C1(
        n9590), .C2(n8056), .ZN(P1_U3327) );
  OAI222_X1 U9726 ( .A1(n5590), .A2(P2_U3151), .B1(n8822), .B2(n8059), .C1(
        n8058), .C2(n8824), .ZN(P2_U3271) );
  AOI22_X1 U9727 ( .A1(n8185), .A2(n10035), .B1(n10040), .B2(n8176), .ZN(n8062) );
  NAND2_X1 U9728 ( .A1(n8060), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8061) );
  OAI211_X1 U9729 ( .C1(n6984), .C2(n8191), .A(n8062), .B(n8061), .ZN(P2_U3172) );
  INV_X1 U9730 ( .A(n6446), .ZN(n8826) );
  OAI222_X1 U9731 ( .A1(n8064), .A2(n8063), .B1(P1_U3086), .B2(n5672), .C1(
        n9590), .C2(n8826), .ZN(P1_U3326) );
  XOR2_X1 U9732 ( .A(n8065), .B(n8066), .Z(n8072) );
  NAND2_X1 U9733 ( .A1(n8200), .A2(n8450), .ZN(n8067) );
  NAND2_X1 U9734 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8472) );
  OAI211_X1 U9735 ( .C1(n8099), .C2(n8202), .A(n8067), .B(n8472), .ZN(n8069)
         );
  NOR2_X1 U9736 ( .A1(n9640), .A2(n8207), .ZN(n8068) );
  AOI211_X1 U9737 ( .C1(n8070), .C2(n8204), .A(n8069), .B(n8068), .ZN(n8071)
         );
  OAI21_X1 U9738 ( .B1(n8072), .B2(n8195), .A(n8071), .ZN(P2_U3155) );
  OAI21_X1 U9739 ( .B1(n8585), .B2(n8074), .A(n8073), .ZN(n8075) );
  NAND2_X1 U9740 ( .A1(n8075), .A2(n8185), .ZN(n8079) );
  AOI22_X1 U9741 ( .A1(n8446), .A2(n8200), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8076) );
  OAI21_X1 U9742 ( .B1(n8620), .B2(n8202), .A(n8076), .ZN(n8077) );
  AOI21_X1 U9743 ( .B1(n8598), .B2(n8204), .A(n8077), .ZN(n8078) );
  OAI211_X1 U9744 ( .C1(n8721), .C2(n8207), .A(n8079), .B(n8078), .ZN(P2_U3156) );
  XOR2_X1 U9745 ( .A(n8081), .B(n8080), .Z(n8086) );
  NAND2_X1 U9746 ( .A1(n8204), .A2(n8646), .ZN(n8083) );
  AOI22_X1 U9747 ( .A1(n8200), .A2(n8448), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3151), .ZN(n8082) );
  OAI211_X1 U9748 ( .C1(n8644), .C2(n8202), .A(n8083), .B(n8082), .ZN(n8084)
         );
  AOI21_X1 U9749 ( .B1(n8735), .B2(n8176), .A(n8084), .ZN(n8085) );
  OAI21_X1 U9750 ( .B1(n8086), .B2(n8195), .A(n8085), .ZN(P2_U3159) );
  XOR2_X1 U9751 ( .A(n8088), .B(n8087), .Z(n8093) );
  NAND2_X1 U9752 ( .A1(n8204), .A2(n8623), .ZN(n8090) );
  AOI22_X1 U9753 ( .A1(n8200), .A2(n8447), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8089) );
  OAI211_X1 U9754 ( .C1(n8645), .C2(n8202), .A(n8090), .B(n8089), .ZN(n8091)
         );
  AOI21_X1 U9755 ( .B1(n8624), .B2(n8176), .A(n8091), .ZN(n8092) );
  OAI21_X1 U9756 ( .B1(n8093), .B2(n8195), .A(n8092), .ZN(P2_U3163) );
  OAI211_X1 U9757 ( .C1(n8094), .C2(n8096), .A(n8095), .B(n8185), .ZN(n8103)
         );
  AOI21_X1 U9758 ( .B1(n8189), .B2(n8454), .A(n8097), .ZN(n8098) );
  OAI21_X1 U9759 ( .B1(n8191), .B2(n8099), .A(n8098), .ZN(n8100) );
  AOI21_X1 U9760 ( .B1(n8101), .B2(n8204), .A(n8100), .ZN(n8102) );
  OAI211_X1 U9761 ( .C1(n10080), .C2(n8207), .A(n8103), .B(n8102), .ZN(
        P2_U3164) );
  OAI21_X1 U9762 ( .B1(n8105), .B2(n8104), .A(n8180), .ZN(n8106) );
  NAND2_X1 U9763 ( .A1(n8106), .A2(n8185), .ZN(n8110) );
  AOI22_X1 U9764 ( .A1(n8445), .A2(n8200), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8107) );
  OAI21_X1 U9765 ( .B1(n8596), .B2(n8202), .A(n8107), .ZN(n8108) );
  AOI21_X1 U9766 ( .B1(n8574), .B2(n8204), .A(n8108), .ZN(n8109) );
  OAI211_X1 U9767 ( .C1(n8714), .C2(n8207), .A(n8110), .B(n8109), .ZN(P2_U3165) );
  OR2_X1 U9768 ( .A1(n8111), .A2(n8113), .ZN(n8121) );
  INV_X1 U9769 ( .A(n8121), .ZN(n8112) );
  AOI21_X1 U9770 ( .B1(n8113), .B2(n8111), .A(n8112), .ZN(n8119) );
  NAND2_X1 U9771 ( .A1(n8200), .A2(n5298), .ZN(n8114) );
  NAND2_X1 U9772 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8509) );
  OAI211_X1 U9773 ( .C1(n8678), .C2(n8202), .A(n8114), .B(n8509), .ZN(n8117)
         );
  NOR2_X1 U9774 ( .A1(n8115), .A2(n8207), .ZN(n8116) );
  AOI211_X1 U9775 ( .C1(n8684), .C2(n8204), .A(n8117), .B(n8116), .ZN(n8118)
         );
  OAI21_X1 U9776 ( .B1(n8119), .B2(n8195), .A(n8118), .ZN(P2_U3166) );
  NAND2_X1 U9777 ( .A1(n8121), .A2(n8120), .ZN(n8123) );
  OAI21_X1 U9778 ( .B1(n8124), .B2(n8123), .A(n8122), .ZN(n8125) );
  NAND2_X1 U9779 ( .A1(n8125), .A2(n8185), .ZN(n8130) );
  AOI22_X1 U9780 ( .A1(n8200), .A2(n8449), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n8126) );
  OAI21_X1 U9781 ( .B1(n8694), .B2(n8202), .A(n8126), .ZN(n8127) );
  AOI21_X1 U9782 ( .B1(n8128), .B2(n8204), .A(n8127), .ZN(n8129) );
  OAI211_X1 U9783 ( .C1(n8131), .C2(n8207), .A(n8130), .B(n8129), .ZN(P2_U3168) );
  INV_X1 U9784 ( .A(n8774), .ZN(n8717) );
  INV_X1 U9785 ( .A(n8073), .ZN(n8134) );
  NOR3_X1 U9786 ( .A1(n8134), .A2(n8133), .A3(n8132), .ZN(n8137) );
  INV_X1 U9787 ( .A(n8135), .ZN(n8136) );
  OAI21_X1 U9788 ( .B1(n8137), .B2(n8136), .A(n8185), .ZN(n8142) );
  NOR2_X1 U9789 ( .A1(n8202), .A2(n8585), .ZN(n8140) );
  OAI22_X1 U9790 ( .A1(n8584), .A2(n8191), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8138), .ZN(n8139) );
  AOI211_X1 U9791 ( .C1(n8586), .C2(n8204), .A(n8140), .B(n8139), .ZN(n8141)
         );
  OAI211_X1 U9792 ( .C1(n8717), .C2(n8207), .A(n8142), .B(n8141), .ZN(P2_U3169) );
  XOR2_X1 U9793 ( .A(n8144), .B(n8143), .Z(n8149) );
  NAND2_X1 U9794 ( .A1(n8204), .A2(n8633), .ZN(n8146) );
  INV_X1 U9795 ( .A(n8632), .ZN(n8606) );
  AOI22_X1 U9796 ( .A1(n8200), .A2(n8606), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8145) );
  OAI211_X1 U9797 ( .C1(n8631), .C2(n8202), .A(n8146), .B(n8145), .ZN(n8147)
         );
  AOI21_X1 U9798 ( .B1(n8731), .B2(n8176), .A(n8147), .ZN(n8148) );
  OAI21_X1 U9799 ( .B1(n8149), .B2(n8195), .A(n8148), .ZN(P2_U3173) );
  INV_X1 U9800 ( .A(n8151), .ZN(n8152) );
  AOI21_X1 U9801 ( .B1(n8153), .B2(n8150), .A(n8152), .ZN(n8161) );
  NAND2_X1 U9802 ( .A1(n8200), .A2(n8451), .ZN(n8155) );
  OAI211_X1 U9803 ( .C1(n8156), .C2(n8202), .A(n8155), .B(n8154), .ZN(n8157)
         );
  AOI21_X1 U9804 ( .B1(n8158), .B2(n8204), .A(n8157), .ZN(n8160) );
  NAND2_X1 U9805 ( .A1(n9646), .A2(n8176), .ZN(n8159) );
  OAI211_X1 U9806 ( .C1(n8161), .C2(n8195), .A(n8160), .B(n8159), .ZN(P2_U3174) );
  XNOR2_X1 U9807 ( .A(n8163), .B(n8447), .ZN(n8164) );
  XNOR2_X1 U9808 ( .A(n8162), .B(n8164), .ZN(n8170) );
  INV_X1 U9809 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8165) );
  OAI22_X1 U9810 ( .A1(n8202), .A2(n8632), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8165), .ZN(n8167) );
  NOR2_X1 U9811 ( .A1(n8191), .A2(n8585), .ZN(n8166) );
  AOI211_X1 U9812 ( .C1(n8610), .C2(n8204), .A(n8167), .B(n8166), .ZN(n8169)
         );
  NAND2_X1 U9813 ( .A1(n8786), .A2(n8176), .ZN(n8168) );
  OAI211_X1 U9814 ( .C1(n8170), .C2(n8195), .A(n8169), .B(n8168), .ZN(P2_U3175) );
  XOR2_X1 U9815 ( .A(n8172), .B(n8171), .Z(n8178) );
  NAND2_X1 U9816 ( .A1(n8204), .A2(n8658), .ZN(n8174) );
  INV_X1 U9817 ( .A(n8631), .ZN(n8654) );
  AOI22_X1 U9818 ( .A1(n8200), .A2(n8654), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        P2_U3151), .ZN(n8173) );
  OAI211_X1 U9819 ( .C1(n8677), .C2(n8202), .A(n8174), .B(n8173), .ZN(n8175)
         );
  AOI21_X1 U9820 ( .B1(n8662), .B2(n8176), .A(n8175), .ZN(n8177) );
  OAI21_X1 U9821 ( .B1(n8178), .B2(n8195), .A(n8177), .ZN(P2_U3178) );
  INV_X1 U9822 ( .A(n8179), .ZN(n8188) );
  INV_X1 U9823 ( .A(n8180), .ZN(n8184) );
  XNOR2_X1 U9824 ( .A(n8181), .B(n8573), .ZN(n8182) );
  OAI211_X1 U9825 ( .C1(n8188), .C2(n8187), .A(n8186), .B(n8185), .ZN(n8194)
         );
  AOI22_X1 U9826 ( .A1(n5451), .A2(n8189), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8190) );
  OAI21_X1 U9827 ( .B1(n8564), .B2(n8191), .A(n8190), .ZN(n8192) );
  AOI21_X1 U9828 ( .B1(n8566), .B2(n8204), .A(n8192), .ZN(n8193) );
  OAI211_X1 U9829 ( .C1(n8711), .C2(n8207), .A(n8194), .B(n8193), .ZN(P2_U3180) );
  AOI21_X1 U9830 ( .B1(n8197), .B2(n8196), .A(n8195), .ZN(n8199) );
  NAND2_X1 U9831 ( .A1(n8199), .A2(n8198), .ZN(n8206) );
  AND2_X1 U9832 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8488) );
  AOI21_X1 U9833 ( .B1(n8200), .B2(n5284), .A(n8488), .ZN(n8201) );
  OAI21_X1 U9834 ( .B1(n8692), .B2(n8202), .A(n8201), .ZN(n8203) );
  AOI21_X1 U9835 ( .B1(n8696), .B2(n8204), .A(n8203), .ZN(n8205) );
  OAI211_X1 U9836 ( .C1(n8208), .C2(n8207), .A(n8206), .B(n8205), .ZN(P2_U3181) );
  INV_X1 U9837 ( .A(n8442), .ZN(n8352) );
  OR2_X1 U9838 ( .A1(n4997), .A2(n8820), .ZN(n8211) );
  AOI21_X1 U9839 ( .B1(n8352), .B2(n8355), .A(n8754), .ZN(n8212) );
  AOI21_X1 U9840 ( .B1(n4275), .B2(n8442), .A(n8212), .ZN(n8365) );
  MUX2_X1 U9841 ( .A(n8344), .B(n4611), .S(n4275), .Z(n8213) );
  NOR2_X1 U9842 ( .A1(n8407), .A2(n8213), .ZN(n8351) );
  OAI211_X1 U9843 ( .C1(n8375), .C2(n8446), .A(n8717), .B(n4275), .ZN(n8216)
         );
  NAND3_X1 U9844 ( .A1(n8774), .A2(n8596), .A3(n8355), .ZN(n8215) );
  NAND3_X1 U9845 ( .A1(n8375), .A2(n4275), .A3(n8446), .ZN(n8214) );
  NAND3_X1 U9846 ( .A1(n8216), .A2(n8215), .A3(n8214), .ZN(n8331) );
  INV_X1 U9847 ( .A(n8377), .ZN(n8336) );
  INV_X1 U9848 ( .A(n8299), .ZN(n8302) );
  OAI211_X1 U9849 ( .C1(n8218), .C2(n6975), .A(n5527), .B(n8217), .ZN(n8221)
         );
  NAND2_X1 U9850 ( .A1(n8219), .A2(n8222), .ZN(n8220) );
  MUX2_X1 U9851 ( .A(n8221), .B(n8220), .S(n4275), .Z(n8225) );
  MUX2_X1 U9852 ( .A(n8222), .B(n5527), .S(n4275), .Z(n8223) );
  NAND3_X1 U9853 ( .A1(n8225), .A2(n8224), .A3(n8223), .ZN(n8232) );
  NAND2_X1 U9854 ( .A1(n8237), .A2(n8226), .ZN(n8229) );
  NAND2_X1 U9855 ( .A1(n8243), .A2(n8227), .ZN(n8228) );
  MUX2_X1 U9856 ( .A(n8229), .B(n8228), .S(n8355), .Z(n8230) );
  INV_X1 U9857 ( .A(n8230), .ZN(n8231) );
  NAND2_X1 U9858 ( .A1(n8232), .A2(n8231), .ZN(n8236) );
  OAI211_X1 U9859 ( .C1(n4275), .C2(n8234), .A(n8233), .B(n8244), .ZN(n8235)
         );
  INV_X1 U9860 ( .A(n8237), .ZN(n8239) );
  OAI21_X1 U9861 ( .B1(n8246), .B2(n8239), .A(n8238), .ZN(n8242) );
  INV_X1 U9862 ( .A(n8240), .ZN(n8241) );
  AOI21_X1 U9863 ( .B1(n8242), .B2(n8389), .A(n8241), .ZN(n8252) );
  INV_X1 U9864 ( .A(n8248), .ZN(n8249) );
  AOI21_X1 U9865 ( .B1(n8250), .B2(n8382), .A(n8249), .ZN(n8251) );
  MUX2_X1 U9866 ( .A(n8252), .B(n8251), .S(n4275), .Z(n8258) );
  NAND2_X1 U9867 ( .A1(n8264), .A2(n8263), .ZN(n8255) );
  NAND2_X1 U9868 ( .A1(n8260), .A2(n8253), .ZN(n8254) );
  MUX2_X1 U9869 ( .A(n8255), .B(n8254), .S(n4275), .Z(n8266) );
  NOR2_X1 U9870 ( .A1(n8266), .A2(n8256), .ZN(n8257) );
  NAND2_X1 U9871 ( .A1(n8258), .A2(n8257), .ZN(n8271) );
  INV_X1 U9872 ( .A(n8259), .ZN(n8274) );
  OAI211_X1 U9873 ( .C1(n8266), .C2(n8261), .A(n8274), .B(n8260), .ZN(n8268)
         );
  AND2_X1 U9874 ( .A1(n8263), .A2(n8262), .ZN(n8265) );
  OAI211_X1 U9875 ( .C1(n8266), .C2(n8265), .A(n8264), .B(n8272), .ZN(n8267)
         );
  MUX2_X1 U9876 ( .A(n8268), .B(n8267), .S(n4275), .Z(n8269) );
  INV_X1 U9877 ( .A(n8269), .ZN(n8270) );
  NAND2_X1 U9878 ( .A1(n8271), .A2(n8270), .ZN(n8276) );
  NAND3_X1 U9879 ( .A1(n8276), .A2(n8272), .A3(n8277), .ZN(n8273) );
  NAND2_X1 U9880 ( .A1(n8273), .A2(n8275), .ZN(n8280) );
  NAND3_X1 U9881 ( .A1(n8276), .A2(n8275), .A3(n8274), .ZN(n8278) );
  NAND2_X1 U9882 ( .A1(n8278), .A2(n8277), .ZN(n8279) );
  MUX2_X1 U9883 ( .A(n8282), .B(n8281), .S(n4275), .Z(n8283) );
  INV_X1 U9884 ( .A(n8285), .ZN(n8286) );
  MUX2_X1 U9885 ( .A(n8287), .B(n8286), .S(n4275), .Z(n8288) );
  NOR2_X1 U9886 ( .A1(n8289), .A2(n8288), .ZN(n8290) );
  MUX2_X1 U9887 ( .A(n8292), .B(n8291), .S(n4275), .Z(n8293) );
  NAND2_X1 U9888 ( .A1(n8294), .A2(n8690), .ZN(n8304) );
  NAND3_X1 U9889 ( .A1(n8304), .A2(n8295), .A3(n8305), .ZN(n8296) );
  NAND2_X1 U9890 ( .A1(n8299), .A2(n8666), .ZN(n8378) );
  NAND2_X1 U9891 ( .A1(n8378), .A2(n4275), .ZN(n8300) );
  NAND3_X1 U9892 ( .A1(n8308), .A2(n8311), .A3(n8402), .ZN(n8301) );
  MUX2_X1 U9893 ( .A(n8302), .B(n8301), .S(n4275), .Z(n8318) );
  NAND2_X1 U9894 ( .A1(n8304), .A2(n8303), .ZN(n8306) );
  NAND3_X1 U9895 ( .A1(n8306), .A2(n8355), .A3(n8305), .ZN(n8307) );
  NAND2_X1 U9896 ( .A1(n8308), .A2(n8307), .ZN(n8309) );
  NAND3_X1 U9897 ( .A1(n8309), .A2(n8663), .A3(n8402), .ZN(n8310) );
  NAND2_X1 U9898 ( .A1(n8310), .A2(n8312), .ZN(n8317) );
  NAND2_X1 U9899 ( .A1(n8320), .A2(n8311), .ZN(n8314) );
  INV_X1 U9900 ( .A(n8312), .ZN(n8313) );
  MUX2_X1 U9901 ( .A(n8314), .B(n8313), .S(n4275), .Z(n8315) );
  NOR2_X1 U9902 ( .A1(n8315), .A2(n4602), .ZN(n8316) );
  OAI21_X1 U9903 ( .B1(n8318), .B2(n8317), .A(n8316), .ZN(n8324) );
  AND2_X1 U9904 ( .A1(n8326), .A2(n8319), .ZN(n8322) );
  AND2_X1 U9905 ( .A1(n8332), .A2(n8320), .ZN(n8321) );
  MUX2_X1 U9906 ( .A(n8322), .B(n8321), .S(n4275), .Z(n8323) );
  NAND2_X1 U9907 ( .A1(n8324), .A2(n8323), .ZN(n8333) );
  NAND3_X1 U9908 ( .A1(n8333), .A2(n8604), .A3(n8326), .ZN(n8329) );
  AND2_X1 U9909 ( .A1(n8327), .A2(n4275), .ZN(n8328) );
  NAND4_X1 U9910 ( .A1(n8336), .A2(n8329), .A3(n8337), .A4(n8328), .ZN(n8330)
         );
  NAND2_X1 U9911 ( .A1(n8331), .A2(n8330), .ZN(n8340) );
  NAND3_X1 U9912 ( .A1(n8333), .A2(n8604), .A3(n8332), .ZN(n8335) );
  NAND3_X1 U9913 ( .A1(n8335), .A2(n8375), .A3(n8334), .ZN(n8338) );
  NAND4_X1 U9914 ( .A1(n8338), .A2(n8355), .A3(n8337), .A4(n8336), .ZN(n8339)
         );
  AOI21_X1 U9915 ( .B1(n8340), .B2(n8339), .A(n8571), .ZN(n8348) );
  MUX2_X1 U9916 ( .A(n8342), .B(n8341), .S(n4275), .Z(n8343) );
  INV_X1 U9917 ( .A(n8343), .ZN(n8347) );
  INV_X1 U9918 ( .A(n8344), .ZN(n8346) );
  MUX2_X1 U9919 ( .A(n4368), .B(n8349), .S(n8355), .Z(n8350) );
  MUX2_X1 U9920 ( .A(n8443), .B(n8358), .S(n8355), .Z(n8362) );
  NAND2_X1 U9921 ( .A1(n8417), .A2(n8420), .ZN(n8411) );
  NAND2_X1 U9922 ( .A1(n8754), .A2(n8352), .ZN(n8354) );
  NAND2_X1 U9923 ( .A1(n8354), .A2(n8353), .ZN(n8421) );
  INV_X1 U9924 ( .A(n8356), .ZN(n8357) );
  MUX2_X1 U9925 ( .A(n8443), .B(n8358), .S(n4275), .Z(n8359) );
  AOI211_X2 U9926 ( .C1(n8363), .C2(n8362), .A(n8361), .B(n8360), .ZN(n8364)
         );
  MUX2_X1 U9927 ( .A(n8365), .B(n4275), .S(n8364), .Z(n8415) );
  INV_X1 U9928 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8366) );
  OAI22_X1 U9929 ( .A1(n9591), .A2(n5039), .B1(n8366), .B2(n4997), .ZN(n8416)
         );
  NAND2_X1 U9930 ( .A1(n8367), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8371) );
  NAND2_X1 U9931 ( .A1(n5513), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8370) );
  NAND2_X1 U9932 ( .A1(n8368), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8369) );
  AND3_X1 U9933 ( .A1(n8371), .A2(n8370), .A3(n8369), .ZN(n8372) );
  NOR2_X1 U9934 ( .A1(n8416), .A2(n8418), .ZN(n8429) );
  INV_X1 U9935 ( .A(n8375), .ZN(n8376) );
  NOR2_X1 U9936 ( .A1(n8377), .A2(n8376), .ZN(n8593) );
  INV_X1 U9937 ( .A(n8629), .ZN(n8404) );
  INV_X1 U9938 ( .A(n8378), .ZN(n8401) );
  NOR4_X1 U9939 ( .A1(n8381), .A2(n8380), .A3(n10035), .A4(n8379), .ZN(n8390)
         );
  INV_X1 U9940 ( .A(n8382), .ZN(n8385) );
  NOR4_X1 U9941 ( .A1(n8386), .A2(n8385), .A3(n8384), .A4(n8383), .ZN(n8387)
         );
  NAND4_X1 U9942 ( .A1(n8390), .A2(n8389), .A3(n8388), .A4(n8387), .ZN(n8394)
         );
  NOR4_X1 U9943 ( .A1(n8394), .A2(n8393), .A3(n8392), .A4(n8391), .ZN(n8395)
         );
  NAND4_X1 U9944 ( .A1(n8397), .A2(n5540), .A3(n8396), .A4(n8395), .ZN(n8398)
         );
  NAND4_X1 U9945 ( .A1(n8402), .A2(n8401), .A3(n8400), .A4(n8663), .ZN(n8403)
         );
  NAND4_X1 U9946 ( .A1(n8582), .A2(n8604), .A3(n8593), .A4(n8405), .ZN(n8406)
         );
  NAND2_X1 U9947 ( .A1(n8409), .A2(n8408), .ZN(n8410) );
  NOR4_X1 U9948 ( .A1(n8429), .A2(n8411), .A3(n8421), .A4(n8410), .ZN(n8413)
         );
  INV_X1 U9949 ( .A(n8416), .ZN(n8753) );
  INV_X1 U9950 ( .A(n8417), .ZN(n8419) );
  NOR2_X1 U9951 ( .A1(n8419), .A2(n8418), .ZN(n8428) );
  INV_X1 U9952 ( .A(n8420), .ZN(n8424) );
  INV_X1 U9953 ( .A(n8421), .ZN(n8423) );
  AOI21_X1 U9954 ( .B1(n8753), .B2(n8754), .A(n8429), .ZN(n8422) );
  OAI211_X1 U9955 ( .C1(n8753), .C2(n8428), .A(n8427), .B(n6974), .ZN(n8432)
         );
  INV_X1 U9956 ( .A(n8429), .ZN(n8431) );
  NAND4_X1 U9957 ( .A1(n8437), .A2(n8436), .A3(n8435), .A4(n8434), .ZN(n8438)
         );
  OAI211_X1 U9958 ( .C1(n8439), .C2(n8441), .A(n8438), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8440) );
  MUX2_X1 U9959 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8539), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9960 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8442), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9961 ( .A(n8443), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8463), .Z(
        P2_U3519) );
  MUX2_X1 U9962 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8444), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9963 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8445), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9964 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n5451), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9965 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8446), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9966 ( .A(n8607), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8463), .Z(
        P2_U3514) );
  MUX2_X1 U9967 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8447), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9968 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8606), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9969 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8448), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9970 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8654), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9971 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8449), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9972 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n5298), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9973 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n5284), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9974 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8450), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9975 ( .A(n8451), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8463), .Z(
        P2_U3505) );
  MUX2_X1 U9976 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8452), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9977 ( .A(n8453), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8463), .Z(
        P2_U3503) );
  MUX2_X1 U9978 ( .A(n8454), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8463), .Z(
        P2_U3502) );
  MUX2_X1 U9979 ( .A(n8455), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8463), .Z(
        P2_U3501) );
  MUX2_X1 U9980 ( .A(n8456), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8463), .Z(
        P2_U3500) );
  MUX2_X1 U9981 ( .A(n5090), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8463), .Z(
        P2_U3499) );
  MUX2_X1 U9982 ( .A(n8457), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8463), .Z(
        P2_U3498) );
  MUX2_X1 U9983 ( .A(n8458), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8463), .Z(
        P2_U3497) );
  MUX2_X1 U9984 ( .A(n8459), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8463), .Z(
        P2_U3496) );
  MUX2_X1 U9985 ( .A(n8460), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8463), .Z(
        P2_U3495) );
  MUX2_X1 U9986 ( .A(n8461), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8463), .Z(
        P2_U3494) );
  MUX2_X1 U9987 ( .A(n8462), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8463), .Z(
        P2_U3493) );
  MUX2_X1 U9988 ( .A(n6985), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8463), .Z(
        P2_U3492) );
  MUX2_X1 U9989 ( .A(n8464), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8463), .Z(
        P2_U3491) );
  AOI21_X1 U9990 ( .B1(n4403), .B2(n8466), .A(n8465), .ZN(n8481) );
  INV_X1 U9991 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8473) );
  OAI21_X1 U9992 ( .B1(n8469), .B2(n8468), .A(n8467), .ZN(n8470) );
  NAND2_X1 U9993 ( .A1(n8470), .A2(n10031), .ZN(n8471) );
  OAI211_X1 U9994 ( .C1(n10010), .C2(n8473), .A(n8472), .B(n8471), .ZN(n8478)
         );
  AOI21_X1 U9995 ( .B1(n4404), .B2(n8475), .A(n8474), .ZN(n8476) );
  NOR2_X1 U9996 ( .A1(n8476), .A2(n10026), .ZN(n8477) );
  AOI211_X1 U9997 ( .C1(n8528), .C2(n8479), .A(n8478), .B(n8477), .ZN(n8480)
         );
  OAI21_X1 U9998 ( .B1(n8481), .B2(n10020), .A(n8480), .ZN(P2_U3196) );
  AOI21_X1 U9999 ( .B1(n8484), .B2(n8483), .A(n8482), .ZN(n8499) );
  OAI21_X1 U10000 ( .B1(n8487), .B2(n8486), .A(n8485), .ZN(n8489) );
  AOI21_X1 U10001 ( .B1(n8489), .B2(n10031), .A(n8488), .ZN(n8490) );
  OAI21_X1 U10002 ( .B1(n8491), .B2(n10010), .A(n8490), .ZN(n8496) );
  AOI21_X1 U10003 ( .B1(n9298), .B2(n8493), .A(n8492), .ZN(n8494) );
  NOR2_X1 U10004 ( .A1(n8494), .A2(n10020), .ZN(n8495) );
  AOI211_X1 U10005 ( .C1(n8528), .C2(n8497), .A(n8496), .B(n8495), .ZN(n8498)
         );
  OAI21_X1 U10006 ( .B1(n8499), .B2(n10026), .A(n8498), .ZN(P2_U3197) );
  INV_X1 U10007 ( .A(n8500), .ZN(n8501) );
  AOI21_X1 U10008 ( .B1(n8503), .B2(n8502), .A(n8501), .ZN(n8519) );
  INV_X1 U10009 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8510) );
  OAI21_X1 U10010 ( .B1(n8506), .B2(n8505), .A(n8504), .ZN(n8507) );
  NAND2_X1 U10011 ( .A1(n8507), .A2(n10031), .ZN(n8508) );
  OAI211_X1 U10012 ( .C1(n10010), .C2(n8510), .A(n8509), .B(n8508), .ZN(n8516)
         );
  NAND2_X1 U10013 ( .A1(n8512), .A2(n8511), .ZN(n8513) );
  AOI21_X1 U10014 ( .B1(n8514), .B2(n8513), .A(n10020), .ZN(n8515) );
  AOI211_X1 U10015 ( .C1(n8528), .C2(n8517), .A(n8516), .B(n8515), .ZN(n8518)
         );
  OAI21_X1 U10016 ( .B1(n8519), .B2(n10026), .A(n8518), .ZN(P2_U3198) );
  AOI21_X1 U10017 ( .B1(n8522), .B2(n8521), .A(n8520), .ZN(n8537) );
  INV_X1 U10018 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8535) );
  INV_X1 U10019 ( .A(n8529), .ZN(n8527) );
  NAND2_X1 U10020 ( .A1(n10031), .A2(n8527), .ZN(n8532) );
  AOI21_X1 U10021 ( .B1(P2_U3893), .B2(n8529), .A(n8528), .ZN(n8531) );
  MUX2_X1 U10022 ( .A(n8532), .B(n8531), .S(n8530), .Z(n8534) );
  NAND2_X1 U10023 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3151), .ZN(n8533) );
  OAI211_X1 U10024 ( .C1(n10010), .C2(n8535), .A(n8534), .B(n8533), .ZN(n8536)
         );
  NOR2_X1 U10025 ( .A1(n8540), .A2(n8698), .ZN(n8548) );
  AOI21_X1 U10026 ( .B1(n8751), .B2(n8699), .A(n8548), .ZN(n8542) );
  NAND2_X1 U10027 ( .A1(n8701), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8541) );
  OAI211_X1 U10028 ( .C1(n8753), .C2(n8545), .A(n8542), .B(n8541), .ZN(
        P2_U3202) );
  NAND2_X1 U10029 ( .A1(n8754), .A2(n8702), .ZN(n8543) );
  OAI211_X1 U10030 ( .C1(n8682), .C2(n9399), .A(n8543), .B(n8542), .ZN(
        P2_U3203) );
  NAND2_X1 U10031 ( .A1(n8544), .A2(n8699), .ZN(n8550) );
  NOR2_X1 U10032 ( .A1(n8546), .A2(n8545), .ZN(n8547) );
  AOI211_X1 U10033 ( .C1(n8701), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8548), .B(
        n8547), .ZN(n8549) );
  OAI211_X1 U10034 ( .C1(n8552), .C2(n8551), .A(n8550), .B(n8549), .ZN(
        P2_U3204) );
  OAI21_X1 U10035 ( .B1(n8554), .B2(n8698), .A(n8553), .ZN(n8555) );
  NAND2_X1 U10036 ( .A1(n8555), .A2(n8699), .ZN(n8558) );
  AOI22_X1 U10037 ( .A1(n8556), .A2(n8702), .B1(n8701), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8557) );
  OAI211_X1 U10038 ( .C1(n8559), .C2(n8705), .A(n8558), .B(n8557), .ZN(
        P2_U3206) );
  XNOR2_X1 U10039 ( .A(n8560), .B(n8561), .ZN(n8763) );
  INV_X1 U10040 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8565) );
  XNOR2_X1 U10041 ( .A(n8562), .B(n8561), .ZN(n8563) );
  INV_X1 U10042 ( .A(n8710), .ZN(n8758) );
  MUX2_X1 U10043 ( .A(n8565), .B(n8758), .S(n8682), .Z(n8568) );
  AOI22_X1 U10044 ( .A1(n8760), .A2(n8702), .B1(n8685), .B2(n8566), .ZN(n8567)
         );
  OAI211_X1 U10045 ( .C1(n8763), .C2(n8705), .A(n8568), .B(n8567), .ZN(
        P2_U3207) );
  XNOR2_X1 U10046 ( .A(n8569), .B(n4689), .ZN(n8770) );
  XOR2_X1 U10047 ( .A(n8571), .B(n8570), .Z(n8572) );
  OAI222_X1 U10048 ( .A1(n8693), .A2(n8596), .B1(n8695), .B2(n8573), .C1(
        n10037), .C2(n8572), .ZN(n8764) );
  INV_X1 U10049 ( .A(n8574), .ZN(n8575) );
  OAI22_X1 U10050 ( .A1(n8714), .A2(n8588), .B1(n8575), .B2(n8698), .ZN(n8576)
         );
  OAI21_X1 U10051 ( .B1(n8764), .B2(n8576), .A(n8699), .ZN(n8578) );
  NAND2_X1 U10052 ( .A1(n8701), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8577) );
  OAI211_X1 U10053 ( .C1(n8770), .C2(n8705), .A(n8578), .B(n8577), .ZN(
        P2_U3208) );
  INV_X1 U10054 ( .A(n8582), .ZN(n8579) );
  XNOR2_X1 U10055 ( .A(n8580), .B(n8579), .ZN(n8777) );
  XOR2_X1 U10056 ( .A(n8582), .B(n8581), .Z(n8583) );
  OAI222_X1 U10057 ( .A1(n8693), .A2(n8585), .B1(n8695), .B2(n8584), .C1(
        n10037), .C2(n8583), .ZN(n8771) );
  INV_X1 U10058 ( .A(n8586), .ZN(n8587) );
  OAI22_X1 U10059 ( .A1(n8717), .A2(n8588), .B1(n8587), .B2(n8698), .ZN(n8589)
         );
  OAI21_X1 U10060 ( .B1(n8771), .B2(n8589), .A(n8699), .ZN(n8591) );
  NAND2_X1 U10061 ( .A1(n8701), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8590) );
  OAI211_X1 U10062 ( .C1(n8777), .C2(n8705), .A(n8591), .B(n8590), .ZN(
        P2_U3209) );
  XNOR2_X1 U10063 ( .A(n8592), .B(n8593), .ZN(n8783) );
  INV_X1 U10064 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8597) );
  XNOR2_X1 U10065 ( .A(n8594), .B(n8593), .ZN(n8595) );
  OAI222_X1 U10066 ( .A1(n8695), .A2(n8596), .B1(n8693), .B2(n8620), .C1(
        n10037), .C2(n8595), .ZN(n8720) );
  INV_X1 U10067 ( .A(n8720), .ZN(n8778) );
  MUX2_X1 U10068 ( .A(n8597), .B(n8778), .S(n8682), .Z(n8600) );
  AOI22_X1 U10069 ( .A1(n8780), .A2(n8702), .B1(n8685), .B2(n8598), .ZN(n8599)
         );
  OAI211_X1 U10070 ( .C1(n8783), .C2(n8705), .A(n8600), .B(n8599), .ZN(
        P2_U3210) );
  XNOR2_X1 U10071 ( .A(n8601), .B(n8604), .ZN(n8789) );
  INV_X1 U10072 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8609) );
  NAND3_X1 U10073 ( .A1(n8614), .A2(n8604), .A3(n8603), .ZN(n8605) );
  NAND2_X1 U10074 ( .A1(n8602), .A2(n8605), .ZN(n8608) );
  AOI222_X1 U10075 ( .A1(n8657), .A2(n8608), .B1(n8607), .B2(n8653), .C1(n8606), .C2(n8655), .ZN(n8784) );
  MUX2_X1 U10076 ( .A(n8609), .B(n8784), .S(n8682), .Z(n8612) );
  AOI22_X1 U10077 ( .A1(n8786), .A2(n8702), .B1(n8685), .B2(n8610), .ZN(n8611)
         );
  OAI211_X1 U10078 ( .C1(n8789), .C2(n8705), .A(n8612), .B(n8611), .ZN(
        P2_U3211) );
  XNOR2_X1 U10079 ( .A(n8613), .B(n8615), .ZN(n8793) );
  INV_X1 U10080 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8622) );
  INV_X1 U10081 ( .A(n8614), .ZN(n8618) );
  NOR3_X1 U10082 ( .A1(n4343), .A2(n8616), .A3(n8615), .ZN(n8617) );
  NOR2_X1 U10083 ( .A1(n8618), .A2(n8617), .ZN(n8619) );
  OAI222_X1 U10084 ( .A1(n8693), .A2(n8645), .B1(n8695), .B2(n8620), .C1(
        n10037), .C2(n8619), .ZN(n8790) );
  INV_X1 U10085 ( .A(n8790), .ZN(n8621) );
  MUX2_X1 U10086 ( .A(n8622), .B(n8621), .S(n8682), .Z(n8626) );
  AOI22_X1 U10087 ( .A1(n8624), .A2(n8702), .B1(n8685), .B2(n8623), .ZN(n8625)
         );
  OAI211_X1 U10088 ( .C1(n8793), .C2(n8705), .A(n8626), .B(n8625), .ZN(
        P2_U3212) );
  XNOR2_X1 U10089 ( .A(n8627), .B(n8629), .ZN(n8799) );
  AOI21_X1 U10090 ( .B1(n8629), .B2(n8628), .A(n4343), .ZN(n8630) );
  OAI222_X1 U10091 ( .A1(n8695), .A2(n8632), .B1(n8693), .B2(n8631), .C1(
        n10037), .C2(n8630), .ZN(n8730) );
  NAND2_X1 U10092 ( .A1(n8730), .A2(n8699), .ZN(n8638) );
  INV_X1 U10093 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8635) );
  INV_X1 U10094 ( .A(n8633), .ZN(n8634) );
  OAI22_X1 U10095 ( .A1(n8682), .A2(n8635), .B1(n8634), .B2(n8698), .ZN(n8636)
         );
  AOI21_X1 U10096 ( .B1(n8731), .B2(n8702), .A(n8636), .ZN(n8637) );
  OAI211_X1 U10097 ( .C1(n8799), .C2(n8705), .A(n8638), .B(n8637), .ZN(
        P2_U3213) );
  OAI21_X1 U10098 ( .B1(n8640), .B2(n8641), .A(n8639), .ZN(n8802) );
  XNOR2_X1 U10099 ( .A(n8642), .B(n8641), .ZN(n8643) );
  OAI222_X1 U10100 ( .A1(n8695), .A2(n8645), .B1(n8693), .B2(n8644), .C1(n8643), .C2(n10037), .ZN(n8734) );
  NAND2_X1 U10101 ( .A1(n8734), .A2(n8699), .ZN(n8651) );
  INV_X1 U10102 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8648) );
  INV_X1 U10103 ( .A(n8646), .ZN(n8647) );
  OAI22_X1 U10104 ( .A1(n8682), .A2(n8648), .B1(n8647), .B2(n8698), .ZN(n8649)
         );
  AOI21_X1 U10105 ( .B1(n8735), .B2(n8702), .A(n8649), .ZN(n8650) );
  OAI211_X1 U10106 ( .C1(n8802), .C2(n8705), .A(n8651), .B(n8650), .ZN(
        P2_U3214) );
  XOR2_X1 U10107 ( .A(n8668), .B(n8652), .Z(n8656) );
  AOI222_X1 U10108 ( .A1(n8657), .A2(n8656), .B1(n5298), .B2(n8655), .C1(n8654), .C2(n8653), .ZN(n8741) );
  INV_X1 U10109 ( .A(n8658), .ZN(n8659) );
  OAI22_X1 U10110 ( .A1(n8682), .A2(n8660), .B1(n8659), .B2(n8698), .ZN(n8661)
         );
  AOI21_X1 U10111 ( .B1(n8662), .B2(n8702), .A(n8661), .ZN(n8671) );
  NAND2_X1 U10112 ( .A1(n8664), .A2(n8663), .ZN(n8667) );
  NAND2_X1 U10113 ( .A1(n8667), .A2(n8665), .ZN(n8739) );
  NAND2_X1 U10114 ( .A1(n8667), .A2(n8666), .ZN(n8669) );
  NAND2_X1 U10115 ( .A1(n8669), .A2(n8668), .ZN(n8738) );
  NAND3_X1 U10116 ( .A1(n8739), .A2(n8738), .A3(n7211), .ZN(n8670) );
  OAI211_X1 U10117 ( .C1(n8741), .C2(n8701), .A(n8671), .B(n8670), .ZN(
        P2_U3215) );
  XOR2_X1 U10118 ( .A(n8672), .B(n8674), .Z(n8810) );
  INV_X1 U10119 ( .A(n8673), .ZN(n8676) );
  INV_X1 U10120 ( .A(n8674), .ZN(n8675) );
  AOI21_X1 U10121 ( .B1(n8676), .B2(n8675), .A(n10037), .ZN(n8681) );
  OAI22_X1 U10122 ( .A1(n8678), .A2(n8693), .B1(n8677), .B2(n8695), .ZN(n8679)
         );
  AOI21_X1 U10123 ( .B1(n8681), .B2(n8680), .A(n8679), .ZN(n8804) );
  MUX2_X1 U10124 ( .A(n8683), .B(n8804), .S(n8682), .Z(n8687) );
  AOI22_X1 U10125 ( .A1(n8807), .A2(n8702), .B1(n8685), .B2(n8684), .ZN(n8686)
         );
  OAI211_X1 U10126 ( .C1(n8810), .C2(n8705), .A(n8687), .B(n8686), .ZN(
        P2_U3217) );
  XNOR2_X1 U10127 ( .A(n8688), .B(n8690), .ZN(n8815) );
  XNOR2_X1 U10128 ( .A(n8689), .B(n8690), .ZN(n8691) );
  OAI222_X1 U10129 ( .A1(n8695), .A2(n8694), .B1(n8693), .B2(n8692), .C1(
        n10037), .C2(n8691), .ZN(n8747) );
  INV_X1 U10130 ( .A(n8696), .ZN(n8697) );
  NOR2_X1 U10131 ( .A1(n8698), .A2(n8697), .ZN(n8700) );
  OAI21_X1 U10132 ( .B1(n8747), .B2(n8700), .A(n8699), .ZN(n8704) );
  AOI22_X1 U10133 ( .A1(n8748), .A2(n8702), .B1(P2_REG2_REG_15__SCAN_IN), .B2(
        n8701), .ZN(n8703) );
  OAI211_X1 U10134 ( .C1(n8815), .C2(n8705), .A(n8704), .B(n8703), .ZN(
        P2_U3218) );
  NAND2_X1 U10135 ( .A1(n8751), .A2(n10103), .ZN(n8707) );
  NAND2_X1 U10136 ( .A1(n10100), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8706) );
  OAI211_X1 U10137 ( .C1(n8753), .C2(n8727), .A(n8707), .B(n8706), .ZN(
        P2_U3490) );
  INV_X1 U10138 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U10139 ( .A1(n8754), .A2(n8744), .ZN(n8708) );
  OAI211_X1 U10140 ( .C1(n10103), .C2(n8709), .A(n8708), .B(n8707), .ZN(
        P2_U3489) );
  MUX2_X1 U10141 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8710), .S(n10103), .Z(
        n8713) );
  OAI22_X1 U10142 ( .A1(n8763), .A2(n8750), .B1(n8711), .B2(n8727), .ZN(n8712)
         );
  OR2_X1 U10143 ( .A1(n8713), .A2(n8712), .ZN(P2_U3485) );
  MUX2_X1 U10144 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8764), .S(n10103), .Z(
        n8716) );
  OAI22_X1 U10145 ( .A1(n8770), .A2(n8750), .B1(n8714), .B2(n8727), .ZN(n8715)
         );
  OR2_X1 U10146 ( .A1(n8716), .A2(n8715), .ZN(P2_U3484) );
  MUX2_X1 U10147 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8771), .S(n10103), .Z(
        n8719) );
  OAI22_X1 U10148 ( .A1(n8777), .A2(n8750), .B1(n8717), .B2(n8727), .ZN(n8718)
         );
  OR2_X1 U10149 ( .A1(n8719), .A2(n8718), .ZN(P2_U3483) );
  MUX2_X1 U10150 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8720), .S(n10103), .Z(
        n8723) );
  OAI22_X1 U10151 ( .A1(n8783), .A2(n8750), .B1(n8721), .B2(n8727), .ZN(n8722)
         );
  OR2_X1 U10152 ( .A1(n8723), .A2(n8722), .ZN(P2_U3482) );
  INV_X1 U10153 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8724) );
  MUX2_X1 U10154 ( .A(n8724), .B(n8784), .S(n10103), .Z(n8726) );
  NAND2_X1 U10155 ( .A1(n8786), .A2(n8744), .ZN(n8725) );
  OAI211_X1 U10156 ( .C1(n8789), .C2(n8750), .A(n8726), .B(n8725), .ZN(
        P2_U3481) );
  MUX2_X1 U10157 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8790), .S(n10103), .Z(
        n8729) );
  OAI22_X1 U10158 ( .A1(n8793), .A2(n8750), .B1(n8792), .B2(n8727), .ZN(n8728)
         );
  OR2_X1 U10159 ( .A1(n8729), .A2(n8728), .ZN(P2_U3480) );
  INV_X1 U10160 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8732) );
  AOI21_X1 U10161 ( .B1(n10066), .B2(n8731), .A(n8730), .ZN(n8796) );
  MUX2_X1 U10162 ( .A(n8732), .B(n8796), .S(n10103), .Z(n8733) );
  OAI21_X1 U10163 ( .B1(n8799), .B2(n8750), .A(n8733), .ZN(P2_U3479) );
  INV_X1 U10164 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8736) );
  AOI21_X1 U10165 ( .B1(n10066), .B2(n8735), .A(n8734), .ZN(n8800) );
  MUX2_X1 U10166 ( .A(n8736), .B(n8800), .S(n10103), .Z(n8737) );
  OAI21_X1 U10167 ( .B1(n8750), .B2(n8802), .A(n8737), .ZN(P2_U3478) );
  NAND3_X1 U10168 ( .A1(n8739), .A2(n10049), .A3(n8738), .ZN(n8740) );
  OAI211_X1 U10169 ( .C1(n8742), .C2(n10079), .A(n8741), .B(n8740), .ZN(n8803)
         );
  MUX2_X1 U10170 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8803), .S(n10103), .Z(
        P2_U3477) );
  MUX2_X1 U10171 ( .A(n8743), .B(n8804), .S(n10103), .Z(n8746) );
  NAND2_X1 U10172 ( .A1(n8807), .A2(n8744), .ZN(n8745) );
  OAI211_X1 U10173 ( .C1(n8810), .C2(n8750), .A(n8746), .B(n8745), .ZN(
        P2_U3475) );
  AOI21_X1 U10174 ( .B1(n10066), .B2(n8748), .A(n8747), .ZN(n8811) );
  MUX2_X1 U10175 ( .A(n9298), .B(n8811), .S(n10103), .Z(n8749) );
  OAI21_X1 U10176 ( .B1(n8750), .B2(n8815), .A(n8749), .ZN(P2_U3474) );
  NAND2_X1 U10177 ( .A1(n8751), .A2(n10085), .ZN(n8755) );
  NAND2_X1 U10178 ( .A1(n10087), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8752) );
  OAI211_X1 U10179 ( .C1(n8753), .C2(n8791), .A(n8755), .B(n8752), .ZN(
        P2_U3458) );
  INV_X1 U10180 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8757) );
  NAND2_X1 U10181 ( .A1(n8754), .A2(n8806), .ZN(n8756) );
  OAI211_X1 U10182 ( .C1(n8757), .C2(n10085), .A(n8756), .B(n8755), .ZN(
        P2_U3457) );
  MUX2_X1 U10183 ( .A(n8759), .B(n8758), .S(n10085), .Z(n8762) );
  NAND2_X1 U10184 ( .A1(n8760), .A2(n8806), .ZN(n8761) );
  OAI211_X1 U10185 ( .C1(n8763), .C2(n8814), .A(n8762), .B(n8761), .ZN(
        P2_U3453) );
  INV_X1 U10186 ( .A(n8764), .ZN(n8765) );
  MUX2_X1 U10187 ( .A(n8766), .B(n8765), .S(n10085), .Z(n8769) );
  NAND2_X1 U10188 ( .A1(n8767), .A2(n8806), .ZN(n8768) );
  OAI211_X1 U10189 ( .C1(n8770), .C2(n8814), .A(n8769), .B(n8768), .ZN(
        P2_U3452) );
  INV_X1 U10190 ( .A(n8771), .ZN(n8772) );
  MUX2_X1 U10191 ( .A(n8773), .B(n8772), .S(n10085), .Z(n8776) );
  NAND2_X1 U10192 ( .A1(n8774), .A2(n8806), .ZN(n8775) );
  OAI211_X1 U10193 ( .C1(n8777), .C2(n8814), .A(n8776), .B(n8775), .ZN(
        P2_U3451) );
  MUX2_X1 U10194 ( .A(n8779), .B(n8778), .S(n10085), .Z(n8782) );
  NAND2_X1 U10195 ( .A1(n8780), .A2(n8806), .ZN(n8781) );
  OAI211_X1 U10196 ( .C1(n8783), .C2(n8814), .A(n8782), .B(n8781), .ZN(
        P2_U3450) );
  MUX2_X1 U10197 ( .A(n8785), .B(n8784), .S(n10085), .Z(n8788) );
  NAND2_X1 U10198 ( .A1(n8786), .A2(n8806), .ZN(n8787) );
  OAI211_X1 U10199 ( .C1(n8789), .C2(n8814), .A(n8788), .B(n8787), .ZN(
        P2_U3449) );
  MUX2_X1 U10200 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8790), .S(n10085), .Z(
        n8795) );
  OAI22_X1 U10201 ( .A1(n8793), .A2(n8814), .B1(n8792), .B2(n8791), .ZN(n8794)
         );
  OR2_X1 U10202 ( .A1(n8795), .A2(n8794), .ZN(P2_U3448) );
  INV_X1 U10203 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8797) );
  MUX2_X1 U10204 ( .A(n8797), .B(n8796), .S(n10085), .Z(n8798) );
  OAI21_X1 U10205 ( .B1(n8799), .B2(n8814), .A(n8798), .ZN(P2_U3447) );
  INV_X1 U10206 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9388) );
  MUX2_X1 U10207 ( .A(n9388), .B(n8800), .S(n10085), .Z(n8801) );
  OAI21_X1 U10208 ( .B1(n8802), .B2(n8814), .A(n8801), .ZN(P2_U3446) );
  MUX2_X1 U10209 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8803), .S(n10085), .Z(
        P2_U3444) );
  INV_X1 U10210 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8805) );
  MUX2_X1 U10211 ( .A(n8805), .B(n8804), .S(n10085), .Z(n8809) );
  NAND2_X1 U10212 ( .A1(n8807), .A2(n8806), .ZN(n8808) );
  OAI211_X1 U10213 ( .C1(n8810), .C2(n8814), .A(n8809), .B(n8808), .ZN(
        P2_U3438) );
  INV_X1 U10214 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8812) );
  MUX2_X1 U10215 ( .A(n8812), .B(n8811), .S(n10085), .Z(n8813) );
  OAI21_X1 U10216 ( .B1(n8815), .B2(n8814), .A(n8813), .ZN(P2_U3435) );
  NOR4_X1 U10217 ( .A1(n4926), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n8816), .ZN(n8817) );
  AOI21_X1 U10218 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n8818), .A(n8817), .ZN(
        n8819) );
  OAI21_X1 U10219 ( .B1(n9591), .B2(n8822), .A(n8819), .ZN(P2_U3264) );
  OAI222_X1 U10220 ( .A1(n8823), .A2(P2_U3151), .B1(n8822), .B2(n8821), .C1(
        n8820), .C2(n8824), .ZN(P2_U3265) );
  OAI222_X1 U10221 ( .A1(P2_U3151), .A2(n8827), .B1(n8822), .B2(n8826), .C1(
        n8825), .C2(n8824), .ZN(P2_U3266) );
  MUX2_X1 U10222 ( .A(n8828), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10223 ( .A1(n9125), .A2(n8928), .ZN(n8830) );
  NAND2_X1 U10224 ( .A1(n9130), .A2(n8929), .ZN(n8829) );
  NAND2_X1 U10225 ( .A1(n8830), .A2(n8829), .ZN(n9262) );
  AOI22_X1 U10226 ( .A1(n8948), .A2(n9262), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n8831) );
  OAI21_X1 U10227 ( .B1(n8944), .B2(n9255), .A(n8831), .ZN(n8838) );
  INV_X1 U10228 ( .A(n6181), .ZN(n8836) );
  NAND3_X1 U10229 ( .A1(n8832), .A2(n8834), .A3(n8833), .ZN(n8835) );
  AOI21_X1 U10230 ( .B1(n8836), .B2(n8835), .A(n8923), .ZN(n8837) );
  AOI211_X1 U10231 ( .C1(n9539), .C2(n8934), .A(n8838), .B(n8837), .ZN(n8839)
         );
  INV_X1 U10232 ( .A(n8839), .ZN(P1_U3216) );
  OAI21_X1 U10233 ( .B1(n8841), .B2(n8840), .A(n7024), .ZN(n8842) );
  NAND2_X1 U10234 ( .A1(n8842), .A2(n8941), .ZN(n8846) );
  AOI22_X1 U10235 ( .A1(n8934), .A2(n4271), .B1(n8843), .B2(n8948), .ZN(n8845)
         );
  MUX2_X1 U10236 ( .A(n8944), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n8844) );
  NAND3_X1 U10237 ( .A1(n8846), .A2(n8845), .A3(n8844), .ZN(P1_U3218) );
  XNOR2_X1 U10238 ( .A(n8848), .B(n8847), .ZN(n8849) );
  XNOR2_X1 U10239 ( .A(n8850), .B(n8849), .ZN(n8856) );
  NOR2_X1 U10240 ( .A1(n8944), .A2(n9468), .ZN(n8854) );
  AND2_X1 U10241 ( .A1(n8958), .A2(n8928), .ZN(n8851) );
  AOI21_X1 U10242 ( .B1(n9118), .B2(n8929), .A(n8851), .ZN(n9466) );
  OAI22_X1 U10243 ( .A1(n9466), .A2(n8918), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8852), .ZN(n8853) );
  AOI211_X1 U10244 ( .C1(n9561), .C2(n8934), .A(n8854), .B(n8853), .ZN(n8855)
         );
  OAI21_X1 U10245 ( .B1(n8856), .B2(n8923), .A(n8855), .ZN(P1_U3219) );
  AOI21_X1 U10246 ( .B1(n4316), .B2(n8858), .A(n8857), .ZN(n8864) );
  NAND2_X1 U10247 ( .A1(n9118), .A2(n8928), .ZN(n8860) );
  NAND2_X1 U10248 ( .A1(n9125), .A2(n8929), .ZN(n8859) );
  NAND2_X1 U10249 ( .A1(n8860), .A2(n8859), .ZN(n9285) );
  AOI22_X1 U10250 ( .A1(n9285), .A2(n8948), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n8861) );
  OAI21_X1 U10251 ( .B1(n8944), .B2(n9289), .A(n8861), .ZN(n8862) );
  AOI21_X1 U10252 ( .B1(n9551), .B2(n8934), .A(n8862), .ZN(n8863) );
  OAI21_X1 U10253 ( .B1(n8864), .B2(n8923), .A(n8863), .ZN(P1_U3223) );
  NAND2_X1 U10254 ( .A1(n9530), .A2(n8934), .ZN(n8871) );
  NAND2_X1 U10255 ( .A1(n9130), .A2(n8928), .ZN(n8869) );
  NAND2_X1 U10256 ( .A1(n8957), .A2(n8929), .ZN(n8868) );
  NAND2_X1 U10257 ( .A1(n8869), .A2(n8868), .ZN(n9227) );
  AOI22_X1 U10258 ( .A1(n8948), .A2(n9227), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n8870) );
  OAI211_X1 U10259 ( .C1(n8944), .C2(n9221), .A(n8871), .B(n8870), .ZN(n8872)
         );
  AOI21_X1 U10260 ( .B1(n8873), .B2(n8941), .A(n8872), .ZN(n8874) );
  INV_X1 U10261 ( .A(n8874), .ZN(P1_U3225) );
  OAI21_X1 U10262 ( .B1(n8877), .B2(n8876), .A(n8875), .ZN(n8878) );
  NAND2_X1 U10263 ( .A1(n8878), .A2(n8941), .ZN(n8883) );
  NAND2_X1 U10264 ( .A1(n8959), .A2(n8928), .ZN(n8880) );
  NAND2_X1 U10265 ( .A1(n9112), .A2(n8929), .ZN(n8879) );
  NAND2_X1 U10266 ( .A1(n8880), .A2(n8879), .ZN(n9665) );
  AND2_X1 U10267 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9040) );
  NOR2_X1 U10268 ( .A1(n8944), .A2(n9675), .ZN(n8881) );
  AOI211_X1 U10269 ( .C1(n8948), .C2(n9665), .A(n9040), .B(n8881), .ZN(n8882)
         );
  OAI211_X1 U10270 ( .C1(n9683), .C2(n8951), .A(n8883), .B(n8882), .ZN(
        P1_U3226) );
  INV_X1 U10271 ( .A(n8884), .ZN(n8889) );
  AOI21_X1 U10272 ( .B1(n8886), .B2(n8888), .A(n8885), .ZN(n8887) );
  AOI21_X1 U10273 ( .B1(n8889), .B2(n8888), .A(n8887), .ZN(n8895) );
  NAND2_X1 U10274 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9066) );
  NAND2_X1 U10275 ( .A1(n8958), .A2(n8929), .ZN(n8891) );
  NAND2_X1 U10276 ( .A1(n9111), .A2(n8928), .ZN(n8890) );
  NAND2_X1 U10277 ( .A1(n8891), .A2(n8890), .ZN(n9491) );
  NAND2_X1 U10278 ( .A1(n8948), .A2(n9491), .ZN(n8892) );
  OAI211_X1 U10279 ( .C1(n8944), .C2(n9496), .A(n9066), .B(n8892), .ZN(n8893)
         );
  AOI21_X1 U10280 ( .B1(n9502), .B2(n8934), .A(n8893), .ZN(n8894) );
  OAI21_X1 U10281 ( .B1(n8895), .B2(n8923), .A(n8894), .ZN(P1_U3228) );
  AOI21_X1 U10282 ( .B1(n8896), .B2(n8898), .A(n8897), .ZN(n8903) );
  NOR2_X1 U10283 ( .A1(n8944), .A2(n9452), .ZN(n8901) );
  AND2_X1 U10284 ( .A1(n9115), .A2(n8928), .ZN(n8899) );
  AOI21_X1 U10285 ( .B1(n9121), .B2(n8929), .A(n8899), .ZN(n9447) );
  OAI22_X1 U10286 ( .A1(n9447), .A2(n8918), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9387), .ZN(n8900) );
  AOI211_X1 U10287 ( .C1(n9556), .C2(n8934), .A(n8901), .B(n8900), .ZN(n8902)
         );
  OAI21_X1 U10288 ( .B1(n8903), .B2(n8923), .A(n8902), .ZN(P1_U3233) );
  OAI21_X1 U10289 ( .B1(n8905), .B2(n8904), .A(n8832), .ZN(n8906) );
  NAND2_X1 U10290 ( .A1(n8906), .A2(n8941), .ZN(n8912) );
  INV_X1 U10291 ( .A(n8907), .ZN(n9275) );
  AND2_X1 U10292 ( .A1(n9129), .A2(n8929), .ZN(n8908) );
  AOI21_X1 U10293 ( .B1(n9121), .B2(n8928), .A(n8908), .ZN(n9271) );
  INV_X1 U10294 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8909) );
  OAI22_X1 U10295 ( .A1(n9271), .A2(n8918), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8909), .ZN(n8910) );
  AOI21_X1 U10296 ( .B1(n9275), .B2(n8921), .A(n8910), .ZN(n8911) );
  OAI211_X1 U10297 ( .C1(n9278), .C2(n8951), .A(n8912), .B(n8911), .ZN(
        P1_U3235) );
  XNOR2_X1 U10298 ( .A(n8914), .B(n8913), .ZN(n8915) );
  XNOR2_X1 U10299 ( .A(n8916), .B(n8915), .ZN(n8924) );
  AOI22_X1 U10300 ( .A1(n9115), .A2(n8929), .B1(n9112), .B2(n8928), .ZN(n9477)
         );
  INV_X1 U10301 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8917) );
  OAI22_X1 U10302 ( .A1(n9477), .A2(n8918), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8917), .ZN(n8920) );
  NOR2_X1 U10303 ( .A1(n9485), .A2(n8951), .ZN(n8919) );
  AOI211_X1 U10304 ( .C1(n9482), .C2(n8921), .A(n8920), .B(n8919), .ZN(n8922)
         );
  OAI21_X1 U10305 ( .B1(n8924), .B2(n8923), .A(n8922), .ZN(P1_U3238) );
  NAND2_X1 U10306 ( .A1(n8925), .A2(n8941), .ZN(n8937) );
  AOI21_X1 U10307 ( .B1(n8865), .B2(n8927), .A(n8926), .ZN(n8936) );
  NAND2_X1 U10308 ( .A1(n9132), .A2(n8928), .ZN(n8931) );
  NAND2_X1 U10309 ( .A1(n8956), .A2(n8929), .ZN(n8930) );
  NAND2_X1 U10310 ( .A1(n8931), .A2(n8930), .ZN(n9214) );
  AOI22_X1 U10311 ( .A1(n8948), .A2(n9214), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n8932) );
  OAI21_X1 U10312 ( .B1(n8944), .B2(n9207), .A(n8932), .ZN(n8933) );
  AOI21_X1 U10313 ( .B1(n9525), .B2(n8934), .A(n8933), .ZN(n8935) );
  OAI21_X1 U10314 ( .B1(n8937), .B2(n8936), .A(n8935), .ZN(P1_U3240) );
  OAI21_X1 U10315 ( .B1(n8940), .B2(n8939), .A(n8938), .ZN(n8942) );
  NAND2_X1 U10316 ( .A1(n8942), .A2(n8941), .ZN(n8950) );
  NAND2_X1 U10317 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9785) );
  INV_X1 U10318 ( .A(n9785), .ZN(n8946) );
  NOR2_X1 U10319 ( .A1(n8944), .A2(n8943), .ZN(n8945) );
  AOI211_X1 U10320 ( .C1(n8948), .C2(n8947), .A(n8946), .B(n8945), .ZN(n8949)
         );
  OAI211_X1 U10321 ( .C1(n9689), .C2(n8951), .A(n8950), .B(n8949), .ZN(
        P1_U3241) );
  MUX2_X1 U10322 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n8952), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10323 ( .A(n8953), .B(P1_DATAO_REG_30__SCAN_IN), .S(n8974), .Z(
        P1_U3584) );
  MUX2_X1 U10324 ( .A(n8954), .B(P1_DATAO_REG_29__SCAN_IN), .S(n8974), .Z(
        P1_U3583) );
  MUX2_X1 U10325 ( .A(n8955), .B(P1_DATAO_REG_28__SCAN_IN), .S(n8974), .Z(
        P1_U3582) );
  MUX2_X1 U10326 ( .A(n8956), .B(P1_DATAO_REG_27__SCAN_IN), .S(n8974), .Z(
        P1_U3581) );
  MUX2_X1 U10327 ( .A(n8957), .B(P1_DATAO_REG_26__SCAN_IN), .S(n8974), .Z(
        P1_U3580) );
  MUX2_X1 U10328 ( .A(n9132), .B(P1_DATAO_REG_25__SCAN_IN), .S(n8974), .Z(
        P1_U3579) );
  MUX2_X1 U10329 ( .A(n9130), .B(P1_DATAO_REG_24__SCAN_IN), .S(n8974), .Z(
        P1_U3578) );
  MUX2_X1 U10330 ( .A(n9129), .B(P1_DATAO_REG_23__SCAN_IN), .S(n8974), .Z(
        P1_U3577) );
  MUX2_X1 U10331 ( .A(n9125), .B(P1_DATAO_REG_22__SCAN_IN), .S(n8974), .Z(
        P1_U3576) );
  MUX2_X1 U10332 ( .A(n9121), .B(P1_DATAO_REG_21__SCAN_IN), .S(n8974), .Z(
        P1_U3575) );
  MUX2_X1 U10333 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9118), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10334 ( .A(n9115), .B(P1_DATAO_REG_19__SCAN_IN), .S(n8974), .Z(
        P1_U3573) );
  MUX2_X1 U10335 ( .A(n8958), .B(P1_DATAO_REG_18__SCAN_IN), .S(n8974), .Z(
        P1_U3572) );
  MUX2_X1 U10336 ( .A(n9112), .B(P1_DATAO_REG_17__SCAN_IN), .S(n8974), .Z(
        P1_U3571) );
  MUX2_X1 U10337 ( .A(n9111), .B(P1_DATAO_REG_16__SCAN_IN), .S(n8974), .Z(
        P1_U3570) );
  MUX2_X1 U10338 ( .A(n8959), .B(P1_DATAO_REG_15__SCAN_IN), .S(n8974), .Z(
        P1_U3569) );
  MUX2_X1 U10339 ( .A(n8960), .B(P1_DATAO_REG_14__SCAN_IN), .S(n8974), .Z(
        P1_U3568) );
  MUX2_X1 U10340 ( .A(n8961), .B(P1_DATAO_REG_13__SCAN_IN), .S(n8974), .Z(
        P1_U3567) );
  MUX2_X1 U10341 ( .A(n8962), .B(P1_DATAO_REG_12__SCAN_IN), .S(n8974), .Z(
        P1_U3566) );
  MUX2_X1 U10342 ( .A(n8963), .B(P1_DATAO_REG_11__SCAN_IN), .S(n8974), .Z(
        P1_U3565) );
  MUX2_X1 U10343 ( .A(n8964), .B(P1_DATAO_REG_10__SCAN_IN), .S(n8974), .Z(
        P1_U3564) );
  MUX2_X1 U10344 ( .A(n8965), .B(P1_DATAO_REG_9__SCAN_IN), .S(n8974), .Z(
        P1_U3563) );
  MUX2_X1 U10345 ( .A(n8966), .B(P1_DATAO_REG_8__SCAN_IN), .S(n8974), .Z(
        P1_U3562) );
  MUX2_X1 U10346 ( .A(n8967), .B(P1_DATAO_REG_7__SCAN_IN), .S(n8974), .Z(
        P1_U3561) );
  MUX2_X1 U10347 ( .A(n8968), .B(P1_DATAO_REG_6__SCAN_IN), .S(n8974), .Z(
        P1_U3560) );
  MUX2_X1 U10348 ( .A(n8969), .B(P1_DATAO_REG_5__SCAN_IN), .S(n8974), .Z(
        P1_U3559) );
  MUX2_X1 U10349 ( .A(n8970), .B(P1_DATAO_REG_4__SCAN_IN), .S(n8974), .Z(
        P1_U3558) );
  MUX2_X1 U10350 ( .A(n8971), .B(P1_DATAO_REG_3__SCAN_IN), .S(n8974), .Z(
        P1_U3557) );
  MUX2_X1 U10351 ( .A(n8972), .B(P1_DATAO_REG_2__SCAN_IN), .S(n8974), .Z(
        P1_U3556) );
  MUX2_X1 U10352 ( .A(n8973), .B(P1_DATAO_REG_1__SCAN_IN), .S(n8974), .Z(
        P1_U3555) );
  MUX2_X1 U10353 ( .A(n8975), .B(P1_DATAO_REG_0__SCAN_IN), .S(n8974), .Z(
        P1_U3554) );
  INV_X1 U10354 ( .A(n9773), .ZN(n9801) );
  OAI22_X1 U10355 ( .A1(n9805), .A2(n7393), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8976), .ZN(n8977) );
  AOI21_X1 U10356 ( .B1(n9801), .B2(n8978), .A(n8977), .ZN(n8986) );
  OAI211_X1 U10357 ( .C1(n8981), .C2(n8980), .A(n9763), .B(n8979), .ZN(n8985)
         );
  OAI211_X1 U10358 ( .C1(n8988), .C2(n8983), .A(n9086), .B(n8982), .ZN(n8984)
         );
  NAND3_X1 U10359 ( .A1(n8986), .A2(n8985), .A3(n8984), .ZN(P1_U3244) );
  MUX2_X1 U10360 ( .A(n8989), .B(n8988), .S(n8987), .Z(n8991) );
  NAND2_X1 U10361 ( .A1(n8991), .A2(n8990), .ZN(n8992) );
  OAI211_X1 U10362 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n8993), .A(n8992), .B(
        P1_U3973), .ZN(n9032) );
  INV_X1 U10363 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8994) );
  OAI22_X1 U10364 ( .A1(n9805), .A2(n8994), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9878), .ZN(n8995) );
  AOI21_X1 U10365 ( .B1(n9801), .B2(n8996), .A(n8995), .ZN(n9006) );
  OAI21_X1 U10366 ( .B1(n8999), .B2(n8998), .A(n8997), .ZN(n9000) );
  OR2_X1 U10367 ( .A1(n9795), .A2(n9000), .ZN(n9005) );
  OAI211_X1 U10368 ( .C1(n9003), .C2(n9002), .A(n9763), .B(n9001), .ZN(n9004)
         );
  NAND4_X1 U10369 ( .A1(n9032), .A2(n9006), .A3(n9005), .A4(n9004), .ZN(
        P1_U3245) );
  NAND2_X1 U10370 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9007) );
  OAI21_X1 U10371 ( .B1(n9805), .B2(n9008), .A(n9007), .ZN(n9009) );
  AOI21_X1 U10372 ( .B1(n9801), .B2(n9010), .A(n9009), .ZN(n9019) );
  OAI211_X1 U10373 ( .C1(n9013), .C2(n9012), .A(n9086), .B(n9011), .ZN(n9018)
         );
  OAI211_X1 U10374 ( .C1(n9016), .C2(n9015), .A(n9763), .B(n9014), .ZN(n9017)
         );
  NAND3_X1 U10375 ( .A1(n9019), .A2(n9018), .A3(n9017), .ZN(P1_U3246) );
  INV_X1 U10376 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9020) );
  OAI22_X1 U10377 ( .A1(n9805), .A2(n9020), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9309), .ZN(n9021) );
  AOI21_X1 U10378 ( .B1(n9801), .B2(n9022), .A(n9021), .ZN(n9031) );
  OAI211_X1 U10379 ( .C1(n9025), .C2(n9024), .A(n9763), .B(n9023), .ZN(n9030)
         );
  OAI211_X1 U10380 ( .C1(n9028), .C2(n9027), .A(n9086), .B(n9026), .ZN(n9029)
         );
  NAND4_X1 U10381 ( .A1(n9032), .A2(n9031), .A3(n9030), .A4(n9029), .ZN(
        P1_U3247) );
  MUX2_X1 U10382 ( .A(n9033), .B(P1_REG1_REG_13__SCAN_IN), .S(n9754), .Z(n9747) );
  OAI21_X1 U10383 ( .B1(n9045), .B2(P1_REG1_REG_12__SCAN_IN), .A(n9034), .ZN(
        n9748) );
  NOR2_X1 U10384 ( .A1(n9747), .A2(n9748), .ZN(n9746) );
  AOI21_X1 U10385 ( .B1(n9754), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9746), .ZN(
        n9760) );
  MUX2_X1 U10386 ( .A(n9035), .B(P1_REG1_REG_14__SCAN_IN), .S(n9758), .Z(n9761) );
  NOR2_X1 U10387 ( .A1(n9760), .A2(n9761), .ZN(n9759) );
  AOI21_X1 U10388 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9758), .A(n9759), .ZN(
        n9036) );
  NOR2_X1 U10389 ( .A1(n9036), .A2(n9048), .ZN(n9037) );
  XNOR2_X1 U10390 ( .A(n9048), .B(n9036), .ZN(n9779) );
  NOR2_X1 U10391 ( .A1(n6014), .A2(n9779), .ZN(n9778) );
  NOR2_X1 U10392 ( .A1(n9037), .A2(n9778), .ZN(n9039) );
  AOI22_X1 U10393 ( .A1(n9059), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n6034), .B2(
        n9042), .ZN(n9038) );
  NAND2_X1 U10394 ( .A1(n9038), .A2(n9039), .ZN(n9058) );
  OAI21_X1 U10395 ( .B1(n9039), .B2(n9038), .A(n9058), .ZN(n9055) );
  AOI21_X1 U10396 ( .B1(n9064), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n9040), .ZN(
        n9041) );
  OAI21_X1 U10397 ( .B1(n9042), .B2(n9773), .A(n9041), .ZN(n9054) );
  NAND2_X1 U10398 ( .A1(n9754), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9043) );
  OAI21_X1 U10399 ( .B1(n9754), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9043), .ZN(
        n9750) );
  OAI21_X1 U10400 ( .B1(n9045), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9044), .ZN(
        n9751) );
  NOR2_X1 U10401 ( .A1(n9750), .A2(n9751), .ZN(n9749) );
  NAND2_X1 U10402 ( .A1(n9758), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9046) );
  OAI21_X1 U10403 ( .B1(n9758), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9046), .ZN(
        n9765) );
  NOR2_X1 U10404 ( .A1(n9764), .A2(n9765), .ZN(n9766) );
  NOR2_X1 U10405 ( .A1(n9047), .A2(n9048), .ZN(n9049) );
  XNOR2_X1 U10406 ( .A(n9048), .B(n9047), .ZN(n9781) );
  NOR2_X1 U10407 ( .A1(n7787), .A2(n9781), .ZN(n9780) );
  NAND2_X1 U10408 ( .A1(n9059), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9050) );
  OAI21_X1 U10409 ( .B1(n9059), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9050), .ZN(
        n9051) );
  NOR2_X1 U10410 ( .A1(n9052), .A2(n9051), .ZN(n9057) );
  AOI211_X1 U10411 ( .C1(n9052), .C2(n9051), .A(n9057), .B(n9795), .ZN(n9053)
         );
  AOI211_X1 U10412 ( .C1(n9763), .C2(n9055), .A(n9054), .B(n9053), .ZN(n9056)
         );
  INV_X1 U10413 ( .A(n9056), .ZN(P1_U3259) );
  XNOR2_X1 U10414 ( .A(n9079), .B(n9497), .ZN(n9072) );
  XOR2_X1 U10415 ( .A(n9072), .B(n9073), .Z(n9071) );
  OAI21_X1 U10416 ( .B1(n9059), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9058), .ZN(
        n9063) );
  NOR2_X1 U10417 ( .A1(n9067), .A2(n9060), .ZN(n9061) );
  AOI21_X1 U10418 ( .B1(n9060), .B2(n9067), .A(n9061), .ZN(n9062) );
  NAND2_X1 U10419 ( .A1(n9063), .A2(n9062), .ZN(n9078) );
  OAI21_X1 U10420 ( .B1(n9063), .B2(n9062), .A(n9078), .ZN(n9069) );
  NAND2_X1 U10421 ( .A1(n9064), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9065) );
  OAI211_X1 U10422 ( .C1(n9773), .C2(n9067), .A(n9066), .B(n9065), .ZN(n9068)
         );
  AOI21_X1 U10423 ( .B1(n9069), .B2(n9763), .A(n9068), .ZN(n9070) );
  OAI21_X1 U10424 ( .B1(n9071), .B2(n9795), .A(n9070), .ZN(P1_U3260) );
  NAND2_X1 U10425 ( .A1(n9073), .A2(n9072), .ZN(n9075) );
  OR2_X1 U10426 ( .A1(n9079), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9074) );
  NAND2_X1 U10427 ( .A1(n9075), .A2(n9074), .ZN(n9796) );
  NAND2_X1 U10428 ( .A1(n9800), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9076) );
  OAI21_X1 U10429 ( .B1(n9800), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9076), .ZN(
        n9797) );
  NAND2_X1 U10430 ( .A1(n9793), .A2(n9076), .ZN(n9077) );
  XNOR2_X1 U10431 ( .A(n9077), .B(n9461), .ZN(n9083) );
  OAI21_X1 U10432 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9079), .A(n9078), .ZN(
        n9792) );
  NAND2_X1 U10433 ( .A1(n9800), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9080) );
  OAI21_X1 U10434 ( .B1(n9800), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9080), .ZN(
        n9791) );
  OR2_X1 U10435 ( .A1(n9792), .A2(n9791), .ZN(n9788) );
  NAND2_X1 U10436 ( .A1(n9788), .A2(n9080), .ZN(n9082) );
  XNOR2_X1 U10437 ( .A(n9082), .B(n9081), .ZN(n9084) );
  AOI22_X1 U10438 ( .A1(n9083), .A2(n9086), .B1(n9763), .B2(n9084), .ZN(n9089)
         );
  INV_X1 U10439 ( .A(n9083), .ZN(n9087) );
  INV_X1 U10440 ( .A(n9763), .ZN(n9790) );
  OAI21_X1 U10441 ( .B1(n9084), .B2(n9790), .A(n9773), .ZN(n9085) );
  AOI21_X1 U10442 ( .B1(n9087), .B2(n9086), .A(n9085), .ZN(n9088) );
  NAND2_X1 U10443 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9090) );
  OAI211_X1 U10444 ( .C1(n4935), .C2(n9805), .A(n9091), .B(n9090), .ZN(
        P1_U3262) );
  INV_X1 U10445 ( .A(n9525), .ZN(n9210) );
  NOR2_X2 U10446 ( .A1(n9479), .A2(n9561), .ZN(n9449) );
  NAND2_X1 U10447 ( .A1(n9210), .A2(n9220), .ZN(n9204) );
  NOR2_X2 U10448 ( .A1(n9204), .A2(n9521), .ZN(n9176) );
  NAND2_X1 U10449 ( .A1(n9508), .A2(n9142), .ZN(n9102) );
  INV_X1 U10450 ( .A(P1_B_REG_SCAN_IN), .ZN(n9096) );
  OR2_X1 U10451 ( .A1(n6707), .A2(n9096), .ZN(n9097) );
  NAND2_X1 U10452 ( .A1(n8929), .A2(n9097), .ZN(n9166) );
  OR2_X1 U10453 ( .A1(n9098), .A2(n9166), .ZN(n9506) );
  NOR2_X1 U10454 ( .A1(n9506), .A2(n9881), .ZN(n9104) );
  NOR2_X1 U10455 ( .A1(n9094), .A2(n9883), .ZN(n9100) );
  AOI211_X1 U10456 ( .C1(n9881), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9104), .B(
        n9100), .ZN(n9101) );
  OAI21_X1 U10457 ( .B1(n9505), .B2(n9499), .A(n9101), .ZN(P1_U3263) );
  OAI211_X1 U10458 ( .C1(n9508), .C2(n9142), .A(n9888), .B(n9102), .ZN(n9507)
         );
  AND2_X1 U10459 ( .A1(n9881), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9103) );
  NOR2_X1 U10460 ( .A1(n9104), .A2(n9103), .ZN(n9107) );
  NAND2_X1 U10461 ( .A1(n9105), .A2(n9835), .ZN(n9106) );
  OAI211_X1 U10462 ( .C1(n9507), .C2(n9499), .A(n9107), .B(n9106), .ZN(
        P1_U3264) );
  NAND2_X1 U10463 ( .A1(n9495), .A2(n9494), .ZN(n9493) );
  INV_X1 U10464 ( .A(n9561), .ZN(n9462) );
  NAND2_X1 U10465 ( .A1(n9462), .A2(n9114), .ZN(n9117) );
  NAND2_X1 U10466 ( .A1(n9442), .A2(n9445), .ZN(n9441) );
  NAND2_X1 U10467 ( .A1(n9441), .A2(n9119), .ZN(n9281) );
  INV_X1 U10468 ( .A(n9551), .ZN(n9293) );
  NAND2_X1 U10469 ( .A1(n9281), .A2(n4901), .ZN(n9123) );
  NAND2_X1 U10470 ( .A1(n9123), .A2(n9122), .ZN(n9268) );
  NAND2_X1 U10471 ( .A1(n9268), .A2(n4900), .ZN(n9127) );
  NAND2_X1 U10472 ( .A1(n9530), .A2(n9132), .ZN(n9135) );
  INV_X1 U10473 ( .A(n9530), .ZN(n9224) );
  INV_X1 U10474 ( .A(n9136), .ZN(n9137) );
  NAND2_X1 U10475 ( .A1(n9515), .A2(n8955), .ZN(n9140) );
  NAND2_X1 U10476 ( .A1(n9174), .A2(n9140), .ZN(n9141) );
  INV_X1 U10477 ( .A(n9510), .ZN(n9146) );
  INV_X1 U10478 ( .A(n9143), .ZN(n9144) );
  AOI22_X1 U10479 ( .A1(n9881), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9144), .B2(
        n9847), .ZN(n9145) );
  OAI21_X1 U10480 ( .B1(n9146), .B2(n9883), .A(n9145), .ZN(n9147) );
  AOI21_X1 U10481 ( .B1(n9509), .B2(n9892), .A(n9147), .ZN(n9173) );
  INV_X1 U10482 ( .A(n9148), .ZN(n9149) );
  INV_X1 U10483 ( .A(n9150), .ZN(n9151) );
  NAND2_X1 U10484 ( .A1(n9245), .A2(n9154), .ZN(n9244) );
  INV_X1 U10485 ( .A(n9156), .ZN(n9157) );
  INV_X1 U10486 ( .A(n9161), .ZN(n9162) );
  XNOR2_X1 U10487 ( .A(n9164), .B(n9163), .ZN(n9171) );
  INV_X1 U10488 ( .A(n9169), .ZN(n9170) );
  NAND2_X1 U10489 ( .A1(n9512), .A2(n9671), .ZN(n9172) );
  OAI211_X1 U10490 ( .C1(n9513), .C2(n9488), .A(n9173), .B(n9172), .ZN(
        P1_U3356) );
  OAI21_X1 U10491 ( .B1(n9175), .B2(n9181), .A(n9174), .ZN(n9518) );
  AOI211_X1 U10492 ( .C1(n9515), .C2(n9196), .A(n9481), .B(n4359), .ZN(n9514)
         );
  INV_X1 U10493 ( .A(n9177), .ZN(n9178) );
  AOI22_X1 U10494 ( .A1(n9881), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9178), .B2(
        n9847), .ZN(n9179) );
  OAI21_X1 U10495 ( .B1(n9093), .B2(n9883), .A(n9179), .ZN(n9185) );
  AOI211_X1 U10496 ( .C1(n9181), .C2(n9180), .A(n9828), .B(n4363), .ZN(n9183)
         );
  NOR2_X1 U10497 ( .A1(n9183), .A2(n9182), .ZN(n9517) );
  NOR2_X1 U10498 ( .A1(n9517), .A2(n9881), .ZN(n9184) );
  AOI211_X1 U10499 ( .C1(n9514), .C2(n9892), .A(n9185), .B(n9184), .ZN(n9186)
         );
  OAI21_X1 U10500 ( .B1(n9518), .B2(n9488), .A(n9186), .ZN(P1_U3265) );
  XNOR2_X1 U10501 ( .A(n9187), .B(n9191), .ZN(n9523) );
  INV_X1 U10502 ( .A(n9189), .ZN(n9190) );
  AOI211_X1 U10503 ( .C1(n9188), .C2(n9192), .A(n9191), .B(n9190), .ZN(n9193)
         );
  OAI21_X1 U10504 ( .B1(n9195), .B2(n9828), .A(n9194), .ZN(n9519) );
  AOI211_X1 U10505 ( .C1(n9521), .C2(n9204), .A(n9481), .B(n9176), .ZN(n9520)
         );
  NAND2_X1 U10506 ( .A1(n9520), .A2(n9892), .ZN(n9199) );
  AOI22_X1 U10507 ( .A1(n9881), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9197), .B2(
        n9847), .ZN(n9198) );
  OAI211_X1 U10508 ( .C1(n9200), .C2(n9883), .A(n9199), .B(n9198), .ZN(n9201)
         );
  AOI21_X1 U10509 ( .B1(n9519), .B2(n9671), .A(n9201), .ZN(n9202) );
  OAI21_X1 U10510 ( .B1(n9523), .B2(n9488), .A(n9202), .ZN(P1_U3266) );
  XOR2_X1 U10511 ( .A(n9213), .B(n9203), .Z(n9528) );
  INV_X1 U10512 ( .A(n9220), .ZN(n9206) );
  INV_X1 U10513 ( .A(n9204), .ZN(n9205) );
  AOI211_X1 U10514 ( .C1(n9525), .C2(n9206), .A(n9481), .B(n9205), .ZN(n9524)
         );
  INV_X1 U10515 ( .A(n9207), .ZN(n9208) );
  AOI22_X1 U10516 ( .A1(n9881), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9208), .B2(
        n9847), .ZN(n9209) );
  OAI21_X1 U10517 ( .B1(n9210), .B2(n9883), .A(n9209), .ZN(n9217) );
  NOR2_X1 U10518 ( .A1(n9188), .A2(n9211), .ZN(n9212) );
  XOR2_X1 U10519 ( .A(n9213), .B(n9212), .Z(n9215) );
  AOI21_X1 U10520 ( .B1(n9215), .B2(n9876), .A(n9214), .ZN(n9527) );
  NOR2_X1 U10521 ( .A1(n9527), .A2(n9881), .ZN(n9216) );
  AOI211_X1 U10522 ( .C1(n9524), .C2(n9892), .A(n9217), .B(n9216), .ZN(n9218)
         );
  OAI21_X1 U10523 ( .B1(n9528), .B2(n9488), .A(n9218), .ZN(P1_U3267) );
  XNOR2_X1 U10524 ( .A(n9219), .B(n9226), .ZN(n9533) );
  AOI211_X1 U10525 ( .C1(n9530), .C2(n9237), .A(n9481), .B(n9220), .ZN(n9529)
         );
  INV_X1 U10526 ( .A(n9221), .ZN(n9222) );
  AOI22_X1 U10527 ( .A1(n9896), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9222), .B2(
        n9847), .ZN(n9223) );
  OAI21_X1 U10528 ( .B1(n9224), .B2(n9883), .A(n9223), .ZN(n9230) );
  XOR2_X1 U10529 ( .A(n9226), .B(n9225), .Z(n9228) );
  AOI21_X1 U10530 ( .B1(n9228), .B2(n9876), .A(n9227), .ZN(n9532) );
  NOR2_X1 U10531 ( .A1(n9532), .A2(n9896), .ZN(n9229) );
  AOI211_X1 U10532 ( .C1(n9529), .C2(n9892), .A(n9230), .B(n9229), .ZN(n9231)
         );
  OAI21_X1 U10533 ( .B1(n9533), .B2(n9488), .A(n9231), .ZN(P1_U3268) );
  OAI21_X1 U10534 ( .B1(n9234), .B2(n9233), .A(n9232), .ZN(n9235) );
  INV_X1 U10535 ( .A(n9235), .ZN(n9538) );
  INV_X1 U10536 ( .A(n9237), .ZN(n9238) );
  AOI211_X1 U10537 ( .C1(n9536), .C2(n9254), .A(n9481), .B(n9238), .ZN(n9535)
         );
  INV_X1 U10538 ( .A(n9536), .ZN(n9239) );
  NOR2_X1 U10539 ( .A1(n9239), .A2(n9883), .ZN(n9243) );
  OAI22_X1 U10540 ( .A1(n9671), .A2(n9241), .B1(n9240), .B2(n9879), .ZN(n9242)
         );
  AOI211_X1 U10541 ( .C1(n9535), .C2(n9892), .A(n9243), .B(n9242), .ZN(n9252)
         );
  NAND2_X1 U10542 ( .A1(n9244), .A2(n9876), .ZN(n9250) );
  AOI21_X1 U10543 ( .B1(n9259), .B2(n4340), .A(n9246), .ZN(n9249) );
  INV_X1 U10544 ( .A(n9247), .ZN(n9248) );
  OAI21_X1 U10545 ( .B1(n9250), .B2(n9249), .A(n9248), .ZN(n9534) );
  NAND2_X1 U10546 ( .A1(n9534), .A2(n9671), .ZN(n9251) );
  OAI211_X1 U10547 ( .C1(n9538), .C2(n9488), .A(n9252), .B(n9251), .ZN(
        P1_U3269) );
  XNOR2_X1 U10548 ( .A(n9253), .B(n9260), .ZN(n9543) );
  AOI21_X1 U10549 ( .B1(n9539), .B2(n9273), .A(n9236), .ZN(n9540) );
  INV_X1 U10550 ( .A(n9255), .ZN(n9256) );
  AOI22_X1 U10551 ( .A1(n9896), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9256), .B2(
        n9847), .ZN(n9257) );
  OAI21_X1 U10552 ( .B1(n9258), .B2(n9883), .A(n9257), .ZN(n9265) );
  OAI21_X1 U10553 ( .B1(n9261), .B2(n9260), .A(n9259), .ZN(n9263) );
  AOI21_X1 U10554 ( .B1(n9263), .B2(n9876), .A(n9262), .ZN(n9542) );
  NOR2_X1 U10555 ( .A1(n9542), .A2(n9881), .ZN(n9264) );
  AOI211_X1 U10556 ( .C1(n9540), .C2(n9266), .A(n9265), .B(n9264), .ZN(n9267)
         );
  OAI21_X1 U10557 ( .B1(n9488), .B2(n9543), .A(n9267), .ZN(P1_U3270) );
  XOR2_X1 U10558 ( .A(n9268), .B(n9270), .Z(n9548) );
  XOR2_X1 U10559 ( .A(n9270), .B(n9269), .Z(n9272) );
  OAI21_X1 U10560 ( .B1(n9272), .B2(n9828), .A(n9271), .ZN(n9544) );
  INV_X1 U10561 ( .A(n9273), .ZN(n9274) );
  AOI211_X1 U10562 ( .C1(n9546), .C2(n4576), .A(n9481), .B(n9274), .ZN(n9545)
         );
  NAND2_X1 U10563 ( .A1(n9545), .A2(n9892), .ZN(n9277) );
  AOI22_X1 U10564 ( .A1(n9896), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9275), .B2(
        n9847), .ZN(n9276) );
  OAI211_X1 U10565 ( .C1(n9278), .C2(n9883), .A(n9277), .B(n9276), .ZN(n9279)
         );
  AOI21_X1 U10566 ( .B1(n9544), .B2(n9671), .A(n9279), .ZN(n9280) );
  OAI21_X1 U10567 ( .B1(n9548), .B2(n9488), .A(n9280), .ZN(P1_U3271) );
  XOR2_X1 U10568 ( .A(n9283), .B(n9281), .Z(n9553) );
  AOI21_X1 U10569 ( .B1(n9284), .B2(n9283), .A(n9282), .ZN(n9287) );
  INV_X1 U10570 ( .A(n9285), .ZN(n9286) );
  OAI21_X1 U10571 ( .B1(n9287), .B2(n9828), .A(n9286), .ZN(n9549) );
  AOI211_X1 U10572 ( .C1(n9551), .C2(n9450), .A(n9481), .B(n9288), .ZN(n9550)
         );
  NAND2_X1 U10573 ( .A1(n9550), .A2(n9892), .ZN(n9292) );
  INV_X1 U10574 ( .A(n9289), .ZN(n9290) );
  AOI22_X1 U10575 ( .A1(n9290), .A2(n9847), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9896), .ZN(n9291) );
  OAI211_X1 U10576 ( .C1(n9293), .C2(n9883), .A(n9292), .B(n9291), .ZN(n9294)
         );
  AOI21_X1 U10577 ( .B1(n9549), .B2(n9671), .A(n9294), .ZN(n9295) );
  OAI21_X1 U10578 ( .B1(n9553), .B2(n9488), .A(n9295), .ZN(n9440) );
  AOI22_X1 U10579 ( .A1(n6252), .A2(keyinput33), .B1(n9241), .B2(keyinput27), 
        .ZN(n9296) );
  OAI221_X1 U10580 ( .B1(n6252), .B2(keyinput33), .C1(n9241), .C2(keyinput27), 
        .A(n9296), .ZN(n9307) );
  INV_X1 U10581 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n9898) );
  AOI22_X1 U10582 ( .A1(n9298), .A2(keyinput26), .B1(n9898), .B2(keyinput5), 
        .ZN(n9297) );
  OAI221_X1 U10583 ( .B1(n9298), .B2(keyinput26), .C1(n9898), .C2(keyinput5), 
        .A(n9297), .ZN(n9306) );
  AOI22_X1 U10584 ( .A1(n9300), .A2(keyinput20), .B1(n5854), .B2(keyinput19), 
        .ZN(n9299) );
  OAI221_X1 U10585 ( .B1(n9300), .B2(keyinput20), .C1(n5854), .C2(keyinput19), 
        .A(n9299), .ZN(n9305) );
  AOI22_X1 U10586 ( .A1(n9303), .A2(keyinput2), .B1(n9302), .B2(keyinput51), 
        .ZN(n9301) );
  OAI221_X1 U10587 ( .B1(n9303), .B2(keyinput2), .C1(n9302), .C2(keyinput51), 
        .A(n9301), .ZN(n9304) );
  NOR4_X1 U10588 ( .A1(n9307), .A2(n9306), .A3(n9305), .A4(n9304), .ZN(n9351)
         );
  AOI22_X1 U10589 ( .A1(n9310), .A2(keyinput55), .B1(keyinput1), .B2(n9309), 
        .ZN(n9308) );
  OAI221_X1 U10590 ( .B1(n9310), .B2(keyinput55), .C1(n9309), .C2(keyinput1), 
        .A(n9308), .ZN(n9314) );
  INV_X1 U10591 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9897) );
  AOI22_X1 U10592 ( .A1(n9897), .A2(keyinput22), .B1(keyinput60), .B2(n9312), 
        .ZN(n9311) );
  OAI221_X1 U10593 ( .B1(n9897), .B2(keyinput22), .C1(n9312), .C2(keyinput60), 
        .A(n9311), .ZN(n9313) );
  NOR2_X1 U10594 ( .A1(n9314), .A2(n9313), .ZN(n9350) );
  INV_X1 U10595 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9899) );
  AOI22_X1 U10596 ( .A1(n9899), .A2(keyinput15), .B1(keyinput58), .B2(n9316), 
        .ZN(n9315) );
  OAI221_X1 U10597 ( .B1(n9899), .B2(keyinput15), .C1(n9316), .C2(keyinput58), 
        .A(n9315), .ZN(n9326) );
  INV_X1 U10598 ( .A(keyinput61), .ZN(n9317) );
  XOR2_X1 U10599 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(n9317), .Z(n9321) );
  XNOR2_X1 U10600 ( .A(keyinput3), .B(P2_REG2_REG_18__SCAN_IN), .ZN(n9320) );
  XNOR2_X1 U10601 ( .A(P1_REG1_REG_30__SCAN_IN), .B(keyinput32), .ZN(n9319) );
  XNOR2_X1 U10602 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput21), .ZN(n9318) );
  NAND4_X1 U10603 ( .A1(n9321), .A2(n9320), .A3(n9319), .A4(n9318), .ZN(n9325)
         );
  AOI22_X1 U10604 ( .A1(n6892), .A2(keyinput34), .B1(n9323), .B2(keyinput11), 
        .ZN(n9322) );
  OAI221_X1 U10605 ( .B1(n6892), .B2(keyinput34), .C1(n9323), .C2(keyinput11), 
        .A(n9322), .ZN(n9324) );
  NOR3_X1 U10606 ( .A1(n9326), .A2(n9325), .A3(n9324), .ZN(n9349) );
  XNOR2_X1 U10607 ( .A(P2_IR_REG_23__SCAN_IN), .B(keyinput35), .ZN(n9330) );
  XNOR2_X1 U10608 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput36), .ZN(n9329) );
  XNOR2_X1 U10609 ( .A(P2_REG0_REG_31__SCAN_IN), .B(keyinput7), .ZN(n9328) );
  XNOR2_X1 U10610 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput44), .ZN(n9327) );
  NAND4_X1 U10611 ( .A1(n9330), .A2(n9329), .A3(n9328), .A4(n9327), .ZN(n9347)
         );
  XOR2_X1 U10612 ( .A(n8041), .B(keyinput57), .Z(n9335) );
  XOR2_X1 U10613 ( .A(n9331), .B(keyinput38), .Z(n9334) );
  INV_X1 U10614 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10091) );
  XOR2_X1 U10615 ( .A(n10091), .B(keyinput13), .Z(n9333) );
  XNOR2_X1 U10616 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput41), .ZN(n9332) );
  NAND4_X1 U10617 ( .A1(n9335), .A2(n9334), .A3(n9333), .A4(n9332), .ZN(n9346)
         );
  XNOR2_X1 U10618 ( .A(P2_REG2_REG_0__SCAN_IN), .B(keyinput39), .ZN(n9339) );
  XNOR2_X1 U10619 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput48), .ZN(n9338) );
  XNOR2_X1 U10620 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput49), .ZN(n9337)
         );
  XNOR2_X1 U10621 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput9), .ZN(n9336) );
  NAND4_X1 U10622 ( .A1(n9339), .A2(n9338), .A3(n9337), .A4(n9336), .ZN(n9345)
         );
  XNOR2_X1 U10623 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput28), .ZN(n9343) );
  XNOR2_X1 U10624 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput46), .ZN(n9342) );
  XNOR2_X1 U10625 ( .A(P2_REG0_REG_17__SCAN_IN), .B(keyinput50), .ZN(n9341) );
  XNOR2_X1 U10626 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput23), .ZN(n9340) );
  NAND4_X1 U10627 ( .A1(n9343), .A2(n9342), .A3(n9341), .A4(n9340), .ZN(n9344)
         );
  NOR4_X1 U10628 ( .A1(n9347), .A2(n9346), .A3(n9345), .A4(n9344), .ZN(n9348)
         );
  NAND4_X1 U10629 ( .A1(n9351), .A2(n9350), .A3(n9349), .A4(n9348), .ZN(n9425)
         );
  NOR3_X1 U10630 ( .A1(keyinput6), .A2(keyinput40), .A3(keyinput26), .ZN(n9357) );
  NAND2_X1 U10631 ( .A1(keyinput15), .A2(keyinput3), .ZN(n9352) );
  NOR3_X1 U10632 ( .A1(keyinput36), .A2(keyinput58), .A3(n9352), .ZN(n9356) );
  NAND3_X1 U10633 ( .A1(keyinput44), .A2(keyinput61), .A3(keyinput21), .ZN(
        n9354) );
  NAND3_X1 U10634 ( .A1(keyinput56), .A2(keyinput47), .A3(keyinput51), .ZN(
        n9353) );
  NOR4_X1 U10635 ( .A1(keyinput7), .A2(keyinput2), .A3(n9354), .A4(n9353), 
        .ZN(n9355) );
  NAND4_X1 U10636 ( .A1(keyinput5), .A2(n9357), .A3(n9356), .A4(n9355), .ZN(
        n9380) );
  NOR4_X1 U10637 ( .A1(keyinput13), .A2(keyinput28), .A3(keyinput29), .A4(
        keyinput42), .ZN(n9362) );
  NOR3_X1 U10638 ( .A1(keyinput12), .A2(keyinput24), .A3(keyinput41), .ZN(
        n9361) );
  NAND4_X1 U10639 ( .A1(keyinput49), .A2(keyinput9), .A3(keyinput23), .A4(
        keyinput46), .ZN(n9359) );
  NAND2_X1 U10640 ( .A1(keyinput16), .A2(keyinput33), .ZN(n9358) );
  NOR4_X1 U10641 ( .A1(keyinput27), .A2(keyinput59), .A3(n9359), .A4(n9358), 
        .ZN(n9360) );
  NAND4_X1 U10642 ( .A1(n9362), .A2(keyinput57), .A3(n9361), .A4(n9360), .ZN(
        n9379) );
  NOR3_X1 U10643 ( .A1(keyinput50), .A2(keyinput48), .A3(keyinput25), .ZN(
        n9365) );
  INV_X1 U10644 ( .A(keyinput14), .ZN(n9363) );
  NOR3_X1 U10645 ( .A1(keyinput54), .A2(keyinput62), .A3(n9363), .ZN(n9364) );
  AND4_X1 U10646 ( .A1(keyinput30), .A2(n9365), .A3(keyinput43), .A4(n9364), 
        .ZN(n9373) );
  NOR2_X1 U10647 ( .A1(keyinput45), .A2(keyinput17), .ZN(n9366) );
  NAND3_X1 U10648 ( .A1(keyinput52), .A2(keyinput63), .A3(n9366), .ZN(n9368)
         );
  NAND3_X1 U10649 ( .A1(keyinput31), .A2(keyinput22), .A3(keyinput60), .ZN(
        n9367) );
  NOR3_X1 U10650 ( .A1(n9368), .A2(n9367), .A3(keyinput18), .ZN(n9372) );
  NOR3_X1 U10651 ( .A1(keyinput0), .A2(keyinput38), .A3(keyinput35), .ZN(n9370) );
  NOR3_X1 U10652 ( .A1(keyinput32), .A2(keyinput4), .A3(keyinput8), .ZN(n9369)
         );
  AND4_X1 U10653 ( .A1(keyinput53), .A2(n9370), .A3(keyinput39), .A4(n9369), 
        .ZN(n9371) );
  NAND3_X1 U10654 ( .A1(n9373), .A2(n9372), .A3(n9371), .ZN(n9378) );
  NOR2_X1 U10655 ( .A1(keyinput55), .A2(keyinput20), .ZN(n9376) );
  NAND2_X1 U10656 ( .A1(keyinput37), .A2(keyinput34), .ZN(n9374) );
  NOR3_X1 U10657 ( .A1(keyinput11), .A2(keyinput10), .A3(n9374), .ZN(n9375) );
  NAND4_X1 U10658 ( .A1(keyinput1), .A2(keyinput19), .A3(n9376), .A4(n9375), 
        .ZN(n9377) );
  NOR4_X1 U10659 ( .A1(n9380), .A2(n9379), .A3(n9378), .A4(n9377), .ZN(n9424)
         );
  INV_X1 U10660 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9382) );
  AOI22_X1 U10661 ( .A1(n7507), .A2(keyinput30), .B1(keyinput25), .B2(n9382), 
        .ZN(n9381) );
  OAI221_X1 U10662 ( .B1(n7507), .B2(keyinput30), .C1(n9382), .C2(keyinput25), 
        .A(n9381), .ZN(n9391) );
  AOI22_X1 U10663 ( .A1(n9385), .A2(keyinput16), .B1(n9384), .B2(keyinput59), 
        .ZN(n9383) );
  OAI221_X1 U10664 ( .B1(n9385), .B2(keyinput16), .C1(n9384), .C2(keyinput59), 
        .A(n9383), .ZN(n9390) );
  AOI22_X1 U10665 ( .A1(n9388), .A2(keyinput56), .B1(n9387), .B2(keyinput47), 
        .ZN(n9386) );
  OAI221_X1 U10666 ( .B1(n9388), .B2(keyinput56), .C1(n9387), .C2(keyinput47), 
        .A(n9386), .ZN(n9389) );
  NOR3_X1 U10667 ( .A1(n9391), .A2(n9390), .A3(n9389), .ZN(n9422) );
  INV_X1 U10668 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9393) );
  AOI22_X1 U10669 ( .A1(n9393), .A2(keyinput31), .B1(keyinput18), .B2(n4948), 
        .ZN(n9392) );
  OAI221_X1 U10670 ( .B1(n9393), .B2(keyinput31), .C1(n4948), .C2(keyinput18), 
        .A(n9392), .ZN(n9402) );
  AOI22_X1 U10671 ( .A1(n9396), .A2(keyinput4), .B1(n9395), .B2(keyinput8), 
        .ZN(n9394) );
  OAI221_X1 U10672 ( .B1(n9396), .B2(keyinput4), .C1(n9395), .C2(keyinput8), 
        .A(n9394), .ZN(n9401) );
  AOI22_X1 U10673 ( .A1(n9399), .A2(keyinput53), .B1(n9398), .B2(keyinput0), 
        .ZN(n9397) );
  OAI221_X1 U10674 ( .B1(n9399), .B2(keyinput53), .C1(n9398), .C2(keyinput0), 
        .A(n9397), .ZN(n9400) );
  NOR3_X1 U10675 ( .A1(n9402), .A2(n9401), .A3(n9400), .ZN(n9421) );
  INV_X1 U10676 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9405) );
  INV_X1 U10677 ( .A(keyinput12), .ZN(n9404) );
  AOI22_X1 U10678 ( .A1(n9405), .A2(keyinput24), .B1(P2_ADDR_REG_17__SCAN_IN), 
        .B2(n9404), .ZN(n9403) );
  OAI221_X1 U10679 ( .B1(n9405), .B2(keyinput24), .C1(n9404), .C2(
        P2_ADDR_REG_17__SCAN_IN), .A(n9403), .ZN(n9410) );
  INV_X1 U10680 ( .A(keyinput42), .ZN(n9407) );
  AOI22_X1 U10681 ( .A1(n9408), .A2(keyinput29), .B1(P2_ADDR_REG_5__SCAN_IN), 
        .B2(n9407), .ZN(n9406) );
  OAI221_X1 U10682 ( .B1(n9408), .B2(keyinput29), .C1(n9407), .C2(
        P2_ADDR_REG_5__SCAN_IN), .A(n9406), .ZN(n9409) );
  NOR2_X1 U10683 ( .A1(n9410), .A2(n9409), .ZN(n9420) );
  INV_X1 U10684 ( .A(keyinput40), .ZN(n9412) );
  AOI22_X1 U10685 ( .A1(n9413), .A2(keyinput6), .B1(P1_ADDR_REG_17__SCAN_IN), 
        .B2(n9412), .ZN(n9411) );
  OAI221_X1 U10686 ( .B1(n9413), .B2(keyinput6), .C1(n9412), .C2(
        P1_ADDR_REG_17__SCAN_IN), .A(n9411), .ZN(n9418) );
  INV_X1 U10687 ( .A(keyinput37), .ZN(n9415) );
  AOI22_X1 U10688 ( .A1(n9416), .A2(keyinput10), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n9415), .ZN(n9414) );
  OAI221_X1 U10689 ( .B1(n9416), .B2(keyinput10), .C1(n9415), .C2(
        P1_ADDR_REG_15__SCAN_IN), .A(n9414), .ZN(n9417) );
  NOR2_X1 U10690 ( .A1(n9418), .A2(n9417), .ZN(n9419) );
  NAND4_X1 U10691 ( .A1(n9422), .A2(n9421), .A3(n9420), .A4(n9419), .ZN(n9423)
         );
  NOR3_X1 U10692 ( .A1(n9425), .A2(n9424), .A3(n9423), .ZN(n9438) );
  INV_X1 U10693 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9428) );
  INV_X1 U10694 ( .A(SI_28_), .ZN(n9427) );
  AOI22_X1 U10695 ( .A1(n9428), .A2(keyinput63), .B1(n9427), .B2(keyinput17), 
        .ZN(n9426) );
  OAI221_X1 U10696 ( .B1(n9428), .B2(keyinput63), .C1(n9427), .C2(keyinput17), 
        .A(n9426), .ZN(n9436) );
  AOI22_X1 U10697 ( .A1(n5740), .A2(keyinput52), .B1(n6033), .B2(keyinput45), 
        .ZN(n9429) );
  OAI221_X1 U10698 ( .B1(n5740), .B2(keyinput52), .C1(n6033), .C2(keyinput45), 
        .A(n9429), .ZN(n9435) );
  AOI22_X1 U10699 ( .A1(n9431), .A2(keyinput14), .B1(keyinput62), .B2(n7298), 
        .ZN(n9430) );
  OAI221_X1 U10700 ( .B1(n9431), .B2(keyinput14), .C1(n7298), .C2(keyinput62), 
        .A(n9430), .ZN(n9434) );
  AOI22_X1 U10701 ( .A1(n5588), .A2(keyinput43), .B1(n6141), .B2(keyinput54), 
        .ZN(n9432) );
  OAI221_X1 U10702 ( .B1(n5588), .B2(keyinput43), .C1(n6141), .C2(keyinput54), 
        .A(n9432), .ZN(n9433) );
  NOR4_X1 U10703 ( .A1(n9436), .A2(n9435), .A3(n9434), .A4(n9433), .ZN(n9437)
         );
  NAND2_X1 U10704 ( .A1(n9438), .A2(n9437), .ZN(n9439) );
  XNOR2_X1 U10705 ( .A(n9440), .B(n9439), .ZN(P1_U3272) );
  OAI21_X1 U10706 ( .B1(n9442), .B2(n9445), .A(n9441), .ZN(n9443) );
  INV_X1 U10707 ( .A(n9443), .ZN(n9558) );
  AOI21_X1 U10708 ( .B1(n9446), .B2(n9445), .A(n9444), .ZN(n9448) );
  OAI21_X1 U10709 ( .B1(n9448), .B2(n9828), .A(n9447), .ZN(n9554) );
  INV_X1 U10710 ( .A(n9450), .ZN(n9451) );
  AOI211_X1 U10711 ( .C1(n9556), .C2(n9459), .A(n9481), .B(n9451), .ZN(n9555)
         );
  NAND2_X1 U10712 ( .A1(n9555), .A2(n9892), .ZN(n9455) );
  INV_X1 U10713 ( .A(n9452), .ZN(n9453) );
  AOI22_X1 U10714 ( .A1(n9453), .A2(n9847), .B1(P1_REG2_REG_20__SCAN_IN), .B2(
        n9881), .ZN(n9454) );
  OAI211_X1 U10715 ( .C1(n9092), .C2(n9883), .A(n9455), .B(n9454), .ZN(n9456)
         );
  AOI21_X1 U10716 ( .B1(n9554), .B2(n9671), .A(n9456), .ZN(n9457) );
  OAI21_X1 U10717 ( .B1(n9558), .B2(n9488), .A(n9457), .ZN(P1_U3273) );
  XOR2_X1 U10718 ( .A(n9458), .B(n9465), .Z(n9563) );
  AOI21_X1 U10719 ( .B1(n9561), .B2(n9479), .A(n9481), .ZN(n9460) );
  AND2_X1 U10720 ( .A1(n9460), .A2(n9459), .ZN(n9560) );
  OAI22_X1 U10721 ( .A1(n9462), .A2(n9883), .B1(n9461), .B2(n9671), .ZN(n9463)
         );
  AOI21_X1 U10722 ( .B1(n9560), .B2(n9892), .A(n9463), .ZN(n9471) );
  XOR2_X1 U10723 ( .A(n9465), .B(n9464), .Z(n9467) );
  OAI21_X1 U10724 ( .B1(n9467), .B2(n9828), .A(n9466), .ZN(n9559) );
  NOR2_X1 U10725 ( .A1(n9468), .A2(n9879), .ZN(n9469) );
  OAI21_X1 U10726 ( .B1(n9559), .B2(n9469), .A(n9671), .ZN(n9470) );
  OAI211_X1 U10727 ( .C1(n9563), .C2(n9488), .A(n9471), .B(n9470), .ZN(
        P1_U3274) );
  XOR2_X1 U10728 ( .A(n9472), .B(n9475), .Z(n9568) );
  NOR2_X1 U10729 ( .A1(n9474), .A2(n4542), .ZN(n9476) );
  XNOR2_X1 U10730 ( .A(n9476), .B(n9475), .ZN(n9478) );
  OAI21_X1 U10731 ( .B1(n9478), .B2(n9828), .A(n9477), .ZN(n9564) );
  INV_X1 U10732 ( .A(n9479), .ZN(n9480) );
  AOI211_X1 U10733 ( .C1(n9566), .C2(n4399), .A(n9481), .B(n9480), .ZN(n9565)
         );
  NAND2_X1 U10734 ( .A1(n9565), .A2(n9892), .ZN(n9484) );
  AOI22_X1 U10735 ( .A1(n9896), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9482), .B2(
        n9847), .ZN(n9483) );
  OAI211_X1 U10736 ( .C1(n9485), .C2(n9883), .A(n9484), .B(n9483), .ZN(n9486)
         );
  AOI21_X1 U10737 ( .B1(n9671), .B2(n9564), .A(n9486), .ZN(n9487) );
  OAI21_X1 U10738 ( .B1(n9568), .B2(n9488), .A(n9487), .ZN(P1_U3275) );
  INV_X1 U10739 ( .A(n9494), .ZN(n9489) );
  XNOR2_X1 U10740 ( .A(n9490), .B(n9489), .ZN(n9492) );
  AOI21_X1 U10741 ( .B1(n9492), .B2(n9876), .A(n9491), .ZN(n9677) );
  OAI21_X1 U10742 ( .B1(n9495), .B2(n9494), .A(n9493), .ZN(n9679) );
  NAND2_X1 U10743 ( .A1(n9679), .A2(n9893), .ZN(n9504) );
  OAI22_X1 U10744 ( .A1(n9671), .A2(n9497), .B1(n9496), .B2(n9879), .ZN(n9501)
         );
  INV_X1 U10745 ( .A(n9657), .ZN(n9498) );
  OAI211_X1 U10746 ( .C1(n4580), .C2(n9498), .A(n4399), .B(n9888), .ZN(n9676)
         );
  NOR2_X1 U10747 ( .A1(n9676), .A2(n9499), .ZN(n9500) );
  AOI211_X1 U10748 ( .C1(n9835), .C2(n9502), .A(n9501), .B(n9500), .ZN(n9503)
         );
  OAI211_X1 U10749 ( .C1(n9881), .C2(n9677), .A(n9504), .B(n9503), .ZN(
        P1_U3276) );
  OAI211_X1 U10750 ( .C1(n9094), .C2(n9983), .A(n9505), .B(n9506), .ZN(n9570)
         );
  MUX2_X1 U10751 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9570), .S(n9569), .Z(
        P1_U3553) );
  OAI211_X1 U10752 ( .C1(n9508), .C2(n9983), .A(n9507), .B(n9506), .ZN(n9571)
         );
  MUX2_X1 U10753 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9571), .S(n10008), .Z(
        P1_U3552) );
  AOI21_X1 U10754 ( .B1(n9933), .B2(n9515), .A(n9514), .ZN(n9516) );
  OAI211_X1 U10755 ( .C1(n9518), .C2(n9937), .A(n9517), .B(n9516), .ZN(n9572)
         );
  MUX2_X1 U10756 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9572), .S(n10008), .Z(
        P1_U3550) );
  OAI21_X1 U10757 ( .B1(n9523), .B2(n9937), .A(n9522), .ZN(n9573) );
  MUX2_X1 U10758 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9573), .S(n9569), .Z(
        P1_U3549) );
  AOI21_X1 U10759 ( .B1(n9933), .B2(n9525), .A(n9524), .ZN(n9526) );
  OAI211_X1 U10760 ( .C1(n9528), .C2(n9937), .A(n9527), .B(n9526), .ZN(n9574)
         );
  MUX2_X1 U10761 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9574), .S(n9569), .Z(
        P1_U3548) );
  AOI21_X1 U10762 ( .B1(n9933), .B2(n9530), .A(n9529), .ZN(n9531) );
  OAI211_X1 U10763 ( .C1(n9533), .C2(n9937), .A(n9532), .B(n9531), .ZN(n9575)
         );
  MUX2_X1 U10764 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9575), .S(n9569), .Z(
        P1_U3547) );
  AOI211_X1 U10765 ( .C1(n9933), .C2(n9536), .A(n9535), .B(n9534), .ZN(n9537)
         );
  OAI21_X1 U10766 ( .B1(n9538), .B2(n9937), .A(n9537), .ZN(n9576) );
  MUX2_X1 U10767 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9576), .S(n9569), .Z(
        P1_U3546) );
  AOI22_X1 U10768 ( .A1(n9540), .A2(n9888), .B1(n9933), .B2(n9539), .ZN(n9541)
         );
  OAI211_X1 U10769 ( .C1(n9543), .C2(n9937), .A(n9542), .B(n9541), .ZN(n9577)
         );
  MUX2_X1 U10770 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9577), .S(n9569), .Z(
        P1_U3545) );
  AOI211_X1 U10771 ( .C1(n9933), .C2(n9546), .A(n9545), .B(n9544), .ZN(n9547)
         );
  OAI21_X1 U10772 ( .B1(n9548), .B2(n9937), .A(n9547), .ZN(n9578) );
  MUX2_X1 U10773 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9578), .S(n9569), .Z(
        P1_U3544) );
  AOI211_X1 U10774 ( .C1(n9933), .C2(n9551), .A(n9550), .B(n9549), .ZN(n9552)
         );
  OAI21_X1 U10775 ( .B1(n9553), .B2(n9937), .A(n9552), .ZN(n9579) );
  MUX2_X1 U10776 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9579), .S(n9569), .Z(
        P1_U3543) );
  AOI211_X1 U10777 ( .C1(n9933), .C2(n9556), .A(n9555), .B(n9554), .ZN(n9557)
         );
  OAI21_X1 U10778 ( .B1(n9558), .B2(n9937), .A(n9557), .ZN(n9580) );
  MUX2_X1 U10779 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9580), .S(n9569), .Z(
        P1_U3542) );
  AOI211_X1 U10780 ( .C1(n9933), .C2(n9561), .A(n9560), .B(n9559), .ZN(n9562)
         );
  OAI21_X1 U10781 ( .B1(n9563), .B2(n9937), .A(n9562), .ZN(n9581) );
  MUX2_X1 U10782 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9581), .S(n9569), .Z(
        P1_U3541) );
  AOI211_X1 U10783 ( .C1(n9933), .C2(n9566), .A(n9565), .B(n9564), .ZN(n9567)
         );
  OAI21_X1 U10784 ( .B1(n9568), .B2(n9937), .A(n9567), .ZN(n9582) );
  MUX2_X1 U10785 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9582), .S(n9569), .Z(
        P1_U3540) );
  MUX2_X1 U10786 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9570), .S(n9991), .Z(
        P1_U3521) );
  MUX2_X1 U10787 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9571), .S(n9991), .Z(
        P1_U3520) );
  MUX2_X1 U10788 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9572), .S(n9991), .Z(
        P1_U3518) );
  MUX2_X1 U10789 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9573), .S(n9991), .Z(
        P1_U3517) );
  MUX2_X1 U10790 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9574), .S(n9991), .Z(
        P1_U3516) );
  MUX2_X1 U10791 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9575), .S(n9991), .Z(
        P1_U3515) );
  MUX2_X1 U10792 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9576), .S(n9991), .Z(
        P1_U3514) );
  MUX2_X1 U10793 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9577), .S(n9991), .Z(
        P1_U3513) );
  MUX2_X1 U10794 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9578), .S(n9991), .Z(
        P1_U3512) );
  MUX2_X1 U10795 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9579), .S(n9991), .Z(
        P1_U3511) );
  MUX2_X1 U10796 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9580), .S(n9991), .Z(
        P1_U3510) );
  MUX2_X1 U10797 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9581), .S(n9991), .Z(
        P1_U3509) );
  MUX2_X1 U10798 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9582), .S(n9991), .Z(
        P1_U3507) );
  MUX2_X1 U10799 ( .A(n9583), .B(P1_D_REG_1__SCAN_IN), .S(n9901), .Z(P1_U3440)
         );
  MUX2_X1 U10800 ( .A(n9584), .B(P1_D_REG_0__SCAN_IN), .S(n9901), .Z(P1_U3439)
         );
  NOR4_X1 U10801 ( .A1(n9586), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5892), .A4(
        P1_U3086), .ZN(n9587) );
  AOI21_X1 U10802 ( .B1(n9588), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9587), .ZN(
        n9589) );
  OAI21_X1 U10803 ( .B1(n9591), .B2(n9590), .A(n9589), .ZN(P1_U3324) );
  INV_X1 U10804 ( .A(n9592), .ZN(n9593) );
  MUX2_X1 U10805 ( .A(n9593), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI211_X1 U10806 ( .C1(n9596), .C2(n9595), .A(n9594), .B(n9790), .ZN(n9601)
         );
  AOI211_X1 U10807 ( .C1(n9599), .C2(n9598), .A(n9597), .B(n9795), .ZN(n9600)
         );
  AOI211_X1 U10808 ( .C1(n9801), .C2(n9602), .A(n9601), .B(n9600), .ZN(n9604)
         );
  OAI211_X1 U10809 ( .C1(n9805), .C2(n9605), .A(n9604), .B(n9603), .ZN(
        P1_U3253) );
  AOI21_X1 U10810 ( .B1(n9608), .B2(n9607), .A(n9606), .ZN(n9609) );
  NAND2_X1 U10811 ( .A1(n9763), .A2(n9609), .ZN(n9617) );
  INV_X1 U10812 ( .A(n9610), .ZN(n9614) );
  NAND2_X1 U10813 ( .A1(n9612), .A2(n9611), .ZN(n9613) );
  NAND2_X1 U10814 ( .A1(n9614), .A2(n9613), .ZN(n9615) );
  OR2_X1 U10815 ( .A1(n9795), .A2(n9615), .ZN(n9616) );
  OAI211_X1 U10816 ( .C1(n9773), .C2(n9618), .A(n9617), .B(n9616), .ZN(n9619)
         );
  INV_X1 U10817 ( .A(n9619), .ZN(n9621) );
  NAND2_X1 U10818 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9620) );
  OAI211_X1 U10819 ( .C1(n9805), .C2(n9622), .A(n9621), .B(n9620), .ZN(
        P1_U3250) );
  AOI21_X1 U10820 ( .B1(n9625), .B2(n9624), .A(n9623), .ZN(n9626) );
  NAND2_X1 U10821 ( .A1(n9763), .A2(n9626), .ZN(n9634) );
  NAND2_X1 U10822 ( .A1(n9628), .A2(n9627), .ZN(n9631) );
  INV_X1 U10823 ( .A(n9629), .ZN(n9630) );
  NAND2_X1 U10824 ( .A1(n9631), .A2(n9630), .ZN(n9632) );
  OR2_X1 U10825 ( .A1(n9795), .A2(n9632), .ZN(n9633) );
  OAI211_X1 U10826 ( .C1(n9773), .C2(n9635), .A(n9634), .B(n9633), .ZN(n9636)
         );
  INV_X1 U10827 ( .A(n9636), .ZN(n9638) );
  NAND2_X1 U10828 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9637) );
  OAI211_X1 U10829 ( .C1(n9805), .C2(n9639), .A(n9638), .B(n9637), .ZN(
        P1_U3251) );
  NOR2_X1 U10830 ( .A1(n9640), .A2(n10079), .ZN(n9642) );
  AOI211_X1 U10831 ( .C1(n9643), .C2(n10049), .A(n9642), .B(n9641), .ZN(n9651)
         );
  AOI22_X1 U10832 ( .A1(n10103), .A2(n9651), .B1(n9644), .B2(n10100), .ZN(
        P2_U3473) );
  AND2_X1 U10833 ( .A1(n9645), .A2(n10049), .ZN(n9648) );
  AND2_X1 U10834 ( .A1(n9646), .A2(n10066), .ZN(n9647) );
  NOR3_X1 U10835 ( .A1(n9649), .A2(n9648), .A3(n9647), .ZN(n9653) );
  AOI22_X1 U10836 ( .A1(n10103), .A2(n9653), .B1(n9650), .B2(n10100), .ZN(
        P2_U3472) );
  INV_X1 U10837 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9652) );
  AOI22_X1 U10838 ( .A1(n10087), .A2(n9652), .B1(n9651), .B2(n10085), .ZN(
        P2_U3432) );
  INV_X1 U10839 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9654) );
  AOI22_X1 U10840 ( .A1(n10087), .A2(n9654), .B1(n9653), .B2(n10085), .ZN(
        P2_U3429) );
  NAND2_X1 U10841 ( .A1(n9655), .A2(n9668), .ZN(n9656) );
  NAND3_X1 U10842 ( .A1(n9657), .A2(n9888), .A3(n9656), .ZN(n9682) );
  INV_X1 U10843 ( .A(n9682), .ZN(n9658) );
  AOI22_X1 U10844 ( .A1(n9658), .A2(n9892), .B1(P1_REG2_REG_16__SCAN_IN), .B2(
        n9881), .ZN(n9674) );
  XNOR2_X1 U10845 ( .A(n9659), .B(n9662), .ZN(n9680) );
  NAND3_X1 U10846 ( .A1(n9662), .A2(n9661), .A3(n9660), .ZN(n9663) );
  NAND2_X1 U10847 ( .A1(n9664), .A2(n9663), .ZN(n9666) );
  AOI21_X1 U10848 ( .B1(n9666), .B2(n9876), .A(n9665), .ZN(n9681) );
  NAND2_X1 U10849 ( .A1(n9668), .A2(n9667), .ZN(n9669) );
  OAI211_X1 U10850 ( .C1(n9680), .C2(n9670), .A(n9681), .B(n9669), .ZN(n9672)
         );
  NAND2_X1 U10851 ( .A1(n9672), .A2(n9671), .ZN(n9673) );
  OAI211_X1 U10852 ( .C1(n9675), .C2(n9879), .A(n9674), .B(n9673), .ZN(
        P1_U3277) );
  OAI211_X1 U10853 ( .C1(n4580), .C2(n9983), .A(n9677), .B(n9676), .ZN(n9678)
         );
  AOI21_X1 U10854 ( .B1(n9679), .B2(n9979), .A(n9678), .ZN(n9692) );
  AOI22_X1 U10855 ( .A1(n10008), .A2(n9692), .B1(n9060), .B2(n10006), .ZN(
        P1_U3539) );
  INV_X1 U10856 ( .A(n9680), .ZN(n9686) );
  INV_X1 U10857 ( .A(n9681), .ZN(n9685) );
  OAI21_X1 U10858 ( .B1(n9683), .B2(n9983), .A(n9682), .ZN(n9684) );
  AOI211_X1 U10859 ( .C1(n9686), .C2(n9979), .A(n9685), .B(n9684), .ZN(n9693)
         );
  AOI22_X1 U10860 ( .A1(n10008), .A2(n9693), .B1(n6034), .B2(n10006), .ZN(
        P1_U3538) );
  OAI211_X1 U10861 ( .C1(n9689), .C2(n9983), .A(n9688), .B(n9687), .ZN(n9690)
         );
  AOI21_X1 U10862 ( .B1(n9691), .B2(n9979), .A(n9690), .ZN(n9695) );
  AOI22_X1 U10863 ( .A1(n10008), .A2(n9695), .B1(n6014), .B2(n10006), .ZN(
        P1_U3537) );
  AOI22_X1 U10864 ( .A1(n9991), .A2(n9692), .B1(n6053), .B2(n9990), .ZN(
        P1_U3504) );
  AOI22_X1 U10865 ( .A1(n9991), .A2(n9693), .B1(n6033), .B2(n9990), .ZN(
        P1_U3501) );
  INV_X1 U10866 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9694) );
  AOI22_X1 U10867 ( .A1(n9991), .A2(n9695), .B1(n9694), .B2(n9990), .ZN(
        P1_U3498) );
  XNOR2_X1 U10868 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10869 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OAI211_X1 U10870 ( .C1(n9698), .C2(n9697), .A(n9763), .B(n9696), .ZN(n9705)
         );
  NOR2_X1 U10871 ( .A1(n9700), .A2(n9699), .ZN(n9701) );
  OR2_X1 U10872 ( .A1(n9702), .A2(n9701), .ZN(n9703) );
  OR2_X1 U10873 ( .A1(n9795), .A2(n9703), .ZN(n9704) );
  OAI211_X1 U10874 ( .C1(n9773), .C2(n9706), .A(n9705), .B(n9704), .ZN(n9707)
         );
  INV_X1 U10875 ( .A(n9707), .ZN(n9709) );
  NAND2_X1 U10876 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9708) );
  OAI211_X1 U10877 ( .C1(n9805), .C2(n9710), .A(n9709), .B(n9708), .ZN(
        P1_U3248) );
  AOI21_X1 U10878 ( .B1(n9713), .B2(n9712), .A(n9711), .ZN(n9714) );
  NAND2_X1 U10879 ( .A1(n9763), .A2(n9714), .ZN(n9722) );
  NAND2_X1 U10880 ( .A1(n9716), .A2(n9715), .ZN(n9719) );
  INV_X1 U10881 ( .A(n9717), .ZN(n9718) );
  NAND2_X1 U10882 ( .A1(n9719), .A2(n9718), .ZN(n9720) );
  OR2_X1 U10883 ( .A1(n9795), .A2(n9720), .ZN(n9721) );
  OAI211_X1 U10884 ( .C1(n9773), .C2(n9723), .A(n9722), .B(n9721), .ZN(n9724)
         );
  INV_X1 U10885 ( .A(n9724), .ZN(n9726) );
  OAI211_X1 U10886 ( .C1(n9805), .C2(n9727), .A(n9726), .B(n9725), .ZN(
        P1_U3249) );
  INV_X1 U10887 ( .A(n9728), .ZN(n9741) );
  AOI21_X1 U10888 ( .B1(n9731), .B2(n9730), .A(n9729), .ZN(n9732) );
  NAND2_X1 U10889 ( .A1(n9763), .A2(n9732), .ZN(n9740) );
  NAND2_X1 U10890 ( .A1(n9734), .A2(n9733), .ZN(n9737) );
  INV_X1 U10891 ( .A(n9735), .ZN(n9736) );
  NAND2_X1 U10892 ( .A1(n9737), .A2(n9736), .ZN(n9738) );
  OR2_X1 U10893 ( .A1(n9795), .A2(n9738), .ZN(n9739) );
  OAI211_X1 U10894 ( .C1(n9773), .C2(n9741), .A(n9740), .B(n9739), .ZN(n9742)
         );
  INV_X1 U10895 ( .A(n9742), .ZN(n9744) );
  OAI211_X1 U10896 ( .C1(n9805), .C2(n9745), .A(n9744), .B(n9743), .ZN(
        P1_U3254) );
  AOI211_X1 U10897 ( .C1(n9748), .C2(n9747), .A(n9746), .B(n9790), .ZN(n9753)
         );
  AOI211_X1 U10898 ( .C1(n9751), .C2(n9750), .A(n9749), .B(n9795), .ZN(n9752)
         );
  AOI211_X1 U10899 ( .C1(n9801), .C2(n9754), .A(n9753), .B(n9752), .ZN(n9756)
         );
  OAI211_X1 U10900 ( .C1(n9805), .C2(n9757), .A(n9756), .B(n9755), .ZN(
        P1_U3256) );
  INV_X1 U10901 ( .A(n9758), .ZN(n9772) );
  AOI21_X1 U10902 ( .B1(n9761), .B2(n9760), .A(n9759), .ZN(n9762) );
  NAND2_X1 U10903 ( .A1(n9763), .A2(n9762), .ZN(n9771) );
  NAND2_X1 U10904 ( .A1(n9765), .A2(n9764), .ZN(n9768) );
  INV_X1 U10905 ( .A(n9766), .ZN(n9767) );
  NAND2_X1 U10906 ( .A1(n9768), .A2(n9767), .ZN(n9769) );
  OR2_X1 U10907 ( .A1(n9795), .A2(n9769), .ZN(n9770) );
  OAI211_X1 U10908 ( .C1(n9773), .C2(n9772), .A(n9771), .B(n9770), .ZN(n9774)
         );
  INV_X1 U10909 ( .A(n9774), .ZN(n9776) );
  OAI211_X1 U10910 ( .C1(n9805), .C2(n9777), .A(n9776), .B(n9775), .ZN(
        P1_U3257) );
  AOI211_X1 U10911 ( .C1(n9779), .C2(n6014), .A(n9778), .B(n9790), .ZN(n9783)
         );
  AOI211_X1 U10912 ( .C1(n9781), .C2(n7787), .A(n9780), .B(n9795), .ZN(n9782)
         );
  AOI211_X1 U10913 ( .C1(n9801), .C2(n9784), .A(n9783), .B(n9782), .ZN(n9786)
         );
  OAI211_X1 U10914 ( .C1(n9787), .C2(n9805), .A(n9786), .B(n9785), .ZN(
        P1_U3258) );
  INV_X1 U10915 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9804) );
  INV_X1 U10916 ( .A(n9788), .ZN(n9789) );
  AOI211_X1 U10917 ( .C1(n9792), .C2(n9791), .A(n9790), .B(n9789), .ZN(n9799)
         );
  INV_X1 U10918 ( .A(n9793), .ZN(n9794) );
  AOI211_X1 U10919 ( .C1(n9797), .C2(n9796), .A(n9795), .B(n9794), .ZN(n9798)
         );
  AOI211_X1 U10920 ( .C1(n9801), .C2(n9800), .A(n9799), .B(n9798), .ZN(n9803)
         );
  NAND2_X1 U10921 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9802) );
  OAI211_X1 U10922 ( .C1(n9805), .C2(n9804), .A(n9803), .B(n9802), .ZN(
        P1_U3261) );
  XNOR2_X1 U10923 ( .A(n9806), .B(n9808), .ZN(n9988) );
  INV_X1 U10924 ( .A(n9807), .ZN(n9812) );
  AOI21_X1 U10925 ( .B1(n9810), .B2(n9809), .A(n9808), .ZN(n9811) );
  NOR3_X1 U10926 ( .A1(n9812), .A2(n9811), .A3(n9828), .ZN(n9814) );
  AOI211_X1 U10927 ( .C1(n9988), .C2(n9833), .A(n9814), .B(n9813), .ZN(n9985)
         );
  INV_X1 U10928 ( .A(n9815), .ZN(n9816) );
  AOI222_X1 U10929 ( .A1(n9817), .A2(n9835), .B1(P1_REG2_REG_14__SCAN_IN), 
        .B2(n9896), .C1(n9847), .C2(n9816), .ZN(n9823) );
  INV_X1 U10930 ( .A(n9818), .ZN(n9819) );
  OAI211_X1 U10931 ( .C1(n9984), .C2(n9820), .A(n9819), .B(n9888), .ZN(n9982)
         );
  INV_X1 U10932 ( .A(n9982), .ZN(n9821) );
  AOI22_X1 U10933 ( .A1(n9988), .A2(n9840), .B1(n9892), .B2(n9821), .ZN(n9822)
         );
  OAI211_X1 U10934 ( .C1(n9896), .C2(n9985), .A(n9823), .B(n9822), .ZN(
        P1_U3279) );
  XNOR2_X1 U10935 ( .A(n9824), .B(n9830), .ZN(n9950) );
  INV_X1 U10936 ( .A(n9825), .ZN(n9832) );
  INV_X1 U10937 ( .A(n9826), .ZN(n9827) );
  AOI211_X1 U10938 ( .C1(n9830), .C2(n9829), .A(n9828), .B(n9827), .ZN(n9831)
         );
  AOI211_X1 U10939 ( .C1(n9833), .C2(n9950), .A(n9832), .B(n9831), .ZN(n9947)
         );
  AOI222_X1 U10940 ( .A1(n9836), .A2(n9835), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n9896), .C1(n9847), .C2(n9834), .ZN(n9842) );
  OAI211_X1 U10941 ( .C1(n9946), .C2(n9838), .A(n9837), .B(n9888), .ZN(n9945)
         );
  INV_X1 U10942 ( .A(n9945), .ZN(n9839) );
  AOI22_X1 U10943 ( .A1(n9950), .A2(n9840), .B1(n9892), .B2(n9839), .ZN(n9841)
         );
  OAI211_X1 U10944 ( .C1(n9896), .C2(n9947), .A(n9842), .B(n9841), .ZN(
        P1_U3285) );
  XNOR2_X1 U10945 ( .A(n9843), .B(n9852), .ZN(n9846) );
  INV_X1 U10946 ( .A(n9844), .ZN(n9845) );
  AOI21_X1 U10947 ( .B1(n9846), .B2(n9876), .A(n9845), .ZN(n9941) );
  AOI22_X1 U10948 ( .A1(n9881), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n9848), .B2(
        n9847), .ZN(n9849) );
  OAI21_X1 U10949 ( .B1(n9883), .B2(n9940), .A(n9849), .ZN(n9850) );
  INV_X1 U10950 ( .A(n9850), .ZN(n9858) );
  XNOR2_X1 U10951 ( .A(n4301), .B(n9852), .ZN(n9944) );
  INV_X1 U10952 ( .A(n9853), .ZN(n9855) );
  OAI211_X1 U10953 ( .C1(n9940), .C2(n9855), .A(n9854), .B(n9888), .ZN(n9939)
         );
  INV_X1 U10954 ( .A(n9939), .ZN(n9856) );
  AOI22_X1 U10955 ( .A1(n9944), .A2(n9893), .B1(n9892), .B2(n9856), .ZN(n9857)
         );
  OAI211_X1 U10956 ( .C1(n9896), .C2(n9941), .A(n9858), .B(n9857), .ZN(
        P1_U3287) );
  XNOR2_X1 U10957 ( .A(n9859), .B(n9860), .ZN(n9862) );
  AOI21_X1 U10958 ( .B1(n9862), .B2(n9876), .A(n9861), .ZN(n9926) );
  NOR2_X1 U10959 ( .A1(n9879), .A2(n9863), .ZN(n9864) );
  AOI21_X1 U10960 ( .B1(n9881), .B2(P1_REG2_REG_4__SCAN_IN), .A(n9864), .ZN(
        n9865) );
  OAI21_X1 U10961 ( .B1(n9883), .B2(n9925), .A(n9865), .ZN(n9866) );
  INV_X1 U10962 ( .A(n9866), .ZN(n9873) );
  XNOR2_X1 U10963 ( .A(n9867), .B(n9868), .ZN(n9929) );
  OAI211_X1 U10964 ( .C1(n9870), .C2(n9925), .A(n9888), .B(n9869), .ZN(n9924)
         );
  INV_X1 U10965 ( .A(n9924), .ZN(n9871) );
  AOI22_X1 U10966 ( .A1(n9929), .A2(n9893), .B1(n9892), .B2(n9871), .ZN(n9872)
         );
  OAI211_X1 U10967 ( .C1(n9896), .C2(n9926), .A(n9873), .B(n9872), .ZN(
        P1_U3289) );
  XNOR2_X1 U10968 ( .A(n9874), .B(n9886), .ZN(n9877) );
  AOI21_X1 U10969 ( .B1(n9877), .B2(n9876), .A(n9875), .ZN(n9914) );
  NOR2_X1 U10970 ( .A1(n9879), .A2(n9878), .ZN(n9880) );
  AOI21_X1 U10971 ( .B1(n9881), .B2(P1_REG2_REG_2__SCAN_IN), .A(n9880), .ZN(
        n9882) );
  OAI21_X1 U10972 ( .B1(n9883), .B2(n9913), .A(n9882), .ZN(n9884) );
  INV_X1 U10973 ( .A(n9884), .ZN(n9895) );
  XNOR2_X1 U10974 ( .A(n9885), .B(n9886), .ZN(n9917) );
  INV_X1 U10975 ( .A(n9887), .ZN(n9890) );
  OAI211_X1 U10976 ( .C1(n9913), .C2(n9890), .A(n9889), .B(n9888), .ZN(n9912)
         );
  INV_X1 U10977 ( .A(n9912), .ZN(n9891) );
  AOI22_X1 U10978 ( .A1(n9917), .A2(n9893), .B1(n9892), .B2(n9891), .ZN(n9894)
         );
  OAI211_X1 U10979 ( .C1(n9896), .C2(n9914), .A(n9895), .B(n9894), .ZN(
        P1_U3291) );
  AND2_X1 U10980 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9901), .ZN(P1_U3294) );
  AND2_X1 U10981 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9901), .ZN(P1_U3295) );
  AND2_X1 U10982 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9901), .ZN(P1_U3296) );
  AND2_X1 U10983 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9901), .ZN(P1_U3297) );
  AND2_X1 U10984 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9901), .ZN(P1_U3298) );
  AND2_X1 U10985 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9901), .ZN(P1_U3299) );
  AND2_X1 U10986 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9901), .ZN(P1_U3300) );
  AND2_X1 U10987 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9901), .ZN(P1_U3301) );
  AND2_X1 U10988 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9901), .ZN(P1_U3302) );
  AND2_X1 U10989 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9901), .ZN(P1_U3303) );
  AND2_X1 U10990 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9901), .ZN(P1_U3304) );
  AND2_X1 U10991 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9901), .ZN(P1_U3305) );
  AND2_X1 U10992 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9901), .ZN(P1_U3306) );
  AND2_X1 U10993 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9901), .ZN(P1_U3307) );
  AND2_X1 U10994 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9901), .ZN(P1_U3308) );
  AND2_X1 U10995 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9901), .ZN(P1_U3309) );
  AND2_X1 U10996 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9901), .ZN(P1_U3310) );
  AND2_X1 U10997 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9901), .ZN(P1_U3311) );
  INV_X1 U10998 ( .A(n9901), .ZN(n9900) );
  NOR2_X1 U10999 ( .A1(n9900), .A2(n9897), .ZN(P1_U3312) );
  AND2_X1 U11000 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9901), .ZN(P1_U3313) );
  AND2_X1 U11001 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9901), .ZN(P1_U3314) );
  AND2_X1 U11002 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9901), .ZN(P1_U3315) );
  AND2_X1 U11003 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9901), .ZN(P1_U3316) );
  AND2_X1 U11004 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9901), .ZN(P1_U3317) );
  NOR2_X1 U11005 ( .A1(n9900), .A2(n9898), .ZN(P1_U3318) );
  AND2_X1 U11006 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9901), .ZN(P1_U3319) );
  AND2_X1 U11007 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9901), .ZN(P1_U3320) );
  AND2_X1 U11008 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9901), .ZN(P1_U3321) );
  NOR2_X1 U11009 ( .A1(n9900), .A2(n9899), .ZN(P1_U3322) );
  AND2_X1 U11010 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9901), .ZN(P1_U3323) );
  INV_X1 U11011 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9902) );
  AOI22_X1 U11012 ( .A1(n9991), .A2(n9903), .B1(n9902), .B2(n9990), .ZN(
        P1_U3453) );
  INV_X1 U11013 ( .A(n9904), .ZN(n9989) );
  INV_X1 U11014 ( .A(n9905), .ZN(n9910) );
  OAI21_X1 U11015 ( .B1(n9907), .B2(n9983), .A(n9906), .ZN(n9909) );
  AOI211_X1 U11016 ( .C1(n9989), .C2(n9910), .A(n9909), .B(n9908), .ZN(n9992)
         );
  INV_X1 U11017 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9911) );
  AOI22_X1 U11018 ( .A1(n9991), .A2(n9992), .B1(n9911), .B2(n9990), .ZN(
        P1_U3456) );
  OAI21_X1 U11019 ( .B1(n9913), .B2(n9983), .A(n9912), .ZN(n9916) );
  INV_X1 U11020 ( .A(n9914), .ZN(n9915) );
  AOI211_X1 U11021 ( .C1(n9917), .C2(n9979), .A(n9916), .B(n9915), .ZN(n9993)
         );
  AOI22_X1 U11022 ( .A1(n9991), .A2(n9993), .B1(n5719), .B2(n9990), .ZN(
        P1_U3459) );
  AOI21_X1 U11023 ( .B1(n9933), .B2(n4271), .A(n9918), .ZN(n9921) );
  OAI211_X1 U11024 ( .C1(n9937), .C2(n9922), .A(n9921), .B(n9920), .ZN(n9923)
         );
  INV_X1 U11025 ( .A(n9923), .ZN(n9994) );
  AOI22_X1 U11026 ( .A1(n9991), .A2(n9994), .B1(n5739), .B2(n9990), .ZN(
        P1_U3462) );
  OAI21_X1 U11027 ( .B1(n9925), .B2(n9983), .A(n9924), .ZN(n9928) );
  INV_X1 U11028 ( .A(n9926), .ZN(n9927) );
  AOI211_X1 U11029 ( .C1(n9979), .C2(n9929), .A(n9928), .B(n9927), .ZN(n9995)
         );
  INV_X1 U11030 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9930) );
  AOI22_X1 U11031 ( .A1(n9991), .A2(n9995), .B1(n9930), .B2(n9990), .ZN(
        P1_U3465) );
  AOI21_X1 U11032 ( .B1(n9933), .B2(n9932), .A(n9931), .ZN(n9934) );
  OAI211_X1 U11033 ( .C1(n9937), .C2(n9936), .A(n9935), .B(n9934), .ZN(n9938)
         );
  INV_X1 U11034 ( .A(n9938), .ZN(n9997) );
  AOI22_X1 U11035 ( .A1(n9991), .A2(n9997), .B1(n5784), .B2(n9990), .ZN(
        P1_U3468) );
  OAI21_X1 U11036 ( .B1(n9940), .B2(n9983), .A(n9939), .ZN(n9943) );
  INV_X1 U11037 ( .A(n9941), .ZN(n9942) );
  AOI211_X1 U11038 ( .C1(n9979), .C2(n9944), .A(n9943), .B(n9942), .ZN(n9999)
         );
  AOI22_X1 U11039 ( .A1(n9991), .A2(n9999), .B1(n5811), .B2(n9990), .ZN(
        P1_U3471) );
  OAI21_X1 U11040 ( .B1(n9946), .B2(n9983), .A(n9945), .ZN(n9949) );
  INV_X1 U11041 ( .A(n9947), .ZN(n9948) );
  AOI211_X1 U11042 ( .C1(n9989), .C2(n9950), .A(n9949), .B(n9948), .ZN(n10000)
         );
  AOI22_X1 U11043 ( .A1(n9991), .A2(n10000), .B1(n5854), .B2(n9990), .ZN(
        P1_U3477) );
  OAI21_X1 U11044 ( .B1(n9952), .B2(n9983), .A(n9951), .ZN(n9954) );
  AOI211_X1 U11045 ( .C1(n9979), .C2(n9955), .A(n9954), .B(n9953), .ZN(n10001)
         );
  INV_X1 U11046 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9956) );
  AOI22_X1 U11047 ( .A1(n9991), .A2(n10001), .B1(n9956), .B2(n9990), .ZN(
        P1_U3480) );
  OAI211_X1 U11048 ( .C1(n9959), .C2(n9983), .A(n9958), .B(n9957), .ZN(n9960)
         );
  AOI21_X1 U11049 ( .B1(n9961), .B2(n9979), .A(n9960), .ZN(n10002) );
  INV_X1 U11050 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9962) );
  AOI22_X1 U11051 ( .A1(n9991), .A2(n10002), .B1(n9962), .B2(n9990), .ZN(
        P1_U3483) );
  OAI21_X1 U11052 ( .B1(n9964), .B2(n9983), .A(n9963), .ZN(n9965) );
  AOI21_X1 U11053 ( .B1(n9966), .B2(n9989), .A(n9965), .ZN(n9967) );
  AND2_X1 U11054 ( .A1(n9968), .A2(n9967), .ZN(n10003) );
  INV_X1 U11055 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9969) );
  AOI22_X1 U11056 ( .A1(n9991), .A2(n10003), .B1(n9969), .B2(n9990), .ZN(
        P1_U3486) );
  OAI211_X1 U11057 ( .C1(n4850), .C2(n9983), .A(n9971), .B(n9970), .ZN(n9972)
         );
  AOI21_X1 U11058 ( .B1(n9973), .B2(n9979), .A(n9972), .ZN(n10004) );
  INV_X1 U11059 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9974) );
  AOI22_X1 U11060 ( .A1(n9991), .A2(n10004), .B1(n9974), .B2(n9990), .ZN(
        P1_U3489) );
  OAI211_X1 U11061 ( .C1(n9977), .C2(n9983), .A(n9976), .B(n9975), .ZN(n9978)
         );
  AOI21_X1 U11062 ( .B1(n9980), .B2(n9979), .A(n9978), .ZN(n10005) );
  INV_X1 U11063 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9981) );
  AOI22_X1 U11064 ( .A1(n9991), .A2(n10005), .B1(n9981), .B2(n9990), .ZN(
        P1_U3492) );
  OAI21_X1 U11065 ( .B1(n9984), .B2(n9983), .A(n9982), .ZN(n9987) );
  INV_X1 U11066 ( .A(n9985), .ZN(n9986) );
  AOI211_X1 U11067 ( .C1(n9989), .C2(n9988), .A(n9987), .B(n9986), .ZN(n10007)
         );
  AOI22_X1 U11068 ( .A1(n9991), .A2(n10007), .B1(n5989), .B2(n9990), .ZN(
        P1_U3495) );
  AOI22_X1 U11069 ( .A1(n10008), .A2(n9992), .B1(n5683), .B2(n10006), .ZN(
        P1_U3523) );
  AOI22_X1 U11070 ( .A1(n10008), .A2(n9993), .B1(n5720), .B2(n10006), .ZN(
        P1_U3524) );
  AOI22_X1 U11071 ( .A1(n10008), .A2(n9994), .B1(n5740), .B2(n10006), .ZN(
        P1_U3525) );
  AOI22_X1 U11072 ( .A1(n10008), .A2(n9995), .B1(n5755), .B2(n10006), .ZN(
        P1_U3526) );
  INV_X1 U11073 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9996) );
  AOI22_X1 U11074 ( .A1(n10008), .A2(n9997), .B1(n9996), .B2(n10006), .ZN(
        P1_U3527) );
  INV_X1 U11075 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9998) );
  AOI22_X1 U11076 ( .A1(n10008), .A2(n9999), .B1(n9998), .B2(n10006), .ZN(
        P1_U3528) );
  AOI22_X1 U11077 ( .A1(n10008), .A2(n10000), .B1(n5853), .B2(n10006), .ZN(
        P1_U3530) );
  AOI22_X1 U11078 ( .A1(n10008), .A2(n10001), .B1(n5868), .B2(n10006), .ZN(
        P1_U3531) );
  AOI22_X1 U11079 ( .A1(n10008), .A2(n10002), .B1(n6874), .B2(n10006), .ZN(
        P1_U3532) );
  AOI22_X1 U11080 ( .A1(n10008), .A2(n10003), .B1(n6877), .B2(n10006), .ZN(
        P1_U3533) );
  AOI22_X1 U11081 ( .A1(n10008), .A2(n10004), .B1(n5941), .B2(n10006), .ZN(
        P1_U3534) );
  AOI22_X1 U11082 ( .A1(n10008), .A2(n10005), .B1(n9033), .B2(n10006), .ZN(
        P1_U3535) );
  AOI22_X1 U11083 ( .A1(n10008), .A2(n10007), .B1(n9035), .B2(n10006), .ZN(
        P1_U3536) );
  INV_X1 U11084 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10009) );
  OAI22_X1 U11085 ( .A1(n10012), .A2(n10011), .B1(n10010), .B2(n10009), .ZN(
        n10013) );
  INV_X1 U11086 ( .A(n10013), .ZN(n10033) );
  OAI21_X1 U11087 ( .B1(n10016), .B2(n10015), .A(n10014), .ZN(n10030) );
  AOI21_X1 U11088 ( .B1(n10025), .B2(n10024), .A(n10023), .ZN(n10027) );
  NOR2_X1 U11089 ( .A1(n10027), .A2(n10026), .ZN(n10028) );
  AOI211_X1 U11090 ( .C1(n10031), .C2(n10030), .A(n10029), .B(n10028), .ZN(
        n10032) );
  OAI211_X1 U11091 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10034), .A(n10033), .B(
        n10032), .ZN(P2_U3199) );
  INV_X1 U11092 ( .A(n10035), .ZN(n10036) );
  AOI21_X1 U11093 ( .B1(n10037), .B2(n10081), .A(n10036), .ZN(n10038) );
  AOI211_X1 U11094 ( .C1(n10066), .C2(n10040), .A(n10039), .B(n10038), .ZN(
        n10088) );
  AOI22_X1 U11095 ( .A1(n10087), .A2(n4928), .B1(n10088), .B2(n10085), .ZN(
        P2_U3390) );
  OAI22_X1 U11096 ( .A1(n10041), .A2(n10069), .B1(n6979), .B2(n10079), .ZN(
        n10042) );
  NOR2_X1 U11097 ( .A1(n10043), .A2(n10042), .ZN(n10089) );
  AOI22_X1 U11098 ( .A1(n10087), .A2(n4584), .B1(n10089), .B2(n10085), .ZN(
        P2_U3396) );
  INV_X1 U11099 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10050) );
  INV_X1 U11100 ( .A(n10044), .ZN(n10048) );
  OAI21_X1 U11101 ( .B1(n10046), .B2(n10079), .A(n10045), .ZN(n10047) );
  AOI21_X1 U11102 ( .B1(n10049), .B2(n10048), .A(n10047), .ZN(n10090) );
  AOI22_X1 U11103 ( .A1(n10087), .A2(n10050), .B1(n10090), .B2(n10085), .ZN(
        P2_U3408) );
  INV_X1 U11104 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10055) );
  OAI22_X1 U11105 ( .A1(n10052), .A2(n10069), .B1(n10051), .B2(n10079), .ZN(
        n10053) );
  NOR2_X1 U11106 ( .A1(n10054), .A2(n10053), .ZN(n10092) );
  AOI22_X1 U11107 ( .A1(n10087), .A2(n10055), .B1(n10092), .B2(n10085), .ZN(
        P2_U3411) );
  INV_X1 U11108 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10061) );
  NOR2_X1 U11109 ( .A1(n10056), .A2(n10081), .ZN(n10059) );
  INV_X1 U11110 ( .A(n10057), .ZN(n10058) );
  AOI211_X1 U11111 ( .C1(n10066), .C2(n10060), .A(n10059), .B(n10058), .ZN(
        n10093) );
  AOI22_X1 U11112 ( .A1(n10087), .A2(n10061), .B1(n10093), .B2(n10085), .ZN(
        P2_U3414) );
  INV_X1 U11113 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10067) );
  NOR2_X1 U11114 ( .A1(n10062), .A2(n10069), .ZN(n10064) );
  AOI211_X1 U11115 ( .C1(n10066), .C2(n10065), .A(n10064), .B(n10063), .ZN(
        n10095) );
  AOI22_X1 U11116 ( .A1(n10087), .A2(n10067), .B1(n10095), .B2(n10085), .ZN(
        P2_U3417) );
  INV_X1 U11117 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10073) );
  OAI22_X1 U11118 ( .A1(n10070), .A2(n10069), .B1(n10068), .B2(n10079), .ZN(
        n10071) );
  NOR2_X1 U11119 ( .A1(n10072), .A2(n10071), .ZN(n10097) );
  AOI22_X1 U11120 ( .A1(n10087), .A2(n10073), .B1(n10097), .B2(n10085), .ZN(
        P2_U3420) );
  INV_X1 U11121 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10078) );
  OAI22_X1 U11122 ( .A1(n10075), .A2(n10081), .B1(n10074), .B2(n10079), .ZN(
        n10076) );
  NOR2_X1 U11123 ( .A1(n10077), .A2(n10076), .ZN(n10099) );
  AOI22_X1 U11124 ( .A1(n10087), .A2(n10078), .B1(n10099), .B2(n10085), .ZN(
        P2_U3423) );
  INV_X1 U11125 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10086) );
  OAI22_X1 U11126 ( .A1(n10082), .A2(n10081), .B1(n10080), .B2(n10079), .ZN(
        n10083) );
  NOR2_X1 U11127 ( .A1(n10084), .A2(n10083), .ZN(n10102) );
  AOI22_X1 U11128 ( .A1(n10087), .A2(n10086), .B1(n10102), .B2(n10085), .ZN(
        P2_U3426) );
  AOI22_X1 U11129 ( .A1(n10103), .A2(n10088), .B1(n6244), .B2(n10100), .ZN(
        P2_U3459) );
  AOI22_X1 U11130 ( .A1(n10103), .A2(n10089), .B1(n6247), .B2(n10100), .ZN(
        P2_U3461) );
  AOI22_X1 U11131 ( .A1(n10103), .A2(n10090), .B1(n6255), .B2(n10100), .ZN(
        P2_U3465) );
  AOI22_X1 U11132 ( .A1(n10103), .A2(n10092), .B1(n10091), .B2(n10100), .ZN(
        P2_U3466) );
  AOI22_X1 U11133 ( .A1(n10103), .A2(n10093), .B1(n6257), .B2(n10100), .ZN(
        P2_U3467) );
  AOI22_X1 U11134 ( .A1(n10103), .A2(n10095), .B1(n10094), .B2(n10100), .ZN(
        P2_U3468) );
  INV_X1 U11135 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10096) );
  AOI22_X1 U11136 ( .A1(n10103), .A2(n10097), .B1(n10096), .B2(n10100), .ZN(
        P2_U3469) );
  AOI22_X1 U11137 ( .A1(n10103), .A2(n10099), .B1(n10098), .B2(n10100), .ZN(
        P2_U3470) );
  AOI22_X1 U11138 ( .A1(n10103), .A2(n10102), .B1(n10101), .B2(n10100), .ZN(
        P2_U3471) );
  NOR2_X1 U11139 ( .A1(n10105), .A2(n10104), .ZN(n10106) );
  XOR2_X1 U11140 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10106), .Z(ADD_1068_U5) );
  XOR2_X1 U11141 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11142 ( .A1(n10108), .A2(n10107), .ZN(n10109) );
  XOR2_X1 U11143 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10109), .Z(ADD_1068_U55)
         );
  XNOR2_X1 U11144 ( .A(n10111), .B(n10110), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11145 ( .A(n10113), .B(n10112), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11146 ( .A(n10115), .B(n10114), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11147 ( .A(n10117), .B(n10116), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11148 ( .A(n10119), .B(n10118), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11149 ( .A(n10121), .B(n10120), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11150 ( .A(n10123), .B(n10122), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11151 ( .A(n10125), .B(n10124), .ZN(ADD_1068_U63) );
  XNOR2_X1 U11152 ( .A(n10127), .B(n10126), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11153 ( .A(n10129), .B(n10128), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11154 ( .A(n10131), .B(n10130), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11155 ( .A(n10133), .B(n10132), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11156 ( .A(n10135), .B(n10134), .ZN(ADD_1068_U48) );
  XOR2_X1 U11157 ( .A(n10137), .B(n10136), .Z(ADD_1068_U54) );
  XOR2_X1 U11158 ( .A(n10139), .B(n10138), .Z(ADD_1068_U53) );
  XNOR2_X1 U11159 ( .A(n10141), .B(n10140), .ZN(ADD_1068_U52) );
  INV_X1 U4785 ( .A(n6505), .ZN(n6111) );
  BUF_X1 U4855 ( .A(n4971), .Z(n5513) );
  BUF_X1 U5387 ( .A(n5647), .Z(n7232) );
  CLKBUF_X1 U4797 ( .A(n5673), .Z(n5675) );
  CLKBUF_X2 U4840 ( .A(n5718), .Z(n4273) );
  CLKBUF_X1 U4858 ( .A(n9919), .Z(n4271) );
  AND4_X1 U4989 ( .A1(n5760), .A2(n4804), .A3(n5622), .A4(n5725), .ZN(n10145)
         );
endmodule

