

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4380, n4381, n4382, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281;

  INV_X4 U4885 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U4886 ( .A(n6452), .ZN(n6460) );
  INV_X1 U4887 ( .A(n5180), .ZN(n7963) );
  CLKBUF_X1 U4888 ( .A(n5039), .Z(n5666) );
  AND3_X1 U4889 ( .A1(n5845), .A2(n5844), .A3(n5843), .ZN(n7316) );
  BUF_X2 U4891 ( .A(n5747), .Z(n6177) );
  CLKBUF_X2 U4892 ( .A(n7964), .Z(n4380) );
  CLKBUF_X2 U4893 ( .A(n5793), .Z(n8300) );
  NOR2_X1 U4894 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5011) );
  OAI211_X1 U4895 ( .C1(n6713), .C2(n6786), .A(n5837), .B(n5836), .ZN(n7273)
         );
  INV_X1 U4896 ( .A(n6456), .ZN(n6445) );
  INV_X1 U4897 ( .A(n6447), .ZN(n6462) );
  OR2_X1 U4899 ( .A1(n7105), .A2(n7106), .ZN(n7103) );
  INV_X1 U4900 ( .A(n5783), .ZN(n6609) );
  INV_X1 U4901 ( .A(n8540), .ZN(n9911) );
  AND2_X2 U4902 ( .A1(n7128), .A2(n6456), .ZN(n6447) );
  BUF_X1 U4903 ( .A(n5040), .Z(n5667) );
  NAND2_X1 U4904 ( .A1(n4982), .A2(n4981), .ZN(n5539) );
  NAND2_X1 U4905 ( .A1(n4438), .A2(n4632), .ZN(n5582) );
  OAI21_X1 U4906 ( .B1(n7305), .B2(n6344), .A(n6343), .ZN(n7550) );
  CLKBUF_X3 U4907 ( .A(n5072), .Z(n6553) );
  INV_X2 U4908 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  AOI21_X2 U4909 ( .B1(n8512), .B2(n8513), .A(n6165), .ZN(n6231) );
  NAND2_X1 U4910 ( .A1(n5026), .A2(n5741), .ZN(n7964) );
  NOR2_X2 U4911 ( .A1(n8863), .A2(n9037), .ZN(n8862) );
  AOI211_X2 U4912 ( .C1(n8178), .C2(n8177), .A(n8176), .B(n8175), .ZN(n8233)
         );
  AOI21_X2 U4913 ( .B1(n7344), .B2(n8396), .A(n7343), .ZN(n7372) );
  AND2_X1 U4914 ( .A1(n4470), .A2(n4468), .ZN(n4467) );
  AOI21_X1 U4915 ( .B1(n9290), .B2(n9586), .A(n4652), .ZN(n9436) );
  OR2_X1 U4916 ( .A1(n6493), .A2(n4946), .ZN(n6494) );
  OR2_X1 U4917 ( .A1(n7952), .A2(n4658), .ZN(n4657) );
  NOR2_X1 U4918 ( .A1(n8087), .A2(n8086), .ZN(n8203) );
  OAI22_X1 U4919 ( .A1(n9170), .A2(n9171), .B1(n6437), .B2(n6436), .ZN(n9162)
         );
  NAND2_X1 U4920 ( .A1(n8076), .A2(n4415), .ZN(n8073) );
  NAND2_X1 U4921 ( .A1(n8892), .A2(n8891), .ZN(n8890) );
  NOR2_X1 U4922 ( .A1(n9293), .A2(n9431), .ZN(n5663) );
  OR2_X1 U4923 ( .A1(n7581), .A2(n7578), .ZN(n6379) );
  NAND2_X1 U4924 ( .A1(n7713), .A2(n7712), .ZN(n7711) );
  NAND2_X1 U4925 ( .A1(n6357), .A2(n6356), .ZN(n7523) );
  NAND2_X1 U4926 ( .A1(n5203), .A2(n8005), .ZN(n9575) );
  AND2_X1 U4927 ( .A1(n7032), .A2(n7034), .ZN(n6305) );
  NAND2_X2 U4928 ( .A1(n7189), .A2(n9776), .ZN(n9785) );
  AND2_X1 U4929 ( .A1(n7435), .A2(n9812), .ZN(n7433) );
  XNOR2_X1 U4930 ( .A(n6286), .B(n6452), .ZN(n7415) );
  NOR2_X1 U4931 ( .A1(n7186), .A2(n9773), .ZN(n7435) );
  NAND2_X2 U4932 ( .A1(n6219), .A2(n8934), .ZN(n8629) );
  INV_X1 U4933 ( .A(n7209), .ZN(n9796) );
  NAND2_X1 U4934 ( .A1(n8315), .A2(n8352), .ZN(n7231) );
  NAND4_X1 U4935 ( .A1(n4999), .A2(n4998), .A3(n4997), .A4(n4996), .ZN(n9235)
         );
  INV_X1 U4936 ( .A(n5771), .ZN(n5792) );
  NAND2_X2 U4937 ( .A1(n6249), .A2(n6891), .ZN(n6452) );
  AND2_X2 U4938 ( .A1(n6249), .A2(n6478), .ZN(n6456) );
  AND2_X1 U4939 ( .A1(n6226), .A2(n6856), .ZN(n5771) );
  INV_X1 U4940 ( .A(n6922), .ZN(n6832) );
  OAI211_X1 U4941 ( .C1(n7060), .C2(n5767), .A(n4849), .B(n5768), .ZN(n8663)
         );
  BUF_X2 U4942 ( .A(n5079), .Z(n5561) );
  NOR2_X1 U4943 ( .A1(n5701), .A2(n5700), .ZN(n7115) );
  INV_X2 U4944 ( .A(n4385), .ZN(n4382) );
  INV_X1 U4945 ( .A(n6035), .ZN(n8855) );
  AOI21_X1 U4946 ( .B1(n5071), .B2(n5070), .A(n4954), .ZN(n5128) );
  CLKBUF_X1 U4947 ( .A(n5558), .Z(n4384) );
  OR2_X1 U4948 ( .A1(n4409), .A2(n4978), .ZN(n4984) );
  XNOR2_X1 U4949 ( .A(n5358), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9349) );
  NAND2_X2 U4950 ( .A1(n5694), .A2(n5698), .ZN(n5766) );
  NAND2_X1 U4951 ( .A1(n4465), .A2(n5034), .ZN(n5048) );
  NAND2_X1 U4952 ( .A1(n6715), .A2(n6233), .ZN(n5773) );
  INV_X1 U4953 ( .A(n5698), .ZN(n7788) );
  XNOR2_X1 U4954 ( .A(n5714), .B(n5713), .ZN(n6233) );
  INV_X2 U4955 ( .A(n9535), .ZN(n7920) );
  NAND2_X1 U4956 ( .A1(n5712), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5714) );
  NAND2_X1 U4957 ( .A1(n5690), .A2(n5706), .ZN(n5691) );
  NAND2_X1 U4958 ( .A1(n4904), .A2(n4972), .ZN(n4903) );
  NOR2_X1 U4959 ( .A1(n4964), .A2(n4963), .ZN(n5356) );
  AND3_X1 U4960 ( .A1(n4922), .A2(n4924), .A3(n5683), .ZN(n5882) );
  AND2_X1 U4961 ( .A1(n4924), .A2(n4832), .ZN(n4831) );
  AND2_X1 U4962 ( .A1(n5707), .A2(n5689), .ZN(n5711) );
  NAND2_X1 U4963 ( .A1(n4439), .A2(n4906), .ZN(n4905) );
  NAND2_X2 U4964 ( .A1(n4586), .A2(n4987), .ZN(n5134) );
  AND4_X1 U4965 ( .A1(n4851), .A2(n4955), .A3(n5011), .A4(n4850), .ZN(n5061)
         );
  AND2_X1 U4966 ( .A1(n5686), .A2(n6186), .ZN(n6182) );
  AND2_X1 U4967 ( .A1(n4511), .A2(n4510), .ZN(n5796) );
  INV_X1 U4968 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5715) );
  NOR2_X1 U4969 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4955) );
  NOR2_X1 U4970 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5831) );
  NOR2_X1 U4971 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n6186) );
  NOR2_X2 U4972 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7706) );
  INV_X1 U4973 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5721) );
  INV_X1 U4974 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5948) );
  NAND2_X1 U4975 ( .A1(n5231), .A2(n5230), .ZN(n5263) );
  OAI21_X1 U4976 ( .B1(n5691), .B2(n4719), .A(n4717), .ZN(n4716) );
  NAND2_X1 U4977 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(n4720), .ZN(n4719) );
  INV_X1 U4978 ( .A(n4718), .ZN(n4717) );
  OAI22_X1 U4979 ( .A1(n4721), .A2(n4720), .B1(P2_IR_REG_31__SCAN_IN), .B2(
        n9124), .ZN(n4718) );
  INV_X1 U4980 ( .A(n6291), .ZN(n4547) );
  OAI21_X1 U4981 ( .B1(n8121), .B2(n4885), .A(n4888), .ZN(n4884) );
  NAND2_X1 U4982 ( .A1(n4889), .A2(n9312), .ZN(n4888) );
  OR2_X1 U4983 ( .A1(n9438), .A2(n9312), .ZN(n8182) );
  NAND2_X1 U4984 ( .A1(n4749), .A2(n4748), .ZN(n5228) );
  AOI21_X1 U4985 ( .B1(n4387), .B2(n4754), .A(n4437), .ZN(n4749) );
  AND2_X1 U4986 ( .A1(n4981), .A2(n7919), .ZN(n5039) );
  OR2_X1 U4987 ( .A1(n5492), .A2(n9978), .ZN(n5523) );
  NAND2_X1 U4988 ( .A1(n8159), .A2(n8079), .ZN(n4502) );
  NAND2_X1 U4989 ( .A1(n8028), .A2(n4491), .ZN(n8027) );
  AND2_X1 U4990 ( .A1(n8946), .A2(n8947), .ZN(n8282) );
  OR2_X1 U4991 ( .A1(n4540), .A2(n4538), .ZN(n4537) );
  NOR2_X1 U4992 ( .A1(n4756), .A2(n4539), .ZN(n4538) );
  NAND2_X1 U4993 ( .A1(n9156), .A2(n9192), .ZN(n4756) );
  NAND2_X1 U4994 ( .A1(n4430), .A2(n4388), .ZN(n4865) );
  INV_X1 U4995 ( .A(n4583), .ZN(n4582) );
  OR2_X1 U4996 ( .A1(n9052), .A2(n8786), .ZN(n8448) );
  OR2_X1 U4997 ( .A1(n9083), .A2(n7896), .ZN(n8433) );
  INV_X1 U4998 ( .A(n8324), .ZN(n4711) );
  NOR2_X1 U4999 ( .A1(n8662), .A2(n7152), .ZN(n8311) );
  NAND2_X1 U5000 ( .A1(n6922), .A2(n6833), .ZN(n8360) );
  AND2_X1 U5001 ( .A1(n6035), .A2(n8501), .ZN(n8337) );
  NAND2_X1 U5002 ( .A1(n5773), .A2(n6553), .ZN(n5793) );
  AND2_X1 U5003 ( .A1(n5687), .A2(n6182), .ZN(n5707) );
  INV_X1 U5004 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5687) );
  AND2_X1 U5005 ( .A1(n4921), .A2(n5795), .ZN(n4922) );
  AND2_X1 U5006 ( .A1(n5685), .A2(n5833), .ZN(n4921) );
  INV_X1 U5007 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5685) );
  INV_X1 U5008 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U5009 ( .A1(n5722), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U5010 ( .A1(n4939), .A2(n5720), .ZN(n4938) );
  INV_X1 U5011 ( .A(n4940), .ZN(n4939) );
  AND2_X1 U5012 ( .A1(n6326), .A2(n4785), .ZN(n4784) );
  NAND2_X1 U5013 ( .A1(n7521), .A2(n7524), .ZN(n4765) );
  OR2_X1 U5014 ( .A1(n8088), .A2(n5565), .ZN(n8238) );
  NOR2_X1 U5015 ( .A1(n8121), .A2(n4887), .ZN(n4886) );
  INV_X1 U5016 ( .A(n5649), .ZN(n4887) );
  OR2_X1 U5017 ( .A1(n9434), .A2(n9139), .ZN(n8129) );
  NAND2_X1 U5018 ( .A1(n5653), .A2(n9778), .ZN(n6891) );
  XNOR2_X1 U5019 ( .A(n7957), .B(n7956), .ZN(n7954) );
  AND2_X1 U5020 ( .A1(n5517), .A2(n5516), .ZN(n5532) );
  AOI21_X1 U5021 ( .B1(n4608), .B2(n4606), .A(n4462), .ZN(n4605) );
  NAND2_X1 U5022 ( .A1(n5552), .A2(n5551), .ZN(n4553) );
  NAND2_X1 U5023 ( .A1(n5352), .A2(n5351), .ZN(n5367) );
  NAND2_X1 U5024 ( .A1(n5349), .A2(n5348), .ZN(n5352) );
  NAND2_X1 U5025 ( .A1(n5286), .A2(n5273), .ZN(n5287) );
  NAND2_X1 U5026 ( .A1(n5269), .A2(n5268), .ZN(n5288) );
  NAND2_X1 U5027 ( .A1(n4483), .A2(n4479), .ZN(n4478) );
  NAND2_X1 U5028 ( .A1(n4486), .A2(n4480), .ZN(n4479) );
  AOI21_X1 U5029 ( .B1(n4488), .B2(n4485), .A(n4484), .ZN(n4483) );
  INV_X1 U5030 ( .A(n5263), .ZN(n4484) );
  INV_X1 U5031 ( .A(n5226), .ZN(n4485) );
  AND2_X1 U5032 ( .A1(n5263), .A2(n5233), .ZN(n5246) );
  AND2_X1 U5033 ( .A1(n4574), .A2(n5187), .ZN(n5185) );
  NAND2_X1 U5034 ( .A1(n4575), .A2(SI_10_), .ZN(n4574) );
  INV_X1 U5035 ( .A(n4576), .ZN(n4575) );
  NAND2_X1 U5036 ( .A1(n5179), .A2(n5155), .ZN(n5157) );
  NAND2_X1 U5037 ( .A1(n5125), .A2(n5124), .ZN(n5130) );
  INV_X1 U5038 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4851) );
  NAND2_X1 U5039 ( .A1(n5002), .A2(n5705), .ZN(n5016) );
  NAND2_X1 U5040 ( .A1(n7929), .A2(n7788), .ZN(n5736) );
  AND2_X1 U5041 ( .A1(n4739), .A2(n4736), .ZN(n4731) );
  AND2_X1 U5042 ( .A1(n4737), .A2(n6216), .ZN(n4736) );
  AOI21_X1 U5043 ( .B1(n4436), .B2(n6216), .A(n4733), .ZN(n4732) );
  INV_X1 U5044 ( .A(n4735), .ZN(n4733) );
  OAI211_X1 U5045 ( .C1(n8491), .C2(n4385), .A(n6216), .B(n4619), .ZN(n4735)
         );
  INV_X1 U5046 ( .A(n5753), .ZN(n6234) );
  NAND2_X1 U5048 ( .A1(n8695), .A2(n4521), .ZN(n4520) );
  OR2_X1 U5049 ( .A1(n9037), .A2(n8883), .ZN(n8846) );
  XNOR2_X1 U5050 ( .A(n9045), .B(n8647), .ZN(n8891) );
  AOI21_X1 U5051 ( .B1(n4697), .B2(n4695), .A(n4428), .ZN(n4694) );
  INV_X1 U5052 ( .A(n8780), .ZN(n4695) );
  OR2_X1 U5053 ( .A1(n9079), .A2(n8996), .ZN(n8776) );
  INV_X1 U5054 ( .A(n5794), .ZN(n8299) );
  INV_X1 U5055 ( .A(n8300), .ZN(n6036) );
  INV_X1 U5056 ( .A(n6713), .ZN(n6590) );
  INV_X1 U5057 ( .A(n7091), .ZN(n8381) );
  NAND2_X1 U5058 ( .A1(n4679), .A2(n4678), .ZN(n7280) );
  AND2_X1 U5059 ( .A1(n8381), .A2(n4411), .ZN(n4678) );
  AND2_X1 U5060 ( .A1(n8383), .A2(n8384), .ZN(n7091) );
  NAND2_X1 U5062 ( .A1(n8662), .A2(n7152), .ZN(n6948) );
  CLKBUF_X1 U5063 ( .A(n6035), .Z(n8342) );
  NAND2_X1 U5064 ( .A1(n5691), .A2(n4714), .ZN(n4713) );
  INV_X1 U5065 ( .A(n4721), .ZN(n4714) );
  NAND2_X1 U5066 ( .A1(n5691), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5692) );
  AND2_X1 U5067 ( .A1(n4546), .A2(n4544), .ZN(n7031) );
  NAND2_X1 U5068 ( .A1(n4547), .A2(n4545), .ZN(n4544) );
  INV_X1 U5069 ( .A(n7253), .ZN(n4545) );
  INV_X1 U5070 ( .A(n9320), .ZN(n9135) );
  AOI21_X1 U5071 ( .B1(n4558), .B2(n4562), .A(n4556), .ZN(n4555) );
  INV_X1 U5072 ( .A(n4558), .ZN(n4557) );
  INV_X1 U5073 ( .A(n7906), .ZN(n4556) );
  NAND2_X1 U5074 ( .A1(n6252), .A2(n4952), .ZN(n6687) );
  NAND2_X1 U5075 ( .A1(n7520), .A2(n4765), .ZN(n6340) );
  OR2_X1 U5076 ( .A1(n9426), .A2(n8084), .ZN(n8204) );
  INV_X1 U5077 ( .A(n8252), .ZN(n4475) );
  AND2_X1 U5078 ( .A1(n8182), .A2(n8185), .ZN(n8121) );
  AOI21_X1 U5079 ( .B1(n9137), .B2(n5512), .A(n5511), .ZN(n9312) );
  OR2_X1 U5080 ( .A1(n5571), .A2(n9217), .ZN(n5648) );
  OAI21_X1 U5081 ( .B1(n7777), .B2(n5635), .A(n5634), .ZN(n7855) );
  INV_X1 U5082 ( .A(n4381), .ZN(n5359) );
  NAND2_X1 U5083 ( .A1(n5557), .A2(n9586), .ZN(n5570) );
  NAND2_X1 U5084 ( .A1(n4977), .A2(n4976), .ZN(n4982) );
  OR2_X1 U5085 ( .A1(n4979), .A2(n4978), .ZN(n4980) );
  NAND2_X1 U5086 ( .A1(n5538), .A2(n5537), .ZN(n9431) );
  NAND2_X1 U5087 ( .A1(n8009), .A2(n8081), .ZN(n4504) );
  NAND2_X1 U5088 ( .A1(n8015), .A2(n8004), .ZN(n8013) );
  INV_X1 U5089 ( .A(n8069), .ZN(n4499) );
  NAND2_X1 U5090 ( .A1(n8059), .A2(n8079), .ZN(n4501) );
  NAND2_X1 U5091 ( .A1(n8060), .A2(n8081), .ZN(n4500) );
  INV_X1 U5092 ( .A(n8068), .ZN(n4497) );
  INV_X1 U5093 ( .A(n9288), .ZN(n4496) );
  OAI21_X1 U5094 ( .B1(n4728), .B2(n8461), .A(n4724), .ZN(n4723) );
  AOI21_X1 U5095 ( .B1(n4729), .B2(n4382), .A(n8460), .ZN(n4728) );
  OAI21_X1 U5096 ( .B1(n4727), .B2(n4725), .A(n4385), .ZN(n4724) );
  AND2_X1 U5097 ( .A1(n8871), .A2(n4449), .ZN(n4722) );
  NAND2_X1 U5098 ( .A1(n4600), .A2(n4598), .ZN(n8490) );
  NOR2_X1 U5099 ( .A1(n8764), .A2(n4599), .ZN(n4598) );
  INV_X1 U5100 ( .A(n8301), .ZN(n4599) );
  NOR2_X1 U5101 ( .A1(n4757), .A2(n4755), .ZN(n4543) );
  INV_X1 U5102 ( .A(n9192), .ZN(n4755) );
  INV_X1 U5103 ( .A(n4593), .ZN(n4592) );
  NAND2_X1 U5104 ( .A1(n5287), .A2(n5286), .ZN(n4597) );
  NAND2_X1 U5105 ( .A1(n4482), .A2(n4488), .ZN(n5265) );
  NAND2_X1 U5106 ( .A1(n5228), .A2(n5226), .ZN(n4482) );
  NAND2_X1 U5107 ( .A1(n4576), .A2(n5158), .ZN(n5187) );
  AOI21_X1 U5108 ( .B1(n4918), .B2(n4920), .A(n4432), .ZN(n4916) );
  AND2_X1 U5109 ( .A1(n8797), .A2(n4441), .ZN(n4737) );
  NOR2_X1 U5110 ( .A1(n4623), .A2(n9020), .ZN(n4622) );
  INV_X1 U5111 ( .A(n4624), .ZN(n4623) );
  AND2_X1 U5112 ( .A1(n8833), .A2(n8834), .ZN(n8285) );
  NOR2_X1 U5113 ( .A1(n9025), .A2(n9031), .ZN(n4624) );
  NOR2_X1 U5114 ( .A1(n8830), .A2(n8646), .ZN(n8468) );
  OR2_X1 U5115 ( .A1(n9031), .A2(n8837), .ZN(n8467) );
  NOR2_X1 U5116 ( .A1(n9068), .A2(n9072), .ZN(n4630) );
  INV_X1 U5117 ( .A(n8437), .ZN(n4844) );
  AND2_X1 U5118 ( .A1(n4844), .A2(n8326), .ZN(n4843) );
  NOR2_X1 U5119 ( .A1(n8436), .A2(n4846), .ZN(n4845) );
  OR2_X1 U5120 ( .A1(n7841), .A2(n7898), .ZN(n8420) );
  OR2_X1 U5121 ( .A1(n9089), .A2(n7838), .ZN(n8414) );
  NAND2_X1 U5122 ( .A1(n5811), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U5123 ( .A1(n7325), .A2(n8661), .ZN(n8366) );
  NAND2_X1 U5124 ( .A1(n6832), .A2(n8550), .ZN(n8310) );
  OR2_X1 U5125 ( .A1(n5794), .A2(n5775), .ZN(n5777) );
  NAND2_X1 U5126 ( .A1(n7706), .A2(n4986), .ZN(n4586) );
  INV_X1 U5127 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4986) );
  NAND2_X1 U5128 ( .A1(n7705), .A2(n4985), .ZN(n4987) );
  INV_X1 U5129 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4985) );
  NOR2_X1 U5130 ( .A1(n6405), .A2(n7883), .ZN(n4773) );
  INV_X1 U5131 ( .A(n6451), .ZN(n4779) );
  NAND2_X1 U5132 ( .A1(n4762), .A2(n4761), .ZN(n4760) );
  NAND2_X1 U5133 ( .A1(n6427), .A2(n6426), .ZN(n4761) );
  NAND2_X1 U5134 ( .A1(n9156), .A2(n4763), .ZN(n4762) );
  NOR2_X1 U5135 ( .A1(n4767), .A2(n4766), .ZN(n4774) );
  INV_X1 U5136 ( .A(n6399), .ZN(n4766) );
  INV_X1 U5137 ( .A(n7824), .ZN(n4767) );
  INV_X1 U5138 ( .A(n4807), .ZN(n9240) );
  INV_X1 U5139 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4962) );
  AND2_X1 U5140 ( .A1(n5140), .A2(n4569), .ZN(n4568) );
  INV_X1 U5141 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4569) );
  OAI21_X1 U5142 ( .B1(n9319), .B2(n5482), .A(n8180), .ZN(n9308) );
  INV_X1 U5143 ( .A(n9323), .ZN(n5482) );
  OR2_X1 U5144 ( .A1(n9443), .A2(n9135), .ZN(n8181) );
  NAND2_X1 U5145 ( .A1(n9455), .A2(n7968), .ZN(n4901) );
  AND2_X1 U5146 ( .A1(n4901), .A2(n4899), .ZN(n4892) );
  OR2_X1 U5147 ( .A1(n5571), .A2(n9341), .ZN(n8180) );
  NAND2_X1 U5148 ( .A1(n5445), .A2(n5444), .ZN(n8258) );
  OR2_X1 U5149 ( .A1(n9460), .A2(n9340), .ZN(n8173) );
  INV_X1 U5150 ( .A(n9394), .ZN(n4645) );
  NOR2_X1 U5151 ( .A1(n9379), .A2(n4648), .ZN(n4647) );
  NAND2_X1 U5152 ( .A1(n8114), .A2(n5640), .ZN(n4857) );
  INV_X1 U5153 ( .A(n5640), .ZN(n4854) );
  OR2_X1 U5154 ( .A1(n9476), .A2(n5388), .ZN(n8034) );
  AND2_X1 U5155 ( .A1(n7846), .A2(n9221), .ZN(n8150) );
  OR2_X1 U5156 ( .A1(n7751), .A2(n5259), .ZN(n8015) );
  AOI21_X1 U5157 ( .B1(n4865), .B2(n4863), .A(n4435), .ZN(n4862) );
  INV_X1 U5158 ( .A(n4399), .ZN(n4863) );
  INV_X1 U5159 ( .A(n4865), .ZN(n4864) );
  OR2_X1 U5160 ( .A1(n9594), .A2(n9501), .ZN(n7746) );
  OR2_X1 U5161 ( .A1(n7574), .A2(n7935), .ZN(n7999) );
  NOR2_X1 U5162 ( .A1(n9303), .A2(n9438), .ZN(n9292) );
  NAND2_X1 U5163 ( .A1(n4581), .A2(n4579), .ZN(n7957) );
  AOI21_X1 U5164 ( .B1(n4583), .B2(n4580), .A(n4461), .ZN(n4579) );
  OR2_X1 U5165 ( .A1(n5532), .A2(n4582), .ZN(n4581) );
  AND2_X1 U5166 ( .A1(n4983), .A2(n4391), .ZN(n4635) );
  NAND2_X1 U5167 ( .A1(n4969), .A2(n4908), .ZN(n4907) );
  INV_X1 U5168 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4969) );
  INV_X1 U5169 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4908) );
  AOI21_X1 U5170 ( .B1(n4613), .B2(n4445), .A(n4612), .ZN(n4611) );
  NOR2_X1 U5171 ( .A1(n5410), .A2(n4618), .ZN(n4617) );
  INV_X1 U5172 ( .A(n5391), .ZN(n4618) );
  NAND2_X1 U5173 ( .A1(n5550), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5552) );
  AND2_X1 U5174 ( .A1(n5391), .A2(n5375), .ZN(n5389) );
  AOI21_X1 U5175 ( .B1(n4402), .B2(n4595), .A(n4594), .ZN(n4593) );
  INV_X1 U5176 ( .A(n5310), .ZN(n4594) );
  INV_X1 U5177 ( .A(n5286), .ZN(n4595) );
  INV_X1 U5178 ( .A(n4402), .ZN(n4596) );
  OR2_X1 U5179 ( .A1(n5766), .A2(n7248), .ZN(n5696) );
  NAND2_X1 U5180 ( .A1(n5936), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U5181 ( .A1(n4931), .A2(n5889), .ZN(n4930) );
  INV_X1 U5182 ( .A(n7609), .ZN(n4931) );
  AND2_X1 U5183 ( .A1(n6018), .A2(n6002), .ZN(n4934) );
  INV_X1 U5184 ( .A(n6506), .ZN(n6018) );
  AND4_X1 U5185 ( .A1(n6059), .A2(n6058), .A3(n6057), .A4(n6056), .ZN(n8648)
         );
  OR2_X1 U5186 ( .A1(n6767), .A2(n6766), .ZN(n4531) );
  OR2_X1 U5187 ( .A1(n6796), .A2(n6795), .ZN(n4529) );
  NAND2_X1 U5188 ( .A1(n8718), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4525) );
  AOI21_X1 U5189 ( .B1(n8729), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8728), .ZN(
        n8747) );
  AOI21_X1 U5190 ( .B1(n8755), .B2(n9853), .A(n8342), .ZN(n4519) );
  NOR2_X1 U5191 ( .A1(n8800), .A2(n8768), .ZN(n8767) );
  NAND2_X1 U5192 ( .A1(n8813), .A2(n8808), .ZN(n8819) );
  XNOR2_X1 U5193 ( .A(n9020), .B(n8795), .ZN(n8808) );
  NAND2_X1 U5194 ( .A1(n9031), .A2(n8837), .ZN(n8834) );
  NAND2_X1 U5195 ( .A1(n8862), .A2(n8763), .ZN(n8852) );
  OR2_X1 U5196 ( .A1(n9031), .A2(n8789), .ZN(n8790) );
  NAND2_X1 U5197 ( .A1(n8890), .A2(n4413), .ZN(n8885) );
  AND4_X1 U5198 ( .A1(n6134), .A2(n6133), .A3(n6132), .A4(n6131), .ZN(n8883)
         );
  NOR2_X1 U5199 ( .A1(n8284), .A2(n4705), .ZN(n4703) );
  INV_X1 U5200 ( .A(n8891), .ZN(n8903) );
  INV_X1 U5201 ( .A(n4838), .ZN(n4837) );
  AOI21_X1 U5202 ( .B1(n4836), .B2(n4838), .A(n4835), .ZN(n4834) );
  NOR2_X1 U5203 ( .A1(n8930), .A2(n4839), .ZN(n4838) );
  OR2_X1 U5204 ( .A1(n9057), .A2(n8783), .ZN(n8784) );
  AND2_X1 U5205 ( .A1(n8453), .A2(n8449), .ZN(n8946) );
  OR2_X1 U5206 ( .A1(n9068), .A2(n8994), .ZN(n4699) );
  INV_X1 U5207 ( .A(n8946), .ZN(n8940) );
  OR2_X1 U5208 ( .A1(n7821), .A2(n4682), .ZN(n8777) );
  NAND2_X1 U5209 ( .A1(n8436), .A2(n4683), .ZN(n4682) );
  INV_X1 U5210 ( .A(n4687), .ZN(n4683) );
  AND2_X1 U5211 ( .A1(n7794), .A2(n4684), .ZN(n7821) );
  NOR2_X1 U5212 ( .A1(n8326), .A2(n4685), .ZN(n4684) );
  INV_X1 U5213 ( .A(n7793), .ZN(n4685) );
  NAND2_X1 U5214 ( .A1(n7792), .A2(n8326), .ZN(n7810) );
  NAND2_X1 U5215 ( .A1(n4826), .A2(n7535), .ZN(n4822) );
  NOR2_X1 U5216 ( .A1(n8416), .A2(n4825), .ZN(n4824) );
  OAI21_X1 U5217 ( .B1(n7371), .B2(n4708), .A(n4706), .ZN(n7635) );
  INV_X1 U5218 ( .A(n4709), .ZN(n4708) );
  AOI21_X1 U5219 ( .B1(n4709), .B2(n4707), .A(n4425), .ZN(n4706) );
  NOR2_X1 U5220 ( .A1(n7498), .A2(n9089), .ZN(n7540) );
  AND2_X1 U5221 ( .A1(n7491), .A2(n4712), .ZN(n4709) );
  NAND2_X1 U5222 ( .A1(n7371), .A2(n4400), .ZN(n4710) );
  AND2_X1 U5223 ( .A1(n8402), .A2(n8396), .ZN(n8395) );
  AND4_X1 U5224 ( .A1(n5881), .A2(n5880), .A3(n5879), .A4(n5878), .ZN(n7286)
         );
  NAND2_X1 U5225 ( .A1(n4821), .A2(n4460), .ZN(n4819) );
  AND2_X1 U5226 ( .A1(n7091), .A2(n8379), .ZN(n4815) );
  NAND2_X1 U5227 ( .A1(n4681), .A2(n4680), .ZN(n6943) );
  AND2_X1 U5228 ( .A1(n4951), .A2(n6842), .ZN(n4680) );
  NAND2_X1 U5229 ( .A1(n7155), .A2(n7156), .ZN(n4681) );
  AND3_X1 U5230 ( .A1(n5800), .A2(n5799), .A3(n5798), .ZN(n7152) );
  OR2_X1 U5231 ( .A1(n5794), .A2(n10255), .ZN(n5799) );
  INV_X1 U5232 ( .A(n8663), .ZN(n7144) );
  INV_X1 U5233 ( .A(n8970), .ZN(n8998) );
  OR2_X1 U5234 ( .A1(n7115), .A2(n9872), .ZN(n7121) );
  NAND2_X1 U5235 ( .A1(n7115), .A2(n8507), .ZN(n7247) );
  NAND2_X1 U5236 ( .A1(n6078), .A2(n6077), .ZN(n9052) );
  NAND2_X1 U5237 ( .A1(n6006), .A2(n6005), .ZN(n9079) );
  INV_X1 U5238 ( .A(n7325), .ZN(n8586) );
  OR2_X1 U5239 ( .A1(n5793), .A2(n6556), .ZN(n5746) );
  OR2_X1 U5240 ( .A1(n5794), .A2(n6555), .ZN(n5745) );
  AND2_X1 U5241 ( .A1(n5713), .A2(n5711), .ZN(n5690) );
  AND3_X1 U5242 ( .A1(n5682), .A2(n4410), .A3(n5681), .ZN(n5684) );
  AND2_X1 U5243 ( .A1(n5680), .A2(n5679), .ZN(n5681) );
  AND4_X1 U5244 ( .A1(n5948), .A2(n4941), .A3(n5715), .A4(n5718), .ZN(n5682)
         );
  XNOR2_X1 U5245 ( .A(n5724), .B(n5723), .ZN(n6215) );
  NAND2_X1 U5246 ( .A1(n5727), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5724) );
  AND2_X1 U5247 ( .A1(n5728), .A2(n5727), .ZN(n6035) );
  NAND2_X1 U5248 ( .A1(n5719), .A2(n4941), .ZN(n4940) );
  INV_X1 U5249 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4511) );
  INV_X1 U5250 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4510) );
  AND2_X1 U5251 ( .A1(n4768), .A2(n4559), .ZN(n4558) );
  OR2_X1 U5252 ( .A1(n4773), .A2(n4560), .ZN(n4559) );
  AND2_X1 U5253 ( .A1(n4769), .A2(n4771), .ZN(n4768) );
  NAND2_X1 U5254 ( .A1(n7826), .A2(n4561), .ZN(n4560) );
  OR2_X1 U5255 ( .A1(n4773), .A2(n4563), .ZN(n4562) );
  INV_X1 U5256 ( .A(n7826), .ZN(n4563) );
  NOR2_X1 U5257 ( .A1(n4779), .A2(n4777), .ZN(n4776) );
  INV_X1 U5258 ( .A(n9163), .ZN(n4777) );
  OR2_X1 U5259 ( .A1(n4780), .A2(n4779), .ZN(n4778) );
  NAND2_X1 U5260 ( .A1(n6306), .A2(n7031), .ZN(n7161) );
  AND2_X1 U5261 ( .A1(n6305), .A2(n6304), .ZN(n6306) );
  AOI21_X1 U5262 ( .B1(n7031), .B2(n6305), .A(n6301), .ZN(n6303) );
  OR2_X1 U5263 ( .A1(n5381), .A2(n5380), .ZN(n5397) );
  INV_X1 U5264 ( .A(n6340), .ZN(n6337) );
  NAND2_X1 U5265 ( .A1(n4760), .A2(n4758), .ZN(n4759) );
  OR2_X1 U5266 ( .A1(n6411), .A2(n6410), .ZN(n6412) );
  NOR2_X1 U5267 ( .A1(n4407), .A2(n4539), .ZN(n4540) );
  NOR2_X1 U5268 ( .A1(n4760), .A2(n4758), .ZN(n4757) );
  NAND2_X1 U5269 ( .A1(n9178), .A2(n9179), .ZN(n9177) );
  NAND3_X1 U5270 ( .A1(n7162), .A2(n4532), .A3(n7163), .ZN(n7932) );
  INV_X1 U5271 ( .A(n7934), .ZN(n4532) );
  NAND2_X1 U5272 ( .A1(n4774), .A2(n6404), .ZN(n7885) );
  OAI22_X1 U5273 ( .A1(n7022), .A2(n6444), .B1(n9812), .B2(n6445), .ZN(n6281)
         );
  AND2_X1 U5274 ( .A1(n9205), .A2(n4781), .ZN(n4780) );
  NAND2_X1 U5275 ( .A1(n5254), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5281) );
  INV_X1 U5276 ( .A(n5255), .ZN(n5254) );
  NAND2_X1 U5277 ( .A1(n5548), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U5278 ( .A1(n5102), .A2(n4566), .ZN(n5548) );
  NOR2_X1 U5279 ( .A1(n5357), .A2(n4567), .ZN(n4566) );
  NAND2_X1 U5280 ( .A1(n4568), .A2(n5547), .ZN(n4567) );
  AND2_X1 U5281 ( .A1(n4982), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4871) );
  NAND2_X1 U5282 ( .A1(n9634), .A2(n4812), .ZN(n4811) );
  NAND2_X1 U5283 ( .A1(n9628), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4812) );
  INV_X1 U5284 ( .A(n6703), .ZN(n4801) );
  AOI21_X1 U5285 ( .B1(n6702), .B2(n4806), .A(n9646), .ZN(n4802) );
  NOR2_X1 U5286 ( .A1(n6814), .A2(n4799), .ZN(n6818) );
  AND2_X1 U5287 ( .A1(n6815), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4799) );
  OR2_X1 U5288 ( .A1(n6818), .A2(n6817), .ZN(n4798) );
  OAI21_X1 U5289 ( .B1(n9713), .B2(n4790), .A(n4789), .ZN(n9724) );
  NAND2_X1 U5290 ( .A1(n4793), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4790) );
  NAND2_X1 U5291 ( .A1(n9243), .A2(n4793), .ZN(n4789) );
  INV_X1 U5292 ( .A(n9725), .ZN(n4793) );
  OR2_X1 U5293 ( .A1(n9713), .A2(n5283), .ZN(n4792) );
  INV_X1 U5294 ( .A(n4568), .ZN(n4565) );
  OAI21_X1 U5295 ( .B1(n5445), .B2(n4640), .A(n4637), .ZN(n9319) );
  AOI21_X1 U5296 ( .B1(n4639), .B2(n8260), .A(n4638), .ZN(n4637) );
  INV_X1 U5297 ( .A(n7970), .ZN(n4638) );
  NOR2_X1 U5298 ( .A1(n5647), .A2(n4900), .ZN(n4899) );
  INV_X1 U5299 ( .A(n4902), .ZN(n4900) );
  AOI21_X1 U5300 ( .B1(n4898), .B2(n4897), .A(n4896), .ZN(n4895) );
  INV_X1 U5301 ( .A(n8049), .ZN(n4896) );
  INV_X1 U5302 ( .A(n5647), .ZN(n4898) );
  AND2_X1 U5303 ( .A1(n5646), .A2(n4902), .ZN(n4897) );
  OR2_X1 U5304 ( .A1(n9465), .A2(n9366), .ZN(n4902) );
  AOI21_X1 U5305 ( .B1(n9355), .B2(n5645), .A(n4945), .ZN(n8266) );
  NAND2_X1 U5306 ( .A1(n9395), .A2(n9394), .ZN(n4649) );
  OR2_X1 U5307 ( .A1(n9388), .A2(n9476), .ZN(n9372) );
  AND2_X1 U5308 ( .A1(n8029), .A2(n8165), .ZN(n9394) );
  NAND2_X1 U5309 ( .A1(n4858), .A2(n9412), .ZN(n9404) );
  OAI21_X1 U5310 ( .B1(n7779), .B2(n8150), .A(n8156), .ZN(n7856) );
  OAI22_X1 U5311 ( .A1(n7739), .A2(n5633), .B1(n9222), .B2(n7751), .ZN(n7777)
         );
  OAI21_X1 U5312 ( .B1(n9575), .B2(n5225), .A(n8007), .ZN(n7772) );
  OR2_X1 U5313 ( .A1(n9592), .A2(n9593), .ZN(n9594) );
  NAND2_X1 U5314 ( .A1(n7386), .A2(n7385), .ZN(n7403) );
  NAND2_X1 U5315 ( .A1(n7177), .A2(n4852), .ZN(n7019) );
  AND2_X1 U5316 ( .A1(n5620), .A2(n5619), .ZN(n4852) );
  NAND2_X1 U5317 ( .A1(n7178), .A2(n7180), .ZN(n7177) );
  XNOR2_X1 U5318 ( .A(n6258), .B(n7333), .ZN(n6885) );
  INV_X1 U5319 ( .A(n6885), .ZN(n8096) );
  AND2_X2 U5320 ( .A1(n5010), .A2(n5009), .ZN(n6268) );
  INV_X1 U5321 ( .A(n9577), .ZN(n9417) );
  NOR2_X1 U5322 ( .A1(n4876), .A2(n4875), .ZN(n5650) );
  INV_X1 U5323 ( .A(n4877), .ZN(n4875) );
  NOR2_X1 U5324 ( .A1(n9301), .A2(n4879), .ZN(n4876) );
  NAND2_X1 U5325 ( .A1(n5361), .A2(n5360), .ZN(n9480) );
  NAND2_X1 U5326 ( .A1(n5298), .A2(n5297), .ZN(n9497) );
  NAND2_X1 U5327 ( .A1(n6474), .A2(n5665), .ZN(n9500) );
  NAND2_X1 U5328 ( .A1(n5608), .A2(n5581), .ZN(n6478) );
  INV_X1 U5329 ( .A(n4905), .ZN(n4904) );
  XNOR2_X1 U5330 ( .A(n5506), .B(n5505), .ZN(n7709) );
  NAND2_X1 U5331 ( .A1(n4604), .A2(n4608), .ZN(n5515) );
  XNOR2_X1 U5332 ( .A(n5501), .B(n5500), .ZN(n7645) );
  OAI21_X1 U5333 ( .B1(n5485), .B2(n5484), .A(n5483), .ZN(n5501) );
  NAND2_X1 U5334 ( .A1(n4488), .A2(n5262), .ZN(n4481) );
  OAI21_X1 U5335 ( .B1(n4483), .B2(n5262), .A(n4478), .ZN(n4477) );
  NAND2_X1 U5336 ( .A1(n4487), .A2(n5226), .ZN(n5247) );
  OR2_X1 U5337 ( .A1(n5228), .A2(n5227), .ZN(n4487) );
  NAND2_X1 U5338 ( .A1(n4750), .A2(n4751), .ZN(n5207) );
  NAND2_X1 U5339 ( .A1(n5128), .A2(n4418), .ZN(n4747) );
  AND2_X1 U5340 ( .A1(n5151), .A2(n5138), .ZN(n5147) );
  AND2_X1 U5341 ( .A1(n5106), .A2(n5108), .ZN(n5129) );
  INV_X1 U5342 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5062) );
  INV_X1 U5343 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4850) );
  XNOR2_X1 U5344 ( .A(n5073), .B(n10127), .ZN(n5126) );
  NAND2_X1 U5345 ( .A1(n5018), .A2(n5017), .ZN(n5031) );
  INV_X1 U5346 ( .A(n8830), .ZN(n9025) );
  NAND2_X1 U5347 ( .A1(n6094), .A2(n6093), .ZN(n9045) );
  NAND2_X1 U5348 ( .A1(n5919), .A2(n5918), .ZN(n9924) );
  AND4_X1 U5349 ( .A1(n6030), .A2(n6029), .A3(n6028), .A4(n6027), .ZN(n8779)
         );
  INV_X1 U5350 ( .A(n8880), .ZN(n9040) );
  AND4_X1 U5351 ( .A1(n6012), .A2(n6011), .A3(n6010), .A4(n6009), .ZN(n8649)
         );
  AND4_X1 U5352 ( .A1(n5981), .A2(n5980), .A3(n5979), .A4(n5978), .ZN(n7896)
         );
  NAND2_X1 U5353 ( .A1(n5994), .A2(n5993), .ZN(n7901) );
  INV_X1 U5354 ( .A(n9865), .ZN(n8497) );
  NAND2_X1 U5355 ( .A1(n4572), .A2(n4571), .ZN(n4570) );
  NAND2_X1 U5356 ( .A1(n4573), .A2(n4738), .ZN(n4572) );
  OR2_X1 U5357 ( .A1(n8495), .A2(n8494), .ZN(n4571) );
  INV_X1 U5358 ( .A(n6727), .ZN(n9542) );
  AOI21_X1 U5359 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n6769), .A(n6764), .ZN(
        n6767) );
  NAND2_X1 U5360 ( .A1(n5974), .A2(n5973), .ZN(n9083) );
  AND2_X1 U5361 ( .A1(n4679), .A2(n4411), .ZN(n7087) );
  INV_X1 U5362 ( .A(n5026), .ZN(n6501) );
  NAND2_X1 U5363 ( .A1(n7932), .A2(n6353), .ZN(n7305) );
  AND3_X1 U5364 ( .A1(n5043), .A2(n5042), .A3(n5041), .ZN(n7258) );
  AND2_X1 U5365 ( .A1(n5523), .A2(n5493), .ZN(n9305) );
  NAND2_X1 U5366 ( .A1(n4473), .A2(n9349), .ZN(n4471) );
  INV_X1 U5367 ( .A(n4469), .ZN(n4468) );
  OAI21_X1 U5368 ( .B1(n4474), .B2(n4389), .A(n8251), .ZN(n4469) );
  OR2_X1 U5369 ( .A1(n5085), .A2(n5084), .ZN(n9231) );
  NAND2_X1 U5370 ( .A1(n6647), .A2(n6514), .ZN(n9631) );
  NAND2_X1 U5371 ( .A1(n7966), .A2(n7965), .ZN(n9426) );
  NAND2_X1 U5372 ( .A1(n5662), .A2(n5661), .ZN(n8088) );
  NAND2_X1 U5373 ( .A1(n4406), .A2(n4949), .ZN(n5613) );
  NAND2_X1 U5374 ( .A1(n5519), .A2(n5518), .ZN(n9434) );
  NAND2_X1 U5375 ( .A1(n4882), .A2(n4880), .ZN(n9283) );
  AND2_X1 U5376 ( .A1(n4882), .A2(n4881), .ZN(n9282) );
  OAI22_X1 U5377 ( .A1(n8189), .A2(n9577), .B1(n9312), .B2(n5559), .ZN(n4652)
         );
  INV_X1 U5378 ( .A(n4885), .ZN(n4883) );
  NAND2_X1 U5379 ( .A1(n4448), .A2(n4659), .ZN(n4658) );
  NAND2_X1 U5380 ( .A1(n9320), .A2(n9419), .ZN(n4659) );
  INV_X1 U5381 ( .A(n5653), .ZN(n8205) );
  NAND2_X1 U5382 ( .A1(n4403), .A2(n4492), .ZN(n4490) );
  AND2_X1 U5383 ( .A1(n8029), .A2(n8026), .ZN(n4491) );
  NOR2_X1 U5384 ( .A1(n8968), .A2(n4416), .ZN(n4741) );
  OAI21_X1 U5385 ( .B1(n8432), .B2(n4745), .A(n4686), .ZN(n4744) );
  NAND2_X1 U5386 ( .A1(n8326), .A2(n4746), .ZN(n4745) );
  INV_X1 U5387 ( .A(n8431), .ZN(n4746) );
  INV_X1 U5388 ( .A(n8040), .ZN(n4507) );
  NAND2_X1 U5389 ( .A1(n4742), .A2(n4740), .ZN(n8441) );
  OAI21_X1 U5390 ( .B1(n4744), .B2(n8434), .A(n4743), .ZN(n4742) );
  OAI21_X1 U5391 ( .B1(n4744), .B2(n4846), .A(n4741), .ZN(n4740) );
  AOI21_X1 U5392 ( .B1(n9079), .B2(n8649), .A(n4382), .ZN(n4743) );
  NAND2_X1 U5393 ( .A1(n4503), .A2(n4423), .ZN(n8159) );
  INV_X1 U5394 ( .A(n8013), .ZN(n4503) );
  AND2_X1 U5395 ( .A1(n8044), .A2(n8043), .ZN(n8170) );
  NOR3_X1 U5396 ( .A1(n8452), .A2(n8903), .A3(n8455), .ZN(n4727) );
  NAND2_X1 U5397 ( .A1(n8343), .A2(n4726), .ZN(n4725) );
  NAND2_X1 U5398 ( .A1(n8898), .A2(n8647), .ZN(n4726) );
  OAI21_X1 U5399 ( .B1(n8459), .B2(n8903), .A(n8458), .ZN(n4729) );
  AND2_X1 U5400 ( .A1(n8555), .A2(n4919), .ZN(n4918) );
  OR2_X1 U5401 ( .A1(n8604), .A2(n4920), .ZN(n4919) );
  INV_X1 U5402 ( .A(n6063), .ZN(n4920) );
  INV_X1 U5403 ( .A(n8410), .ZN(n4830) );
  INV_X1 U5404 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4720) );
  NAND2_X1 U5405 ( .A1(n4787), .A2(n4788), .ZN(n4785) );
  INV_X1 U5406 ( .A(n5215), .ZN(n4788) );
  AOI21_X1 U5407 ( .B1(n5215), .B2(n5180), .A(n6445), .ZN(n4787) );
  INV_X1 U5408 ( .A(n9181), .ZN(n4763) );
  AOI21_X1 U5409 ( .B1(n4498), .B2(n4495), .A(n4494), .ZN(n8076) );
  INV_X1 U5410 ( .A(n8070), .ZN(n4494) );
  NOR2_X1 U5411 ( .A1(n4497), .A2(n4496), .ZN(n4495) );
  INV_X1 U5412 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4960) );
  INV_X1 U5413 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n4961) );
  INV_X1 U5414 ( .A(n5531), .ZN(n4580) );
  NOR2_X1 U5415 ( .A1(n4584), .A2(n5659), .ZN(n4583) );
  INV_X1 U5416 ( .A(n5535), .ZN(n4584) );
  NOR2_X1 U5417 ( .A1(n4607), .A2(n4603), .ZN(n4602) );
  INV_X1 U5418 ( .A(n5465), .ZN(n4603) );
  INV_X1 U5419 ( .A(n4608), .ZN(n4607) );
  INV_X1 U5420 ( .A(n5483), .ZN(n4606) );
  OR2_X1 U5421 ( .A1(n5462), .A2(n5461), .ZN(n5466) );
  INV_X1 U5422 ( .A(n5446), .ZN(n4612) );
  INV_X1 U5423 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U5424 ( .A1(n4596), .A2(n5324), .ZN(n4589) );
  NOR2_X1 U5425 ( .A1(n4592), .A2(n5328), .ZN(n4591) );
  INV_X1 U5426 ( .A(n5262), .ZN(n4480) );
  NAND2_X1 U5427 ( .A1(n4578), .A2(n4577), .ZN(n4576) );
  NAND2_X1 U5428 ( .A1(n6553), .A2(n6579), .ZN(n4577) );
  OR2_X1 U5429 ( .A1(n6553), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n4578) );
  INV_X1 U5430 ( .A(n7478), .ZN(n4932) );
  OR2_X1 U5431 ( .A1(n5771), .A2(n6832), .ZN(n5750) );
  NAND2_X1 U5432 ( .A1(n4723), .A2(n4722), .ZN(n8463) );
  OR2_X1 U5433 ( .A1(n8492), .A2(n4382), .ZN(n4619) );
  INV_X1 U5434 ( .A(n8488), .ZN(n4739) );
  NAND2_X1 U5435 ( .A1(n9005), .A2(n8764), .ZN(n8489) );
  NOR2_X1 U5436 ( .A1(n8481), .A2(n4848), .ZN(n4847) );
  INV_X1 U5437 ( .A(n8287), .ZN(n4848) );
  AND2_X1 U5438 ( .A1(n8490), .A2(n8478), .ZN(n8485) );
  INV_X1 U5439 ( .A(n8848), .ZN(n8788) );
  NOR2_X1 U5440 ( .A1(n9025), .A2(n8817), .ZN(n8286) );
  INV_X1 U5441 ( .A(n8282), .ZN(n4836) );
  INV_X1 U5442 ( .A(n8451), .ZN(n4835) );
  INV_X1 U5443 ( .A(n4694), .ZN(n4692) );
  AND2_X1 U5444 ( .A1(n9062), .A2(n8781), .ZN(n8782) );
  INV_X1 U5445 ( .A(n6053), .ZN(n6054) );
  INV_X1 U5446 ( .A(n4828), .ZN(n4825) );
  INV_X1 U5447 ( .A(n4400), .ZN(n4707) );
  NOR2_X1 U5448 ( .A1(n4830), .A2(n4829), .ZN(n4828) );
  INV_X1 U5449 ( .A(n8406), .ZN(n4829) );
  OAI21_X1 U5450 ( .B1(n8405), .B2(n4830), .A(n4827), .ZN(n4826) );
  AND2_X1 U5451 ( .A1(n8397), .A2(n8406), .ZN(n8323) );
  NOR2_X1 U5452 ( .A1(n5893), .A2(n10187), .ZN(n5921) );
  AND2_X1 U5453 ( .A1(n9911), .A2(n7316), .ZN(n4625) );
  AND2_X1 U5454 ( .A1(n6950), .A2(n7089), .ZN(n4814) );
  AND2_X1 U5455 ( .A1(n6948), .A2(n8366), .ZN(n8313) );
  NAND2_X1 U5456 ( .A1(n8664), .A2(n9885), .ZN(n8315) );
  OR2_X1 U5457 ( .A1(n6923), .A2(n6828), .ZN(n7048) );
  NAND2_X1 U5458 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n9124), .ZN(n4721) );
  OR2_X1 U5459 ( .A1(n6181), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n6191) );
  INV_X1 U5460 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5686) );
  INV_X1 U5461 ( .A(n6391), .ZN(n4561) );
  OR2_X1 U5462 ( .A1(n4773), .A2(n6399), .ZN(n4769) );
  OR2_X1 U5463 ( .A1(n6404), .A2(n4772), .ZN(n4771) );
  INV_X1 U5464 ( .A(n7883), .ZN(n4772) );
  NAND2_X1 U5465 ( .A1(n4536), .A2(n4534), .ZN(n4542) );
  NOR2_X1 U5466 ( .A1(n4543), .A2(n4535), .ZN(n4534) );
  INV_X1 U5467 ( .A(n4759), .ZN(n4535) );
  OR2_X1 U5468 ( .A1(n6959), .A2(n6290), .ZN(n7253) );
  OR2_X1 U5469 ( .A1(n9685), .A2(n4808), .ZN(n4807) );
  AND2_X1 U5470 ( .A1(n9684), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4808) );
  NOR2_X1 U5471 ( .A1(n9346), .A2(n5571), .ZN(n9302) );
  NAND2_X1 U5472 ( .A1(n4677), .A2(n8256), .ZN(n4676) );
  NOR2_X1 U5473 ( .A1(n9465), .A2(n9471), .ZN(n4677) );
  NOR2_X1 U5474 ( .A1(n9497), .A2(n7778), .ZN(n4671) );
  AND2_X1 U5475 ( .A1(n4671), .A2(n4670), .ZN(n4669) );
  INV_X1 U5476 ( .A(n5300), .ZN(n5299) );
  NAND2_X1 U5477 ( .A1(n4861), .A2(n4865), .ZN(n9581) );
  NAND2_X1 U5478 ( .A1(n7403), .A2(n4399), .ZN(n4861) );
  NAND2_X1 U5479 ( .A1(n5054), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U5480 ( .A1(n5093), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5117) );
  INV_X1 U5481 ( .A(n5095), .ZN(n5093) );
  INV_X1 U5482 ( .A(n6249), .ZN(n6890) );
  OAI22_X1 U5483 ( .A1(n5077), .A2(n6530), .B1(n4631), .B2(n5539), .ZN(n5005)
         );
  INV_X1 U5484 ( .A(n4881), .ZN(n4879) );
  AOI21_X1 U5485 ( .B1(n4881), .B2(n4878), .A(n4431), .ZN(n4877) );
  INV_X1 U5486 ( .A(n4886), .ZN(n4878) );
  NAND2_X1 U5487 ( .A1(n7781), .A2(n7846), .ZN(n7860) );
  OR2_X1 U5488 ( .A1(n7220), .A2(n7192), .ZN(n7186) );
  NOR2_X1 U5489 ( .A1(n7205), .A2(n7209), .ZN(n7218) );
  NAND2_X1 U5490 ( .A1(n7333), .A2(n8210), .ZN(n7205) );
  NAND2_X1 U5491 ( .A1(n5485), .A2(n5483), .ZN(n4604) );
  AND2_X1 U5492 ( .A1(n4609), .A2(n5500), .ZN(n4608) );
  NAND2_X1 U5493 ( .A1(n5484), .A2(n5483), .ZN(n4609) );
  NAND2_X1 U5494 ( .A1(n4590), .A2(n4587), .ZN(n5349) );
  INV_X1 U5495 ( .A(n4588), .ZN(n4587) );
  NAND2_X1 U5496 ( .A1(n5288), .A2(n4591), .ZN(n4590) );
  OAI21_X1 U5497 ( .B1(n4592), .B2(n4589), .A(n5327), .ZN(n4588) );
  INV_X1 U5498 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5312) );
  INV_X1 U5499 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4956) );
  OR2_X1 U5500 ( .A1(n5248), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5295) );
  NAND2_X1 U5501 ( .A1(n5227), .A2(n5226), .ZN(n4489) );
  NAND2_X1 U5502 ( .A1(n5209), .A2(n10018), .ZN(n5226) );
  AOI21_X1 U5503 ( .B1(n5185), .B2(n4753), .A(n4752), .ZN(n4751) );
  INV_X1 U5504 ( .A(n5156), .ZN(n4753) );
  INV_X1 U5505 ( .A(n5187), .ZN(n4752) );
  INV_X1 U5506 ( .A(n5185), .ZN(n4754) );
  INV_X1 U5507 ( .A(n4913), .ZN(n4912) );
  OAI21_X1 U5508 ( .B1(n8561), .B2(n4914), .A(n8635), .ZN(n4913) );
  NAND2_X1 U5509 ( .A1(n7711), .A2(n4421), .ZN(n7832) );
  INV_X1 U5510 ( .A(n7835), .ZN(n5964) );
  INV_X1 U5511 ( .A(n6040), .ZN(n6041) );
  NAND2_X1 U5512 ( .A1(n6041), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6053) );
  AND2_X1 U5513 ( .A1(n8506), .A2(n5735), .ZN(n8547) );
  OR2_X1 U5514 ( .A1(n8507), .A2(n5747), .ZN(n5735) );
  NAND2_X1 U5515 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(n6054), .ZN(n6068) );
  AOI21_X1 U5516 ( .B1(n4928), .B2(n4930), .A(n4927), .ZN(n4926) );
  INV_X1 U5517 ( .A(n8620), .ZN(n4927) );
  NAND2_X1 U5518 ( .A1(n4933), .A2(n4932), .ZN(n7476) );
  NAND2_X1 U5519 ( .A1(n6066), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6082) );
  INV_X1 U5520 ( .A(n6068), .ZN(n6066) );
  INV_X1 U5521 ( .A(n6024), .ZN(n6025) );
  NAND2_X1 U5522 ( .A1(n4734), .A2(n4464), .ZN(n4573) );
  NAND2_X1 U5523 ( .A1(n4732), .A2(n4730), .ZN(n4734) );
  AND4_X1 U5524 ( .A1(n5828), .A2(n5827), .A3(n5826), .A4(n5825), .ZN(n6945)
         );
  NOR2_X1 U5525 ( .A1(n9540), .A2(n9539), .ZN(n9538) );
  AOI21_X1 U5526 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7451), .A(n7450), .ZN(
        n8668) );
  NOR2_X1 U5527 ( .A1(n7598), .A2(n4458), .ZN(n7602) );
  NAND2_X1 U5528 ( .A1(n7602), .A2(n7601), .ZN(n7654) );
  NAND2_X1 U5529 ( .A1(n7654), .A2(n4512), .ZN(n7656) );
  NAND2_X1 U5530 ( .A1(n7651), .A2(n7499), .ZN(n4512) );
  NAND2_X1 U5531 ( .A1(n7656), .A2(n7657), .ZN(n8680) );
  NAND2_X1 U5532 ( .A1(n8862), .A2(n4620), .ZN(n8800) );
  NOR2_X1 U5533 ( .A1(n8804), .A2(n4621), .ZN(n4620) );
  INV_X1 U5534 ( .A(n4622), .ZN(n4621) );
  NAND2_X1 U5535 ( .A1(n8295), .A2(n8294), .ZN(n8768) );
  AND2_X1 U5536 ( .A1(n8309), .A2(n8479), .ZN(n8797) );
  NAND2_X1 U5537 ( .A1(n8862), .A2(n4624), .ZN(n8825) );
  NOR2_X1 U5538 ( .A1(n8468), .A2(n8286), .ZN(n8833) );
  CLKBUF_X1 U5539 ( .A(n8832), .Z(n8847) );
  AND2_X1 U5540 ( .A1(n8467), .A2(n8834), .ZN(n8848) );
  INV_X1 U5541 ( .A(n6116), .ZN(n6100) );
  OR2_X1 U5542 ( .A1(n8896), .A2(n9040), .ZN(n8863) );
  AND2_X1 U5543 ( .A1(n8846), .A2(n8464), .ZN(n8871) );
  NAND2_X1 U5544 ( .A1(n4702), .A2(n4700), .ZN(n8861) );
  NAND2_X1 U5545 ( .A1(n4701), .A2(n4401), .ZN(n4700) );
  INV_X1 U5546 ( .A(n4703), .ZN(n4701) );
  OR2_X1 U5547 ( .A1(n8910), .A2(n9045), .ZN(n8896) );
  AND2_X1 U5548 ( .A1(n8980), .A2(n4626), .ZN(n8909) );
  NOR2_X1 U5549 ( .A1(n9057), .A2(n4628), .ZN(n4626) );
  NAND2_X1 U5550 ( .A1(n8909), .A2(n8916), .ZN(n8910) );
  INV_X1 U5551 ( .A(n4690), .ZN(n8926) );
  OAI21_X1 U5552 ( .B1(n8979), .B2(n4693), .A(n4691), .ZN(n4690) );
  NAND2_X1 U5553 ( .A1(n8940), .A2(n4697), .ZN(n4693) );
  AOI21_X1 U5554 ( .B1(n8940), .B2(n4692), .A(n8782), .ZN(n4691) );
  AND4_X1 U5555 ( .A1(n6045), .A2(n6044), .A3(n6043), .A4(n6042), .ZN(n8953)
         );
  AND2_X1 U5556 ( .A1(n8990), .A2(n8778), .ZN(n8968) );
  NAND2_X1 U5557 ( .A1(n8980), .A2(n4630), .ZN(n8961) );
  NAND2_X1 U5558 ( .A1(n4842), .A2(n4840), .ZN(n8992) );
  NAND2_X1 U5559 ( .A1(n4841), .A2(n4844), .ZN(n4840) );
  INV_X1 U5560 ( .A(n4845), .ZN(n4841) );
  NAND2_X1 U5561 ( .A1(n8980), .A2(n8990), .ZN(n8981) );
  NOR2_X1 U5562 ( .A1(n10210), .A2(n5986), .ZN(n6007) );
  AND2_X1 U5563 ( .A1(n9083), .A2(n8650), .ZN(n4687) );
  NOR2_X1 U5564 ( .A1(n7803), .A2(n9083), .ZN(n7814) );
  AND2_X1 U5565 ( .A1(n7814), .A2(n7816), .ZN(n8980) );
  OR2_X1 U5566 ( .A1(n7637), .A2(n7901), .ZN(n7803) );
  AND2_X1 U5567 ( .A1(n8420), .A2(n8421), .ZN(n8327) );
  AND4_X1 U5568 ( .A1(n5963), .A2(n5962), .A3(n5961), .A4(n5960), .ZN(n7898)
         );
  NAND2_X1 U5569 ( .A1(n7490), .A2(n8405), .ZN(n7492) );
  OR2_X1 U5570 ( .A1(n7375), .A2(n9924), .ZN(n7498) );
  NAND2_X1 U5571 ( .A1(n7372), .A2(n8406), .ZN(n7490) );
  AOI21_X1 U5572 ( .B1(n7282), .B2(n8319), .A(n4424), .ZN(n4688) );
  AND3_X1 U5573 ( .A1(n4394), .A2(n9917), .A3(n6952), .ZN(n7347) );
  AND4_X1 U5574 ( .A1(n5863), .A2(n5862), .A3(n5861), .A4(n5860), .ZN(n7482)
         );
  NAND2_X1 U5575 ( .A1(n6952), .A2(n4625), .ZN(n7360) );
  NAND2_X1 U5576 ( .A1(n6952), .A2(n7316), .ZN(n7097) );
  AND2_X1 U5577 ( .A1(n7089), .A2(n8379), .ZN(n8376) );
  NAND2_X1 U5578 ( .A1(n7265), .A2(n8374), .ZN(n4820) );
  NAND2_X1 U5579 ( .A1(n7264), .A2(n6950), .ZN(n4821) );
  OR2_X1 U5580 ( .A1(n5794), .A2(n5835), .ZN(n5837) );
  NOR2_X1 U5581 ( .A1(n7149), .A2(n8586), .ZN(n7271) );
  OR2_X1 U5582 ( .A1(n7147), .A2(n9897), .ZN(n7149) );
  OR2_X1 U5583 ( .A1(n6841), .A2(n8311), .ZN(n7156) );
  NOR2_X1 U5584 ( .A1(n7239), .A2(n7234), .ZN(n7236) );
  INV_X1 U5585 ( .A(n8314), .ZN(n8356) );
  NAND2_X1 U5586 ( .A1(n6833), .A2(n9872), .ZN(n7234) );
  NAND2_X1 U5587 ( .A1(n6180), .A2(n6179), .ZN(n9020) );
  NAND2_X1 U5588 ( .A1(n8945), .A2(n8453), .ZN(n8931) );
  NAND2_X1 U5589 ( .A1(n5934), .A2(n5933), .ZN(n9089) );
  INV_X1 U5590 ( .A(n9927), .ZN(n9899) );
  INV_X1 U5591 ( .A(n9925), .ZN(n9898) );
  NOR2_X2 U5592 ( .A1(n5774), .A2(n5778), .ZN(n9891) );
  NAND2_X1 U5593 ( .A1(n5777), .A2(n5776), .ZN(n5778) );
  NAND2_X1 U5594 ( .A1(n7797), .A2(n9103), .ZN(n9931) );
  AND3_X2 U5595 ( .A1(n5684), .A2(n4831), .A3(n4922), .ZN(n5706) );
  AND2_X1 U5596 ( .A1(n5683), .A2(n5731), .ZN(n4832) );
  INV_X1 U5597 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5713) );
  INV_X1 U5598 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5688) );
  INV_X1 U5599 ( .A(n5706), .ZN(n6181) );
  NAND2_X1 U5600 ( .A1(n4937), .A2(n4936), .ZN(n4935) );
  INV_X1 U5601 ( .A(n4938), .ZN(n4937) );
  AND2_X1 U5602 ( .A1(n5795), .A2(n5833), .ZN(n4923) );
  NAND2_X1 U5603 ( .A1(n6448), .A2(n6450), .ZN(n6451) );
  INV_X1 U5604 ( .A(n6449), .ZN(n6450) );
  INV_X1 U5605 ( .A(n4765), .ZN(n6350) );
  NAND2_X1 U5606 ( .A1(n5395), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U5607 ( .A1(n6331), .A2(n6330), .ZN(n7521) );
  NAND2_X1 U5608 ( .A1(n7756), .A2(n6391), .ZN(n7825) );
  NAND2_X1 U5609 ( .A1(n7825), .A2(n7826), .ZN(n7824) );
  OR2_X1 U5610 ( .A1(n5240), .A2(n5239), .ZN(n5255) );
  OR2_X1 U5611 ( .A1(n5173), .A2(n6811), .ZN(n5197) );
  AND2_X1 U5612 ( .A1(n6377), .A2(n6372), .ZN(n6373) );
  AND2_X1 U5613 ( .A1(n8126), .A2(n8125), .ZN(n8128) );
  OR3_X1 U5614 ( .A1(n8208), .A2(n8241), .A3(n8124), .ZN(n8126) );
  AND3_X1 U5615 ( .A1(n5224), .A2(n5223), .A3(n5222), .ZN(n7551) );
  AND2_X1 U5616 ( .A1(n5169), .A2(n5168), .ZN(n7935) );
  AND3_X1 U5617 ( .A1(n5123), .A2(n5122), .A3(n5121), .ZN(n6309) );
  NOR2_X1 U5618 ( .A1(n6703), .A2(n6702), .ZN(n6701) );
  AND2_X1 U5619 ( .A1(n4798), .A2(n4797), .ZN(n6872) );
  NAND2_X1 U5620 ( .A1(n6871), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4797) );
  NAND2_X1 U5621 ( .A1(n6872), .A2(n6873), .ZN(n9237) );
  NOR2_X1 U5622 ( .A1(n9670), .A2(n4809), .ZN(n9686) );
  AND2_X1 U5623 ( .A1(n9675), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4809) );
  NOR2_X1 U5624 ( .A1(n9686), .A2(n9687), .ZN(n9685) );
  XNOR2_X1 U5625 ( .A(n4807), .B(n9699), .ZN(n9701) );
  NOR2_X1 U5626 ( .A1(n9735), .A2(n4796), .ZN(n9754) );
  AND2_X1 U5627 ( .A1(n9739), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4796) );
  NOR2_X1 U5628 ( .A1(n9754), .A2(n9755), .ZN(n9756) );
  XNOR2_X1 U5629 ( .A(n4794), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9270) );
  OR2_X1 U5630 ( .A1(n9756), .A2(n4795), .ZN(n4794) );
  AND2_X1 U5631 ( .A1(n9752), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4795) );
  NOR2_X1 U5632 ( .A1(n4884), .A2(n9288), .ZN(n4881) );
  INV_X1 U5633 ( .A(n4884), .ZN(n4880) );
  AND2_X1 U5634 ( .A1(n8129), .A2(n8184), .ZN(n9288) );
  NAND2_X1 U5635 ( .A1(n9307), .A2(n9135), .ZN(n4885) );
  INV_X1 U5636 ( .A(n7950), .ZN(n9286) );
  AND2_X1 U5637 ( .A1(n8181), .A2(n8186), .ZN(n9309) );
  NAND2_X1 U5638 ( .A1(n5452), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5475) );
  INV_X1 U5639 ( .A(n5453), .ZN(n5452) );
  NAND2_X1 U5640 ( .A1(n4891), .A2(n4890), .ZN(n9324) );
  NAND2_X1 U5641 ( .A1(n4393), .A2(n4901), .ZN(n4890) );
  AND2_X1 U5642 ( .A1(n8180), .A2(n8061), .ZN(n9323) );
  NAND2_X1 U5643 ( .A1(n8258), .A2(n8173), .ZN(n9337) );
  NAND2_X1 U5644 ( .A1(n8258), .A2(n4639), .ZN(n9339) );
  NOR2_X1 U5645 ( .A1(n9372), .A2(n4675), .ZN(n8267) );
  INV_X1 U5646 ( .A(n4677), .ZN(n4675) );
  INV_X1 U5647 ( .A(n4647), .ZN(n4646) );
  AND2_X1 U5648 ( .A1(n5405), .A2(n4644), .ZN(n4643) );
  NAND2_X1 U5649 ( .A1(n4647), .A2(n4645), .ZN(n4644) );
  NOR2_X1 U5650 ( .A1(n9372), .A2(n9471), .ZN(n9357) );
  INV_X1 U5651 ( .A(n4856), .ZN(n4855) );
  AOI21_X1 U5652 ( .B1(n4856), .B2(n4854), .A(n4451), .ZN(n4853) );
  AND2_X1 U5653 ( .A1(n4857), .A2(n5641), .ZN(n4856) );
  AND2_X1 U5654 ( .A1(n7781), .A2(n4667), .ZN(n9406) );
  NOR2_X1 U5655 ( .A1(n9486), .A2(n4668), .ZN(n4667) );
  INV_X1 U5656 ( .A(n4669), .ZN(n4668) );
  NAND2_X1 U5657 ( .A1(n7781), .A2(n4671), .ZN(n7868) );
  AOI21_X1 U5658 ( .B1(n4862), .B2(n4864), .A(n4429), .ZN(n4860) );
  NAND2_X1 U5659 ( .A1(n5216), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5240) );
  INV_X1 U5660 ( .A(n5217), .ZN(n5216) );
  NAND2_X1 U5661 ( .A1(n5195), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5217) );
  INV_X1 U5662 ( .A(n5197), .ZN(n5195) );
  NAND2_X1 U5663 ( .A1(n7569), .A2(n9507), .ZN(n9592) );
  INV_X1 U5664 ( .A(n4642), .ZN(n4641) );
  AND2_X1 U5665 ( .A1(n7999), .A2(n7984), .ZN(n8101) );
  AND2_X1 U5666 ( .A1(n7433), .A2(n4665), .ZN(n7569) );
  AND2_X1 U5667 ( .A1(n4392), .A2(n9564), .ZN(n4665) );
  OR2_X1 U5668 ( .A1(n8101), .A2(n7561), .ZN(n7564) );
  NAND2_X1 U5669 ( .A1(n5116), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5171) );
  INV_X1 U5670 ( .A(n5117), .ZN(n5116) );
  OR2_X1 U5671 ( .A1(n5171), .A2(n5170), .ZN(n5173) );
  NAND2_X1 U5672 ( .A1(n7398), .A2(n5146), .ZN(n7557) );
  NAND2_X1 U5673 ( .A1(n7433), .A2(n4386), .ZN(n7625) );
  AND2_X1 U5674 ( .A1(n7982), .A2(n7993), .ZN(n8099) );
  NAND2_X1 U5675 ( .A1(n7433), .A2(n9819), .ZN(n7406) );
  NAND2_X1 U5676 ( .A1(n4446), .A2(n5115), .ZN(n7398) );
  OAI211_X1 U5677 ( .C1(n5026), .C2(n6662), .A(n5076), .B(n5075), .ZN(n7437)
         );
  OR2_X1 U5678 ( .A1(n5180), .A2(n5835), .ZN(n5075) );
  AND2_X1 U5679 ( .A1(n7019), .A2(n5621), .ZN(n7432) );
  AND3_X1 U5680 ( .A1(n5060), .A2(n5059), .A3(n5058), .ZN(n7022) );
  NAND2_X1 U5681 ( .A1(n8140), .A2(n8138), .ZN(n8090) );
  INV_X1 U5682 ( .A(n5615), .ZN(n8092) );
  AND3_X1 U5683 ( .A1(n5025), .A2(n5024), .A3(n5023), .ZN(n7201) );
  NAND2_X1 U5684 ( .A1(n5491), .A2(n5490), .ZN(n9443) );
  INV_X1 U5685 ( .A(n7437), .ZN(n9812) );
  AND2_X1 U5686 ( .A1(n4636), .A2(n4633), .ZN(n4979) );
  NOR2_X1 U5687 ( .A1(n4634), .A2(n4968), .ZN(n4633) );
  XNOR2_X1 U5688 ( .A(n7954), .B(SI_30_), .ZN(n8293) );
  XNOR2_X1 U5689 ( .A(n5660), .B(n5536), .ZN(n8288) );
  NAND2_X1 U5690 ( .A1(n4585), .A2(n5535), .ZN(n5660) );
  NAND2_X1 U5691 ( .A1(n5532), .A2(n5531), .ZN(n4585) );
  XNOR2_X1 U5692 ( .A(n5532), .B(n5531), .ZN(n7789) );
  INV_X1 U5693 ( .A(n4907), .ZN(n4906) );
  INV_X1 U5694 ( .A(n5409), .ZN(n4615) );
  INV_X1 U5695 ( .A(n4614), .ZN(n4613) );
  OAI21_X1 U5696 ( .B1(n4617), .B2(n4445), .A(n5425), .ZN(n4614) );
  NAND2_X1 U5697 ( .A1(n4553), .A2(n4550), .ZN(n4549) );
  NOR2_X1 U5698 ( .A1(n4552), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n4548) );
  NAND2_X1 U5699 ( .A1(n4616), .A2(n5409), .ZN(n5427) );
  OAI21_X1 U5700 ( .B1(n5288), .B2(n4596), .A(n4593), .ZN(n5329) );
  OAI21_X1 U5701 ( .B1(n5288), .B2(n5287), .A(n5286), .ZN(n5309) );
  OR2_X1 U5702 ( .A1(n5234), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U5703 ( .A1(n5157), .A2(n5156), .ZN(n5186) );
  NAND2_X1 U5704 ( .A1(n5156), .A2(n5154), .ZN(n5178) );
  NAND2_X1 U5705 ( .A1(n4466), .A2(n5151), .ZN(n5179) );
  NAND2_X1 U5706 ( .A1(n4747), .A2(n4422), .ZN(n4466) );
  AND2_X1 U5707 ( .A1(n5148), .A2(n5147), .ZN(n5149) );
  OR2_X1 U5708 ( .A1(n5110), .A2(n5109), .ZN(n5125) );
  XNOR2_X1 U5709 ( .A(n5132), .B(SI_7_), .ZN(n5124) );
  NAND2_X1 U5710 ( .A1(n5048), .A2(n5047), .ZN(n5071) );
  XNOR2_X1 U5711 ( .A(n5016), .B(n4990), .ZN(n5015) );
  AND2_X1 U5712 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4989) );
  AND4_X1 U5713 ( .A1(n6147), .A2(n6146), .A3(n6145), .A4(n6144), .ZN(n8837)
         );
  AND4_X1 U5714 ( .A1(n5990), .A2(n5989), .A3(n5988), .A4(n5987), .ZN(n8576)
         );
  NAND2_X1 U5715 ( .A1(n7711), .A2(n5947), .ZN(n7834) );
  NAND2_X1 U5716 ( .A1(n5955), .A2(n5954), .ZN(n7841) );
  AND4_X1 U5717 ( .A1(n6088), .A2(n6087), .A3(n6086), .A4(n6085), .ZN(n8786)
         );
  NAND2_X1 U5718 ( .A1(n7476), .A2(n5889), .ZN(n7608) );
  NAND2_X1 U5719 ( .A1(n6920), .A2(n5765), .ZN(n7070) );
  OR2_X1 U5720 ( .A1(n5766), .A2(n5754), .ZN(n5756) );
  NAND2_X1 U5721 ( .A1(n6038), .A2(n6037), .ZN(n9068) );
  NAND2_X1 U5722 ( .A1(n8603), .A2(n8604), .ZN(n4917) );
  AND4_X1 U5723 ( .A1(n5941), .A2(n5940), .A3(n5939), .A4(n5938), .ZN(n7838)
         );
  NAND2_X1 U5724 ( .A1(n6123), .A2(n6122), .ZN(n8560) );
  NAND2_X1 U5725 ( .A1(n6125), .A2(n6124), .ZN(n9037) );
  NAND2_X1 U5726 ( .A1(n6003), .A2(n6002), .ZN(n6507) );
  OR2_X1 U5727 ( .A1(n5736), .A2(n5693), .ZN(n5697) );
  AND4_X1 U5728 ( .A1(n5926), .A2(n5925), .A3(n5924), .A4(n5923), .ZN(n7715)
         );
  AND4_X1 U5729 ( .A1(n6073), .A2(n6072), .A3(n6071), .A4(n6070), .ZN(n8951)
         );
  NAND2_X1 U5730 ( .A1(n4925), .A2(n4928), .ZN(n8621) );
  OR2_X1 U5731 ( .A1(n4933), .A2(n4930), .ZN(n4925) );
  NAND2_X1 U5732 ( .A1(n6504), .A2(n6019), .ZN(n7915) );
  AND2_X1 U5733 ( .A1(n6242), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8627) );
  NAND2_X1 U5734 ( .A1(n4911), .A2(n6138), .ZN(n8634) );
  NAND2_X1 U5735 ( .A1(n8560), .A2(n8561), .ZN(n4911) );
  INV_X1 U5736 ( .A(n6945), .ZN(n8660) );
  OAI211_X1 U5737 ( .C1(n5810), .C2(n6606), .A(n5812), .B(n4434), .ZN(n8661)
         );
  AND2_X1 U5738 ( .A1(n5769), .A2(n5770), .ZN(n4849) );
  INV_X1 U5739 ( .A(n4953), .ZN(n8664) );
  OR2_X1 U5740 ( .A1(n5766), .A2(n7117), .ZN(n5739) );
  INV_X1 U5741 ( .A(P2_U3966), .ZN(n8665) );
  NOR2_X1 U5742 ( .A1(n9550), .A2(n4943), .ZN(n6742) );
  INV_X1 U5743 ( .A(n4531), .ZN(n6778) );
  AND2_X1 U5744 ( .A1(n4531), .A2(n4530), .ZN(n6796) );
  NAND2_X1 U5745 ( .A1(n6779), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4530) );
  INV_X1 U5746 ( .A(n4529), .ZN(n6794) );
  AND2_X1 U5747 ( .A1(n4529), .A2(n4528), .ZN(n6781) );
  NAND2_X1 U5748 ( .A1(n6783), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4528) );
  NOR2_X1 U5749 ( .A1(n6903), .A2(n4527), .ZN(n6907) );
  AND2_X1 U5750 ( .A1(n6904), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4527) );
  NOR2_X1 U5751 ( .A1(n6907), .A2(n6906), .ZN(n6983) );
  NOR2_X1 U5752 ( .A1(n6983), .A2(n4526), .ZN(n6987) );
  AND2_X1 U5753 ( .A1(n6984), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4526) );
  NOR2_X1 U5754 ( .A1(n6987), .A2(n6986), .ZN(n7450) );
  AND2_X1 U5755 ( .A1(n4524), .A2(n4523), .ZN(n8728) );
  NAND2_X1 U5756 ( .A1(n4516), .A2(n4515), .ZN(n4514) );
  NAND2_X1 U5757 ( .A1(n4519), .A2(n6039), .ZN(n4516) );
  NAND2_X1 U5758 ( .A1(n8759), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n4515) );
  AOI22_X1 U5759 ( .A1(n4519), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n6039), .B2(
        n8759), .ZN(n4518) );
  AOI22_X1 U5760 ( .A1(n4519), .A2(n9549), .B1(n8759), .B2(n9549), .ZN(n4517)
         );
  AND2_X1 U5761 ( .A1(n6154), .A2(n6153), .ZN(n8830) );
  NAND2_X1 U5762 ( .A1(n7645), .A2(n8299), .ZN(n6140) );
  NAND2_X1 U5763 ( .A1(n8890), .A2(n8458), .ZN(n8882) );
  AND2_X1 U5764 ( .A1(n6097), .A2(n6096), .ZN(n8880) );
  NAND2_X1 U5765 ( .A1(n9047), .A2(n4704), .ZN(n8876) );
  NAND2_X1 U5766 ( .A1(n8904), .A2(n8903), .ZN(n9047) );
  INV_X1 U5767 ( .A(n9052), .ZN(n8916) );
  OAI21_X1 U5768 ( .B1(n8979), .B2(n4696), .A(n4694), .ZN(n8941) );
  AND2_X1 U5769 ( .A1(n4698), .A2(n4412), .ZN(n8960) );
  NAND2_X1 U5770 ( .A1(n8979), .A2(n8780), .ZN(n4698) );
  NAND2_X1 U5771 ( .A1(n7810), .A2(n8435), .ZN(n7811) );
  NAND2_X1 U5772 ( .A1(n7794), .A2(n7793), .ZN(n7795) );
  NAND2_X1 U5773 ( .A1(n4710), .A2(n4709), .ZN(n7534) );
  NAND2_X1 U5774 ( .A1(n4710), .A2(n4712), .ZN(n7488) );
  INV_X1 U5775 ( .A(n9094), .ZN(n7369) );
  NAND2_X1 U5776 ( .A1(n7283), .A2(n7282), .ZN(n7342) );
  NAND2_X1 U5777 ( .A1(n4819), .A2(n4818), .ZN(n7090) );
  AND3_X1 U5778 ( .A1(n5809), .A2(n5808), .A3(n5807), .ZN(n7325) );
  INV_X1 U5779 ( .A(n6833), .ZN(n8550) );
  AND2_X1 U5780 ( .A1(n8936), .A2(n7059), .ZN(n8845) );
  INV_X1 U5781 ( .A(n5694), .ZN(n7929) );
  INV_X1 U5782 ( .A(n5864), .ZN(n4833) );
  CLKBUF_X1 U5783 ( .A(n6215), .Z(n6216) );
  NOR2_X1 U5784 ( .A1(n5916), .A2(n4940), .ZN(n5971) );
  NAND2_X1 U5785 ( .A1(n5743), .A2(n5744), .ZN(n6727) );
  NAND2_X1 U5786 ( .A1(n9203), .A2(n6451), .ZN(n9133) );
  NAND2_X1 U5787 ( .A1(n5252), .A2(n5251), .ZN(n7751) );
  NAND2_X1 U5788 ( .A1(n5433), .A2(n5432), .ZN(n9460) );
  NAND2_X1 U5789 ( .A1(n6274), .A2(n6273), .ZN(n6972) );
  AND3_X1 U5790 ( .A1(n5345), .A2(n5344), .A3(n5343), .ZN(n7909) );
  OAI21_X1 U5791 ( .B1(n7756), .B2(n4562), .A(n4558), .ZN(n7905) );
  NAND2_X1 U5792 ( .A1(n4775), .A2(n4427), .ZN(n6493) );
  NAND2_X1 U5793 ( .A1(n6490), .A2(n6489), .ZN(n6491) );
  NAND2_X1 U5794 ( .A1(n9177), .A2(n9181), .ZN(n9155) );
  AND3_X1 U5795 ( .A1(n5307), .A2(n5306), .A3(n5305), .ZN(n7876) );
  NAND2_X1 U5796 ( .A1(n5377), .A2(n5376), .ZN(n9476) );
  CLKBUF_X1 U5797 ( .A(n9199), .Z(n9188) );
  OR2_X1 U5798 ( .A1(n6352), .A2(n6342), .ZN(n6344) );
  NAND2_X1 U5799 ( .A1(n5237), .A2(n5236), .ZN(n9501) );
  INV_X1 U5800 ( .A(n9218), .ZN(n9340) );
  NAND2_X1 U5801 ( .A1(n9178), .A2(n4540), .ZN(n4533) );
  NAND2_X1 U5802 ( .A1(n7885), .A2(n7883), .ZN(n7882) );
  AND3_X1 U5803 ( .A1(n5101), .A2(n5100), .A3(n5099), .ZN(n7427) );
  AND2_X1 U5804 ( .A1(n5481), .A2(n5480), .ZN(n9341) );
  NAND2_X1 U5805 ( .A1(n5499), .A2(n5498), .ZN(n9320) );
  INV_X1 U5806 ( .A(n9381), .ZN(n9219) );
  OR2_X1 U5807 ( .A1(n5387), .A2(n5386), .ZN(n9396) );
  OR2_X1 U5808 ( .A1(n5285), .A2(n5284), .ZN(n9221) );
  OR2_X1 U5809 ( .A1(n5258), .A2(n5257), .ZN(n9222) );
  INV_X1 U5810 ( .A(n6309), .ZN(n9228) );
  NAND2_X1 U5811 ( .A1(n4874), .A2(n4868), .ZN(n6258) );
  NAND2_X1 U5812 ( .A1(n5039), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4874) );
  AND3_X1 U5813 ( .A1(n4872), .A2(n4873), .A3(n4869), .ZN(n4868) );
  OR2_X1 U5814 ( .A1(n5539), .A2(n7126), .ZN(n4997) );
  NAND2_X1 U5815 ( .A1(n6515), .A2(n6516), .ZN(n9634) );
  INV_X1 U5816 ( .A(n4811), .ZN(n6635) );
  NAND2_X1 U5817 ( .A1(n4813), .A2(n4811), .ZN(n6637) );
  INV_X1 U5818 ( .A(n6634), .ZN(n4813) );
  NOR2_X1 U5819 ( .A1(n6701), .A2(n4805), .ZN(n9645) );
  OAI21_X1 U5820 ( .B1(n4801), .B2(n4805), .A(n4802), .ZN(n4804) );
  NAND2_X1 U5821 ( .A1(n4806), .A2(n4803), .ZN(n4800) );
  INV_X1 U5822 ( .A(n4798), .ZN(n6870) );
  INV_X1 U5823 ( .A(n4792), .ZN(n9712) );
  INV_X1 U5824 ( .A(n9243), .ZN(n4791) );
  NOR2_X1 U5825 ( .A1(n5357), .A2(n4565), .ZN(n4564) );
  OR2_X1 U5826 ( .A1(n9432), .A2(n9425), .ZN(n5655) );
  AOI21_X1 U5827 ( .B1(n9439), .B2(n9401), .A(n7953), .ZN(n4655) );
  NAND2_X1 U5828 ( .A1(n4893), .A2(n4895), .ZN(n9335) );
  NAND2_X1 U5829 ( .A1(n8266), .A2(n4899), .ZN(n4893) );
  NAND2_X1 U5830 ( .A1(n5451), .A2(n5450), .ZN(n9344) );
  INV_X1 U5831 ( .A(n9460), .ZN(n8256) );
  NAND2_X1 U5832 ( .A1(n4894), .A2(n4902), .ZN(n8253) );
  OR2_X1 U5833 ( .A1(n8266), .A2(n5646), .ZN(n4894) );
  NAND2_X1 U5834 ( .A1(n4649), .A2(n8165), .ZN(n9378) );
  NAND2_X1 U5835 ( .A1(n9404), .A2(n5640), .ZN(n9387) );
  INV_X1 U5836 ( .A(n9590), .ZN(n9410) );
  NAND2_X1 U5837 ( .A1(n4786), .A2(n5215), .ZN(n9593) );
  INV_X1 U5838 ( .A(n5627), .ZN(n4866) );
  NAND2_X1 U5839 ( .A1(n7403), .A2(n5628), .ZN(n4867) );
  NAND2_X1 U5840 ( .A1(n5194), .A2(n5193), .ZN(n7516) );
  NAND2_X1 U5841 ( .A1(n7177), .A2(n5619), .ZN(n7017) );
  NAND2_X1 U5842 ( .A1(n9837), .A2(n5586), .ZN(n9776) );
  AND2_X1 U5843 ( .A1(n9785), .A2(n9772), .ZN(n9590) );
  NOR2_X1 U5844 ( .A1(n5673), .A2(n5672), .ZN(n9603) );
  NAND2_X1 U5845 ( .A1(n5671), .A2(n9428), .ZN(n5672) );
  NAND2_X1 U5846 ( .A1(n8088), .A2(n9500), .ZN(n5671) );
  NOR2_X1 U5847 ( .A1(n9430), .A2(n4663), .ZN(n4662) );
  OAI21_X1 U5848 ( .B1(n9432), .B2(n9505), .A(n4664), .ZN(n4663) );
  NAND2_X1 U5849 ( .A1(n9431), .A2(n9500), .ZN(n4664) );
  NAND2_X1 U5850 ( .A1(n9436), .A2(n4650), .ZN(n9516) );
  INV_X1 U5851 ( .A(n4651), .ZN(n4650) );
  OAI21_X1 U5852 ( .B1(n9437), .B2(n9505), .A(n9435), .ZN(n4651) );
  INV_X1 U5853 ( .A(n4657), .ZN(n9441) );
  XNOR2_X1 U5854 ( .A(n7962), .B(n7961), .ZN(n8298) );
  INV_X1 U5855 ( .A(n4982), .ZN(n7919) );
  XNOR2_X1 U5856 ( .A(n5447), .B(n5446), .ZN(n7298) );
  OAI21_X1 U5857 ( .B1(n5392), .B2(n4445), .A(n4613), .ZN(n5447) );
  INV_X1 U5858 ( .A(n5652), .ZN(n8125) );
  INV_X1 U5859 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10115) );
  AND2_X1 U5860 ( .A1(n4747), .A2(n5131), .ZN(n5150) );
  INV_X1 U5861 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6561) );
  XNOR2_X1 U5862 ( .A(n4810), .B(n4991), .ZN(n6650) );
  NAND2_X1 U5863 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4810) );
  AND2_X1 U5864 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7705) );
  NAND2_X1 U5865 ( .A1(n4570), .A2(n8496), .ZN(n8503) );
  NAND2_X1 U5866 ( .A1(n8247), .A2(n4473), .ZN(n4472) );
  NAND2_X1 U5867 ( .A1(n4656), .A2(n4653), .ZN(P1_U3264) );
  INV_X1 U5868 ( .A(n4654), .ZN(n4653) );
  NAND2_X1 U5869 ( .A1(n4657), .A2(n9785), .ZN(n4656) );
  OAI21_X1 U5870 ( .B1(n9442), .B2(n9425), .A(n4655), .ZN(n4654) );
  AND2_X1 U5871 ( .A1(n8342), .A2(n8341), .ZN(n4385) );
  INV_X1 U5872 ( .A(n5611), .ZN(n5651) );
  INV_X1 U5873 ( .A(n4870), .ZN(n5040) );
  AND2_X1 U5874 ( .A1(n8394), .A2(n8391), .ZN(n8319) );
  INV_X1 U5875 ( .A(n6267), .ZN(n6328) );
  INV_X2 U5876 ( .A(n6328), .ZN(n6457) );
  INV_X1 U5877 ( .A(n6428), .ZN(n4758) );
  AND2_X1 U5878 ( .A1(n9819), .A2(n9823), .ZN(n4386) );
  AND2_X1 U5879 ( .A1(n4751), .A2(n5204), .ZN(n4387) );
  INV_X1 U5880 ( .A(n9179), .ZN(n4539) );
  OR2_X1 U5881 ( .A1(n7516), .A2(n9225), .ZN(n4388) );
  OR2_X1 U5882 ( .A1(n8201), .A2(n9349), .ZN(n4389) );
  INV_X1 U5883 ( .A(n9057), .ZN(n8928) );
  NAND2_X1 U5884 ( .A1(n6065), .A2(n6064), .ZN(n9057) );
  AND2_X1 U5885 ( .A1(n8153), .A2(n5115), .ZN(n4390) );
  AND2_X1 U5886 ( .A1(n5062), .A2(n5140), .ZN(n4391) );
  AND2_X1 U5887 ( .A1(n4386), .A2(n4666), .ZN(n4392) );
  NAND2_X1 U5888 ( .A1(n4443), .A2(n4895), .ZN(n4393) );
  AND2_X1 U5889 ( .A1(n4625), .A2(n7363), .ZN(n4394) );
  AND3_X1 U5890 ( .A1(n4833), .A2(n5684), .A3(n5683), .ZN(n4395) );
  XNOR2_X1 U5891 ( .A(n5552), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5652) );
  INV_X2 U5892 ( .A(n5736), .ZN(n5783) );
  NAND2_X1 U5893 ( .A1(n5472), .A2(n5471), .ZN(n5571) );
  AND2_X1 U5894 ( .A1(n8862), .A2(n4622), .ZN(n4396) );
  AND2_X1 U5895 ( .A1(n4649), .A2(n4647), .ZN(n4397) );
  OR2_X1 U5896 ( .A1(n5582), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4398) );
  AND2_X1 U5897 ( .A1(n5628), .A2(n4388), .ZN(n4399) );
  AND2_X1 U5898 ( .A1(n4711), .A2(n7370), .ZN(n4400) );
  OR2_X1 U5899 ( .A1(n9040), .A2(n8893), .ZN(n4401) );
  AND2_X1 U5900 ( .A1(n4597), .A2(n5308), .ZN(n4402) );
  INV_X1 U5901 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5970) );
  OR2_X1 U5902 ( .A1(n8021), .A2(n8020), .ZN(n4403) );
  OR3_X1 U5903 ( .A1(n8484), .A2(n8483), .A3(n8482), .ZN(n4404) );
  OR2_X1 U5904 ( .A1(n5142), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n4405) );
  INV_X1 U5905 ( .A(n8165), .ZN(n4648) );
  AND2_X1 U5906 ( .A1(n5570), .A2(n5569), .ZN(n4406) );
  NAND2_X1 U5907 ( .A1(n5145), .A2(n5144), .ZN(n7410) );
  OR2_X1 U5908 ( .A1(n4764), .A2(n6428), .ZN(n4407) );
  INV_X1 U5909 ( .A(n5134), .ZN(n5741) );
  NAND2_X1 U5910 ( .A1(n5277), .A2(n5276), .ZN(n7778) );
  NAND2_X1 U5911 ( .A1(n5026), .A2(n6553), .ZN(n5180) );
  INV_X1 U5912 ( .A(n9156), .ZN(n4764) );
  MUX2_X1 U5913 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9129), .S(n5773), .Z(n8507) );
  OR3_X1 U5914 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4408) );
  NOR2_X1 U5915 ( .A1(n5582), .A2(n4903), .ZN(n4409) );
  NAND2_X1 U5916 ( .A1(n4924), .A2(n4923), .ZN(n5841) );
  AND4_X1 U5917 ( .A1(n5720), .A2(n4936), .A3(n5721), .A4(n5678), .ZN(n4410)
         );
  NAND2_X1 U5918 ( .A1(n7269), .A2(n7316), .ZN(n4411) );
  NAND2_X1 U5919 ( .A1(n8990), .A2(n8779), .ZN(n4412) );
  NAND2_X1 U5920 ( .A1(n8971), .A2(n8282), .ZN(n8945) );
  INV_X1 U5921 ( .A(n7491), .ZN(n4827) );
  NAND2_X1 U5922 ( .A1(n5102), .A2(n5140), .ZN(n5142) );
  AND2_X1 U5923 ( .A1(n8284), .A2(n8458), .ZN(n4413) );
  NAND2_X1 U5924 ( .A1(n4955), .A2(n5011), .ZN(n5044) );
  AND2_X1 U5925 ( .A1(n7516), .A2(n9225), .ZN(n4414) );
  AND2_X1 U5926 ( .A1(n8196), .A2(n8192), .ZN(n4415) );
  OR2_X1 U5927 ( .A1(n8437), .A2(n4385), .ZN(n4416) );
  INV_X1 U5928 ( .A(n9465), .ZN(n8270) );
  NAND2_X1 U5929 ( .A1(n5417), .A2(n5416), .ZN(n9465) );
  AND2_X1 U5930 ( .A1(n5655), .A2(n5654), .ZN(n4417) );
  AND2_X1 U5931 ( .A1(n5127), .A2(n5126), .ZN(n4418) );
  XNOR2_X1 U5932 ( .A(n5205), .B(SI_11_), .ZN(n5204) );
  AND3_X1 U5933 ( .A1(n4994), .A2(n4992), .A3(n4993), .ZN(n7333) );
  INV_X1 U5934 ( .A(n9072), .ZN(n8990) );
  NAND2_X1 U5935 ( .A1(n6022), .A2(n6021), .ZN(n9072) );
  AND2_X1 U5936 ( .A1(n4792), .A2(n4791), .ZN(n4419) );
  AND2_X1 U5937 ( .A1(n4504), .A2(n4502), .ZN(n4420) );
  AND2_X1 U5938 ( .A1(n5964), .A2(n5947), .ZN(n4421) );
  AND2_X1 U5939 ( .A1(n5131), .A2(n5149), .ZN(n4422) );
  NAND2_X1 U5940 ( .A1(n8008), .A2(n8007), .ZN(n4423) );
  AND2_X1 U5941 ( .A1(n7341), .A2(n8656), .ZN(n4424) );
  INV_X1 U5942 ( .A(n4705), .ZN(n4704) );
  AND2_X1 U5943 ( .A1(n9089), .A2(n8653), .ZN(n4425) );
  AND2_X1 U5944 ( .A1(n9047), .A2(n4703), .ZN(n4426) );
  INV_X1 U5945 ( .A(n4770), .ZN(n7884) );
  NOR2_X1 U5946 ( .A1(n4774), .A2(n6404), .ZN(n4770) );
  NAND2_X1 U5947 ( .A1(n6140), .A2(n6139), .ZN(n9031) );
  AND2_X1 U5948 ( .A1(n4778), .A2(n6455), .ZN(n4427) );
  INV_X1 U5949 ( .A(n4697), .ZN(n4696) );
  AND2_X1 U5950 ( .A1(n4699), .A2(n4412), .ZN(n4697) );
  NOR2_X1 U5951 ( .A1(n8966), .A2(n8953), .ZN(n4428) );
  NOR2_X1 U5952 ( .A1(n5632), .A2(n5631), .ZN(n4429) );
  OR2_X1 U5953 ( .A1(n5627), .A2(n4414), .ZN(n4430) );
  AND2_X1 U5954 ( .A1(n9434), .A2(n5568), .ZN(n4431) );
  AND2_X1 U5955 ( .A1(n6076), .A2(n6075), .ZN(n4432) );
  NAND2_X1 U5956 ( .A1(n5652), .A2(n5651), .ZN(n6249) );
  INV_X1 U5957 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4936) );
  INV_X1 U5958 ( .A(n4628), .ZN(n4627) );
  NAND2_X1 U5959 ( .A1(n4629), .A2(n4630), .ZN(n4628) );
  AND2_X1 U5960 ( .A1(n4533), .A2(n4759), .ZN(n4433) );
  AND2_X1 U5961 ( .A1(n5813), .A2(n5814), .ZN(n4434) );
  INV_X1 U5962 ( .A(n4640), .ZN(n4639) );
  NAND2_X1 U5963 ( .A1(n9334), .A2(n8173), .ZN(n4640) );
  NAND2_X1 U5964 ( .A1(n9580), .A2(n5629), .ZN(n4435) );
  AND2_X1 U5965 ( .A1(n8433), .A2(n8435), .ZN(n8326) );
  AND2_X1 U5966 ( .A1(n4739), .A2(n4404), .ZN(n4436) );
  INV_X1 U5967 ( .A(n4474), .ZN(n4473) );
  NAND2_X1 U5968 ( .A1(n8246), .A2(n4475), .ZN(n4474) );
  AND2_X1 U5969 ( .A1(n5206), .A2(SI_11_), .ZN(n4437) );
  INV_X1 U5970 ( .A(n4806), .ZN(n4805) );
  AND2_X1 U5971 ( .A1(n5061), .A2(n4391), .ZN(n4438) );
  INV_X1 U5972 ( .A(n4488), .ZN(n4486) );
  AND2_X1 U5973 ( .A1(n4489), .A2(n5246), .ZN(n4488) );
  INV_X1 U5974 ( .A(n4493), .ZN(n4492) );
  NAND2_X1 U5975 ( .A1(n8024), .A2(n8112), .ZN(n4493) );
  AND2_X1 U5976 ( .A1(n4971), .A2(n4970), .ZN(n4439) );
  XNOR2_X1 U5977 ( .A(n4980), .B(P1_IR_REG_29__SCAN_IN), .ZN(n4981) );
  AND2_X1 U5978 ( .A1(n4483), .A2(n4480), .ZN(n4440) );
  NOR2_X1 U5979 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5795) );
  OAI22_X1 U5980 ( .A1(n4932), .A2(n4930), .B1(n5899), .B2(n5900), .ZN(n4929)
         );
  INV_X1 U5981 ( .A(n4929), .ZN(n4928) );
  AND2_X1 U5982 ( .A1(n5892), .A2(n5891), .ZN(n9917) );
  AND2_X1 U5983 ( .A1(n8475), .A2(n8474), .ZN(n4441) );
  INV_X1 U5984 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5547) );
  AND2_X1 U5985 ( .A1(n4401), .A2(n8903), .ZN(n4442) );
  NAND2_X1 U5986 ( .A1(n4922), .A2(n4924), .ZN(n5864) );
  NAND2_X1 U5987 ( .A1(n9344), .A2(n9321), .ZN(n4443) );
  NAND2_X1 U5988 ( .A1(n5102), .A2(n4564), .ZN(n4444) );
  AND2_X1 U5989 ( .A1(n7995), .A2(n7999), .ZN(n8154) );
  OR2_X1 U5990 ( .A1(n5426), .A2(n4615), .ZN(n4445) );
  AND2_X1 U5991 ( .A1(n5092), .A2(n5091), .ZN(n4446) );
  AND2_X1 U5992 ( .A1(n8980), .A2(n4627), .ZN(n4447) );
  NAND2_X1 U5993 ( .A1(n7772), .A2(n8106), .ZN(n7740) );
  INV_X1 U5994 ( .A(n8435), .ZN(n4846) );
  INV_X1 U5995 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5249) );
  XNOR2_X1 U5996 ( .A(n9079), .B(n8649), .ZN(n8436) );
  INV_X1 U5997 ( .A(n8436), .ZN(n4686) );
  OR2_X1 U5998 ( .A1(n7356), .A2(n8319), .ZN(n7283) );
  OR2_X1 U5999 ( .A1(n9139), .A2(n9577), .ZN(n4448) );
  NAND2_X1 U6000 ( .A1(n4917), .A2(n6063), .ZN(n8554) );
  OAI21_X1 U6001 ( .B1(n5916), .B2(n4935), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6020) );
  OR2_X1 U6002 ( .A1(n8462), .A2(n4382), .ZN(n4449) );
  NAND2_X1 U6003 ( .A1(n5508), .A2(n5507), .ZN(n9438) );
  OR2_X1 U6004 ( .A1(n9062), .A2(n8648), .ZN(n8453) );
  INV_X1 U6005 ( .A(n8453), .ZN(n4839) );
  NOR2_X1 U6006 ( .A1(n7821), .A2(n4687), .ZN(n4450) );
  NAND2_X1 U6007 ( .A1(n5336), .A2(n5335), .ZN(n9486) );
  NAND2_X1 U6008 ( .A1(n7781), .A2(n4669), .ZN(n4672) );
  AND2_X1 U6009 ( .A1(n9480), .A2(n9418), .ZN(n4451) );
  INV_X1 U6010 ( .A(n8804), .ZN(n9014) );
  NAND2_X1 U6011 ( .A1(n8291), .A2(n8290), .ZN(n8804) );
  INV_X1 U6012 ( .A(n4674), .ZN(n9345) );
  NOR2_X1 U6013 ( .A1(n9372), .A2(n4676), .ZN(n4674) );
  NOR3_X1 U6014 ( .A1(n9372), .A2(n9344), .A3(n4676), .ZN(n4673) );
  NAND2_X1 U6015 ( .A1(n6187), .A2(n6186), .ZN(n4452) );
  OR2_X1 U6016 ( .A1(n5916), .A2(n4938), .ZN(n4453) );
  INV_X1 U6017 ( .A(n6138), .ZN(n4914) );
  AND2_X1 U6018 ( .A1(n7810), .A2(n4845), .ZN(n4454) );
  AND2_X1 U6019 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(n4978), .ZN(n4455) );
  XNOR2_X1 U6020 ( .A(n4984), .B(n4983), .ZN(n5558) );
  INV_X1 U6021 ( .A(n8140), .ZN(n4660) );
  NAND2_X1 U6022 ( .A1(n7162), .A2(n7163), .ZN(n7159) );
  NAND2_X1 U6023 ( .A1(n5316), .A2(n5315), .ZN(n9490) );
  INV_X1 U6024 ( .A(n9490), .ZN(n4670) );
  AND2_X1 U6025 ( .A1(n4394), .A2(n6952), .ZN(n4456) );
  AND2_X1 U6026 ( .A1(n7433), .A2(n4392), .ZN(n4457) );
  AND2_X1 U6027 ( .A1(n7599), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4458) );
  NAND2_X1 U6028 ( .A1(n4689), .A2(n4688), .ZN(n7368) );
  AOI21_X1 U6029 ( .B1(n4446), .B2(n4390), .A(n4641), .ZN(n7506) );
  AND2_X1 U6030 ( .A1(n4867), .A2(n4866), .ZN(n7505) );
  NAND2_X1 U6031 ( .A1(n4681), .A2(n6842), .ZN(n6941) );
  AND2_X1 U6032 ( .A1(n4821), .A2(n4820), .ZN(n4459) );
  NAND2_X1 U6033 ( .A1(n6052), .A2(n6051), .ZN(n9062) );
  INV_X1 U6034 ( .A(n9062), .ZN(n4629) );
  NAND2_X1 U6035 ( .A1(n4551), .A2(n4549), .ZN(n5653) );
  AND2_X1 U6036 ( .A1(n8026), .A2(n8167), .ZN(n8114) );
  AND2_X1 U6037 ( .A1(n4820), .A2(n8379), .ZN(n4460) );
  AND2_X1 U6038 ( .A1(n5658), .A2(SI_29_), .ZN(n4461) );
  NAND2_X1 U6039 ( .A1(n5514), .A2(n5513), .ZN(n4462) );
  NAND2_X1 U6040 ( .A1(n8205), .A2(n9349), .ZN(n8079) );
  NAND2_X1 U6041 ( .A1(n5183), .A2(n5182), .ZN(n9830) );
  INV_X1 U6042 ( .A(n9830), .ZN(n4666) );
  NAND2_X1 U6043 ( .A1(n8310), .A2(n8360), .ZN(n7114) );
  INV_X1 U6044 ( .A(n9349), .ZN(n9778) );
  OR2_X1 U6045 ( .A1(n5691), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n4463) );
  NAND2_X1 U6046 ( .A1(n8308), .A2(n9873), .ZN(n4464) );
  INV_X1 U6047 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n4631) );
  NAND2_X1 U6048 ( .A1(n5031), .A2(n5030), .ZN(n4465) );
  OR2_X1 U6049 ( .A1(n8202), .A2(n4471), .ZN(n4470) );
  NAND2_X1 U6050 ( .A1(n4472), .A2(n4467), .ZN(P1_U3240) );
  OAI211_X1 U6051 ( .C1(n5228), .C2(n4481), .A(n4477), .B(n4476), .ZN(n6617)
         );
  NAND2_X1 U6052 ( .A1(n5228), .A2(n4440), .ZN(n4476) );
  OAI211_X1 U6053 ( .C1(n8022), .C2(n4493), .A(n8025), .B(n4490), .ZN(n8028)
         );
  NAND3_X1 U6054 ( .A1(n4501), .A2(n4500), .A3(n4499), .ZN(n4498) );
  NAND3_X1 U6055 ( .A1(n4586), .A2(n4987), .A3(n4988), .ZN(n5705) );
  NAND3_X1 U6056 ( .A1(n4509), .A2(n8051), .A3(n4505), .ZN(n8055) );
  OAI21_X1 U6057 ( .B1(n4508), .B2(n8035), .A(n4506), .ZN(n4505) );
  NOR2_X1 U6058 ( .A1(n8079), .A2(n4507), .ZN(n4506) );
  AOI21_X1 U6059 ( .B1(n8046), .B2(n8034), .A(n8033), .ZN(n4508) );
  NAND3_X1 U6060 ( .A1(n8170), .A2(n8079), .A3(n8047), .ZN(n4509) );
  AND2_X2 U6061 ( .A1(n5796), .A2(n5831), .ZN(n4924) );
  NAND2_X1 U6062 ( .A1(n8750), .A2(n4514), .ZN(n4513) );
  OAI211_X1 U6063 ( .C1(n8750), .C2(n4518), .A(n4517), .B(n4513), .ZN(n8761)
         );
  NAND2_X1 U6064 ( .A1(n4520), .A2(n4525), .ZN(n4524) );
  NAND2_X1 U6065 ( .A1(n8695), .A2(n8696), .ZN(n8699) );
  INV_X1 U6066 ( .A(n4520), .ZN(n8713) );
  NOR2_X1 U6067 ( .A1(n8698), .A2(n4522), .ZN(n4521) );
  INV_X1 U6068 ( .A(n8696), .ZN(n4522) );
  INV_X1 U6069 ( .A(n4524), .ZN(n8716) );
  INV_X1 U6070 ( .A(n8715), .ZN(n4523) );
  MUX2_X1 U6071 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n7118), .S(n6727), .Z(n9540)
         );
  NAND2_X1 U6072 ( .A1(n9178), .A2(n4537), .ZN(n4536) );
  INV_X1 U6073 ( .A(n4542), .ZN(n6431) );
  AND2_X1 U6074 ( .A1(n4542), .A2(n4541), .ZN(n9143) );
  INV_X1 U6075 ( .A(n6430), .ZN(n4541) );
  NAND3_X1 U6076 ( .A1(n6960), .A2(n7252), .A3(n4547), .ZN(n4546) );
  NAND2_X1 U6077 ( .A1(n6972), .A2(n6973), .ZN(n6960) );
  AOI21_X1 U6078 ( .B1(n5552), .B2(n4548), .A(n4455), .ZN(n4551) );
  NOR2_X1 U6079 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(n4978), .ZN(n4550) );
  INV_X1 U6080 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4552) );
  INV_X1 U6081 ( .A(n7756), .ZN(n4554) );
  OAI21_X1 U6082 ( .B1(n4554), .B2(n4557), .A(n4555), .ZN(n7904) );
  NAND2_X1 U6083 ( .A1(n8298), .A2(n8299), .ZN(n4600) );
  NAND2_X1 U6084 ( .A1(n4600), .A2(n8301), .ZN(n9005) );
  NAND2_X1 U6085 ( .A1(n5466), .A2(n4602), .ZN(n4601) );
  NAND2_X1 U6086 ( .A1(n5466), .A2(n5465), .ZN(n5485) );
  NAND2_X1 U6087 ( .A1(n4601), .A2(n4605), .ZN(n5517) );
  NAND2_X1 U6088 ( .A1(n5392), .A2(n4613), .ZN(n4610) );
  NAND2_X1 U6089 ( .A1(n4610), .A2(n4611), .ZN(n5449) );
  NAND2_X1 U6090 ( .A1(n5392), .A2(n4617), .ZN(n4616) );
  NAND2_X1 U6091 ( .A1(n5392), .A2(n5391), .ZN(n5411) );
  AND3_X2 U6092 ( .A1(n5746), .A2(n5745), .A3(n4950), .ZN(n6833) );
  INV_X1 U6093 ( .A(n4968), .ZN(n4632) );
  NAND2_X1 U6094 ( .A1(n5061), .A2(n4635), .ZN(n4634) );
  INV_X1 U6095 ( .A(n4903), .ZN(n4636) );
  AND2_X1 U6096 ( .A1(n5061), .A2(n5062), .ZN(n5102) );
  AOI21_X1 U6097 ( .B1(n8153), .B2(n8131), .A(n8154), .ZN(n4642) );
  OAI21_X1 U6098 ( .B1(n9395), .B2(n4646), .A(n4643), .ZN(n9364) );
  OAI21_X2 U6099 ( .B1(n8148), .B2(n4660), .A(n8138), .ZN(n7179) );
  NAND2_X1 U6100 ( .A1(n7200), .A2(n8214), .ZN(n8148) );
  NAND2_X2 U6101 ( .A1(n5558), .A2(n9619), .ZN(n5026) );
  XNOR2_X2 U6102 ( .A(n4661), .B(n4972), .ZN(n9619) );
  OAI21_X2 U6103 ( .B1(n5582), .B2(n4905), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4661) );
  NAND2_X1 U6104 ( .A1(n4406), .A2(n4662), .ZN(n9515) );
  AOI211_X1 U6105 ( .C1(n9293), .C2(n9431), .A(n9832), .B(n5663), .ZN(n9430)
         );
  INV_X1 U6106 ( .A(n4672), .ZN(n9405) );
  INV_X1 U6107 ( .A(n4673), .ZN(n9346) );
  NAND3_X1 U6108 ( .A1(n6947), .A2(n6946), .A3(n7086), .ZN(n4679) );
  NAND2_X1 U6109 ( .A1(n6947), .A2(n6946), .ZN(n7085) );
  NAND2_X1 U6110 ( .A1(n7356), .A2(n7282), .ZN(n4689) );
  NAND2_X1 U6111 ( .A1(n5706), .A2(n5711), .ZN(n5712) );
  NAND2_X1 U6112 ( .A1(n5709), .A2(n5706), .ZN(n6184) );
  NAND2_X1 U6113 ( .A1(n8904), .A2(n4442), .ZN(n4702) );
  NOR2_X1 U6114 ( .A1(n8898), .A2(n8920), .ZN(n4705) );
  NAND2_X1 U6115 ( .A1(n7371), .A2(n7370), .ZN(n7487) );
  OR2_X1 U6116 ( .A1(n9924), .A2(n8654), .ZN(n4712) );
  INV_X1 U6117 ( .A(n4716), .ZN(n4715) );
  NAND2_X2 U6118 ( .A1(n7929), .A2(n5698), .ZN(n5753) );
  NAND2_X2 U6119 ( .A1(n4715), .A2(n4713), .ZN(n5694) );
  NAND3_X1 U6120 ( .A1(n4732), .A2(n4730), .A3(n8493), .ZN(n4738) );
  NAND2_X1 U6121 ( .A1(n8476), .A2(n4731), .ZN(n4730) );
  OR2_X1 U6122 ( .A1(n5157), .A2(n4754), .ZN(n4750) );
  NAND2_X1 U6123 ( .A1(n5157), .A2(n4387), .ZN(n4748) );
  OAI21_X1 U6124 ( .B1(n9177), .B2(n4764), .A(n4757), .ZN(n9191) );
  NAND2_X1 U6125 ( .A1(n9162), .A2(n9163), .ZN(n4782) );
  NAND2_X1 U6126 ( .A1(n9162), .A2(n4776), .ZN(n4775) );
  NAND2_X1 U6127 ( .A1(n4782), .A2(n4780), .ZN(n9203) );
  AND2_X1 U6128 ( .A1(n4782), .A2(n4781), .ZN(n9206) );
  NAND2_X1 U6129 ( .A1(n6443), .A2(n6442), .ZN(n4781) );
  NAND2_X1 U6130 ( .A1(n6599), .A2(n4787), .ZN(n4783) );
  NAND2_X1 U6131 ( .A1(n4784), .A2(n4783), .ZN(n6327) );
  NAND2_X1 U6132 ( .A1(n6599), .A2(n7963), .ZN(n4786) );
  XNOR2_X1 U6133 ( .A(n9242), .B(n9257), .ZN(n9713) );
  OAI22_X1 U6134 ( .A1(n4801), .A2(n4800), .B1(n4802), .B2(n6519), .ZN(n6659)
         );
  INV_X1 U6135 ( .A(n4804), .ZN(n9644) );
  INV_X1 U6136 ( .A(n6519), .ZN(n4803) );
  NAND2_X1 U6137 ( .A1(n6704), .A2(n6517), .ZN(n4806) );
  MUX2_X1 U6138 ( .A(n6513), .B(P1_REG2_REG_1__SCAN_IN), .S(n6650), .Z(n6647)
         );
  NAND2_X1 U6139 ( .A1(n7264), .A2(n4814), .ZN(n4816) );
  NAND3_X1 U6140 ( .A1(n4816), .A2(n4817), .A3(n4815), .ZN(n7285) );
  NAND3_X1 U6141 ( .A1(n7265), .A2(n8374), .A3(n7089), .ZN(n4817) );
  NAND2_X1 U6142 ( .A1(n8379), .A2(n8380), .ZN(n4818) );
  AOI21_X1 U6143 ( .B1(n7372), .B2(n4828), .A(n4826), .ZN(n7536) );
  NAND2_X1 U6144 ( .A1(n4823), .A2(n4822), .ZN(n7537) );
  NAND2_X1 U6145 ( .A1(n7372), .A2(n4824), .ZN(n4823) );
  OAI21_X2 U6146 ( .B1(n8971), .B2(n4837), .A(n4834), .ZN(n8918) );
  NOR2_X1 U6147 ( .A1(n8918), .A2(n8919), .ZN(n8917) );
  NAND2_X1 U6148 ( .A1(n7792), .A2(n4843), .ZN(n4842) );
  NAND2_X1 U6149 ( .A1(n8819), .A2(n8287), .ZN(n8772) );
  NAND2_X1 U6150 ( .A1(n8819), .A2(n4847), .ZN(n8292) );
  NAND2_X1 U6151 ( .A1(n9891), .A2(n8663), .ZN(n8367) );
  NAND3_X1 U6152 ( .A1(n4851), .A2(n4955), .A3(n5011), .ZN(n5086) );
  OAI21_X1 U6153 ( .B1(n9403), .B2(n4855), .A(n4853), .ZN(n9371) );
  INV_X1 U6154 ( .A(n9403), .ZN(n4858) );
  NAND2_X1 U6155 ( .A1(n7403), .A2(n4862), .ZN(n4859) );
  NAND2_X1 U6156 ( .A1(n4860), .A2(n4859), .ZN(n7739) );
  NAND3_X1 U6157 ( .A1(n4982), .A2(n4981), .A3(P1_REG3_REG_1__SCAN_IN), .ZN(
        n4869) );
  NAND2_X1 U6158 ( .A1(n7919), .A2(n7853), .ZN(n4870) );
  NAND3_X1 U6159 ( .A1(n7919), .A2(n7853), .A3(P1_REG0_REG_1__SCAN_IN), .ZN(
        n4873) );
  NAND2_X1 U6160 ( .A1(n7853), .A2(n4982), .ZN(n5079) );
  NAND2_X1 U6161 ( .A1(n4871), .A2(n7853), .ZN(n4872) );
  NAND2_X1 U6162 ( .A1(n9301), .A2(n4886), .ZN(n4882) );
  AOI21_X1 U6163 ( .B1(n9301), .B2(n5649), .A(n4883), .ZN(n7947) );
  INV_X1 U6164 ( .A(n9438), .ZN(n4889) );
  NAND2_X1 U6165 ( .A1(n8266), .A2(n4892), .ZN(n4891) );
  OR2_X1 U6166 ( .A1(n5582), .A2(n4907), .ZN(n5573) );
  NAND2_X1 U6167 ( .A1(n5764), .A2(n5765), .ZN(n6918) );
  NAND2_X1 U6168 ( .A1(n8545), .A2(n5751), .ZN(n6919) );
  NAND3_X1 U6169 ( .A1(n8545), .A2(n5764), .A3(n4909), .ZN(n6920) );
  AND2_X1 U6170 ( .A1(n5765), .A2(n5751), .ZN(n4909) );
  NAND2_X1 U6171 ( .A1(n4910), .A2(n4912), .ZN(n6152) );
  NAND3_X1 U6172 ( .A1(n6123), .A2(n6122), .A3(n6138), .ZN(n4910) );
  NAND2_X1 U6173 ( .A1(n4915), .A2(n4916), .ZN(n6091) );
  NAND2_X1 U6174 ( .A1(n8603), .A2(n4918), .ZN(n4915) );
  OAI21_X1 U6175 ( .B1(n7475), .B2(n4929), .A(n4926), .ZN(n5915) );
  INV_X1 U6176 ( .A(n7475), .ZN(n4933) );
  NAND2_X1 U6177 ( .A1(n6003), .A2(n4934), .ZN(n6504) );
  NOR2_X1 U6178 ( .A1(n5916), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5932) );
  INV_X1 U6179 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4941) );
  NAND2_X1 U6180 ( .A1(n9406), .A2(n9393), .ZN(n9388) );
  AOI21_X1 U6181 ( .B1(n6447), .B2(n9235), .A(n6256), .ZN(n6688) );
  NAND2_X1 U6182 ( .A1(n6688), .A2(n6687), .ZN(n6690) );
  XNOR2_X1 U6183 ( .A(n5228), .B(n5227), .ZN(n6599) );
  NAND2_X1 U6184 ( .A1(n9292), .A2(n5572), .ZN(n9293) );
  INV_X1 U6185 ( .A(n6268), .ZN(n6974) );
  XNOR2_X1 U6186 ( .A(n6281), .B(n6452), .ZN(n7420) );
  NAND2_X1 U6187 ( .A1(n4979), .A2(n4973), .ZN(n9533) );
  NAND2_X1 U6188 ( .A1(n8345), .A2(n8367), .ZN(n8314) );
  XNOR2_X1 U6189 ( .A(n5546), .B(n8122), .ZN(n5557) );
  INV_X1 U6190 ( .A(n7198), .ZN(n5616) );
  OR2_X1 U6191 ( .A1(n5726), .A2(n5725), .ZN(n5728) );
  OAI222_X1 U6192 ( .A1(P2_U3152), .A2(n7929), .B1(n7928), .B2(n7927), .C1(
        n10118), .C2(n10258), .ZN(P2_U3328) );
  OR2_X1 U6193 ( .A1(n5079), .A2(n4995), .ZN(n4996) );
  XNOR2_X1 U6194 ( .A(n6091), .B(n6089), .ZN(n8611) );
  OR2_X1 U6195 ( .A1(n5763), .A2(n5762), .ZN(n5764) );
  OAI222_X1 U6196 ( .A1(n7924), .A2(n7854), .B1(P1_U3084), .B2(n7853), .C1(
        n7920), .C2(n7852), .ZN(P1_U3324) );
  INV_X1 U6197 ( .A(n4981), .ZN(n7853) );
  XNOR2_X1 U6198 ( .A(n5553), .B(P1_IR_REG_20__SCAN_IN), .ZN(n5611) );
  AND3_X1 U6199 ( .A1(n6471), .A2(n6472), .A3(n9204), .ZN(n4942) );
  INV_X1 U6200 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4972) );
  NOR2_X1 U6201 ( .A1(n5753), .A2(n5699), .ZN(n5700) );
  AND2_X1 U6202 ( .A1(n9554), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4943) );
  OR2_X1 U6203 ( .A1(n5587), .A2(n9776), .ZN(n4944) );
  NOR2_X1 U6204 ( .A1(n5644), .A2(n9362), .ZN(n4945) );
  NAND2_X1 U6205 ( .A1(n6492), .A2(n9204), .ZN(n4946) );
  INV_X1 U6206 ( .A(n8881), .ZN(n8284) );
  AND2_X1 U6207 ( .A1(n8848), .A2(n8846), .ZN(n4947) );
  OR2_X1 U6208 ( .A1(n6478), .A2(n10045), .ZN(n4948) );
  AND2_X1 U6209 ( .A1(n5588), .A2(n4944), .ZN(n4949) );
  AND2_X1 U6210 ( .A1(n5530), .A2(n5529), .ZN(n9139) );
  INV_X1 U6211 ( .A(n9139), .ZN(n5568) );
  OR2_X1 U6212 ( .A1(n5773), .A2(n6727), .ZN(n4950) );
  INV_X1 U6213 ( .A(n8379), .ZN(n7088) );
  OR2_X1 U6214 ( .A1(n8661), .A2(n8586), .ZN(n4951) );
  AND2_X1 U6215 ( .A1(n6251), .A2(n4948), .ZN(n4952) );
  OAI21_X1 U6216 ( .B1(n7635), .B2(n8327), .A(n7634), .ZN(n7636) );
  AND4_X2 U6217 ( .A1(n5758), .A2(n5757), .A3(n5756), .A4(n5755), .ZN(n4953)
         );
  NOR2_X1 U6218 ( .A1(n5069), .A2(n5068), .ZN(n4954) );
  NAND2_X1 U6219 ( .A1(n8053), .A2(n8079), .ZN(n8054) );
  AND2_X1 U6220 ( .A1(n5549), .A2(n5547), .ZN(n4965) );
  AND2_X1 U6221 ( .A1(n4966), .A2(n4965), .ZN(n4967) );
  NAND2_X1 U6222 ( .A1(n5356), .A2(n4967), .ZN(n4968) );
  NAND2_X1 U6223 ( .A1(n6259), .A2(n6456), .ZN(n6260) );
  OAI21_X1 U6224 ( .B1(n8591), .B2(n6110), .A(n6109), .ZN(n6111) );
  AND2_X1 U6225 ( .A1(n5688), .A2(n5729), .ZN(n5689) );
  INV_X1 U6226 ( .A(n7033), .ZN(n6301) );
  INV_X1 U6227 ( .A(n8260), .ZN(n5444) );
  OR2_X1 U6228 ( .A1(n6091), .A2(n6090), .ZN(n6092) );
  INV_X1 U6229 ( .A(n6082), .ZN(n6080) );
  INV_X1 U6230 ( .A(n6114), .ZN(n6099) );
  NOR2_X1 U6231 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5716) );
  NAND2_X1 U6232 ( .A1(n6255), .A2(n6254), .ZN(n6256) );
  AND2_X1 U6233 ( .A1(n9426), .A2(n8084), .ZN(n8241) );
  INV_X1 U6234 ( .A(n5397), .ZN(n5395) );
  INV_X1 U6235 ( .A(n7385), .ZN(n5115) );
  INV_X1 U6236 ( .A(n7020), .ZN(n5620) );
  AND2_X1 U6237 ( .A1(n5263), .A2(n5262), .ZN(n5264) );
  INV_X1 U6238 ( .A(n5178), .ZN(n5155) );
  OR2_X1 U6239 ( .A1(n5958), .A2(n5957), .ZN(n5984) );
  XNOR2_X1 U6240 ( .A(n5747), .B(n8550), .ZN(n5748) );
  AND2_X1 U6241 ( .A1(n5921), .A2(n5920), .ZN(n5936) );
  OR2_X1 U6242 ( .A1(n5875), .A2(n5874), .ZN(n5893) );
  NAND2_X1 U6243 ( .A1(n6080), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U6244 ( .A1(n6025), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6040) );
  OR2_X1 U6245 ( .A1(n5984), .A2(n5983), .ZN(n5986) );
  NAND2_X1 U6246 ( .A1(n6100), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6128) );
  NOR2_X1 U6247 ( .A1(n5849), .A2(n5848), .ZN(n5858) );
  AND2_X1 U6248 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5811) );
  NAND2_X1 U6249 ( .A1(n6099), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6116) );
  INV_X1 U6250 ( .A(n8317), .ZN(n7265) );
  INV_X1 U6251 ( .A(n5339), .ZN(n5337) );
  NAND2_X1 U6252 ( .A1(n5299), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5319) );
  XNOR2_X1 U6253 ( .A(n6279), .B(n6460), .ZN(n6289) );
  OR3_X1 U6254 ( .A1(n5436), .A2(n5435), .A3(n5434), .ZN(n5453) );
  OR2_X1 U6255 ( .A1(n5319), .A2(n5318), .ZN(n5339) );
  INV_X1 U6256 ( .A(n5039), .ZN(n5077) );
  OR2_X1 U6257 ( .A1(n5281), .A2(n5280), .ZN(n5300) );
  AOI21_X1 U6258 ( .B1(n5568), .B2(n9419), .A(n5567), .ZN(n5569) );
  INV_X1 U6259 ( .A(n7778), .ZN(n7846) );
  NAND2_X1 U6260 ( .A1(n5271), .A2(n5270), .ZN(n5286) );
  NAND2_X1 U6261 ( .A1(n5265), .A2(n5264), .ZN(n5269) );
  OR2_X1 U6262 ( .A1(n5130), .A2(n5129), .ZN(n5131) );
  OR2_X1 U6263 ( .A1(n6224), .A2(n6223), .ZN(n6225) );
  AOI21_X1 U6264 ( .B1(n8758), .B2(n9853), .A(n8757), .ZN(n8759) );
  INV_X1 U6265 ( .A(n9020), .ZN(n8812) );
  AND2_X1 U6266 ( .A1(n9072), .A2(n8779), .ZN(n8440) );
  INV_X1 U6267 ( .A(n8376), .ZN(n7086) );
  INV_X1 U6268 ( .A(n8342), .ZN(n8756) );
  NAND2_X1 U6269 ( .A1(n6218), .A2(n8497), .ZN(n8934) );
  AND2_X1 U6270 ( .A1(n8409), .A2(n8410), .ZN(n8324) );
  NAND2_X1 U6271 ( .A1(n6184), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5710) );
  INV_X1 U6272 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10257) );
  NAND2_X1 U6273 ( .A1(n7709), .A2(n7963), .ZN(n5508) );
  NAND2_X1 U6274 ( .A1(n5337), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5381) );
  INV_X1 U6275 ( .A(n9211), .ZN(n9186) );
  INV_X1 U6276 ( .A(n9225), .ZN(n9576) );
  OR2_X1 U6277 ( .A1(n6499), .A2(n6525), .ZN(n9577) );
  INV_X1 U6278 ( .A(n7038), .ZN(n9819) );
  INV_X1 U6279 ( .A(n7223), .ZN(n9801) );
  INV_X1 U6280 ( .A(n9500), .ZN(n9831) );
  NAND2_X1 U6281 ( .A1(n5449), .A2(n5448), .ZN(n5462) );
  NAND2_X1 U6282 ( .A1(n5372), .A2(n5371), .ZN(n5390) );
  AND2_X1 U6283 ( .A1(n5310), .A2(n5293), .ZN(n5308) );
  NAND2_X1 U6284 ( .A1(n5226), .A2(n5211), .ZN(n5227) );
  NAND2_X1 U6285 ( .A1(n5152), .A2(n10088), .ZN(n5156) );
  INV_X1 U6286 ( .A(n8627), .ZN(n8640) );
  AND4_X1 U6287 ( .A1(n6239), .A2(n6238), .A3(n6237), .A4(n6236), .ZN(n8816)
         );
  AND4_X1 U6288 ( .A1(n5910), .A2(n5909), .A3(n5908), .A4(n5907), .ZN(n7671)
         );
  NAND2_X1 U6289 ( .A1(n8448), .A2(n8450), .ZN(n8919) );
  INV_X1 U6290 ( .A(n8323), .ZN(n7367) );
  INV_X1 U6291 ( .A(n8801), .ZN(n9001) );
  INV_X1 U6292 ( .A(n9891), .ZN(n7071) );
  INV_X1 U6293 ( .A(n9931), .ZN(n9874) );
  AND2_X1 U6294 ( .A1(n6216), .A2(n6217), .ZN(n9922) );
  AND2_X1 U6295 ( .A1(n6197), .A2(n6196), .ZN(n9864) );
  INV_X1 U6296 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5833) );
  AND3_X1 U6297 ( .A1(n5404), .A2(n5403), .A3(n5402), .ZN(n9381) );
  AND2_X1 U6298 ( .A1(n8043), .A2(n8040), .ZN(n8271) );
  AND2_X1 U6299 ( .A1(n7973), .A2(n7972), .ZN(n8112) );
  AND2_X1 U6300 ( .A1(n8004), .A2(n8132), .ZN(n8106) );
  AND2_X1 U6301 ( .A1(n8127), .A2(n6525), .ZN(n9419) );
  AND2_X1 U6302 ( .A1(n9582), .A2(n7016), .ZN(n9505) );
  INV_X1 U6303 ( .A(n7016), .ZN(n9837) );
  XNOR2_X1 U6304 ( .A(n5048), .B(n5047), .ZN(n5775) );
  AND2_X1 U6305 ( .A1(n6245), .A2(n6244), .ZN(n6246) );
  INV_X1 U6306 ( .A(n8845), .ZN(n8989) );
  INV_X1 U6307 ( .A(n8905), .ZN(n9003) );
  INV_X1 U6308 ( .A(n9947), .ZN(n9945) );
  INV_X1 U6309 ( .A(n9935), .ZN(n9933) );
  INV_X1 U6310 ( .A(n9866), .ZN(n9868) );
  INV_X1 U6311 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6571) );
  INV_X1 U6312 ( .A(n9443), .ZN(n9307) );
  INV_X1 U6313 ( .A(n9341), .ZN(n9217) );
  OR2_X1 U6314 ( .A1(n5323), .A2(n5322), .ZN(n9420) );
  OR2_X1 U6315 ( .A1(n6883), .A2(n6882), .ZN(n9849) );
  NOR2_X1 U6316 ( .A1(n9840), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5677) );
  OR2_X1 U6317 ( .A1(n6883), .A2(n5676), .ZN(n9838) );
  INV_X1 U6318 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10132) );
  XNOR2_X1 U6319 ( .A(n5029), .B(n5028), .ZN(n6640) );
  AOI21_X1 U6320 ( .B1(n9603), .B2(n9840), .A(n5677), .ZN(P1_U3521) );
  NAND2_X1 U6321 ( .A1(n5249), .A2(n4956), .ZN(n5294) );
  INV_X1 U6322 ( .A(n5294), .ZN(n4959) );
  NOR2_X1 U6323 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4958) );
  NOR2_X1 U6324 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n4957) );
  NAND3_X1 U6325 ( .A1(n4959), .A2(n4958), .A3(n4957), .ZN(n4964) );
  NAND4_X1 U6326 ( .A1(n4962), .A2(n4961), .A3(n5312), .A4(n4960), .ZN(n4963)
         );
  NOR3_X1 U6327 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .A3(
        P1_IR_REG_22__SCAN_IN), .ZN(n4966) );
  INV_X1 U6328 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4971) );
  INV_X1 U6329 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4970) );
  INV_X1 U6330 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4983) );
  INV_X1 U6331 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4973) );
  NAND2_X1 U6332 ( .A1(n9533), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4974) );
  NAND2_X1 U6333 ( .A1(n4974), .A2(P1_IR_REG_30__SCAN_IN), .ZN(n4977) );
  INV_X1 U6334 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4975) );
  AND2_X1 U6335 ( .A1(n4975), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10247) );
  NAND2_X1 U6336 ( .A1(n9533), .A2(n10247), .ZN(n4976) );
  INV_X1 U6337 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4978) );
  INV_X1 U6338 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6513) );
  INV_X1 U6339 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7011) );
  INV_X1 U6340 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6552) );
  OR2_X1 U6341 ( .A1(n4380), .A2(n6552), .ZN(n4994) );
  AND2_X1 U6342 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4988) );
  NAND2_X1 U6343 ( .A1(n5134), .A2(n4989), .ZN(n5002) );
  INV_X1 U6344 ( .A(SI_1_), .ZN(n4990) );
  MUX2_X1 U6345 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5134), .Z(n5014) );
  XNOR2_X1 U6346 ( .A(n5015), .B(n5014), .ZN(n6555) );
  OR2_X1 U6347 ( .A1(n5180), .A2(n6555), .ZN(n4993) );
  INV_X1 U6348 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4991) );
  OR2_X1 U6349 ( .A1(n5026), .A2(n6650), .ZN(n4992) );
  NAND2_X1 U6350 ( .A1(n5039), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4999) );
  NAND2_X1 U6351 ( .A1(n5040), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n4998) );
  INV_X1 U6352 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7126) );
  INV_X1 U6353 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n4995) );
  NAND2_X1 U6354 ( .A1(n6553), .A2(SI_0_), .ZN(n5001) );
  INV_X1 U6355 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5000) );
  NAND2_X1 U6356 ( .A1(n5001), .A2(n5000), .ZN(n5003) );
  AND2_X1 U6357 ( .A1(n5003), .A2(n5002), .ZN(n9537) );
  MUX2_X1 U6358 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9537), .S(n5026), .Z(n7130) );
  INV_X1 U6359 ( .A(n7130), .ZN(n8210) );
  NOR2_X1 U6360 ( .A1(n9235), .A2(n8210), .ZN(n6889) );
  NAND2_X1 U6361 ( .A1(n8096), .A2(n6889), .ZN(n6888) );
  INV_X1 U6362 ( .A(n6258), .ZN(n8212) );
  NAND2_X1 U6363 ( .A1(n8212), .A2(n6259), .ZN(n5004) );
  NAND2_X1 U6364 ( .A1(n6888), .A2(n5004), .ZN(n7199) );
  INV_X1 U6365 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6530) );
  INV_X1 U6366 ( .A(n5005), .ZN(n5010) );
  INV_X1 U6367 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5007) );
  INV_X1 U6368 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6512) );
  OR2_X1 U6369 ( .A1(n5079), .A2(n6512), .ZN(n5006) );
  OAI21_X1 U6370 ( .B1(n4870), .B2(n5007), .A(n5006), .ZN(n5008) );
  INV_X1 U6371 ( .A(n5008), .ZN(n5009) );
  OR2_X1 U6372 ( .A1(n5011), .A2(n4978), .ZN(n5013) );
  INV_X1 U6373 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5012) );
  NAND2_X1 U6374 ( .A1(n5013), .A2(n5012), .ZN(n5027) );
  OAI21_X1 U6375 ( .B1(n5013), .B2(n5012), .A(n5027), .ZN(n9629) );
  INV_X1 U6376 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6565) );
  OR2_X1 U6377 ( .A1(n4380), .A2(n6565), .ZN(n5020) );
  NAND2_X1 U6378 ( .A1(n5015), .A2(n5014), .ZN(n5018) );
  NAND2_X1 U6379 ( .A1(n5016), .A2(SI_1_), .ZN(n5017) );
  INV_X1 U6380 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6570) );
  MUX2_X1 U6381 ( .A(n6570), .B(n6565), .S(n5134), .Z(n5032) );
  XNOR2_X1 U6382 ( .A(n5032), .B(SI_2_), .ZN(n5030) );
  XNOR2_X1 U6383 ( .A(n5031), .B(n5030), .ZN(n6569) );
  OR2_X1 U6384 ( .A1(n5180), .A2(n6569), .ZN(n5019) );
  OAI211_X1 U6385 ( .C1(n5026), .C2(n9629), .A(n5020), .B(n5019), .ZN(n7209)
         );
  NAND2_X1 U6386 ( .A1(n6974), .A2(n9796), .ZN(n8216) );
  NAND2_X1 U6387 ( .A1(n6268), .A2(n7209), .ZN(n8214) );
  NAND2_X1 U6388 ( .A1(n8216), .A2(n8214), .ZN(n5615) );
  NAND2_X1 U6389 ( .A1(n7199), .A2(n8092), .ZN(n7200) );
  OR2_X1 U6390 ( .A1(n5079), .A2(n7217), .ZN(n5022) );
  OR2_X1 U6391 ( .A1(n5539), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5021) );
  AND2_X1 U6392 ( .A1(n5022), .A2(n5021), .ZN(n5025) );
  NAND2_X1 U6393 ( .A1(n5666), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5024) );
  NAND2_X1 U6394 ( .A1(n5667), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5023) );
  NAND2_X1 U6395 ( .A1(n5027), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5029) );
  INV_X1 U6396 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5028) );
  INV_X1 U6397 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6559) );
  OR2_X1 U6398 ( .A1(n4381), .A2(n6559), .ZN(n5036) );
  INV_X1 U6399 ( .A(n5032), .ZN(n5033) );
  NAND2_X1 U6400 ( .A1(n5033), .A2(SI_2_), .ZN(n5034) );
  INV_X1 U6401 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6557) );
  MUX2_X1 U6402 ( .A(n6557), .B(n6559), .S(n5134), .Z(n5049) );
  XNOR2_X1 U6403 ( .A(n5049), .B(SI_3_), .ZN(n5047) );
  OR2_X1 U6404 ( .A1(n5180), .A2(n5775), .ZN(n5035) );
  OAI211_X1 U6405 ( .C1(n5026), .C2(n6640), .A(n5036), .B(n5035), .ZN(n7223)
         );
  NAND2_X1 U6406 ( .A1(n7201), .A2(n7223), .ZN(n8140) );
  INV_X1 U6407 ( .A(n7201), .ZN(n9233) );
  NAND2_X1 U6408 ( .A1(n9233), .A2(n9801), .ZN(n8138) );
  XNOR2_X1 U6409 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7185) );
  OR2_X1 U6410 ( .A1(n5539), .A2(n7185), .ZN(n5038) );
  INV_X1 U6411 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6517) );
  OR2_X1 U6412 ( .A1(n5079), .A2(n6517), .ZN(n5037) );
  AND2_X1 U6413 ( .A1(n5038), .A2(n5037), .ZN(n5043) );
  NAND2_X1 U6414 ( .A1(n5039), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5042) );
  NAND2_X1 U6415 ( .A1(n5040), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5041) );
  NAND2_X1 U6416 ( .A1(n5044), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5045) );
  MUX2_X1 U6417 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5045), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5046) );
  NAND2_X1 U6418 ( .A1(n5046), .A2(n5086), .ZN(n6704) );
  INV_X1 U6419 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6566) );
  OR2_X1 U6420 ( .A1(n4381), .A2(n6566), .ZN(n5053) );
  INV_X1 U6421 ( .A(n5049), .ZN(n5050) );
  NAND2_X1 U6422 ( .A1(n5050), .A2(SI_3_), .ZN(n5066) );
  NAND2_X1 U6423 ( .A1(n5071), .A2(n5066), .ZN(n5051) );
  MUX2_X1 U6424 ( .A(n10257), .B(n6566), .S(n5134), .Z(n5064) );
  XNOR2_X1 U6425 ( .A(n5064), .B(SI_4_), .ZN(n5068) );
  XNOR2_X1 U6426 ( .A(n5051), .B(n5068), .ZN(n10255) );
  OR2_X1 U6427 ( .A1(n5180), .A2(n10255), .ZN(n5052) );
  OAI211_X1 U6428 ( .C1(n5026), .C2(n6704), .A(n5053), .B(n5052), .ZN(n7192)
         );
  NAND2_X1 U6429 ( .A1(n7258), .A2(n7192), .ZN(n8218) );
  NAND2_X1 U6430 ( .A1(n7179), .A2(n8218), .ZN(n7441) );
  INV_X1 U6431 ( .A(n7258), .ZN(n9232) );
  INV_X1 U6432 ( .A(n7192), .ZN(n7187) );
  NAND2_X1 U6433 ( .A1(n9232), .A2(n7187), .ZN(n8139) );
  NAND2_X1 U6434 ( .A1(n7441), .A2(n8139), .ZN(n7021) );
  NAND3_X1 U6435 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5083) );
  INV_X1 U6436 ( .A(n5083), .ZN(n5054) );
  INV_X1 U6437 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6651) );
  NAND2_X1 U6438 ( .A1(n5083), .A2(n6651), .ZN(n5055) );
  NAND2_X1 U6439 ( .A1(n5095), .A2(n5055), .ZN(n7423) );
  OR2_X1 U6440 ( .A1(n5539), .A2(n7423), .ZN(n5057) );
  INV_X1 U6441 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6520) );
  OR2_X1 U6442 ( .A1(n5561), .A2(n6520), .ZN(n5056) );
  AND2_X1 U6443 ( .A1(n5057), .A2(n5056), .ZN(n5060) );
  NAND2_X1 U6444 ( .A1(n5666), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U6445 ( .A1(n5667), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5058) );
  OR2_X1 U6446 ( .A1(n5061), .A2(n4978), .ZN(n5063) );
  XNOR2_X1 U6447 ( .A(n5063), .B(n5062), .ZN(n6662) );
  OR2_X1 U6448 ( .A1(n4380), .A2(n6561), .ZN(n5076) );
  MUX2_X1 U6449 ( .A(n6571), .B(n6561), .S(n5134), .Z(n5104) );
  XNOR2_X1 U6450 ( .A(n5104), .B(SI_6_), .ZN(n5109) );
  INV_X1 U6451 ( .A(n5064), .ZN(n5065) );
  NAND2_X1 U6452 ( .A1(n5065), .A2(SI_4_), .ZN(n5067) );
  AND2_X1 U6453 ( .A1(n5066), .A2(n5067), .ZN(n5070) );
  INV_X1 U6454 ( .A(n5067), .ZN(n5069) );
  INV_X1 U6455 ( .A(n5741), .ZN(n5072) );
  MUX2_X1 U6456 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5072), .Z(n5073) );
  INV_X1 U6457 ( .A(SI_5_), .ZN(n10127) );
  NAND2_X1 U6458 ( .A1(n5128), .A2(n5126), .ZN(n5107) );
  NAND2_X1 U6459 ( .A1(n5073), .A2(SI_5_), .ZN(n5106) );
  NAND2_X1 U6460 ( .A1(n5107), .A2(n5106), .ZN(n5074) );
  XNOR2_X1 U6461 ( .A(n5109), .B(n5074), .ZN(n5835) );
  NAND2_X1 U6462 ( .A1(n7022), .A2(n7437), .ZN(n7978) );
  INV_X1 U6463 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6529) );
  INV_X1 U6464 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5078) );
  OAI22_X1 U6465 ( .A1(n5077), .A2(n6529), .B1(n4870), .B2(n5078), .ZN(n5085)
         );
  INV_X1 U6466 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6518) );
  INV_X1 U6467 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U6468 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5080) );
  NAND2_X1 U6469 ( .A1(n5081), .A2(n5080), .ZN(n5082) );
  NAND2_X1 U6470 ( .A1(n5083), .A2(n5082), .ZN(n9775) );
  OAI22_X1 U6471 ( .A1(n5561), .A2(n6518), .B1(n5539), .B2(n9775), .ZN(n5084)
         );
  INV_X1 U6472 ( .A(n9231), .ZN(n7181) );
  NAND2_X1 U6473 ( .A1(n5086), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5087) );
  XNOR2_X1 U6474 ( .A(n5087), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9643) );
  INV_X1 U6475 ( .A(n9643), .ZN(n6562) );
  XNOR2_X1 U6476 ( .A(n5128), .B(n5126), .ZN(n6567) );
  OR2_X1 U6477 ( .A1(n5180), .A2(n6567), .ZN(n5089) );
  INV_X1 U6478 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6563) );
  OR2_X1 U6479 ( .A1(n4381), .A2(n6563), .ZN(n5088) );
  OAI211_X2 U6480 ( .C1(n5026), .C2(n6562), .A(n5089), .B(n5088), .ZN(n9773)
         );
  NAND2_X1 U6481 ( .A1(n7181), .A2(n9773), .ZN(n7442) );
  AND2_X1 U6482 ( .A1(n7978), .A2(n7442), .ZN(n8219) );
  NAND2_X1 U6483 ( .A1(n7021), .A2(n8219), .ZN(n5092) );
  INV_X1 U6484 ( .A(n9773), .ZN(n5090) );
  AND2_X1 U6485 ( .A1(n9231), .A2(n5090), .ZN(n7439) );
  NAND2_X1 U6486 ( .A1(n7978), .A2(n7439), .ZN(n8137) );
  INV_X1 U6487 ( .A(n7022), .ZN(n9230) );
  NAND2_X1 U6488 ( .A1(n9230), .A2(n9812), .ZN(n7990) );
  AND2_X1 U6489 ( .A1(n8137), .A2(n7990), .ZN(n5091) );
  INV_X1 U6490 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U6491 ( .A1(n5095), .A2(n5094), .ZN(n5096) );
  NAND2_X1 U6492 ( .A1(n5117), .A2(n5096), .ZN(n7387) );
  OR2_X1 U6493 ( .A1(n5539), .A2(n7387), .ZN(n5098) );
  INV_X1 U6494 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7384) );
  OR2_X1 U6495 ( .A1(n5561), .A2(n7384), .ZN(n5097) );
  AND2_X1 U6496 ( .A1(n5098), .A2(n5097), .ZN(n5101) );
  NAND2_X1 U6497 ( .A1(n5667), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5100) );
  NAND2_X1 U6498 ( .A1(n5666), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5099) );
  OR2_X1 U6499 ( .A1(n5102), .A2(n4978), .ZN(n5103) );
  XNOR2_X1 U6500 ( .A(n5103), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6540) );
  INV_X1 U6501 ( .A(n6540), .ZN(n6681) );
  INV_X1 U6502 ( .A(n5104), .ZN(n5105) );
  NAND2_X1 U6503 ( .A1(n5105), .A2(SI_6_), .ZN(n5108) );
  NAND2_X1 U6504 ( .A1(n5107), .A2(n5129), .ZN(n5111) );
  INV_X1 U6505 ( .A(n5108), .ZN(n5110) );
  AND2_X1 U6506 ( .A1(n5111), .A2(n5125), .ZN(n5112) );
  INV_X1 U6507 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6573) );
  INV_X1 U6508 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6560) );
  MUX2_X1 U6509 ( .A(n6573), .B(n6560), .S(n5134), .Z(n5132) );
  XNOR2_X1 U6510 ( .A(n5112), .B(n5124), .ZN(n6572) );
  OR2_X1 U6511 ( .A1(n6572), .A2(n5180), .ZN(n5114) );
  OR2_X1 U6512 ( .A1(n4381), .A2(n6560), .ZN(n5113) );
  OAI211_X1 U6513 ( .C1(n5026), .C2(n6681), .A(n5114), .B(n5113), .ZN(n7038)
         );
  NAND2_X1 U6514 ( .A1(n7427), .A2(n7038), .ZN(n7977) );
  INV_X1 U6515 ( .A(n7427), .ZN(n9229) );
  NAND2_X1 U6516 ( .A1(n9229), .A2(n9819), .ZN(n7991) );
  NAND2_X1 U6517 ( .A1(n7977), .A2(n7991), .ZN(n7385) );
  INV_X1 U6518 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7169) );
  NAND2_X1 U6519 ( .A1(n5117), .A2(n7169), .ZN(n5118) );
  NAND2_X1 U6520 ( .A1(n5171), .A2(n5118), .ZN(n7408) );
  OR2_X1 U6521 ( .A1(n5539), .A2(n7408), .ZN(n5120) );
  INV_X1 U6522 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9659) );
  OR2_X1 U6523 ( .A1(n5561), .A2(n9659), .ZN(n5119) );
  AND2_X1 U6524 ( .A1(n5120), .A2(n5119), .ZN(n5123) );
  NAND2_X1 U6525 ( .A1(n5667), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U6526 ( .A1(n5666), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5121) );
  INV_X1 U6527 ( .A(n5130), .ZN(n5127) );
  INV_X1 U6528 ( .A(n5132), .ZN(n5133) );
  NAND2_X1 U6529 ( .A1(n5133), .A2(SI_7_), .ZN(n5148) );
  NAND2_X1 U6530 ( .A1(n5150), .A2(n5148), .ZN(n5139) );
  INV_X1 U6531 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6554) );
  MUX2_X1 U6532 ( .A(n6554), .B(n10115), .S(n5134), .Z(n5136) );
  INV_X1 U6533 ( .A(SI_8_), .ZN(n5135) );
  NAND2_X1 U6534 ( .A1(n5136), .A2(n5135), .ZN(n5151) );
  INV_X1 U6535 ( .A(n5136), .ZN(n5137) );
  NAND2_X1 U6536 ( .A1(n5137), .A2(SI_8_), .ZN(n5138) );
  XNOR2_X1 U6537 ( .A(n5139), .B(n5147), .ZN(n6564) );
  OR2_X1 U6538 ( .A1(n6564), .A2(n5180), .ZN(n5145) );
  INV_X1 U6539 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5140) );
  NAND2_X1 U6540 ( .A1(n5142), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5141) );
  MUX2_X1 U6541 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5141), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5143) );
  NAND2_X1 U6542 ( .A1(n5143), .A2(n4405), .ZN(n9658) );
  INV_X1 U6543 ( .A(n9658), .ZN(n9656) );
  AOI22_X1 U6544 ( .A1(n5359), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6501), .B2(
        n9656), .ZN(n5144) );
  NAND2_X1 U6545 ( .A1(n6309), .A2(n7410), .ZN(n7982) );
  NAND2_X1 U6546 ( .A1(n7982), .A2(n7977), .ZN(n8131) );
  INV_X1 U6547 ( .A(n8131), .ZN(n5146) );
  INV_X1 U6548 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6575) );
  MUX2_X1 U6549 ( .A(n6575), .B(n10132), .S(n5072), .Z(n5152) );
  INV_X1 U6550 ( .A(SI_9_), .ZN(n10088) );
  INV_X1 U6551 ( .A(n5152), .ZN(n5153) );
  NAND2_X1 U6552 ( .A1(n5153), .A2(SI_9_), .ZN(n5154) );
  INV_X1 U6553 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6581) );
  INV_X1 U6554 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6579) );
  INV_X1 U6555 ( .A(SI_10_), .ZN(n5158) );
  XNOR2_X1 U6556 ( .A(n5186), .B(n5185), .ZN(n6578) );
  NAND2_X1 U6557 ( .A1(n6578), .A2(n7963), .ZN(n5160) );
  NOR2_X1 U6558 ( .A1(n4405), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5213) );
  OR2_X1 U6559 ( .A1(n5213), .A2(n4978), .ZN(n5190) );
  XNOR2_X1 U6560 ( .A(n5190), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6871) );
  AOI22_X1 U6561 ( .A1(n5359), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6501), .B2(
        n6871), .ZN(n5159) );
  NAND2_X1 U6562 ( .A1(n5160), .A2(n5159), .ZN(n7574) );
  INV_X1 U6563 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5163) );
  INV_X1 U6564 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5170) );
  INV_X1 U6565 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6811) );
  NAND2_X1 U6566 ( .A1(n5173), .A2(n6811), .ZN(n5161) );
  NAND2_X1 U6567 ( .A1(n5197), .A2(n5161), .ZN(n7571) );
  OR2_X1 U6568 ( .A1(n5539), .A2(n7571), .ZN(n5162) );
  OAI21_X1 U6569 ( .B1(n5077), .B2(n5163), .A(n5162), .ZN(n5164) );
  INV_X1 U6570 ( .A(n5164), .ZN(n5169) );
  INV_X1 U6571 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5166) );
  INV_X1 U6572 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7572) );
  OR2_X1 U6573 ( .A1(n5561), .A2(n7572), .ZN(n5165) );
  OAI21_X1 U6574 ( .B1(n4870), .B2(n5166), .A(n5165), .ZN(n5167) );
  INV_X1 U6575 ( .A(n5167), .ZN(n5168) );
  NAND2_X1 U6576 ( .A1(n5666), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6577 ( .A1(n5667), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5176) );
  INV_X1 U6578 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7624) );
  OR2_X1 U6579 ( .A1(n5561), .A2(n7624), .ZN(n5175) );
  NAND2_X1 U6580 ( .A1(n5171), .A2(n5170), .ZN(n5172) );
  NAND2_X1 U6581 ( .A1(n5173), .A2(n5172), .ZN(n7939) );
  OR2_X1 U6582 ( .A1(n5539), .A2(n7939), .ZN(n5174) );
  NAND4_X1 U6583 ( .A1(n5177), .A2(n5176), .A3(n5175), .A4(n5174), .ZN(n9227)
         );
  INV_X1 U6584 ( .A(n9227), .ZN(n7401) );
  XNOR2_X1 U6585 ( .A(n5179), .B(n5178), .ZN(n6574) );
  OR2_X1 U6586 ( .A1(n6574), .A2(n5180), .ZN(n5183) );
  NAND2_X1 U6587 ( .A1(n4405), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5181) );
  XNOR2_X1 U6588 ( .A(n5181), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6815) );
  AOI22_X1 U6589 ( .A1(n5359), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6501), .B2(
        n6815), .ZN(n5182) );
  OR2_X1 U6590 ( .A1(n7401), .A2(n9830), .ZN(n7994) );
  NAND2_X1 U6591 ( .A1(n7999), .A2(n7994), .ZN(n7981) );
  INV_X1 U6592 ( .A(n7410), .ZN(n9823) );
  NAND2_X1 U6593 ( .A1(n9228), .A2(n9823), .ZN(n7993) );
  INV_X1 U6594 ( .A(n7993), .ZN(n5184) );
  NOR2_X1 U6595 ( .A1(n7981), .A2(n5184), .ZN(n8153) );
  NAND2_X1 U6596 ( .A1(n7574), .A2(n7935), .ZN(n7984) );
  NAND2_X1 U6597 ( .A1(n9830), .A2(n7401), .ZN(n7983) );
  NAND2_X1 U6598 ( .A1(n7984), .A2(n7983), .ZN(n7995) );
  INV_X1 U6599 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5188) );
  INV_X1 U6600 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10116) );
  MUX2_X1 U6601 ( .A(n5188), .B(n10116), .S(n6553), .Z(n5205) );
  XNOR2_X1 U6602 ( .A(n5207), .B(n5204), .ZN(n6576) );
  NAND2_X1 U6603 ( .A1(n6576), .A2(n7963), .ZN(n5194) );
  INV_X1 U6604 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5189) );
  NAND2_X1 U6605 ( .A1(n5190), .A2(n5189), .ZN(n5191) );
  NAND2_X1 U6606 ( .A1(n5191), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5192) );
  XNOR2_X1 U6607 ( .A(n5192), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9248) );
  AOI22_X1 U6608 ( .A1(n5359), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6501), .B2(
        n9248), .ZN(n5193) );
  NAND2_X1 U6609 ( .A1(n5666), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5202) );
  NAND2_X1 U6610 ( .A1(n5667), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5201) );
  INV_X1 U6611 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7514) );
  OR2_X1 U6612 ( .A1(n5561), .A2(n7514), .ZN(n5200) );
  INV_X1 U6613 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U6614 ( .A1(n5197), .A2(n5196), .ZN(n5198) );
  NAND2_X1 U6615 ( .A1(n5217), .A2(n5198), .ZN(n7513) );
  OR2_X1 U6616 ( .A1(n5539), .A2(n7513), .ZN(n5199) );
  NAND4_X1 U6617 ( .A1(n5202), .A2(n5201), .A3(n5200), .A4(n5199), .ZN(n9225)
         );
  NAND2_X1 U6618 ( .A1(n7516), .A2(n9576), .ZN(n8003) );
  NAND2_X1 U6619 ( .A1(n7506), .A2(n8003), .ZN(n5203) );
  OR2_X1 U6620 ( .A1(n7516), .A2(n9576), .ZN(n8005) );
  INV_X1 U6621 ( .A(n5205), .ZN(n5206) );
  INV_X1 U6622 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6602) );
  INV_X1 U6623 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5208) );
  MUX2_X1 U6624 ( .A(n6602), .B(n5208), .S(n6553), .Z(n5209) );
  INV_X1 U6625 ( .A(SI_12_), .ZN(n10018) );
  INV_X1 U6626 ( .A(n5209), .ZN(n5210) );
  NAND2_X1 U6627 ( .A1(n5210), .A2(SI_12_), .ZN(n5211) );
  NOR2_X1 U6628 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5212) );
  NAND2_X1 U6629 ( .A1(n5213), .A2(n5212), .ZN(n5234) );
  NAND2_X1 U6630 ( .A1(n5234), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5214) );
  XNOR2_X1 U6631 ( .A(n5214), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9675) );
  AOI22_X1 U6632 ( .A1(n5359), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6501), .B2(
        n9675), .ZN(n5215) );
  INV_X1 U6633 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7528) );
  NAND2_X1 U6634 ( .A1(n5217), .A2(n7528), .ZN(n5218) );
  NAND2_X1 U6635 ( .A1(n5240), .A2(n5218), .ZN(n9587) );
  OR2_X1 U6636 ( .A1(n5539), .A2(n9587), .ZN(n5221) );
  INV_X1 U6637 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n5219) );
  OR2_X1 U6638 ( .A1(n5561), .A2(n5219), .ZN(n5220) );
  AND2_X1 U6639 ( .A1(n5221), .A2(n5220), .ZN(n5224) );
  NAND2_X1 U6640 ( .A1(n5666), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5223) );
  NAND2_X1 U6641 ( .A1(n5667), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5222) );
  OR2_X1 U6642 ( .A1(n9593), .A2(n7551), .ZN(n8006) );
  INV_X1 U6643 ( .A(n8006), .ZN(n5225) );
  NAND2_X1 U6644 ( .A1(n9593), .A2(n7551), .ZN(n8007) );
  INV_X1 U6645 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9993) );
  INV_X1 U6646 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5229) );
  MUX2_X1 U6647 ( .A(n9993), .B(n5229), .S(n6553), .Z(n5231) );
  INV_X1 U6648 ( .A(SI_13_), .ZN(n5230) );
  INV_X1 U6649 ( .A(n5231), .ZN(n5232) );
  NAND2_X1 U6650 ( .A1(n5232), .A2(SI_13_), .ZN(n5233) );
  XNOR2_X1 U6651 ( .A(n5247), .B(n5246), .ZN(n6614) );
  NAND2_X1 U6652 ( .A1(n6614), .A2(n7963), .ZN(n5237) );
  NAND2_X1 U6653 ( .A1(n5248), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5235) );
  XNOR2_X1 U6654 ( .A(n5235), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9684) );
  AOI22_X1 U6655 ( .A1(n5359), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6501), .B2(
        n9684), .ZN(n5236) );
  NAND2_X1 U6656 ( .A1(n5666), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5245) );
  NAND2_X1 U6657 ( .A1(n5667), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5244) );
  INV_X1 U6658 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n5238) );
  OR2_X1 U6659 ( .A1(n5561), .A2(n5238), .ZN(n5243) );
  INV_X1 U6660 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6661 ( .A1(n5240), .A2(n5239), .ZN(n5241) );
  NAND2_X1 U6662 ( .A1(n5255), .A2(n5241), .ZN(n7768) );
  OR2_X1 U6663 ( .A1(n5539), .A2(n7768), .ZN(n5242) );
  NAND4_X1 U6664 ( .A1(n5245), .A2(n5244), .A3(n5243), .A4(n5242), .ZN(n9223)
         );
  INV_X1 U6665 ( .A(n9223), .ZN(n9578) );
  OR2_X1 U6666 ( .A1(n9501), .A2(n9578), .ZN(n8004) );
  NAND2_X1 U6667 ( .A1(n9501), .A2(n9578), .ZN(n8132) );
  INV_X1 U6668 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6618) );
  INV_X1 U6669 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6620) );
  MUX2_X1 U6670 ( .A(n6618), .B(n6620), .S(n6553), .Z(n5266) );
  XNOR2_X1 U6671 ( .A(n5266), .B(SI_14_), .ZN(n5262) );
  NAND2_X1 U6672 ( .A1(n6617), .A2(n7963), .ZN(n5252) );
  NAND2_X1 U6673 ( .A1(n5295), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5250) );
  NAND2_X1 U6674 ( .A1(n5250), .A2(n5249), .ZN(n5274) );
  OAI21_X1 U6675 ( .B1(n5250), .B2(n5249), .A(n5274), .ZN(n9255) );
  INV_X1 U6676 ( .A(n9255), .ZN(n9699) );
  AOI22_X1 U6677 ( .A1(n5359), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6501), .B2(
        n9699), .ZN(n5251) );
  INV_X1 U6678 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9254) );
  INV_X1 U6679 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5253) );
  OAI22_X1 U6680 ( .A1(n5077), .A2(n9254), .B1(n4870), .B2(n5253), .ZN(n5258)
         );
  INV_X1 U6681 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7749) );
  INV_X1 U6682 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7582) );
  NAND2_X1 U6683 ( .A1(n5255), .A2(n7582), .ZN(n5256) );
  NAND2_X1 U6684 ( .A1(n5281), .A2(n5256), .ZN(n7748) );
  OAI22_X1 U6685 ( .A1(n5561), .A2(n7749), .B1(n5539), .B2(n7748), .ZN(n5257)
         );
  INV_X1 U6686 ( .A(n9222), .ZN(n5259) );
  NAND2_X1 U6687 ( .A1(n7751), .A2(n5259), .ZN(n8134) );
  NAND2_X1 U6688 ( .A1(n8015), .A2(n8134), .ZN(n8108) );
  INV_X1 U6689 ( .A(n8132), .ZN(n8014) );
  NOR2_X1 U6690 ( .A1(n8108), .A2(n8014), .ZN(n5260) );
  NAND2_X1 U6691 ( .A1(n7740), .A2(n5260), .ZN(n5261) );
  NAND2_X1 U6692 ( .A1(n5261), .A2(n8015), .ZN(n7779) );
  INV_X1 U6693 ( .A(n5266), .ZN(n5267) );
  NAND2_X1 U6694 ( .A1(n5267), .A2(SI_14_), .ZN(n5268) );
  INV_X1 U6695 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10094) );
  INV_X1 U6696 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6623) );
  MUX2_X1 U6697 ( .A(n10094), .B(n6623), .S(n6553), .Z(n5271) );
  INV_X1 U6698 ( .A(SI_15_), .ZN(n5270) );
  INV_X1 U6699 ( .A(n5271), .ZN(n5272) );
  NAND2_X1 U6700 ( .A1(n5272), .A2(SI_15_), .ZN(n5273) );
  XNOR2_X1 U6701 ( .A(n5288), .B(n5287), .ZN(n6621) );
  NAND2_X1 U6702 ( .A1(n6621), .A2(n7963), .ZN(n5277) );
  NAND2_X1 U6703 ( .A1(n5274), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5275) );
  XNOR2_X1 U6704 ( .A(n5275), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9716) );
  AOI22_X1 U6705 ( .A1(n5359), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9716), .B2(
        n6501), .ZN(n5276) );
  INV_X1 U6706 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5279) );
  INV_X1 U6707 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5278) );
  OAI22_X1 U6708 ( .A1(n5077), .A2(n5279), .B1(n4870), .B2(n5278), .ZN(n5285)
         );
  INV_X1 U6709 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n5283) );
  INV_X1 U6710 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U6711 ( .A1(n5281), .A2(n5280), .ZN(n5282) );
  NAND2_X1 U6712 ( .A1(n5300), .A2(n5282), .ZN(n7782) );
  OAI22_X1 U6713 ( .A1(n5561), .A2(n5283), .B1(n5539), .B2(n7782), .ZN(n5284)
         );
  INV_X1 U6714 ( .A(n9221), .ZN(n7858) );
  NAND2_X1 U6715 ( .A1(n7778), .A2(n7858), .ZN(n8156) );
  INV_X1 U6716 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5290) );
  INV_X1 U6717 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5289) );
  MUX2_X1 U6718 ( .A(n5290), .B(n5289), .S(n6553), .Z(n5291) );
  INV_X1 U6719 ( .A(SI_16_), .ZN(n10191) );
  NAND2_X1 U6720 ( .A1(n5291), .A2(n10191), .ZN(n5310) );
  INV_X1 U6721 ( .A(n5291), .ZN(n5292) );
  NAND2_X1 U6722 ( .A1(n5292), .A2(SI_16_), .ZN(n5293) );
  XNOR2_X1 U6723 ( .A(n5309), .B(n5308), .ZN(n6624) );
  NAND2_X1 U6724 ( .A1(n6624), .A2(n7963), .ZN(n5298) );
  NOR2_X1 U6725 ( .A1(n5295), .A2(n5294), .ZN(n5313) );
  OR2_X1 U6726 ( .A1(n5313), .A2(n4978), .ZN(n5296) );
  XNOR2_X1 U6727 ( .A(n5296), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9728) );
  AOI22_X1 U6728 ( .A1(n5359), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9728), .B2(
        n6501), .ZN(n5297) );
  INV_X1 U6729 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n10048) );
  NAND2_X1 U6730 ( .A1(n5300), .A2(n10048), .ZN(n5301) );
  NAND2_X1 U6731 ( .A1(n5319), .A2(n5301), .ZN(n7760) );
  OR2_X1 U6732 ( .A1(n5539), .A2(n7760), .ZN(n5304) );
  INV_X1 U6733 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5302) );
  OR2_X1 U6734 ( .A1(n5561), .A2(n5302), .ZN(n5303) );
  AND2_X1 U6735 ( .A1(n5304), .A2(n5303), .ZN(n5307) );
  NAND2_X1 U6736 ( .A1(n5667), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6737 ( .A1(n5666), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5305) );
  OR2_X1 U6738 ( .A1(n9497), .A2(n7876), .ZN(n8149) );
  NAND2_X1 U6739 ( .A1(n9497), .A2(n7876), .ZN(n8023) );
  NAND2_X1 U6740 ( .A1(n8149), .A2(n8023), .ZN(n8021) );
  INV_X1 U6741 ( .A(n8021), .ZN(n8110) );
  INV_X1 U6742 ( .A(n8023), .ZN(n8161) );
  AOI21_X2 U6743 ( .B1(n7856), .B2(n8110), .A(n8161), .ZN(n7872) );
  INV_X1 U6744 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6667) );
  INV_X1 U6745 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5311) );
  MUX2_X1 U6746 ( .A(n6667), .B(n5311), .S(n6553), .Z(n5325) );
  XNOR2_X1 U6747 ( .A(n5325), .B(SI_17_), .ZN(n5324) );
  XNOR2_X1 U6748 ( .A(n5329), .B(n5324), .ZN(n6663) );
  NAND2_X1 U6749 ( .A1(n6663), .A2(n7963), .ZN(n5316) );
  NAND2_X1 U6750 ( .A1(n5313), .A2(n5312), .ZN(n5314) );
  NAND2_X1 U6751 ( .A1(n5314), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5331) );
  XNOR2_X1 U6752 ( .A(n5331), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9739) );
  AOI22_X1 U6753 ( .A1(n9739), .A2(n6501), .B1(n5359), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n5315) );
  INV_X1 U6754 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9261) );
  INV_X1 U6755 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n5317) );
  OAI22_X1 U6756 ( .A1(n5077), .A2(n9261), .B1(n4870), .B2(n5317), .ZN(n5323)
         );
  INV_X1 U6757 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n5321) );
  INV_X1 U6758 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5318) );
  NAND2_X1 U6759 ( .A1(n5319), .A2(n5318), .ZN(n5320) );
  NAND2_X1 U6760 ( .A1(n5339), .A2(n5320), .ZN(n7869) );
  OAI22_X1 U6761 ( .A1(n5561), .A2(n5321), .B1(n5539), .B2(n7869), .ZN(n5322)
         );
  INV_X1 U6762 ( .A(n9420), .ZN(n7888) );
  OR2_X1 U6763 ( .A1(n9490), .A2(n7888), .ZN(n7973) );
  NAND2_X1 U6764 ( .A1(n9490), .A2(n7888), .ZN(n7972) );
  NAND2_X1 U6765 ( .A1(n7872), .A2(n8112), .ZN(n7873) );
  INV_X1 U6766 ( .A(n5324), .ZN(n5328) );
  INV_X1 U6767 ( .A(n5325), .ZN(n5326) );
  NAND2_X1 U6768 ( .A1(n5326), .A2(SI_17_), .ZN(n5327) );
  MUX2_X1 U6769 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6553), .Z(n5350) );
  XNOR2_X1 U6770 ( .A(n5350), .B(SI_18_), .ZN(n5347) );
  XNOR2_X1 U6771 ( .A(n5349), .B(n5347), .ZN(n6823) );
  NAND2_X1 U6772 ( .A1(n6823), .A2(n7963), .ZN(n5336) );
  INV_X1 U6773 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5330) );
  NAND2_X1 U6774 ( .A1(n5331), .A2(n5330), .ZN(n5332) );
  NAND2_X1 U6775 ( .A1(n5332), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5333) );
  XNOR2_X1 U6776 ( .A(n5333), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9752) );
  INV_X1 U6777 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10004) );
  NOR2_X1 U6778 ( .A1(n4380), .A2(n10004), .ZN(n5334) );
  AOI21_X1 U6779 ( .B1(n9752), .B2(n6501), .A(n5334), .ZN(n5335) );
  INV_X1 U6780 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U6781 ( .A1(n5339), .A2(n5338), .ZN(n5340) );
  NAND2_X1 U6782 ( .A1(n5381), .A2(n5340), .ZN(n9407) );
  OR2_X1 U6783 ( .A1(n5539), .A2(n9407), .ZN(n5342) );
  INV_X1 U6784 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9247) );
  OR2_X1 U6785 ( .A1(n5561), .A2(n9247), .ZN(n5341) );
  AND2_X1 U6786 ( .A1(n5342), .A2(n5341), .ZN(n5345) );
  NAND2_X1 U6787 ( .A1(n5667), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5344) );
  NAND2_X1 U6788 ( .A1(n5666), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5343) );
  OR2_X1 U6789 ( .A1(n9486), .A2(n7909), .ZN(n8026) );
  NAND2_X1 U6790 ( .A1(n9486), .A2(n7909), .ZN(n8167) );
  INV_X1 U6791 ( .A(n8114), .ZN(n9412) );
  INV_X1 U6792 ( .A(n7973), .ZN(n9413) );
  NOR2_X1 U6793 ( .A1(n9412), .A2(n9413), .ZN(n5346) );
  NAND2_X1 U6794 ( .A1(n7873), .A2(n5346), .ZN(n9415) );
  NAND2_X1 U6795 ( .A1(n9415), .A2(n8167), .ZN(n9395) );
  INV_X1 U6796 ( .A(n5347), .ZN(n5348) );
  NAND2_X1 U6797 ( .A1(n5350), .A2(SI_18_), .ZN(n5351) );
  INV_X1 U6798 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7926) );
  INV_X1 U6799 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10050) );
  MUX2_X1 U6800 ( .A(n7926), .B(n10050), .S(n6553), .Z(n5353) );
  INV_X1 U6801 ( .A(SI_19_), .ZN(n10092) );
  NAND2_X1 U6802 ( .A1(n5353), .A2(n10092), .ZN(n5371) );
  INV_X1 U6803 ( .A(n5353), .ZN(n5354) );
  NAND2_X1 U6804 ( .A1(n5354), .A2(SI_19_), .ZN(n5355) );
  NAND2_X1 U6805 ( .A1(n5371), .A2(n5355), .ZN(n5368) );
  XNOR2_X1 U6806 ( .A(n5367), .B(n5368), .ZN(n6917) );
  NAND2_X1 U6807 ( .A1(n6917), .A2(n7963), .ZN(n5361) );
  INV_X1 U6808 ( .A(n5356), .ZN(n5357) );
  NAND2_X1 U6809 ( .A1(n4444), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5358) );
  AOI22_X1 U6810 ( .A1(n5359), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9349), .B2(
        n6501), .ZN(n5360) );
  NAND2_X1 U6811 ( .A1(n5667), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U6812 ( .A1(n5666), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5365) );
  XNOR2_X1 U6813 ( .A(n5381), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n9391) );
  INV_X1 U6814 ( .A(n5539), .ZN(n5512) );
  NAND2_X1 U6815 ( .A1(n9391), .A2(n5512), .ZN(n5364) );
  INV_X1 U6816 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n5362) );
  OR2_X1 U6817 ( .A1(n5561), .A2(n5362), .ZN(n5363) );
  NAND4_X1 U6818 ( .A1(n5366), .A2(n5365), .A3(n5364), .A4(n5363), .ZN(n9418)
         );
  INV_X1 U6819 ( .A(n9418), .ZN(n9380) );
  OR2_X1 U6820 ( .A1(n9480), .A2(n9380), .ZN(n8029) );
  NAND2_X1 U6821 ( .A1(n9480), .A2(n9380), .ZN(n8165) );
  INV_X1 U6822 ( .A(n5367), .ZN(n5370) );
  INV_X1 U6823 ( .A(n5368), .ZN(n5369) );
  NAND2_X1 U6824 ( .A1(n5370), .A2(n5369), .ZN(n5372) );
  INV_X1 U6825 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8278) );
  INV_X1 U6826 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6971) );
  MUX2_X1 U6827 ( .A(n8278), .B(n6971), .S(n6553), .Z(n5373) );
  INV_X1 U6828 ( .A(SI_20_), .ZN(n10101) );
  NAND2_X1 U6829 ( .A1(n5373), .A2(n10101), .ZN(n5391) );
  INV_X1 U6830 ( .A(n5373), .ZN(n5374) );
  NAND2_X1 U6831 ( .A1(n5374), .A2(SI_20_), .ZN(n5375) );
  XNOR2_X1 U6832 ( .A(n5390), .B(n5389), .ZN(n6970) );
  NAND2_X1 U6833 ( .A1(n6970), .A2(n7963), .ZN(n5377) );
  OR2_X1 U6834 ( .A1(n4381), .A2(n6971), .ZN(n5376) );
  INV_X1 U6835 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5379) );
  INV_X1 U6836 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5378) );
  OAI21_X1 U6837 ( .B1(n5381), .B2(n5379), .A(n5378), .ZN(n5382) );
  NAND2_X1 U6838 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5380) );
  NAND2_X1 U6839 ( .A1(n5382), .A2(n5397), .ZN(n9374) );
  INV_X1 U6840 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n5383) );
  OAI22_X1 U6841 ( .A1(n9374), .A2(n5539), .B1(n5561), .B2(n5383), .ZN(n5387)
         );
  INV_X1 U6842 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5385) );
  INV_X1 U6843 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n5384) );
  OAI22_X1 U6844 ( .A1(n5077), .A2(n5385), .B1(n4870), .B2(n5384), .ZN(n5386)
         );
  INV_X1 U6845 ( .A(n9396), .ZN(n5388) );
  NAND2_X1 U6846 ( .A1(n9476), .A2(n5388), .ZN(n8036) );
  NAND2_X1 U6847 ( .A1(n8034), .A2(n8036), .ZN(n9379) );
  NAND2_X1 U6848 ( .A1(n5390), .A2(n5389), .ZN(n5392) );
  INV_X1 U6849 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6982) );
  INV_X1 U6850 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7000) );
  MUX2_X1 U6851 ( .A(n6982), .B(n7000), .S(n6553), .Z(n5407) );
  XNOR2_X1 U6852 ( .A(n5407), .B(SI_21_), .ZN(n5406) );
  XNOR2_X1 U6853 ( .A(n5411), .B(n5406), .ZN(n6981) );
  NAND2_X1 U6854 ( .A1(n6981), .A2(n7963), .ZN(n5394) );
  OR2_X1 U6855 ( .A1(n4380), .A2(n7000), .ZN(n5393) );
  NAND2_X2 U6856 ( .A1(n5394), .A2(n5393), .ZN(n9471) );
  INV_X1 U6857 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U6858 ( .A1(n5397), .A2(n5396), .ZN(n5398) );
  NAND2_X1 U6859 ( .A1(n5436), .A2(n5398), .ZN(n9358) );
  OR2_X1 U6860 ( .A1(n9358), .A2(n5539), .ZN(n5404) );
  INV_X1 U6861 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5399) );
  INV_X1 U6862 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10142) );
  OAI22_X1 U6863 ( .A1(n5077), .A2(n5399), .B1(n4870), .B2(n10142), .ZN(n5400)
         );
  INV_X1 U6864 ( .A(n5400), .ZN(n5403) );
  INV_X1 U6865 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n5401) );
  OR2_X1 U6866 ( .A1(n5561), .A2(n5401), .ZN(n5402) );
  OR2_X1 U6867 ( .A1(n9471), .A2(n9381), .ZN(n8042) );
  NAND2_X1 U6868 ( .A1(n9471), .A2(n9381), .ZN(n8038) );
  NAND2_X1 U6869 ( .A1(n8042), .A2(n8038), .ZN(n9362) );
  INV_X1 U6870 ( .A(n8034), .ZN(n9363) );
  NOR2_X1 U6871 ( .A1(n9362), .A2(n9363), .ZN(n5405) );
  NAND2_X1 U6872 ( .A1(n9364), .A2(n8038), .ZN(n8272) );
  INV_X1 U6873 ( .A(n5406), .ZN(n5410) );
  INV_X1 U6874 ( .A(n5407), .ZN(n5408) );
  NAND2_X1 U6875 ( .A1(n5408), .A2(SI_21_), .ZN(n5409) );
  INV_X1 U6876 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7246) );
  INV_X1 U6877 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7923) );
  MUX2_X1 U6878 ( .A(n7246), .B(n7923), .S(n6553), .Z(n5413) );
  INV_X1 U6879 ( .A(SI_22_), .ZN(n5412) );
  NAND2_X1 U6880 ( .A1(n5413), .A2(n5412), .ZN(n5425) );
  INV_X1 U6881 ( .A(n5413), .ZN(n5414) );
  NAND2_X1 U6882 ( .A1(n5414), .A2(SI_22_), .ZN(n5415) );
  NAND2_X1 U6883 ( .A1(n5425), .A2(n5415), .ZN(n5426) );
  XNOR2_X1 U6884 ( .A(n5427), .B(n5426), .ZN(n7245) );
  NAND2_X1 U6885 ( .A1(n7245), .A2(n7963), .ZN(n5417) );
  OR2_X1 U6886 ( .A1(n4381), .A2(n7923), .ZN(n5416) );
  XNOR2_X1 U6887 ( .A(n5436), .B(P1_REG3_REG_22__SCAN_IN), .ZN(n9195) );
  NAND2_X1 U6888 ( .A1(n9195), .A2(n5512), .ZN(n5423) );
  INV_X1 U6889 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6890 ( .A1(n5667), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U6891 ( .A1(n5666), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5418) );
  OAI211_X1 U6892 ( .C1(n5420), .C2(n5561), .A(n5419), .B(n5418), .ZN(n5421)
         );
  INV_X1 U6893 ( .A(n5421), .ZN(n5422) );
  NAND2_X1 U6894 ( .A1(n5423), .A2(n5422), .ZN(n9366) );
  INV_X1 U6895 ( .A(n9366), .ZN(n9151) );
  OR2_X1 U6896 ( .A1(n9465), .A2(n9151), .ZN(n8043) );
  NAND2_X1 U6897 ( .A1(n9465), .A2(n9151), .ZN(n8040) );
  NAND2_X1 U6898 ( .A1(n8272), .A2(n8271), .ZN(n5424) );
  NAND2_X1 U6899 ( .A1(n5424), .A2(n8040), .ZN(n8257) );
  INV_X1 U6900 ( .A(n8257), .ZN(n5445) );
  INV_X1 U6901 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7297) );
  INV_X1 U6902 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7301) );
  MUX2_X1 U6903 ( .A(n7297), .B(n7301), .S(n6553), .Z(n5429) );
  INV_X1 U6904 ( .A(SI_23_), .ZN(n5428) );
  NAND2_X1 U6905 ( .A1(n5429), .A2(n5428), .ZN(n5448) );
  INV_X1 U6906 ( .A(n5429), .ZN(n5430) );
  NAND2_X1 U6907 ( .A1(n5430), .A2(SI_23_), .ZN(n5431) );
  AND2_X1 U6908 ( .A1(n5448), .A2(n5431), .ZN(n5446) );
  NAND2_X1 U6909 ( .A1(n7298), .A2(n7963), .ZN(n5433) );
  OR2_X1 U6910 ( .A1(n4381), .A2(n7301), .ZN(n5432) );
  INV_X1 U6911 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5435) );
  INV_X1 U6912 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5434) );
  OAI21_X1 U6913 ( .B1(n5436), .B2(n5435), .A(n5434), .ZN(n5437) );
  AND2_X1 U6914 ( .A1(n5437), .A2(n5453), .ZN(n9148) );
  NAND2_X1 U6915 ( .A1(n9148), .A2(n5512), .ZN(n5443) );
  INV_X1 U6916 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U6917 ( .A1(n5666), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U6918 ( .A1(n5667), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5438) );
  OAI211_X1 U6919 ( .C1(n5561), .C2(n5440), .A(n5439), .B(n5438), .ZN(n5441)
         );
  INV_X1 U6920 ( .A(n5441), .ZN(n5442) );
  NAND2_X1 U6921 ( .A1(n5443), .A2(n5442), .ZN(n9218) );
  NAND2_X1 U6922 ( .A1(n9460), .A2(n9340), .ZN(n8178) );
  NAND2_X1 U6923 ( .A1(n8173), .A2(n8178), .ZN(n8260) );
  INV_X1 U6924 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7472) );
  INV_X1 U6925 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7470) );
  MUX2_X1 U6926 ( .A(n7472), .B(n7470), .S(n6553), .Z(n5463) );
  XNOR2_X1 U6927 ( .A(n5463), .B(SI_24_), .ZN(n5460) );
  XNOR2_X1 U6928 ( .A(n5462), .B(n5460), .ZN(n7469) );
  NAND2_X1 U6929 ( .A1(n7469), .A2(n7963), .ZN(n5451) );
  OR2_X1 U6930 ( .A1(n4380), .A2(n7470), .ZN(n5450) );
  INV_X1 U6931 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n10014) );
  NAND2_X1 U6932 ( .A1(n5453), .A2(n10014), .ZN(n5454) );
  NAND2_X1 U6933 ( .A1(n5475), .A2(n5454), .ZN(n9348) );
  OR2_X1 U6934 ( .A1(n9348), .A2(n5539), .ZN(n5459) );
  INV_X1 U6935 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5455) );
  INV_X1 U6936 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n10091) );
  OAI22_X1 U6937 ( .A1(n5077), .A2(n5455), .B1(n5561), .B2(n10091), .ZN(n5457)
         );
  INV_X1 U6938 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10145) );
  NOR2_X1 U6939 ( .A1(n4870), .A2(n10145), .ZN(n5456) );
  NOR2_X1 U6940 ( .A1(n5457), .A2(n5456), .ZN(n5458) );
  NAND2_X1 U6941 ( .A1(n5459), .A2(n5458), .ZN(n9321) );
  INV_X1 U6942 ( .A(n9321), .ZN(n7968) );
  XNOR2_X1 U6943 ( .A(n9344), .B(n7968), .ZN(n9336) );
  NAND2_X1 U6944 ( .A1(n9344), .A2(n7968), .ZN(n7970) );
  INV_X1 U6945 ( .A(n5460), .ZN(n5461) );
  INV_X1 U6946 ( .A(n5463), .ZN(n5464) );
  NAND2_X1 U6947 ( .A1(n5464), .A2(SI_24_), .ZN(n5465) );
  INV_X1 U6948 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7590) );
  INV_X1 U6949 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7593) );
  MUX2_X1 U6950 ( .A(n7590), .B(n7593), .S(n6553), .Z(n5468) );
  INV_X1 U6951 ( .A(SI_25_), .ZN(n5467) );
  NAND2_X1 U6952 ( .A1(n5468), .A2(n5467), .ZN(n5483) );
  INV_X1 U6953 ( .A(n5468), .ZN(n5469) );
  NAND2_X1 U6954 ( .A1(n5469), .A2(SI_25_), .ZN(n5470) );
  NAND2_X1 U6955 ( .A1(n5483), .A2(n5470), .ZN(n5484) );
  XNOR2_X1 U6956 ( .A(n5485), .B(n5484), .ZN(n7588) );
  NAND2_X1 U6957 ( .A1(n7588), .A2(n7963), .ZN(n5472) );
  OR2_X1 U6958 ( .A1(n4380), .A2(n7593), .ZN(n5471) );
  INV_X1 U6959 ( .A(n5475), .ZN(n5473) );
  NAND2_X1 U6960 ( .A1(n5473), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5492) );
  INV_X1 U6961 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U6962 ( .A1(n5475), .A2(n5474), .ZN(n5476) );
  NAND2_X1 U6963 ( .A1(n5492), .A2(n5476), .ZN(n9326) );
  OR2_X1 U6964 ( .A1(n9326), .A2(n5539), .ZN(n5481) );
  INV_X1 U6965 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9325) );
  NAND2_X1 U6966 ( .A1(n5666), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U6967 ( .A1(n5667), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5477) );
  OAI211_X1 U6968 ( .C1(n9325), .C2(n5561), .A(n5478), .B(n5477), .ZN(n5479)
         );
  INV_X1 U6969 ( .A(n5479), .ZN(n5480) );
  NAND2_X1 U6970 ( .A1(n5571), .A2(n9341), .ZN(n8061) );
  INV_X1 U6971 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n10190) );
  INV_X1 U6972 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7647) );
  MUX2_X1 U6973 ( .A(n10190), .B(n7647), .S(n6553), .Z(n5487) );
  INV_X1 U6974 ( .A(SI_26_), .ZN(n5486) );
  NAND2_X1 U6975 ( .A1(n5487), .A2(n5486), .ZN(n5514) );
  INV_X1 U6976 ( .A(n5487), .ZN(n5488) );
  NAND2_X1 U6977 ( .A1(n5488), .A2(SI_26_), .ZN(n5489) );
  AND2_X1 U6978 ( .A1(n5514), .A2(n5489), .ZN(n5500) );
  NAND2_X1 U6979 ( .A1(n7645), .A2(n7963), .ZN(n5491) );
  OR2_X1 U6980 ( .A1(n4380), .A2(n7647), .ZN(n5490) );
  INV_X1 U6981 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9978) );
  NAND2_X1 U6982 ( .A1(n5492), .A2(n9978), .ZN(n5493) );
  NAND2_X1 U6983 ( .A1(n9305), .A2(n5512), .ZN(n5499) );
  INV_X1 U6984 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U6985 ( .A1(n5667), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U6986 ( .A1(n5666), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5494) );
  OAI211_X1 U6987 ( .C1(n5496), .C2(n5561), .A(n5495), .B(n5494), .ZN(n5497)
         );
  INV_X1 U6988 ( .A(n5497), .ZN(n5498) );
  NAND2_X1 U6989 ( .A1(n9443), .A2(n9135), .ZN(n8186) );
  NAND2_X1 U6990 ( .A1(n9308), .A2(n9309), .ZN(n9314) );
  NAND2_X1 U6991 ( .A1(n9314), .A2(n8181), .ZN(n7949) );
  NAND2_X1 U6992 ( .A1(n5515), .A2(n5514), .ZN(n5506) );
  INV_X1 U6993 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7931) );
  INV_X1 U6994 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7710) );
  MUX2_X1 U6995 ( .A(n7931), .B(n7710), .S(n6553), .Z(n5503) );
  INV_X1 U6996 ( .A(SI_27_), .ZN(n5502) );
  NAND2_X1 U6997 ( .A1(n5503), .A2(n5502), .ZN(n5513) );
  INV_X1 U6998 ( .A(n5503), .ZN(n5504) );
  NAND2_X1 U6999 ( .A1(n5504), .A2(SI_27_), .ZN(n5516) );
  AND2_X1 U7000 ( .A1(n5513), .A2(n5516), .ZN(n5505) );
  OR2_X1 U7001 ( .A1(n4381), .A2(n7710), .ZN(n5507) );
  XNOR2_X1 U7002 ( .A(n5523), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9137) );
  INV_X1 U7003 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n10078) );
  NAND2_X1 U7004 ( .A1(n5667), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U7005 ( .A1(n5666), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5509) );
  OAI211_X1 U7006 ( .C1(n10078), .C2(n5561), .A(n5510), .B(n5509), .ZN(n5511)
         );
  NAND2_X1 U7007 ( .A1(n9438), .A2(n9312), .ZN(n8185) );
  NAND2_X1 U7008 ( .A1(n7949), .A2(n8121), .ZN(n7950) );
  INV_X1 U7009 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10188) );
  INV_X1 U7010 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7790) );
  MUX2_X1 U7011 ( .A(n10188), .B(n7790), .S(n6553), .Z(n5534) );
  XNOR2_X1 U7012 ( .A(n5534), .B(SI_28_), .ZN(n5531) );
  NAND2_X1 U7013 ( .A1(n7789), .A2(n7963), .ZN(n5519) );
  OR2_X1 U7014 ( .A1(n4381), .A2(n7790), .ZN(n5518) );
  INV_X1 U7015 ( .A(n5523), .ZN(n5521) );
  AND2_X1 U7016 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5520) );
  NAND2_X1 U7017 ( .A1(n5521), .A2(n5520), .ZN(n5587) );
  INV_X1 U7018 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9134) );
  INV_X1 U7019 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5522) );
  OAI21_X1 U7020 ( .B1(n5523), .B2(n9134), .A(n5522), .ZN(n5524) );
  NAND2_X1 U7021 ( .A1(n5587), .A2(n5524), .ZN(n9297) );
  OR2_X1 U7022 ( .A1(n9297), .A2(n5539), .ZN(n5530) );
  INV_X1 U7023 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U7024 ( .A1(n5666), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U7025 ( .A1(n5667), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5525) );
  OAI211_X1 U7026 ( .C1(n5527), .C2(n5561), .A(n5526), .B(n5525), .ZN(n5528)
         );
  INV_X1 U7027 ( .A(n5528), .ZN(n5529) );
  NAND2_X1 U7028 ( .A1(n9434), .A2(n9139), .ZN(n8184) );
  NAND3_X1 U7029 ( .A1(n7950), .A2(n9288), .A3(n8182), .ZN(n9287) );
  NAND2_X1 U7030 ( .A1(n9287), .A2(n8184), .ZN(n5546) );
  INV_X1 U7031 ( .A(SI_28_), .ZN(n5533) );
  NAND2_X1 U7032 ( .A1(n5534), .A2(n5533), .ZN(n5535) );
  INV_X1 U7033 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8289) );
  INV_X1 U7034 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7854) );
  MUX2_X1 U7035 ( .A(n8289), .B(n7854), .S(n6553), .Z(n5657) );
  XNOR2_X1 U7036 ( .A(n5657), .B(SI_29_), .ZN(n5536) );
  NAND2_X1 U7037 ( .A1(n8288), .A2(n7963), .ZN(n5538) );
  OR2_X1 U7038 ( .A1(n4380), .A2(n7854), .ZN(n5537) );
  OR2_X1 U7039 ( .A1(n5587), .A2(n5539), .ZN(n5545) );
  INV_X1 U7040 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U7041 ( .A1(n5666), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7042 ( .A1(n5667), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5540) );
  OAI211_X1 U7043 ( .C1(n5542), .C2(n5561), .A(n5541), .B(n5540), .ZN(n5543)
         );
  INV_X1 U7044 ( .A(n5543), .ZN(n5544) );
  NAND2_X1 U7045 ( .A1(n5545), .A2(n5544), .ZN(n9291) );
  XNOR2_X1 U7046 ( .A(n9431), .B(n9291), .ZN(n8122) );
  NAND2_X1 U7047 ( .A1(n5553), .A2(n5549), .ZN(n5550) );
  INV_X1 U7048 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U7049 ( .A1(n5653), .A2(n9349), .ZN(n5555) );
  NAND2_X1 U7050 ( .A1(n5652), .A2(n5611), .ZN(n5554) );
  NAND2_X1 U7051 ( .A1(n5555), .A2(n5554), .ZN(n9586) );
  INV_X1 U7052 ( .A(n9586), .ZN(n5556) );
  NAND2_X1 U7053 ( .A1(n5653), .A2(n5652), .ZN(n6499) );
  INV_X1 U7054 ( .A(n6499), .ZN(n8127) );
  INV_X1 U7055 ( .A(n4384), .ZN(n6525) );
  INV_X1 U7056 ( .A(n9419), .ZN(n5559) );
  INV_X1 U7057 ( .A(n9619), .ZN(n8248) );
  AND2_X1 U7058 ( .A1(n8248), .A2(P1_B_REG_SCAN_IN), .ZN(n5560) );
  NOR2_X1 U7059 ( .A1(n9577), .A2(n5560), .ZN(n5670) );
  INV_X1 U7060 ( .A(n5670), .ZN(n5566) );
  INV_X1 U7061 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7062 ( .A1(n5666), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5563) );
  INV_X1 U7063 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n7943) );
  OR2_X1 U7064 ( .A1(n5561), .A2(n7943), .ZN(n5562) );
  OAI211_X1 U7065 ( .C1(n4870), .C2(n5564), .A(n5563), .B(n5562), .ZN(n9215)
         );
  INV_X1 U7066 ( .A(n9215), .ZN(n5565) );
  NOR2_X1 U7067 ( .A1(n5566), .A2(n5565), .ZN(n5567) );
  NAND2_X1 U7068 ( .A1(n7218), .A2(n9801), .ZN(n7220) );
  INV_X1 U7069 ( .A(n7574), .ZN(n9564) );
  INV_X1 U7070 ( .A(n7516), .ZN(n9507) );
  NOR2_X2 U7071 ( .A1(n7746), .A2(n7751), .ZN(n7781) );
  INV_X1 U7072 ( .A(n9486), .ZN(n9411) );
  INV_X1 U7073 ( .A(n9480), .ZN(n9393) );
  NAND2_X1 U7074 ( .A1(n9302), .A2(n9307), .ZN(n9303) );
  INV_X1 U7075 ( .A(n9434), .ZN(n5572) );
  NAND2_X1 U7076 ( .A1(n8205), .A2(n8125), .ZN(n6672) );
  OR2_X1 U7077 ( .A1(n6672), .A2(n5611), .ZN(n9832) );
  NAND2_X1 U7078 ( .A1(n9430), .A2(n9778), .ZN(n5588) );
  OR2_X1 U7079 ( .A1(n8079), .A2(n5611), .ZN(n7016) );
  NAND2_X1 U7080 ( .A1(n5573), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U7081 ( .A1(n5580), .A2(n4971), .ZN(n5574) );
  NAND2_X1 U7082 ( .A1(n5574), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5575) );
  XNOR2_X1 U7083 ( .A(n5575), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U7084 ( .A1(n4398), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5576) );
  MUX2_X1 U7085 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5576), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5577) );
  INV_X1 U7086 ( .A(n5577), .ZN(n5579) );
  INV_X1 U7087 ( .A(n5573), .ZN(n5578) );
  NOR2_X1 U7088 ( .A1(n5579), .A2(n5578), .ZN(n5589) );
  XNOR2_X1 U7089 ( .A(n5580), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5607) );
  AND2_X1 U7090 ( .A1(n5589), .A2(n5607), .ZN(n5581) );
  NAND2_X1 U7091 ( .A1(n5582), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5583) );
  MUX2_X1 U7092 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5583), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n5584) );
  NAND2_X1 U7093 ( .A1(n5584), .A2(n4398), .ZN(n6498) );
  AND2_X1 U7094 ( .A1(n6498), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5585) );
  AND2_X1 U7095 ( .A1(n6478), .A2(n5585), .ZN(n9794) );
  AND2_X1 U7096 ( .A1(n9794), .A2(n8125), .ZN(n5586) );
  INV_X1 U7097 ( .A(n5607), .ZN(n7591) );
  INV_X1 U7098 ( .A(n5589), .ZN(n7471) );
  AND2_X1 U7099 ( .A1(n7471), .A2(P1_B_REG_SCAN_IN), .ZN(n5591) );
  NOR2_X1 U7100 ( .A1(n7471), .A2(P1_B_REG_SCAN_IN), .ZN(n5590) );
  AOI21_X1 U7101 ( .B1(n7591), .B2(n5591), .A(n5590), .ZN(n5592) );
  AND2_X1 U7102 ( .A1(n5592), .A2(n5608), .ZN(n6583) );
  INV_X1 U7103 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6587) );
  NAND2_X1 U7104 ( .A1(n6583), .A2(n6587), .ZN(n5593) );
  INV_X1 U7105 ( .A(n5608), .ZN(n7649) );
  NAND2_X1 U7106 ( .A1(n7649), .A2(n7471), .ZN(n6585) );
  NAND2_X1 U7107 ( .A1(n5593), .A2(n6585), .ZN(n5605) );
  NOR4_X1 U7108 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5597) );
  NOR4_X1 U7109 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n5596) );
  INV_X1 U7110 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10172) );
  INV_X1 U7111 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10062) );
  INV_X1 U7112 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10016) );
  INV_X1 U7113 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10162) );
  NAND4_X1 U7114 ( .A1(n10172), .A2(n10062), .A3(n10016), .A4(n10162), .ZN(
        n5594) );
  NOR2_X1 U7115 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n5594), .ZN(n10217) );
  NOR4_X1 U7116 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n5595) );
  NAND4_X1 U7117 ( .A1(n5597), .A2(n5596), .A3(n10217), .A4(n5595), .ZN(n5602)
         );
  NOR4_X1 U7118 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n5600) );
  NOR4_X1 U7119 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5599) );
  NOR4_X1 U7120 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5598) );
  INV_X1 U7121 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9788) );
  NAND4_X1 U7122 ( .A1(n5600), .A2(n5599), .A3(n5598), .A4(n9788), .ZN(n5601)
         );
  NOR2_X1 U7123 ( .A1(n5602), .A2(n5601), .ZN(n6466) );
  INV_X1 U7124 ( .A(n6466), .ZN(n5603) );
  NAND2_X1 U7125 ( .A1(n6583), .A2(n5603), .ZN(n5604) );
  NAND2_X1 U7126 ( .A1(n5605), .A2(n5604), .ZN(n5676) );
  INV_X1 U7127 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U7128 ( .A1(n6583), .A2(n5606), .ZN(n5610) );
  OR2_X1 U7129 ( .A1(n5608), .A2(n5607), .ZN(n5609) );
  NAND2_X1 U7130 ( .A1(n5610), .A2(n5609), .ZN(n9791) );
  NOR2_X1 U7131 ( .A1(n5676), .A2(n9791), .ZN(n5612) );
  AND2_X1 U7132 ( .A1(n5651), .A2(n9778), .ZN(n6248) );
  OR2_X1 U7133 ( .A1(n6499), .A2(n6248), .ZN(n6477) );
  NAND2_X1 U7134 ( .A1(n6477), .A2(n9794), .ZN(n5674) );
  INV_X1 U7135 ( .A(n5674), .ZN(n7001) );
  NAND2_X1 U7136 ( .A1(n5612), .A2(n7001), .ZN(n7189) );
  NAND2_X1 U7137 ( .A1(n5613), .A2(n9785), .ZN(n5656) );
  INV_X1 U7138 ( .A(n9344), .ZN(n9455) );
  AND2_X1 U7139 ( .A1(n9235), .A2(n7130), .ZN(n6884) );
  NAND2_X1 U7140 ( .A1(n6885), .A2(n6884), .ZN(n6886) );
  NAND2_X1 U7141 ( .A1(n6258), .A2(n6259), .ZN(n5614) );
  NAND2_X1 U7142 ( .A1(n6886), .A2(n5614), .ZN(n7198) );
  NAND2_X1 U7143 ( .A1(n5616), .A2(n5615), .ZN(n7196) );
  NAND2_X1 U7144 ( .A1(n6268), .A2(n9796), .ZN(n5617) );
  NAND2_X1 U7145 ( .A1(n7196), .A2(n5617), .ZN(n7213) );
  NAND2_X1 U7146 ( .A1(n7213), .A2(n8090), .ZN(n7212) );
  NAND2_X1 U7147 ( .A1(n7201), .A2(n9801), .ZN(n5618) );
  NAND2_X1 U7148 ( .A1(n7212), .A2(n5618), .ZN(n7178) );
  NAND2_X1 U7149 ( .A1(n8218), .A2(n8139), .ZN(n7180) );
  NAND2_X1 U7150 ( .A1(n7258), .A2(n7187), .ZN(n5619) );
  XNOR2_X1 U7151 ( .A(n9231), .B(n9773), .ZN(n7020) );
  NAND2_X1 U7152 ( .A1(n9231), .A2(n9773), .ZN(n5621) );
  NAND2_X1 U7153 ( .A1(n7978), .A2(n7990), .ZN(n8095) );
  NAND2_X1 U7154 ( .A1(n7432), .A2(n8095), .ZN(n7431) );
  NAND2_X1 U7155 ( .A1(n7022), .A2(n9812), .ZN(n5622) );
  NAND2_X1 U7156 ( .A1(n7431), .A2(n5622), .ZN(n7386) );
  INV_X1 U7157 ( .A(n7935), .ZN(n9226) );
  OR2_X1 U7158 ( .A1(n7574), .A2(n9226), .ZN(n5623) );
  OR2_X1 U7159 ( .A1(n9830), .A2(n9227), .ZN(n7561) );
  NAND2_X1 U7160 ( .A1(n5623), .A2(n7564), .ZN(n5626) );
  NOR2_X1 U7161 ( .A1(n8099), .A2(n5626), .ZN(n5624) );
  NAND2_X1 U7162 ( .A1(n7427), .A2(n9819), .ZN(n7402) );
  AND2_X1 U7163 ( .A1(n5624), .A2(n7402), .ZN(n5628) );
  NAND2_X1 U7164 ( .A1(n9228), .A2(n7410), .ZN(n7617) );
  NAND2_X1 U7165 ( .A1(n9830), .A2(n9227), .ZN(n5625) );
  AND2_X1 U7166 ( .A1(n7617), .A2(n5625), .ZN(n7560) );
  INV_X1 U7167 ( .A(n8101), .ZN(n7567) );
  AND2_X1 U7168 ( .A1(n7560), .A2(n7567), .ZN(n7563) );
  NOR2_X1 U7169 ( .A1(n5626), .A2(n7563), .ZN(n5627) );
  NAND2_X1 U7170 ( .A1(n8006), .A2(n8007), .ZN(n9580) );
  OR2_X1 U7171 ( .A1(n9501), .A2(n9223), .ZN(n5629) );
  INV_X1 U7172 ( .A(n5629), .ZN(n5632) );
  INV_X1 U7173 ( .A(n7551), .ZN(n9224) );
  NAND2_X1 U7174 ( .A1(n9593), .A2(n9224), .ZN(n7765) );
  NAND2_X1 U7175 ( .A1(n9501), .A2(n9223), .ZN(n5630) );
  AND2_X1 U7176 ( .A1(n7765), .A2(n5630), .ZN(n5631) );
  AND2_X1 U7177 ( .A1(n7751), .A2(n9222), .ZN(n5633) );
  NOR2_X1 U7178 ( .A1(n7778), .A2(n9221), .ZN(n5635) );
  NAND2_X1 U7179 ( .A1(n7778), .A2(n9221), .ZN(n5634) );
  NAND2_X1 U7180 ( .A1(n7855), .A2(n8021), .ZN(n5637) );
  INV_X1 U7181 ( .A(n7876), .ZN(n9220) );
  NAND2_X1 U7182 ( .A1(n9497), .A2(n9220), .ZN(n5636) );
  NAND2_X1 U7183 ( .A1(n5637), .A2(n5636), .ZN(n7867) );
  AND2_X1 U7184 ( .A1(n9490), .A2(n9420), .ZN(n5639) );
  OR2_X1 U7185 ( .A1(n9490), .A2(n9420), .ZN(n5638) );
  OAI21_X1 U7186 ( .B1(n7867), .B2(n5639), .A(n5638), .ZN(n9403) );
  INV_X1 U7187 ( .A(n7909), .ZN(n9397) );
  NAND2_X1 U7188 ( .A1(n9486), .A2(n9397), .ZN(n5640) );
  OR2_X1 U7189 ( .A1(n9480), .A2(n9418), .ZN(n5641) );
  OR2_X1 U7190 ( .A1(n9476), .A2(n9396), .ZN(n5642) );
  NAND2_X1 U7191 ( .A1(n9371), .A2(n5642), .ZN(n9355) );
  NAND2_X1 U7192 ( .A1(n9476), .A2(n9396), .ZN(n9354) );
  NAND2_X1 U7193 ( .A1(n9471), .A2(n9219), .ZN(n5643) );
  AND2_X1 U7194 ( .A1(n9354), .A2(n5643), .ZN(n5645) );
  INV_X1 U7195 ( .A(n5643), .ZN(n5644) );
  AND2_X1 U7196 ( .A1(n9465), .A2(n9366), .ZN(n5646) );
  NOR2_X1 U7197 ( .A1(n9460), .A2(n9218), .ZN(n5647) );
  NAND2_X1 U7198 ( .A1(n9460), .A2(n9218), .ZN(n8049) );
  OAI21_X1 U7199 ( .B1(n9324), .B2(n9323), .A(n5648), .ZN(n9301) );
  NAND2_X1 U7200 ( .A1(n9443), .A2(n9320), .ZN(n5649) );
  INV_X1 U7201 ( .A(n9312), .ZN(n9216) );
  XNOR2_X1 U7202 ( .A(n5650), .B(n8122), .ZN(n9432) );
  OR2_X1 U7203 ( .A1(n6249), .A2(n6891), .ZN(n6668) );
  AND2_X1 U7204 ( .A1(n6668), .A2(n6452), .ZN(n9771) );
  NAND2_X1 U7205 ( .A1(n9785), .A2(n9771), .ZN(n9425) );
  OR2_X1 U7206 ( .A1(n6672), .A2(n5651), .ZN(n6474) );
  INV_X1 U7207 ( .A(n6474), .ZN(n9772) );
  INV_X2 U7208 ( .A(n9785), .ZN(n9787) );
  AOI22_X1 U7209 ( .A1(n9431), .A2(n9590), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9787), .ZN(n5654) );
  NAND2_X1 U7210 ( .A1(n5656), .A2(n4417), .ZN(P1_U3355) );
  INV_X1 U7211 ( .A(n5657), .ZN(n5658) );
  NOR2_X1 U7212 ( .A1(n5658), .A2(SI_29_), .ZN(n5659) );
  MUX2_X1 U7213 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n6553), .Z(n7956) );
  NAND2_X1 U7214 ( .A1(n8293), .A2(n7963), .ZN(n5662) );
  INV_X1 U7215 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7921) );
  OR2_X1 U7216 ( .A1(n4381), .A2(n7921), .ZN(n5661) );
  INV_X1 U7217 ( .A(n8088), .ZN(n5664) );
  NAND2_X1 U7218 ( .A1(n5664), .A2(n5663), .ZN(n9276) );
  OAI21_X1 U7219 ( .B1(n5664), .B2(n5663), .A(n9276), .ZN(n7946) );
  NOR2_X1 U7220 ( .A1(n7946), .A2(n9832), .ZN(n5673) );
  OR2_X1 U7221 ( .A1(n6672), .A2(n9778), .ZN(n5665) );
  INV_X1 U7222 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9277) );
  NAND2_X1 U7223 ( .A1(n5666), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U7224 ( .A1(n5667), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5668) );
  OAI211_X1 U7225 ( .C1(n5561), .C2(n9277), .A(n5669), .B(n5668), .ZN(n8072)
         );
  NAND2_X1 U7226 ( .A1(n8072), .A2(n5670), .ZN(n9428) );
  OAI21_X1 U7227 ( .B1(n7016), .B2(n5652), .A(n9791), .ZN(n5675) );
  OR2_X1 U7228 ( .A1(n5675), .A2(n5674), .ZN(n6883) );
  INV_X2 U7229 ( .A(n9838), .ZN(n9840) );
  INV_X1 U7230 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5718) );
  INV_X1 U7231 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5678) );
  NOR2_X1 U7232 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5680) );
  NOR2_X1 U7233 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5679) );
  INV_X1 U7234 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5683) );
  INV_X1 U7235 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5731) );
  INV_X1 U7236 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9124) );
  XNOR2_X2 U7237 ( .A(n5692), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5698) );
  INV_X1 U7238 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5693) );
  INV_X1 U7239 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7248) );
  NAND2_X2 U7240 ( .A1(n5694), .A2(n7788), .ZN(n5767) );
  INV_X1 U7241 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9855) );
  OR2_X1 U7242 ( .A1(n5767), .A2(n9855), .ZN(n5695) );
  NAND3_X1 U7243 ( .A1(n5697), .A2(n5696), .A3(n5695), .ZN(n5701) );
  INV_X1 U7244 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5699) );
  INV_X1 U7245 ( .A(SI_0_), .ZN(n5703) );
  INV_X1 U7246 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5702) );
  OAI21_X1 U7247 ( .B1(n6553), .B2(n5703), .A(n5702), .ZN(n5704) );
  AND2_X1 U7248 ( .A1(n5705), .A2(n5704), .ZN(n9129) );
  INV_X1 U7249 ( .A(n5707), .ZN(n5708) );
  NOR2_X1 U7250 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(n5708), .ZN(n5709) );
  XNOR2_X1 U7251 ( .A(n5710), .B(n5688), .ZN(n6715) );
  INV_X1 U7252 ( .A(n8507), .ZN(n9872) );
  INV_X1 U7253 ( .A(n7121), .ZN(n5733) );
  NAND2_X1 U7254 ( .A1(n5882), .A2(n5715), .ZN(n5890) );
  INV_X1 U7255 ( .A(n5890), .ZN(n5717) );
  NAND2_X1 U7256 ( .A1(n5717), .A2(n5716), .ZN(n5916) );
  INV_X1 U7257 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5951) );
  AND3_X1 U7258 ( .A1(n5951), .A2(n5948), .A3(n5718), .ZN(n5719) );
  NAND2_X1 U7259 ( .A1(n6020), .A2(n5721), .ZN(n5722) );
  INV_X1 U7260 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U7261 ( .A1(n5726), .A2(n5725), .ZN(n5727) );
  INV_X1 U7262 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5723) );
  AND2_X1 U7263 ( .A1(n6215), .A2(n8855), .ZN(n6226) );
  NAND2_X1 U7264 ( .A1(n6181), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5730) );
  INV_X1 U7265 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5729) );
  XNOR2_X1 U7266 ( .A(n5730), .B(n5729), .ZN(n8340) );
  OR2_X1 U7267 ( .A1(n4395), .A2(n5970), .ZN(n5732) );
  XNOR2_X1 U7268 ( .A(n5732), .B(n5731), .ZN(n8338) );
  NAND2_X1 U7269 ( .A1(n8340), .A2(n8338), .ZN(n9873) );
  INV_X1 U7270 ( .A(n9873), .ZN(n6856) );
  NAND2_X1 U7271 ( .A1(n5733), .A2(n5792), .ZN(n8506) );
  INV_X1 U7272 ( .A(n8340), .ZN(n8501) );
  NAND2_X1 U7273 ( .A1(n9873), .A2(n8338), .ZN(n5734) );
  INV_X1 U7274 ( .A(n8338), .ZN(n8351) );
  NAND2_X1 U7275 ( .A1(n6215), .A2(n8351), .ZN(n7053) );
  OAI21_X2 U7276 ( .B1(n8337), .B2(n5734), .A(n7053), .ZN(n5747) );
  INV_X1 U7277 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7118) );
  OR2_X1 U7278 ( .A1(n5767), .A2(n7118), .ZN(n5740) );
  INV_X1 U7279 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7117) );
  INV_X1 U7280 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6726) );
  OR2_X1 U7281 ( .A1(n5753), .A2(n6726), .ZN(n5738) );
  NAND2_X1 U7282 ( .A1(n5783), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5737) );
  NAND4_X1 U7283 ( .A1(n5740), .A2(n5739), .A3(n5738), .A4(n5737), .ZN(n6922)
         );
  INV_X1 U7284 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6556) );
  NAND2_X2 U7285 ( .A1(n5773), .A2(n5741), .ZN(n5794) );
  NAND2_X1 U7286 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5742) );
  MUX2_X1 U7287 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5742), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5744) );
  INV_X1 U7288 ( .A(n5796), .ZN(n5743) );
  XNOR2_X1 U7289 ( .A(n5750), .B(n5748), .ZN(n8546) );
  NAND2_X1 U7290 ( .A1(n8547), .A2(n8546), .ZN(n8545) );
  INV_X1 U7291 ( .A(n5748), .ZN(n5749) );
  NAND2_X1 U7292 ( .A1(n5750), .A2(n5749), .ZN(n5751) );
  INV_X1 U7293 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5752) );
  OR2_X1 U7294 ( .A1(n5767), .A2(n5752), .ZN(n5758) );
  INV_X1 U7295 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6725) );
  OR2_X1 U7296 ( .A1(n5753), .A2(n6725), .ZN(n5757) );
  INV_X1 U7297 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U7298 ( .A1(n5783), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5755) );
  NOR2_X1 U7299 ( .A1(n4953), .A2(n5771), .ZN(n5763) );
  OR2_X1 U7300 ( .A1(n5796), .A2(n5970), .ZN(n5759) );
  XNOR2_X1 U7301 ( .A(n5759), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9554) );
  INV_X1 U7302 ( .A(n9554), .ZN(n6728) );
  OR2_X1 U7303 ( .A1(n5793), .A2(n6570), .ZN(n5761) );
  OR2_X1 U7304 ( .A1(n5794), .A2(n6569), .ZN(n5760) );
  OAI211_X1 U7305 ( .C1(n6713), .C2(n6728), .A(n5761), .B(n5760), .ZN(n6836)
         );
  INV_X1 U7306 ( .A(n6836), .ZN(n9885) );
  INV_X1 U7307 ( .A(n9885), .ZN(n7239) );
  XNOR2_X1 U7308 ( .A(n7239), .B(n5747), .ZN(n5762) );
  NAND2_X1 U7309 ( .A1(n5763), .A2(n5762), .ZN(n5765) );
  NAND2_X1 U7310 ( .A1(n5783), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5770) );
  INV_X1 U7311 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6724) );
  OR2_X1 U7312 ( .A1(n5753), .A2(n6724), .ZN(n5769) );
  OR2_X1 U7313 ( .A1(n5766), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5768) );
  INV_X1 U7314 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7060) );
  CLKBUF_X3 U7315 ( .A(n5771), .Z(n8504) );
  OR2_X1 U7316 ( .A1(n7144), .A2(n8504), .ZN(n5779) );
  NAND2_X1 U7317 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4408), .ZN(n5772) );
  XNOR2_X1 U7318 ( .A(n5772), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6723) );
  INV_X1 U7319 ( .A(n6723), .ZN(n6750) );
  NOR2_X1 U7320 ( .A1(n5773), .A2(n6750), .ZN(n5774) );
  OR2_X1 U7321 ( .A1(n5793), .A2(n6557), .ZN(n5776) );
  XNOR2_X1 U7322 ( .A(n7071), .B(n5747), .ZN(n5780) );
  XNOR2_X1 U7323 ( .A(n5779), .B(n5780), .ZN(n7069) );
  NAND2_X1 U7324 ( .A1(n7070), .A2(n7069), .ZN(n7068) );
  INV_X1 U7325 ( .A(n5779), .ZN(n5781) );
  NAND2_X1 U7326 ( .A1(n5781), .A2(n5780), .ZN(n5782) );
  NAND2_X1 U7327 ( .A1(n7068), .A2(n5782), .ZN(n6933) );
  NAND2_X1 U7328 ( .A1(n5783), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5791) );
  INV_X1 U7329 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6722) );
  OR2_X1 U7330 ( .A1(n5753), .A2(n6722), .ZN(n5790) );
  INV_X1 U7331 ( .A(n5811), .ZN(n5787) );
  INV_X1 U7332 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5785) );
  INV_X1 U7333 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5784) );
  NAND2_X1 U7334 ( .A1(n5785), .A2(n5784), .ZN(n5786) );
  NAND2_X1 U7335 ( .A1(n5787), .A2(n5786), .ZN(n7150) );
  OR2_X1 U7336 ( .A1(n5766), .A2(n7150), .ZN(n5789) );
  INV_X1 U7337 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7151) );
  OR2_X1 U7338 ( .A1(n5767), .A2(n7151), .ZN(n5788) );
  NAND4_X1 U7339 ( .A1(n5791), .A2(n5790), .A3(n5789), .A4(n5788), .ZN(n8662)
         );
  AND2_X1 U7340 ( .A1(n8662), .A2(n5792), .ZN(n5802) );
  OR2_X1 U7341 ( .A1(n8300), .A2(n10257), .ZN(n5800) );
  NAND2_X1 U7342 ( .A1(n5796), .A2(n5795), .ZN(n5829) );
  NAND2_X1 U7343 ( .A1(n5829), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5797) );
  XNOR2_X1 U7344 ( .A(n5797), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6721) );
  INV_X1 U7345 ( .A(n6721), .ZN(n10254) );
  OR2_X1 U7346 ( .A1(n6713), .A2(n10254), .ZN(n5798) );
  XNOR2_X1 U7347 ( .A(n7152), .B(n6155), .ZN(n5801) );
  AND2_X1 U7348 ( .A1(n5802), .A2(n5801), .ZN(n6930) );
  INV_X1 U7349 ( .A(n5801), .ZN(n5804) );
  INV_X1 U7350 ( .A(n5802), .ZN(n5803) );
  NAND2_X1 U7351 ( .A1(n5804), .A2(n5803), .ZN(n6929) );
  OAI21_X2 U7352 ( .B1(n6933), .B2(n6930), .A(n6929), .ZN(n8582) );
  INV_X1 U7353 ( .A(n8582), .ZN(n5816) );
  INV_X1 U7354 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6568) );
  OR2_X1 U7355 ( .A1(n8300), .A2(n6568), .ZN(n5809) );
  OR2_X1 U7356 ( .A1(n5794), .A2(n6567), .ZN(n5808) );
  OR2_X1 U7357 ( .A1(n5829), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U7358 ( .A1(n5805), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5806) );
  XNOR2_X1 U7359 ( .A(n5806), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6769) );
  INV_X1 U7360 ( .A(n6769), .ZN(n6738) );
  OR2_X1 U7361 ( .A1(n6713), .A2(n6738), .ZN(n5807) );
  XNOR2_X1 U7362 ( .A(n7325), .B(n6177), .ZN(n5818) );
  NAND2_X1 U7363 ( .A1(n5783), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5814) );
  INV_X1 U7364 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5810) );
  INV_X1 U7365 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6731) );
  OR2_X1 U7366 ( .A1(n5753), .A2(n6731), .ZN(n5813) );
  OAI21_X1 U7367 ( .B1(n5811), .B2(P2_REG3_REG_5__SCAN_IN), .A(n5849), .ZN(
        n7323) );
  OR2_X1 U7368 ( .A1(n5766), .A2(n7323), .ZN(n5812) );
  NAND2_X1 U7369 ( .A1(n8661), .A2(n5792), .ZN(n5817) );
  XNOR2_X1 U7370 ( .A(n5818), .B(n5817), .ZN(n8581) );
  INV_X1 U7371 ( .A(n8581), .ZN(n5815) );
  NAND2_X1 U7372 ( .A1(n5816), .A2(n5815), .ZN(n5822) );
  INV_X1 U7373 ( .A(n5817), .ZN(n5820) );
  INV_X1 U7374 ( .A(n5818), .ZN(n5819) );
  NAND2_X1 U7375 ( .A1(n5820), .A2(n5819), .ZN(n5821) );
  NAND2_X1 U7376 ( .A1(n5822), .A2(n5821), .ZN(n7105) );
  INV_X1 U7377 ( .A(n5767), .ZN(n6594) );
  NAND2_X1 U7378 ( .A1(n6594), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5828) );
  INV_X1 U7379 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6787) );
  OR2_X1 U7380 ( .A1(n5753), .A2(n6787), .ZN(n5827) );
  INV_X1 U7381 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5823) );
  XNOR2_X1 U7382 ( .A(n5849), .B(n5823), .ZN(n7107) );
  OR2_X1 U7383 ( .A1(n5766), .A2(n7107), .ZN(n5826) );
  INV_X1 U7384 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5824) );
  OR2_X1 U7385 ( .A1(n6609), .A2(n5824), .ZN(n5825) );
  OR2_X1 U7386 ( .A1(n6945), .A2(n8504), .ZN(n5839) );
  INV_X1 U7387 ( .A(n5829), .ZN(n5830) );
  AND2_X1 U7388 ( .A1(n5831), .A2(n5830), .ZN(n5832) );
  OR2_X1 U7389 ( .A1(n5832), .A2(n5970), .ZN(n5834) );
  XNOR2_X1 U7390 ( .A(n5834), .B(n5833), .ZN(n6786) );
  OR2_X1 U7391 ( .A1(n8300), .A2(n6571), .ZN(n5836) );
  XNOR2_X1 U7392 ( .A(n6155), .B(n7273), .ZN(n5838) );
  NAND2_X1 U7393 ( .A1(n5839), .A2(n5838), .ZN(n5840) );
  OAI21_X1 U7394 ( .B1(n5839), .B2(n5838), .A(n5840), .ZN(n7106) );
  NAND2_X1 U7395 ( .A1(n7103), .A2(n5840), .ZN(n7134) );
  OR2_X1 U7396 ( .A1(n5794), .A2(n6572), .ZN(n5845) );
  OR2_X1 U7397 ( .A1(n8300), .A2(n6573), .ZN(n5844) );
  NAND2_X1 U7398 ( .A1(n5841), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5842) );
  XNOR2_X1 U7399 ( .A(n5842), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6783) );
  INV_X1 U7400 ( .A(n6783), .ZN(n6803) );
  OR2_X1 U7401 ( .A1(n6713), .A2(n6803), .ZN(n5843) );
  XNOR2_X1 U7402 ( .A(n7316), .B(n6177), .ZN(n5856) );
  NAND2_X1 U7403 ( .A1(n5783), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5854) );
  INV_X1 U7404 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6784) );
  OR2_X1 U7405 ( .A1(n5753), .A2(n6784), .ZN(n5853) );
  INV_X1 U7406 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5846) );
  OR2_X1 U7407 ( .A1(n6606), .A2(n5846), .ZN(n5852) );
  INV_X1 U7408 ( .A(n5849), .ZN(n5847) );
  AOI21_X1 U7409 ( .B1(n5847), .B2(P2_REG3_REG_6__SCAN_IN), .A(
        P2_REG3_REG_7__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U7410 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5848) );
  OR2_X1 U7411 ( .A1(n5850), .A2(n5858), .ZN(n7313) );
  OR2_X1 U7412 ( .A1(n5766), .A2(n7313), .ZN(n5851) );
  NAND4_X1 U7413 ( .A1(n5854), .A2(n5853), .A3(n5852), .A4(n5851), .ZN(n8659)
         );
  NAND2_X1 U7414 ( .A1(n8659), .A2(n5792), .ZN(n5855) );
  XNOR2_X1 U7415 ( .A(n5856), .B(n5855), .ZN(n7133) );
  OAI22_X1 U7416 ( .A1(n7134), .A2(n7133), .B1(n5856), .B2(n5855), .ZN(n8535)
         );
  NAND2_X1 U7417 ( .A1(n6234), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5863) );
  INV_X1 U7418 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5857) );
  OR2_X1 U7419 ( .A1(n6609), .A2(n5857), .ZN(n5862) );
  NAND2_X1 U7420 ( .A1(n5858), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5875) );
  OR2_X1 U7421 ( .A1(n5858), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U7422 ( .A1(n5875), .A2(n5859), .ZN(n8538) );
  OR2_X1 U7423 ( .A1(n5766), .A2(n8538), .ZN(n5861) );
  INV_X1 U7424 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7096) );
  OR2_X1 U7425 ( .A1(n6606), .A2(n7096), .ZN(n5860) );
  OR2_X1 U7426 ( .A1(n7482), .A2(n8504), .ZN(n5868) );
  NAND2_X1 U7427 ( .A1(n5864), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5865) );
  XNOR2_X1 U7428 ( .A(n5865), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6904) );
  INV_X1 U7429 ( .A(n6904), .ZN(n6910) );
  OR2_X1 U7430 ( .A1(n5794), .A2(n6564), .ZN(n5867) );
  OR2_X1 U7431 ( .A1(n8300), .A2(n6554), .ZN(n5866) );
  OAI211_X1 U7432 ( .C1(n6713), .C2(n6910), .A(n5867), .B(n5866), .ZN(n8540)
         );
  XNOR2_X1 U7433 ( .A(n8540), .B(n6177), .ZN(n5869) );
  XNOR2_X1 U7434 ( .A(n5868), .B(n5869), .ZN(n8534) );
  NAND2_X1 U7435 ( .A1(n8535), .A2(n8534), .ZN(n5872) );
  INV_X1 U7436 ( .A(n5868), .ZN(n5870) );
  NAND2_X1 U7437 ( .A1(n5870), .A2(n5869), .ZN(n5871) );
  NAND2_X1 U7438 ( .A1(n5872), .A2(n5871), .ZN(n7475) );
  NAND2_X1 U7439 ( .A1(n6234), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5881) );
  INV_X1 U7440 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5873) );
  OR2_X1 U7441 ( .A1(n6606), .A2(n5873), .ZN(n5880) );
  INV_X1 U7442 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7443 ( .A1(n5875), .A2(n5874), .ZN(n5876) );
  NAND2_X1 U7444 ( .A1(n5893), .A2(n5876), .ZN(n7481) );
  OR2_X1 U7445 ( .A1(n5766), .A2(n7481), .ZN(n5879) );
  INV_X1 U7446 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5877) );
  OR2_X1 U7447 ( .A1(n6609), .A2(n5877), .ZN(n5878) );
  OR2_X1 U7448 ( .A1(n7286), .A2(n8504), .ZN(n5888) );
  INV_X1 U7449 ( .A(n5882), .ZN(n5883) );
  NAND2_X1 U7450 ( .A1(n5883), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5884) );
  XNOR2_X1 U7451 ( .A(n5884), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6984) );
  INV_X1 U7452 ( .A(n6984), .ZN(n6991) );
  OR2_X1 U7453 ( .A1(n5794), .A2(n6574), .ZN(n5886) );
  OR2_X1 U7454 ( .A1(n8300), .A2(n6575), .ZN(n5885) );
  OAI211_X1 U7455 ( .C1(n6713), .C2(n6991), .A(n5886), .B(n5885), .ZN(n9099)
         );
  XNOR2_X1 U7456 ( .A(n6155), .B(n9099), .ZN(n5887) );
  NAND2_X1 U7457 ( .A1(n5888), .A2(n5887), .ZN(n5889) );
  OAI21_X1 U7458 ( .B1(n5888), .B2(n5887), .A(n5889), .ZN(n7478) );
  NAND2_X1 U7459 ( .A1(n5890), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5902) );
  XNOR2_X1 U7460 ( .A(n5902), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7451) );
  AOI22_X1 U7461 ( .A1(n6036), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6590), .B2(
        n7451), .ZN(n5892) );
  NAND2_X1 U7462 ( .A1(n6578), .A2(n8299), .ZN(n5891) );
  XNOR2_X1 U7463 ( .A(n9917), .B(n6177), .ZN(n5900) );
  NAND2_X1 U7464 ( .A1(n5783), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5898) );
  INV_X1 U7465 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6992) );
  OR2_X1 U7466 ( .A1(n5753), .A2(n6992), .ZN(n5897) );
  INV_X1 U7467 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7290) );
  OR2_X1 U7468 ( .A1(n6606), .A2(n7290), .ZN(n5896) );
  INV_X1 U7469 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10187) );
  AND2_X1 U7470 ( .A1(n5893), .A2(n10187), .ZN(n5894) );
  OR2_X1 U7471 ( .A1(n5894), .A2(n5921), .ZN(n7610) );
  OR2_X1 U7472 ( .A1(n5766), .A2(n7610), .ZN(n5895) );
  NAND4_X1 U7473 ( .A1(n5898), .A2(n5897), .A3(n5896), .A4(n5895), .ZN(n8656)
         );
  NAND2_X1 U7474 ( .A1(n8656), .A2(n5792), .ZN(n5899) );
  XNOR2_X1 U7475 ( .A(n5900), .B(n5899), .ZN(n7609) );
  NAND2_X1 U7476 ( .A1(n6576), .A2(n8299), .ZN(n5906) );
  INV_X1 U7477 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U7478 ( .A1(n5902), .A2(n5901), .ZN(n5903) );
  NAND2_X1 U7479 ( .A1(n5903), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5904) );
  XNOR2_X1 U7480 ( .A(n5904), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8672) );
  AOI22_X1 U7481 ( .A1(n6036), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6590), .B2(
        n8672), .ZN(n5905) );
  NAND2_X1 U7482 ( .A1(n5906), .A2(n5905), .ZN(n9094) );
  XNOR2_X1 U7483 ( .A(n9094), .B(n6177), .ZN(n5912) );
  NAND2_X1 U7484 ( .A1(n5783), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5910) );
  INV_X1 U7485 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7457) );
  OR2_X1 U7486 ( .A1(n5753), .A2(n7457), .ZN(n5909) );
  XNOR2_X1 U7487 ( .A(n5921), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n8625) );
  OR2_X1 U7488 ( .A1(n5766), .A2(n8625), .ZN(n5908) );
  INV_X1 U7489 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7349) );
  OR2_X1 U7490 ( .A1(n6606), .A2(n7349), .ZN(n5907) );
  OR2_X1 U7491 ( .A1(n7671), .A2(n8504), .ZN(n5911) );
  XNOR2_X1 U7492 ( .A(n5912), .B(n5911), .ZN(n8620) );
  INV_X1 U7493 ( .A(n5911), .ZN(n5913) );
  NAND2_X1 U7494 ( .A1(n5913), .A2(n5912), .ZN(n5914) );
  NAND2_X1 U7495 ( .A1(n5915), .A2(n5914), .ZN(n7667) );
  NAND2_X1 U7496 ( .A1(n6599), .A2(n8299), .ZN(n5919) );
  NAND2_X1 U7497 ( .A1(n5916), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5917) );
  XNOR2_X1 U7498 ( .A(n5917), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7599) );
  AOI22_X1 U7499 ( .A1(n6036), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6590), .B2(
        n7599), .ZN(n5918) );
  XNOR2_X1 U7500 ( .A(n9924), .B(n6155), .ZN(n5927) );
  NAND2_X1 U7501 ( .A1(n5783), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5926) );
  INV_X1 U7502 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7377) );
  OR2_X1 U7503 ( .A1(n6606), .A2(n7377), .ZN(n5925) );
  INV_X1 U7504 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7456) );
  OR2_X1 U7505 ( .A1(n5753), .A2(n7456), .ZN(n5924) );
  AND2_X1 U7506 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n5920) );
  AOI21_X1 U7507 ( .B1(n5921), .B2(P2_REG3_REG_11__SCAN_IN), .A(
        P2_REG3_REG_12__SCAN_IN), .ZN(n5922) );
  OR2_X1 U7508 ( .A1(n5936), .A2(n5922), .ZN(n7670) );
  OR2_X1 U7509 ( .A1(n5766), .A2(n7670), .ZN(n5923) );
  OR2_X1 U7510 ( .A1(n7715), .A2(n8504), .ZN(n5928) );
  NAND2_X1 U7511 ( .A1(n5927), .A2(n5928), .ZN(n7665) );
  NAND2_X1 U7512 ( .A1(n7667), .A2(n7665), .ZN(n5931) );
  INV_X1 U7513 ( .A(n5927), .ZN(n5930) );
  INV_X1 U7514 ( .A(n5928), .ZN(n5929) );
  NAND2_X1 U7515 ( .A1(n5930), .A2(n5929), .ZN(n7666) );
  NAND2_X1 U7516 ( .A1(n5931), .A2(n7666), .ZN(n7713) );
  NAND2_X1 U7517 ( .A1(n6614), .A2(n8299), .ZN(n5934) );
  OR2_X1 U7518 ( .A1(n5932), .A2(n5970), .ZN(n5949) );
  XNOR2_X1 U7519 ( .A(n5949), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7655) );
  AOI22_X1 U7520 ( .A1(n6036), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6590), .B2(
        n7655), .ZN(n5933) );
  XNOR2_X1 U7521 ( .A(n9089), .B(n6177), .ZN(n5942) );
  NAND2_X1 U7522 ( .A1(n5783), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5941) );
  INV_X1 U7523 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7499) );
  OR2_X1 U7524 ( .A1(n6606), .A2(n7499), .ZN(n5940) );
  INV_X1 U7525 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5935) );
  OR2_X1 U7526 ( .A1(n5753), .A2(n5935), .ZN(n5939) );
  OR2_X1 U7527 ( .A1(n5936), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U7528 ( .A1(n5958), .A2(n5937), .ZN(n7714) );
  OR2_X1 U7529 ( .A1(n5766), .A2(n7714), .ZN(n5938) );
  NOR2_X1 U7530 ( .A1(n7838), .A2(n8504), .ZN(n5943) );
  NAND2_X1 U7531 ( .A1(n5942), .A2(n5943), .ZN(n5947) );
  INV_X1 U7532 ( .A(n5942), .ZN(n5945) );
  INV_X1 U7533 ( .A(n5943), .ZN(n5944) );
  NAND2_X1 U7534 ( .A1(n5945), .A2(n5944), .ZN(n5946) );
  AND2_X1 U7535 ( .A1(n5947), .A2(n5946), .ZN(n7712) );
  NAND2_X1 U7536 ( .A1(n6617), .A2(n8299), .ZN(n5955) );
  NAND2_X1 U7537 ( .A1(n5949), .A2(n5948), .ZN(n5950) );
  NAND2_X1 U7538 ( .A1(n5950), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5952) );
  OR2_X1 U7539 ( .A1(n5952), .A2(n5951), .ZN(n5953) );
  NAND2_X1 U7540 ( .A1(n5952), .A2(n5951), .ZN(n5991) );
  AND2_X1 U7541 ( .A1(n5953), .A2(n5991), .ZN(n8681) );
  AOI22_X1 U7542 ( .A1(n6036), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6590), .B2(
        n8681), .ZN(n5954) );
  XNOR2_X1 U7543 ( .A(n7841), .B(n6177), .ZN(n5965) );
  NAND2_X1 U7544 ( .A1(n5783), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5963) );
  INV_X1 U7545 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5956) );
  OR2_X1 U7546 ( .A1(n5753), .A2(n5956), .ZN(n5962) );
  INV_X1 U7547 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U7548 ( .A1(n5958), .A2(n5957), .ZN(n5959) );
  NAND2_X1 U7549 ( .A1(n5984), .A2(n5959), .ZN(n7837) );
  OR2_X1 U7550 ( .A1(n5766), .A2(n7837), .ZN(n5961) );
  INV_X1 U7551 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7541) );
  OR2_X1 U7552 ( .A1(n6606), .A2(n7541), .ZN(n5960) );
  NOR2_X1 U7553 ( .A1(n7898), .A2(n8504), .ZN(n5966) );
  XNOR2_X1 U7554 ( .A(n5965), .B(n5966), .ZN(n7835) );
  INV_X1 U7555 ( .A(n5965), .ZN(n5968) );
  INV_X1 U7556 ( .A(n5966), .ZN(n5967) );
  NAND2_X1 U7557 ( .A1(n5968), .A2(n5967), .ZN(n5969) );
  NAND2_X1 U7558 ( .A1(n7832), .A2(n5969), .ZN(n7893) );
  NAND2_X1 U7559 ( .A1(n6624), .A2(n8299), .ZN(n5974) );
  OR2_X1 U7560 ( .A1(n5971), .A2(n5970), .ZN(n5972) );
  XNOR2_X1 U7561 ( .A(n5972), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8718) );
  AOI22_X1 U7562 ( .A1(n6036), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6590), .B2(
        n8718), .ZN(n5973) );
  XNOR2_X1 U7563 ( .A(n9083), .B(n6177), .ZN(n8572) );
  NAND2_X1 U7564 ( .A1(n5783), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5981) );
  INV_X1 U7565 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7801) );
  OR2_X1 U7566 ( .A1(n6606), .A2(n7801), .ZN(n5980) );
  INV_X1 U7567 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n5975) );
  OR2_X1 U7568 ( .A1(n5753), .A2(n5975), .ZN(n5979) );
  INV_X1 U7569 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5983) );
  INV_X1 U7570 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10210) );
  NAND2_X1 U7571 ( .A1(n5986), .A2(n10210), .ZN(n5977) );
  INV_X1 U7572 ( .A(n6007), .ZN(n5976) );
  NAND2_X1 U7573 ( .A1(n5977), .A2(n5976), .ZN(n8575) );
  OR2_X1 U7574 ( .A1(n5766), .A2(n8575), .ZN(n5978) );
  NOR2_X1 U7575 ( .A1(n7896), .A2(n8504), .ZN(n5997) );
  NAND2_X1 U7576 ( .A1(n5783), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5990) );
  INV_X1 U7577 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7639) );
  OR2_X1 U7578 ( .A1(n5767), .A2(n7639), .ZN(n5989) );
  INV_X1 U7579 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5982) );
  OR2_X1 U7580 ( .A1(n5753), .A2(n5982), .ZN(n5988) );
  NAND2_X1 U7581 ( .A1(n5984), .A2(n5983), .ZN(n5985) );
  NAND2_X1 U7582 ( .A1(n5986), .A2(n5985), .ZN(n7897) );
  OR2_X1 U7583 ( .A1(n5766), .A2(n7897), .ZN(n5987) );
  NOR2_X1 U7584 ( .A1(n8576), .A2(n8504), .ZN(n7894) );
  NAND2_X1 U7585 ( .A1(n6621), .A2(n8299), .ZN(n5994) );
  NAND2_X1 U7586 ( .A1(n5991), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5992) );
  XNOR2_X1 U7587 ( .A(n5992), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8701) );
  AOI22_X1 U7588 ( .A1(n6036), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6590), .B2(
        n8701), .ZN(n5993) );
  XNOR2_X1 U7589 ( .A(n7901), .B(n6177), .ZN(n5996) );
  AOI22_X1 U7590 ( .A1(n8572), .A2(n5997), .B1(n7894), .B2(n5996), .ZN(n5995)
         );
  NAND2_X1 U7591 ( .A1(n7893), .A2(n5995), .ZN(n6003) );
  INV_X1 U7592 ( .A(n8572), .ZN(n6001) );
  OAI21_X1 U7593 ( .B1(n5996), .B2(n7894), .A(n5997), .ZN(n6000) );
  INV_X1 U7594 ( .A(n5996), .ZN(n8570) );
  INV_X1 U7595 ( .A(n7894), .ZN(n5998) );
  INV_X1 U7596 ( .A(n5997), .ZN(n8571) );
  AND3_X1 U7597 ( .A1(n8570), .A2(n5998), .A3(n8571), .ZN(n5999) );
  AOI21_X1 U7598 ( .B1(n6001), .B2(n6000), .A(n5999), .ZN(n6002) );
  NAND2_X1 U7599 ( .A1(n6663), .A2(n8299), .ZN(n6006) );
  NAND2_X1 U7600 ( .A1(n4453), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6004) );
  XNOR2_X1 U7601 ( .A(n6004), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8729) );
  AOI22_X1 U7602 ( .A1(n6036), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6590), .B2(
        n8729), .ZN(n6005) );
  XNOR2_X1 U7603 ( .A(n9079), .B(n6177), .ZN(n6013) );
  NAND2_X1 U7604 ( .A1(n6594), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6012) );
  INV_X1 U7605 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8736) );
  OR2_X1 U7606 ( .A1(n5753), .A2(n8736), .ZN(n6011) );
  NAND2_X1 U7607 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(n6007), .ZN(n6024) );
  OAI21_X1 U7608 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(n6007), .A(n6024), .ZN(
        n7817) );
  OR2_X1 U7609 ( .A1(n5766), .A2(n7817), .ZN(n6010) );
  INV_X1 U7610 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n6008) );
  OR2_X1 U7611 ( .A1(n6609), .A2(n6008), .ZN(n6009) );
  NOR2_X1 U7612 ( .A1(n8649), .A2(n8504), .ZN(n6014) );
  NAND2_X1 U7613 ( .A1(n6013), .A2(n6014), .ZN(n6019) );
  INV_X1 U7614 ( .A(n6013), .ZN(n6016) );
  INV_X1 U7615 ( .A(n6014), .ZN(n6015) );
  NAND2_X1 U7616 ( .A1(n6016), .A2(n6015), .ZN(n6017) );
  NAND2_X1 U7617 ( .A1(n6019), .A2(n6017), .ZN(n6506) );
  NAND2_X1 U7618 ( .A1(n6823), .A2(n8299), .ZN(n6022) );
  XNOR2_X1 U7619 ( .A(n6020), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8745) );
  AOI22_X1 U7620 ( .A1(n6036), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6590), .B2(
        n8745), .ZN(n6021) );
  XNOR2_X1 U7621 ( .A(n9072), .B(n6155), .ZN(n6031) );
  NAND2_X1 U7622 ( .A1(n6234), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6030) );
  INV_X1 U7623 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6023) );
  OR2_X1 U7624 ( .A1(n5767), .A2(n6023), .ZN(n6029) );
  OAI21_X1 U7625 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(n6025), .A(n6040), .ZN(
        n8984) );
  OR2_X1 U7626 ( .A1(n5766), .A2(n8984), .ZN(n6028) );
  INV_X1 U7627 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n6026) );
  OR2_X1 U7628 ( .A1(n6609), .A2(n6026), .ZN(n6027) );
  NOR2_X1 U7629 ( .A1(n8779), .A2(n8504), .ZN(n6032) );
  XNOR2_X1 U7630 ( .A(n6031), .B(n6032), .ZN(n7914) );
  NAND2_X1 U7631 ( .A1(n7915), .A2(n7914), .ZN(n7913) );
  INV_X1 U7632 ( .A(n6031), .ZN(n6033) );
  NAND2_X1 U7633 ( .A1(n6033), .A2(n6032), .ZN(n6034) );
  NAND2_X1 U7634 ( .A1(n7913), .A2(n6034), .ZN(n8528) );
  NAND2_X1 U7635 ( .A1(n6917), .A2(n8299), .ZN(n6038) );
  AOI22_X1 U7636 ( .A1(n6036), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6590), .B2(
        n8342), .ZN(n6037) );
  XNOR2_X1 U7637 ( .A(n9068), .B(n6155), .ZN(n6046) );
  NAND2_X1 U7638 ( .A1(n5783), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6045) );
  INV_X1 U7639 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8753) );
  OR2_X1 U7640 ( .A1(n5753), .A2(n8753), .ZN(n6044) );
  INV_X1 U7641 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6039) );
  OR2_X1 U7642 ( .A1(n6606), .A2(n6039), .ZN(n6043) );
  OAI21_X1 U7643 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(n6041), .A(n6053), .ZN(
        n8963) );
  OR2_X1 U7644 ( .A1(n5766), .A2(n8963), .ZN(n6042) );
  OR2_X1 U7645 ( .A1(n8953), .A2(n8504), .ZN(n6047) );
  NAND2_X1 U7646 ( .A1(n6046), .A2(n6047), .ZN(n8527) );
  NAND2_X1 U7647 ( .A1(n8528), .A2(n8527), .ZN(n6050) );
  INV_X1 U7648 ( .A(n6046), .ZN(n6049) );
  INV_X1 U7649 ( .A(n6047), .ZN(n6048) );
  NAND2_X1 U7650 ( .A1(n6049), .A2(n6048), .ZN(n8526) );
  NAND2_X1 U7651 ( .A1(n6050), .A2(n8526), .ZN(n8603) );
  NAND2_X1 U7652 ( .A1(n6970), .A2(n8299), .ZN(n6052) );
  OR2_X1 U7653 ( .A1(n8300), .A2(n8278), .ZN(n6051) );
  XNOR2_X1 U7654 ( .A(n9062), .B(n6155), .ZN(n6060) );
  NAND2_X1 U7655 ( .A1(n6234), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6059) );
  INV_X1 U7656 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n10036) );
  OR2_X1 U7657 ( .A1(n6609), .A2(n10036), .ZN(n6058) );
  OAI21_X1 U7658 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(n6054), .A(n6068), .ZN(
        n8942) );
  OR2_X1 U7659 ( .A1(n5766), .A2(n8942), .ZN(n6057) );
  INV_X1 U7660 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n6055) );
  OR2_X1 U7661 ( .A1(n6606), .A2(n6055), .ZN(n6056) );
  NOR2_X1 U7662 ( .A1(n8648), .A2(n8504), .ZN(n6061) );
  XNOR2_X1 U7663 ( .A(n6060), .B(n6061), .ZN(n8604) );
  INV_X1 U7664 ( .A(n6060), .ZN(n6062) );
  NAND2_X1 U7665 ( .A1(n6062), .A2(n6061), .ZN(n6063) );
  NAND2_X1 U7666 ( .A1(n6981), .A2(n8299), .ZN(n6065) );
  OR2_X1 U7667 ( .A1(n8300), .A2(n6982), .ZN(n6064) );
  XNOR2_X1 U7668 ( .A(n9057), .B(n6155), .ZN(n6074) );
  NAND2_X1 U7669 ( .A1(n6234), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6073) );
  INV_X1 U7670 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8927) );
  OR2_X1 U7671 ( .A1(n5767), .A2(n8927), .ZN(n6072) );
  INV_X1 U7672 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7673 ( .A1(n6068), .A2(n6067), .ZN(n6069) );
  NAND2_X1 U7674 ( .A1(n6082), .A2(n6069), .ZN(n8935) );
  OR2_X1 U7675 ( .A1(n5766), .A2(n8935), .ZN(n6071) );
  INV_X1 U7676 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n10153) );
  OR2_X1 U7677 ( .A1(n6609), .A2(n10153), .ZN(n6070) );
  NOR2_X1 U7678 ( .A1(n8951), .A2(n8504), .ZN(n6075) );
  XNOR2_X1 U7679 ( .A(n6074), .B(n6075), .ZN(n8555) );
  INV_X1 U7680 ( .A(n6074), .ZN(n6076) );
  NAND2_X1 U7681 ( .A1(n7245), .A2(n8299), .ZN(n6078) );
  OR2_X1 U7682 ( .A1(n8300), .A2(n7246), .ZN(n6077) );
  XNOR2_X1 U7683 ( .A(n9052), .B(n6155), .ZN(n6089) );
  NAND2_X1 U7684 ( .A1(n6234), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6088) );
  INV_X1 U7685 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n6079) );
  OR2_X1 U7686 ( .A1(n6606), .A2(n6079), .ZN(n6087) );
  INV_X1 U7687 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7688 ( .A1(n6082), .A2(n6081), .ZN(n6083) );
  NAND2_X1 U7689 ( .A1(n6114), .A2(n6083), .ZN(n8913) );
  OR2_X1 U7690 ( .A1(n5766), .A2(n8913), .ZN(n6086) );
  INV_X1 U7691 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n6084) );
  OR2_X1 U7692 ( .A1(n6609), .A2(n6084), .ZN(n6085) );
  OR2_X1 U7693 ( .A1(n8786), .A2(n8504), .ZN(n8610) );
  NAND2_X1 U7694 ( .A1(n8611), .A2(n8610), .ZN(n8609) );
  INV_X1 U7695 ( .A(n6089), .ZN(n6090) );
  NAND2_X1 U7696 ( .A1(n8609), .A2(n6092), .ZN(n6113) );
  INV_X1 U7697 ( .A(n6113), .ZN(n6095) );
  NAND2_X1 U7698 ( .A1(n7298), .A2(n8299), .ZN(n6094) );
  OR2_X1 U7699 ( .A1(n8300), .A2(n7297), .ZN(n6093) );
  XNOR2_X1 U7700 ( .A(n9045), .B(n6177), .ZN(n6112) );
  NAND2_X1 U7701 ( .A1(n6095), .A2(n6112), .ZN(n8591) );
  NAND2_X1 U7702 ( .A1(n7469), .A2(n8299), .ZN(n6097) );
  OR2_X1 U7703 ( .A1(n8300), .A2(n7472), .ZN(n6096) );
  XNOR2_X1 U7704 ( .A(n8880), .B(n6177), .ZN(n8595) );
  NAND2_X1 U7705 ( .A1(n6234), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6106) );
  INV_X1 U7706 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6098) );
  OR2_X1 U7707 ( .A1(n6606), .A2(n6098), .ZN(n6105) );
  INV_X1 U7708 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U7709 ( .A1(n6116), .A2(n8598), .ZN(n6101) );
  NAND2_X1 U7710 ( .A1(n6128), .A2(n6101), .ZN(n8877) );
  OR2_X1 U7711 ( .A1(n5766), .A2(n8877), .ZN(n6104) );
  INV_X1 U7712 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n6102) );
  OR2_X1 U7713 ( .A1(n6609), .A2(n6102), .ZN(n6103) );
  NAND4_X1 U7714 ( .A1(n6106), .A2(n6105), .A3(n6104), .A4(n6103), .ZN(n8893)
         );
  NAND2_X1 U7715 ( .A1(n8893), .A2(n5792), .ZN(n6107) );
  AND2_X1 U7716 ( .A1(n8595), .A2(n6107), .ZN(n6110) );
  INV_X1 U7717 ( .A(n8595), .ZN(n6108) );
  INV_X1 U7718 ( .A(n6107), .ZN(n8594) );
  NAND2_X1 U7719 ( .A1(n6108), .A2(n8594), .ZN(n6109) );
  INV_X1 U7720 ( .A(n6111), .ZN(n6123) );
  XNOR2_X1 U7721 ( .A(n6113), .B(n6112), .ZN(n8519) );
  INV_X1 U7722 ( .A(n8893), .ZN(n8521) );
  NAND2_X1 U7723 ( .A1(n6234), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6120) );
  INV_X1 U7724 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8900) );
  OR2_X1 U7725 ( .A1(n5767), .A2(n8900), .ZN(n6119) );
  INV_X1 U7726 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8520) );
  NAND2_X1 U7727 ( .A1(n6114), .A2(n8520), .ZN(n6115) );
  NAND2_X1 U7728 ( .A1(n6116), .A2(n6115), .ZN(n8899) );
  OR2_X1 U7729 ( .A1(n5766), .A2(n8899), .ZN(n6118) );
  INV_X1 U7730 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n10095) );
  OR2_X1 U7731 ( .A1(n6609), .A2(n10095), .ZN(n6117) );
  NAND4_X1 U7732 ( .A1(n6120), .A2(n6119), .A3(n6118), .A4(n6117), .ZN(n8647)
         );
  NAND2_X1 U7733 ( .A1(n8647), .A2(n5792), .ZN(n8592) );
  AOI21_X1 U7734 ( .B1(n8595), .B2(n8521), .A(n8592), .ZN(n6121) );
  NAND2_X1 U7735 ( .A1(n8519), .A2(n6121), .ZN(n6122) );
  NAND2_X1 U7736 ( .A1(n7588), .A2(n8299), .ZN(n6125) );
  OR2_X1 U7737 ( .A1(n8300), .A2(n7590), .ZN(n6124) );
  XNOR2_X1 U7738 ( .A(n9037), .B(n6155), .ZN(n6135) );
  NAND2_X1 U7739 ( .A1(n6234), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6134) );
  INV_X1 U7740 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8866) );
  OR2_X1 U7741 ( .A1(n5767), .A2(n8866), .ZN(n6133) );
  INV_X1 U7742 ( .A(n6128), .ZN(n6126) );
  NAND2_X1 U7743 ( .A1(n6126), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6142) );
  INV_X1 U7744 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7745 ( .A1(n6128), .A2(n6127), .ZN(n6129) );
  NAND2_X1 U7746 ( .A1(n6142), .A2(n6129), .ZN(n8865) );
  OR2_X1 U7747 ( .A1(n5766), .A2(n8865), .ZN(n6132) );
  INV_X1 U7748 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n6130) );
  OR2_X1 U7749 ( .A1(n6609), .A2(n6130), .ZN(n6131) );
  NOR2_X1 U7750 ( .A1(n8883), .A2(n8504), .ZN(n6136) );
  XNOR2_X1 U7751 ( .A(n6135), .B(n6136), .ZN(n8561) );
  INV_X1 U7752 ( .A(n6135), .ZN(n6137) );
  NAND2_X1 U7753 ( .A1(n6137), .A2(n6136), .ZN(n6138) );
  OR2_X1 U7754 ( .A1(n8300), .A2(n10190), .ZN(n6139) );
  XNOR2_X1 U7755 ( .A(n9031), .B(n6155), .ZN(n6148) );
  NAND2_X1 U7756 ( .A1(n6234), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6147) );
  INV_X1 U7757 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n10221) );
  OR2_X1 U7758 ( .A1(n5767), .A2(n10221), .ZN(n6146) );
  INV_X1 U7759 ( .A(n6142), .ZN(n6141) );
  NAND2_X1 U7760 ( .A1(n6141), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6168) );
  INV_X1 U7761 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10160) );
  NAND2_X1 U7762 ( .A1(n6142), .A2(n10160), .ZN(n6143) );
  NAND2_X1 U7763 ( .A1(n6168), .A2(n6143), .ZN(n8857) );
  OR2_X1 U7764 ( .A1(n5766), .A2(n8857), .ZN(n6145) );
  INV_X1 U7765 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n10033) );
  OR2_X1 U7766 ( .A1(n6609), .A2(n10033), .ZN(n6144) );
  NOR2_X1 U7767 ( .A1(n8837), .A2(n8504), .ZN(n6149) );
  XNOR2_X1 U7768 ( .A(n6148), .B(n6149), .ZN(n8635) );
  INV_X1 U7769 ( .A(n6148), .ZN(n6150) );
  NAND2_X1 U7770 ( .A1(n6150), .A2(n6149), .ZN(n6151) );
  NAND2_X1 U7771 ( .A1(n6152), .A2(n6151), .ZN(n8512) );
  NAND2_X1 U7772 ( .A1(n7709), .A2(n8299), .ZN(n6154) );
  OR2_X1 U7773 ( .A1(n8300), .A2(n7931), .ZN(n6153) );
  XNOR2_X1 U7774 ( .A(n8830), .B(n6155), .ZN(n6164) );
  NAND2_X1 U7775 ( .A1(n6234), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6161) );
  INV_X1 U7776 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6156) );
  OR2_X1 U7777 ( .A1(n6606), .A2(n6156), .ZN(n6160) );
  INV_X1 U7778 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8514) );
  XNOR2_X1 U7779 ( .A(n6168), .B(n8514), .ZN(n8827) );
  OR2_X1 U7780 ( .A1(n5766), .A2(n8827), .ZN(n6159) );
  INV_X1 U7781 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6157) );
  OR2_X1 U7782 ( .A1(n6609), .A2(n6157), .ZN(n6158) );
  NAND4_X1 U7783 ( .A1(n6161), .A2(n6160), .A3(n6159), .A4(n6158), .ZN(n8646)
         );
  NAND2_X1 U7784 ( .A1(n8646), .A2(n5792), .ZN(n6162) );
  XNOR2_X1 U7785 ( .A(n6164), .B(n6162), .ZN(n8513) );
  INV_X1 U7786 ( .A(n6162), .ZN(n6163) );
  AND2_X1 U7787 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  NAND2_X1 U7788 ( .A1(n6594), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6176) );
  INV_X1 U7789 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6166) );
  OR2_X1 U7790 ( .A1(n5753), .A2(n6166), .ZN(n6175) );
  INV_X1 U7791 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6167) );
  OAI21_X1 U7792 ( .B1(n6168), .B2(n8514), .A(n6167), .ZN(n6171) );
  INV_X1 U7793 ( .A(n6168), .ZN(n6170) );
  AND2_X1 U7794 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6169) );
  NAND2_X1 U7795 ( .A1(n6170), .A2(n6169), .ZN(n8799) );
  NAND2_X1 U7796 ( .A1(n6171), .A2(n8799), .ZN(n6243) );
  OR2_X1 U7797 ( .A1(n5766), .A2(n6243), .ZN(n6174) );
  INV_X1 U7798 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6172) );
  OR2_X1 U7799 ( .A1(n6609), .A2(n6172), .ZN(n6173) );
  NAND4_X1 U7800 ( .A1(n6176), .A2(n6175), .A3(n6174), .A4(n6173), .ZN(n8795)
         );
  NAND2_X1 U7801 ( .A1(n8795), .A2(n5792), .ZN(n6178) );
  XNOR2_X1 U7802 ( .A(n6178), .B(n6177), .ZN(n6221) );
  INV_X1 U7803 ( .A(n6221), .ZN(n6222) );
  NAND2_X1 U7804 ( .A1(n7789), .A2(n8299), .ZN(n6180) );
  OR2_X1 U7805 ( .A1(n8300), .A2(n10188), .ZN(n6179) );
  INV_X1 U7806 ( .A(n6191), .ZN(n6187) );
  NAND2_X1 U7807 ( .A1(n6182), .A2(n6187), .ZN(n6189) );
  NAND2_X1 U7808 ( .A1(n6189), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6183) );
  MUX2_X1 U7809 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6183), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6185) );
  NAND2_X1 U7810 ( .A1(n6185), .A2(n6184), .ZN(n7646) );
  INV_X1 U7811 ( .A(n7646), .ZN(n6197) );
  NAND2_X1 U7812 ( .A1(n4452), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6188) );
  MUX2_X1 U7813 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6188), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6190) );
  NAND2_X1 U7814 ( .A1(n6190), .A2(n6189), .ZN(n7589) );
  NAND2_X1 U7815 ( .A1(n6191), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6210) );
  INV_X1 U7816 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U7817 ( .A1(n6210), .A2(n6192), .ZN(n6212) );
  NAND2_X1 U7818 ( .A1(n6212), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6194) );
  INV_X1 U7819 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6193) );
  XNOR2_X1 U7820 ( .A(n6194), .B(n6193), .ZN(n7474) );
  XNOR2_X1 U7821 ( .A(n7474), .B(P2_B_REG_SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7822 ( .A1(n7589), .A2(n6195), .ZN(n6196) );
  INV_X1 U7823 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9869) );
  AND2_X1 U7824 ( .A1(n7646), .A2(n7589), .ZN(n9871) );
  AOI21_X1 U7825 ( .B1(n9864), .B2(n9869), .A(n9871), .ZN(n7049) );
  NOR4_X1 U7826 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6201) );
  NOR4_X1 U7827 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6200) );
  NOR4_X1 U7828 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6199) );
  NOR4_X1 U7829 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6198) );
  NAND4_X1 U7830 ( .A1(n6201), .A2(n6200), .A3(n6199), .A4(n6198), .ZN(n6207)
         );
  NOR2_X1 U7831 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .ZN(
        n6205) );
  NOR4_X1 U7832 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6204) );
  NOR4_X1 U7833 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6203) );
  NOR4_X1 U7834 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n6202) );
  NAND4_X1 U7835 ( .A1(n6205), .A2(n6204), .A3(n6203), .A4(n6202), .ZN(n6206)
         );
  OAI21_X1 U7836 ( .B1(n6207), .B2(n6206), .A(n9864), .ZN(n6827) );
  NAND2_X1 U7837 ( .A1(n7049), .A2(n6827), .ZN(n6240) );
  INV_X1 U7838 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10008) );
  AND2_X1 U7839 ( .A1(n7646), .A2(n7474), .ZN(n9867) );
  AOI21_X1 U7840 ( .B1(n9864), .B2(n10008), .A(n9867), .ZN(n6860) );
  NOR2_X1 U7841 ( .A1(n7646), .A2(n7589), .ZN(n6209) );
  INV_X1 U7842 ( .A(n7474), .ZN(n6208) );
  NAND2_X1 U7843 ( .A1(n6209), .A2(n6208), .ZN(n6503) );
  INV_X1 U7844 ( .A(n6210), .ZN(n6211) );
  NAND2_X1 U7845 ( .A1(n6211), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n6213) );
  AND2_X1 U7846 ( .A1(n6213), .A2(n6212), .ZN(n6588) );
  NOR2_X1 U7847 ( .A1(n6588), .A2(P2_U3152), .ZN(n9870) );
  NAND2_X1 U7848 ( .A1(n6503), .A2(n9870), .ZN(n9865) );
  NAND2_X1 U7849 ( .A1(n6860), .A2(n8497), .ZN(n6214) );
  NOR2_X1 U7850 ( .A1(n6240), .A2(n6214), .ZN(n6232) );
  INV_X1 U7851 ( .A(n6216), .ZN(n6852) );
  NOR2_X1 U7852 ( .A1(n6216), .A2(n9873), .ZN(n7059) );
  NAND2_X1 U7853 ( .A1(n6232), .A2(n7059), .ZN(n6219) );
  AND2_X1 U7854 ( .A1(n8342), .A2(n8340), .ZN(n6217) );
  NAND2_X1 U7855 ( .A1(n9922), .A2(n8338), .ZN(n6830) );
  INV_X1 U7856 ( .A(n6830), .ZN(n6218) );
  NOR3_X1 U7857 ( .A1(n8812), .A2(n6222), .A3(n8629), .ZN(n6220) );
  AOI21_X1 U7858 ( .B1(n6222), .B2(n8812), .A(n6220), .ZN(n6230) );
  NOR3_X1 U7859 ( .A1(n8812), .A2(n6221), .A3(n8629), .ZN(n6224) );
  NOR2_X1 U7860 ( .A1(n9020), .A2(n6222), .ZN(n6223) );
  NAND2_X1 U7861 ( .A1(n6231), .A2(n6225), .ZN(n6229) );
  INV_X1 U7862 ( .A(n8629), .ZN(n8619) );
  OR2_X1 U7863 ( .A1(n6226), .A2(n9873), .ZN(n9925) );
  AND2_X1 U7864 ( .A1(n8501), .A2(n8351), .ZN(n6843) );
  INV_X1 U7865 ( .A(n6843), .ZN(n6591) );
  AND2_X1 U7866 ( .A1(n9925), .A2(n6591), .ZN(n6227) );
  NAND2_X1 U7867 ( .A1(n6232), .A2(n6227), .ZN(n8643) );
  OAI21_X1 U7868 ( .B1(n8812), .B2(n8619), .A(n8643), .ZN(n6228) );
  OAI211_X1 U7869 ( .C1(n6231), .C2(n6230), .A(n6229), .B(n6228), .ZN(n6247)
         );
  AND2_X1 U7870 ( .A1(n6232), .A2(n6226), .ZN(n8638) );
  INV_X1 U7871 ( .A(n6233), .ZN(n6716) );
  AND2_X1 U7872 ( .A1(n6716), .A2(n6843), .ZN(n8995) );
  AND2_X1 U7873 ( .A1(n8638), .A2(n8995), .ZN(n8628) );
  AOI22_X1 U7874 ( .A1(n8628), .A2(n8646), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6245) );
  AND2_X1 U7875 ( .A1(n6233), .A2(n6843), .ZN(n8993) );
  AND2_X1 U7876 ( .A1(n8638), .A2(n8993), .ZN(n8624) );
  NAND2_X1 U7877 ( .A1(n6234), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6239) );
  OR2_X1 U7878 ( .A1(n5767), .A2(n10174), .ZN(n6238) );
  OR2_X1 U7879 ( .A1(n5766), .A2(n8799), .ZN(n6237) );
  INV_X1 U7880 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6235) );
  OR2_X1 U7881 ( .A1(n6609), .A2(n6235), .ZN(n6236) );
  INV_X1 U7882 ( .A(n8816), .ZN(n8645) );
  INV_X1 U7883 ( .A(n6860), .ZN(n7050) );
  OAI21_X1 U7884 ( .B1(n6240), .B2(n7050), .A(n6830), .ZN(n6925) );
  INV_X1 U7885 ( .A(n6588), .ZN(n6241) );
  OR2_X1 U7886 ( .A1(n6226), .A2(n6591), .ZN(n6826) );
  NAND4_X1 U7887 ( .A1(n6925), .A2(n6503), .A3(n6241), .A4(n6826), .ZN(n6242)
         );
  INV_X1 U7888 ( .A(n6243), .ZN(n8810) );
  AOI22_X1 U7889 ( .A1(n8624), .A2(n8645), .B1(n8627), .B2(n8810), .ZN(n6244)
         );
  NAND2_X1 U7890 ( .A1(n6247), .A2(n6246), .ZN(P2_U3222) );
  AND2_X2 U7891 ( .A1(n6890), .A2(n6478), .ZN(n6267) );
  NAND2_X1 U7892 ( .A1(n8205), .A2(n6248), .ZN(n7128) );
  AOI22_X1 U7893 ( .A1(n9460), .A2(n6457), .B1(n6447), .B2(n9218), .ZN(n9146)
         );
  OAI22_X1 U7894 ( .A1(n8270), .A2(n6445), .B1(n9151), .B2(n6444), .ZN(n6250)
         );
  XOR2_X1 U7895 ( .A(n6452), .B(n6250), .Z(n9192) );
  NAND2_X1 U7896 ( .A1(n9235), .A2(n6267), .ZN(n6252) );
  NAND2_X1 U7897 ( .A1(n7130), .A2(n6456), .ZN(n6251) );
  INV_X1 U7898 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10045) );
  INV_X1 U7899 ( .A(n6687), .ZN(n6253) );
  NAND2_X1 U7900 ( .A1(n6253), .A2(n6452), .ZN(n6257) );
  NAND2_X1 U7901 ( .A1(n7130), .A2(n6267), .ZN(n6255) );
  INV_X1 U7902 ( .A(n6478), .ZN(n6497) );
  NAND2_X1 U7903 ( .A1(n6497), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U7904 ( .A1(n6257), .A2(n6690), .ZN(n6265) );
  NAND2_X1 U7905 ( .A1(n6258), .A2(n6267), .ZN(n6261) );
  INV_X1 U7906 ( .A(n7333), .ZN(n6259) );
  NAND2_X1 U7907 ( .A1(n6261), .A2(n6260), .ZN(n6262) );
  XNOR2_X1 U7908 ( .A(n6262), .B(n6452), .ZN(n6263) );
  XNOR2_X1 U7909 ( .A(n6265), .B(n6263), .ZN(n7003) );
  AOI22_X1 U7910 ( .A1(n6258), .A2(n6447), .B1(n6259), .B2(n6457), .ZN(n7005)
         );
  NAND2_X1 U7911 ( .A1(n7003), .A2(n7005), .ZN(n7004) );
  INV_X1 U7912 ( .A(n6263), .ZN(n6264) );
  NAND2_X1 U7913 ( .A1(n6265), .A2(n6264), .ZN(n6266) );
  NAND2_X1 U7914 ( .A1(n7004), .A2(n6266), .ZN(n7079) );
  INV_X1 U7915 ( .A(n6267), .ZN(n6444) );
  OAI22_X1 U7916 ( .A1(n6268), .A2(n6444), .B1(n9796), .B2(n6445), .ZN(n6269)
         );
  XNOR2_X1 U7917 ( .A(n6269), .B(n6460), .ZN(n6270) );
  OAI22_X1 U7918 ( .A1(n6268), .A2(n6462), .B1(n9796), .B2(n6444), .ZN(n6271)
         );
  XNOR2_X1 U7919 ( .A(n6270), .B(n6271), .ZN(n7078) );
  NAND2_X1 U7920 ( .A1(n7079), .A2(n7078), .ZN(n6274) );
  INV_X1 U7921 ( .A(n6270), .ZN(n6272) );
  OR2_X1 U7922 ( .A1(n6272), .A2(n6271), .ZN(n6273) );
  OAI22_X1 U7923 ( .A1(n7201), .A2(n6444), .B1(n9801), .B2(n6445), .ZN(n6275)
         );
  XNOR2_X1 U7924 ( .A(n6275), .B(n6460), .ZN(n6278) );
  OAI22_X1 U7925 ( .A1(n7201), .A2(n6462), .B1(n9801), .B2(n6444), .ZN(n6276)
         );
  XNOR2_X1 U7926 ( .A(n6278), .B(n6276), .ZN(n6973) );
  INV_X1 U7927 ( .A(n6276), .ZN(n6277) );
  NAND2_X1 U7928 ( .A1(n6278), .A2(n6277), .ZN(n6961) );
  OAI22_X1 U7929 ( .A1(n7258), .A2(n6444), .B1(n7187), .B2(n6445), .ZN(n6279)
         );
  OAI22_X1 U7930 ( .A1(n7258), .A2(n6462), .B1(n7187), .B2(n6444), .ZN(n6288)
         );
  INV_X1 U7931 ( .A(n6288), .ZN(n6280) );
  NAND2_X1 U7932 ( .A1(n6289), .A2(n6280), .ZN(n6287) );
  AND2_X1 U7933 ( .A1(n6961), .A2(n6287), .ZN(n7252) );
  OAI22_X1 U7934 ( .A1(n7022), .A2(n6462), .B1(n9812), .B2(n6444), .ZN(n6293)
         );
  NAND2_X1 U7935 ( .A1(n9231), .A2(n6447), .ZN(n6283) );
  NAND2_X1 U7936 ( .A1(n9773), .A2(n6457), .ZN(n6282) );
  NAND2_X1 U7937 ( .A1(n6283), .A2(n6282), .ZN(n7255) );
  NAND2_X1 U7938 ( .A1(n9231), .A2(n6457), .ZN(n6285) );
  NAND2_X1 U7939 ( .A1(n9773), .A2(n6456), .ZN(n6284) );
  NAND2_X1 U7940 ( .A1(n6285), .A2(n6284), .ZN(n6286) );
  OAI22_X1 U7941 ( .A1(n7420), .A2(n6293), .B1(n7255), .B2(n7415), .ZN(n6291)
         );
  INV_X1 U7942 ( .A(n6287), .ZN(n6290) );
  XNOR2_X1 U7943 ( .A(n6289), .B(n6288), .ZN(n6959) );
  NAND2_X1 U7944 ( .A1(n7415), .A2(n7255), .ZN(n6292) );
  INV_X1 U7945 ( .A(n6293), .ZN(n7419) );
  NAND2_X1 U7946 ( .A1(n6292), .A2(n7419), .ZN(n6295) );
  INV_X1 U7947 ( .A(n6292), .ZN(n6294) );
  AOI22_X1 U7948 ( .A1(n7420), .A2(n6295), .B1(n6294), .B2(n6293), .ZN(n7032)
         );
  OAI22_X1 U7949 ( .A1(n7427), .A2(n6444), .B1(n9819), .B2(n6445), .ZN(n6296)
         );
  XNOR2_X1 U7950 ( .A(n6296), .B(n6460), .ZN(n6300) );
  INV_X1 U7951 ( .A(n6300), .ZN(n6297) );
  OAI22_X1 U7952 ( .A1(n7427), .A2(n6462), .B1(n9819), .B2(n6444), .ZN(n6298)
         );
  NAND2_X1 U7953 ( .A1(n6297), .A2(n6298), .ZN(n7034) );
  INV_X1 U7954 ( .A(n6298), .ZN(n6299) );
  NAND2_X1 U7955 ( .A1(n6300), .A2(n6299), .ZN(n7033) );
  NAND2_X1 U7956 ( .A1(n7410), .A2(n6457), .ZN(n6302) );
  OAI21_X1 U7957 ( .B1(n6309), .B2(n6462), .A(n6302), .ZN(n6307) );
  NAND2_X1 U7958 ( .A1(n6303), .A2(n6307), .ZN(n7163) );
  INV_X1 U7959 ( .A(n6307), .ZN(n6304) );
  OR2_X1 U7960 ( .A1(n6307), .A2(n7033), .ZN(n7160) );
  NAND2_X1 U7961 ( .A1(n7410), .A2(n6456), .ZN(n6308) );
  OAI21_X1 U7962 ( .B1(n6309), .B2(n6444), .A(n6308), .ZN(n6310) );
  XNOR2_X1 U7963 ( .A(n6310), .B(n6452), .ZN(n7165) );
  AND2_X1 U7964 ( .A1(n7160), .A2(n7165), .ZN(n6311) );
  NAND2_X1 U7965 ( .A1(n7161), .A2(n6311), .ZN(n7162) );
  NAND2_X1 U7966 ( .A1(n9830), .A2(n6456), .ZN(n6313) );
  NAND2_X1 U7967 ( .A1(n9227), .A2(n6457), .ZN(n6312) );
  NAND2_X1 U7968 ( .A1(n6313), .A2(n6312), .ZN(n6314) );
  XNOR2_X1 U7969 ( .A(n6314), .B(n6460), .ZN(n6316) );
  AOI22_X1 U7970 ( .A1(n9830), .A2(n6457), .B1(n6447), .B2(n9227), .ZN(n6315)
         );
  XNOR2_X1 U7971 ( .A(n6316), .B(n6315), .ZN(n7934) );
  NAND2_X1 U7972 ( .A1(n6316), .A2(n6315), .ZN(n6353) );
  NAND2_X1 U7973 ( .A1(n7574), .A2(n6456), .ZN(n6318) );
  NAND2_X1 U7974 ( .A1(n9226), .A2(n6457), .ZN(n6317) );
  NAND2_X1 U7975 ( .A1(n6318), .A2(n6317), .ZN(n6319) );
  XNOR2_X1 U7976 ( .A(n6319), .B(n6460), .ZN(n7303) );
  NOR2_X1 U7977 ( .A1(n7935), .A2(n6462), .ZN(n6320) );
  AOI21_X1 U7978 ( .B1(n7574), .B2(n6457), .A(n6320), .ZN(n7302) );
  AND2_X1 U7979 ( .A1(n7303), .A2(n7302), .ZN(n6352) );
  NAND2_X1 U7980 ( .A1(n7516), .A2(n6456), .ZN(n6322) );
  NAND2_X1 U7981 ( .A1(n9225), .A2(n6457), .ZN(n6321) );
  NAND2_X1 U7982 ( .A1(n6322), .A2(n6321), .ZN(n6323) );
  XNOR2_X1 U7983 ( .A(n6323), .B(n6452), .ZN(n6335) );
  AND2_X1 U7984 ( .A1(n9225), .A2(n6447), .ZN(n6324) );
  AOI21_X1 U7985 ( .B1(n7516), .B2(n6457), .A(n6324), .ZN(n6334) );
  INV_X1 U7986 ( .A(n6334), .ZN(n6325) );
  NAND2_X1 U7987 ( .A1(n6335), .A2(n6325), .ZN(n7524) );
  NAND2_X1 U7988 ( .A1(n9224), .A2(n6457), .ZN(n6326) );
  XNOR2_X1 U7989 ( .A(n6327), .B(n6460), .ZN(n6333) );
  INV_X1 U7990 ( .A(n6333), .ZN(n6331) );
  NOR2_X1 U7991 ( .A1(n7551), .A2(n6462), .ZN(n6329) );
  AOI21_X1 U7992 ( .B1(n9593), .B2(n6457), .A(n6329), .ZN(n6332) );
  INV_X1 U7993 ( .A(n6332), .ZN(n6330) );
  NAND2_X1 U7994 ( .A1(n6333), .A2(n6332), .ZN(n7520) );
  XNOR2_X1 U7995 ( .A(n6335), .B(n6334), .ZN(n7522) );
  AND2_X1 U7996 ( .A1(n7522), .A2(n7520), .ZN(n6336) );
  NOR2_X1 U7997 ( .A1(n6337), .A2(n6336), .ZN(n6342) );
  INV_X1 U7998 ( .A(n7303), .ZN(n6339) );
  INV_X1 U7999 ( .A(n7302), .ZN(n6338) );
  NAND2_X1 U8000 ( .A1(n6339), .A2(n6338), .ZN(n6356) );
  AND2_X1 U8001 ( .A1(n6356), .A2(n6340), .ZN(n6341) );
  OR2_X1 U8002 ( .A1(n6342), .A2(n6341), .ZN(n6343) );
  NAND2_X1 U8003 ( .A1(n9501), .A2(n6456), .ZN(n6346) );
  NAND2_X1 U8004 ( .A1(n9223), .A2(n6457), .ZN(n6345) );
  NAND2_X1 U8005 ( .A1(n6346), .A2(n6345), .ZN(n6347) );
  XNOR2_X1 U8006 ( .A(n6347), .B(n6452), .ZN(n7547) );
  NAND2_X1 U8007 ( .A1(n9501), .A2(n6457), .ZN(n6349) );
  NAND2_X1 U8008 ( .A1(n9223), .A2(n6447), .ZN(n6348) );
  NAND2_X1 U8009 ( .A1(n6349), .A2(n6348), .ZN(n7548) );
  OAI21_X1 U8010 ( .B1(n7550), .B2(n7547), .A(n7548), .ZN(n6362) );
  AND2_X1 U8011 ( .A1(n7520), .A2(n7547), .ZN(n6358) );
  INV_X1 U8012 ( .A(n6358), .ZN(n6351) );
  OR2_X1 U8013 ( .A1(n6351), .A2(n6350), .ZN(n6361) );
  INV_X1 U8014 ( .A(n6352), .ZN(n6354) );
  AND2_X1 U8015 ( .A1(n6354), .A2(n6353), .ZN(n6355) );
  NAND2_X1 U8016 ( .A1(n7932), .A2(n6355), .ZN(n6357) );
  AND2_X1 U8017 ( .A1(n7522), .A2(n6358), .ZN(n6359) );
  NAND2_X1 U8018 ( .A1(n7523), .A2(n6359), .ZN(n6360) );
  NAND3_X1 U8019 ( .A1(n6362), .A2(n6361), .A3(n6360), .ZN(n7581) );
  NAND2_X1 U8020 ( .A1(n7751), .A2(n6457), .ZN(n6364) );
  NAND2_X1 U8021 ( .A1(n9222), .A2(n6447), .ZN(n6363) );
  NAND2_X1 U8022 ( .A1(n6364), .A2(n6363), .ZN(n7578) );
  NAND2_X1 U8023 ( .A1(n7751), .A2(n6456), .ZN(n6366) );
  NAND2_X1 U8024 ( .A1(n9222), .A2(n6457), .ZN(n6365) );
  NAND2_X1 U8025 ( .A1(n6366), .A2(n6365), .ZN(n6367) );
  XNOR2_X1 U8026 ( .A(n6367), .B(n6460), .ZN(n7579) );
  INV_X1 U8027 ( .A(n7579), .ZN(n6368) );
  NAND2_X1 U8028 ( .A1(n6379), .A2(n6368), .ZN(n6374) );
  NAND2_X1 U8029 ( .A1(n7581), .A2(n7578), .ZN(n6377) );
  NAND2_X1 U8030 ( .A1(n7778), .A2(n6456), .ZN(n6370) );
  NAND2_X1 U8031 ( .A1(n9221), .A2(n6457), .ZN(n6369) );
  NAND2_X1 U8032 ( .A1(n6370), .A2(n6369), .ZN(n6371) );
  XNOR2_X1 U8033 ( .A(n6371), .B(n6452), .ZN(n6378) );
  INV_X1 U8034 ( .A(n6378), .ZN(n6372) );
  NAND2_X1 U8035 ( .A1(n6374), .A2(n6373), .ZN(n7731) );
  NAND2_X1 U8036 ( .A1(n7778), .A2(n6267), .ZN(n6376) );
  NAND2_X1 U8037 ( .A1(n9221), .A2(n6447), .ZN(n6375) );
  NAND2_X1 U8038 ( .A1(n6376), .A2(n6375), .ZN(n7733) );
  NAND2_X1 U8039 ( .A1(n7731), .A2(n7733), .ZN(n7758) );
  NAND2_X1 U8040 ( .A1(n6377), .A2(n7579), .ZN(n6380) );
  NAND3_X1 U8041 ( .A1(n6380), .A2(n6379), .A3(n6378), .ZN(n7730) );
  NAND2_X1 U8042 ( .A1(n9497), .A2(n6456), .ZN(n6382) );
  NAND2_X1 U8043 ( .A1(n9220), .A2(n6457), .ZN(n6381) );
  NAND2_X1 U8044 ( .A1(n6382), .A2(n6381), .ZN(n6383) );
  XNOR2_X1 U8045 ( .A(n6383), .B(n6460), .ZN(n6385) );
  NOR2_X1 U8046 ( .A1(n7876), .A2(n6462), .ZN(n6384) );
  AOI21_X1 U8047 ( .B1(n9497), .B2(n6457), .A(n6384), .ZN(n6386) );
  NAND2_X1 U8048 ( .A1(n6385), .A2(n6386), .ZN(n6391) );
  INV_X1 U8049 ( .A(n6385), .ZN(n6388) );
  INV_X1 U8050 ( .A(n6386), .ZN(n6387) );
  NAND2_X1 U8051 ( .A1(n6388), .A2(n6387), .ZN(n6389) );
  AND2_X1 U8052 ( .A1(n6391), .A2(n6389), .ZN(n7757) );
  AND2_X1 U8053 ( .A1(n7730), .A2(n7757), .ZN(n6390) );
  NAND2_X1 U8054 ( .A1(n7758), .A2(n6390), .ZN(n7756) );
  NAND2_X1 U8055 ( .A1(n9490), .A2(n6456), .ZN(n6393) );
  NAND2_X1 U8056 ( .A1(n9420), .A2(n6457), .ZN(n6392) );
  NAND2_X1 U8057 ( .A1(n6393), .A2(n6392), .ZN(n6394) );
  XNOR2_X1 U8058 ( .A(n6394), .B(n6452), .ZN(n6396) );
  AND2_X1 U8059 ( .A1(n9420), .A2(n6447), .ZN(n6395) );
  AOI21_X1 U8060 ( .B1(n9490), .B2(n6457), .A(n6395), .ZN(n6397) );
  XNOR2_X1 U8061 ( .A(n6396), .B(n6397), .ZN(n7826) );
  INV_X1 U8062 ( .A(n6396), .ZN(n6398) );
  NAND2_X1 U8063 ( .A1(n6398), .A2(n6397), .ZN(n6399) );
  NAND2_X1 U8064 ( .A1(n9486), .A2(n6456), .ZN(n6401) );
  NAND2_X1 U8065 ( .A1(n9397), .A2(n6457), .ZN(n6400) );
  NAND2_X1 U8066 ( .A1(n6401), .A2(n6400), .ZN(n6402) );
  XNOR2_X1 U8067 ( .A(n6402), .B(n6452), .ZN(n6404) );
  NOR2_X1 U8068 ( .A1(n7909), .A2(n6462), .ZN(n6403) );
  AOI21_X1 U8069 ( .B1(n9486), .B2(n6457), .A(n6403), .ZN(n7883) );
  INV_X1 U8070 ( .A(n6404), .ZN(n6405) );
  NAND2_X1 U8071 ( .A1(n9480), .A2(n6456), .ZN(n6407) );
  NAND2_X1 U8072 ( .A1(n9418), .A2(n6457), .ZN(n6406) );
  NAND2_X1 U8073 ( .A1(n6407), .A2(n6406), .ZN(n6408) );
  XNOR2_X1 U8074 ( .A(n6408), .B(n6452), .ZN(n6411) );
  AOI22_X1 U8075 ( .A1(n9480), .A2(n6267), .B1(n6447), .B2(n9418), .ZN(n6409)
         );
  XNOR2_X1 U8076 ( .A(n6411), .B(n6409), .ZN(n7906) );
  INV_X1 U8077 ( .A(n6409), .ZN(n6410) );
  NAND2_X1 U8078 ( .A1(n7904), .A2(n6412), .ZN(n9178) );
  NAND2_X1 U8079 ( .A1(n9476), .A2(n6456), .ZN(n6414) );
  NAND2_X1 U8080 ( .A1(n9396), .A2(n6457), .ZN(n6413) );
  NAND2_X1 U8081 ( .A1(n6414), .A2(n6413), .ZN(n6415) );
  XNOR2_X1 U8082 ( .A(n6415), .B(n6452), .ZN(n6418) );
  NAND2_X1 U8083 ( .A1(n9476), .A2(n6457), .ZN(n6417) );
  NAND2_X1 U8084 ( .A1(n9396), .A2(n6447), .ZN(n6416) );
  NAND2_X1 U8085 ( .A1(n6417), .A2(n6416), .ZN(n6419) );
  NAND2_X1 U8086 ( .A1(n6418), .A2(n6419), .ZN(n9179) );
  INV_X1 U8087 ( .A(n6418), .ZN(n6421) );
  INV_X1 U8088 ( .A(n6419), .ZN(n6420) );
  NAND2_X1 U8089 ( .A1(n6421), .A2(n6420), .ZN(n9181) );
  NAND2_X1 U8090 ( .A1(n9471), .A2(n6456), .ZN(n6423) );
  NAND2_X1 U8091 ( .A1(n9219), .A2(n6457), .ZN(n6422) );
  NAND2_X1 U8092 ( .A1(n6423), .A2(n6422), .ZN(n6424) );
  XNOR2_X1 U8093 ( .A(n6424), .B(n6452), .ZN(n6425) );
  AOI22_X1 U8094 ( .A1(n9471), .A2(n6457), .B1(n6447), .B2(n9219), .ZN(n6426)
         );
  XNOR2_X1 U8095 ( .A(n6425), .B(n6426), .ZN(n9156) );
  INV_X1 U8096 ( .A(n6425), .ZN(n6427) );
  OAI22_X1 U8097 ( .A1(n8270), .A2(n6444), .B1(n9151), .B2(n6462), .ZN(n6428)
         );
  OAI22_X1 U8098 ( .A1(n8256), .A2(n6445), .B1(n9340), .B2(n6444), .ZN(n6429)
         );
  XNOR2_X1 U8099 ( .A(n6429), .B(n6452), .ZN(n6430) );
  NAND2_X1 U8100 ( .A1(n6431), .A2(n6430), .ZN(n9144) );
  AOI21_X1 U8101 ( .B1(n9146), .B2(n9144), .A(n9143), .ZN(n9170) );
  AOI22_X1 U8102 ( .A1(n9344), .A2(n6267), .B1(n6447), .B2(n9321), .ZN(n6435)
         );
  NAND2_X1 U8103 ( .A1(n9344), .A2(n6456), .ZN(n6433) );
  NAND2_X1 U8104 ( .A1(n9321), .A2(n6457), .ZN(n6432) );
  NAND2_X1 U8105 ( .A1(n6433), .A2(n6432), .ZN(n6434) );
  XNOR2_X1 U8106 ( .A(n6434), .B(n6452), .ZN(n6437) );
  XOR2_X1 U8107 ( .A(n6435), .B(n6437), .Z(n9171) );
  INV_X1 U8108 ( .A(n6435), .ZN(n6436) );
  NAND2_X1 U8109 ( .A1(n5571), .A2(n6456), .ZN(n6439) );
  NAND2_X1 U8110 ( .A1(n9217), .A2(n6457), .ZN(n6438) );
  NAND2_X1 U8111 ( .A1(n6439), .A2(n6438), .ZN(n6440) );
  XNOR2_X1 U8112 ( .A(n6440), .B(n6452), .ZN(n6441) );
  AOI22_X1 U8113 ( .A1(n5571), .A2(n6457), .B1(n6447), .B2(n9217), .ZN(n6442)
         );
  XNOR2_X1 U8114 ( .A(n6441), .B(n6442), .ZN(n9163) );
  INV_X1 U8115 ( .A(n6441), .ZN(n6443) );
  OAI22_X1 U8116 ( .A1(n9307), .A2(n6445), .B1(n9135), .B2(n6444), .ZN(n6446)
         );
  XNOR2_X1 U8117 ( .A(n6446), .B(n6452), .ZN(n6448) );
  AOI22_X1 U8118 ( .A1(n9443), .A2(n6457), .B1(n6447), .B2(n9320), .ZN(n6449)
         );
  XNOR2_X1 U8119 ( .A(n6448), .B(n6449), .ZN(n9205) );
  AOI22_X1 U8120 ( .A1(n9438), .A2(n6456), .B1(n6267), .B2(n9216), .ZN(n6453)
         );
  XNOR2_X1 U8121 ( .A(n6453), .B(n6452), .ZN(n9130) );
  NOR2_X1 U8122 ( .A1(n9312), .A2(n6462), .ZN(n6454) );
  AOI21_X1 U8123 ( .B1(n9438), .B2(n6267), .A(n6454), .ZN(n9131) );
  NAND2_X1 U8124 ( .A1(n9130), .A2(n9131), .ZN(n6455) );
  NAND2_X1 U8125 ( .A1(n9434), .A2(n6456), .ZN(n6459) );
  NAND2_X1 U8126 ( .A1(n5568), .A2(n6457), .ZN(n6458) );
  NAND2_X1 U8127 ( .A1(n6459), .A2(n6458), .ZN(n6461) );
  XNOR2_X1 U8128 ( .A(n6461), .B(n6460), .ZN(n6465) );
  NOR2_X1 U8129 ( .A1(n9139), .A2(n6462), .ZN(n6463) );
  AOI21_X1 U8130 ( .B1(n9434), .B2(n6267), .A(n6463), .ZN(n6464) );
  XNOR2_X1 U8131 ( .A(n6465), .B(n6464), .ZN(n6492) );
  INV_X1 U8132 ( .A(n6492), .ZN(n6471) );
  OR2_X1 U8133 ( .A1(n9130), .A2(n9131), .ZN(n6472) );
  NAND2_X1 U8134 ( .A1(n6466), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U8135 ( .A1(n6583), .A2(n6467), .ZN(n6468) );
  NAND2_X1 U8136 ( .A1(n6468), .A2(n6585), .ZN(n6882) );
  OR2_X1 U8137 ( .A1(n9791), .A2(n6882), .ZN(n6476) );
  INV_X1 U8138 ( .A(n9794), .ZN(n6469) );
  NOR2_X1 U8139 ( .A1(n6476), .A2(n6469), .ZN(n6485) );
  NOR2_X1 U8140 ( .A1(n9500), .A2(n8127), .ZN(n6470) );
  NAND2_X1 U8141 ( .A1(n6485), .A2(n6470), .ZN(n9201) );
  INV_X1 U8142 ( .A(n9201), .ZN(n9204) );
  INV_X1 U8143 ( .A(n6472), .ZN(n6473) );
  NAND3_X1 U8144 ( .A1(n6492), .A2(n9204), .A3(n6473), .ZN(n6490) );
  NAND3_X1 U8145 ( .A1(n6476), .A2(n9794), .A3(n9772), .ZN(n6481) );
  NAND2_X1 U8146 ( .A1(n6481), .A2(n7001), .ZN(n9165) );
  NOR2_X1 U8147 ( .A1(n9165), .A2(n9831), .ZN(n9199) );
  INV_X1 U8148 ( .A(n6476), .ZN(n7002) );
  NAND2_X1 U8149 ( .A1(n9794), .A2(n6525), .ZN(n6475) );
  NOR2_X1 U8150 ( .A1(n6475), .A2(n6668), .ZN(n8249) );
  NAND2_X1 U8151 ( .A1(n7002), .A2(n8249), .ZN(n9207) );
  INV_X1 U8152 ( .A(n9297), .ZN(n6483) );
  NAND2_X1 U8153 ( .A1(n6476), .A2(n9831), .ZN(n6479) );
  NAND4_X1 U8154 ( .A1(n6479), .A2(n6498), .A3(n6478), .A4(n6477), .ZN(n6480)
         );
  NAND2_X1 U8155 ( .A1(n6480), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6482) );
  NAND2_X1 U8156 ( .A1(n6482), .A2(n6481), .ZN(n9211) );
  AOI22_X1 U8157 ( .A1(n6483), .A2(n9211), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6487) );
  NOR2_X1 U8158 ( .A1(n6668), .A2(n6525), .ZN(n6484) );
  NAND2_X1 U8159 ( .A1(n6485), .A2(n6484), .ZN(n9208) );
  INV_X1 U8160 ( .A(n9208), .ZN(n9183) );
  NAND2_X1 U8161 ( .A1(n9291), .A2(n9183), .ZN(n6486) );
  OAI211_X1 U8162 ( .C1(n9312), .C2(n9207), .A(n6487), .B(n6486), .ZN(n6488)
         );
  AOI21_X1 U8163 ( .B1(n9434), .B2(n9199), .A(n6488), .ZN(n6489) );
  AOI21_X1 U8164 ( .B1(n6493), .B2(n4942), .A(n6491), .ZN(n6495) );
  NAND2_X1 U8165 ( .A1(n6495), .A2(n6494), .ZN(P1_U3218) );
  NAND2_X1 U8166 ( .A1(n6497), .A2(n6498), .ZN(n6694) );
  INV_X1 U8167 ( .A(n6498), .ZN(n7299) );
  OR2_X1 U8168 ( .A1(n6499), .A2(n7299), .ZN(n6500) );
  NAND2_X1 U8169 ( .A1(n6694), .A2(n6500), .ZN(n9624) );
  OR2_X1 U8170 ( .A1(n9624), .A2(n6501), .ZN(n6502) );
  NAND2_X1 U8171 ( .A1(n6502), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  OR2_X2 U8172 ( .A1(n6694), .A2(P1_U3084), .ZN(n9234) );
  INV_X1 U8173 ( .A(n9234), .ZN(P1_U4006) );
  OR2_X1 U8174 ( .A1(n6503), .A2(P2_U3152), .ZN(n6712) );
  NOR2_X2 U8175 ( .A1(n6712), .A2(n6588), .ZN(P2_U3966) );
  INV_X1 U8176 ( .A(n6504), .ZN(n6505) );
  AOI211_X1 U8177 ( .C1(n6507), .C2(n6506), .A(n8643), .B(n6505), .ZN(n6511)
         );
  INV_X1 U8178 ( .A(n9079), .ZN(n7816) );
  NOR2_X1 U8179 ( .A1(n7816), .A2(n8619), .ZN(n6510) );
  INV_X1 U8180 ( .A(n8624), .ZN(n8613) );
  INV_X1 U8181 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10065) );
  OAI22_X1 U8182 ( .A1(n8613), .A2(n8779), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10065), .ZN(n6509) );
  INV_X1 U8183 ( .A(n8628), .ZN(n8614) );
  OAI22_X1 U8184 ( .A1(n8614), .A2(n7896), .B1(n8640), .B2(n7817), .ZN(n6508)
         );
  OR4_X1 U8185 ( .A1(n6511), .A2(n6510), .A3(n6509), .A4(n6508), .ZN(P2_U3230)
         );
  AND2_X1 U8186 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7937) );
  MUX2_X1 U8187 ( .A(n7384), .B(P1_REG2_REG_7__SCAN_IN), .S(n6540), .Z(n6679)
         );
  NOR2_X1 U8188 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9643), .ZN(n6519) );
  INV_X1 U8189 ( .A(n9629), .ZN(n9628) );
  MUX2_X1 U8190 ( .A(n6512), .B(P1_REG2_REG_2__SCAN_IN), .S(n9629), .Z(n6516)
         );
  AND2_X1 U8191 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6514) );
  OR2_X1 U8192 ( .A1(n6650), .A2(n6513), .ZN(n9630) );
  NAND2_X1 U8193 ( .A1(n9631), .A2(n9630), .ZN(n6515) );
  INV_X1 U8194 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7217) );
  MUX2_X1 U8195 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n7217), .S(n6640), .Z(n6634)
         );
  OAI21_X1 U8196 ( .B1(n6640), .B2(n7217), .A(n6637), .ZN(n6703) );
  MUX2_X1 U8197 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6517), .S(n6704), .Z(n6702)
         );
  MUX2_X1 U8198 ( .A(n6518), .B(P1_REG2_REG_5__SCAN_IN), .S(n9643), .Z(n9646)
         );
  MUX2_X1 U8199 ( .A(n6520), .B(P1_REG2_REG_6__SCAN_IN), .S(n6662), .Z(n6658)
         );
  NAND2_X1 U8200 ( .A1(n6659), .A2(n6658), .ZN(n6657) );
  OAI21_X1 U8201 ( .B1(n6662), .B2(n6520), .A(n6657), .ZN(n6680) );
  NOR2_X1 U8202 ( .A1(n6679), .A2(n6680), .ZN(n6678) );
  AOI21_X1 U8203 ( .B1(n6681), .B2(n7384), .A(n6678), .ZN(n9662) );
  NAND2_X1 U8204 ( .A1(n9658), .A2(n9659), .ZN(n6521) );
  AOI22_X1 U8205 ( .A1(n9662), .A2(n6521), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n9656), .ZN(n6527) );
  NAND2_X1 U8206 ( .A1(n6815), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6522) );
  OAI21_X1 U8207 ( .B1(n6815), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6522), .ZN(
        n6526) );
  NOR2_X1 U8208 ( .A1(n6527), .A2(n6526), .ZN(n6814) );
  INV_X1 U8209 ( .A(n9624), .ZN(n6523) );
  AND2_X1 U8210 ( .A1(n6523), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6545) );
  INV_X1 U8211 ( .A(n6545), .ZN(n6524) );
  NOR2_X1 U8212 ( .A1(n6524), .A2(n9619), .ZN(n6547) );
  AND2_X1 U8213 ( .A1(n6547), .A2(n6525), .ZN(n9758) );
  INV_X1 U8214 ( .A(n9758), .ZN(n9723) );
  AOI211_X1 U8215 ( .C1(n6527), .C2(n6526), .A(n6814), .B(n9723), .ZN(n6551)
         );
  INV_X1 U8216 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9847) );
  MUX2_X1 U8217 ( .A(n9847), .B(P1_REG1_REG_8__SCAN_IN), .S(n9658), .Z(n9664)
         );
  INV_X1 U8218 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6528) );
  AND2_X1 U8219 ( .A1(n6662), .A2(n6528), .ZN(n6539) );
  NAND2_X1 U8220 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9643), .ZN(n6537) );
  MUX2_X1 U8221 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6529), .S(n9643), .Z(n9649)
         );
  INV_X1 U8222 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6536) );
  MUX2_X1 U8223 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6536), .S(n6704), .Z(n6698)
         );
  INV_X1 U8224 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6535) );
  MUX2_X1 U8225 ( .A(n6530), .B(P1_REG1_REG_2__SCAN_IN), .S(n9629), .Z(n9639)
         );
  INV_X1 U8226 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6531) );
  MUX2_X1 U8227 ( .A(n6531), .B(P1_REG1_REG_1__SCAN_IN), .S(n6650), .Z(n6642)
         );
  AND2_X1 U8228 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6643) );
  NAND2_X1 U8229 ( .A1(n6642), .A2(n6643), .ZN(n6641) );
  OR2_X1 U8230 ( .A1(n6650), .A2(n6531), .ZN(n6532) );
  NAND2_X1 U8231 ( .A1(n6641), .A2(n6532), .ZN(n9640) );
  NAND2_X1 U8232 ( .A1(n9639), .A2(n9640), .ZN(n9638) );
  OR2_X1 U8233 ( .A1(n9629), .A2(n6530), .ZN(n6628) );
  NAND2_X1 U8234 ( .A1(n9638), .A2(n6628), .ZN(n6534) );
  MUX2_X1 U8235 ( .A(n6535), .B(P1_REG1_REG_3__SCAN_IN), .S(n6640), .Z(n6533)
         );
  NAND2_X1 U8236 ( .A1(n6534), .A2(n6533), .ZN(n6631) );
  OAI21_X1 U8237 ( .B1(n6640), .B2(n6535), .A(n6631), .ZN(n6699) );
  NOR2_X1 U8238 ( .A1(n6698), .A2(n6699), .ZN(n6697) );
  AOI21_X1 U8239 ( .B1(n6704), .B2(n6536), .A(n6697), .ZN(n9650) );
  NAND2_X1 U8240 ( .A1(n9649), .A2(n9650), .ZN(n9648) );
  NAND2_X1 U8241 ( .A1(n6537), .A2(n9648), .ZN(n6654) );
  NOR2_X1 U8242 ( .A1(n6662), .A2(n6528), .ZN(n6538) );
  OR2_X1 U8243 ( .A1(n6539), .A2(n6538), .ZN(n6653) );
  NOR2_X1 U8244 ( .A1(n6654), .A2(n6653), .ZN(n6652) );
  NOR2_X1 U8245 ( .A1(n6539), .A2(n6652), .ZN(n6677) );
  INV_X1 U8246 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9845) );
  AOI22_X1 U8247 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6681), .B1(n6540), .B2(
        n9845), .ZN(n6676) );
  NOR2_X1 U8248 ( .A1(n6677), .A2(n6676), .ZN(n6675) );
  NOR2_X1 U8249 ( .A1(n6540), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6541) );
  NOR2_X1 U8250 ( .A1(n6675), .A2(n6541), .ZN(n9665) );
  NAND2_X1 U8251 ( .A1(n9664), .A2(n9665), .ZN(n9663) );
  OAI21_X1 U8252 ( .B1(n9847), .B2(n9658), .A(n9663), .ZN(n6543) );
  INV_X1 U8253 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9850) );
  INV_X1 U8254 ( .A(n6815), .ZN(n6558) );
  AOI22_X1 U8255 ( .A1(n6815), .A2(n9850), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6558), .ZN(n6542) );
  NOR2_X1 U8256 ( .A1(n6543), .A2(n6542), .ZN(n6806) );
  AOI21_X1 U8257 ( .B1(n6543), .B2(n6542), .A(n6806), .ZN(n6546) );
  NOR2_X1 U8258 ( .A1(n4384), .A2(n8248), .ZN(n6544) );
  NAND2_X1 U8259 ( .A1(n6545), .A2(n6544), .ZN(n9765) );
  NOR2_X1 U8260 ( .A1(n6546), .A2(n9765), .ZN(n6550) );
  AND2_X1 U8261 ( .A1(n6547), .A2(n4384), .ZN(n9753) );
  INV_X1 U8262 ( .A(n9753), .ZN(n6876) );
  INV_X1 U8263 ( .A(n6694), .ZN(n6548) );
  NOR2_X1 U8264 ( .A1(P1_U3083), .A2(n6548), .ZN(n9655) );
  INV_X1 U8265 ( .A(n9655), .ZN(n9769) );
  INV_X1 U8266 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10274) );
  OAI22_X1 U8267 ( .A1(n6558), .A2(n6876), .B1(n9769), .B2(n10274), .ZN(n6549)
         );
  OR4_X1 U8268 ( .A1(n7937), .A2(n6551), .A3(n6550), .A4(n6549), .ZN(P1_U3250)
         );
  XNOR2_X1 U8269 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OR2_X1 U8270 ( .A1(n6553), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7924) );
  AND2_X1 U8271 ( .A1(n6553), .A2(P1_U3084), .ZN(n9535) );
  OAI222_X1 U8272 ( .A1(n7924), .A2(n6552), .B1(n7920), .B2(n6555), .C1(
        P1_U3084), .C2(n6650), .ZN(P1_U3352) );
  NAND2_X1 U8273 ( .A1(n6553), .A2(P2_U3152), .ZN(n8511) );
  INV_X1 U8274 ( .A(n8511), .ZN(n6824) );
  INV_X1 U8275 ( .A(n6824), .ZN(n10258) );
  OR2_X1 U8276 ( .A1(n6553), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7928) );
  OAI222_X1 U8277 ( .A1(n10258), .A2(n6554), .B1(n7928), .B2(n6564), .C1(
        P2_U3152), .C2(n6910), .ZN(P2_U3350) );
  OAI222_X1 U8278 ( .A1(n10258), .A2(n6556), .B1(n7928), .B2(n6555), .C1(
        P2_U3152), .C2(n6727), .ZN(P2_U3357) );
  OAI222_X1 U8279 ( .A1(n10258), .A2(n6557), .B1(n7928), .B2(n5775), .C1(
        P2_U3152), .C2(n6750), .ZN(P2_U3355) );
  OAI222_X1 U8280 ( .A1(n7924), .A2(n10132), .B1(n7920), .B2(n6574), .C1(n6558), .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U8281 ( .A(n7924), .ZN(n6664) );
  INV_X1 U8282 ( .A(n6664), .ZN(n9531) );
  OAI222_X1 U8283 ( .A1(n9531), .A2(n6559), .B1(n7920), .B2(n5775), .C1(
        P1_U3084), .C2(n6640), .ZN(P1_U3350) );
  OAI222_X1 U8284 ( .A1(n9531), .A2(n6560), .B1(n7920), .B2(n6572), .C1(
        P1_U3084), .C2(n6681), .ZN(P1_U3346) );
  OAI222_X1 U8285 ( .A1(n9531), .A2(n6561), .B1(n7920), .B2(n5835), .C1(
        P1_U3084), .C2(n6662), .ZN(P1_U3347) );
  OAI222_X1 U8286 ( .A1(n9531), .A2(n6563), .B1(n7920), .B2(n6567), .C1(
        P1_U3084), .C2(n6562), .ZN(P1_U3348) );
  OAI222_X1 U8287 ( .A1(n9531), .A2(n10115), .B1(n7920), .B2(n6564), .C1(
        P1_U3084), .C2(n9658), .ZN(P1_U3345) );
  OAI222_X1 U8288 ( .A1(n9531), .A2(n6565), .B1(n7920), .B2(n6569), .C1(
        P1_U3084), .C2(n9629), .ZN(P1_U3351) );
  OAI222_X1 U8289 ( .A1(n9531), .A2(n6566), .B1(n7920), .B2(n10255), .C1(
        P1_U3084), .C2(n6704), .ZN(P1_U3349) );
  INV_X1 U8290 ( .A(n7928), .ZN(n9127) );
  INV_X1 U8291 ( .A(n9127), .ZN(n10256) );
  OAI222_X1 U8292 ( .A1(n10258), .A2(n6568), .B1(n10256), .B2(n6567), .C1(
        P2_U3152), .C2(n6738), .ZN(P2_U3353) );
  OAI222_X1 U8293 ( .A1(n10258), .A2(n6570), .B1(n10256), .B2(n6569), .C1(
        P2_U3152), .C2(n6728), .ZN(P2_U3356) );
  OAI222_X1 U8294 ( .A1(n10258), .A2(n6571), .B1(n10256), .B2(n5835), .C1(
        P2_U3152), .C2(n6786), .ZN(P2_U3352) );
  OAI222_X1 U8295 ( .A1(n10258), .A2(n6573), .B1(n10256), .B2(n6572), .C1(
        P2_U3152), .C2(n6803), .ZN(P2_U3351) );
  OAI222_X1 U8296 ( .A1(n8511), .A2(n6575), .B1(n10256), .B2(n6574), .C1(n6991), .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8297 ( .A(n6576), .ZN(n6582) );
  AOI22_X1 U8298 ( .A1(n8672), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n6824), .ZN(n6577) );
  OAI21_X1 U8299 ( .B1(n6582), .B2(n10256), .A(n6577), .ZN(P2_U3347) );
  INV_X1 U8300 ( .A(n6578), .ZN(n6580) );
  INV_X1 U8301 ( .A(n6871), .ZN(n6808) );
  OAI222_X1 U8302 ( .A1(n7924), .A2(n6579), .B1(n7920), .B2(n6580), .C1(n6808), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U8303 ( .A(n7451), .ZN(n7459) );
  OAI222_X1 U8304 ( .A1(n8511), .A2(n6581), .B1(n7928), .B2(n6580), .C1(n7459), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8305 ( .A(n9248), .ZN(n6875) );
  OAI222_X1 U8306 ( .A1(n7924), .A2(n10116), .B1(n7920), .B2(n6582), .C1(n6875), .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U8307 ( .A(n6583), .ZN(n6584) );
  NAND2_X1 U8308 ( .A1(n6584), .A2(n9794), .ZN(n9790) );
  INV_X1 U8309 ( .A(n9790), .ZN(n9789) );
  OAI21_X1 U8310 ( .B1(n9789), .B2(P1_D_REG_0__SCAN_IN), .A(n6585), .ZN(n6586)
         );
  OAI21_X1 U8311 ( .B1(n9794), .B2(n6587), .A(n6586), .ZN(P1_U3440) );
  AND2_X1 U8312 ( .A1(n6588), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8496) );
  INV_X1 U8313 ( .A(n8496), .ZN(n8500) );
  NAND2_X1 U8314 ( .A1(n9865), .A2(n8500), .ZN(n6589) );
  NAND2_X1 U8315 ( .A1(n6590), .A2(n6589), .ZN(n6593) );
  OR2_X1 U8316 ( .A1(n9865), .A2(n6591), .ZN(n6592) );
  NAND2_X1 U8317 ( .A1(n6593), .A2(n6592), .ZN(n9854) );
  NOR2_X1 U8318 ( .A1(n9854), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8319 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6598) );
  INV_X1 U8320 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n10146) );
  NAND2_X1 U8321 ( .A1(n5783), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6596) );
  NAND2_X1 U8322 ( .A1(n6594), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6595) );
  OAI211_X1 U8323 ( .C1(n5753), .C2(n10146), .A(n6596), .B(n6595), .ZN(n8302)
         );
  NAND2_X1 U8324 ( .A1(n8302), .A2(P2_U3966), .ZN(n6597) );
  OAI21_X1 U8325 ( .B1(P2_U3966), .B2(n6598), .A(n6597), .ZN(P2_U3583) );
  INV_X1 U8326 ( .A(n6599), .ZN(n6601) );
  AOI22_X1 U8327 ( .A1(n9675), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n6664), .ZN(n6600) );
  OAI21_X1 U8328 ( .B1(n6601), .B2(n7920), .A(n6600), .ZN(P1_U3341) );
  INV_X1 U8329 ( .A(n7599), .ZN(n7595) );
  OAI222_X1 U8330 ( .A1(n8511), .A2(n6602), .B1(n7928), .B2(n6601), .C1(
        P2_U3152), .C2(n7595), .ZN(P2_U3346) );
  INV_X1 U8331 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6604) );
  NAND2_X1 U8332 ( .A1(n8072), .A2(P1_U4006), .ZN(n6603) );
  OAI21_X1 U8333 ( .B1(P1_U4006), .B2(n6604), .A(n6603), .ZN(P1_U3586) );
  INV_X1 U8334 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6605) );
  OR2_X1 U8335 ( .A1(n6606), .A2(n6605), .ZN(n6612) );
  INV_X1 U8336 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6607) );
  OR2_X1 U8337 ( .A1(n5753), .A2(n6607), .ZN(n6611) );
  INV_X1 U8338 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6608) );
  OR2_X1 U8339 ( .A1(n6609), .A2(n6608), .ZN(n6610) );
  AND3_X1 U8340 ( .A1(n6612), .A2(n6611), .A3(n6610), .ZN(n8774) );
  NAND2_X1 U8341 ( .A1(n8665), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6613) );
  OAI21_X1 U8342 ( .B1(n8774), .B2(n8665), .A(n6613), .ZN(P2_U3582) );
  INV_X1 U8343 ( .A(n6614), .ZN(n6616) );
  AOI22_X1 U8344 ( .A1(n9684), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n6664), .ZN(n6615) );
  OAI21_X1 U8345 ( .B1(n6616), .B2(n7920), .A(n6615), .ZN(P1_U3340) );
  INV_X1 U8346 ( .A(n7655), .ZN(n7651) );
  OAI222_X1 U8347 ( .A1(n8511), .A2(n9993), .B1(n7928), .B2(n6616), .C1(n7651), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8348 ( .A(n6617), .ZN(n6619) );
  INV_X1 U8349 ( .A(n8681), .ZN(n8687) );
  OAI222_X1 U8350 ( .A1(n8511), .A2(n6618), .B1(n7928), .B2(n6619), .C1(n8687), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  OAI222_X1 U8351 ( .A1(n7924), .A2(n6620), .B1(n7920), .B2(n6619), .C1(n9255), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8352 ( .A(n6621), .ZN(n6622) );
  INV_X1 U8353 ( .A(n8701), .ZN(n8694) );
  OAI222_X1 U8354 ( .A1(n8511), .A2(n10094), .B1(n10256), .B2(n6622), .C1(
        P2_U3152), .C2(n8694), .ZN(P2_U3343) );
  INV_X1 U8355 ( .A(n9716), .ZN(n9257) );
  OAI222_X1 U8356 ( .A1(n7924), .A2(n6623), .B1(n7920), .B2(n6622), .C1(
        P1_U3084), .C2(n9257), .ZN(P1_U3338) );
  INV_X1 U8357 ( .A(n6624), .ZN(n6627) );
  AOI22_X1 U8358 ( .A1(n9728), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n6664), .ZN(n6625) );
  OAI21_X1 U8359 ( .B1(n6627), .B2(n7920), .A(n6625), .ZN(P1_U3337) );
  AOI22_X1 U8360 ( .A1(n8718), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n6824), .ZN(n6626) );
  OAI21_X1 U8361 ( .B1(n6627), .B2(n10256), .A(n6626), .ZN(P2_U3342) );
  MUX2_X1 U8362 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6535), .S(n6640), .Z(n6629)
         );
  NAND3_X1 U8363 ( .A1(n6629), .A2(n9638), .A3(n6628), .ZN(n6630) );
  NAND2_X1 U8364 ( .A1(n6631), .A2(n6630), .ZN(n6632) );
  NAND2_X1 U8365 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6975) );
  OAI21_X1 U8366 ( .B1(n9765), .B2(n6632), .A(n6975), .ZN(n6633) );
  AOI21_X1 U8367 ( .B1(n9655), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6633), .ZN(
        n6639) );
  NAND2_X1 U8368 ( .A1(n6635), .A2(n6634), .ZN(n6636) );
  NAND3_X1 U8369 ( .A1(n9758), .A2(n6637), .A3(n6636), .ZN(n6638) );
  OAI211_X1 U8370 ( .C1(n6876), .C2(n6640), .A(n6639), .B(n6638), .ZN(P1_U3244) );
  OAI21_X1 U8371 ( .B1(n6643), .B2(n6642), .A(n6641), .ZN(n6645) );
  NAND2_X1 U8372 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(P1_U3084), .ZN(n6644) );
  OAI21_X1 U8373 ( .B1(n9765), .B2(n6645), .A(n6644), .ZN(n6646) );
  AOI21_X1 U8374 ( .B1(n9655), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n6646), .ZN(
        n6649) );
  NAND2_X1 U8375 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6691) );
  OAI211_X1 U8376 ( .C1(n6514), .C2(n6647), .A(n9758), .B(n9631), .ZN(n6648)
         );
  OAI211_X1 U8377 ( .C1(n6876), .C2(n6650), .A(n6649), .B(n6648), .ZN(P1_U3242) );
  NOR2_X1 U8378 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6651), .ZN(n7424) );
  AOI21_X1 U8379 ( .B1(n6654), .B2(n6653), .A(n6652), .ZN(n6655) );
  NOR2_X1 U8380 ( .A1(n9765), .A2(n6655), .ZN(n6656) );
  AOI211_X1 U8381 ( .C1(n9655), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n7424), .B(
        n6656), .ZN(n6661) );
  OAI211_X1 U8382 ( .C1(n6659), .C2(n6658), .A(n9758), .B(n6657), .ZN(n6660)
         );
  OAI211_X1 U8383 ( .C1(n6876), .C2(n6662), .A(n6661), .B(n6660), .ZN(P1_U3247) );
  INV_X1 U8384 ( .A(n6663), .ZN(n6666) );
  AOI22_X1 U8385 ( .A1(n9739), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n6664), .ZN(n6665) );
  OAI21_X1 U8386 ( .B1(n6666), .B2(n7920), .A(n6665), .ZN(P1_U3336) );
  INV_X1 U8387 ( .A(n8729), .ZN(n8735) );
  OAI222_X1 U8388 ( .A1(n8511), .A2(n6667), .B1(n10256), .B2(n6666), .C1(n8735), .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8389 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6674) );
  XNOR2_X1 U8390 ( .A(n9235), .B(n7130), .ZN(n8091) );
  INV_X1 U8391 ( .A(n6668), .ZN(n6670) );
  INV_X1 U8392 ( .A(n6672), .ZN(n6669) );
  NOR3_X1 U8393 ( .A1(n8091), .A2(n6670), .A3(n6669), .ZN(n6671) );
  AOI21_X1 U8394 ( .B1(n9417), .B2(n6258), .A(n6671), .ZN(n7125) );
  OAI21_X1 U8395 ( .B1(n8210), .B2(n6672), .A(n7125), .ZN(n9513) );
  NAND2_X1 U8396 ( .A1(n9513), .A2(n9840), .ZN(n6673) );
  OAI21_X1 U8397 ( .B1(n9840), .B2(n6674), .A(n6673), .ZN(P1_U3454) );
  AOI21_X1 U8398 ( .B1(n6677), .B2(n6676), .A(n6675), .ZN(n6686) );
  AOI21_X1 U8399 ( .B1(n6680), .B2(n6679), .A(n6678), .ZN(n6682) );
  OAI22_X1 U8400 ( .A1(n6682), .A2(n9723), .B1(n6876), .B2(n6681), .ZN(n6683)
         );
  INV_X1 U8401 ( .A(n6683), .ZN(n6685) );
  NOR2_X1 U8402 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5094), .ZN(n7037) );
  AOI21_X1 U8403 ( .B1(n9655), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n7037), .ZN(
        n6684) );
  OAI211_X1 U8404 ( .C1(n6686), .C2(n9765), .A(n6685), .B(n6684), .ZN(P1_U3248) );
  OR2_X1 U8405 ( .A1(n6688), .A2(n6687), .ZN(n6689) );
  NAND2_X1 U8406 ( .A1(n6690), .A2(n6689), .ZN(n7012) );
  MUX2_X1 U8407 ( .A(n7012), .B(n6691), .S(n8248), .Z(n6696) );
  NOR2_X1 U8408 ( .A1(n9619), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6692) );
  OR2_X1 U8409 ( .A1(n4384), .A2(n6692), .ZN(n9621) );
  INV_X1 U8410 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10074) );
  NAND2_X1 U8411 ( .A1(n9621), .A2(n10074), .ZN(n6693) );
  NAND2_X1 U8412 ( .A1(n6693), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9623) );
  NOR2_X1 U8413 ( .A1(n9623), .A2(n6694), .ZN(n6695) );
  OAI21_X1 U8414 ( .B1(n6696), .B2(n4384), .A(n6695), .ZN(n9637) );
  AOI21_X1 U8415 ( .B1(n6699), .B2(n6698), .A(n6697), .ZN(n6700) );
  NAND2_X1 U8416 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n6963) );
  OAI21_X1 U8417 ( .B1(n9765), .B2(n6700), .A(n6963), .ZN(n6707) );
  AOI21_X1 U8418 ( .B1(n6703), .B2(n6702), .A(n6701), .ZN(n6705) );
  OAI22_X1 U8419 ( .A1(n6705), .A2(n9723), .B1(n6876), .B2(n6704), .ZN(n6706)
         );
  AOI211_X1 U8420 ( .C1(n9655), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n6707), .B(
        n6706), .ZN(n6708) );
  NAND2_X1 U8421 ( .A1(n9637), .A2(n6708), .ZN(P1_U3245) );
  NAND2_X1 U8422 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9539) );
  AOI21_X1 U8423 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n9542), .A(n9538), .ZN(
        n9552) );
  AOI22_X1 U8424 ( .A1(n9554), .A2(n5752), .B1(P2_REG2_REG_2__SCAN_IN), .B2(
        n6728), .ZN(n9551) );
  NOR2_X1 U8425 ( .A1(n9552), .A2(n9551), .ZN(n9550) );
  NAND2_X1 U8426 ( .A1(n6723), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6709) );
  OAI21_X1 U8427 ( .B1(n6723), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6709), .ZN(
        n6743) );
  NOR2_X1 U8428 ( .A1(n6742), .A2(n6743), .ZN(n6741) );
  AOI21_X1 U8429 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n6723), .A(n6741), .ZN(
        n6755) );
  NAND2_X1 U8430 ( .A1(n6721), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6710) );
  OAI21_X1 U8431 ( .B1(n6721), .B2(P2_REG2_REG_4__SCAN_IN), .A(n6710), .ZN(
        n6754) );
  NOR2_X1 U8432 ( .A1(n6755), .A2(n6754), .ZN(n6753) );
  AOI21_X1 U8433 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n6721), .A(n6753), .ZN(
        n6718) );
  NAND2_X1 U8434 ( .A1(n6769), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6711) );
  OAI21_X1 U8435 ( .B1(n6769), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6711), .ZN(
        n6717) );
  NOR2_X1 U8436 ( .A1(n6718), .A2(n6717), .ZN(n6764) );
  OAI211_X1 U8437 ( .C1(n9865), .C2(n6843), .A(n8500), .B(n6712), .ZN(n6714)
         );
  NAND2_X1 U8438 ( .A1(n6714), .A2(n6713), .ZN(n6732) );
  NAND2_X1 U8439 ( .A1(n8665), .A2(n6732), .ZN(n6719) );
  INV_X1 U8440 ( .A(n6715), .ZN(n8498) );
  NAND3_X1 U8441 ( .A1(n6719), .A2(n6716), .A3(n8498), .ZN(n9549) );
  AOI211_X1 U8442 ( .C1(n6718), .C2(n6717), .A(n6764), .B(n9549), .ZN(n6740)
         );
  AND2_X1 U8443 ( .A1(n6233), .A2(n6719), .ZN(n9555) );
  INV_X1 U8444 ( .A(n9555), .ZN(n9857) );
  INV_X1 U8445 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10047) );
  NOR2_X1 U8446 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10047), .ZN(n6720) );
  AOI21_X1 U8447 ( .B1(n9854), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6720), .ZN(
        n6737) );
  NAND2_X1 U8448 ( .A1(n6721), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6730) );
  MUX2_X1 U8449 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6722), .S(n6721), .Z(n6758)
         );
  NAND2_X1 U8450 ( .A1(n6723), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6729) );
  MUX2_X1 U8451 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6724), .S(n6723), .Z(n6746)
         );
  MUX2_X1 U8452 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6725), .S(n9554), .Z(n9557)
         );
  MUX2_X1 U8453 ( .A(n6726), .B(P2_REG1_REG_1__SCAN_IN), .S(n6727), .Z(n9544)
         );
  NAND3_X1 U8454 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n9544), .ZN(n9543) );
  OAI21_X1 U8455 ( .B1(n6727), .B2(n6726), .A(n9543), .ZN(n9558) );
  NAND2_X1 U8456 ( .A1(n9557), .A2(n9558), .ZN(n9556) );
  OAI21_X1 U8457 ( .B1(n6728), .B2(n6725), .A(n9556), .ZN(n6747) );
  NAND2_X1 U8458 ( .A1(n6746), .A2(n6747), .ZN(n6745) );
  NAND2_X1 U8459 ( .A1(n6729), .A2(n6745), .ZN(n6759) );
  NAND2_X1 U8460 ( .A1(n6758), .A2(n6759), .ZN(n6757) );
  NAND2_X1 U8461 ( .A1(n6730), .A2(n6757), .ZN(n6735) );
  MUX2_X1 U8462 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6731), .S(n6769), .Z(n6734)
         );
  INV_X1 U8463 ( .A(n6732), .ZN(n6733) );
  AND2_X1 U8464 ( .A1(n6715), .A2(n6733), .ZN(n9853) );
  NAND2_X1 U8465 ( .A1(n6734), .A2(n6735), .ZN(n6770) );
  OAI211_X1 U8466 ( .C1(n6735), .C2(n6734), .A(n9853), .B(n6770), .ZN(n6736)
         );
  OAI211_X1 U8467 ( .C1(n9857), .C2(n6738), .A(n6737), .B(n6736), .ZN(n6739)
         );
  OR2_X1 U8468 ( .A1(n6740), .A2(n6739), .ZN(P2_U3250) );
  AOI211_X1 U8469 ( .C1(n6743), .C2(n6742), .A(n6741), .B(n9549), .ZN(n6752)
         );
  NOR2_X1 U8470 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5785), .ZN(n6744) );
  AOI21_X1 U8471 ( .B1(n9854), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6744), .ZN(
        n6749) );
  OAI211_X1 U8472 ( .C1(n6747), .C2(n6746), .A(n9853), .B(n6745), .ZN(n6748)
         );
  OAI211_X1 U8473 ( .C1(n9857), .C2(n6750), .A(n6749), .B(n6748), .ZN(n6751)
         );
  OR2_X1 U8474 ( .A1(n6752), .A2(n6751), .ZN(P2_U3248) );
  AOI211_X1 U8475 ( .C1(n6755), .C2(n6754), .A(n6753), .B(n9549), .ZN(n6763)
         );
  NAND2_X1 U8476 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n6934) );
  INV_X1 U8477 ( .A(n6934), .ZN(n6756) );
  AOI21_X1 U8478 ( .B1(n9854), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6756), .ZN(
        n6761) );
  OAI211_X1 U8479 ( .C1(n6759), .C2(n6758), .A(n9853), .B(n6757), .ZN(n6760)
         );
  OAI211_X1 U8480 ( .C1(n9857), .C2(n10254), .A(n6761), .B(n6760), .ZN(n6762)
         );
  OR2_X1 U8481 ( .A1(n6763), .A2(n6762), .ZN(P2_U3249) );
  INV_X1 U8482 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6765) );
  XNOR2_X1 U8483 ( .A(n6786), .B(n6765), .ZN(n6766) );
  AOI211_X1 U8484 ( .C1(n6767), .C2(n6766), .A(n6778), .B(n9549), .ZN(n6777)
         );
  NAND2_X1 U8485 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7108) );
  INV_X1 U8486 ( .A(n7108), .ZN(n6768) );
  AOI21_X1 U8487 ( .B1(n9854), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6768), .ZN(
        n6775) );
  NAND2_X1 U8488 ( .A1(n6769), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6771) );
  NAND2_X1 U8489 ( .A1(n6771), .A2(n6770), .ZN(n6773) );
  MUX2_X1 U8490 ( .A(n6787), .B(P2_REG1_REG_6__SCAN_IN), .S(n6786), .Z(n6772)
         );
  NAND2_X1 U8491 ( .A1(n6773), .A2(n6772), .ZN(n6785) );
  OAI211_X1 U8492 ( .C1(n6773), .C2(n6772), .A(n9853), .B(n6785), .ZN(n6774)
         );
  OAI211_X1 U8493 ( .C1(n9857), .C2(n6786), .A(n6775), .B(n6774), .ZN(n6776)
         );
  OR2_X1 U8494 ( .A1(n6777), .A2(n6776), .ZN(P2_U3251) );
  INV_X1 U8495 ( .A(n6786), .ZN(n6779) );
  AOI22_X1 U8496 ( .A1(n6783), .A2(n5846), .B1(P2_REG2_REG_7__SCAN_IN), .B2(
        n6803), .ZN(n6795) );
  AOI22_X1 U8497 ( .A1(n6904), .A2(n7096), .B1(P2_REG2_REG_8__SCAN_IN), .B2(
        n6910), .ZN(n6780) );
  NOR2_X1 U8498 ( .A1(n6781), .A2(n6780), .ZN(n6903) );
  AOI211_X1 U8499 ( .C1(n6781), .C2(n6780), .A(n6903), .B(n9549), .ZN(n6793)
         );
  INV_X1 U8500 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10051) );
  NOR2_X1 U8501 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10051), .ZN(n6782) );
  AOI21_X1 U8502 ( .B1(n9854), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6782), .ZN(
        n6791) );
  MUX2_X1 U8503 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6784), .S(n6783), .Z(n6799)
         );
  OAI21_X1 U8504 ( .B1(n6787), .B2(n6786), .A(n6785), .ZN(n6800) );
  NAND2_X1 U8505 ( .A1(n6799), .A2(n6800), .ZN(n6798) );
  OAI21_X1 U8506 ( .B1(n6803), .B2(n6784), .A(n6798), .ZN(n6789) );
  MUX2_X1 U8507 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9942), .S(n6904), .Z(n6788)
         );
  NAND2_X1 U8508 ( .A1(n6788), .A2(n6789), .ZN(n6909) );
  OAI211_X1 U8509 ( .C1(n6789), .C2(n6788), .A(n9853), .B(n6909), .ZN(n6790)
         );
  OAI211_X1 U8510 ( .C1(n9857), .C2(n6910), .A(n6791), .B(n6790), .ZN(n6792)
         );
  OR2_X1 U8511 ( .A1(n6793), .A2(n6792), .ZN(P2_U3253) );
  AOI211_X1 U8512 ( .C1(n6796), .C2(n6795), .A(n6794), .B(n9549), .ZN(n6805)
         );
  INV_X1 U8513 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6797) );
  NOR2_X1 U8514 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6797), .ZN(n7136) );
  AOI21_X1 U8515 ( .B1(n9854), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7136), .ZN(
        n6802) );
  OAI211_X1 U8516 ( .C1(n6800), .C2(n6799), .A(n9853), .B(n6798), .ZN(n6801)
         );
  OAI211_X1 U8517 ( .C1(n9857), .C2(n6803), .A(n6802), .B(n6801), .ZN(n6804)
         );
  OR2_X1 U8518 ( .A1(n6805), .A2(n6804), .ZN(P2_U3252) );
  NOR2_X1 U8519 ( .A1(n6815), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6807) );
  NOR2_X1 U8520 ( .A1(n6807), .A2(n6806), .ZN(n6810) );
  AOI22_X1 U8521 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6808), .B1(n6871), .B2(
        n5163), .ZN(n6809) );
  NOR2_X1 U8522 ( .A1(n6810), .A2(n6809), .ZN(n6864) );
  AOI21_X1 U8523 ( .B1(n6810), .B2(n6809), .A(n6864), .ZN(n6822) );
  INV_X1 U8524 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6813) );
  NOR2_X1 U8525 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6811), .ZN(n7307) );
  INV_X1 U8526 ( .A(n7307), .ZN(n6812) );
  OAI21_X1 U8527 ( .B1(n9769), .B2(n6813), .A(n6812), .ZN(n6820) );
  NAND2_X1 U8528 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n6871), .ZN(n6816) );
  OAI21_X1 U8529 ( .B1(n6871), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6816), .ZN(
        n6817) );
  AOI211_X1 U8530 ( .C1(n6818), .C2(n6817), .A(n6870), .B(n9723), .ZN(n6819)
         );
  AOI211_X1 U8531 ( .C1(n9753), .C2(n6871), .A(n6820), .B(n6819), .ZN(n6821)
         );
  OAI21_X1 U8532 ( .B1(n6822), .B2(n9765), .A(n6821), .ZN(P1_U3251) );
  INV_X1 U8533 ( .A(n6823), .ZN(n6881) );
  AOI22_X1 U8534 ( .A1(n8745), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n6824), .ZN(n6825) );
  OAI21_X1 U8535 ( .B1(n6881), .B2(n10256), .A(n6825), .ZN(P2_U3340) );
  NAND2_X1 U8536 ( .A1(n6826), .A2(n8497), .ZN(n6923) );
  INV_X1 U8537 ( .A(n6827), .ZN(n6828) );
  INV_X1 U8538 ( .A(n7049), .ZN(n6829) );
  NAND2_X1 U8539 ( .A1(n6830), .A2(n6829), .ZN(n6831) );
  NOR2_X1 U8540 ( .A1(n7048), .A2(n6831), .ZN(n6861) );
  AND2_X2 U8541 ( .A1(n6861), .A2(n7050), .ZN(n9935) );
  INV_X1 U8542 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6859) );
  NAND2_X1 U8543 ( .A1(n7114), .A2(n7121), .ZN(n6835) );
  NAND2_X1 U8544 ( .A1(n6832), .A2(n6833), .ZN(n6834) );
  NAND2_X1 U8545 ( .A1(n6835), .A2(n6834), .ZN(n7227) );
  NAND2_X1 U8546 ( .A1(n4953), .A2(n6836), .ZN(n8352) );
  NAND2_X1 U8547 ( .A1(n7227), .A2(n7231), .ZN(n6838) );
  NAND2_X1 U8548 ( .A1(n4953), .A2(n9885), .ZN(n6837) );
  NAND2_X1 U8549 ( .A1(n6838), .A2(n6837), .ZN(n7047) );
  NAND2_X1 U8550 ( .A1(n7144), .A2(n7071), .ZN(n8345) );
  NAND2_X1 U8551 ( .A1(n7047), .A2(n8314), .ZN(n6840) );
  NAND2_X1 U8552 ( .A1(n7144), .A2(n9891), .ZN(n6839) );
  NAND2_X1 U8553 ( .A1(n6840), .A2(n6839), .ZN(n7155) );
  INV_X1 U8554 ( .A(n6948), .ZN(n6841) );
  INV_X1 U8555 ( .A(n8662), .ZN(n7073) );
  NAND2_X1 U8556 ( .A1(n7073), .A2(n7152), .ZN(n6842) );
  INV_X1 U8557 ( .A(n8661), .ZN(n7268) );
  NAND2_X1 U8558 ( .A1(n7268), .A2(n8586), .ZN(n8347) );
  NAND2_X1 U8559 ( .A1(n8347), .A2(n8366), .ZN(n6850) );
  XOR2_X1 U8560 ( .A(n6941), .B(n6850), .Z(n7326) );
  AOI21_X1 U8561 ( .B1(n7053), .B2(n8340), .A(n8342), .ZN(n6845) );
  NAND2_X1 U8562 ( .A1(n6226), .A2(n6843), .ZN(n6844) );
  NAND2_X1 U8563 ( .A1(n6845), .A2(n6844), .ZN(n7797) );
  INV_X1 U8564 ( .A(n9922), .ZN(n9103) );
  NAND2_X1 U8565 ( .A1(n8310), .A2(n7247), .ZN(n8350) );
  NAND2_X1 U8566 ( .A1(n8350), .A2(n8360), .ZN(n7230) );
  INV_X1 U8567 ( .A(n7230), .ZN(n6847) );
  INV_X1 U8568 ( .A(n7231), .ZN(n6846) );
  NAND2_X1 U8569 ( .A1(n6847), .A2(n6846), .ZN(n7228) );
  NAND2_X1 U8570 ( .A1(n7228), .A2(n8352), .ZN(n7055) );
  NAND2_X1 U8571 ( .A1(n7055), .A2(n8356), .ZN(n6848) );
  NAND2_X1 U8572 ( .A1(n6848), .A2(n8345), .ZN(n7142) );
  INV_X1 U8573 ( .A(n7142), .ZN(n6849) );
  NAND2_X1 U8574 ( .A1(n6849), .A2(n8312), .ZN(n6949) );
  NAND2_X1 U8575 ( .A1(n6949), .A2(n6948), .ZN(n6851) );
  XNOR2_X1 U8576 ( .A(n6851), .B(n6850), .ZN(n6855) );
  AND2_X1 U8577 ( .A1(n6852), .A2(n8351), .ZN(n8307) );
  NOR2_X2 U8578 ( .A1(n8307), .A2(n8337), .ZN(n8970) );
  INV_X1 U8579 ( .A(n8993), .ZN(n8950) );
  OR2_X1 U8580 ( .A1(n6945), .A2(n8950), .ZN(n6854) );
  NAND2_X1 U8581 ( .A1(n8662), .A2(n8995), .ZN(n6853) );
  NAND2_X1 U8582 ( .A1(n6854), .A2(n6853), .ZN(n8584) );
  AOI21_X1 U8583 ( .B1(n6855), .B2(n8998), .A(n8584), .ZN(n7331) );
  NAND2_X1 U8584 ( .A1(n7236), .A2(n9891), .ZN(n7147) );
  INV_X1 U8585 ( .A(n7152), .ZN(n9897) );
  NAND2_X1 U8586 ( .A1(n6216), .A2(n6856), .ZN(n9927) );
  AOI211_X1 U8587 ( .C1(n8586), .C2(n7149), .A(n9927), .B(n7271), .ZN(n7329)
         );
  AOI21_X1 U8588 ( .B1(n9898), .B2(n8586), .A(n7329), .ZN(n6857) );
  OAI211_X1 U8589 ( .C1(n7326), .C2(n9874), .A(n7331), .B(n6857), .ZN(n6862)
         );
  NAND2_X1 U8590 ( .A1(n6862), .A2(n9935), .ZN(n6858) );
  OAI21_X1 U8591 ( .B1(n9935), .B2(n6859), .A(n6858), .ZN(P2_U3466) );
  AND2_X2 U8592 ( .A1(n6861), .A2(n6860), .ZN(n9947) );
  NAND2_X1 U8593 ( .A1(n6862), .A2(n9947), .ZN(n6863) );
  OAI21_X1 U8594 ( .B1(n9947), .B2(n6731), .A(n6863), .ZN(P2_U3525) );
  NOR2_X1 U8595 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6871), .ZN(n6865) );
  NOR2_X1 U8596 ( .A1(n6865), .A2(n6864), .ZN(n6868) );
  INV_X1 U8597 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6866) );
  AOI22_X1 U8598 ( .A1(n9248), .A2(n6866), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n6875), .ZN(n6867) );
  NOR2_X1 U8599 ( .A1(n6868), .A2(n6867), .ZN(n9250) );
  AOI21_X1 U8600 ( .B1(n6868), .B2(n6867), .A(n9250), .ZN(n6880) );
  NOR2_X1 U8601 ( .A1(n9248), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6869) );
  AOI21_X1 U8602 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9248), .A(n6869), .ZN(
        n6873) );
  OAI21_X1 U8603 ( .B1(n6873), .B2(n6872), .A(n9237), .ZN(n6878) );
  AND2_X1 U8604 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7393) );
  AOI21_X1 U8605 ( .B1(n9655), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n7393), .ZN(
        n6874) );
  OAI21_X1 U8606 ( .B1(n6876), .B2(n6875), .A(n6874), .ZN(n6877) );
  AOI21_X1 U8607 ( .B1(n6878), .B2(n9758), .A(n6877), .ZN(n6879) );
  OAI21_X1 U8608 ( .B1(n6880), .B2(n9765), .A(n6879), .ZN(P1_U3252) );
  INV_X1 U8609 ( .A(n9752), .ZN(n9263) );
  OAI222_X1 U8610 ( .A1(n7924), .A2(n10004), .B1(n7920), .B2(n6881), .C1(
        P1_U3084), .C2(n9263), .ZN(P1_U3335) );
  OR2_X1 U8611 ( .A1(n6885), .A2(n6884), .ZN(n6887) );
  NAND2_X1 U8612 ( .A1(n6887), .A2(n6886), .ZN(n7332) );
  OAI21_X1 U8613 ( .B1(n8096), .B2(n6889), .A(n6888), .ZN(n6896) );
  INV_X1 U8614 ( .A(n9235), .ZN(n7007) );
  OAI22_X1 U8615 ( .A1(n7007), .A2(n5559), .B1(n6268), .B2(n9577), .ZN(n6895)
         );
  OR2_X1 U8616 ( .A1(n6891), .A2(n6890), .ZN(n6893) );
  OR2_X1 U8617 ( .A1(n7128), .A2(n8125), .ZN(n6892) );
  AND2_X1 U8618 ( .A1(n6893), .A2(n6892), .ZN(n9582) );
  NOR2_X1 U8619 ( .A1(n7332), .A2(n9582), .ZN(n6894) );
  AOI211_X1 U8620 ( .C1(n9586), .C2(n6896), .A(n6895), .B(n6894), .ZN(n7336)
         );
  INV_X1 U8621 ( .A(n7205), .ZN(n6897) );
  AOI211_X1 U8622 ( .C1(n7130), .C2(n6259), .A(n9832), .B(n6897), .ZN(n7334)
         );
  AOI21_X1 U8623 ( .B1(n6259), .B2(n9500), .A(n7334), .ZN(n6898) );
  OAI211_X1 U8624 ( .C1(n7016), .C2(n7332), .A(n7336), .B(n6898), .ZN(n6900)
         );
  NAND2_X1 U8625 ( .A1(n6900), .A2(n9852), .ZN(n6899) );
  OAI21_X1 U8626 ( .B1(n9852), .B2(n6531), .A(n6899), .ZN(P1_U3524) );
  INV_X1 U8627 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6902) );
  NAND2_X1 U8628 ( .A1(n6900), .A2(n9840), .ZN(n6901) );
  OAI21_X1 U8629 ( .B1(n9840), .B2(n6902), .A(n6901), .ZN(P1_U3457) );
  NAND2_X1 U8630 ( .A1(n6984), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6905) );
  OAI21_X1 U8631 ( .B1(n6984), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6905), .ZN(
        n6906) );
  AOI211_X1 U8632 ( .C1(n6907), .C2(n6906), .A(n6983), .B(n9549), .ZN(n6916)
         );
  NAND2_X1 U8633 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7479) );
  INV_X1 U8634 ( .A(n7479), .ZN(n6908) );
  AOI21_X1 U8635 ( .B1(n9854), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n6908), .ZN(
        n6914) );
  INV_X1 U8636 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9942) );
  OAI21_X1 U8637 ( .B1(n6910), .B2(n9942), .A(n6909), .ZN(n6912) );
  MUX2_X1 U8638 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6990), .S(n6984), .Z(n6911)
         );
  NAND2_X1 U8639 ( .A1(n6911), .A2(n6912), .ZN(n6989) );
  OAI211_X1 U8640 ( .C1(n6912), .C2(n6911), .A(n9853), .B(n6989), .ZN(n6913)
         );
  OAI211_X1 U8641 ( .C1(n9857), .C2(n6991), .A(n6914), .B(n6913), .ZN(n6915)
         );
  OR2_X1 U8642 ( .A1(n6916), .A2(n6915), .ZN(P2_U3254) );
  INV_X1 U8643 ( .A(n6917), .ZN(n7925) );
  OAI222_X1 U8644 ( .A1(n7924), .A2(n10050), .B1(n7920), .B2(n7925), .C1(n9778), .C2(P1_U3084), .ZN(P1_U3334) );
  AOI21_X1 U8645 ( .B1(n6919), .B2(n6918), .A(n8643), .ZN(n6921) );
  NAND2_X1 U8646 ( .A1(n6921), .A2(n6920), .ZN(n6928) );
  AOI22_X1 U8647 ( .A1(n8993), .A2(n8663), .B1(n6922), .B2(n8995), .ZN(n7232)
         );
  INV_X1 U8648 ( .A(n7232), .ZN(n6926) );
  INV_X1 U8649 ( .A(n6923), .ZN(n6924) );
  NAND2_X1 U8650 ( .A1(n6925), .A2(n6924), .ZN(n8549) );
  AOI22_X1 U8651 ( .A1(n6926), .A2(n8638), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n8549), .ZN(n6927) );
  OAI211_X1 U8652 ( .C1(n9885), .C2(n8619), .A(n6928), .B(n6927), .ZN(P2_U3239) );
  INV_X1 U8653 ( .A(n6929), .ZN(n6931) );
  NOR2_X1 U8654 ( .A1(n6931), .A2(n6930), .ZN(n6932) );
  XNOR2_X1 U8655 ( .A(n6933), .B(n6932), .ZN(n6940) );
  INV_X1 U8656 ( .A(n7150), .ZN(n6938) );
  NAND2_X1 U8657 ( .A1(n8629), .A2(n9897), .ZN(n6935) );
  NAND2_X1 U8658 ( .A1(n6935), .A2(n6934), .ZN(n6937) );
  OAI22_X1 U8659 ( .A1(n7144), .A2(n8614), .B1(n8613), .B2(n7268), .ZN(n6936)
         );
  AOI211_X1 U8660 ( .C1(n6938), .C2(n8627), .A(n6937), .B(n6936), .ZN(n6939)
         );
  OAI21_X1 U8661 ( .B1(n6940), .B2(n8643), .A(n6939), .ZN(P2_U3232) );
  INV_X1 U8662 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6956) );
  NAND2_X1 U8663 ( .A1(n8661), .A2(n8586), .ZN(n6942) );
  NAND2_X1 U8664 ( .A1(n6943), .A2(n6942), .ZN(n7263) );
  NAND2_X1 U8665 ( .A1(n6945), .A2(n7273), .ZN(n8374) );
  INV_X2 U8666 ( .A(n7273), .ZN(n6944) );
  NAND2_X1 U8667 ( .A1(n8660), .A2(n6944), .ZN(n8373) );
  AND2_X1 U8668 ( .A1(n8374), .A2(n8373), .ZN(n8317) );
  NAND2_X1 U8669 ( .A1(n7263), .A2(n7265), .ZN(n6947) );
  OR2_X1 U8670 ( .A1(n6945), .A2(n6944), .ZN(n6946) );
  NOR2_X1 U8671 ( .A1(n8659), .A2(n7316), .ZN(n8380) );
  NAND2_X1 U8672 ( .A1(n8659), .A2(n7316), .ZN(n8379) );
  XNOR2_X1 U8673 ( .A(n7085), .B(n7086), .ZN(n7322) );
  NAND2_X1 U8674 ( .A1(n6949), .A2(n8313), .ZN(n7264) );
  AND2_X1 U8675 ( .A1(n8347), .A2(n8374), .ZN(n6950) );
  XNOR2_X1 U8676 ( .A(n4459), .B(n8376), .ZN(n6951) );
  INV_X1 U8677 ( .A(n7482), .ZN(n8658) );
  AOI222_X1 U8678 ( .A1(n8998), .A2(n6951), .B1(n8658), .B2(n8993), .C1(n8660), 
        .C2(n8995), .ZN(n7317) );
  INV_X1 U8679 ( .A(n7316), .ZN(n7137) );
  AND2_X1 U8680 ( .A1(n7271), .A2(n6944), .ZN(n6952) );
  INV_X1 U8681 ( .A(n6952), .ZN(n7270) );
  INV_X1 U8682 ( .A(n7097), .ZN(n6953) );
  AOI21_X1 U8683 ( .B1(n7137), .B2(n7270), .A(n6953), .ZN(n7320) );
  AOI22_X1 U8684 ( .A1(n7320), .A2(n9899), .B1(n9898), .B2(n7137), .ZN(n6954)
         );
  OAI211_X1 U8685 ( .C1(n9874), .C2(n7322), .A(n7317), .B(n6954), .ZN(n6957)
         );
  NAND2_X1 U8686 ( .A1(n6957), .A2(n9935), .ZN(n6955) );
  OAI21_X1 U8687 ( .B1(n9935), .B2(n6956), .A(n6955), .ZN(P2_U3472) );
  NAND2_X1 U8688 ( .A1(n6957), .A2(n9947), .ZN(n6958) );
  OAI21_X1 U8689 ( .B1(n9947), .B2(n6784), .A(n6958), .ZN(P2_U3527) );
  NAND2_X1 U8690 ( .A1(n6960), .A2(n6961), .ZN(n6962) );
  XOR2_X1 U8691 ( .A(n6959), .B(n6962), .Z(n6969) );
  INV_X1 U8692 ( .A(n7185), .ZN(n6967) );
  NAND2_X1 U8693 ( .A1(n7192), .A2(n9500), .ZN(n9806) );
  NOR2_X1 U8694 ( .A1(n9165), .A2(n9806), .ZN(n6966) );
  NAND2_X1 U8695 ( .A1(n9183), .A2(n9231), .ZN(n6964) );
  OAI211_X1 U8696 ( .C1(n7201), .C2(n9207), .A(n6964), .B(n6963), .ZN(n6965)
         );
  AOI211_X1 U8697 ( .C1(n6967), .C2(n9211), .A(n6966), .B(n6965), .ZN(n6968)
         );
  OAI21_X1 U8698 ( .B1(n6969), .B2(n9201), .A(n6968), .ZN(P1_U3228) );
  INV_X1 U8699 ( .A(n6970), .ZN(n8277) );
  OAI222_X1 U8700 ( .A1(P1_U3084), .A2(n5651), .B1(n7920), .B2(n8277), .C1(
        n6971), .C2(n9531), .ZN(P1_U3333) );
  XOR2_X1 U8701 ( .A(n6973), .B(n6972), .Z(n6980) );
  INV_X1 U8702 ( .A(n9207), .ZN(n9194) );
  NAND2_X1 U8703 ( .A1(n6974), .A2(n9194), .ZN(n6976) );
  OAI211_X1 U8704 ( .C1(n7258), .C2(n9208), .A(n6976), .B(n6975), .ZN(n6978)
         );
  NOR2_X1 U8705 ( .A1(n9186), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6977) );
  AOI211_X1 U8706 ( .C1(n9188), .C2(n7223), .A(n6978), .B(n6977), .ZN(n6979)
         );
  OAI21_X1 U8707 ( .B1(n6980), .B2(n9201), .A(n6979), .ZN(P1_U3216) );
  INV_X1 U8708 ( .A(n6981), .ZN(n6999) );
  OAI222_X1 U8709 ( .A1(n8511), .A2(n6982), .B1(n7928), .B2(n6999), .C1(n8338), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  NAND2_X1 U8710 ( .A1(n7451), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6985) );
  OAI21_X1 U8711 ( .B1(n7451), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6985), .ZN(
        n6986) );
  AOI211_X1 U8712 ( .C1(n6987), .C2(n6986), .A(n7450), .B(n9549), .ZN(n6998)
         );
  NOR2_X1 U8713 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10187), .ZN(n6988) );
  AOI21_X1 U8714 ( .B1(n9854), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n6988), .ZN(
        n6996) );
  INV_X1 U8715 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6990) );
  OAI21_X1 U8716 ( .B1(n6991), .B2(n6990), .A(n6989), .ZN(n6994) );
  MUX2_X1 U8717 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6992), .S(n7451), .Z(n6993)
         );
  NAND2_X1 U8718 ( .A1(n6993), .A2(n6994), .ZN(n7458) );
  OAI211_X1 U8719 ( .C1(n6994), .C2(n6993), .A(n9853), .B(n7458), .ZN(n6995)
         );
  OAI211_X1 U8720 ( .C1(n9857), .C2(n7459), .A(n6996), .B(n6995), .ZN(n6997)
         );
  OR2_X1 U8721 ( .A1(n6998), .A2(n6997), .ZN(P2_U3255) );
  OAI222_X1 U8722 ( .A1(n9531), .A2(n7000), .B1(P1_U3084), .B2(n8125), .C1(
        n7920), .C2(n6999), .ZN(P1_U3332) );
  AOI21_X1 U8723 ( .B1(n7002), .B2(n7001), .A(n9188), .ZN(n7082) );
  INV_X1 U8724 ( .A(n7082), .ZN(n7015) );
  OAI21_X1 U8725 ( .B1(n7005), .B2(n7003), .A(n7004), .ZN(n7006) );
  NAND2_X1 U8726 ( .A1(n7006), .A2(n9204), .ZN(n7010) );
  OAI22_X1 U8727 ( .A1(n7007), .A2(n9207), .B1(n6268), .B2(n9208), .ZN(n7008)
         );
  AOI21_X1 U8728 ( .B1(n9188), .B2(n6259), .A(n7008), .ZN(n7009) );
  OAI211_X1 U8729 ( .C1(n7015), .C2(n7011), .A(n7010), .B(n7009), .ZN(P1_U3220) );
  AOI22_X1 U8730 ( .A1(n9188), .A2(n7130), .B1(n9183), .B2(n6258), .ZN(n7014)
         );
  NAND2_X1 U8731 ( .A1(n7012), .A2(n9204), .ZN(n7013) );
  OAI211_X1 U8732 ( .C1(n7015), .C2(n7126), .A(n7014), .B(n7013), .ZN(P1_U3230) );
  NAND2_X1 U8733 ( .A1(n7017), .A2(n7020), .ZN(n7018) );
  NAND2_X1 U8734 ( .A1(n7019), .A2(n7018), .ZN(n9782) );
  XNOR2_X1 U8735 ( .A(n7021), .B(n5620), .ZN(n7024) );
  OAI22_X1 U8736 ( .A1(n7022), .A2(n9577), .B1(n7258), .B2(n5559), .ZN(n7023)
         );
  AOI21_X1 U8737 ( .B1(n7024), .B2(n9586), .A(n7023), .ZN(n9781) );
  NAND2_X1 U8738 ( .A1(n7186), .A2(n9773), .ZN(n7025) );
  INV_X1 U8739 ( .A(n9832), .ZN(n9595) );
  NAND2_X1 U8740 ( .A1(n7025), .A2(n9595), .ZN(n7026) );
  NOR2_X1 U8741 ( .A1(n7435), .A2(n7026), .ZN(n9779) );
  AOI21_X1 U8742 ( .B1(n9773), .B2(n9500), .A(n9779), .ZN(n7027) );
  OAI211_X1 U8743 ( .C1(n9505), .C2(n9782), .A(n9781), .B(n7027), .ZN(n7029)
         );
  NAND2_X1 U8744 ( .A1(n7029), .A2(n9852), .ZN(n7028) );
  OAI21_X1 U8745 ( .B1(n9852), .B2(n6529), .A(n7028), .ZN(P1_U3528) );
  NAND2_X1 U8746 ( .A1(n7029), .A2(n9840), .ZN(n7030) );
  OAI21_X1 U8747 ( .B1(n9840), .B2(n5078), .A(n7030), .ZN(P1_U3469) );
  NAND2_X1 U8748 ( .A1(n7031), .A2(n7032), .ZN(n7036) );
  NAND2_X1 U8749 ( .A1(n7034), .A2(n7033), .ZN(n7035) );
  XNOR2_X1 U8750 ( .A(n7036), .B(n7035), .ZN(n7045) );
  AOI21_X1 U8751 ( .B1(n9230), .B2(n9194), .A(n7037), .ZN(n7043) );
  NAND2_X1 U8752 ( .A1(n9188), .A2(n7038), .ZN(n7042) );
  INV_X1 U8753 ( .A(n7387), .ZN(n7039) );
  NAND2_X1 U8754 ( .A1(n9211), .A2(n7039), .ZN(n7041) );
  NAND2_X1 U8755 ( .A1(n9228), .A2(n9183), .ZN(n7040) );
  NAND4_X1 U8756 ( .A1(n7043), .A2(n7042), .A3(n7041), .A4(n7040), .ZN(n7044)
         );
  AOI21_X1 U8757 ( .B1(n7045), .B2(n9204), .A(n7044), .ZN(n7046) );
  INV_X1 U8758 ( .A(n7046), .ZN(P1_U3211) );
  XNOR2_X1 U8759 ( .A(n7047), .B(n8356), .ZN(n9890) );
  INV_X1 U8760 ( .A(n7048), .ZN(n7052) );
  AND2_X1 U8761 ( .A1(n7050), .A2(n7049), .ZN(n7051) );
  NAND2_X1 U8762 ( .A1(n7052), .A2(n7051), .ZN(n7062) );
  NAND2_X2 U8763 ( .A1(n7062), .A2(n8934), .ZN(n8936) );
  NOR2_X1 U8764 ( .A1(n7053), .A2(n8756), .ZN(n7054) );
  NAND2_X1 U8765 ( .A1(n8936), .A2(n7054), .ZN(n7807) );
  XNOR2_X1 U8766 ( .A(n7055), .B(n8356), .ZN(n7057) );
  INV_X1 U8767 ( .A(n8995), .ZN(n8952) );
  OAI22_X1 U8768 ( .A1(n7073), .A2(n8950), .B1(n4953), .B2(n8952), .ZN(n7056)
         );
  AOI21_X1 U8769 ( .B1(n7057), .B2(n8998), .A(n7056), .ZN(n7058) );
  OAI21_X1 U8770 ( .B1(n9890), .B2(n7797), .A(n7058), .ZN(n9893) );
  NAND2_X1 U8771 ( .A1(n9893), .A2(n8936), .ZN(n7067) );
  OAI22_X1 U8772 ( .A1(n8936), .A2(n7060), .B1(n8934), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n7065) );
  OR2_X1 U8773 ( .A1(n7236), .A2(n9891), .ZN(n7061) );
  NAND2_X1 U8774 ( .A1(n7147), .A2(n7061), .ZN(n9892) );
  INV_X1 U8775 ( .A(n7062), .ZN(n7063) );
  NAND2_X1 U8776 ( .A1(n7063), .A2(n8504), .ZN(n8801) );
  NOR2_X1 U8777 ( .A1(n9892), .A2(n8801), .ZN(n7064) );
  AOI211_X1 U8778 ( .C1(n8845), .C2(n7071), .A(n7065), .B(n7064), .ZN(n7066)
         );
  OAI211_X1 U8779 ( .C1(n9890), .C2(n7807), .A(n7067), .B(n7066), .ZN(P2_U3293) );
  INV_X1 U8780 ( .A(n8643), .ZN(n8622) );
  OAI211_X1 U8781 ( .C1(n7070), .C2(n7069), .A(n7068), .B(n8622), .ZN(n7077)
         );
  NAND2_X1 U8782 ( .A1(n8629), .A2(n7071), .ZN(n7072) );
  OAI21_X1 U8783 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n5785), .A(n7072), .ZN(n7075) );
  OAI22_X1 U8784 ( .A1(n4953), .A2(n8614), .B1(n8613), .B2(n7073), .ZN(n7074)
         );
  AOI211_X1 U8785 ( .C1(n8627), .C2(n5785), .A(n7075), .B(n7074), .ZN(n7076)
         );
  NAND2_X1 U8786 ( .A1(n7077), .A2(n7076), .ZN(P2_U3220) );
  XOR2_X1 U8787 ( .A(n7079), .B(n7078), .Z(n7084) );
  INV_X1 U8788 ( .A(n9199), .ZN(n9214) );
  AOI22_X1 U8789 ( .A1(n9233), .A2(n9183), .B1(n9194), .B2(n6258), .ZN(n7080)
         );
  OAI21_X1 U8790 ( .B1(n9214), .B2(n9796), .A(n7080), .ZN(n7081) );
  AOI21_X1 U8791 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n7082), .A(n7081), .ZN(
        n7083) );
  OAI21_X1 U8792 ( .B1(n7084), .B2(n9201), .A(n7083), .ZN(P1_U3235) );
  INV_X1 U8793 ( .A(n8659), .ZN(n7269) );
  NAND2_X1 U8794 ( .A1(n7482), .A2(n8540), .ZN(n8383) );
  NAND2_X1 U8795 ( .A1(n8658), .A2(n9911), .ZN(n8384) );
  OAI21_X1 U8796 ( .B1(n7087), .B2(n8381), .A(n7280), .ZN(n9910) );
  INV_X1 U8797 ( .A(n8380), .ZN(n7089) );
  OAI21_X1 U8798 ( .B1(n7091), .B2(n7090), .A(n7285), .ZN(n7094) );
  OR2_X1 U8799 ( .A1(n7286), .A2(n8950), .ZN(n7093) );
  NAND2_X1 U8800 ( .A1(n8659), .A2(n8995), .ZN(n7092) );
  NAND2_X1 U8801 ( .A1(n7093), .A2(n7092), .ZN(n8537) );
  AOI21_X1 U8802 ( .B1(n7094), .B2(n8998), .A(n8537), .ZN(n7095) );
  OAI21_X1 U8803 ( .B1(n9910), .B2(n7797), .A(n7095), .ZN(n9913) );
  NAND2_X1 U8804 ( .A1(n9913), .A2(n8936), .ZN(n7102) );
  OAI22_X1 U8805 ( .A1(n8936), .A2(n7096), .B1(n8538), .B2(n8934), .ZN(n7100)
         );
  NAND2_X1 U8806 ( .A1(n7097), .A2(n8540), .ZN(n7098) );
  NAND2_X1 U8807 ( .A1(n7360), .A2(n7098), .ZN(n9912) );
  NOR2_X1 U8808 ( .A1(n9912), .A2(n8801), .ZN(n7099) );
  AOI211_X1 U8809 ( .C1(n8845), .C2(n8540), .A(n7100), .B(n7099), .ZN(n7101)
         );
  OAI211_X1 U8810 ( .C1(n9910), .C2(n7807), .A(n7102), .B(n7101), .ZN(P2_U3288) );
  INV_X1 U8811 ( .A(n7103), .ZN(n7104) );
  AOI21_X1 U8812 ( .B1(n7106), .B2(n7105), .A(n7104), .ZN(n7113) );
  INV_X1 U8813 ( .A(n7107), .ZN(n7272) );
  NAND2_X1 U8814 ( .A1(n8629), .A2(n7273), .ZN(n7109) );
  NAND2_X1 U8815 ( .A1(n7109), .A2(n7108), .ZN(n7111) );
  OAI22_X1 U8816 ( .A1(n7268), .A2(n8614), .B1(n8613), .B2(n7269), .ZN(n7110)
         );
  AOI211_X1 U8817 ( .C1(n7272), .C2(n8627), .A(n7111), .B(n7110), .ZN(n7112)
         );
  OAI21_X1 U8818 ( .B1(n7113), .B2(n8643), .A(n7112), .ZN(P2_U3241) );
  XNOR2_X1 U8819 ( .A(n7114), .B(n7247), .ZN(n7116) );
  INV_X1 U8820 ( .A(n7115), .ZN(n8666) );
  AOI222_X1 U8821 ( .A1(n8998), .A2(n7116), .B1(n8664), .B2(n8993), .C1(n8666), 
        .C2(n8995), .ZN(n9879) );
  OAI21_X1 U8822 ( .B1(n6833), .B2(n9872), .A(n7234), .ZN(n9878) );
  NOR2_X1 U8823 ( .A1(n8801), .A2(n9878), .ZN(n7120) );
  OAI22_X1 U8824 ( .A1(n8936), .A2(n7118), .B1(n7117), .B2(n8934), .ZN(n7119)
         );
  AOI211_X1 U8825 ( .C1(n8845), .C2(n8550), .A(n7120), .B(n7119), .ZN(n7124)
         );
  XNOR2_X1 U8826 ( .A(n7121), .B(n7114), .ZN(n9882) );
  INV_X1 U8827 ( .A(n7797), .ZN(n7497) );
  NAND2_X1 U8828 ( .A1(n8936), .A2(n7497), .ZN(n7122) );
  NAND2_X1 U8829 ( .A1(n7807), .A2(n7122), .ZN(n8905) );
  NAND2_X1 U8830 ( .A1(n9882), .A2(n8905), .ZN(n7123) );
  OAI211_X1 U8831 ( .C1(n9879), .C2(n8956), .A(n7124), .B(n7123), .ZN(P2_U3295) );
  OAI21_X1 U8832 ( .B1(n7126), .B2(n9776), .A(n7125), .ZN(n7127) );
  NAND2_X1 U8833 ( .A1(n7127), .A2(n9785), .ZN(n7132) );
  NOR2_X1 U8834 ( .A1(n7128), .A2(n5652), .ZN(n7129) );
  AND2_X1 U8835 ( .A1(n9785), .A2(n7129), .ZN(n9401) );
  OAI21_X1 U8836 ( .B1(n9590), .B2(n9401), .A(n7130), .ZN(n7131) );
  OAI211_X1 U8837 ( .C1(n4995), .C2(n9785), .A(n7132), .B(n7131), .ZN(P1_U3291) );
  XNOR2_X1 U8838 ( .A(n7134), .B(n7133), .ZN(n7140) );
  AOI22_X1 U8839 ( .A1(n8628), .A2(n8660), .B1(n8624), .B2(n8658), .ZN(n7139)
         );
  NOR2_X1 U8840 ( .A1(n8640), .A2(n7313), .ZN(n7135) );
  AOI211_X1 U8841 ( .C1(n7137), .C2(n8629), .A(n7136), .B(n7135), .ZN(n7138)
         );
  OAI211_X1 U8842 ( .C1(n7140), .C2(n8643), .A(n7139), .B(n7138), .ZN(P2_U3215) );
  INV_X1 U8843 ( .A(n7156), .ZN(n7141) );
  XNOR2_X1 U8844 ( .A(n7142), .B(n7141), .ZN(n7146) );
  NAND2_X1 U8845 ( .A1(n8661), .A2(n8993), .ZN(n7143) );
  OAI21_X1 U8846 ( .B1(n7144), .B2(n8952), .A(n7143), .ZN(n7145) );
  AOI21_X1 U8847 ( .B1(n7146), .B2(n8998), .A(n7145), .ZN(n9904) );
  NAND2_X1 U8848 ( .A1(n7147), .A2(n9897), .ZN(n7148) );
  AND2_X1 U8849 ( .A1(n7149), .A2(n7148), .ZN(n9900) );
  OAI22_X1 U8850 ( .A1(n8936), .A2(n7151), .B1(n7150), .B2(n8934), .ZN(n7154)
         );
  NOR2_X1 U8851 ( .A1(n8989), .A2(n7152), .ZN(n7153) );
  AOI211_X1 U8852 ( .C1(n9900), .C2(n9001), .A(n7154), .B(n7153), .ZN(n7158)
         );
  XNOR2_X1 U8853 ( .A(n7155), .B(n7156), .ZN(n9901) );
  NAND2_X1 U8854 ( .A1(n9901), .A2(n8905), .ZN(n7157) );
  OAI211_X1 U8855 ( .C1(n9904), .C2(n8956), .A(n7158), .B(n7157), .ZN(P2_U3292) );
  INV_X1 U8856 ( .A(n7159), .ZN(n7168) );
  AND2_X1 U8857 ( .A1(n7161), .A2(n7160), .ZN(n7167) );
  INV_X1 U8858 ( .A(n7162), .ZN(n7164) );
  NAND2_X1 U8859 ( .A1(n7164), .A2(n7163), .ZN(n7166) );
  AOI22_X1 U8860 ( .A1(n7168), .A2(n7167), .B1(n7166), .B2(n7165), .ZN(n7176)
         );
  NOR2_X1 U8861 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7169), .ZN(n9657) );
  AOI21_X1 U8862 ( .B1(n9229), .B2(n9194), .A(n9657), .ZN(n7174) );
  NAND2_X1 U8863 ( .A1(n9188), .A2(n7410), .ZN(n7173) );
  INV_X1 U8864 ( .A(n7408), .ZN(n7170) );
  NAND2_X1 U8865 ( .A1(n9211), .A2(n7170), .ZN(n7172) );
  NAND2_X1 U8866 ( .A1(n9183), .A2(n9227), .ZN(n7171) );
  AND4_X1 U8867 ( .A1(n7174), .A2(n7173), .A3(n7172), .A4(n7171), .ZN(n7175)
         );
  OAI21_X1 U8868 ( .B1(n7176), .B2(n9201), .A(n7175), .ZN(P1_U3219) );
  OAI21_X1 U8869 ( .B1(n7178), .B2(n7180), .A(n7177), .ZN(n9810) );
  INV_X1 U8870 ( .A(n9810), .ZN(n7195) );
  INV_X1 U8871 ( .A(n7180), .ZN(n8093) );
  XNOR2_X1 U8872 ( .A(n7179), .B(n8093), .ZN(n7184) );
  INV_X1 U8873 ( .A(n9582), .ZN(n7511) );
  OAI22_X1 U8874 ( .A1(n7181), .A2(n9577), .B1(n7201), .B2(n5559), .ZN(n7182)
         );
  AOI21_X1 U8875 ( .B1(n9810), .B2(n7511), .A(n7182), .ZN(n7183) );
  OAI21_X1 U8876 ( .B1(n5556), .B2(n7184), .A(n7183), .ZN(n9808) );
  NAND2_X1 U8877 ( .A1(n9808), .A2(n9785), .ZN(n7194) );
  OAI22_X1 U8878 ( .A1(n9785), .A2(n6517), .B1(n7185), .B2(n9776), .ZN(n7191)
         );
  INV_X1 U8879 ( .A(n7220), .ZN(n7188) );
  OAI211_X1 U8880 ( .C1(n7188), .C2(n7187), .A(n9595), .B(n7186), .ZN(n9807)
         );
  NOR2_X1 U8881 ( .A1(n7189), .A2(n9349), .ZN(n9598) );
  INV_X1 U8882 ( .A(n9598), .ZN(n9329) );
  NOR2_X1 U8883 ( .A1(n9807), .A2(n9329), .ZN(n7190) );
  AOI211_X1 U8884 ( .C1(n9590), .C2(n7192), .A(n7191), .B(n7190), .ZN(n7193)
         );
  OAI211_X1 U8885 ( .C1(n7195), .C2(n9425), .A(n7194), .B(n7193), .ZN(P1_U3287) );
  INV_X1 U8886 ( .A(n7196), .ZN(n7197) );
  AOI21_X1 U8887 ( .B1(n8092), .B2(n7198), .A(n7197), .ZN(n9795) );
  OAI21_X1 U8888 ( .B1(n8092), .B2(n7199), .A(n7200), .ZN(n7203) );
  OAI22_X1 U8889 ( .A1(n8212), .A2(n5559), .B1(n7201), .B2(n9577), .ZN(n7202)
         );
  AOI21_X1 U8890 ( .B1(n7203), .B2(n9586), .A(n7202), .ZN(n7204) );
  OAI21_X1 U8891 ( .B1(n9795), .B2(n9582), .A(n7204), .ZN(n9798) );
  NAND2_X1 U8892 ( .A1(n9798), .A2(n9785), .ZN(n7211) );
  OAI22_X1 U8893 ( .A1(n9785), .A2(n6512), .B1(n4631), .B2(n9776), .ZN(n7208)
         );
  AND2_X1 U8894 ( .A1(n7209), .A2(n7205), .ZN(n7206) );
  OR2_X1 U8895 ( .A1(n7206), .A2(n7218), .ZN(n9797) );
  INV_X1 U8896 ( .A(n9401), .ZN(n9281) );
  NOR2_X1 U8897 ( .A1(n9797), .A2(n9281), .ZN(n7207) );
  AOI211_X1 U8898 ( .C1(n9590), .C2(n7209), .A(n7208), .B(n7207), .ZN(n7210)
         );
  OAI211_X1 U8899 ( .C1(n9795), .C2(n9425), .A(n7211), .B(n7210), .ZN(P1_U3289) );
  OAI21_X1 U8900 ( .B1(n7213), .B2(n8090), .A(n7212), .ZN(n9805) );
  INV_X1 U8901 ( .A(n9805), .ZN(n7226) );
  XNOR2_X1 U8902 ( .A(n8148), .B(n8090), .ZN(n7216) );
  OAI22_X1 U8903 ( .A1(n7258), .A2(n9577), .B1(n6268), .B2(n5559), .ZN(n7214)
         );
  AOI21_X1 U8904 ( .B1(n9805), .B2(n7511), .A(n7214), .ZN(n7215) );
  OAI21_X1 U8905 ( .B1(n5556), .B2(n7216), .A(n7215), .ZN(n9803) );
  NAND2_X1 U8906 ( .A1(n9803), .A2(n9785), .ZN(n7225) );
  OAI22_X1 U8907 ( .A1(n9785), .A2(n7217), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9776), .ZN(n7222) );
  OR2_X1 U8908 ( .A1(n7218), .A2(n9801), .ZN(n7219) );
  NAND2_X1 U8909 ( .A1(n7220), .A2(n7219), .ZN(n9802) );
  NOR2_X1 U8910 ( .A1(n9802), .A2(n9281), .ZN(n7221) );
  AOI211_X1 U8911 ( .C1(n9590), .C2(n7223), .A(n7222), .B(n7221), .ZN(n7224)
         );
  OAI211_X1 U8912 ( .C1(n7226), .C2(n9425), .A(n7225), .B(n7224), .ZN(P1_U3288) );
  XNOR2_X1 U8913 ( .A(n7231), .B(n7227), .ZN(n9888) );
  INV_X1 U8914 ( .A(n9888), .ZN(n7244) );
  INV_X1 U8915 ( .A(n7228), .ZN(n7229) );
  AOI21_X1 U8916 ( .B1(n7231), .B2(n7230), .A(n7229), .ZN(n7233) );
  OAI21_X1 U8917 ( .B1(n7233), .B2(n8970), .A(n7232), .ZN(n9886) );
  NAND2_X1 U8918 ( .A1(n7234), .A2(n7239), .ZN(n7235) );
  NAND2_X1 U8919 ( .A1(n7235), .A2(n9899), .ZN(n7237) );
  OR2_X1 U8920 ( .A1(n7237), .A2(n7236), .ZN(n9884) );
  OAI22_X1 U8921 ( .A1(n8801), .A2(n9884), .B1(n5754), .B2(n8934), .ZN(n7238)
         );
  INV_X1 U8922 ( .A(n7238), .ZN(n7241) );
  NAND2_X1 U8923 ( .A1(n8845), .A2(n7239), .ZN(n7240) );
  OAI211_X1 U8924 ( .C1(n5752), .C2(n8936), .A(n7241), .B(n7240), .ZN(n7242)
         );
  AOI21_X1 U8925 ( .B1(n9886), .B2(n8936), .A(n7242), .ZN(n7243) );
  OAI21_X1 U8926 ( .B1(n9003), .B2(n7244), .A(n7243), .ZN(P2_U3294) );
  INV_X1 U8927 ( .A(n7245), .ZN(n7922) );
  OAI222_X1 U8928 ( .A1(n8511), .A2(n7246), .B1(n7928), .B2(n7922), .C1(
        P2_U3152), .C2(n8340), .ZN(P2_U3336) );
  NAND2_X1 U8929 ( .A1(n8666), .A2(n9872), .ZN(n8359) );
  AND2_X1 U8930 ( .A1(n7247), .A2(n8359), .ZN(n9875) );
  OAI22_X1 U8931 ( .A1(n9875), .A2(n8970), .B1(n6832), .B2(n8950), .ZN(n9877)
         );
  OAI22_X1 U8932 ( .A1(n8936), .A2(n9855), .B1(n7248), .B2(n8934), .ZN(n7250)
         );
  AOI21_X1 U8933 ( .B1(n8989), .B2(n8801), .A(n9872), .ZN(n7249) );
  AOI211_X1 U8934 ( .C1(n8936), .C2(n9877), .A(n7250), .B(n7249), .ZN(n7251)
         );
  OAI21_X1 U8935 ( .B1(n9875), .B2(n9003), .A(n7251), .ZN(P2_U3296) );
  NAND2_X1 U8936 ( .A1(n6960), .A2(n7252), .ZN(n7254) );
  AND2_X1 U8937 ( .A1(n7254), .A2(n7253), .ZN(n7417) );
  XOR2_X1 U8938 ( .A(n7415), .B(n7417), .Z(n7256) );
  NOR2_X1 U8939 ( .A1(n7256), .A2(n7255), .ZN(n7416) );
  AOI21_X1 U8940 ( .B1(n7256), .B2(n7255), .A(n7416), .ZN(n7262) );
  NAND2_X1 U8941 ( .A1(n9230), .A2(n9183), .ZN(n7257) );
  OR2_X1 U8942 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5081), .ZN(n9653) );
  OAI211_X1 U8943 ( .C1(n7258), .C2(n9207), .A(n7257), .B(n9653), .ZN(n7260)
         );
  NOR2_X1 U8944 ( .A1(n9186), .A2(n9775), .ZN(n7259) );
  AOI211_X1 U8945 ( .C1(n9188), .C2(n9773), .A(n7260), .B(n7259), .ZN(n7261)
         );
  OAI21_X1 U8946 ( .B1(n7262), .B2(n9201), .A(n7261), .ZN(P1_U3225) );
  XNOR2_X1 U8947 ( .A(n7263), .B(n8317), .ZN(n9909) );
  INV_X1 U8948 ( .A(n9909), .ZN(n7278) );
  NAND2_X1 U8949 ( .A1(n7264), .A2(n8347), .ZN(n7266) );
  XNOR2_X1 U8950 ( .A(n7266), .B(n7265), .ZN(n7267) );
  OAI222_X1 U8951 ( .A1(n8950), .A2(n7269), .B1(n8952), .B2(n7268), .C1(n7267), 
        .C2(n8970), .ZN(n9907) );
  OAI21_X1 U8952 ( .B1(n6944), .B2(n7271), .A(n7270), .ZN(n9906) );
  INV_X1 U8953 ( .A(n8936), .ZN(n8987) );
  INV_X1 U8954 ( .A(n8934), .ZN(n8985) );
  AOI22_X1 U8955 ( .A1(n8987), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n7272), .B2(
        n8985), .ZN(n7275) );
  NAND2_X1 U8956 ( .A1(n8845), .A2(n7273), .ZN(n7274) );
  OAI211_X1 U8957 ( .C1(n9906), .C2(n8801), .A(n7275), .B(n7274), .ZN(n7276)
         );
  AOI21_X1 U8958 ( .B1(n9907), .B2(n8936), .A(n7276), .ZN(n7277) );
  OAI21_X1 U8959 ( .B1(n9003), .B2(n7278), .A(n7277), .ZN(P2_U3290) );
  OR2_X1 U8960 ( .A1(n7482), .A2(n9911), .ZN(n7279) );
  NAND2_X1 U8961 ( .A1(n7280), .A2(n7279), .ZN(n7356) );
  NAND2_X1 U8962 ( .A1(n7286), .A2(n9099), .ZN(n8394) );
  INV_X1 U8963 ( .A(n7286), .ZN(n8657) );
  INV_X1 U8964 ( .A(n9099), .ZN(n7363) );
  NAND2_X1 U8965 ( .A1(n8657), .A2(n7363), .ZN(n8391) );
  NAND2_X1 U8966 ( .A1(n7286), .A2(n7363), .ZN(n7281) );
  AND2_X1 U8967 ( .A1(n7283), .A2(n7281), .ZN(n7284) );
  NOR2_X1 U8968 ( .A1(n8656), .A2(n9917), .ZN(n7343) );
  INV_X1 U8969 ( .A(n7343), .ZN(n8402) );
  NAND2_X1 U8970 ( .A1(n8656), .A2(n9917), .ZN(n8396) );
  INV_X1 U8971 ( .A(n8395), .ZN(n8321) );
  AND2_X1 U8972 ( .A1(n8321), .A2(n7281), .ZN(n7282) );
  OAI21_X1 U8973 ( .B1(n7284), .B2(n8321), .A(n7342), .ZN(n9916) );
  NAND2_X1 U8974 ( .A1(n7285), .A2(n8383), .ZN(n7354) );
  NAND2_X1 U8975 ( .A1(n7354), .A2(n8319), .ZN(n7353) );
  NAND2_X1 U8976 ( .A1(n7353), .A2(n8394), .ZN(n7344) );
  XNOR2_X1 U8977 ( .A(n7344), .B(n8395), .ZN(n7288) );
  OAI22_X1 U8978 ( .A1(n7286), .A2(n8952), .B1(n7671), .B2(n8950), .ZN(n7287)
         );
  AOI21_X1 U8979 ( .B1(n7288), .B2(n8998), .A(n7287), .ZN(n7289) );
  OAI21_X1 U8980 ( .B1(n9916), .B2(n7797), .A(n7289), .ZN(n9919) );
  NAND2_X1 U8981 ( .A1(n9919), .A2(n8936), .ZN(n7295) );
  INV_X1 U8982 ( .A(n9917), .ZN(n7341) );
  OAI22_X1 U8983 ( .A1(n8936), .A2(n7290), .B1(n7610), .B2(n8934), .ZN(n7293)
         );
  INV_X1 U8984 ( .A(n7347), .ZN(n7291) );
  OAI21_X1 U8985 ( .B1(n9917), .B2(n4456), .A(n7291), .ZN(n9918) );
  NOR2_X1 U8986 ( .A1(n9918), .A2(n8801), .ZN(n7292) );
  AOI211_X1 U8987 ( .C1(n8845), .C2(n7341), .A(n7293), .B(n7292), .ZN(n7294)
         );
  OAI211_X1 U8988 ( .C1(n9916), .C2(n7807), .A(n7295), .B(n7294), .ZN(P2_U3286) );
  NAND2_X1 U8989 ( .A1(n7298), .A2(n9127), .ZN(n7296) );
  OAI211_X1 U8990 ( .C1(n7297), .C2(n10258), .A(n7296), .B(n8500), .ZN(
        P2_U3335) );
  NAND2_X1 U8991 ( .A1(n7298), .A2(n9535), .ZN(n7300) );
  NAND2_X1 U8992 ( .A1(n7299), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8252) );
  OAI211_X1 U8993 ( .C1(n7301), .C2(n9531), .A(n7300), .B(n8252), .ZN(P1_U3330) );
  XNOR2_X1 U8994 ( .A(n7303), .B(n7302), .ZN(n7304) );
  XNOR2_X1 U8995 ( .A(n7305), .B(n7304), .ZN(n7312) );
  INV_X1 U8996 ( .A(n7571), .ZN(n7306) );
  NAND2_X1 U8997 ( .A1(n9211), .A2(n7306), .ZN(n7309) );
  AOI21_X1 U8998 ( .B1(n9194), .B2(n9227), .A(n7307), .ZN(n7308) );
  OAI211_X1 U8999 ( .C1(n9576), .C2(n9208), .A(n7309), .B(n7308), .ZN(n7310)
         );
  AOI21_X1 U9000 ( .B1(n9199), .B2(n7574), .A(n7310), .ZN(n7311) );
  OAI21_X1 U9001 ( .B1(n7312), .B2(n9201), .A(n7311), .ZN(P1_U3215) );
  INV_X1 U9002 ( .A(n7313), .ZN(n7314) );
  AOI22_X1 U9003 ( .A1(n8987), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n7314), .B2(
        n8985), .ZN(n7315) );
  OAI21_X1 U9004 ( .B1(n8989), .B2(n7316), .A(n7315), .ZN(n7319) );
  INV_X1 U9005 ( .A(n8936), .ZN(n8956) );
  NOR2_X1 U9006 ( .A1(n7317), .A2(n8956), .ZN(n7318) );
  AOI211_X1 U9007 ( .C1(n7320), .C2(n9001), .A(n7319), .B(n7318), .ZN(n7321)
         );
  OAI21_X1 U9008 ( .B1(n9003), .B2(n7322), .A(n7321), .ZN(P2_U3289) );
  NOR2_X1 U9009 ( .A1(n8987), .A2(n8342), .ZN(n8977) );
  INV_X1 U9010 ( .A(n7323), .ZN(n8585) );
  AOI22_X1 U9011 ( .A1(n8987), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n8585), .B2(
        n8985), .ZN(n7324) );
  OAI21_X1 U9012 ( .B1(n8989), .B2(n7325), .A(n7324), .ZN(n7328) );
  NOR2_X1 U9013 ( .A1(n7326), .A2(n9003), .ZN(n7327) );
  AOI211_X1 U9014 ( .C1(n7329), .C2(n8977), .A(n7328), .B(n7327), .ZN(n7330)
         );
  OAI21_X1 U9015 ( .B1(n8956), .B2(n7331), .A(n7330), .ZN(P2_U3291) );
  INV_X1 U9016 ( .A(n7332), .ZN(n7339) );
  INV_X1 U9017 ( .A(n9425), .ZN(n9599) );
  OAI22_X1 U9018 ( .A1(n9410), .A2(n7333), .B1(n6513), .B2(n9785), .ZN(n7338)
         );
  INV_X1 U9019 ( .A(n9776), .ZN(n9588) );
  AOI22_X1 U9020 ( .A1(n7334), .A2(n9778), .B1(n9588), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n7335) );
  AOI21_X1 U9021 ( .B1(n7336), .B2(n7335), .A(n9787), .ZN(n7337) );
  AOI211_X1 U9022 ( .C1(n7339), .C2(n9599), .A(n7338), .B(n7337), .ZN(n7340)
         );
  INV_X1 U9023 ( .A(n7340), .ZN(P1_U3290) );
  INV_X1 U9024 ( .A(n7671), .ZN(n8655) );
  NAND2_X1 U9025 ( .A1(n7369), .A2(n8655), .ZN(n8397) );
  NAND2_X1 U9026 ( .A1(n7671), .A2(n9094), .ZN(n8406) );
  XNOR2_X1 U9027 ( .A(n7368), .B(n7367), .ZN(n9098) );
  XNOR2_X1 U9028 ( .A(n7372), .B(n7367), .ZN(n7345) );
  INV_X1 U9029 ( .A(n7715), .ZN(n8654) );
  AOI222_X1 U9030 ( .A1(n8998), .A2(n7345), .B1(n8654), .B2(n8993), .C1(n8656), 
        .C2(n8995), .ZN(n9097) );
  OAI21_X1 U9031 ( .B1(n8625), .B2(n8934), .A(n9097), .ZN(n7346) );
  NAND2_X1 U9032 ( .A1(n7346), .A2(n8936), .ZN(n7352) );
  OR2_X1 U9033 ( .A1(n7347), .A2(n7369), .ZN(n7348) );
  NAND2_X1 U9034 ( .A1(n7347), .A2(n7369), .ZN(n7375) );
  AND2_X1 U9035 ( .A1(n7348), .A2(n7375), .ZN(n9095) );
  OAI22_X1 U9036 ( .A1(n8989), .A2(n7369), .B1(n8936), .B2(n7349), .ZN(n7350)
         );
  AOI21_X1 U9037 ( .B1(n9095), .B2(n9001), .A(n7350), .ZN(n7351) );
  OAI211_X1 U9038 ( .C1(n9003), .C2(n9098), .A(n7352), .B(n7351), .ZN(P2_U3285) );
  OAI21_X1 U9039 ( .B1(n8319), .B2(n7354), .A(n7353), .ZN(n7359) );
  INV_X1 U9040 ( .A(n8656), .ZN(n7480) );
  OAI22_X1 U9041 ( .A1(n7480), .A2(n8950), .B1(n7482), .B2(n8952), .ZN(n7358)
         );
  INV_X1 U9042 ( .A(n7283), .ZN(n7355) );
  AOI21_X1 U9043 ( .B1(n8319), .B2(n7356), .A(n7355), .ZN(n9104) );
  NOR2_X1 U9044 ( .A1(n9104), .A2(n7797), .ZN(n7357) );
  AOI211_X1 U9045 ( .C1(n8998), .C2(n7359), .A(n7358), .B(n7357), .ZN(n9102)
         );
  AOI21_X1 U9046 ( .B1(n9099), .B2(n7360), .A(n4456), .ZN(n9100) );
  INV_X1 U9047 ( .A(n7481), .ZN(n7361) );
  AOI22_X1 U9048 ( .A1(n8987), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7361), .B2(
        n8985), .ZN(n7362) );
  OAI21_X1 U9049 ( .B1(n8989), .B2(n7363), .A(n7362), .ZN(n7365) );
  NOR2_X1 U9050 ( .A1(n9104), .A2(n7807), .ZN(n7364) );
  AOI211_X1 U9051 ( .C1(n9100), .C2(n9001), .A(n7365), .B(n7364), .ZN(n7366)
         );
  OAI21_X1 U9052 ( .B1(n9102), .B2(n8956), .A(n7366), .ZN(P2_U3287) );
  NAND2_X1 U9053 ( .A1(n7368), .A2(n7367), .ZN(n7371) );
  OR2_X1 U9054 ( .A1(n7369), .A2(n7671), .ZN(n7370) );
  OR2_X1 U9055 ( .A1(n9924), .A2(n7715), .ZN(n8409) );
  NAND2_X1 U9056 ( .A1(n9924), .A2(n7715), .ZN(n8410) );
  XNOR2_X1 U9057 ( .A(n7487), .B(n8324), .ZN(n9932) );
  INV_X1 U9058 ( .A(n9932), .ZN(n7382) );
  NAND2_X1 U9059 ( .A1(n7490), .A2(n8397), .ZN(n7373) );
  XNOR2_X1 U9060 ( .A(n7373), .B(n8324), .ZN(n7374) );
  OAI222_X1 U9061 ( .A1(n8950), .A2(n7838), .B1(n8952), .B2(n7671), .C1(n8970), 
        .C2(n7374), .ZN(n9929) );
  NAND2_X1 U9062 ( .A1(n7375), .A2(n9924), .ZN(n7376) );
  NAND2_X1 U9063 ( .A1(n7498), .A2(n7376), .ZN(n9928) );
  OAI22_X1 U9064 ( .A1(n8936), .A2(n7377), .B1(n7670), .B2(n8934), .ZN(n7378)
         );
  AOI21_X1 U9065 ( .B1(n8845), .B2(n9924), .A(n7378), .ZN(n7379) );
  OAI21_X1 U9066 ( .B1(n9928), .B2(n8801), .A(n7379), .ZN(n7380) );
  AOI21_X1 U9067 ( .B1(n9929), .B2(n8936), .A(n7380), .ZN(n7381) );
  OAI21_X1 U9068 ( .B1(n9003), .B2(n7382), .A(n7381), .ZN(P2_U3284) );
  OAI21_X1 U9069 ( .B1(n4446), .B2(n5115), .A(n7398), .ZN(n7383) );
  AOI222_X1 U9070 ( .A1(n9586), .A2(n7383), .B1(n9228), .B2(n9417), .C1(n9230), 
        .C2(n9419), .ZN(n9818) );
  MUX2_X1 U9071 ( .A(n7384), .B(n9818), .S(n9785), .Z(n7391) );
  OAI21_X1 U9072 ( .B1(n7386), .B2(n7385), .A(n7403), .ZN(n9821) );
  OAI211_X1 U9073 ( .C1(n7433), .C2(n9819), .A(n9595), .B(n7406), .ZN(n9817)
         );
  NOR2_X1 U9074 ( .A1(n9817), .A2(n9329), .ZN(n7389) );
  OAI22_X1 U9075 ( .A1(n9410), .A2(n9819), .B1(n7387), .B2(n9776), .ZN(n7388)
         );
  AOI211_X1 U9076 ( .C1(n9821), .C2(n9599), .A(n7389), .B(n7388), .ZN(n7390)
         );
  NAND2_X1 U9077 ( .A1(n7391), .A2(n7390), .ZN(P1_U3284) );
  XNOR2_X1 U9078 ( .A(n7523), .B(n7522), .ZN(n7397) );
  NOR2_X1 U9079 ( .A1(n7935), .A2(n9207), .ZN(n7392) );
  AOI211_X1 U9080 ( .C1(n9183), .C2(n9224), .A(n7393), .B(n7392), .ZN(n7394)
         );
  OAI21_X1 U9081 ( .B1(n9186), .B2(n7513), .A(n7394), .ZN(n7395) );
  AOI21_X1 U9082 ( .B1(n9199), .B2(n7516), .A(n7395), .ZN(n7396) );
  OAI21_X1 U9083 ( .B1(n7397), .B2(n9201), .A(n7396), .ZN(P1_U3234) );
  NAND2_X1 U9084 ( .A1(n7398), .A2(n7977), .ZN(n7399) );
  XOR2_X1 U9085 ( .A(n8099), .B(n7399), .Z(n7400) );
  OAI222_X1 U9086 ( .A1(n9577), .A2(n7401), .B1(n5559), .B2(n7427), .C1(n7400), 
        .C2(n5556), .ZN(n9825) );
  INV_X1 U9087 ( .A(n9825), .ZN(n7414) );
  NAND2_X1 U9088 ( .A1(n7403), .A2(n7402), .ZN(n7405) );
  OR2_X1 U9089 ( .A1(n7405), .A2(n8099), .ZN(n7618) );
  INV_X1 U9090 ( .A(n7618), .ZN(n7404) );
  AOI21_X1 U9091 ( .B1(n8099), .B2(n7405), .A(n7404), .ZN(n9828) );
  NAND2_X1 U9092 ( .A1(n7406), .A2(n7410), .ZN(n7407) );
  NAND2_X1 U9093 ( .A1(n7625), .A2(n7407), .ZN(n9824) );
  OAI22_X1 U9094 ( .A1(n9785), .A2(n9659), .B1(n7408), .B2(n9776), .ZN(n7409)
         );
  AOI21_X1 U9095 ( .B1(n9590), .B2(n7410), .A(n7409), .ZN(n7411) );
  OAI21_X1 U9096 ( .B1(n9824), .B2(n9281), .A(n7411), .ZN(n7412) );
  AOI21_X1 U9097 ( .B1(n9828), .B2(n9599), .A(n7412), .ZN(n7413) );
  OAI21_X1 U9098 ( .B1(n9787), .B2(n7414), .A(n7413), .ZN(P1_U3283) );
  INV_X1 U9099 ( .A(n7415), .ZN(n7418) );
  AOI21_X1 U9100 ( .B1(n7418), .B2(n7417), .A(n7416), .ZN(n7422) );
  XNOR2_X1 U9101 ( .A(n7420), .B(n7419), .ZN(n7421) );
  XNOR2_X1 U9102 ( .A(n7422), .B(n7421), .ZN(n7430) );
  INV_X1 U9103 ( .A(n7423), .ZN(n7436) );
  NAND2_X1 U9104 ( .A1(n9188), .A2(n7437), .ZN(n7426) );
  AOI21_X1 U9105 ( .B1(n9194), .B2(n9231), .A(n7424), .ZN(n7425) );
  OAI211_X1 U9106 ( .C1(n7427), .C2(n9208), .A(n7426), .B(n7425), .ZN(n7428)
         );
  AOI21_X1 U9107 ( .B1(n7436), .B2(n9211), .A(n7428), .ZN(n7429) );
  OAI21_X1 U9108 ( .B1(n7430), .B2(n9201), .A(n7429), .ZN(P1_U3237) );
  OAI21_X1 U9109 ( .B1(n7432), .B2(n8095), .A(n7431), .ZN(n9816) );
  INV_X1 U9110 ( .A(n7433), .ZN(n7434) );
  OAI21_X1 U9111 ( .B1(n9812), .B2(n7435), .A(n7434), .ZN(n9813) );
  AOI22_X1 U9112 ( .A1(n9590), .A2(n7437), .B1(n7436), .B2(n9588), .ZN(n7438)
         );
  OAI21_X1 U9113 ( .B1(n9813), .B2(n9281), .A(n7438), .ZN(n7448) );
  INV_X1 U9114 ( .A(n7439), .ZN(n7440) );
  AND2_X1 U9115 ( .A1(n7440), .A2(n8139), .ZN(n8142) );
  NAND2_X1 U9116 ( .A1(n7441), .A2(n8142), .ZN(n7443) );
  NAND2_X1 U9117 ( .A1(n7443), .A2(n7442), .ZN(n7976) );
  OR2_X1 U9118 ( .A1(n7976), .A2(n8095), .ZN(n7992) );
  NAND2_X1 U9119 ( .A1(n7976), .A2(n8095), .ZN(n7444) );
  NAND3_X1 U9120 ( .A1(n7992), .A2(n9586), .A3(n7444), .ZN(n7446) );
  AOI22_X1 U9121 ( .A1(n9229), .A2(n9417), .B1(n9419), .B2(n9231), .ZN(n7445)
         );
  NAND2_X1 U9122 ( .A1(n7446), .A2(n7445), .ZN(n9814) );
  MUX2_X1 U9123 ( .A(n9814), .B(P1_REG2_REG_6__SCAN_IN), .S(n9787), .Z(n7447)
         );
  AOI211_X1 U9124 ( .C1(n9599), .C2(n9816), .A(n7448), .B(n7447), .ZN(n7449)
         );
  INV_X1 U9125 ( .A(n7449), .ZN(P1_U3285) );
  NOR2_X1 U9126 ( .A1(n8672), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7452) );
  AOI21_X1 U9127 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n8672), .A(n7452), .ZN(
        n8669) );
  NAND2_X1 U9128 ( .A1(n8668), .A2(n8669), .ZN(n8667) );
  OAI21_X1 U9129 ( .B1(n8672), .B2(P2_REG2_REG_11__SCAN_IN), .A(n8667), .ZN(
        n7455) );
  NAND2_X1 U9130 ( .A1(n7599), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7453) );
  OAI21_X1 U9131 ( .B1(n7599), .B2(P2_REG2_REG_12__SCAN_IN), .A(n7453), .ZN(
        n7454) );
  NOR2_X1 U9132 ( .A1(n7454), .A2(n7455), .ZN(n7598) );
  AOI211_X1 U9133 ( .C1(n7455), .C2(n7454), .A(n7598), .B(n9549), .ZN(n7468)
         );
  INV_X1 U9134 ( .A(n9853), .ZN(n9859) );
  MUX2_X1 U9135 ( .A(n7456), .B(P2_REG1_REG_12__SCAN_IN), .S(n7599), .Z(n7462)
         );
  NAND2_X1 U9136 ( .A1(n8672), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7460) );
  MUX2_X1 U9137 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7457), .S(n8672), .Z(n8674)
         );
  OAI21_X1 U9138 ( .B1(n7459), .B2(n6992), .A(n7458), .ZN(n8675) );
  NAND2_X1 U9139 ( .A1(n8674), .A2(n8675), .ZN(n8673) );
  NAND2_X1 U9140 ( .A1(n7460), .A2(n8673), .ZN(n7461) );
  NOR2_X1 U9141 ( .A1(n7461), .A2(n7462), .ZN(n7594) );
  AOI21_X1 U9142 ( .B1(n7462), .B2(n7461), .A(n7594), .ZN(n7466) );
  NAND2_X1 U9143 ( .A1(n9555), .A2(n7599), .ZN(n7465) );
  NAND2_X1 U9144 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7669) );
  INV_X1 U9145 ( .A(n7669), .ZN(n7463) );
  AOI21_X1 U9146 ( .B1(n9854), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7463), .ZN(
        n7464) );
  OAI211_X1 U9147 ( .C1(n9859), .C2(n7466), .A(n7465), .B(n7464), .ZN(n7467)
         );
  OR2_X1 U9148 ( .A1(n7468), .A2(n7467), .ZN(P2_U3257) );
  INV_X1 U9149 ( .A(n7469), .ZN(n7473) );
  OAI222_X1 U9150 ( .A1(n7471), .A2(P1_U3084), .B1(n7920), .B2(n7473), .C1(
        n7470), .C2(n7924), .ZN(P1_U3329) );
  OAI222_X1 U9151 ( .A1(P2_U3152), .A2(n7474), .B1(n7928), .B2(n7473), .C1(
        n7472), .C2(n10258), .ZN(P2_U3334) );
  INV_X1 U9152 ( .A(n7476), .ZN(n7477) );
  AOI21_X1 U9153 ( .B1(n7475), .B2(n7478), .A(n7477), .ZN(n7486) );
  OAI21_X1 U9154 ( .B1(n8613), .B2(n7480), .A(n7479), .ZN(n7484) );
  OAI22_X1 U9155 ( .A1(n8614), .A2(n7482), .B1(n8640), .B2(n7481), .ZN(n7483)
         );
  AOI211_X1 U9156 ( .C1(n9099), .C2(n8629), .A(n7484), .B(n7483), .ZN(n7485)
         );
  OAI21_X1 U9157 ( .B1(n7486), .B2(n8643), .A(n7485), .ZN(P2_U3233) );
  NAND2_X1 U9158 ( .A1(n9089), .A2(n7838), .ZN(n7535) );
  NAND2_X1 U9159 ( .A1(n8414), .A2(n7535), .ZN(n7491) );
  NAND2_X1 U9160 ( .A1(n7488), .A2(n4827), .ZN(n7489) );
  AND2_X1 U9161 ( .A1(n7534), .A2(n7489), .ZN(n9088) );
  OAI22_X1 U9162 ( .A1(n7715), .A2(n8952), .B1(n7898), .B2(n8950), .ZN(n7496)
         );
  AND2_X1 U9163 ( .A1(n8409), .A2(n8397), .ZN(n8405) );
  INV_X1 U9164 ( .A(n7536), .ZN(n7494) );
  NAND3_X1 U9165 ( .A1(n7492), .A2(n7491), .A3(n8410), .ZN(n7493) );
  AOI21_X1 U9166 ( .B1(n7494), .B2(n7493), .A(n8970), .ZN(n7495) );
  AOI211_X1 U9167 ( .C1(n9088), .C2(n7497), .A(n7496), .B(n7495), .ZN(n9092)
         );
  AOI21_X1 U9168 ( .B1(n9089), .B2(n7498), .A(n7540), .ZN(n9090) );
  INV_X1 U9169 ( .A(n9089), .ZN(n7720) );
  NOR2_X1 U9170 ( .A1(n8989), .A2(n7720), .ZN(n7501) );
  OAI22_X1 U9171 ( .A1(n8936), .A2(n7499), .B1(n7714), .B2(n8934), .ZN(n7500)
         );
  AOI211_X1 U9172 ( .C1(n9090), .C2(n9001), .A(n7501), .B(n7500), .ZN(n7504)
         );
  INV_X1 U9173 ( .A(n7807), .ZN(n7502) );
  NAND2_X1 U9174 ( .A1(n9088), .A2(n7502), .ZN(n7503) );
  OAI211_X1 U9175 ( .C1(n9092), .C2(n8956), .A(n7504), .B(n7503), .ZN(P2_U3283) );
  XNOR2_X1 U9176 ( .A(n7516), .B(n9576), .ZN(n8010) );
  XNOR2_X1 U9177 ( .A(n7505), .B(n8010), .ZN(n9510) );
  INV_X1 U9178 ( .A(n8010), .ZN(n8104) );
  XNOR2_X1 U9179 ( .A(n7506), .B(n8104), .ZN(n7509) );
  OAI22_X1 U9180 ( .A1(n7551), .A2(n9577), .B1(n7935), .B2(n5559), .ZN(n7507)
         );
  INV_X1 U9181 ( .A(n7507), .ZN(n7508) );
  OAI21_X1 U9182 ( .B1(n7509), .B2(n5556), .A(n7508), .ZN(n7510) );
  AOI21_X1 U9183 ( .B1(n9510), .B2(n7511), .A(n7510), .ZN(n9512) );
  OR2_X1 U9184 ( .A1(n7569), .A2(n9507), .ZN(n7512) );
  NAND2_X1 U9185 ( .A1(n9592), .A2(n7512), .ZN(n9508) );
  OAI22_X1 U9186 ( .A1(n9785), .A2(n7514), .B1(n7513), .B2(n9776), .ZN(n7515)
         );
  AOI21_X1 U9187 ( .B1(n7516), .B2(n9590), .A(n7515), .ZN(n7517) );
  OAI21_X1 U9188 ( .B1(n9508), .B2(n9281), .A(n7517), .ZN(n7518) );
  AOI21_X1 U9189 ( .B1(n9510), .B2(n9599), .A(n7518), .ZN(n7519) );
  OAI21_X1 U9190 ( .B1(n9512), .B2(n9787), .A(n7519), .ZN(P1_U3280) );
  NAND2_X1 U9191 ( .A1(n7521), .A2(n7520), .ZN(n7527) );
  NAND2_X1 U9192 ( .A1(n7523), .A2(n7522), .ZN(n7525) );
  NAND2_X1 U9193 ( .A1(n7525), .A2(n7524), .ZN(n7526) );
  XOR2_X1 U9194 ( .A(n7527), .B(n7526), .Z(n7533) );
  NOR2_X1 U9195 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7528), .ZN(n9674) );
  NOR2_X1 U9196 ( .A1(n9578), .A2(n9208), .ZN(n7529) );
  AOI211_X1 U9197 ( .C1(n9194), .C2(n9225), .A(n9674), .B(n7529), .ZN(n7530)
         );
  OAI21_X1 U9198 ( .B1(n9186), .B2(n9587), .A(n7530), .ZN(n7531) );
  AOI21_X1 U9199 ( .B1(n9199), .B2(n9593), .A(n7531), .ZN(n7532) );
  OAI21_X1 U9200 ( .B1(n7533), .B2(n9201), .A(n7532), .ZN(P1_U3222) );
  INV_X1 U9201 ( .A(n7838), .ZN(n8653) );
  NAND2_X1 U9202 ( .A1(n7841), .A2(n7898), .ZN(n8421) );
  XNOR2_X1 U9203 ( .A(n7635), .B(n8327), .ZN(n9572) );
  INV_X1 U9204 ( .A(n9572), .ZN(n7546) );
  INV_X1 U9205 ( .A(n7535), .ZN(n8416) );
  NAND2_X1 U9206 ( .A1(n7537), .A2(n8327), .ZN(n7631) );
  OAI211_X1 U9207 ( .C1(n7537), .C2(n8327), .A(n7631), .B(n8998), .ZN(n7539)
         );
  INV_X1 U9208 ( .A(n8576), .ZN(n8651) );
  AOI22_X1 U9209 ( .A1(n8993), .A2(n8651), .B1(n8653), .B2(n8995), .ZN(n7538)
         );
  NAND2_X1 U9210 ( .A1(n7539), .A2(n7538), .ZN(n9570) );
  INV_X1 U9211 ( .A(n7841), .ZN(n9568) );
  NAND2_X1 U9212 ( .A1(n7540), .A2(n9568), .ZN(n7637) );
  OAI21_X1 U9213 ( .B1(n7540), .B2(n9568), .A(n7637), .ZN(n9569) );
  OAI22_X1 U9214 ( .A1(n8936), .A2(n7541), .B1(n7837), .B2(n8934), .ZN(n7542)
         );
  AOI21_X1 U9215 ( .B1(n7841), .B2(n8845), .A(n7542), .ZN(n7543) );
  OAI21_X1 U9216 ( .B1(n9569), .B2(n8801), .A(n7543), .ZN(n7544) );
  AOI21_X1 U9217 ( .B1(n9570), .B2(n8936), .A(n7544), .ZN(n7545) );
  OAI21_X1 U9218 ( .B1(n7546), .B2(n9003), .A(n7545), .ZN(P2_U3282) );
  XOR2_X1 U9219 ( .A(n7548), .B(n7547), .Z(n7549) );
  XNOR2_X1 U9220 ( .A(n7550), .B(n7549), .ZN(n7556) );
  AND2_X1 U9221 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9683) );
  NOR2_X1 U9222 ( .A1(n7551), .A2(n9207), .ZN(n7552) );
  AOI211_X1 U9223 ( .C1(n9183), .C2(n9222), .A(n9683), .B(n7552), .ZN(n7553)
         );
  OAI21_X1 U9224 ( .B1(n9186), .B2(n7768), .A(n7553), .ZN(n7554) );
  AOI21_X1 U9225 ( .B1(n9501), .B2(n9199), .A(n7554), .ZN(n7555) );
  OAI21_X1 U9226 ( .B1(n7556), .B2(n9201), .A(n7555), .ZN(P1_U3232) );
  NAND2_X1 U9227 ( .A1(n7557), .A2(n7993), .ZN(n7621) );
  AND2_X1 U9228 ( .A1(n7994), .A2(n7983), .ZN(n8100) );
  NAND2_X1 U9229 ( .A1(n7621), .A2(n8100), .ZN(n7620) );
  NAND2_X1 U9230 ( .A1(n7620), .A2(n7994), .ZN(n7558) );
  XOR2_X1 U9231 ( .A(n8101), .B(n7558), .Z(n7559) );
  AOI222_X1 U9232 ( .A1(n9586), .A2(n7559), .B1(n9225), .B2(n9417), .C1(n9227), 
        .C2(n9419), .ZN(n9563) );
  NAND2_X1 U9233 ( .A1(n7618), .A2(n7560), .ZN(n7562) );
  NAND2_X1 U9234 ( .A1(n7562), .A2(n7561), .ZN(n7568) );
  NAND2_X1 U9235 ( .A1(n7618), .A2(n7563), .ZN(n7565) );
  AND2_X1 U9236 ( .A1(n7565), .A2(n7564), .ZN(n7566) );
  OAI21_X1 U9237 ( .B1(n7568), .B2(n7567), .A(n7566), .ZN(n9566) );
  OAI21_X1 U9238 ( .B1(n4457), .B2(n9564), .A(n9595), .ZN(n7570) );
  OR2_X1 U9239 ( .A1(n7570), .A2(n7569), .ZN(n9562) );
  OAI22_X1 U9240 ( .A1(n9785), .A2(n7572), .B1(n7571), .B2(n9776), .ZN(n7573)
         );
  AOI21_X1 U9241 ( .B1(n7574), .B2(n9590), .A(n7573), .ZN(n7575) );
  OAI21_X1 U9242 ( .B1(n9562), .B2(n9329), .A(n7575), .ZN(n7576) );
  AOI21_X1 U9243 ( .B1(n9566), .B2(n9599), .A(n7576), .ZN(n7577) );
  OAI21_X1 U9244 ( .B1(n9563), .B2(n9787), .A(n7577), .ZN(P1_U3281) );
  XNOR2_X1 U9245 ( .A(n7579), .B(n7578), .ZN(n7580) );
  XNOR2_X1 U9246 ( .A(n7581), .B(n7580), .ZN(n7587) );
  NOR2_X1 U9247 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7582), .ZN(n9698) );
  NOR2_X1 U9248 ( .A1(n7858), .A2(n9208), .ZN(n7583) );
  AOI211_X1 U9249 ( .C1(n9194), .C2(n9223), .A(n9698), .B(n7583), .ZN(n7584)
         );
  OAI21_X1 U9250 ( .B1(n9186), .B2(n7748), .A(n7584), .ZN(n7585) );
  AOI21_X1 U9251 ( .B1(n7751), .B2(n9199), .A(n7585), .ZN(n7586) );
  OAI21_X1 U9252 ( .B1(n7587), .B2(n9201), .A(n7586), .ZN(P1_U3213) );
  INV_X1 U9253 ( .A(n7588), .ZN(n7592) );
  OAI222_X1 U9254 ( .A1(n8511), .A2(n7590), .B1(n7928), .B2(n7592), .C1(
        P2_U3152), .C2(n7589), .ZN(P2_U3333) );
  OAI222_X1 U9255 ( .A1(n7924), .A2(n7593), .B1(n7920), .B2(n7592), .C1(n7591), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  AOI21_X1 U9256 ( .B1(n7595), .B2(n7456), .A(n7594), .ZN(n7597) );
  AOI22_X1 U9257 ( .A1(n7655), .A2(n5935), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7651), .ZN(n7596) );
  NOR2_X1 U9258 ( .A1(n7597), .A2(n7596), .ZN(n7650) );
  AOI21_X1 U9259 ( .B1(n7597), .B2(n7596), .A(n7650), .ZN(n7607) );
  NOR2_X1 U9260 ( .A1(n7655), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7600) );
  AOI21_X1 U9261 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n7655), .A(n7600), .ZN(
        n7601) );
  OAI21_X1 U9262 ( .B1(n7602), .B2(n7601), .A(n7654), .ZN(n7603) );
  INV_X1 U9263 ( .A(n9549), .ZN(n9856) );
  NAND2_X1 U9264 ( .A1(n7603), .A2(n9856), .ZN(n7606) );
  INV_X1 U9265 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n9980) );
  NOR2_X1 U9266 ( .A1(n9980), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7717) );
  NOR2_X1 U9267 ( .A1(n9857), .A2(n7651), .ZN(n7604) );
  AOI211_X1 U9268 ( .C1(P2_ADDR_REG_13__SCAN_IN), .C2(n9854), .A(n7717), .B(
        n7604), .ZN(n7605) );
  OAI211_X1 U9269 ( .C1(n7607), .C2(n9859), .A(n7606), .B(n7605), .ZN(P2_U3258) );
  XOR2_X1 U9270 ( .A(n7608), .B(n7609), .Z(n7615) );
  INV_X1 U9271 ( .A(n7610), .ZN(n7611) );
  AOI22_X1 U9272 ( .A1(n8628), .A2(n8657), .B1(n8627), .B2(n7611), .ZN(n7613)
         );
  AOI22_X1 U9273 ( .A1(n8624), .A2(n8655), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n7612) );
  OAI211_X1 U9274 ( .C1(n9917), .C2(n8619), .A(n7613), .B(n7612), .ZN(n7614)
         );
  AOI21_X1 U9275 ( .B1(n7615), .B2(n8622), .A(n7614), .ZN(n7616) );
  INV_X1 U9276 ( .A(n7616), .ZN(P2_U3219) );
  NAND2_X1 U9277 ( .A1(n7618), .A2(n7617), .ZN(n7619) );
  XOR2_X1 U9278 ( .A(n8100), .B(n7619), .Z(n9829) );
  AOI22_X1 U9279 ( .A1(n9419), .A2(n9228), .B1(n9226), .B2(n9417), .ZN(n7623)
         );
  OAI211_X1 U9280 ( .C1(n7621), .C2(n8100), .A(n7620), .B(n9586), .ZN(n7622)
         );
  OAI211_X1 U9281 ( .C1(n9829), .C2(n9582), .A(n7623), .B(n7622), .ZN(n9834)
         );
  NAND2_X1 U9282 ( .A1(n9834), .A2(n9785), .ZN(n7630) );
  OAI22_X1 U9283 ( .A1(n9785), .A2(n7624), .B1(n7939), .B2(n9776), .ZN(n7628)
         );
  AND2_X1 U9284 ( .A1(n7625), .A2(n9830), .ZN(n7626) );
  OR2_X1 U9285 ( .A1(n7626), .A2(n4457), .ZN(n9833) );
  NOR2_X1 U9286 ( .A1(n9833), .A2(n9281), .ZN(n7627) );
  AOI211_X1 U9287 ( .C1(n9590), .C2(n9830), .A(n7628), .B(n7627), .ZN(n7629)
         );
  OAI211_X1 U9288 ( .C1(n9829), .C2(n9425), .A(n7630), .B(n7629), .ZN(P1_U3282) );
  NAND2_X1 U9289 ( .A1(n7631), .A2(n8420), .ZN(n7791) );
  NOR2_X1 U9290 ( .A1(n7901), .A2(n8576), .ZN(n8428) );
  INV_X1 U9291 ( .A(n8428), .ZN(n7632) );
  NAND2_X1 U9292 ( .A1(n7901), .A2(n8576), .ZN(n8427) );
  NAND2_X1 U9293 ( .A1(n7632), .A2(n8427), .ZN(n8424) );
  XOR2_X1 U9294 ( .A(n7791), .B(n8424), .Z(n7633) );
  OAI222_X1 U9295 ( .A1(n8952), .A2(n7898), .B1(n8950), .B2(n7896), .C1(n8970), 
        .C2(n7633), .ZN(n7723) );
  INV_X1 U9296 ( .A(n7723), .ZN(n7644) );
  INV_X1 U9297 ( .A(n7898), .ZN(n8652) );
  OR2_X1 U9298 ( .A1(n7841), .A2(n8652), .ZN(n7634) );
  NAND2_X1 U9299 ( .A1(n7636), .A2(n8424), .ZN(n7794) );
  OAI21_X1 U9300 ( .B1(n7636), .B2(n8424), .A(n7794), .ZN(n7725) );
  NAND2_X1 U9301 ( .A1(n7637), .A2(n7901), .ZN(n7638) );
  NAND2_X1 U9302 ( .A1(n7803), .A2(n7638), .ZN(n7722) );
  OAI22_X1 U9303 ( .A1(n8936), .A2(n7639), .B1(n7897), .B2(n8934), .ZN(n7640)
         );
  AOI21_X1 U9304 ( .B1(n7901), .B2(n8845), .A(n7640), .ZN(n7641) );
  OAI21_X1 U9305 ( .B1(n7722), .B2(n8801), .A(n7641), .ZN(n7642) );
  AOI21_X1 U9306 ( .B1(n7725), .B2(n8905), .A(n7642), .ZN(n7643) );
  OAI21_X1 U9307 ( .B1(n7644), .B2(n8956), .A(n7643), .ZN(P2_U3281) );
  INV_X1 U9308 ( .A(n7645), .ZN(n7648) );
  OAI222_X1 U9309 ( .A1(P2_U3152), .A2(n7646), .B1(n7928), .B2(n7648), .C1(
        n10190), .C2(n10258), .ZN(P2_U3332) );
  OAI222_X1 U9310 ( .A1(n7649), .A2(P1_U3084), .B1(n7920), .B2(n7648), .C1(
        n7647), .C2(n7924), .ZN(P1_U3327) );
  AOI21_X1 U9311 ( .B1(n7651), .B2(n5935), .A(n7650), .ZN(n7653) );
  AOI22_X1 U9312 ( .A1(n8681), .A2(n5956), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n8687), .ZN(n7652) );
  NOR2_X1 U9313 ( .A1(n7653), .A2(n7652), .ZN(n8686) );
  AOI21_X1 U9314 ( .B1(n7653), .B2(n7652), .A(n8686), .ZN(n7664) );
  AOI22_X1 U9315 ( .A1(n8681), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7541), .B2(
        n8687), .ZN(n7657) );
  OAI21_X1 U9316 ( .B1(n7657), .B2(n7656), .A(n8680), .ZN(n7658) );
  NAND2_X1 U9317 ( .A1(n7658), .A2(n9856), .ZN(n7663) );
  INV_X1 U9318 ( .A(n9854), .ZN(n7660) );
  INV_X1 U9319 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7659) );
  NAND2_X1 U9320 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7836) );
  OAI21_X1 U9321 ( .B1(n7660), .B2(n7659), .A(n7836), .ZN(n7661) );
  AOI21_X1 U9322 ( .B1(n8681), .B2(n9555), .A(n7661), .ZN(n7662) );
  OAI211_X1 U9323 ( .C1(n7664), .C2(n9859), .A(n7663), .B(n7662), .ZN(P2_U3259) );
  NAND2_X1 U9324 ( .A1(n7666), .A2(n7665), .ZN(n7668) );
  XOR2_X1 U9325 ( .A(n7668), .B(n7667), .Z(n7675) );
  OAI21_X1 U9326 ( .B1(n8613), .B2(n7838), .A(n7669), .ZN(n7673) );
  OAI22_X1 U9327 ( .A1(n8614), .A2(n7671), .B1(n8640), .B2(n7670), .ZN(n7672)
         );
  AOI211_X1 U9328 ( .C1(n9924), .C2(n8629), .A(n7673), .B(n7672), .ZN(n7674)
         );
  OAI21_X1 U9329 ( .B1(n7675), .B2(n8643), .A(n7674), .ZN(P2_U3226) );
  INV_X1 U9330 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10270) );
  NOR2_X1 U9331 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7676) );
  AOI21_X1 U9332 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7676), .ZN(n9955) );
  NOR2_X1 U9333 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7677) );
  AOI21_X1 U9334 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7677), .ZN(n9958) );
  NOR2_X1 U9335 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7678) );
  AOI21_X1 U9336 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7678), .ZN(n9961) );
  NOR2_X1 U9337 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7679) );
  AOI21_X1 U9338 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7679), .ZN(n9964) );
  NOR2_X1 U9339 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7680) );
  AOI21_X1 U9340 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7680), .ZN(n9967) );
  NOR2_X1 U9341 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7687) );
  XNOR2_X1 U9342 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10281) );
  NAND2_X1 U9343 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7685) );
  XOR2_X1 U9344 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10279) );
  NAND2_X1 U9345 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7683) );
  XOR2_X1 U9346 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10277) );
  AOI21_X1 U9347 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9948) );
  INV_X1 U9348 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7681) );
  NAND3_X1 U9349 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9950) );
  OAI21_X1 U9350 ( .B1(n9948), .B2(n7681), .A(n9950), .ZN(n10276) );
  NAND2_X1 U9351 ( .A1(n10277), .A2(n10276), .ZN(n7682) );
  NAND2_X1 U9352 ( .A1(n7683), .A2(n7682), .ZN(n10278) );
  NAND2_X1 U9353 ( .A1(n10279), .A2(n10278), .ZN(n7684) );
  NAND2_X1 U9354 ( .A1(n7685), .A2(n7684), .ZN(n10280) );
  NOR2_X1 U9355 ( .A1(n10281), .A2(n10280), .ZN(n7686) );
  NOR2_X1 U9356 ( .A1(n7687), .A2(n7686), .ZN(n7688) );
  NOR2_X1 U9357 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7688), .ZN(n10266) );
  AND2_X1 U9358 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7688), .ZN(n10265) );
  NOR2_X1 U9359 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10265), .ZN(n7689) );
  NOR2_X1 U9360 ( .A1(n10266), .A2(n7689), .ZN(n7690) );
  NAND2_X1 U9361 ( .A1(n7690), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7692) );
  XOR2_X1 U9362 ( .A(n7690), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10264) );
  NAND2_X1 U9363 ( .A1(n10264), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7691) );
  NAND2_X1 U9364 ( .A1(n7692), .A2(n7691), .ZN(n7693) );
  NAND2_X1 U9365 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7693), .ZN(n7695) );
  XOR2_X1 U9366 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7693), .Z(n10263) );
  NAND2_X1 U9367 ( .A1(n10263), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7694) );
  NAND2_X1 U9368 ( .A1(n7695), .A2(n7694), .ZN(n7696) );
  NAND2_X1 U9369 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7696), .ZN(n7698) );
  XOR2_X1 U9370 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7696), .Z(n10275) );
  NAND2_X1 U9371 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10275), .ZN(n7697) );
  NAND2_X1 U9372 ( .A1(n7698), .A2(n7697), .ZN(n7699) );
  AND2_X1 U9373 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7699), .ZN(n7700) );
  XNOR2_X1 U9374 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7699), .ZN(n10273) );
  NOR2_X1 U9375 ( .A1(n10274), .A2(n10273), .ZN(n10272) );
  NOR2_X1 U9376 ( .A1(n7700), .A2(n10272), .ZN(n9976) );
  NAND2_X1 U9377 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7701) );
  OAI21_X1 U9378 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7701), .ZN(n9975) );
  NOR2_X1 U9379 ( .A1(n9976), .A2(n9975), .ZN(n9974) );
  AOI21_X1 U9380 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9974), .ZN(n9973) );
  NAND2_X1 U9381 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7702) );
  OAI21_X1 U9382 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7702), .ZN(n9972) );
  NOR2_X1 U9383 ( .A1(n9973), .A2(n9972), .ZN(n9971) );
  AOI21_X1 U9384 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9971), .ZN(n9970) );
  NOR2_X1 U9385 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7703) );
  AOI21_X1 U9386 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7703), .ZN(n9969) );
  NAND2_X1 U9387 ( .A1(n9970), .A2(n9969), .ZN(n9968) );
  OAI21_X1 U9388 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9968), .ZN(n9966) );
  NAND2_X1 U9389 ( .A1(n9967), .A2(n9966), .ZN(n9965) );
  OAI21_X1 U9390 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9965), .ZN(n9963) );
  NAND2_X1 U9391 ( .A1(n9964), .A2(n9963), .ZN(n9962) );
  OAI21_X1 U9392 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9962), .ZN(n9960) );
  NAND2_X1 U9393 ( .A1(n9961), .A2(n9960), .ZN(n9959) );
  OAI21_X1 U9394 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9959), .ZN(n9957) );
  NAND2_X1 U9395 ( .A1(n9958), .A2(n9957), .ZN(n9956) );
  OAI21_X1 U9396 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9956), .ZN(n9954) );
  NAND2_X1 U9397 ( .A1(n9955), .A2(n9954), .ZN(n9953) );
  OAI21_X1 U9398 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9953), .ZN(n10269) );
  NOR2_X1 U9399 ( .A1(n10270), .A2(n10269), .ZN(n7704) );
  NAND2_X1 U9400 ( .A1(n10270), .A2(n10269), .ZN(n10268) );
  OAI21_X1 U9401 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7704), .A(n10268), .ZN(
        n7708) );
  NOR2_X1 U9402 ( .A1(n7706), .A2(n7705), .ZN(n7707) );
  XNOR2_X1 U9403 ( .A(n7708), .B(n7707), .ZN(ADD_1071_U4) );
  INV_X1 U9404 ( .A(n7709), .ZN(n7930) );
  OAI222_X1 U9405 ( .A1(n7924), .A2(n7710), .B1(P1_U3084), .B2(n9619), .C1(
        n7920), .C2(n7930), .ZN(P1_U3326) );
  OAI211_X1 U9406 ( .C1(n7713), .C2(n7712), .A(n7711), .B(n8622), .ZN(n7719)
         );
  OAI22_X1 U9407 ( .A1(n8614), .A2(n7715), .B1(n8640), .B2(n7714), .ZN(n7716)
         );
  AOI211_X1 U9408 ( .C1(n8624), .C2(n8652), .A(n7717), .B(n7716), .ZN(n7718)
         );
  OAI211_X1 U9409 ( .C1(n7720), .C2(n8619), .A(n7719), .B(n7718), .ZN(P2_U3236) );
  INV_X1 U9410 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7726) );
  INV_X1 U9411 ( .A(n7901), .ZN(n7721) );
  OAI22_X1 U9412 ( .A1(n7722), .A2(n9927), .B1(n7721), .B2(n9925), .ZN(n7724)
         );
  AOI211_X1 U9413 ( .C1(n9931), .C2(n7725), .A(n7724), .B(n7723), .ZN(n7728)
         );
  MUX2_X1 U9414 ( .A(n7726), .B(n7728), .S(n9935), .Z(n7727) );
  INV_X1 U9415 ( .A(n7727), .ZN(P2_U3496) );
  MUX2_X1 U9416 ( .A(n5982), .B(n7728), .S(n9947), .Z(n7729) );
  INV_X1 U9417 ( .A(n7729), .ZN(P2_U3535) );
  NAND2_X1 U9418 ( .A1(n7730), .A2(n7731), .ZN(n7732) );
  XOR2_X1 U9419 ( .A(n7733), .B(n7732), .Z(n7738) );
  AND2_X1 U9420 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9715) );
  NOR2_X1 U9421 ( .A1(n7876), .A2(n9208), .ZN(n7734) );
  AOI211_X1 U9422 ( .C1(n9194), .C2(n9222), .A(n9715), .B(n7734), .ZN(n7735)
         );
  OAI21_X1 U9423 ( .B1(n9186), .B2(n7782), .A(n7735), .ZN(n7736) );
  AOI21_X1 U9424 ( .B1(n7778), .B2(n9199), .A(n7736), .ZN(n7737) );
  OAI21_X1 U9425 ( .B1(n7738), .B2(n9201), .A(n7737), .ZN(P1_U3239) );
  XOR2_X1 U9426 ( .A(n8108), .B(n7739), .Z(n9608) );
  INV_X1 U9427 ( .A(n9608), .ZN(n7755) );
  NAND2_X1 U9428 ( .A1(n7740), .A2(n8132), .ZN(n7742) );
  INV_X1 U9429 ( .A(n8108), .ZN(n7741) );
  XNOR2_X1 U9430 ( .A(n7742), .B(n7741), .ZN(n7743) );
  NAND2_X1 U9431 ( .A1(n7743), .A2(n9586), .ZN(n7745) );
  AOI22_X1 U9432 ( .A1(n9417), .A2(n9221), .B1(n9223), .B2(n9419), .ZN(n7744)
         );
  NAND2_X1 U9433 ( .A1(n7745), .A2(n7744), .ZN(n9607) );
  INV_X1 U9434 ( .A(n7751), .ZN(n9605) );
  INV_X1 U9435 ( .A(n7746), .ZN(n7767) );
  INV_X1 U9436 ( .A(n7781), .ZN(n7747) );
  OAI211_X1 U9437 ( .C1(n9605), .C2(n7767), .A(n7747), .B(n9595), .ZN(n9604)
         );
  OAI22_X1 U9438 ( .A1(n9785), .A2(n7749), .B1(n7748), .B2(n9776), .ZN(n7750)
         );
  AOI21_X1 U9439 ( .B1(n7751), .B2(n9590), .A(n7750), .ZN(n7752) );
  OAI21_X1 U9440 ( .B1(n9604), .B2(n9329), .A(n7752), .ZN(n7753) );
  AOI21_X1 U9441 ( .B1(n9607), .B2(n9785), .A(n7753), .ZN(n7754) );
  OAI21_X1 U9442 ( .B1(n7755), .B2(n9425), .A(n7754), .ZN(P1_U3277) );
  INV_X1 U9443 ( .A(n9497), .ZN(n7864) );
  AOI21_X1 U9444 ( .B1(n7758), .B2(n7730), .A(n7757), .ZN(n7759) );
  OAI21_X1 U9445 ( .B1(n4554), .B2(n7759), .A(n9204), .ZN(n7764) );
  INV_X1 U9446 ( .A(n7760), .ZN(n7861) );
  NAND2_X1 U9447 ( .A1(n9194), .A2(n9221), .ZN(n7761) );
  NAND2_X1 U9448 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9722) );
  OAI211_X1 U9449 ( .C1(n7888), .C2(n9208), .A(n7761), .B(n9722), .ZN(n7762)
         );
  AOI21_X1 U9450 ( .B1(n7861), .B2(n9211), .A(n7762), .ZN(n7763) );
  OAI211_X1 U9451 ( .C1(n7864), .C2(n9214), .A(n7764), .B(n7763), .ZN(P1_U3224) );
  NAND2_X1 U9452 ( .A1(n9581), .A2(n9580), .ZN(n9579) );
  NAND2_X1 U9453 ( .A1(n9579), .A2(n7765), .ZN(n7766) );
  XOR2_X1 U9454 ( .A(n8106), .B(n7766), .Z(n9506) );
  AOI21_X1 U9455 ( .B1(n9501), .B2(n9594), .A(n7767), .ZN(n9502) );
  INV_X1 U9456 ( .A(n9501), .ZN(n7771) );
  INV_X1 U9457 ( .A(n7768), .ZN(n7769) );
  AOI22_X1 U9458 ( .A1(n9787), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7769), .B2(
        n9588), .ZN(n7770) );
  OAI21_X1 U9459 ( .B1(n7771), .B2(n9410), .A(n7770), .ZN(n7775) );
  OAI21_X1 U9460 ( .B1(n8106), .B2(n7772), .A(n7740), .ZN(n7773) );
  AOI222_X1 U9461 ( .A1(n9586), .A2(n7773), .B1(n9224), .B2(n9419), .C1(n9222), 
        .C2(n9417), .ZN(n9504) );
  NOR2_X1 U9462 ( .A1(n9504), .A2(n9787), .ZN(n7774) );
  AOI211_X1 U9463 ( .C1(n9502), .C2(n9401), .A(n7775), .B(n7774), .ZN(n7776)
         );
  OAI21_X1 U9464 ( .B1(n9425), .B2(n9506), .A(n7776), .ZN(P1_U3278) );
  INV_X1 U9465 ( .A(n8156), .ZN(n8136) );
  OR2_X1 U9466 ( .A1(n8150), .A2(n8136), .ZN(n8012) );
  XNOR2_X1 U9467 ( .A(n7777), .B(n8012), .ZN(n7848) );
  INV_X1 U9468 ( .A(n7848), .ZN(n7787) );
  AOI22_X1 U9469 ( .A1(n7778), .A2(n9590), .B1(P1_REG2_REG_15__SCAN_IN), .B2(
        n9787), .ZN(n7786) );
  XNOR2_X1 U9470 ( .A(n7779), .B(n8012), .ZN(n7780) );
  AOI222_X1 U9471 ( .A1(n9586), .A2(n7780), .B1(n9220), .B2(n9417), .C1(n9222), 
        .C2(n9419), .ZN(n7845) );
  INV_X1 U9472 ( .A(n7845), .ZN(n7784) );
  OAI211_X1 U9473 ( .C1(n7781), .C2(n7846), .A(n7860), .B(n9595), .ZN(n7844)
         );
  OAI22_X1 U9474 ( .A1(n7844), .A2(n9349), .B1(n9776), .B2(n7782), .ZN(n7783)
         );
  OAI21_X1 U9475 ( .B1(n7784), .B2(n7783), .A(n9785), .ZN(n7785) );
  OAI211_X1 U9476 ( .C1(n7787), .C2(n9425), .A(n7786), .B(n7785), .ZN(P1_U3276) );
  INV_X1 U9477 ( .A(n8288), .ZN(n7852) );
  OAI222_X1 U9478 ( .A1(n7788), .A2(P2_U3152), .B1(n7928), .B2(n7852), .C1(
        n8289), .C2(n10258), .ZN(P2_U3329) );
  INV_X1 U9479 ( .A(n7789), .ZN(n8510) );
  OAI222_X1 U9480 ( .A1(n7924), .A2(n7790), .B1(P1_U3084), .B2(n4384), .C1(
        n7920), .C2(n8510), .ZN(P1_U3325) );
  NAND2_X1 U9481 ( .A1(n9083), .A2(n7896), .ZN(n8435) );
  OAI21_X2 U9482 ( .B1(n7791), .B2(n8428), .A(n8427), .ZN(n7792) );
  OAI21_X1 U9483 ( .B1(n8326), .B2(n7792), .A(n7810), .ZN(n7800) );
  OAI22_X1 U9484 ( .A1(n8576), .A2(n8952), .B1(n8649), .B2(n8950), .ZN(n7799)
         );
  OR2_X1 U9485 ( .A1(n7901), .A2(n8651), .ZN(n7793) );
  AND2_X1 U9486 ( .A1(n7795), .A2(n8326), .ZN(n7796) );
  OR2_X1 U9487 ( .A1(n7796), .A2(n7821), .ZN(n9087) );
  NOR2_X1 U9488 ( .A1(n9087), .A2(n7797), .ZN(n7798) );
  AOI211_X1 U9489 ( .C1(n8998), .C2(n7800), .A(n7799), .B(n7798), .ZN(n9086)
         );
  OAI22_X1 U9490 ( .A1(n8936), .A2(n7801), .B1(n8575), .B2(n8934), .ZN(n7802)
         );
  AOI21_X1 U9491 ( .B1(n9083), .B2(n8845), .A(n7802), .ZN(n7806) );
  AND2_X1 U9492 ( .A1(n7803), .A2(n9083), .ZN(n7804) );
  NOR2_X1 U9493 ( .A1(n7814), .A2(n7804), .ZN(n9084) );
  NAND2_X1 U9494 ( .A1(n9084), .A2(n9001), .ZN(n7805) );
  OAI211_X1 U9495 ( .C1(n9087), .C2(n7807), .A(n7806), .B(n7805), .ZN(n7808)
         );
  INV_X1 U9496 ( .A(n7808), .ZN(n7809) );
  OAI21_X1 U9497 ( .B1(n9086), .B2(n8956), .A(n7809), .ZN(P2_U3280) );
  AOI211_X1 U9498 ( .C1(n8436), .C2(n7811), .A(n8970), .B(n4454), .ZN(n7813)
         );
  OAI22_X1 U9499 ( .A1(n8779), .A2(n8950), .B1(n7896), .B2(n8952), .ZN(n7812)
         );
  NOR2_X1 U9500 ( .A1(n7813), .A2(n7812), .ZN(n9081) );
  INV_X1 U9501 ( .A(n7814), .ZN(n7815) );
  AOI211_X1 U9502 ( .C1(n9079), .C2(n7815), .A(n9927), .B(n8980), .ZN(n9078)
         );
  NOR2_X1 U9503 ( .A1(n7816), .A2(n8989), .ZN(n7820) );
  INV_X1 U9504 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7818) );
  OAI22_X1 U9505 ( .A1(n8936), .A2(n7818), .B1(n7817), .B2(n8934), .ZN(n7819)
         );
  AOI211_X1 U9506 ( .C1(n9078), .C2(n8977), .A(n7820), .B(n7819), .ZN(n7823)
         );
  INV_X1 U9507 ( .A(n7896), .ZN(n8650) );
  OAI21_X1 U9508 ( .B1(n4450), .B2(n8436), .A(n8777), .ZN(n9077) );
  NAND2_X1 U9509 ( .A1(n9077), .A2(n8905), .ZN(n7822) );
  OAI211_X1 U9510 ( .C1(n9081), .C2(n8956), .A(n7823), .B(n7822), .ZN(P2_U3279) );
  OAI21_X1 U9511 ( .B1(n7826), .B2(n7825), .A(n7824), .ZN(n7827) );
  NAND2_X1 U9512 ( .A1(n7827), .A2(n9204), .ZN(n7831) );
  NAND2_X1 U9513 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9740) );
  OAI21_X1 U9514 ( .B1(n7876), .B2(n9207), .A(n9740), .ZN(n7829) );
  NOR2_X1 U9515 ( .A1(n9186), .A2(n7869), .ZN(n7828) );
  AOI211_X1 U9516 ( .C1(n9183), .C2(n9397), .A(n7829), .B(n7828), .ZN(n7830)
         );
  OAI211_X1 U9517 ( .C1(n4670), .C2(n9214), .A(n7831), .B(n7830), .ZN(P1_U3226) );
  INV_X1 U9518 ( .A(n7832), .ZN(n7833) );
  AOI21_X1 U9519 ( .B1(n7835), .B2(n7834), .A(n7833), .ZN(n7843) );
  OAI21_X1 U9520 ( .B1(n8613), .B2(n8576), .A(n7836), .ZN(n7840) );
  OAI22_X1 U9521 ( .A1(n8614), .A2(n7838), .B1(n8640), .B2(n7837), .ZN(n7839)
         );
  AOI211_X1 U9522 ( .C1(n7841), .C2(n8629), .A(n7840), .B(n7839), .ZN(n7842)
         );
  OAI21_X1 U9523 ( .B1(n7843), .B2(n8643), .A(n7842), .ZN(P2_U3217) );
  INV_X1 U9524 ( .A(n9505), .ZN(n9827) );
  OAI211_X1 U9525 ( .C1(n7846), .C2(n9831), .A(n7845), .B(n7844), .ZN(n7847)
         );
  AOI21_X1 U9526 ( .B1(n7848), .B2(n9827), .A(n7847), .ZN(n7850) );
  MUX2_X1 U9527 ( .A(n5279), .B(n7850), .S(n9852), .Z(n7849) );
  INV_X1 U9528 ( .A(n7849), .ZN(P1_U3538) );
  MUX2_X1 U9529 ( .A(n5278), .B(n7850), .S(n9840), .Z(n7851) );
  INV_X1 U9530 ( .A(n7851), .ZN(P1_U3499) );
  XNOR2_X1 U9531 ( .A(n7855), .B(n8021), .ZN(n9499) );
  XNOR2_X1 U9532 ( .A(n7856), .B(n8021), .ZN(n7857) );
  OAI222_X1 U9533 ( .A1(n9577), .A2(n7888), .B1(n5559), .B2(n7858), .C1(n7857), 
        .C2(n5556), .ZN(n9495) );
  INV_X1 U9534 ( .A(n7868), .ZN(n7859) );
  AOI211_X1 U9535 ( .C1(n9497), .C2(n7860), .A(n9832), .B(n7859), .ZN(n9496)
         );
  NAND2_X1 U9536 ( .A1(n9496), .A2(n9598), .ZN(n7863) );
  AOI22_X1 U9537 ( .A1(n9787), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n7861), .B2(
        n9588), .ZN(n7862) );
  OAI211_X1 U9538 ( .C1(n7864), .C2(n9410), .A(n7863), .B(n7862), .ZN(n7865)
         );
  AOI21_X1 U9539 ( .B1(n9495), .B2(n9785), .A(n7865), .ZN(n7866) );
  OAI21_X1 U9540 ( .B1(n9499), .B2(n9425), .A(n7866), .ZN(P1_U3275) );
  XOR2_X1 U9541 ( .A(n7867), .B(n8112), .Z(n9494) );
  AOI21_X1 U9542 ( .B1(n9490), .B2(n7868), .A(n9405), .ZN(n9491) );
  INV_X1 U9543 ( .A(n7869), .ZN(n7870) );
  AOI22_X1 U9544 ( .A1(n9787), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n7870), .B2(
        n9588), .ZN(n7871) );
  OAI21_X1 U9545 ( .B1(n4670), .B2(n9410), .A(n7871), .ZN(n7880) );
  INV_X1 U9546 ( .A(n8112), .ZN(n7875) );
  INV_X1 U9547 ( .A(n7872), .ZN(n7874) );
  INV_X1 U9548 ( .A(n7873), .ZN(n9414) );
  AOI211_X1 U9549 ( .C1(n7875), .C2(n7874), .A(n5556), .B(n9414), .ZN(n7878)
         );
  OAI22_X1 U9550 ( .A1(n7876), .A2(n5559), .B1(n7909), .B2(n9577), .ZN(n7877)
         );
  NOR2_X1 U9551 ( .A1(n7878), .A2(n7877), .ZN(n9493) );
  NOR2_X1 U9552 ( .A1(n9493), .A2(n9787), .ZN(n7879) );
  AOI211_X1 U9553 ( .C1(n9491), .C2(n9401), .A(n7880), .B(n7879), .ZN(n7881)
         );
  OAI21_X1 U9554 ( .B1(n9425), .B2(n9494), .A(n7881), .ZN(P1_U3274) );
  NOR2_X1 U9555 ( .A1(n7882), .A2(n4770), .ZN(n7887) );
  AOI21_X1 U9556 ( .B1(n7885), .B2(n7884), .A(n7883), .ZN(n7886) );
  OAI21_X1 U9557 ( .B1(n7887), .B2(n7886), .A(n9204), .ZN(n7892) );
  NAND2_X1 U9558 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9750) );
  OAI21_X1 U9559 ( .B1(n7888), .B2(n9207), .A(n9750), .ZN(n7890) );
  NOR2_X1 U9560 ( .A1(n9186), .A2(n9407), .ZN(n7889) );
  AOI211_X1 U9561 ( .C1(n9183), .C2(n9418), .A(n7890), .B(n7889), .ZN(n7891)
         );
  OAI211_X1 U9562 ( .C1(n9411), .C2(n9214), .A(n7892), .B(n7891), .ZN(P1_U3236) );
  XNOR2_X1 U9563 ( .A(n7893), .B(n8570), .ZN(n7895) );
  NOR2_X1 U9564 ( .A1(n7895), .A2(n7894), .ZN(n8569) );
  AOI21_X1 U9565 ( .B1(n7895), .B2(n7894), .A(n8569), .ZN(n7903) );
  NAND2_X1 U9566 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n8684) );
  OAI21_X1 U9567 ( .B1(n8613), .B2(n7896), .A(n8684), .ZN(n7900) );
  OAI22_X1 U9568 ( .A1(n8614), .A2(n7898), .B1(n8640), .B2(n7897), .ZN(n7899)
         );
  AOI211_X1 U9569 ( .C1(n7901), .C2(n8629), .A(n7900), .B(n7899), .ZN(n7902)
         );
  OAI21_X1 U9570 ( .B1(n7903), .B2(n8643), .A(n7902), .ZN(P2_U3243) );
  OAI21_X1 U9571 ( .B1(n7906), .B2(n7905), .A(n7904), .ZN(n7907) );
  NAND2_X1 U9572 ( .A1(n7907), .A2(n9204), .ZN(n7912) );
  NAND2_X1 U9573 ( .A1(n9183), .A2(n9396), .ZN(n7908) );
  NAND2_X1 U9574 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9273) );
  OAI211_X1 U9575 ( .C1(n7909), .C2(n9207), .A(n7908), .B(n9273), .ZN(n7910)
         );
  AOI21_X1 U9576 ( .B1(n9391), .B2(n9211), .A(n7910), .ZN(n7911) );
  OAI211_X1 U9577 ( .C1(n9393), .C2(n9214), .A(n7912), .B(n7911), .ZN(P1_U3217) );
  OAI211_X1 U9578 ( .C1(n7915), .C2(n7914), .A(n7913), .B(n8622), .ZN(n7918)
         );
  INV_X1 U9579 ( .A(n8953), .ZN(n8994) );
  AND2_X1 U9580 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3152), .ZN(n8732) );
  OAI22_X1 U9581 ( .A1(n8614), .A2(n8649), .B1(n8640), .B2(n8984), .ZN(n7916)
         );
  AOI211_X1 U9582 ( .C1(n8624), .C2(n8994), .A(n8732), .B(n7916), .ZN(n7917)
         );
  OAI211_X1 U9583 ( .C1(n8990), .C2(n8619), .A(n7918), .B(n7917), .ZN(P2_U3240) );
  INV_X1 U9584 ( .A(n8293), .ZN(n7927) );
  OAI222_X1 U9585 ( .A1(n7921), .A2(n7924), .B1(n7920), .B2(n7927), .C1(
        P1_U3084), .C2(n7919), .ZN(P1_U3323) );
  OAI222_X1 U9586 ( .A1(n7924), .A2(n7923), .B1(n7920), .B2(n7922), .C1(
        P1_U3084), .C2(n8205), .ZN(P1_U3331) );
  OAI222_X1 U9587 ( .A1(n8511), .A2(n7926), .B1(n7928), .B2(n7925), .C1(
        P2_U3152), .C2(n8855), .ZN(P2_U3339) );
  INV_X1 U9588 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n10118) );
  OAI222_X1 U9589 ( .A1(n8511), .A2(n7931), .B1(n10256), .B2(n7930), .C1(n6715), .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U9590 ( .A(n7932), .ZN(n7933) );
  AOI21_X1 U9591 ( .B1(n7934), .B2(n7159), .A(n7933), .ZN(n7942) );
  NOR2_X1 U9592 ( .A1(n7935), .A2(n9208), .ZN(n7936) );
  AOI211_X1 U9593 ( .C1(n9194), .C2(n9228), .A(n7937), .B(n7936), .ZN(n7938)
         );
  OAI21_X1 U9594 ( .B1(n9186), .B2(n7939), .A(n7938), .ZN(n7940) );
  AOI21_X1 U9595 ( .B1(n9188), .B2(n9830), .A(n7940), .ZN(n7941) );
  OAI21_X1 U9596 ( .B1(n7942), .B2(n9201), .A(n7941), .ZN(P1_U3229) );
  NOR2_X1 U9597 ( .A1(n9785), .A2(n7943), .ZN(n7944) );
  NOR2_X1 U9598 ( .A1(n9787), .A2(n9428), .ZN(n9278) );
  AOI211_X1 U9599 ( .C1(n8088), .C2(n9590), .A(n7944), .B(n9278), .ZN(n7945)
         );
  OAI21_X1 U9600 ( .B1(n7946), .B2(n9281), .A(n7945), .ZN(P1_U3262) );
  XOR2_X1 U9601 ( .A(n8121), .B(n7947), .Z(n9442) );
  AOI21_X1 U9602 ( .B1(n9438), .B2(n9303), .A(n9292), .ZN(n9439) );
  AOI22_X1 U9603 ( .A1(n9137), .A2(n9588), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9787), .ZN(n7948) );
  OAI21_X1 U9604 ( .B1(n4889), .B2(n9410), .A(n7948), .ZN(n7953) );
  INV_X1 U9605 ( .A(n7949), .ZN(n7951) );
  INV_X1 U9606 ( .A(n8121), .ZN(n8236) );
  AOI211_X1 U9607 ( .C1(n7951), .C2(n8236), .A(n5556), .B(n9286), .ZN(n7952)
         );
  NAND2_X1 U9608 ( .A1(n8238), .A2(n8072), .ZN(n7967) );
  INV_X1 U9609 ( .A(n7954), .ZN(n7955) );
  NAND2_X1 U9610 ( .A1(n7955), .A2(SI_30_), .ZN(n7959) );
  NAND2_X1 U9611 ( .A1(n7957), .A2(n7956), .ZN(n7958) );
  NAND2_X1 U9612 ( .A1(n7959), .A2(n7958), .ZN(n7962) );
  MUX2_X1 U9613 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6553), .Z(n7960) );
  XNOR2_X1 U9614 ( .A(n7960), .B(SI_31_), .ZN(n7961) );
  NAND2_X1 U9615 ( .A1(n8298), .A2(n7963), .ZN(n7966) );
  OR2_X1 U9616 ( .A1(n4380), .A2(n6598), .ZN(n7965) );
  NAND2_X1 U9617 ( .A1(n7967), .A2(n9426), .ZN(n8196) );
  OR2_X1 U9618 ( .A1(n9344), .A2(n7968), .ZN(n8174) );
  AND2_X1 U9619 ( .A1(n8174), .A2(n7970), .ZN(n8048) );
  MUX2_X1 U9620 ( .A(n9340), .B(n8256), .S(n8079), .Z(n7969) );
  NAND2_X1 U9621 ( .A1(n8048), .A2(n7969), .ZN(n8052) );
  AND2_X1 U9622 ( .A1(n8061), .A2(n7970), .ZN(n8230) );
  OAI21_X1 U9623 ( .B1(n8256), .B2(n8052), .A(n8230), .ZN(n7971) );
  INV_X1 U9624 ( .A(n8079), .ZN(n8081) );
  NAND2_X1 U9625 ( .A1(n7971), .A2(n8081), .ZN(n8056) );
  NAND2_X1 U9626 ( .A1(n8167), .A2(n7972), .ZN(n8160) );
  NAND2_X1 U9627 ( .A1(n8026), .A2(n7973), .ZN(n8166) );
  MUX2_X1 U9628 ( .A(n8160), .B(n8166), .S(n8079), .Z(n7974) );
  INV_X1 U9629 ( .A(n7974), .ZN(n8025) );
  INV_X1 U9630 ( .A(n8095), .ZN(n7975) );
  NAND2_X1 U9631 ( .A1(n7976), .A2(n7975), .ZN(n7979) );
  NAND3_X1 U9632 ( .A1(n7979), .A2(n7978), .A3(n7977), .ZN(n7980) );
  NAND3_X1 U9633 ( .A1(n7980), .A2(n8153), .A3(n7991), .ZN(n7989) );
  INV_X1 U9634 ( .A(n7981), .ZN(n7987) );
  NAND2_X1 U9635 ( .A1(n7983), .A2(n7982), .ZN(n7986) );
  INV_X1 U9636 ( .A(n7984), .ZN(n7985) );
  AOI21_X1 U9637 ( .B1(n7987), .B2(n7986), .A(n7985), .ZN(n7988) );
  NAND3_X1 U9638 ( .A1(n7989), .A2(n7988), .A3(n8007), .ZN(n8002) );
  AND2_X1 U9639 ( .A1(n7991), .A2(n7990), .ZN(n8145) );
  AOI21_X1 U9640 ( .B1(n7992), .B2(n8145), .A(n8131), .ZN(n7998) );
  NAND2_X1 U9641 ( .A1(n7994), .A2(n7993), .ZN(n7997) );
  INV_X1 U9642 ( .A(n7995), .ZN(n7996) );
  OAI21_X1 U9643 ( .B1(n7998), .B2(n7997), .A(n7996), .ZN(n8000) );
  NAND3_X1 U9644 ( .A1(n8000), .A2(n7999), .A3(n8006), .ZN(n8001) );
  MUX2_X1 U9645 ( .A(n8002), .B(n8001), .S(n8081), .Z(n8011) );
  AND2_X1 U9646 ( .A1(n8007), .A2(n8003), .ZN(n8152) );
  OAI211_X1 U9647 ( .C1(n8152), .C2(n5225), .A(n8134), .B(n8132), .ZN(n8009)
         );
  NAND2_X1 U9648 ( .A1(n8006), .A2(n8005), .ZN(n8008) );
  OAI21_X1 U9649 ( .B1(n8011), .B2(n8010), .A(n4420), .ZN(n8019) );
  INV_X1 U9650 ( .A(n8012), .ZN(n8111) );
  NAND2_X1 U9651 ( .A1(n8013), .A2(n8134), .ZN(n8017) );
  NAND2_X1 U9652 ( .A1(n8015), .A2(n8014), .ZN(n8016) );
  AND2_X1 U9653 ( .A1(n8016), .A2(n8134), .ZN(n8157) );
  MUX2_X1 U9654 ( .A(n8017), .B(n8157), .S(n8079), .Z(n8018) );
  NAND3_X1 U9655 ( .A1(n8019), .A2(n8111), .A3(n8018), .ZN(n8022) );
  MUX2_X1 U9656 ( .A(n8136), .B(n8150), .S(n8079), .Z(n8020) );
  MUX2_X1 U9657 ( .A(n8149), .B(n8023), .S(n8079), .Z(n8024) );
  NAND3_X1 U9658 ( .A1(n8027), .A2(n8165), .A3(n8036), .ZN(n8032) );
  NAND3_X1 U9659 ( .A1(n8028), .A2(n8167), .A3(n8165), .ZN(n8030) );
  AND2_X1 U9660 ( .A1(n8034), .A2(n8029), .ZN(n8172) );
  NAND2_X1 U9661 ( .A1(n8030), .A2(n8172), .ZN(n8031) );
  MUX2_X1 U9662 ( .A(n8032), .B(n8031), .S(n8079), .Z(n8046) );
  INV_X1 U9663 ( .A(n8038), .ZN(n8033) );
  NAND2_X1 U9664 ( .A1(n8043), .A2(n8042), .ZN(n8035) );
  INV_X1 U9665 ( .A(n8036), .ZN(n8037) );
  NAND2_X1 U9666 ( .A1(n8042), .A2(n8037), .ZN(n8039) );
  AND2_X1 U9667 ( .A1(n8039), .A2(n8038), .ZN(n8041) );
  AND2_X1 U9668 ( .A1(n8041), .A2(n8040), .ZN(n8045) );
  INV_X1 U9669 ( .A(n8045), .ZN(n8171) );
  OR2_X1 U9670 ( .A1(n8171), .A2(n8042), .ZN(n8044) );
  NAND2_X1 U9671 ( .A1(n8046), .A2(n8045), .ZN(n8047) );
  INV_X1 U9672 ( .A(n8048), .ZN(n8050) );
  OAI21_X1 U9673 ( .B1(n8050), .B2(n8049), .A(n8052), .ZN(n8051) );
  OAI211_X1 U9674 ( .C1(n8052), .C2(n9340), .A(n8180), .B(n8174), .ZN(n8053)
         );
  NAND3_X1 U9675 ( .A1(n8056), .A2(n8055), .A3(n8054), .ZN(n8065) );
  NAND2_X1 U9676 ( .A1(n8065), .A2(n8180), .ZN(n8057) );
  AOI21_X1 U9677 ( .B1(n8057), .B2(n9307), .A(n9320), .ZN(n8060) );
  NAND2_X1 U9678 ( .A1(n8065), .A2(n8061), .ZN(n8058) );
  AOI21_X1 U9679 ( .B1(n8058), .B2(n9135), .A(n9443), .ZN(n8059) );
  NAND2_X1 U9680 ( .A1(n8061), .A2(n9320), .ZN(n8064) );
  NAND2_X1 U9681 ( .A1(n9443), .A2(n8180), .ZN(n8062) );
  AND2_X1 U9682 ( .A1(n8185), .A2(n8062), .ZN(n8063) );
  MUX2_X1 U9683 ( .A(n8064), .B(n8063), .S(n8081), .Z(n8067) );
  INV_X1 U9684 ( .A(n8065), .ZN(n8066) );
  AOI22_X1 U9685 ( .A1(n8182), .A2(n8067), .B1(n8066), .B2(n8121), .ZN(n8069)
         );
  MUX2_X1 U9686 ( .A(n8182), .B(n8185), .S(n8079), .Z(n8068) );
  MUX2_X1 U9687 ( .A(n8184), .B(n8129), .S(n8079), .Z(n8070) );
  NAND2_X1 U9688 ( .A1(n8072), .A2(n9215), .ZN(n8071) );
  NAND2_X1 U9689 ( .A1(n8088), .A2(n8071), .ZN(n8192) );
  INV_X1 U9690 ( .A(n9291), .ZN(n8189) );
  OAI21_X1 U9691 ( .B1(n8073), .B2(n8189), .A(n8196), .ZN(n8075) );
  INV_X1 U9692 ( .A(n9431), .ZN(n8077) );
  INV_X1 U9693 ( .A(n8072), .ZN(n8084) );
  OAI22_X1 U9694 ( .A1(n8073), .A2(n8077), .B1(n8241), .B2(n8192), .ZN(n8074)
         );
  MUX2_X1 U9695 ( .A(n8075), .B(n8074), .S(n8079), .Z(n8087) );
  INV_X1 U9696 ( .A(n8076), .ZN(n8078) );
  NAND3_X1 U9697 ( .A1(n8078), .A2(n8077), .A3(n8189), .ZN(n8083) );
  AND2_X1 U9698 ( .A1(n9291), .A2(n8079), .ZN(n8080) );
  AOI21_X1 U9699 ( .B1(n9431), .B2(n8081), .A(n8080), .ZN(n8082) );
  NAND4_X1 U9700 ( .A1(n8196), .A2(n8083), .A3(n8082), .A4(n8192), .ZN(n8085)
         );
  NAND2_X1 U9701 ( .A1(n8085), .A2(n8204), .ZN(n8086) );
  NAND2_X1 U9702 ( .A1(n8088), .A2(n5565), .ZN(n8089) );
  NAND2_X1 U9703 ( .A1(n8204), .A2(n8089), .ZN(n8208) );
  INV_X1 U9704 ( .A(n9362), .ZN(n8117) );
  INV_X1 U9705 ( .A(n8090), .ZN(n8094) );
  AND4_X1 U9706 ( .A1(n8094), .A2(n8093), .A3(n8092), .A4(n8091), .ZN(n8098)
         );
  NOR2_X1 U9707 ( .A1(n5620), .A2(n8095), .ZN(n8097) );
  AND4_X1 U9708 ( .A1(n8098), .A2(n5115), .A3(n8097), .A4(n8096), .ZN(n8102)
         );
  NAND4_X1 U9709 ( .A1(n8102), .A2(n8101), .A3(n8100), .A4(n8099), .ZN(n8103)
         );
  NOR2_X1 U9710 ( .A1(n9580), .A2(n8103), .ZN(n8105) );
  NAND3_X1 U9711 ( .A1(n8106), .A2(n8105), .A3(n8104), .ZN(n8107) );
  NOR2_X1 U9712 ( .A1(n8108), .A2(n8107), .ZN(n8109) );
  AND4_X1 U9713 ( .A1(n8112), .A2(n8111), .A3(n8110), .A4(n8109), .ZN(n8113)
         );
  NAND3_X1 U9714 ( .A1(n9394), .A2(n8114), .A3(n8113), .ZN(n8115) );
  NOR2_X1 U9715 ( .A1(n9379), .A2(n8115), .ZN(n8116) );
  NAND3_X1 U9716 ( .A1(n8271), .A2(n8117), .A3(n8116), .ZN(n8118) );
  NOR2_X1 U9717 ( .A1(n8260), .A2(n8118), .ZN(n8119) );
  INV_X1 U9718 ( .A(n9336), .ZN(n9334) );
  AND4_X1 U9719 ( .A1(n9309), .A2(n9323), .A3(n8119), .A4(n9334), .ZN(n8120)
         );
  AND4_X1 U9720 ( .A1(n8122), .A2(n9288), .A3(n8121), .A4(n8120), .ZN(n8123)
         );
  NAND2_X1 U9721 ( .A1(n8238), .A2(n8123), .ZN(n8124) );
  AOI21_X1 U9722 ( .B1(n8203), .B2(n8127), .A(n8128), .ZN(n8202) );
  INV_X1 U9723 ( .A(n8128), .ZN(n8200) );
  OR2_X1 U9724 ( .A1(n9431), .A2(n8189), .ZN(n8130) );
  NAND2_X1 U9725 ( .A1(n8130), .A2(n8129), .ZN(n8237) );
  INV_X1 U9726 ( .A(n8237), .ZN(n8195) );
  NOR2_X1 U9727 ( .A1(n8154), .A2(n8131), .ZN(n8133) );
  NAND4_X1 U9728 ( .A1(n8134), .A2(n8152), .A3(n8133), .A4(n8132), .ZN(n8135)
         );
  NOR4_X1 U9729 ( .A1(n8160), .A2(n8136), .A3(n8161), .A4(n8135), .ZN(n8222)
         );
  NAND2_X1 U9730 ( .A1(n8145), .A2(n8137), .ZN(n8209) );
  NAND2_X1 U9731 ( .A1(n8139), .A2(n8138), .ZN(n8220) );
  NOR2_X1 U9732 ( .A1(n8209), .A2(n8220), .ZN(n8147) );
  INV_X1 U9733 ( .A(n8218), .ZN(n8141) );
  NOR2_X1 U9734 ( .A1(n4660), .A2(n8141), .ZN(n8144) );
  INV_X1 U9735 ( .A(n8142), .ZN(n8143) );
  OAI21_X1 U9736 ( .B1(n8144), .B2(n8143), .A(n8219), .ZN(n8146) );
  AOI22_X1 U9737 ( .A1(n8148), .A2(n8147), .B1(n8146), .B2(n8145), .ZN(n8164)
         );
  INV_X1 U9738 ( .A(n8149), .ZN(n8151) );
  NOR2_X1 U9739 ( .A1(n8151), .A2(n8150), .ZN(n8163) );
  INV_X1 U9740 ( .A(n8152), .ZN(n8155) );
  NOR3_X1 U9741 ( .A1(n8155), .A2(n8154), .A3(n8153), .ZN(n8158) );
  OAI211_X1 U9742 ( .C1(n8159), .C2(n8158), .A(n8157), .B(n8156), .ZN(n8162)
         );
  AOI211_X1 U9743 ( .C1(n8163), .C2(n8162), .A(n8161), .B(n8160), .ZN(n8229)
         );
  AOI21_X1 U9744 ( .B1(n8222), .B2(n8164), .A(n8229), .ZN(n8179) );
  NOR2_X1 U9745 ( .A1(n8171), .A2(n4648), .ZN(n8168) );
  NAND2_X1 U9746 ( .A1(n8178), .A2(n8168), .ZN(n8226) );
  NAND3_X1 U9747 ( .A1(n8168), .A2(n8167), .A3(n8166), .ZN(n8169) );
  OAI211_X1 U9748 ( .C1(n8172), .C2(n8171), .A(n8170), .B(n8169), .ZN(n8177)
         );
  INV_X1 U9749 ( .A(n8173), .ZN(n8176) );
  INV_X1 U9750 ( .A(n8174), .ZN(n8175) );
  OAI21_X1 U9751 ( .B1(n8179), .B2(n8226), .A(n8233), .ZN(n8183) );
  NAND2_X1 U9752 ( .A1(n8181), .A2(n8180), .ZN(n8234) );
  INV_X1 U9753 ( .A(n8182), .ZN(n9285) );
  AOI211_X1 U9754 ( .C1(n8230), .C2(n8183), .A(n8234), .B(n9285), .ZN(n8194)
         );
  OAI211_X1 U9755 ( .C1(n9285), .C2(n8186), .A(n8185), .B(n8184), .ZN(n8187)
         );
  INV_X1 U9756 ( .A(n8187), .ZN(n8188) );
  OR2_X1 U9757 ( .A1(n8237), .A2(n8188), .ZN(n8191) );
  NAND2_X1 U9758 ( .A1(n9431), .A2(n8189), .ZN(n8190) );
  NAND2_X1 U9759 ( .A1(n8191), .A2(n8190), .ZN(n8239) );
  INV_X1 U9760 ( .A(n8192), .ZN(n8193) );
  AOI211_X1 U9761 ( .C1(n8195), .C2(n8194), .A(n8239), .B(n8193), .ZN(n8198)
         );
  INV_X1 U9762 ( .A(n8196), .ZN(n8197) );
  OAI211_X1 U9763 ( .C1(n8198), .C2(n8197), .A(n5652), .B(n8204), .ZN(n8199)
         );
  NAND2_X1 U9764 ( .A1(n8200), .A2(n8199), .ZN(n8201) );
  INV_X1 U9765 ( .A(n8203), .ZN(n8206) );
  NAND4_X1 U9766 ( .A1(n8206), .A2(n8205), .A3(n8204), .A4(n5652), .ZN(n8207)
         );
  NAND2_X1 U9767 ( .A1(n8207), .A2(n5611), .ZN(n8247) );
  INV_X1 U9768 ( .A(n8208), .ZN(n8243) );
  INV_X1 U9769 ( .A(n8209), .ZN(n8225) );
  INV_X1 U9770 ( .A(n7199), .ZN(n8215) );
  NAND2_X1 U9771 ( .A1(n9235), .A2(n8210), .ZN(n8211) );
  OAI211_X1 U9772 ( .C1(n8212), .C2(n6259), .A(n5652), .B(n8211), .ZN(n8213)
         );
  NAND3_X1 U9773 ( .A1(n8215), .A2(n8214), .A3(n8213), .ZN(n8217) );
  AOI21_X1 U9774 ( .B1(n8217), .B2(n8216), .A(n4660), .ZN(n8221) );
  OAI211_X1 U9775 ( .C1(n8221), .C2(n8220), .A(n8219), .B(n8218), .ZN(n8224)
         );
  INV_X1 U9776 ( .A(n8222), .ZN(n8223) );
  AOI21_X1 U9777 ( .B1(n8225), .B2(n8224), .A(n8223), .ZN(n8228) );
  INV_X1 U9778 ( .A(n8226), .ZN(n8227) );
  OAI21_X1 U9779 ( .B1(n8229), .B2(n8228), .A(n8227), .ZN(n8232) );
  INV_X1 U9780 ( .A(n8230), .ZN(n8231) );
  AOI21_X1 U9781 ( .B1(n8233), .B2(n8232), .A(n8231), .ZN(n8235) );
  NOR4_X1 U9782 ( .A1(n8237), .A2(n8236), .A3(n8235), .A4(n8234), .ZN(n8240)
         );
  OAI21_X1 U9783 ( .B1(n8240), .B2(n8239), .A(n8238), .ZN(n8242) );
  AOI21_X1 U9784 ( .B1(n8243), .B2(n8242), .A(n8241), .ZN(n8244) );
  XNOR2_X1 U9785 ( .A(n8244), .B(n9349), .ZN(n8245) );
  NAND2_X1 U9786 ( .A1(n8245), .A2(n5651), .ZN(n8246) );
  NAND2_X1 U9787 ( .A1(n8249), .A2(n8248), .ZN(n8250) );
  OAI211_X1 U9788 ( .C1(n5653), .C2(n8252), .A(n8250), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8251) );
  XOR2_X1 U9789 ( .A(n8260), .B(n8253), .Z(n9464) );
  INV_X1 U9790 ( .A(n8267), .ZN(n8254) );
  AOI21_X1 U9791 ( .B1(n9460), .B2(n8254), .A(n4674), .ZN(n9461) );
  AOI22_X1 U9792 ( .A1(P1_REG2_REG_23__SCAN_IN), .A2(n9787), .B1(n9148), .B2(
        n9588), .ZN(n8255) );
  OAI21_X1 U9793 ( .B1(n8256), .B2(n9410), .A(n8255), .ZN(n8264) );
  AND2_X1 U9794 ( .A1(n9321), .A2(n9417), .ZN(n8262) );
  INV_X1 U9795 ( .A(n8258), .ZN(n8259) );
  AOI211_X1 U9796 ( .C1(n8260), .C2(n8257), .A(n5556), .B(n8259), .ZN(n8261)
         );
  AOI211_X1 U9797 ( .C1(n9419), .C2(n9366), .A(n8262), .B(n8261), .ZN(n9463)
         );
  NOR2_X1 U9798 ( .A1(n9463), .A2(n9787), .ZN(n8263) );
  AOI211_X1 U9799 ( .C1(n9461), .C2(n9401), .A(n8264), .B(n8263), .ZN(n8265)
         );
  OAI21_X1 U9800 ( .B1(n9464), .B2(n9425), .A(n8265), .ZN(P1_U3268) );
  XOR2_X1 U9801 ( .A(n8266), .B(n8271), .Z(n9469) );
  INV_X1 U9802 ( .A(n9357), .ZN(n8268) );
  AOI21_X1 U9803 ( .B1(n9465), .B2(n8268), .A(n8267), .ZN(n9466) );
  AOI22_X1 U9804 ( .A1(n9787), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9195), .B2(
        n9588), .ZN(n8269) );
  OAI21_X1 U9805 ( .B1(n8270), .B2(n9410), .A(n8269), .ZN(n8275) );
  XNOR2_X1 U9806 ( .A(n8272), .B(n8271), .ZN(n8273) );
  AOI222_X1 U9807 ( .A1(n9586), .A2(n8273), .B1(n9218), .B2(n9417), .C1(n9219), 
        .C2(n9419), .ZN(n9468) );
  NOR2_X1 U9808 ( .A1(n9468), .A2(n9787), .ZN(n8274) );
  AOI211_X1 U9809 ( .C1(n9466), .C2(n9401), .A(n8275), .B(n8274), .ZN(n8276)
         );
  OAI21_X1 U9810 ( .B1(n9469), .B2(n9425), .A(n8276), .ZN(P1_U3269) );
  OAI222_X1 U9811 ( .A1(n8511), .A2(n8278), .B1(n10256), .B2(n8277), .C1(n6216), .C2(P2_U3152), .ZN(P2_U3338) );
  NOR2_X1 U9812 ( .A1(n9079), .A2(n8649), .ZN(n8437) );
  NOR2_X1 U9813 ( .A1(n8992), .A2(n8440), .ZN(n8969) );
  OR2_X1 U9814 ( .A1(n9068), .A2(n8953), .ZN(n8442) );
  NAND2_X1 U9815 ( .A1(n9068), .A2(n8953), .ZN(n8947) );
  NAND2_X1 U9816 ( .A1(n8442), .A2(n8947), .ZN(n8967) );
  INV_X1 U9817 ( .A(n8967), .ZN(n8280) );
  INV_X1 U9818 ( .A(n8779), .ZN(n8778) );
  INV_X1 U9819 ( .A(n8968), .ZN(n8279) );
  NAND2_X1 U9820 ( .A1(n8280), .A2(n8279), .ZN(n8281) );
  OR2_X2 U9821 ( .A1(n8969), .A2(n8281), .ZN(n8971) );
  NAND2_X1 U9822 ( .A1(n9062), .A2(n8648), .ZN(n8449) );
  XNOR2_X1 U9823 ( .A(n9057), .B(n8951), .ZN(n8930) );
  NAND2_X1 U9824 ( .A1(n9057), .A2(n8951), .ZN(n8451) );
  NAND2_X1 U9825 ( .A1(n9052), .A2(n8786), .ZN(n8450) );
  INV_X1 U9826 ( .A(n8448), .ZN(n8283) );
  NOR2_X2 U9827 ( .A1(n8917), .A2(n8283), .ZN(n8892) );
  INV_X1 U9828 ( .A(n8647), .ZN(n8920) );
  NAND2_X1 U9829 ( .A1(n9045), .A2(n8920), .ZN(n8458) );
  NAND2_X1 U9830 ( .A1(n8880), .A2(n8893), .ZN(n8343) );
  NAND2_X1 U9831 ( .A1(n9040), .A2(n8521), .ZN(n8462) );
  NAND2_X1 U9832 ( .A1(n8343), .A2(n8462), .ZN(n8881) );
  NAND2_X1 U9833 ( .A1(n8885), .A2(n8343), .ZN(n8870) );
  NAND2_X1 U9834 ( .A1(n9037), .A2(n8883), .ZN(n8464) );
  NAND2_X1 U9835 ( .A1(n8870), .A2(n8871), .ZN(n8869) );
  NAND2_X1 U9836 ( .A1(n8869), .A2(n4947), .ZN(n8832) );
  INV_X1 U9837 ( .A(n8646), .ZN(n8817) );
  NAND2_X1 U9838 ( .A1(n8832), .A2(n8285), .ZN(n8831) );
  INV_X1 U9839 ( .A(n8286), .ZN(n8470) );
  NAND2_X1 U9840 ( .A1(n8831), .A2(n8470), .ZN(n8813) );
  NAND2_X1 U9841 ( .A1(n8812), .A2(n8795), .ZN(n8287) );
  NAND2_X1 U9842 ( .A1(n8288), .A2(n8299), .ZN(n8291) );
  OR2_X1 U9843 ( .A1(n8300), .A2(n8289), .ZN(n8290) );
  NOR2_X1 U9844 ( .A1(n8804), .A2(n8816), .ZN(n8481) );
  NAND2_X1 U9845 ( .A1(n8804), .A2(n8816), .ZN(n8479) );
  NAND2_X1 U9846 ( .A1(n8292), .A2(n8479), .ZN(n8297) );
  NAND2_X1 U9847 ( .A1(n8293), .A2(n8299), .ZN(n8295) );
  OR2_X1 U9848 ( .A1(n8300), .A2(n10118), .ZN(n8294) );
  OR2_X1 U9849 ( .A1(n8768), .A2(n8774), .ZN(n8477) );
  NOR2_X1 U9850 ( .A1(n8302), .A2(n8338), .ZN(n8296) );
  AOI21_X1 U9851 ( .B1(n8297), .B2(n8477), .A(n8296), .ZN(n8304) );
  NOR2_X1 U9852 ( .A1(n8297), .A2(n8768), .ZN(n8303) );
  OR2_X1 U9853 ( .A1(n8300), .A2(n6604), .ZN(n8301) );
  INV_X1 U9854 ( .A(n8302), .ZN(n8764) );
  NAND2_X1 U9855 ( .A1(n8768), .A2(n8774), .ZN(n8478) );
  OAI21_X1 U9856 ( .B1(n8304), .B2(n8303), .A(n8485), .ZN(n8305) );
  NAND2_X1 U9857 ( .A1(n8305), .A2(n8489), .ZN(n8306) );
  XNOR2_X1 U9858 ( .A(n8306), .B(n8855), .ZN(n8495) );
  NOR2_X1 U9859 ( .A1(n8504), .A2(n8307), .ZN(n8494) );
  INV_X1 U9860 ( .A(n8337), .ZN(n8308) );
  NAND2_X1 U9861 ( .A1(n8489), .A2(n8477), .ZN(n8486) );
  INV_X1 U9862 ( .A(n8486), .ZN(n8335) );
  INV_X1 U9863 ( .A(n8481), .ZN(n8309) );
  INV_X1 U9864 ( .A(n8797), .ZN(n8333) );
  INV_X1 U9865 ( .A(n8833), .ZN(n8792) );
  NOR2_X1 U9866 ( .A1(n8968), .A2(n8440), .ZN(n8991) );
  NAND2_X1 U9867 ( .A1(n8352), .A2(n8310), .ZN(n8358) );
  INV_X1 U9868 ( .A(n8311), .ZN(n8312) );
  NAND2_X1 U9869 ( .A1(n8347), .A2(n8312), .ZN(n8344) );
  INV_X1 U9870 ( .A(n8313), .ZN(n8368) );
  NOR4_X1 U9871 ( .A1(n8358), .A2(n8344), .A3(n8314), .A4(n8368), .ZN(n8318)
         );
  NAND2_X1 U9872 ( .A1(n8360), .A2(n8315), .ZN(n8353) );
  NOR3_X1 U9873 ( .A1(n7086), .A2(n8353), .A3(n6216), .ZN(n8316) );
  NAND4_X1 U9874 ( .A1(n8318), .A2(n8317), .A3(n9875), .A4(n8316), .ZN(n8322)
         );
  INV_X1 U9875 ( .A(n8319), .ZN(n8320) );
  NOR4_X1 U9876 ( .A1(n8322), .A2(n8321), .A3(n8320), .A4(n8381), .ZN(n8325)
         );
  NAND4_X1 U9877 ( .A1(n8325), .A2(n4827), .A3(n8324), .A4(n8323), .ZN(n8328)
         );
  INV_X1 U9878 ( .A(n8326), .ZN(n8430) );
  INV_X1 U9879 ( .A(n8327), .ZN(n8417) );
  NOR4_X1 U9880 ( .A1(n8328), .A2(n8430), .A3(n8424), .A4(n8417), .ZN(n8329)
         );
  NAND4_X1 U9881 ( .A1(n8280), .A2(n8991), .A3(n8329), .A4(n4686), .ZN(n8330)
         );
  NOR4_X1 U9882 ( .A1(n8919), .A2(n8930), .A3(n8940), .A4(n8330), .ZN(n8331)
         );
  NAND4_X1 U9883 ( .A1(n8871), .A2(n8284), .A3(n8331), .A4(n8891), .ZN(n8332)
         );
  NOR4_X1 U9884 ( .A1(n8333), .A2(n8792), .A3(n8788), .A4(n8332), .ZN(n8334)
         );
  NAND4_X1 U9885 ( .A1(n8485), .A2(n8335), .A3(n8334), .A4(n8808), .ZN(n8336)
         );
  XOR2_X1 U9886 ( .A(n8855), .B(n8336), .Z(n8339) );
  AOI22_X1 U9887 ( .A1(n8339), .A2(n8338), .B1(n8337), .B2(n6216), .ZN(n8493)
         );
  AND2_X1 U9888 ( .A1(n8340), .A2(n8351), .ZN(n8341) );
  INV_X1 U9889 ( .A(n9045), .ZN(n8898) );
  INV_X1 U9890 ( .A(n8343), .ZN(n8461) );
  MUX2_X1 U9891 ( .A(n8344), .B(n8368), .S(n4382), .Z(n8355) );
  INV_X1 U9892 ( .A(n8344), .ZN(n8346) );
  AOI22_X1 U9893 ( .A1(n8355), .A2(n8347), .B1(n8346), .B2(n8345), .ZN(n8349)
         );
  INV_X1 U9894 ( .A(n8374), .ZN(n8348) );
  OAI21_X1 U9895 ( .B1(n8349), .B2(n8348), .A(n4382), .ZN(n8365) );
  AOI21_X1 U9896 ( .B1(n8351), .B2(n8359), .A(n8350), .ZN(n8354) );
  OAI211_X1 U9897 ( .C1(n8354), .C2(n8353), .A(n8352), .B(n4382), .ZN(n8357)
         );
  INV_X1 U9898 ( .A(n8355), .ZN(n8371) );
  NAND3_X1 U9899 ( .A1(n8357), .A2(n8371), .A3(n8356), .ZN(n8364) );
  AOI21_X1 U9900 ( .B1(n8360), .B2(n8359), .A(n8358), .ZN(n8362) );
  INV_X1 U9901 ( .A(n8315), .ZN(n8361) );
  NOR3_X1 U9902 ( .A1(n8362), .A2(n8361), .A3(n4382), .ZN(n8363) );
  AOI21_X1 U9903 ( .B1(n8365), .B2(n8364), .A(n8363), .ZN(n8378) );
  INV_X1 U9904 ( .A(n8366), .ZN(n8370) );
  INV_X1 U9905 ( .A(n8367), .ZN(n8369) );
  OAI22_X1 U9906 ( .A1(n8371), .A2(n8370), .B1(n8369), .B2(n8368), .ZN(n8372)
         );
  AOI21_X1 U9907 ( .B1(n8372), .B2(n8373), .A(n4382), .ZN(n8377) );
  MUX2_X1 U9908 ( .A(n8374), .B(n8373), .S(n4382), .Z(n8375) );
  OAI211_X1 U9909 ( .C1(n8378), .C2(n8377), .A(n8376), .B(n8375), .ZN(n8390)
         );
  MUX2_X1 U9910 ( .A(n7088), .B(n8380), .S(n4382), .Z(n8382) );
  NOR2_X1 U9911 ( .A1(n8382), .A2(n8381), .ZN(n8389) );
  INV_X1 U9912 ( .A(n8394), .ZN(n8388) );
  INV_X1 U9913 ( .A(n8383), .ZN(n8386) );
  NAND2_X1 U9914 ( .A1(n8391), .A2(n8384), .ZN(n8385) );
  MUX2_X1 U9915 ( .A(n8386), .B(n8385), .S(n4382), .Z(n8387) );
  AOI211_X1 U9916 ( .C1(n8390), .C2(n8389), .A(n8388), .B(n8387), .ZN(n8399)
         );
  INV_X1 U9917 ( .A(n8396), .ZN(n8393) );
  INV_X1 U9918 ( .A(n8391), .ZN(n8392) );
  NOR3_X1 U9919 ( .A1(n8399), .A2(n8393), .A3(n8392), .ZN(n8401) );
  NAND2_X1 U9920 ( .A1(n8395), .A2(n8394), .ZN(n8398) );
  OAI211_X1 U9921 ( .C1(n8399), .C2(n8398), .A(n8397), .B(n8396), .ZN(n8400)
         );
  MUX2_X1 U9922 ( .A(n8401), .B(n8400), .S(n4382), .Z(n8404) );
  AOI21_X1 U9923 ( .B1(n8406), .B2(n8402), .A(n4382), .ZN(n8403) );
  NOR2_X1 U9924 ( .A1(n8404), .A2(n8403), .ZN(n8413) );
  INV_X1 U9925 ( .A(n8405), .ZN(n8408) );
  NAND2_X1 U9926 ( .A1(n8410), .A2(n8406), .ZN(n8407) );
  MUX2_X1 U9927 ( .A(n8408), .B(n8407), .S(n4382), .Z(n8412) );
  MUX2_X1 U9928 ( .A(n8410), .B(n8409), .S(n4382), .Z(n8411) );
  OAI21_X1 U9929 ( .B1(n8413), .B2(n8412), .A(n8411), .ZN(n8419) );
  INV_X1 U9930 ( .A(n8414), .ZN(n8415) );
  MUX2_X1 U9931 ( .A(n8416), .B(n8415), .S(n4382), .Z(n8418) );
  AOI211_X1 U9932 ( .C1(n8419), .C2(n4827), .A(n8418), .B(n8417), .ZN(n8426)
         );
  INV_X1 U9933 ( .A(n8420), .ZN(n8423) );
  INV_X1 U9934 ( .A(n8421), .ZN(n8422) );
  MUX2_X1 U9935 ( .A(n8423), .B(n8422), .S(n4382), .Z(n8425) );
  NOR3_X1 U9936 ( .A1(n8426), .A2(n8425), .A3(n8424), .ZN(n8432) );
  INV_X1 U9937 ( .A(n8427), .ZN(n8429) );
  MUX2_X1 U9938 ( .A(n8429), .B(n8428), .S(n4382), .Z(n8431) );
  INV_X1 U9939 ( .A(n8433), .ZN(n8434) );
  INV_X1 U9940 ( .A(n8440), .ZN(n8438) );
  OAI211_X1 U9941 ( .C1(n8441), .C2(n8968), .A(n8438), .B(n8947), .ZN(n8439)
         );
  NAND3_X1 U9942 ( .A1(n8439), .A2(n8453), .A3(n8442), .ZN(n8446) );
  NOR2_X1 U9943 ( .A1(n8441), .A2(n8440), .ZN(n8444) );
  INV_X1 U9944 ( .A(n8442), .ZN(n8443) );
  OAI211_X1 U9945 ( .C1(n8444), .C2(n8443), .A(n8449), .B(n8947), .ZN(n8445)
         );
  MUX2_X1 U9946 ( .A(n8446), .B(n8445), .S(n4382), .Z(n8457) );
  OR2_X1 U9947 ( .A1(n9057), .A2(n8951), .ZN(n8447) );
  NAND2_X1 U9948 ( .A1(n8448), .A2(n8447), .ZN(n8454) );
  AOI21_X1 U9949 ( .B1(n8457), .B2(n8449), .A(n8454), .ZN(n8452) );
  OAI21_X1 U9950 ( .B1(n8454), .B2(n8451), .A(n8450), .ZN(n8455) );
  NOR2_X1 U9951 ( .A1(n8454), .A2(n4839), .ZN(n8456) );
  AOI21_X1 U9952 ( .B1(n8457), .B2(n8456), .A(n8455), .ZN(n8459) );
  INV_X1 U9953 ( .A(n8462), .ZN(n8460) );
  OAI211_X1 U9954 ( .C1(n8846), .C2(n4382), .A(n8463), .B(n8467), .ZN(n8466)
         );
  NAND2_X1 U9955 ( .A1(n8834), .A2(n8464), .ZN(n8465) );
  AOI22_X1 U9956 ( .A1(n8466), .A2(n8834), .B1(n4382), .B2(n8465), .ZN(n8473)
         );
  OAI21_X1 U9957 ( .B1(n4385), .B2(n8467), .A(n8833), .ZN(n8472) );
  INV_X1 U9958 ( .A(n8468), .ZN(n8469) );
  MUX2_X1 U9959 ( .A(n8470), .B(n8469), .S(n4382), .Z(n8471) );
  OAI211_X1 U9960 ( .C1(n8473), .C2(n8472), .A(n8808), .B(n8471), .ZN(n8476)
         );
  NAND3_X1 U9961 ( .A1(n8812), .A2(n8795), .A3(n4382), .ZN(n8475) );
  INV_X1 U9962 ( .A(n8795), .ZN(n8838) );
  NAND3_X1 U9963 ( .A1(n9020), .A2(n8838), .A3(n4385), .ZN(n8474) );
  INV_X1 U9964 ( .A(n8477), .ZN(n8484) );
  INV_X1 U9965 ( .A(n8478), .ZN(n8483) );
  INV_X1 U9966 ( .A(n8479), .ZN(n8480) );
  MUX2_X1 U9967 ( .A(n8481), .B(n8480), .S(n4382), .Z(n8482) );
  INV_X1 U9968 ( .A(n8485), .ZN(n8487) );
  MUX2_X1 U9969 ( .A(n8487), .B(n8486), .S(n4382), .Z(n8488) );
  INV_X1 U9970 ( .A(n8489), .ZN(n8492) );
  INV_X1 U9971 ( .A(n8490), .ZN(n8491) );
  NAND4_X1 U9972 ( .A1(n6226), .A2(n8498), .A3(n8497), .A4(n8995), .ZN(n8499)
         );
  OAI211_X1 U9973 ( .C1(n8501), .C2(n8500), .A(n8499), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8502) );
  NAND2_X1 U9974 ( .A1(n8503), .A2(n8502), .ZN(P2_U3244) );
  OAI21_X1 U9975 ( .B1(n7115), .B2(n8504), .A(n9872), .ZN(n8505) );
  NAND3_X1 U9976 ( .A1(n8506), .A2(n8622), .A3(n8505), .ZN(n8509) );
  AOI22_X1 U9977 ( .A1(n8629), .A2(n8507), .B1(n8549), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n8508) );
  OAI211_X1 U9978 ( .C1(n6832), .C2(n8613), .A(n8509), .B(n8508), .ZN(P2_U3234) );
  OAI222_X1 U9979 ( .A1(n8511), .A2(n10188), .B1(n10256), .B2(n8510), .C1(
        n6233), .C2(P2_U3152), .ZN(P2_U3330) );
  XNOR2_X1 U9980 ( .A(n8512), .B(n8513), .ZN(n8518) );
  OAI22_X1 U9981 ( .A1(n8613), .A2(n8838), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8514), .ZN(n8516) );
  OAI22_X1 U9982 ( .A1(n8614), .A2(n8837), .B1(n8640), .B2(n8827), .ZN(n8515)
         );
  AOI211_X1 U9983 ( .C1(n9025), .C2(n8629), .A(n8516), .B(n8515), .ZN(n8517)
         );
  OAI21_X1 U9984 ( .B1(n8518), .B2(n8643), .A(n8517), .ZN(P2_U3216) );
  INV_X1 U9985 ( .A(n8519), .ZN(n8593) );
  XNOR2_X1 U9986 ( .A(n8593), .B(n8592), .ZN(n8525) );
  OAI22_X1 U9987 ( .A1(n8613), .A2(n8521), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8520), .ZN(n8523) );
  OAI22_X1 U9988 ( .A1(n8614), .A2(n8786), .B1(n8640), .B2(n8899), .ZN(n8522)
         );
  AOI211_X1 U9989 ( .C1(n9045), .C2(n8629), .A(n8523), .B(n8522), .ZN(n8524)
         );
  OAI21_X1 U9990 ( .B1(n8525), .B2(n8643), .A(n8524), .ZN(P2_U3218) );
  NAND2_X1 U9991 ( .A1(n8527), .A2(n8526), .ZN(n8529) );
  XOR2_X1 U9992 ( .A(n8529), .B(n8528), .Z(n8533) );
  OAI22_X1 U9993 ( .A1(n8779), .A2(n8952), .B1(n8648), .B2(n8950), .ZN(n8973)
         );
  AOI22_X1 U9994 ( .A1(n8973), .A2(n8638), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n8530) );
  OAI21_X1 U9995 ( .B1(n8963), .B2(n8640), .A(n8530), .ZN(n8531) );
  AOI21_X1 U9996 ( .B1(n9068), .B2(n8629), .A(n8531), .ZN(n8532) );
  OAI21_X1 U9997 ( .B1(n8533), .B2(n8643), .A(n8532), .ZN(P2_U3221) );
  XOR2_X1 U9998 ( .A(n8535), .B(n8534), .Z(n8536) );
  NAND2_X1 U9999 ( .A1(n8536), .A2(n8622), .ZN(n8544) );
  AOI22_X1 U10000 ( .A1(n8537), .A2(n8638), .B1(P2_REG3_REG_8__SCAN_IN), .B2(
        P2_U3152), .ZN(n8543) );
  INV_X1 U10001 ( .A(n8538), .ZN(n8539) );
  NAND2_X1 U10002 ( .A1(n8627), .A2(n8539), .ZN(n8542) );
  NAND2_X1 U10003 ( .A1(n8629), .A2(n8540), .ZN(n8541) );
  NAND4_X1 U10004 ( .A1(n8544), .A2(n8543), .A3(n8542), .A4(n8541), .ZN(
        P2_U3223) );
  OAI21_X1 U10005 ( .B1(n8547), .B2(n8546), .A(n8545), .ZN(n8548) );
  NAND2_X1 U10006 ( .A1(n8548), .A2(n8622), .ZN(n8553) );
  AOI22_X1 U10007 ( .A1(n8629), .A2(n8550), .B1(n8549), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n8552) );
  AOI22_X1 U10008 ( .A1(n8628), .A2(n8666), .B1(n8624), .B2(n8664), .ZN(n8551)
         );
  NAND3_X1 U10009 ( .A1(n8553), .A2(n8552), .A3(n8551), .ZN(P2_U3224) );
  XNOR2_X1 U10010 ( .A(n8554), .B(n8555), .ZN(n8559) );
  OAI22_X1 U10011 ( .A1(n8648), .A2(n8952), .B1(n8786), .B2(n8950), .ZN(n8932)
         );
  AOI22_X1 U10012 ( .A1(n8932), .A2(n8638), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8556) );
  OAI21_X1 U10013 ( .B1(n8935), .B2(n8640), .A(n8556), .ZN(n8557) );
  AOI21_X1 U10014 ( .B1(n9057), .B2(n8629), .A(n8557), .ZN(n8558) );
  OAI21_X1 U10015 ( .B1(n8559), .B2(n8643), .A(n8558), .ZN(P2_U3225) );
  XNOR2_X1 U10016 ( .A(n8560), .B(n8561), .ZN(n8568) );
  OR2_X1 U10017 ( .A1(n8837), .A2(n8950), .ZN(n8563) );
  NAND2_X1 U10018 ( .A1(n8893), .A2(n8995), .ZN(n8562) );
  AND2_X1 U10019 ( .A1(n8563), .A2(n8562), .ZN(n8872) );
  INV_X1 U10020 ( .A(n8872), .ZN(n8564) );
  AOI22_X1 U10021 ( .A1(n8564), .A2(n8638), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8565) );
  OAI21_X1 U10022 ( .B1(n8865), .B2(n8640), .A(n8565), .ZN(n8566) );
  AOI21_X1 U10023 ( .B1(n9037), .B2(n8629), .A(n8566), .ZN(n8567) );
  OAI21_X1 U10024 ( .B1(n8568), .B2(n8643), .A(n8567), .ZN(P2_U3227) );
  AOI21_X1 U10025 ( .B1(n8570), .B2(n7893), .A(n8569), .ZN(n8574) );
  XNOR2_X1 U10026 ( .A(n8572), .B(n8571), .ZN(n8573) );
  XNOR2_X1 U10027 ( .A(n8574), .B(n8573), .ZN(n8580) );
  NAND2_X1 U10028 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8706) );
  OAI21_X1 U10029 ( .B1(n8613), .B2(n8649), .A(n8706), .ZN(n8578) );
  OAI22_X1 U10030 ( .A1(n8614), .A2(n8576), .B1(n8640), .B2(n8575), .ZN(n8577)
         );
  AOI211_X1 U10031 ( .C1(n9083), .C2(n8629), .A(n8578), .B(n8577), .ZN(n8579)
         );
  OAI21_X1 U10032 ( .B1(n8580), .B2(n8643), .A(n8579), .ZN(P2_U3228) );
  XOR2_X1 U10033 ( .A(n8582), .B(n8581), .Z(n8583) );
  NAND2_X1 U10034 ( .A1(n8583), .A2(n8622), .ZN(n8590) );
  AOI22_X1 U10035 ( .A1(n8584), .A2(n8638), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n8589) );
  NAND2_X1 U10036 ( .A1(n8627), .A2(n8585), .ZN(n8588) );
  NAND2_X1 U10037 ( .A1(n8629), .A2(n8586), .ZN(n8587) );
  NAND4_X1 U10038 ( .A1(n8590), .A2(n8589), .A3(n8588), .A4(n8587), .ZN(
        P2_U3229) );
  OAI21_X1 U10039 ( .B1(n8593), .B2(n8592), .A(n8591), .ZN(n8597) );
  XNOR2_X1 U10040 ( .A(n8595), .B(n8594), .ZN(n8596) );
  XNOR2_X1 U10041 ( .A(n8597), .B(n8596), .ZN(n8602) );
  OAI22_X1 U10042 ( .A1(n8613), .A2(n8883), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8598), .ZN(n8600) );
  OAI22_X1 U10043 ( .A1(n8614), .A2(n8920), .B1(n8640), .B2(n8877), .ZN(n8599)
         );
  AOI211_X1 U10044 ( .C1(n9040), .C2(n8629), .A(n8600), .B(n8599), .ZN(n8601)
         );
  OAI21_X1 U10045 ( .B1(n8602), .B2(n8643), .A(n8601), .ZN(P2_U3231) );
  XNOR2_X1 U10046 ( .A(n8603), .B(n8604), .ZN(n8608) );
  INV_X1 U10047 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10211) );
  OAI22_X1 U10048 ( .A1(n8613), .A2(n8951), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10211), .ZN(n8606) );
  OAI22_X1 U10049 ( .A1(n8614), .A2(n8953), .B1(n8640), .B2(n8942), .ZN(n8605)
         );
  AOI211_X1 U10050 ( .C1(n9062), .C2(n8629), .A(n8606), .B(n8605), .ZN(n8607)
         );
  OAI21_X1 U10051 ( .B1(n8608), .B2(n8643), .A(n8607), .ZN(P2_U3235) );
  OAI21_X1 U10052 ( .B1(n8611), .B2(n8610), .A(n8609), .ZN(n8612) );
  NAND2_X1 U10053 ( .A1(n8612), .A2(n8622), .ZN(n8618) );
  NOR2_X1 U10054 ( .A1(n8613), .A2(n8920), .ZN(n8616) );
  OAI22_X1 U10055 ( .A1(n8614), .A2(n8951), .B1(n8640), .B2(n8913), .ZN(n8615)
         );
  AOI211_X1 U10056 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3152), .A(n8616), 
        .B(n8615), .ZN(n8617) );
  OAI211_X1 U10057 ( .C1(n8916), .C2(n8619), .A(n8618), .B(n8617), .ZN(
        P2_U3237) );
  XOR2_X1 U10058 ( .A(n8621), .B(n8620), .Z(n8623) );
  NAND2_X1 U10059 ( .A1(n8623), .A2(n8622), .ZN(n8633) );
  INV_X1 U10060 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10128) );
  NOR2_X1 U10061 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10128), .ZN(n8671) );
  AOI21_X1 U10062 ( .B1(n8624), .B2(n8654), .A(n8671), .ZN(n8632) );
  INV_X1 U10063 ( .A(n8625), .ZN(n8626) );
  AOI22_X1 U10064 ( .A1(n8628), .A2(n8656), .B1(n8627), .B2(n8626), .ZN(n8631)
         );
  NAND2_X1 U10065 ( .A1(n8629), .A2(n9094), .ZN(n8630) );
  NAND4_X1 U10066 ( .A1(n8633), .A2(n8632), .A3(n8631), .A4(n8630), .ZN(
        P2_U3238) );
  XNOR2_X1 U10067 ( .A(n8634), .B(n8635), .ZN(n8644) );
  OR2_X1 U10068 ( .A1(n8883), .A2(n8952), .ZN(n8637) );
  NAND2_X1 U10069 ( .A1(n8646), .A2(n8993), .ZN(n8636) );
  NAND2_X1 U10070 ( .A1(n8637), .A2(n8636), .ZN(n8850) );
  AOI22_X1 U10071 ( .A1(n8850), .A2(n8638), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8639) );
  OAI21_X1 U10072 ( .B1(n8857), .B2(n8640), .A(n8639), .ZN(n8641) );
  AOI21_X1 U10073 ( .B1(n9031), .B2(n8629), .A(n8641), .ZN(n8642) );
  OAI21_X1 U10074 ( .B1(n8644), .B2(n8643), .A(n8642), .ZN(P2_U3242) );
  MUX2_X1 U10075 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8645), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U10076 ( .A(n8795), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8665), .Z(
        P2_U3580) );
  MUX2_X1 U10077 ( .A(n8646), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8665), .Z(
        P2_U3579) );
  INV_X1 U10078 ( .A(n8837), .ZN(n8789) );
  MUX2_X1 U10079 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8789), .S(P2_U3966), .Z(
        P2_U3578) );
  INV_X1 U10080 ( .A(n8883), .ZN(n8787) );
  MUX2_X1 U10081 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8787), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U10082 ( .A(n8893), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8665), .Z(
        P2_U3576) );
  MUX2_X1 U10083 ( .A(n8647), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8665), .Z(
        P2_U3575) );
  INV_X1 U10084 ( .A(n8786), .ZN(n8894) );
  MUX2_X1 U10085 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8894), .S(P2_U3966), .Z(
        P2_U3574) );
  INV_X1 U10086 ( .A(n8951), .ZN(n8783) );
  MUX2_X1 U10087 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8783), .S(P2_U3966), .Z(
        P2_U3573) );
  INV_X1 U10088 ( .A(n8648), .ZN(n8781) );
  MUX2_X1 U10089 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8781), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10090 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8994), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10091 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8778), .S(P2_U3966), .Z(
        P2_U3570) );
  INV_X1 U10092 ( .A(n8649), .ZN(n8996) );
  MUX2_X1 U10093 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8996), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10094 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8650), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10095 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8651), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10096 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8652), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10097 ( .A(n8653), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8665), .Z(
        P2_U3565) );
  MUX2_X1 U10098 ( .A(n8654), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8665), .Z(
        P2_U3564) );
  MUX2_X1 U10099 ( .A(n8655), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8665), .Z(
        P2_U3563) );
  MUX2_X1 U10100 ( .A(n8656), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8665), .Z(
        P2_U3562) );
  MUX2_X1 U10101 ( .A(n8657), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8665), .Z(
        P2_U3561) );
  MUX2_X1 U10102 ( .A(n8658), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8665), .Z(
        P2_U3560) );
  MUX2_X1 U10103 ( .A(n8659), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8665), .Z(
        P2_U3559) );
  MUX2_X1 U10104 ( .A(n8660), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8665), .Z(
        P2_U3558) );
  MUX2_X1 U10105 ( .A(n8661), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8665), .Z(
        P2_U3557) );
  MUX2_X1 U10106 ( .A(n8662), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8665), .Z(
        P2_U3556) );
  MUX2_X1 U10107 ( .A(n8663), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8665), .Z(
        P2_U3555) );
  MUX2_X1 U10108 ( .A(n8664), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8665), .Z(
        P2_U3554) );
  MUX2_X1 U10109 ( .A(n6922), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8665), .Z(
        P2_U3553) );
  MUX2_X1 U10110 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8666), .S(P2_U3966), .Z(
        P2_U3552) );
  OAI21_X1 U10111 ( .B1(n8669), .B2(n8668), .A(n8667), .ZN(n8670) );
  NAND2_X1 U10112 ( .A1(n9856), .A2(n8670), .ZN(n8679) );
  AOI21_X1 U10113 ( .B1(n9854), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8671), .ZN(
        n8678) );
  NAND2_X1 U10114 ( .A1(n9555), .A2(n8672), .ZN(n8677) );
  OAI211_X1 U10115 ( .C1(n8675), .C2(n8674), .A(n9853), .B(n8673), .ZN(n8676)
         );
  NAND4_X1 U10116 ( .A1(n8679), .A2(n8678), .A3(n8677), .A4(n8676), .ZN(
        P2_U3256) );
  OAI21_X1 U10117 ( .B1(n8681), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8680), .ZN(
        n8693) );
  XNOR2_X1 U10118 ( .A(n8701), .B(n8693), .ZN(n8682) );
  NAND2_X1 U10119 ( .A1(n8682), .A2(n7639), .ZN(n8695) );
  OAI21_X1 U10120 ( .B1(n8682), .B2(n7639), .A(n8695), .ZN(n8683) );
  NAND2_X1 U10121 ( .A1(n8683), .A2(n9856), .ZN(n8692) );
  INV_X1 U10122 ( .A(n8684), .ZN(n8685) );
  AOI21_X1 U10123 ( .B1(n9854), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8685), .ZN(
        n8691) );
  AOI21_X1 U10124 ( .B1(n8687), .B2(n5956), .A(n8686), .ZN(n8700) );
  XNOR2_X1 U10125 ( .A(n8700), .B(n8694), .ZN(n8688) );
  NAND2_X1 U10126 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8688), .ZN(n8702) );
  OAI211_X1 U10127 ( .C1(n8688), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9853), .B(
        n8702), .ZN(n8690) );
  NAND2_X1 U10128 ( .A1(n9555), .A2(n8701), .ZN(n8689) );
  NAND4_X1 U10129 ( .A1(n8692), .A2(n8691), .A3(n8690), .A4(n8689), .ZN(
        P2_U3260) );
  NAND2_X1 U10130 ( .A1(n8694), .A2(n8693), .ZN(n8696) );
  NAND2_X1 U10131 ( .A1(n8718), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8697) );
  OAI21_X1 U10132 ( .B1(n8718), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8697), .ZN(
        n8698) );
  AOI211_X1 U10133 ( .C1(n8699), .C2(n8698), .A(n8713), .B(n9549), .ZN(n8712)
         );
  NAND2_X1 U10134 ( .A1(n8701), .A2(n8700), .ZN(n8703) );
  NAND2_X1 U10135 ( .A1(n8703), .A2(n8702), .ZN(n8705) );
  XNOR2_X1 U10136 ( .A(n8718), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8704) );
  NOR2_X1 U10137 ( .A1(n8704), .A2(n8705), .ZN(n8719) );
  AOI21_X1 U10138 ( .B1(n8705), .B2(n8704), .A(n8719), .ZN(n8710) );
  INV_X1 U10139 ( .A(n8706), .ZN(n8707) );
  AOI21_X1 U10140 ( .B1(n9854), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8707), .ZN(
        n8709) );
  NAND2_X1 U10141 ( .A1(n9555), .A2(n8718), .ZN(n8708) );
  OAI211_X1 U10142 ( .C1(n8710), .C2(n9859), .A(n8709), .B(n8708), .ZN(n8711)
         );
  OR2_X1 U10143 ( .A1(n8712), .A2(n8711), .ZN(P2_U3261) );
  NAND2_X1 U10144 ( .A1(n8729), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8714) );
  OAI21_X1 U10145 ( .B1(n8729), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8714), .ZN(
        n8715) );
  AOI211_X1 U10146 ( .C1(n8716), .C2(n8715), .A(n8728), .B(n9549), .ZN(n8727)
         );
  NOR2_X1 U10147 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10065), .ZN(n8717) );
  AOI21_X1 U10148 ( .B1(n9854), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8717), .ZN(
        n8725) );
  XNOR2_X1 U10149 ( .A(n8735), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8723) );
  OR2_X1 U10150 ( .A1(n8718), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8721) );
  INV_X1 U10151 ( .A(n8719), .ZN(n8720) );
  AND2_X1 U10152 ( .A1(n8721), .A2(n8720), .ZN(n8722) );
  NAND2_X1 U10153 ( .A1(n8723), .A2(n8722), .ZN(n8734) );
  OAI211_X1 U10154 ( .C1(n8723), .C2(n8722), .A(n9853), .B(n8734), .ZN(n8724)
         );
  OAI211_X1 U10155 ( .C1(n9857), .C2(n8735), .A(n8725), .B(n8724), .ZN(n8726)
         );
  OR2_X1 U10156 ( .A1(n8727), .A2(n8726), .ZN(P2_U3262) );
  XNOR2_X1 U10157 ( .A(n8747), .B(n8745), .ZN(n8730) );
  NAND2_X1 U10158 ( .A1(n8730), .A2(n6023), .ZN(n8749) );
  OAI21_X1 U10159 ( .B1(n8730), .B2(n6023), .A(n8749), .ZN(n8731) );
  NAND2_X1 U10160 ( .A1(n8731), .A2(n9856), .ZN(n8744) );
  AOI21_X1 U10161 ( .B1(n9854), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8732), .ZN(
        n8743) );
  NAND2_X1 U10162 ( .A1(n9555), .A2(n8745), .ZN(n8742) );
  OR2_X1 U10163 ( .A1(n8745), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8751) );
  NAND2_X1 U10164 ( .A1(n8745), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8733) );
  AND2_X1 U10165 ( .A1(n8751), .A2(n8733), .ZN(n8739) );
  OAI21_X1 U10166 ( .B1(n8736), .B2(n8735), .A(n8734), .ZN(n8737) );
  INV_X1 U10167 ( .A(n8737), .ZN(n8738) );
  NAND2_X1 U10168 ( .A1(n8739), .A2(n8738), .ZN(n8752) );
  OAI21_X1 U10169 ( .B1(n8739), .B2(n8738), .A(n8752), .ZN(n8740) );
  NAND2_X1 U10170 ( .A1(n9853), .A2(n8740), .ZN(n8741) );
  NAND4_X1 U10171 ( .A1(n8744), .A2(n8743), .A3(n8742), .A4(n8741), .ZN(
        P2_U3263) );
  INV_X1 U10172 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8762) );
  INV_X1 U10173 ( .A(n8745), .ZN(n8746) );
  NAND2_X1 U10174 ( .A1(n8747), .A2(n8746), .ZN(n8748) );
  NAND2_X1 U10175 ( .A1(n8749), .A2(n8748), .ZN(n8750) );
  NAND2_X1 U10176 ( .A1(n8752), .A2(n8751), .ZN(n8754) );
  XNOR2_X1 U10177 ( .A(n8754), .B(n8753), .ZN(n8758) );
  INV_X1 U10178 ( .A(n8758), .ZN(n8755) );
  OR2_X1 U10179 ( .A1(n9555), .A2(n8756), .ZN(n8757) );
  NAND2_X1 U10180 ( .A1(n9854), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8760) );
  OAI211_X1 U10181 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n8762), .A(n8761), .B(
        n8760), .ZN(P2_U3264) );
  INV_X1 U10182 ( .A(n9031), .ZN(n8763) );
  XOR2_X1 U10183 ( .A(n9005), .B(n8767), .Z(n9007) );
  INV_X1 U10184 ( .A(P2_B_REG_SCAN_IN), .ZN(n10037) );
  OAI21_X1 U10185 ( .B1(n6715), .B2(n10037), .A(n8993), .ZN(n8775) );
  NOR2_X1 U10186 ( .A1(n8764), .A2(n8775), .ZN(n9004) );
  INV_X1 U10187 ( .A(n9004), .ZN(n9010) );
  NOR2_X1 U10188 ( .A1(n8956), .A2(n9010), .ZN(n8769) );
  AOI21_X1 U10189 ( .B1(n8956), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8769), .ZN(
        n8766) );
  NAND2_X1 U10190 ( .A1(n9005), .A2(n8845), .ZN(n8765) );
  OAI211_X1 U10191 ( .C1(n9007), .C2(n8801), .A(n8766), .B(n8765), .ZN(
        P2_U3265) );
  INV_X1 U10192 ( .A(n8768), .ZN(n9012) );
  INV_X1 U10193 ( .A(n8767), .ZN(n9009) );
  NAND2_X1 U10194 ( .A1(n8800), .A2(n8768), .ZN(n9008) );
  NAND3_X1 U10195 ( .A1(n9009), .A2(n9001), .A3(n9008), .ZN(n8771) );
  AOI21_X1 U10196 ( .B1(n8956), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8769), .ZN(
        n8770) );
  OAI211_X1 U10197 ( .C1(n9012), .C2(n8989), .A(n8771), .B(n8770), .ZN(
        P2_U3266) );
  XNOR2_X1 U10198 ( .A(n8772), .B(n8797), .ZN(n8773) );
  OAI222_X1 U10199 ( .A1(n8952), .A2(n8838), .B1(n8775), .B2(n8774), .C1(n8773), .C2(n8970), .ZN(n9017) );
  INV_X1 U10200 ( .A(n9017), .ZN(n8807) );
  NAND2_X1 U10201 ( .A1(n8777), .A2(n8776), .ZN(n8979) );
  NAND2_X1 U10202 ( .A1(n9072), .A2(n8778), .ZN(n8780) );
  INV_X1 U10203 ( .A(n9068), .ZN(n8966) );
  OAI21_X1 U10204 ( .B1(n8928), .B2(n8951), .A(n8926), .ZN(n8785) );
  NAND2_X1 U10205 ( .A1(n8785), .A2(n8784), .ZN(n8908) );
  AOI22_X1 U10206 ( .A1(n8908), .A2(n8919), .B1(n8916), .B2(n8786), .ZN(n8904)
         );
  OAI22_X1 U10207 ( .A1(n8861), .A2(n8871), .B1(n9037), .B2(n8787), .ZN(n8844)
         );
  NAND2_X1 U10208 ( .A1(n8844), .A2(n8788), .ZN(n8791) );
  NAND2_X1 U10209 ( .A1(n8791), .A2(n8790), .ZN(n8824) );
  NAND2_X1 U10210 ( .A1(n8824), .A2(n8792), .ZN(n8794) );
  NAND2_X1 U10211 ( .A1(n8830), .A2(n8817), .ZN(n8793) );
  NAND2_X1 U10212 ( .A1(n8794), .A2(n8793), .ZN(n8809) );
  INV_X1 U10213 ( .A(n8808), .ZN(n8814) );
  NOR2_X1 U10214 ( .A1(n9020), .A2(n8795), .ZN(n8796) );
  AOI21_X1 U10215 ( .B1(n8809), .B2(n8814), .A(n8796), .ZN(n8798) );
  XNOR2_X1 U10216 ( .A(n8798), .B(n8797), .ZN(n9013) );
  NAND2_X1 U10217 ( .A1(n9013), .A2(n8905), .ZN(n8806) );
  OAI22_X1 U10218 ( .A1(n8936), .A2(n10174), .B1(n8799), .B2(n8934), .ZN(n8803) );
  OAI21_X1 U10219 ( .B1(n4396), .B2(n9014), .A(n8800), .ZN(n9015) );
  NOR2_X1 U10220 ( .A1(n9015), .A2(n8801), .ZN(n8802) );
  AOI211_X1 U10221 ( .C1(n8845), .C2(n8804), .A(n8803), .B(n8802), .ZN(n8805)
         );
  OAI211_X1 U10222 ( .C1(n8807), .C2(n8956), .A(n8806), .B(n8805), .ZN(
        P2_U3267) );
  XNOR2_X1 U10223 ( .A(n8809), .B(n8808), .ZN(n9024) );
  AOI21_X1 U10224 ( .B1(n9020), .B2(n8825), .A(n4396), .ZN(n9021) );
  AOI22_X1 U10225 ( .A1(n8987), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8810), .B2(
        n8985), .ZN(n8811) );
  OAI21_X1 U10226 ( .B1(n8812), .B2(n8989), .A(n8811), .ZN(n8822) );
  INV_X1 U10227 ( .A(n8813), .ZN(n8815) );
  AOI21_X1 U10228 ( .B1(n8815), .B2(n8814), .A(n8970), .ZN(n8820) );
  OAI22_X1 U10229 ( .A1(n8817), .A2(n8952), .B1(n8816), .B2(n8950), .ZN(n8818)
         );
  AOI21_X1 U10230 ( .B1(n8820), .B2(n8819), .A(n8818), .ZN(n9023) );
  NOR2_X1 U10231 ( .A1(n9023), .A2(n8956), .ZN(n8821) );
  AOI211_X1 U10232 ( .C1(n9001), .C2(n9021), .A(n8822), .B(n8821), .ZN(n8823)
         );
  OAI21_X1 U10233 ( .B1(n9003), .B2(n9024), .A(n8823), .ZN(P2_U3268) );
  XNOR2_X1 U10234 ( .A(n8824), .B(n8833), .ZN(n9029) );
  INV_X1 U10235 ( .A(n8825), .ZN(n8826) );
  AOI21_X1 U10236 ( .B1(n9025), .B2(n8852), .A(n8826), .ZN(n9026) );
  INV_X1 U10237 ( .A(n8827), .ZN(n8828) );
  AOI22_X1 U10238 ( .A1(n8987), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8828), .B2(
        n8985), .ZN(n8829) );
  OAI21_X1 U10239 ( .B1(n8830), .B2(n8989), .A(n8829), .ZN(n8842) );
  INV_X1 U10240 ( .A(n8831), .ZN(n8836) );
  AOI21_X1 U10241 ( .B1(n8847), .B2(n8834), .A(n8833), .ZN(n8835) );
  NOR3_X1 U10242 ( .A1(n8836), .A2(n8835), .A3(n8970), .ZN(n8840) );
  OAI22_X1 U10243 ( .A1(n8838), .A2(n8950), .B1(n8837), .B2(n8952), .ZN(n8839)
         );
  NOR2_X1 U10244 ( .A1(n8840), .A2(n8839), .ZN(n9028) );
  NOR2_X1 U10245 ( .A1(n9028), .A2(n8956), .ZN(n8841) );
  AOI211_X1 U10246 ( .C1(n9001), .C2(n9026), .A(n8842), .B(n8841), .ZN(n8843)
         );
  OAI21_X1 U10247 ( .B1(n9029), .B2(n9003), .A(n8843), .ZN(P2_U3269) );
  XNOR2_X1 U10248 ( .A(n8844), .B(n8848), .ZN(n9034) );
  AOI22_X1 U10249 ( .A1(n9031), .A2(n8845), .B1(n8956), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8860) );
  AND2_X1 U10250 ( .A1(n8869), .A2(n8846), .ZN(n8849) );
  OAI21_X1 U10251 ( .B1(n8849), .B2(n8848), .A(n8847), .ZN(n8851) );
  AOI21_X1 U10252 ( .B1(n8851), .B2(n8998), .A(n8850), .ZN(n9033) );
  INV_X1 U10253 ( .A(n8862), .ZN(n8854) );
  INV_X1 U10254 ( .A(n8852), .ZN(n8853) );
  AOI211_X1 U10255 ( .C1(n9031), .C2(n8854), .A(n9927), .B(n8853), .ZN(n9030)
         );
  NAND2_X1 U10256 ( .A1(n9030), .A2(n8855), .ZN(n8856) );
  OAI211_X1 U10257 ( .C1(n8934), .C2(n8857), .A(n9033), .B(n8856), .ZN(n8858)
         );
  NAND2_X1 U10258 ( .A1(n8858), .A2(n8936), .ZN(n8859) );
  OAI211_X1 U10259 ( .C1(n9034), .C2(n9003), .A(n8860), .B(n8859), .ZN(
        P2_U3270) );
  XOR2_X1 U10260 ( .A(n8871), .B(n8861), .Z(n9039) );
  AOI211_X1 U10261 ( .C1(n9037), .C2(n8863), .A(n9927), .B(n8862), .ZN(n9036)
         );
  INV_X1 U10262 ( .A(n9037), .ZN(n8864) );
  NOR2_X1 U10263 ( .A1(n8864), .A2(n8989), .ZN(n8868) );
  OAI22_X1 U10264 ( .A1(n8936), .A2(n8866), .B1(n8865), .B2(n8934), .ZN(n8867)
         );
  AOI211_X1 U10265 ( .C1(n9036), .C2(n8977), .A(n8868), .B(n8867), .ZN(n8875)
         );
  OAI211_X1 U10266 ( .C1(n8871), .C2(n8870), .A(n8869), .B(n8998), .ZN(n8873)
         );
  NAND2_X1 U10267 ( .A1(n8873), .A2(n8872), .ZN(n9035) );
  NAND2_X1 U10268 ( .A1(n9035), .A2(n8936), .ZN(n8874) );
  OAI211_X1 U10269 ( .C1(n9039), .C2(n9003), .A(n8875), .B(n8874), .ZN(
        P2_U3271) );
  AOI21_X1 U10270 ( .B1(n8284), .B2(n8876), .A(n4426), .ZN(n9044) );
  XNOR2_X1 U10271 ( .A(n8896), .B(n8880), .ZN(n9041) );
  INV_X1 U10272 ( .A(n8877), .ZN(n8878) );
  AOI22_X1 U10273 ( .A1(n8987), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8878), .B2(
        n8985), .ZN(n8879) );
  OAI21_X1 U10274 ( .B1(n8880), .B2(n8989), .A(n8879), .ZN(n8888) );
  AOI21_X1 U10275 ( .B1(n8882), .B2(n8881), .A(n8970), .ZN(n8886) );
  OAI22_X1 U10276 ( .A1(n8920), .A2(n8952), .B1(n8883), .B2(n8950), .ZN(n8884)
         );
  AOI21_X1 U10277 ( .B1(n8886), .B2(n8885), .A(n8884), .ZN(n9043) );
  NOR2_X1 U10278 ( .A1(n9043), .A2(n8956), .ZN(n8887) );
  AOI211_X1 U10279 ( .C1(n9041), .C2(n9001), .A(n8888), .B(n8887), .ZN(n8889)
         );
  OAI21_X1 U10280 ( .B1(n9003), .B2(n9044), .A(n8889), .ZN(P2_U3272) );
  OAI21_X1 U10281 ( .B1(n8892), .B2(n8891), .A(n8890), .ZN(n8895) );
  AOI222_X1 U10282 ( .A1(n8998), .A2(n8895), .B1(n8894), .B2(n8995), .C1(n8893), .C2(n8993), .ZN(n9051) );
  INV_X1 U10283 ( .A(n8896), .ZN(n8897) );
  AOI21_X1 U10284 ( .B1(n9045), .B2(n8910), .A(n8897), .ZN(n9046) );
  NOR2_X1 U10285 ( .A1(n8898), .A2(n8989), .ZN(n8902) );
  OAI22_X1 U10286 ( .A1(n8936), .A2(n8900), .B1(n8899), .B2(n8934), .ZN(n8901)
         );
  AOI211_X1 U10287 ( .C1(n9046), .C2(n9001), .A(n8902), .B(n8901), .ZN(n8907)
         );
  OR2_X1 U10288 ( .A1(n8904), .A2(n8903), .ZN(n9048) );
  NAND3_X1 U10289 ( .A1(n9048), .A2(n9047), .A3(n8905), .ZN(n8906) );
  OAI211_X1 U10290 ( .C1(n9051), .C2(n8956), .A(n8907), .B(n8906), .ZN(
        P2_U3273) );
  XOR2_X1 U10291 ( .A(n8908), .B(n8919), .Z(n9056) );
  INV_X1 U10292 ( .A(n8909), .ZN(n8912) );
  INV_X1 U10293 ( .A(n8910), .ZN(n8911) );
  AOI21_X1 U10294 ( .B1(n9052), .B2(n8912), .A(n8911), .ZN(n9053) );
  INV_X1 U10295 ( .A(n8913), .ZN(n8914) );
  AOI22_X1 U10296 ( .A1(n8987), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8914), .B2(
        n8985), .ZN(n8915) );
  OAI21_X1 U10297 ( .B1(n8916), .B2(n8989), .A(n8915), .ZN(n8924) );
  AOI211_X1 U10298 ( .C1(n8919), .C2(n8918), .A(n8970), .B(n8917), .ZN(n8922)
         );
  OAI22_X1 U10299 ( .A1(n8920), .A2(n8950), .B1(n8951), .B2(n8952), .ZN(n8921)
         );
  NOR2_X1 U10300 ( .A1(n8922), .A2(n8921), .ZN(n9055) );
  NOR2_X1 U10301 ( .A1(n9055), .A2(n8956), .ZN(n8923) );
  AOI211_X1 U10302 ( .C1(n9053), .C2(n9001), .A(n8924), .B(n8923), .ZN(n8925)
         );
  OAI21_X1 U10303 ( .B1(n9003), .B2(n9056), .A(n8925), .ZN(P2_U3274) );
  XOR2_X1 U10304 ( .A(n8926), .B(n8930), .Z(n9061) );
  XNOR2_X1 U10305 ( .A(n4447), .B(n9057), .ZN(n9058) );
  OAI22_X1 U10306 ( .A1(n8928), .A2(n8989), .B1(n8936), .B2(n8927), .ZN(n8929)
         );
  AOI21_X1 U10307 ( .B1(n9058), .B2(n9001), .A(n8929), .ZN(n8939) );
  XNOR2_X1 U10308 ( .A(n8931), .B(n8930), .ZN(n8933) );
  AOI21_X1 U10309 ( .B1(n8933), .B2(n8998), .A(n8932), .ZN(n9060) );
  OAI21_X1 U10310 ( .B1(n8935), .B2(n8934), .A(n9060), .ZN(n8937) );
  NAND2_X1 U10311 ( .A1(n8937), .A2(n8936), .ZN(n8938) );
  OAI211_X1 U10312 ( .C1(n9061), .C2(n9003), .A(n8939), .B(n8938), .ZN(
        P2_U3275) );
  XNOR2_X1 U10313 ( .A(n8941), .B(n8940), .ZN(n9066) );
  AOI21_X1 U10314 ( .B1(n9062), .B2(n8961), .A(n4447), .ZN(n9063) );
  INV_X1 U10315 ( .A(n8942), .ZN(n8943) );
  AOI22_X1 U10316 ( .A1(n8987), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8943), .B2(
        n8985), .ZN(n8944) );
  OAI21_X1 U10317 ( .B1(n4629), .B2(n8989), .A(n8944), .ZN(n8958) );
  INV_X1 U10318 ( .A(n8945), .ZN(n8949) );
  AOI21_X1 U10319 ( .B1(n8971), .B2(n8947), .A(n8946), .ZN(n8948) );
  NOR3_X1 U10320 ( .A1(n8949), .A2(n8948), .A3(n8970), .ZN(n8955) );
  OAI22_X1 U10321 ( .A1(n8953), .A2(n8952), .B1(n8951), .B2(n8950), .ZN(n8954)
         );
  NOR2_X1 U10322 ( .A1(n8955), .A2(n8954), .ZN(n9065) );
  NOR2_X1 U10323 ( .A1(n9065), .A2(n8956), .ZN(n8957) );
  AOI211_X1 U10324 ( .C1(n9063), .C2(n9001), .A(n8958), .B(n8957), .ZN(n8959)
         );
  OAI21_X1 U10325 ( .B1(n9003), .B2(n9066), .A(n8959), .ZN(P2_U3276) );
  XNOR2_X1 U10326 ( .A(n8960), .B(n8967), .ZN(n9071) );
  INV_X1 U10327 ( .A(n8961), .ZN(n8962) );
  AOI211_X1 U10328 ( .C1(n9068), .C2(n8981), .A(n9927), .B(n8962), .ZN(n9067)
         );
  INV_X1 U10329 ( .A(n8963), .ZN(n8964) );
  AOI22_X1 U10330 ( .A1(n8987), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8964), .B2(
        n8985), .ZN(n8965) );
  OAI21_X1 U10331 ( .B1(n8966), .B2(n8989), .A(n8965), .ZN(n8976) );
  OAI21_X1 U10332 ( .B1(n8969), .B2(n8968), .A(n8967), .ZN(n8972) );
  AOI21_X1 U10333 ( .B1(n8972), .B2(n8971), .A(n8970), .ZN(n8974) );
  NOR2_X1 U10334 ( .A1(n8974), .A2(n8973), .ZN(n9070) );
  NOR2_X1 U10335 ( .A1(n9070), .A2(n8956), .ZN(n8975) );
  AOI211_X1 U10336 ( .C1(n9067), .C2(n8977), .A(n8976), .B(n8975), .ZN(n8978)
         );
  OAI21_X1 U10337 ( .B1(n9003), .B2(n9071), .A(n8978), .ZN(P2_U3277) );
  XNOR2_X1 U10338 ( .A(n8979), .B(n8991), .ZN(n9076) );
  INV_X1 U10339 ( .A(n8980), .ZN(n8983) );
  INV_X1 U10340 ( .A(n8981), .ZN(n8982) );
  AOI21_X1 U10341 ( .B1(n9072), .B2(n8983), .A(n8982), .ZN(n9073) );
  INV_X1 U10342 ( .A(n8984), .ZN(n8986) );
  AOI22_X1 U10343 ( .A1(n8987), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8986), .B2(
        n8985), .ZN(n8988) );
  OAI21_X1 U10344 ( .B1(n8990), .B2(n8989), .A(n8988), .ZN(n9000) );
  XNOR2_X1 U10345 ( .A(n8992), .B(n8991), .ZN(n8997) );
  AOI222_X1 U10346 ( .A1(n8998), .A2(n8997), .B1(n8996), .B2(n8995), .C1(n8994), .C2(n8993), .ZN(n9075) );
  NOR2_X1 U10347 ( .A1(n9075), .A2(n8956), .ZN(n8999) );
  AOI211_X1 U10348 ( .C1(n9073), .C2(n9001), .A(n9000), .B(n8999), .ZN(n9002)
         );
  OAI21_X1 U10349 ( .B1(n9003), .B2(n9076), .A(n9002), .ZN(P2_U3278) );
  AOI21_X1 U10350 ( .B1(n9005), .B2(n9898), .A(n9004), .ZN(n9006) );
  OAI21_X1 U10351 ( .B1(n9007), .B2(n9927), .A(n9006), .ZN(n9105) );
  MUX2_X1 U10352 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9105), .S(n9947), .Z(
        P2_U3551) );
  NAND3_X1 U10353 ( .A1(n9009), .A2(n9899), .A3(n9008), .ZN(n9011) );
  OAI211_X1 U10354 ( .C1(n9012), .C2(n9925), .A(n9011), .B(n9010), .ZN(n9106)
         );
  MUX2_X1 U10355 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9106), .S(n9947), .Z(
        P2_U3550) );
  NAND2_X1 U10356 ( .A1(n9013), .A2(n9931), .ZN(n9019) );
  OAI22_X1 U10357 ( .A1(n9015), .A2(n9927), .B1(n9014), .B2(n9925), .ZN(n9016)
         );
  NOR2_X1 U10358 ( .A1(n9017), .A2(n9016), .ZN(n9018) );
  NAND2_X1 U10359 ( .A1(n9019), .A2(n9018), .ZN(n9107) );
  MUX2_X1 U10360 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9107), .S(n9947), .Z(
        P2_U3549) );
  AOI22_X1 U10361 ( .A1(n9021), .A2(n9899), .B1(n9898), .B2(n9020), .ZN(n9022)
         );
  OAI211_X1 U10362 ( .C1(n9024), .C2(n9874), .A(n9023), .B(n9022), .ZN(n9108)
         );
  MUX2_X1 U10363 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9108), .S(n9947), .Z(
        P2_U3548) );
  AOI22_X1 U10364 ( .A1(n9026), .A2(n9899), .B1(n9898), .B2(n9025), .ZN(n9027)
         );
  OAI211_X1 U10365 ( .C1(n9029), .C2(n9874), .A(n9028), .B(n9027), .ZN(n9109)
         );
  MUX2_X1 U10366 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9109), .S(n9947), .Z(
        P2_U3547) );
  AOI21_X1 U10367 ( .B1(n9898), .B2(n9031), .A(n9030), .ZN(n9032) );
  OAI211_X1 U10368 ( .C1(n9034), .C2(n9874), .A(n9033), .B(n9032), .ZN(n9110)
         );
  MUX2_X1 U10369 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9110), .S(n9947), .Z(
        P2_U3546) );
  AOI211_X1 U10370 ( .C1(n9898), .C2(n9037), .A(n9036), .B(n9035), .ZN(n9038)
         );
  OAI21_X1 U10371 ( .B1(n9039), .B2(n9874), .A(n9038), .ZN(n9111) );
  MUX2_X1 U10372 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9111), .S(n9947), .Z(
        P2_U3545) );
  AOI22_X1 U10373 ( .A1(n9041), .A2(n9899), .B1(n9898), .B2(n9040), .ZN(n9042)
         );
  OAI211_X1 U10374 ( .C1(n9044), .C2(n9874), .A(n9043), .B(n9042), .ZN(n9112)
         );
  MUX2_X1 U10375 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9112), .S(n9947), .Z(
        P2_U3544) );
  AOI22_X1 U10376 ( .A1(n9046), .A2(n9899), .B1(n9898), .B2(n9045), .ZN(n9050)
         );
  NAND3_X1 U10377 ( .A1(n9048), .A2(n9047), .A3(n9931), .ZN(n9049) );
  NAND3_X1 U10378 ( .A1(n9051), .A2(n9050), .A3(n9049), .ZN(n9113) );
  MUX2_X1 U10379 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9113), .S(n9947), .Z(
        P2_U3543) );
  AOI22_X1 U10380 ( .A1(n9053), .A2(n9899), .B1(n9898), .B2(n9052), .ZN(n9054)
         );
  OAI211_X1 U10381 ( .C1(n9056), .C2(n9874), .A(n9055), .B(n9054), .ZN(n9114)
         );
  MUX2_X1 U10382 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9114), .S(n9947), .Z(
        P2_U3542) );
  AOI22_X1 U10383 ( .A1(n9058), .A2(n9899), .B1(n9898), .B2(n9057), .ZN(n9059)
         );
  OAI211_X1 U10384 ( .C1(n9061), .C2(n9874), .A(n9060), .B(n9059), .ZN(n9115)
         );
  MUX2_X1 U10385 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9115), .S(n9947), .Z(
        P2_U3541) );
  AOI22_X1 U10386 ( .A1(n9063), .A2(n9899), .B1(n9898), .B2(n9062), .ZN(n9064)
         );
  OAI211_X1 U10387 ( .C1(n9066), .C2(n9874), .A(n9065), .B(n9064), .ZN(n9116)
         );
  MUX2_X1 U10388 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9116), .S(n9947), .Z(
        P2_U3540) );
  AOI21_X1 U10389 ( .B1(n9898), .B2(n9068), .A(n9067), .ZN(n9069) );
  OAI211_X1 U10390 ( .C1(n9071), .C2(n9874), .A(n9070), .B(n9069), .ZN(n9117)
         );
  MUX2_X1 U10391 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9117), .S(n9947), .Z(
        P2_U3539) );
  AOI22_X1 U10392 ( .A1(n9073), .A2(n9899), .B1(n9898), .B2(n9072), .ZN(n9074)
         );
  OAI211_X1 U10393 ( .C1(n9874), .C2(n9076), .A(n9075), .B(n9074), .ZN(n9118)
         );
  MUX2_X1 U10394 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9118), .S(n9947), .Z(
        P2_U3538) );
  INV_X1 U10395 ( .A(n9077), .ZN(n9082) );
  AOI21_X1 U10396 ( .B1(n9898), .B2(n9079), .A(n9078), .ZN(n9080) );
  OAI211_X1 U10397 ( .C1(n9874), .C2(n9082), .A(n9081), .B(n9080), .ZN(n9119)
         );
  MUX2_X1 U10398 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9119), .S(n9947), .Z(
        P2_U3537) );
  AOI22_X1 U10399 ( .A1(n9084), .A2(n9899), .B1(n9898), .B2(n9083), .ZN(n9085)
         );
  OAI211_X1 U10400 ( .C1(n9103), .C2(n9087), .A(n9086), .B(n9085), .ZN(n9120)
         );
  MUX2_X1 U10401 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9120), .S(n9947), .Z(
        P2_U3536) );
  INV_X1 U10402 ( .A(n9088), .ZN(n9093) );
  AOI22_X1 U10403 ( .A1(n9090), .A2(n9899), .B1(n9898), .B2(n9089), .ZN(n9091)
         );
  OAI211_X1 U10404 ( .C1(n9103), .C2(n9093), .A(n9092), .B(n9091), .ZN(n9121)
         );
  MUX2_X1 U10405 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9121), .S(n9947), .Z(
        P2_U3533) );
  AOI22_X1 U10406 ( .A1(n9095), .A2(n9899), .B1(n9898), .B2(n9094), .ZN(n9096)
         );
  OAI211_X1 U10407 ( .C1(n9874), .C2(n9098), .A(n9097), .B(n9096), .ZN(n9122)
         );
  MUX2_X1 U10408 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9122), .S(n9947), .Z(
        P2_U3531) );
  AOI22_X1 U10409 ( .A1(n9100), .A2(n9899), .B1(n9898), .B2(n9099), .ZN(n9101)
         );
  OAI211_X1 U10410 ( .C1(n9104), .C2(n9103), .A(n9102), .B(n9101), .ZN(n9123)
         );
  MUX2_X1 U10411 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n9123), .S(n9947), .Z(
        P2_U3529) );
  MUX2_X1 U10412 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9105), .S(n9935), .Z(
        P2_U3519) );
  MUX2_X1 U10413 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9106), .S(n9935), .Z(
        P2_U3518) );
  MUX2_X1 U10414 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9107), .S(n9935), .Z(
        P2_U3517) );
  MUX2_X1 U10415 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9108), .S(n9935), .Z(
        P2_U3516) );
  MUX2_X1 U10416 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9109), .S(n9935), .Z(
        P2_U3515) );
  MUX2_X1 U10417 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9110), .S(n9935), .Z(
        P2_U3514) );
  MUX2_X1 U10418 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9111), .S(n9935), .Z(
        P2_U3513) );
  MUX2_X1 U10419 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9112), .S(n9935), .Z(
        P2_U3512) );
  MUX2_X1 U10420 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9113), .S(n9935), .Z(
        P2_U3511) );
  MUX2_X1 U10421 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9114), .S(n9935), .Z(
        P2_U3510) );
  MUX2_X1 U10422 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9115), .S(n9935), .Z(
        P2_U3509) );
  MUX2_X1 U10423 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9116), .S(n9935), .Z(
        P2_U3508) );
  MUX2_X1 U10424 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9117), .S(n9935), .Z(
        P2_U3507) );
  MUX2_X1 U10425 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9118), .S(n9935), .Z(
        P2_U3505) );
  MUX2_X1 U10426 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9119), .S(n9935), .Z(
        P2_U3502) );
  MUX2_X1 U10427 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9120), .S(n9935), .Z(
        P2_U3499) );
  MUX2_X1 U10428 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9121), .S(n9935), .Z(
        P2_U3490) );
  MUX2_X1 U10429 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n9122), .S(n9935), .Z(
        P2_U3484) );
  MUX2_X1 U10430 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n9123), .S(n9935), .Z(
        P2_U3478) );
  NAND3_X1 U10431 ( .A1(n9124), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n9125) );
  OAI22_X1 U10432 ( .A1(n4463), .A2(n9125), .B1(n6604), .B2(n10258), .ZN(n9126) );
  AOI21_X1 U10433 ( .B1(n8298), .B2(n9127), .A(n9126), .ZN(n9128) );
  INV_X1 U10434 ( .A(n9128), .ZN(P2_U3327) );
  MUX2_X1 U10435 ( .A(n9129), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XOR2_X1 U10436 ( .A(n9131), .B(n9130), .Z(n9132) );
  XNOR2_X1 U10437 ( .A(n9133), .B(n9132), .ZN(n9142) );
  OAI22_X1 U10438 ( .A1(n9135), .A2(n9207), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9134), .ZN(n9136) );
  AOI21_X1 U10439 ( .B1(n9137), .B2(n9211), .A(n9136), .ZN(n9138) );
  OAI21_X1 U10440 ( .B1(n9139), .B2(n9208), .A(n9138), .ZN(n9140) );
  AOI21_X1 U10441 ( .B1(n9438), .B2(n9199), .A(n9140), .ZN(n9141) );
  OAI21_X1 U10442 ( .B1(n9142), .B2(n9201), .A(n9141), .ZN(P1_U3212) );
  INV_X1 U10443 ( .A(n9143), .ZN(n9145) );
  NAND2_X1 U10444 ( .A1(n9145), .A2(n9144), .ZN(n9147) );
  XNOR2_X1 U10445 ( .A(n9147), .B(n9146), .ZN(n9154) );
  AOI22_X1 U10446 ( .A1(n9321), .A2(n9183), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9150) );
  NAND2_X1 U10447 ( .A1(n9211), .A2(n9148), .ZN(n9149) );
  OAI211_X1 U10448 ( .C1(n9151), .C2(n9207), .A(n9150), .B(n9149), .ZN(n9152)
         );
  AOI21_X1 U10449 ( .B1(n9460), .B2(n9188), .A(n9152), .ZN(n9153) );
  OAI21_X1 U10450 ( .B1(n9154), .B2(n9201), .A(n9153), .ZN(P1_U3214) );
  XOR2_X1 U10451 ( .A(n9156), .B(n9155), .Z(n9161) );
  AOI22_X1 U10452 ( .A1(n9396), .A2(n9194), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9158) );
  NAND2_X1 U10453 ( .A1(n9366), .A2(n9183), .ZN(n9157) );
  OAI211_X1 U10454 ( .C1(n9186), .C2(n9358), .A(n9158), .B(n9157), .ZN(n9159)
         );
  AOI21_X1 U10455 ( .B1(n9471), .B2(n9188), .A(n9159), .ZN(n9160) );
  OAI21_X1 U10456 ( .B1(n9161), .B2(n9201), .A(n9160), .ZN(P1_U3221) );
  XOR2_X1 U10457 ( .A(n9163), .B(n9162), .Z(n9169) );
  AOI22_X1 U10458 ( .A1(n9321), .A2(n9194), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9164) );
  OAI21_X1 U10459 ( .B1(n9186), .B2(n9326), .A(n9164), .ZN(n9167) );
  NAND2_X1 U10460 ( .A1(n5571), .A2(n9500), .ZN(n9450) );
  NOR2_X1 U10461 ( .A1(n9450), .A2(n9165), .ZN(n9166) );
  AOI211_X1 U10462 ( .C1(n9183), .C2(n9320), .A(n9167), .B(n9166), .ZN(n9168)
         );
  OAI21_X1 U10463 ( .B1(n9169), .B2(n9201), .A(n9168), .ZN(P1_U3223) );
  XOR2_X1 U10464 ( .A(n9171), .B(n9170), .Z(n9176) );
  OAI22_X1 U10465 ( .A1(n9340), .A2(n9207), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10014), .ZN(n9172) );
  AOI21_X1 U10466 ( .B1(n9217), .B2(n9183), .A(n9172), .ZN(n9173) );
  OAI21_X1 U10467 ( .B1(n9186), .B2(n9348), .A(n9173), .ZN(n9174) );
  AOI21_X1 U10468 ( .B1(n9344), .B2(n9188), .A(n9174), .ZN(n9175) );
  OAI21_X1 U10469 ( .B1(n9176), .B2(n9201), .A(n9175), .ZN(P1_U3227) );
  INV_X1 U10470 ( .A(n9177), .ZN(n9182) );
  AOI21_X1 U10471 ( .B1(n9179), .B2(n9181), .A(n9178), .ZN(n9180) );
  AOI21_X1 U10472 ( .B1(n9182), .B2(n9181), .A(n9180), .ZN(n9190) );
  NAND2_X1 U10473 ( .A1(n9219), .A2(n9183), .ZN(n9185) );
  AOI22_X1 U10474 ( .A1(n9194), .A2(n9418), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9184) );
  OAI211_X1 U10475 ( .C1(n9186), .C2(n9374), .A(n9185), .B(n9184), .ZN(n9187)
         );
  AOI21_X1 U10476 ( .B1(n9476), .B2(n9188), .A(n9187), .ZN(n9189) );
  OAI21_X1 U10477 ( .B1(n9190), .B2(n9201), .A(n9189), .ZN(P1_U3231) );
  NAND2_X1 U10478 ( .A1(n4433), .A2(n9191), .ZN(n9193) );
  XNOR2_X1 U10479 ( .A(n9193), .B(n9192), .ZN(n9202) );
  AOI22_X1 U10480 ( .A1(n9219), .A2(n9194), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9197) );
  NAND2_X1 U10481 ( .A1(n9211), .A2(n9195), .ZN(n9196) );
  OAI211_X1 U10482 ( .C1(n9340), .C2(n9208), .A(n9197), .B(n9196), .ZN(n9198)
         );
  AOI21_X1 U10483 ( .B1(n9465), .B2(n9199), .A(n9198), .ZN(n9200) );
  OAI21_X1 U10484 ( .B1(n9202), .B2(n9201), .A(n9200), .ZN(P1_U3233) );
  OAI211_X1 U10485 ( .C1(n9206), .C2(n9205), .A(n9203), .B(n9204), .ZN(n9213)
         );
  OAI22_X1 U10486 ( .A1(n9341), .A2(n9207), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9978), .ZN(n9210) );
  NOR2_X1 U10487 ( .A1(n9312), .A2(n9208), .ZN(n9209) );
  AOI211_X1 U10488 ( .C1(n9305), .C2(n9211), .A(n9210), .B(n9209), .ZN(n9212)
         );
  OAI211_X1 U10489 ( .C1(n9307), .C2(n9214), .A(n9213), .B(n9212), .ZN(
        P1_U3238) );
  MUX2_X1 U10490 ( .A(n9215), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9234), .Z(
        P1_U3585) );
  MUX2_X1 U10491 ( .A(n9291), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9234), .Z(
        P1_U3584) );
  MUX2_X1 U10492 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n5568), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10493 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9216), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10494 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9320), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10495 ( .A(n9217), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9234), .Z(
        P1_U3580) );
  MUX2_X1 U10496 ( .A(n9321), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9234), .Z(
        P1_U3579) );
  MUX2_X1 U10497 ( .A(n9218), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9234), .Z(
        P1_U3578) );
  MUX2_X1 U10498 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9366), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10499 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9219), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10500 ( .A(n9396), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9234), .Z(
        P1_U3575) );
  MUX2_X1 U10501 ( .A(n9418), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9234), .Z(
        P1_U3574) );
  MUX2_X1 U10502 ( .A(n9397), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9234), .Z(
        P1_U3573) );
  MUX2_X1 U10503 ( .A(n9420), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9234), .Z(
        P1_U3572) );
  MUX2_X1 U10504 ( .A(n9220), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9234), .Z(
        P1_U3571) );
  MUX2_X1 U10505 ( .A(n9221), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9234), .Z(
        P1_U3570) );
  MUX2_X1 U10506 ( .A(n9222), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9234), .Z(
        P1_U3569) );
  MUX2_X1 U10507 ( .A(n9223), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9234), .Z(
        P1_U3568) );
  MUX2_X1 U10508 ( .A(n9224), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9234), .Z(
        P1_U3567) );
  MUX2_X1 U10509 ( .A(n9225), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9234), .Z(
        P1_U3566) );
  MUX2_X1 U10510 ( .A(n9226), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9234), .Z(
        P1_U3565) );
  MUX2_X1 U10511 ( .A(n9227), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9234), .Z(
        P1_U3564) );
  MUX2_X1 U10512 ( .A(n9228), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9234), .Z(
        P1_U3563) );
  MUX2_X1 U10513 ( .A(n9229), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9234), .Z(
        P1_U3562) );
  MUX2_X1 U10514 ( .A(n9230), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9234), .Z(
        P1_U3561) );
  MUX2_X1 U10515 ( .A(n9231), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9234), .Z(
        P1_U3560) );
  MUX2_X1 U10516 ( .A(n9232), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9234), .Z(
        P1_U3559) );
  MUX2_X1 U10517 ( .A(n9233), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9234), .Z(
        P1_U3558) );
  MUX2_X1 U10518 ( .A(n6974), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9234), .Z(
        P1_U3557) );
  MUX2_X1 U10519 ( .A(n6258), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9234), .Z(
        P1_U3556) );
  MUX2_X1 U10520 ( .A(n9235), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9234), .Z(
        P1_U3555) );
  INV_X1 U10521 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9275) );
  NAND2_X1 U10522 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9675), .ZN(n9236) );
  OAI21_X1 U10523 ( .B1(n9675), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9236), .ZN(
        n9671) );
  OAI21_X1 U10524 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9248), .A(n9237), .ZN(
        n9672) );
  NOR2_X1 U10525 ( .A1(n9671), .A2(n9672), .ZN(n9670) );
  OR2_X1 U10526 ( .A1(n9684), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9239) );
  NAND2_X1 U10527 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n9684), .ZN(n9238) );
  NAND2_X1 U10528 ( .A1(n9239), .A2(n9238), .ZN(n9687) );
  NOR2_X1 U10529 ( .A1(n9240), .A2(n9255), .ZN(n9241) );
  NOR2_X1 U10530 ( .A1(n7749), .A2(n9701), .ZN(n9700) );
  NOR2_X1 U10531 ( .A1(n9241), .A2(n9700), .ZN(n9242) );
  NOR2_X1 U10532 ( .A1(n9242), .A2(n9257), .ZN(n9243) );
  NAND2_X1 U10533 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9728), .ZN(n9244) );
  OAI21_X1 U10534 ( .B1(n9728), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9244), .ZN(
        n9725) );
  AOI21_X1 U10535 ( .B1(n9728), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9724), .ZN(
        n9736) );
  OR2_X1 U10536 ( .A1(n9739), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9246) );
  NAND2_X1 U10537 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9739), .ZN(n9245) );
  NAND2_X1 U10538 ( .A1(n9246), .A2(n9245), .ZN(n9737) );
  NOR2_X1 U10539 ( .A1(n9736), .A2(n9737), .ZN(n9735) );
  MUX2_X1 U10540 ( .A(n9247), .B(P1_REG2_REG_18__SCAN_IN), .S(n9752), .Z(n9755) );
  INV_X1 U10541 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9264) );
  XNOR2_X1 U10542 ( .A(n9752), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9764) );
  INV_X1 U10543 ( .A(n9739), .ZN(n9262) );
  XNOR2_X1 U10544 ( .A(n9262), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9746) );
  INV_X1 U10545 ( .A(n9728), .ZN(n9260) );
  INV_X1 U10546 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9259) );
  XOR2_X1 U10547 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9728), .Z(n9730) );
  INV_X1 U10548 ( .A(n9684), .ZN(n9253) );
  INV_X1 U10549 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9252) );
  INV_X1 U10550 ( .A(n9675), .ZN(n9251) );
  INV_X1 U10551 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9615) );
  NOR2_X1 U10552 ( .A1(n9248), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9249) );
  NOR2_X1 U10553 ( .A1(n9250), .A2(n9249), .ZN(n9678) );
  MUX2_X1 U10554 ( .A(n9615), .B(P1_REG1_REG_12__SCAN_IN), .S(n9675), .Z(n9677) );
  NOR2_X1 U10555 ( .A1(n9678), .A2(n9677), .ZN(n9676) );
  AOI21_X1 U10556 ( .B1(n9251), .B2(n9615), .A(n9676), .ZN(n9692) );
  MUX2_X1 U10557 ( .A(n9252), .B(P1_REG1_REG_13__SCAN_IN), .S(n9684), .Z(n9693) );
  NOR2_X1 U10558 ( .A1(n9692), .A2(n9693), .ZN(n9691) );
  AOI21_X1 U10559 ( .B1(n9253), .B2(n9252), .A(n9691), .ZN(n9706) );
  MUX2_X1 U10560 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9254), .S(n9255), .Z(n9707) );
  NOR2_X1 U10561 ( .A1(n9706), .A2(n9707), .ZN(n9705) );
  AOI21_X1 U10562 ( .B1(n9255), .B2(n9254), .A(n9705), .ZN(n9256) );
  NAND2_X1 U10563 ( .A1(n9716), .A2(n9256), .ZN(n9258) );
  XNOR2_X1 U10564 ( .A(n9257), .B(n9256), .ZN(n9718) );
  NAND2_X1 U10565 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9718), .ZN(n9717) );
  NAND2_X1 U10566 ( .A1(n9258), .A2(n9717), .ZN(n9731) );
  NAND2_X1 U10567 ( .A1(n9730), .A2(n9731), .ZN(n9729) );
  OAI21_X1 U10568 ( .B1(n9260), .B2(n9259), .A(n9729), .ZN(n9745) );
  NAND2_X1 U10569 ( .A1(n9746), .A2(n9745), .ZN(n9744) );
  OAI21_X1 U10570 ( .B1(n9262), .B2(n9261), .A(n9744), .ZN(n9763) );
  NOR2_X1 U10571 ( .A1(n9764), .A2(n9763), .ZN(n9762) );
  AOI21_X1 U10572 ( .B1(n9264), .B2(n9263), .A(n9762), .ZN(n9265) );
  XNOR2_X1 U10573 ( .A(n9265), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9267) );
  OAI22_X1 U10574 ( .A1(n9270), .A2(n9723), .B1(n9267), .B2(n9765), .ZN(n9266)
         );
  INV_X1 U10575 ( .A(n9266), .ZN(n9272) );
  INV_X1 U10576 ( .A(n9267), .ZN(n9268) );
  NOR2_X1 U10577 ( .A1(n9268), .A2(n9765), .ZN(n9269) );
  AOI211_X1 U10578 ( .C1(n9270), .C2(n9758), .A(n9753), .B(n9269), .ZN(n9271)
         );
  MUX2_X1 U10579 ( .A(n9272), .B(n9271), .S(n9349), .Z(n9274) );
  OAI211_X1 U10580 ( .C1(n9275), .C2(n9769), .A(n9274), .B(n9273), .ZN(
        P1_U3260) );
  XNOR2_X1 U10581 ( .A(n9276), .B(n9426), .ZN(n9429) );
  NOR2_X1 U10582 ( .A1(n9785), .A2(n9277), .ZN(n9279) );
  AOI211_X1 U10583 ( .C1(n9426), .C2(n9590), .A(n9279), .B(n9278), .ZN(n9280)
         );
  OAI21_X1 U10584 ( .B1(n9429), .B2(n9281), .A(n9280), .ZN(P1_U3261) );
  AOI21_X1 U10585 ( .B1(n9288), .B2(n9283), .A(n9282), .ZN(n9284) );
  INV_X1 U10586 ( .A(n9284), .ZN(n9437) );
  AOI22_X1 U10587 ( .A1(n9434), .A2(n9590), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9787), .ZN(n9300) );
  NOR2_X1 U10588 ( .A1(n9286), .A2(n9285), .ZN(n9289) );
  OAI21_X1 U10589 ( .B1(n9289), .B2(n9288), .A(n9287), .ZN(n9290) );
  INV_X1 U10590 ( .A(n9292), .ZN(n9295) );
  INV_X1 U10591 ( .A(n9293), .ZN(n9294) );
  AOI211_X1 U10592 ( .C1(n9434), .C2(n9295), .A(n9832), .B(n9294), .ZN(n9433)
         );
  NAND2_X1 U10593 ( .A1(n9433), .A2(n9778), .ZN(n9296) );
  OAI211_X1 U10594 ( .C1(n9776), .C2(n9297), .A(n9436), .B(n9296), .ZN(n9298)
         );
  NAND2_X1 U10595 ( .A1(n9298), .A2(n9785), .ZN(n9299) );
  OAI211_X1 U10596 ( .C1(n9437), .C2(n9425), .A(n9300), .B(n9299), .ZN(
        P1_U3263) );
  XNOR2_X1 U10597 ( .A(n9301), .B(n9309), .ZN(n9447) );
  INV_X1 U10598 ( .A(n9302), .ZN(n9327) );
  INV_X1 U10599 ( .A(n9303), .ZN(n9304) );
  AOI21_X1 U10600 ( .B1(n9443), .B2(n9327), .A(n9304), .ZN(n9444) );
  AOI22_X1 U10601 ( .A1(n9305), .A2(n9588), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9787), .ZN(n9306) );
  OAI21_X1 U10602 ( .B1(n9307), .B2(n9410), .A(n9306), .ZN(n9317) );
  INV_X1 U10603 ( .A(n9308), .ZN(n9311) );
  INV_X1 U10604 ( .A(n9309), .ZN(n9310) );
  AOI21_X1 U10605 ( .B1(n9311), .B2(n9310), .A(n5556), .ZN(n9315) );
  OAI22_X1 U10606 ( .A1(n9312), .A2(n9577), .B1(n9341), .B2(n5559), .ZN(n9313)
         );
  AOI21_X1 U10607 ( .B1(n9315), .B2(n9314), .A(n9313), .ZN(n9446) );
  NOR2_X1 U10608 ( .A1(n9446), .A2(n9787), .ZN(n9316) );
  AOI211_X1 U10609 ( .C1(n9401), .C2(n9444), .A(n9317), .B(n9316), .ZN(n9318)
         );
  OAI21_X1 U10610 ( .B1(n9447), .B2(n9425), .A(n9318), .ZN(P1_U3265) );
  XNOR2_X1 U10611 ( .A(n9319), .B(n9323), .ZN(n9322) );
  AOI222_X1 U10612 ( .A1(n9586), .A2(n9322), .B1(n9321), .B2(n9419), .C1(n9320), .C2(n9417), .ZN(n9451) );
  XNOR2_X1 U10613 ( .A(n9324), .B(n9323), .ZN(n9448) );
  NAND2_X1 U10614 ( .A1(n9448), .A2(n9599), .ZN(n9333) );
  OAI22_X1 U10615 ( .A1(n9326), .A2(n9776), .B1(n9325), .B2(n9785), .ZN(n9331)
         );
  INV_X1 U10616 ( .A(n5571), .ZN(n9328) );
  OAI211_X1 U10617 ( .C1(n9328), .C2(n4673), .A(n9327), .B(n9595), .ZN(n9449)
         );
  NOR2_X1 U10618 ( .A1(n9449), .A2(n9329), .ZN(n9330) );
  AOI211_X1 U10619 ( .C1(n9590), .C2(n5571), .A(n9331), .B(n9330), .ZN(n9332)
         );
  OAI211_X1 U10620 ( .C1(n9787), .C2(n9451), .A(n9333), .B(n9332), .ZN(
        P1_U3266) );
  XNOR2_X1 U10621 ( .A(n9335), .B(n9334), .ZN(n9453) );
  INV_X1 U10622 ( .A(n9453), .ZN(n9353) );
  AOI22_X1 U10623 ( .A1(n9344), .A2(n9590), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9787), .ZN(n9352) );
  NAND2_X1 U10624 ( .A1(n9337), .A2(n9336), .ZN(n9338) );
  AOI21_X1 U10625 ( .B1(n9339), .B2(n9338), .A(n5556), .ZN(n9343) );
  OAI22_X1 U10626 ( .A1(n9341), .A2(n9577), .B1(n9340), .B2(n5559), .ZN(n9342)
         );
  OR2_X1 U10627 ( .A1(n9343), .A2(n9342), .ZN(n9457) );
  AOI21_X1 U10628 ( .B1(n9345), .B2(n9344), .A(n9832), .ZN(n9347) );
  NAND2_X1 U10629 ( .A1(n9347), .A2(n9346), .ZN(n9454) );
  OAI22_X1 U10630 ( .A1(n9454), .A2(n9349), .B1(n9776), .B2(n9348), .ZN(n9350)
         );
  OAI21_X1 U10631 ( .B1(n9457), .B2(n9350), .A(n9785), .ZN(n9351) );
  OAI211_X1 U10632 ( .C1(n9353), .C2(n9425), .A(n9352), .B(n9351), .ZN(
        P1_U3267) );
  NAND2_X1 U10633 ( .A1(n9355), .A2(n9354), .ZN(n9356) );
  XNOR2_X1 U10634 ( .A(n9356), .B(n9362), .ZN(n9474) );
  AOI211_X1 U10635 ( .C1(n9471), .C2(n9372), .A(n9832), .B(n9357), .ZN(n9470)
         );
  INV_X1 U10636 ( .A(n9471), .ZN(n9361) );
  INV_X1 U10637 ( .A(n9358), .ZN(n9359) );
  AOI22_X1 U10638 ( .A1(n9787), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9359), .B2(
        n9588), .ZN(n9360) );
  OAI21_X1 U10639 ( .B1(n9361), .B2(n9410), .A(n9360), .ZN(n9369) );
  OAI21_X1 U10640 ( .B1(n4397), .B2(n9363), .A(n9362), .ZN(n9365) );
  NAND2_X1 U10641 ( .A1(n9365), .A2(n9364), .ZN(n9367) );
  AOI222_X1 U10642 ( .A1(n9586), .A2(n9367), .B1(n9366), .B2(n9417), .C1(n9396), .C2(n9419), .ZN(n9473) );
  NOR2_X1 U10643 ( .A1(n9473), .A2(n9787), .ZN(n9368) );
  AOI211_X1 U10644 ( .C1(n9470), .C2(n9598), .A(n9369), .B(n9368), .ZN(n9370)
         );
  OAI21_X1 U10645 ( .B1(n9425), .B2(n9474), .A(n9370), .ZN(P1_U3270) );
  XNOR2_X1 U10646 ( .A(n9371), .B(n9379), .ZN(n9479) );
  INV_X1 U10647 ( .A(n9372), .ZN(n9373) );
  AOI211_X1 U10648 ( .C1(n9476), .C2(n9388), .A(n9832), .B(n9373), .ZN(n9475)
         );
  INV_X1 U10649 ( .A(n9476), .ZN(n9377) );
  INV_X1 U10650 ( .A(n9374), .ZN(n9375) );
  AOI22_X1 U10651 ( .A1(n9787), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9375), .B2(
        n9588), .ZN(n9376) );
  OAI21_X1 U10652 ( .B1(n9377), .B2(n9410), .A(n9376), .ZN(n9385) );
  AOI211_X1 U10653 ( .C1(n9379), .C2(n9378), .A(n5556), .B(n4397), .ZN(n9383)
         );
  OAI22_X1 U10654 ( .A1(n9381), .A2(n9577), .B1(n9380), .B2(n5559), .ZN(n9382)
         );
  NOR2_X1 U10655 ( .A1(n9383), .A2(n9382), .ZN(n9478) );
  NOR2_X1 U10656 ( .A1(n9478), .A2(n9787), .ZN(n9384) );
  AOI211_X1 U10657 ( .C1(n9475), .C2(n9598), .A(n9385), .B(n9384), .ZN(n9386)
         );
  OAI21_X1 U10658 ( .B1(n9425), .B2(n9479), .A(n9386), .ZN(P1_U3271) );
  XOR2_X1 U10659 ( .A(n9387), .B(n9394), .Z(n9484) );
  INV_X1 U10660 ( .A(n9406), .ZN(n9390) );
  INV_X1 U10661 ( .A(n9388), .ZN(n9389) );
  AOI21_X1 U10662 ( .B1(n9480), .B2(n9390), .A(n9389), .ZN(n9481) );
  AOI22_X1 U10663 ( .A1(n9787), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9391), .B2(
        n9588), .ZN(n9392) );
  OAI21_X1 U10664 ( .B1(n9393), .B2(n9410), .A(n9392), .ZN(n9400) );
  XNOR2_X1 U10665 ( .A(n9395), .B(n9394), .ZN(n9398) );
  AOI222_X1 U10666 ( .A1(n9586), .A2(n9398), .B1(n9397), .B2(n9419), .C1(n9396), .C2(n9417), .ZN(n9483) );
  NOR2_X1 U10667 ( .A1(n9483), .A2(n9787), .ZN(n9399) );
  AOI211_X1 U10668 ( .C1(n9481), .C2(n9401), .A(n9400), .B(n9399), .ZN(n9402)
         );
  OAI21_X1 U10669 ( .B1(n9484), .B2(n9425), .A(n9402), .ZN(P1_U3272) );
  OAI21_X1 U10670 ( .B1(n4858), .B2(n9412), .A(n9404), .ZN(n9489) );
  AOI211_X1 U10671 ( .C1(n9486), .C2(n4672), .A(n9832), .B(n9406), .ZN(n9485)
         );
  INV_X1 U10672 ( .A(n9407), .ZN(n9408) );
  AOI22_X1 U10673 ( .A1(n9787), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9408), .B2(
        n9588), .ZN(n9409) );
  OAI21_X1 U10674 ( .B1(n9411), .B2(n9410), .A(n9409), .ZN(n9423) );
  OAI21_X1 U10675 ( .B1(n9414), .B2(n9413), .A(n9412), .ZN(n9416) );
  NAND2_X1 U10676 ( .A1(n9416), .A2(n9415), .ZN(n9421) );
  AOI222_X1 U10677 ( .A1(n9586), .A2(n9421), .B1(n9420), .B2(n9419), .C1(n9418), .C2(n9417), .ZN(n9488) );
  NOR2_X1 U10678 ( .A1(n9488), .A2(n9787), .ZN(n9422) );
  AOI211_X1 U10679 ( .C1(n9485), .C2(n9598), .A(n9423), .B(n9422), .ZN(n9424)
         );
  OAI21_X1 U10680 ( .B1(n9425), .B2(n9489), .A(n9424), .ZN(P1_U3273) );
  NAND2_X1 U10681 ( .A1(n9426), .A2(n9500), .ZN(n9427) );
  OAI211_X1 U10682 ( .C1(n9429), .C2(n9832), .A(n9428), .B(n9427), .ZN(n9514)
         );
  MUX2_X1 U10683 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9514), .S(n9852), .Z(
        P1_U3554) );
  INV_X2 U10684 ( .A(n9849), .ZN(n9852) );
  MUX2_X1 U10685 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9515), .S(n9852), .Z(
        P1_U3552) );
  AOI21_X1 U10686 ( .B1(n9434), .B2(n9500), .A(n9433), .ZN(n9435) );
  MUX2_X1 U10687 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9516), .S(n9852), .Z(
        P1_U3551) );
  AOI22_X1 U10688 ( .A1(n9439), .A2(n9595), .B1(n9438), .B2(n9500), .ZN(n9440)
         );
  OAI211_X1 U10689 ( .C1(n9442), .C2(n9505), .A(n9441), .B(n9440), .ZN(n9517)
         );
  MUX2_X1 U10690 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9517), .S(n9852), .Z(
        P1_U3550) );
  AOI22_X1 U10691 ( .A1(n9444), .A2(n9595), .B1(n9443), .B2(n9500), .ZN(n9445)
         );
  OAI211_X1 U10692 ( .C1(n9447), .C2(n9505), .A(n9446), .B(n9445), .ZN(n9518)
         );
  MUX2_X1 U10693 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9518), .S(n9852), .Z(
        P1_U3549) );
  NAND2_X1 U10694 ( .A1(n9448), .A2(n9827), .ZN(n9452) );
  NAND4_X1 U10695 ( .A1(n9452), .A2(n9451), .A3(n9450), .A4(n9449), .ZN(n9519)
         );
  MUX2_X1 U10696 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9519), .S(n9852), .Z(
        P1_U3548) );
  NAND2_X1 U10697 ( .A1(n9453), .A2(n9827), .ZN(n9459) );
  OAI21_X1 U10698 ( .B1(n9455), .B2(n9831), .A(n9454), .ZN(n9456) );
  NOR2_X1 U10699 ( .A1(n9457), .A2(n9456), .ZN(n9458) );
  NAND2_X1 U10700 ( .A1(n9459), .A2(n9458), .ZN(n9520) );
  MUX2_X1 U10701 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9520), .S(n9852), .Z(
        P1_U3547) );
  AOI22_X1 U10702 ( .A1(n9461), .A2(n9595), .B1(n9460), .B2(n9500), .ZN(n9462)
         );
  OAI211_X1 U10703 ( .C1(n9464), .C2(n9505), .A(n9463), .B(n9462), .ZN(n9521)
         );
  MUX2_X1 U10704 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9521), .S(n9852), .Z(
        P1_U3546) );
  AOI22_X1 U10705 ( .A1(n9466), .A2(n9595), .B1(n9465), .B2(n9500), .ZN(n9467)
         );
  OAI211_X1 U10706 ( .C1(n9469), .C2(n9505), .A(n9468), .B(n9467), .ZN(n9522)
         );
  MUX2_X1 U10707 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9522), .S(n9852), .Z(
        P1_U3545) );
  AOI21_X1 U10708 ( .B1(n9471), .B2(n9500), .A(n9470), .ZN(n9472) );
  OAI211_X1 U10709 ( .C1(n9474), .C2(n9505), .A(n9473), .B(n9472), .ZN(n9523)
         );
  MUX2_X1 U10710 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9523), .S(n9852), .Z(
        P1_U3544) );
  AOI21_X1 U10711 ( .B1(n9476), .B2(n9500), .A(n9475), .ZN(n9477) );
  OAI211_X1 U10712 ( .C1(n9479), .C2(n9505), .A(n9478), .B(n9477), .ZN(n9524)
         );
  MUX2_X1 U10713 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9524), .S(n9852), .Z(
        P1_U3543) );
  AOI22_X1 U10714 ( .A1(n9481), .A2(n9595), .B1(n9480), .B2(n9500), .ZN(n9482)
         );
  OAI211_X1 U10715 ( .C1(n9484), .C2(n9505), .A(n9483), .B(n9482), .ZN(n9525)
         );
  MUX2_X1 U10716 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9525), .S(n9852), .Z(
        P1_U3542) );
  AOI21_X1 U10717 ( .B1(n9486), .B2(n9500), .A(n9485), .ZN(n9487) );
  OAI211_X1 U10718 ( .C1(n9489), .C2(n9505), .A(n9488), .B(n9487), .ZN(n9526)
         );
  MUX2_X1 U10719 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9526), .S(n9852), .Z(
        P1_U3541) );
  AOI22_X1 U10720 ( .A1(n9491), .A2(n9595), .B1(n9490), .B2(n9500), .ZN(n9492)
         );
  OAI211_X1 U10721 ( .C1(n9494), .C2(n9505), .A(n9493), .B(n9492), .ZN(n9527)
         );
  MUX2_X1 U10722 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9527), .S(n9852), .Z(
        P1_U3540) );
  AOI211_X1 U10723 ( .C1(n9497), .C2(n9500), .A(n9496), .B(n9495), .ZN(n9498)
         );
  OAI21_X1 U10724 ( .B1(n9499), .B2(n9505), .A(n9498), .ZN(n9528) );
  MUX2_X1 U10725 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9528), .S(n9852), .Z(
        P1_U3539) );
  AOI22_X1 U10726 ( .A1(n9502), .A2(n9595), .B1(n9501), .B2(n9500), .ZN(n9503)
         );
  OAI211_X1 U10727 ( .C1(n9506), .C2(n9505), .A(n9504), .B(n9503), .ZN(n9529)
         );
  MUX2_X1 U10728 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9529), .S(n9852), .Z(
        P1_U3536) );
  OAI22_X1 U10729 ( .A1(n9508), .A2(n9832), .B1(n9507), .B2(n9831), .ZN(n9509)
         );
  AOI21_X1 U10730 ( .B1(n9510), .B2(n9837), .A(n9509), .ZN(n9511) );
  NAND2_X1 U10731 ( .A1(n9512), .A2(n9511), .ZN(n9530) );
  MUX2_X1 U10732 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9530), .S(n9852), .Z(
        P1_U3534) );
  MUX2_X1 U10733 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9513), .S(n9852), .Z(
        P1_U3523) );
  MUX2_X1 U10734 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9514), .S(n9840), .Z(
        P1_U3522) );
  MUX2_X1 U10735 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9515), .S(n9840), .Z(
        P1_U3520) );
  MUX2_X1 U10736 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9516), .S(n9840), .Z(
        P1_U3519) );
  MUX2_X1 U10737 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9517), .S(n9840), .Z(
        P1_U3518) );
  MUX2_X1 U10738 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9518), .S(n9840), .Z(
        P1_U3517) );
  MUX2_X1 U10739 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9519), .S(n9840), .Z(
        P1_U3516) );
  MUX2_X1 U10740 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9520), .S(n9840), .Z(
        P1_U3515) );
  MUX2_X1 U10741 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9521), .S(n9840), .Z(
        P1_U3514) );
  MUX2_X1 U10742 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9522), .S(n9840), .Z(
        P1_U3513) );
  MUX2_X1 U10743 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9523), .S(n9840), .Z(
        P1_U3512) );
  MUX2_X1 U10744 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9524), .S(n9840), .Z(
        P1_U3511) );
  MUX2_X1 U10745 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9525), .S(n9840), .Z(
        P1_U3510) );
  MUX2_X1 U10746 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9526), .S(n9840), .Z(
        P1_U3508) );
  MUX2_X1 U10747 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9527), .S(n9840), .Z(
        P1_U3505) );
  MUX2_X1 U10748 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9528), .S(n9840), .Z(
        P1_U3502) );
  MUX2_X1 U10749 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9529), .S(n9840), .Z(
        P1_U3493) );
  MUX2_X1 U10750 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n9530), .S(n9840), .Z(
        P1_U3487) );
  NAND2_X1 U10751 ( .A1(n10247), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9532) );
  OAI22_X1 U10752 ( .A1(n9533), .A2(n9532), .B1(n6598), .B2(n9531), .ZN(n9534)
         );
  AOI21_X1 U10753 ( .B1(n8298), .B2(n9535), .A(n9534), .ZN(n9536) );
  INV_X1 U10754 ( .A(n9536), .ZN(P1_U3322) );
  MUX2_X1 U10755 ( .A(n9537), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10756 ( .A1(n9854), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9548) );
  AOI211_X1 U10757 ( .C1(n9540), .C2(n9539), .A(n9538), .B(n9549), .ZN(n9541)
         );
  AOI21_X1 U10758 ( .B1(n9555), .B2(n9542), .A(n9541), .ZN(n9547) );
  AND2_X1 U10759 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9545) );
  OAI211_X1 U10760 ( .C1(n9545), .C2(n9544), .A(n9853), .B(n9543), .ZN(n9546)
         );
  NAND3_X1 U10761 ( .A1(n9548), .A2(n9547), .A3(n9546), .ZN(P2_U3246) );
  AOI22_X1 U10762 ( .A1(n9854), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9561) );
  AOI211_X1 U10763 ( .C1(n9552), .C2(n9551), .A(n9550), .B(n9549), .ZN(n9553)
         );
  AOI21_X1 U10764 ( .B1(n9555), .B2(n9554), .A(n9553), .ZN(n9560) );
  OAI211_X1 U10765 ( .C1(n9558), .C2(n9557), .A(n9853), .B(n9556), .ZN(n9559)
         );
  NAND3_X1 U10766 ( .A1(n9561), .A2(n9560), .A3(n9559), .ZN(P2_U3247) );
  OAI211_X1 U10767 ( .C1(n9564), .C2(n9831), .A(n9563), .B(n9562), .ZN(n9565)
         );
  AOI21_X1 U10768 ( .B1(n9827), .B2(n9566), .A(n9565), .ZN(n9567) );
  AOI22_X1 U10769 ( .A1(n9840), .A2(n9567), .B1(n5166), .B2(n9838), .ZN(
        P1_U3484) );
  AOI22_X1 U10770 ( .A1(n9852), .A2(n9567), .B1(n5163), .B2(n9849), .ZN(
        P1_U3533) );
  OAI22_X1 U10771 ( .A1(n9569), .A2(n9927), .B1(n9568), .B2(n9925), .ZN(n9571)
         );
  AOI211_X1 U10772 ( .C1(n9572), .C2(n9931), .A(n9571), .B(n9570), .ZN(n9574)
         );
  AOI22_X1 U10773 ( .A1(n9947), .A2(n9574), .B1(n5956), .B2(n9945), .ZN(
        P2_U3534) );
  INV_X1 U10774 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9573) );
  AOI22_X1 U10775 ( .A1(n9935), .A2(n9574), .B1(n9573), .B2(n9933), .ZN(
        P2_U3493) );
  XNOR2_X1 U10776 ( .A(n9575), .B(n9580), .ZN(n9585) );
  OAI22_X1 U10777 ( .A1(n9578), .A2(n9577), .B1(n9576), .B2(n5559), .ZN(n9584)
         );
  OAI21_X1 U10778 ( .B1(n9581), .B2(n9580), .A(n9579), .ZN(n9591) );
  NOR2_X1 U10779 ( .A1(n9591), .A2(n9582), .ZN(n9583) );
  AOI211_X1 U10780 ( .C1(n9586), .C2(n9585), .A(n9584), .B(n9583), .ZN(n9611)
         );
  INV_X1 U10781 ( .A(n9587), .ZN(n9589) );
  AOI222_X1 U10782 ( .A1(n9593), .A2(n9590), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n9787), .C1(n9589), .C2(n9588), .ZN(n9601) );
  INV_X1 U10783 ( .A(n9591), .ZN(n9614) );
  INV_X1 U10784 ( .A(n9592), .ZN(n9596) );
  INV_X1 U10785 ( .A(n9593), .ZN(n9610) );
  OAI211_X1 U10786 ( .C1(n9596), .C2(n9610), .A(n9595), .B(n9594), .ZN(n9609)
         );
  INV_X1 U10787 ( .A(n9609), .ZN(n9597) );
  AOI22_X1 U10788 ( .A1(n9614), .A2(n9599), .B1(n9598), .B2(n9597), .ZN(n9600)
         );
  OAI211_X1 U10789 ( .C1(n9787), .C2(n9611), .A(n9601), .B(n9600), .ZN(
        P1_U3279) );
  INV_X1 U10790 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9602) );
  AOI22_X1 U10791 ( .A1(n9852), .A2(n9603), .B1(n9602), .B2(n9849), .ZN(
        P1_U3553) );
  OAI21_X1 U10792 ( .B1(n9605), .B2(n9831), .A(n9604), .ZN(n9606) );
  AOI211_X1 U10793 ( .C1(n9608), .C2(n9827), .A(n9607), .B(n9606), .ZN(n9616)
         );
  AOI22_X1 U10794 ( .A1(n9852), .A2(n9616), .B1(n9254), .B2(n9849), .ZN(
        P1_U3537) );
  OAI21_X1 U10795 ( .B1(n9610), .B2(n9831), .A(n9609), .ZN(n9613) );
  INV_X1 U10796 ( .A(n9611), .ZN(n9612) );
  AOI211_X1 U10797 ( .C1(n9837), .C2(n9614), .A(n9613), .B(n9612), .ZN(n9618)
         );
  AOI22_X1 U10798 ( .A1(n9852), .A2(n9618), .B1(n9615), .B2(n9849), .ZN(
        P1_U3535) );
  AOI22_X1 U10799 ( .A1(n9840), .A2(n9616), .B1(n5253), .B2(n9838), .ZN(
        P1_U3496) );
  INV_X1 U10800 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9617) );
  AOI22_X1 U10801 ( .A1(n9840), .A2(n9618), .B1(n9617), .B2(n9838), .ZN(
        P1_U3490) );
  XNOR2_X1 U10802 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  AOI21_X1 U10803 ( .B1(n9619), .B2(n10045), .A(P1_IR_REG_0__SCAN_IN), .ZN(
        n9620) );
  OAI21_X1 U10804 ( .B1(n9621), .B2(n9620), .A(n5026), .ZN(n9622) );
  NOR3_X1 U10805 ( .A1(n9624), .A2(n9623), .A3(n9622), .ZN(n9626) );
  NOR3_X1 U10806 ( .A1(n9765), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n10074), .ZN(
        n9625) );
  AOI211_X1 U10807 ( .C1(P1_ADDR_REG_0__SCAN_IN), .C2(n9655), .A(n9626), .B(
        n9625), .ZN(n9627) );
  OAI21_X1 U10808 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7126), .A(n9627), .ZN(
        P1_U3241) );
  AOI22_X1 U10809 ( .A1(n9753), .A2(n9628), .B1(n9655), .B2(
        P1_ADDR_REG_2__SCAN_IN), .ZN(n9636) );
  MUX2_X1 U10810 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6512), .S(n9629), .Z(n9632)
         );
  NAND3_X1 U10811 ( .A1(n9632), .A2(n9631), .A3(n9630), .ZN(n9633) );
  NAND3_X1 U10812 ( .A1(n9758), .A2(n9634), .A3(n9633), .ZN(n9635) );
  AND3_X1 U10813 ( .A1(n9637), .A2(n9636), .A3(n9635), .ZN(n9642) );
  INV_X1 U10814 ( .A(n9765), .ZN(n9743) );
  OAI211_X1 U10815 ( .C1(n9640), .C2(n9639), .A(n9743), .B(n9638), .ZN(n9641)
         );
  OAI211_X1 U10816 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n4631), .A(n9642), .B(
        n9641), .ZN(P1_U3243) );
  AOI22_X1 U10817 ( .A1(n9753), .A2(n9643), .B1(n9655), .B2(
        P1_ADDR_REG_5__SCAN_IN), .ZN(n9654) );
  AOI21_X1 U10818 ( .B1(n9646), .B2(n9645), .A(n9644), .ZN(n9647) );
  OR2_X1 U10819 ( .A1(n9723), .A2(n9647), .ZN(n9652) );
  OAI211_X1 U10820 ( .C1(n9650), .C2(n9649), .A(n9743), .B(n9648), .ZN(n9651)
         );
  NAND4_X1 U10821 ( .A1(n9654), .A2(n9653), .A3(n9652), .A4(n9651), .ZN(
        P1_U3246) );
  AOI22_X1 U10822 ( .A1(n9753), .A2(n9656), .B1(n9655), .B2(
        P1_ADDR_REG_8__SCAN_IN), .ZN(n9669) );
  INV_X1 U10823 ( .A(n9657), .ZN(n9668) );
  MUX2_X1 U10824 ( .A(n9659), .B(P1_REG2_REG_8__SCAN_IN), .S(n9658), .Z(n9661)
         );
  AOI21_X1 U10825 ( .B1(n9662), .B2(n9661), .A(n9723), .ZN(n9660) );
  OAI21_X1 U10826 ( .B1(n9662), .B2(n9661), .A(n9660), .ZN(n9667) );
  OAI211_X1 U10827 ( .C1(n9665), .C2(n9664), .A(n9743), .B(n9663), .ZN(n9666)
         );
  NAND4_X1 U10828 ( .A1(n9669), .A2(n9668), .A3(n9667), .A4(n9666), .ZN(
        P1_U3249) );
  INV_X1 U10829 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9682) );
  AOI211_X1 U10830 ( .C1(n9672), .C2(n9671), .A(n9670), .B(n9723), .ZN(n9673)
         );
  AOI211_X1 U10831 ( .C1(n9753), .C2(n9675), .A(n9674), .B(n9673), .ZN(n9681)
         );
  AOI21_X1 U10832 ( .B1(n9678), .B2(n9677), .A(n9676), .ZN(n9679) );
  OR2_X1 U10833 ( .A1(n9679), .A2(n9765), .ZN(n9680) );
  OAI211_X1 U10834 ( .C1(n9682), .C2(n9769), .A(n9681), .B(n9680), .ZN(
        P1_U3253) );
  INV_X1 U10835 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9697) );
  AOI21_X1 U10836 ( .B1(n9753), .B2(n9684), .A(n9683), .ZN(n9690) );
  AOI21_X1 U10837 ( .B1(n9687), .B2(n9686), .A(n9685), .ZN(n9688) );
  NAND2_X1 U10838 ( .A1(n9758), .A2(n9688), .ZN(n9689) );
  AND2_X1 U10839 ( .A1(n9690), .A2(n9689), .ZN(n9696) );
  AOI21_X1 U10840 ( .B1(n9693), .B2(n9692), .A(n9691), .ZN(n9694) );
  OR2_X1 U10841 ( .A1(n9765), .A2(n9694), .ZN(n9695) );
  OAI211_X1 U10842 ( .C1(n9697), .C2(n9769), .A(n9696), .B(n9695), .ZN(
        P1_U3254) );
  INV_X1 U10843 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9711) );
  AOI21_X1 U10844 ( .B1(n9753), .B2(n9699), .A(n9698), .ZN(n9704) );
  AOI21_X1 U10845 ( .B1(n9701), .B2(n7749), .A(n9700), .ZN(n9702) );
  NAND2_X1 U10846 ( .A1(n9758), .A2(n9702), .ZN(n9703) );
  AND2_X1 U10847 ( .A1(n9704), .A2(n9703), .ZN(n9710) );
  AOI21_X1 U10848 ( .B1(n9707), .B2(n9706), .A(n9705), .ZN(n9708) );
  OR2_X1 U10849 ( .A1(n9765), .A2(n9708), .ZN(n9709) );
  OAI211_X1 U10850 ( .C1(n9711), .C2(n9769), .A(n9710), .B(n9709), .ZN(
        P1_U3255) );
  INV_X1 U10851 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9721) );
  AOI211_X1 U10852 ( .C1(n9713), .C2(n5283), .A(n9712), .B(n9723), .ZN(n9714)
         );
  AOI211_X1 U10853 ( .C1(n9753), .C2(n9716), .A(n9715), .B(n9714), .ZN(n9720)
         );
  OAI211_X1 U10854 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9718), .A(n9743), .B(
        n9717), .ZN(n9719) );
  OAI211_X1 U10855 ( .C1(n9721), .C2(n9769), .A(n9720), .B(n9719), .ZN(
        P1_U3256) );
  INV_X1 U10856 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9734) );
  INV_X1 U10857 ( .A(n9722), .ZN(n9727) );
  AOI211_X1 U10858 ( .C1(n4419), .C2(n9725), .A(n9724), .B(n9723), .ZN(n9726)
         );
  AOI211_X1 U10859 ( .C1(n9753), .C2(n9728), .A(n9727), .B(n9726), .ZN(n9733)
         );
  OAI211_X1 U10860 ( .C1(n9731), .C2(n9730), .A(n9743), .B(n9729), .ZN(n9732)
         );
  OAI211_X1 U10861 ( .C1(n9734), .C2(n9769), .A(n9733), .B(n9732), .ZN(
        P1_U3257) );
  INV_X1 U10862 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9749) );
  AOI21_X1 U10863 ( .B1(n9737), .B2(n9736), .A(n9735), .ZN(n9738) );
  NAND2_X1 U10864 ( .A1(n9758), .A2(n9738), .ZN(n9742) );
  NAND2_X1 U10865 ( .A1(n9753), .A2(n9739), .ZN(n9741) );
  AND3_X1 U10866 ( .A1(n9742), .A2(n9741), .A3(n9740), .ZN(n9748) );
  OAI211_X1 U10867 ( .C1(n9746), .C2(n9745), .A(n9744), .B(n9743), .ZN(n9747)
         );
  OAI211_X1 U10868 ( .C1(n9749), .C2(n9769), .A(n9748), .B(n9747), .ZN(
        P1_U3258) );
  INV_X1 U10869 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9770) );
  INV_X1 U10870 ( .A(n9750), .ZN(n9751) );
  AOI21_X1 U10871 ( .B1(n9753), .B2(n9752), .A(n9751), .ZN(n9761) );
  NAND2_X1 U10872 ( .A1(n9755), .A2(n9754), .ZN(n9759) );
  INV_X1 U10873 ( .A(n9756), .ZN(n9757) );
  NAND3_X1 U10874 ( .A1(n9759), .A2(n9758), .A3(n9757), .ZN(n9760) );
  AND2_X1 U10875 ( .A1(n9761), .A2(n9760), .ZN(n9768) );
  AOI21_X1 U10876 ( .B1(n9764), .B2(n9763), .A(n9762), .ZN(n9766) );
  OR2_X1 U10877 ( .A1(n9766), .A2(n9765), .ZN(n9767) );
  OAI211_X1 U10878 ( .C1(n9770), .C2(n9769), .A(n9768), .B(n9767), .ZN(
        P1_U3259) );
  INV_X1 U10879 ( .A(n9771), .ZN(n9783) );
  NAND2_X1 U10880 ( .A1(n9773), .A2(n9772), .ZN(n9774) );
  OAI21_X1 U10881 ( .B1(n9776), .B2(n9775), .A(n9774), .ZN(n9777) );
  AOI21_X1 U10882 ( .B1(n9779), .B2(n9778), .A(n9777), .ZN(n9780) );
  OAI211_X1 U10883 ( .C1(n9783), .C2(n9782), .A(n9781), .B(n9780), .ZN(n9784)
         );
  INV_X1 U10884 ( .A(n9784), .ZN(n9786) );
  AOI22_X1 U10885 ( .A1(n9787), .A2(n6518), .B1(n9786), .B2(n9785), .ZN(
        P1_U3286) );
  NOR2_X1 U10886 ( .A1(n9789), .A2(n10162), .ZN(P1_U3292) );
  AND2_X1 U10887 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9790), .ZN(P1_U3293) );
  AND2_X1 U10888 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9790), .ZN(P1_U3294) );
  AND2_X1 U10889 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9790), .ZN(P1_U3295) );
  INV_X1 U10890 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9991) );
  NOR2_X1 U10891 ( .A1(n9789), .A2(n9991), .ZN(P1_U3296) );
  NOR2_X1 U10892 ( .A1(n9789), .A2(n9788), .ZN(P1_U3297) );
  INV_X1 U10893 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10125) );
  NOR2_X1 U10894 ( .A1(n9789), .A2(n10125), .ZN(P1_U3298) );
  AND2_X1 U10895 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9790), .ZN(P1_U3299) );
  AND2_X1 U10896 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9790), .ZN(P1_U3300) );
  AND2_X1 U10897 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9790), .ZN(P1_U3301) );
  INV_X1 U10898 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10178) );
  NOR2_X1 U10899 ( .A1(n9789), .A2(n10178), .ZN(P1_U3302) );
  AND2_X1 U10900 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9790), .ZN(P1_U3303) );
  AND2_X1 U10901 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9790), .ZN(P1_U3304) );
  AND2_X1 U10902 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9790), .ZN(P1_U3305) );
  AND2_X1 U10903 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9790), .ZN(P1_U3306) );
  INV_X1 U10904 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10034) );
  NOR2_X1 U10905 ( .A1(n9789), .A2(n10034), .ZN(P1_U3307) );
  NOR2_X1 U10906 ( .A1(n9789), .A2(n10172), .ZN(P1_U3308) );
  AND2_X1 U10907 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9790), .ZN(P1_U3309) );
  AND2_X1 U10908 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9790), .ZN(P1_U3310) );
  AND2_X1 U10909 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9790), .ZN(P1_U3311) );
  AND2_X1 U10910 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9790), .ZN(P1_U3312) );
  INV_X1 U10911 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10184) );
  NOR2_X1 U10912 ( .A1(n9789), .A2(n10184), .ZN(P1_U3313) );
  AND2_X1 U10913 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9790), .ZN(P1_U3314) );
  NOR2_X1 U10914 ( .A1(n9789), .A2(n10062), .ZN(P1_U3315) );
  INV_X1 U10915 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10061) );
  NOR2_X1 U10916 ( .A1(n9789), .A2(n10061), .ZN(P1_U3316) );
  INV_X1 U10917 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10185) );
  NOR2_X1 U10918 ( .A1(n9789), .A2(n10185), .ZN(P1_U3317) );
  NOR2_X1 U10919 ( .A1(n9789), .A2(n10016), .ZN(P1_U3318) );
  INV_X1 U10920 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10103) );
  NOR2_X1 U10921 ( .A1(n9789), .A2(n10103), .ZN(P1_U3319) );
  AND2_X1 U10922 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9790), .ZN(P1_U3320) );
  AND2_X1 U10923 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9790), .ZN(P1_U3321) );
  INV_X1 U10924 ( .A(n9791), .ZN(n9792) );
  NAND2_X1 U10925 ( .A1(n9792), .A2(n9794), .ZN(n9793) );
  OAI21_X1 U10926 ( .B1(n9794), .B2(n5606), .A(n9793), .ZN(P1_U3441) );
  INV_X1 U10927 ( .A(n9795), .ZN(n9800) );
  OAI22_X1 U10928 ( .A1(n9797), .A2(n9832), .B1(n9796), .B2(n9831), .ZN(n9799)
         );
  AOI211_X1 U10929 ( .C1(n9837), .C2(n9800), .A(n9799), .B(n9798), .ZN(n9841)
         );
  AOI22_X1 U10930 ( .A1(n9840), .A2(n9841), .B1(n5007), .B2(n9838), .ZN(
        P1_U3460) );
  OAI22_X1 U10931 ( .A1(n9802), .A2(n9832), .B1(n9801), .B2(n9831), .ZN(n9804)
         );
  AOI211_X1 U10932 ( .C1(n9837), .C2(n9805), .A(n9804), .B(n9803), .ZN(n9842)
         );
  INV_X1 U10933 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10002) );
  AOI22_X1 U10934 ( .A1(n9840), .A2(n9842), .B1(n10002), .B2(n9838), .ZN(
        P1_U3463) );
  NAND2_X1 U10935 ( .A1(n9807), .A2(n9806), .ZN(n9809) );
  AOI211_X1 U10936 ( .C1(n9837), .C2(n9810), .A(n9809), .B(n9808), .ZN(n9843)
         );
  INV_X1 U10937 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9811) );
  AOI22_X1 U10938 ( .A1(n9840), .A2(n9843), .B1(n9811), .B2(n9838), .ZN(
        P1_U3466) );
  OAI22_X1 U10939 ( .A1(n9813), .A2(n9832), .B1(n9812), .B2(n9831), .ZN(n9815)
         );
  AOI211_X1 U10940 ( .C1(n9816), .C2(n9827), .A(n9815), .B(n9814), .ZN(n9844)
         );
  INV_X1 U10941 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9983) );
  AOI22_X1 U10942 ( .A1(n9840), .A2(n9844), .B1(n9983), .B2(n9838), .ZN(
        P1_U3472) );
  OAI211_X1 U10943 ( .C1(n9819), .C2(n9831), .A(n9818), .B(n9817), .ZN(n9820)
         );
  AOI21_X1 U10944 ( .B1(n9827), .B2(n9821), .A(n9820), .ZN(n9846) );
  INV_X1 U10945 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9822) );
  AOI22_X1 U10946 ( .A1(n9840), .A2(n9846), .B1(n9822), .B2(n9838), .ZN(
        P1_U3475) );
  OAI22_X1 U10947 ( .A1(n9824), .A2(n9832), .B1(n9823), .B2(n9831), .ZN(n9826)
         );
  AOI211_X1 U10948 ( .C1(n9828), .C2(n9827), .A(n9826), .B(n9825), .ZN(n9848)
         );
  INV_X1 U10949 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10064) );
  AOI22_X1 U10950 ( .A1(n9840), .A2(n9848), .B1(n10064), .B2(n9838), .ZN(
        P1_U3478) );
  INV_X1 U10951 ( .A(n9829), .ZN(n9836) );
  OAI22_X1 U10952 ( .A1(n9833), .A2(n9832), .B1(n4666), .B2(n9831), .ZN(n9835)
         );
  AOI211_X1 U10953 ( .C1(n9837), .C2(n9836), .A(n9835), .B(n9834), .ZN(n9851)
         );
  INV_X1 U10954 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9839) );
  AOI22_X1 U10955 ( .A1(n9840), .A2(n9851), .B1(n9839), .B2(n9838), .ZN(
        P1_U3481) );
  AOI22_X1 U10956 ( .A1(n9852), .A2(n9841), .B1(n6530), .B2(n9849), .ZN(
        P1_U3525) );
  AOI22_X1 U10957 ( .A1(n9852), .A2(n9842), .B1(n6535), .B2(n9849), .ZN(
        P1_U3526) );
  AOI22_X1 U10958 ( .A1(n9852), .A2(n9843), .B1(n6536), .B2(n9849), .ZN(
        P1_U3527) );
  AOI22_X1 U10959 ( .A1(n9852), .A2(n9844), .B1(n6528), .B2(n9849), .ZN(
        P1_U3529) );
  AOI22_X1 U10960 ( .A1(n9852), .A2(n9846), .B1(n9845), .B2(n9849), .ZN(
        P1_U3530) );
  AOI22_X1 U10961 ( .A1(n9852), .A2(n9848), .B1(n9847), .B2(n9849), .ZN(
        P1_U3531) );
  AOI22_X1 U10962 ( .A1(n9852), .A2(n9851), .B1(n9850), .B2(n9849), .ZN(
        P1_U3532) );
  AOI22_X1 U10963 ( .A1(n9856), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9853), .ZN(n9863) );
  AOI22_X1 U10964 ( .A1(n9854), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9862) );
  NAND2_X1 U10965 ( .A1(n9856), .A2(n9855), .ZN(n9858) );
  OAI211_X1 U10966 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n9859), .A(n9858), .B(
        n9857), .ZN(n9860) );
  NAND2_X1 U10967 ( .A1(n9860), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9861) );
  OAI211_X1 U10968 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9863), .A(n9862), .B(
        n9861), .ZN(P2_U3245) );
  NOR2_X1 U10969 ( .A1(n9865), .A2(n9864), .ZN(n9866) );
  AND2_X1 U10970 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9868), .ZN(P2_U3297) );
  AND2_X1 U10971 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9868), .ZN(P2_U3298) );
  AND2_X1 U10972 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9868), .ZN(P2_U3299) );
  AND2_X1 U10973 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9868), .ZN(P2_U3300) );
  AND2_X1 U10974 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9868), .ZN(P2_U3301) );
  AND2_X1 U10975 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9868), .ZN(P2_U3302) );
  INV_X1 U10976 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10150) );
  NOR2_X1 U10977 ( .A1(n9866), .A2(n10150), .ZN(P2_U3303) );
  AND2_X1 U10978 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9868), .ZN(P2_U3304) );
  AND2_X1 U10979 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9868), .ZN(P2_U3305) );
  AND2_X1 U10980 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9868), .ZN(P2_U3306) );
  INV_X1 U10981 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10130) );
  NOR2_X1 U10982 ( .A1(n9866), .A2(n10130), .ZN(P2_U3307) );
  AND2_X1 U10983 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9868), .ZN(P2_U3308) );
  AND2_X1 U10984 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9868), .ZN(P2_U3309) );
  AND2_X1 U10985 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9868), .ZN(P2_U3310) );
  AND2_X1 U10986 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9868), .ZN(P2_U3311) );
  AND2_X1 U10987 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9868), .ZN(P2_U3312) );
  AND2_X1 U10988 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9868), .ZN(P2_U3313) );
  AND2_X1 U10989 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9868), .ZN(P2_U3314) );
  INV_X1 U10990 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10031) );
  NOR2_X1 U10991 ( .A1(n9866), .A2(n10031), .ZN(P2_U3315) );
  AND2_X1 U10992 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9868), .ZN(P2_U3316) );
  AND2_X1 U10993 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9868), .ZN(P2_U3317) );
  AND2_X1 U10994 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9868), .ZN(P2_U3318) );
  AND2_X1 U10995 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9868), .ZN(P2_U3319) );
  AND2_X1 U10996 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9868), .ZN(P2_U3320) );
  AND2_X1 U10997 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9868), .ZN(P2_U3321) );
  AND2_X1 U10998 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9868), .ZN(P2_U3322) );
  AND2_X1 U10999 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9868), .ZN(P2_U3323) );
  AND2_X1 U11000 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9868), .ZN(P2_U3324) );
  AND2_X1 U11001 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9868), .ZN(P2_U3325) );
  AND2_X1 U11002 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9868), .ZN(P2_U3326) );
  AOI22_X1 U11003 ( .A1(n9867), .A2(n9870), .B1(n10008), .B2(n9868), .ZN(
        P2_U3437) );
  AOI22_X1 U11004 ( .A1(n9871), .A2(n9870), .B1(n9869), .B2(n9868), .ZN(
        P2_U3438) );
  OAI22_X1 U11005 ( .A1(n9875), .A2(n9874), .B1(n9873), .B2(n9872), .ZN(n9876)
         );
  NOR2_X1 U11006 ( .A1(n9877), .A2(n9876), .ZN(n9936) );
  AOI22_X1 U11007 ( .A1(n9935), .A2(n9936), .B1(n5693), .B2(n9933), .ZN(
        P2_U3451) );
  OAI22_X1 U11008 ( .A1(n9878), .A2(n9927), .B1(n6833), .B2(n9925), .ZN(n9881)
         );
  INV_X1 U11009 ( .A(n9879), .ZN(n9880) );
  AOI211_X1 U11010 ( .C1(n9931), .C2(n9882), .A(n9881), .B(n9880), .ZN(n9937)
         );
  INV_X1 U11011 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9883) );
  AOI22_X1 U11012 ( .A1(n9935), .A2(n9937), .B1(n9883), .B2(n9933), .ZN(
        P2_U3454) );
  OAI21_X1 U11013 ( .B1(n9885), .B2(n9925), .A(n9884), .ZN(n9887) );
  AOI211_X1 U11014 ( .C1(n9931), .C2(n9888), .A(n9887), .B(n9886), .ZN(n9938)
         );
  INV_X1 U11015 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9889) );
  AOI22_X1 U11016 ( .A1(n9935), .A2(n9938), .B1(n9889), .B2(n9933), .ZN(
        P2_U3457) );
  INV_X1 U11017 ( .A(n9890), .ZN(n9895) );
  OAI22_X1 U11018 ( .A1(n9892), .A2(n9927), .B1(n9891), .B2(n9925), .ZN(n9894)
         );
  AOI211_X1 U11019 ( .C1(n9922), .C2(n9895), .A(n9894), .B(n9893), .ZN(n9939)
         );
  INV_X1 U11020 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9896) );
  AOI22_X1 U11021 ( .A1(n9935), .A2(n9939), .B1(n9896), .B2(n9933), .ZN(
        P2_U3460) );
  AOI22_X1 U11022 ( .A1(n9900), .A2(n9899), .B1(n9898), .B2(n9897), .ZN(n9903)
         );
  NAND2_X1 U11023 ( .A1(n9901), .A2(n9931), .ZN(n9902) );
  AND3_X1 U11024 ( .A1(n9904), .A2(n9903), .A3(n9902), .ZN(n9940) );
  INV_X1 U11025 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9905) );
  AOI22_X1 U11026 ( .A1(n9935), .A2(n9940), .B1(n9905), .B2(n9933), .ZN(
        P2_U3463) );
  OAI22_X1 U11027 ( .A1(n9906), .A2(n9927), .B1(n6944), .B2(n9925), .ZN(n9908)
         );
  AOI211_X1 U11028 ( .C1(n9909), .C2(n9931), .A(n9908), .B(n9907), .ZN(n9941)
         );
  AOI22_X1 U11029 ( .A1(n9935), .A2(n9941), .B1(n5824), .B2(n9933), .ZN(
        P2_U3469) );
  INV_X1 U11030 ( .A(n9910), .ZN(n9915) );
  OAI22_X1 U11031 ( .A1(n9912), .A2(n9927), .B1(n9911), .B2(n9925), .ZN(n9914)
         );
  AOI211_X1 U11032 ( .C1(n9922), .C2(n9915), .A(n9914), .B(n9913), .ZN(n9943)
         );
  AOI22_X1 U11033 ( .A1(n9935), .A2(n9943), .B1(n5857), .B2(n9933), .ZN(
        P2_U3475) );
  INV_X1 U11034 ( .A(n9916), .ZN(n9921) );
  OAI22_X1 U11035 ( .A1(n9918), .A2(n9927), .B1(n9917), .B2(n9925), .ZN(n9920)
         );
  AOI211_X1 U11036 ( .C1(n9922), .C2(n9921), .A(n9920), .B(n9919), .ZN(n9944)
         );
  INV_X1 U11037 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9923) );
  AOI22_X1 U11038 ( .A1(n9935), .A2(n9944), .B1(n9923), .B2(n9933), .ZN(
        P2_U3481) );
  INV_X1 U11039 ( .A(n9924), .ZN(n9926) );
  OAI22_X1 U11040 ( .A1(n9928), .A2(n9927), .B1(n9926), .B2(n9925), .ZN(n9930)
         );
  AOI211_X1 U11041 ( .C1(n9932), .C2(n9931), .A(n9930), .B(n9929), .ZN(n9946)
         );
  INV_X1 U11042 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9934) );
  AOI22_X1 U11043 ( .A1(n9935), .A2(n9946), .B1(n9934), .B2(n9933), .ZN(
        P2_U3487) );
  AOI22_X1 U11044 ( .A1(n9947), .A2(n9936), .B1(n5699), .B2(n9945), .ZN(
        P2_U3520) );
  AOI22_X1 U11045 ( .A1(n9947), .A2(n9937), .B1(n6726), .B2(n9945), .ZN(
        P2_U3521) );
  AOI22_X1 U11046 ( .A1(n9947), .A2(n9938), .B1(n6725), .B2(n9945), .ZN(
        P2_U3522) );
  AOI22_X1 U11047 ( .A1(n9947), .A2(n9939), .B1(n6724), .B2(n9945), .ZN(
        P2_U3523) );
  AOI22_X1 U11048 ( .A1(n9947), .A2(n9940), .B1(n6722), .B2(n9945), .ZN(
        P2_U3524) );
  AOI22_X1 U11049 ( .A1(n9947), .A2(n9941), .B1(n6787), .B2(n9945), .ZN(
        P2_U3526) );
  AOI22_X1 U11050 ( .A1(n9947), .A2(n9943), .B1(n9942), .B2(n9945), .ZN(
        P2_U3528) );
  AOI22_X1 U11051 ( .A1(n9947), .A2(n9944), .B1(n6992), .B2(n9945), .ZN(
        P2_U3530) );
  AOI22_X1 U11052 ( .A1(n9947), .A2(n9946), .B1(n7456), .B2(n9945), .ZN(
        P2_U3532) );
  INV_X1 U11053 ( .A(n9948), .ZN(n9949) );
  NAND2_X1 U11054 ( .A1(n9950), .A2(n9949), .ZN(n9951) );
  XNOR2_X1 U11055 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9951), .ZN(ADD_1071_U5) );
  INV_X1 U11056 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10076) );
  INV_X1 U11057 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9952) );
  AOI22_X1 U11058 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n10076), .B2(n9952), .ZN(ADD_1071_U46) );
  OAI21_X1 U11059 ( .B1(n9955), .B2(n9954), .A(n9953), .ZN(ADD_1071_U56) );
  OAI21_X1 U11060 ( .B1(n9958), .B2(n9957), .A(n9956), .ZN(ADD_1071_U57) );
  OAI21_X1 U11061 ( .B1(n9961), .B2(n9960), .A(n9959), .ZN(ADD_1071_U58) );
  OAI21_X1 U11062 ( .B1(n9964), .B2(n9963), .A(n9962), .ZN(ADD_1071_U59) );
  OAI21_X1 U11063 ( .B1(n9967), .B2(n9966), .A(n9965), .ZN(ADD_1071_U60) );
  OAI21_X1 U11064 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(ADD_1071_U61) );
  AOI21_X1 U11065 ( .B1(n9973), .B2(n9972), .A(n9971), .ZN(ADD_1071_U62) );
  AOI21_X1 U11066 ( .B1(n9976), .B2(n9975), .A(n9974), .ZN(ADD_1071_U63) );
  AOI22_X1 U11067 ( .A1(n9978), .A2(keyinput9), .B1(keyinput48), .B2(n6726), 
        .ZN(n9977) );
  OAI221_X1 U11068 ( .B1(n9978), .B2(keyinput9), .C1(n6726), .C2(keyinput48), 
        .A(n9977), .ZN(n9989) );
  AOI22_X1 U11069 ( .A1(n5857), .A2(keyinput123), .B1(n9980), .B2(keyinput4), 
        .ZN(n9979) );
  OAI221_X1 U11070 ( .B1(n5857), .B2(keyinput123), .C1(n9980), .C2(keyinput4), 
        .A(n9979), .ZN(n9988) );
  INV_X1 U11071 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9982) );
  AOI22_X1 U11072 ( .A1(n9983), .A2(keyinput91), .B1(n9982), .B2(keyinput61), 
        .ZN(n9981) );
  OAI221_X1 U11073 ( .B1(n9983), .B2(keyinput91), .C1(n9982), .C2(keyinput61), 
        .A(n9981), .ZN(n9987) );
  XNOR2_X1 U11074 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput95), .ZN(n9985) );
  XNOR2_X1 U11075 ( .A(P1_REG0_REG_22__SCAN_IN), .B(keyinput113), .ZN(n9984)
         );
  NAND2_X1 U11076 ( .A1(n9985), .A2(n9984), .ZN(n9986) );
  NOR4_X1 U11077 ( .A1(n9989), .A2(n9988), .A3(n9987), .A4(n9986), .ZN(n10029)
         );
  AOI22_X1 U11078 ( .A1(P1_U3084), .A2(keyinput53), .B1(keyinput103), .B2(
        n9991), .ZN(n9990) );
  OAI221_X1 U11079 ( .B1(P1_U3084), .B2(keyinput53), .C1(n9991), .C2(
        keyinput103), .A(n9990), .ZN(n10000) );
  AOI22_X1 U11080 ( .A1(n9993), .A2(keyinput46), .B1(keyinput38), .B2(n10257), 
        .ZN(n9992) );
  OAI221_X1 U11081 ( .B1(n9993), .B2(keyinput46), .C1(n10257), .C2(keyinput38), 
        .A(n9992), .ZN(n9999) );
  XNOR2_X1 U11082 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput112), .ZN(n9997) );
  XNOR2_X1 U11083 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput60), .ZN(n9996) );
  XNOR2_X1 U11084 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput67), .ZN(n9995) );
  XNOR2_X1 U11085 ( .A(keyinput68), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9994) );
  NAND4_X1 U11086 ( .A1(n9997), .A2(n9996), .A3(n9995), .A4(n9994), .ZN(n9998)
         );
  NOR3_X1 U11087 ( .A1(n10000), .A2(n9999), .A3(n9998), .ZN(n10028) );
  AOI22_X1 U11088 ( .A1(n10002), .A2(keyinput80), .B1(n5081), .B2(keyinput124), 
        .ZN(n10001) );
  OAI221_X1 U11089 ( .B1(n10002), .B2(keyinput80), .C1(n5081), .C2(keyinput124), .A(n10001), .ZN(n10012) );
  AOI22_X1 U11090 ( .A1(n10004), .A2(keyinput87), .B1(keyinput118), .B2(n5877), 
        .ZN(n10003) );
  OAI221_X1 U11091 ( .B1(n10004), .B2(keyinput87), .C1(n5877), .C2(keyinput118), .A(n10003), .ZN(n10011) );
  INV_X1 U11092 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n10006) );
  AOI22_X1 U11093 ( .A1(n5606), .A2(keyinput22), .B1(keyinput76), .B2(n10006), 
        .ZN(n10005) );
  OAI221_X1 U11094 ( .B1(n5606), .B2(keyinput22), .C1(n10006), .C2(keyinput76), 
        .A(n10005), .ZN(n10010) );
  AOI22_X1 U11095 ( .A1(n10008), .A2(keyinput70), .B1(keyinput88), .B2(n6023), 
        .ZN(n10007) );
  OAI221_X1 U11096 ( .B1(n10008), .B2(keyinput70), .C1(n6023), .C2(keyinput88), 
        .A(n10007), .ZN(n10009) );
  NOR4_X1 U11097 ( .A1(n10012), .A2(n10011), .A3(n10010), .A4(n10009), .ZN(
        n10027) );
  AOI22_X1 U11098 ( .A1(n10014), .A2(keyinput63), .B1(keyinput30), .B2(n6167), 
        .ZN(n10013) );
  OAI221_X1 U11099 ( .B1(n10014), .B2(keyinput63), .C1(n6167), .C2(keyinput30), 
        .A(n10013), .ZN(n10025) );
  INV_X1 U11100 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10237) );
  AOI22_X1 U11101 ( .A1(n10016), .A2(keyinput105), .B1(keyinput65), .B2(n10237), .ZN(n10015) );
  OAI221_X1 U11102 ( .B1(n10016), .B2(keyinput105), .C1(n10237), .C2(
        keyinput65), .A(n10015), .ZN(n10024) );
  AOI22_X1 U11103 ( .A1(n10018), .A2(keyinput7), .B1(keyinput114), .B2(n7096), 
        .ZN(n10017) );
  OAI221_X1 U11104 ( .B1(n10018), .B2(keyinput7), .C1(n7096), .C2(keyinput114), 
        .A(n10017), .ZN(n10023) );
  INV_X1 U11105 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10021) );
  INV_X1 U11106 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n10020) );
  AOI22_X1 U11107 ( .A1(n10021), .A2(keyinput45), .B1(n10020), .B2(keyinput79), 
        .ZN(n10019) );
  OAI221_X1 U11108 ( .B1(n10021), .B2(keyinput45), .C1(n10020), .C2(keyinput79), .A(n10019), .ZN(n10022) );
  NOR4_X1 U11109 ( .A1(n10025), .A2(n10024), .A3(n10023), .A4(n10022), .ZN(
        n10026) );
  NAND4_X1 U11110 ( .A1(n10029), .A2(n10028), .A3(n10027), .A4(n10026), .ZN(
        n10205) );
  AOI22_X1 U11111 ( .A1(n10270), .A2(keyinput90), .B1(n10031), .B2(keyinput69), 
        .ZN(n10030) );
  OAI221_X1 U11112 ( .B1(n10270), .B2(keyinput90), .C1(n10031), .C2(keyinput69), .A(n10030), .ZN(n10043) );
  AOI22_X1 U11113 ( .A1(n10034), .A2(keyinput3), .B1(keyinput41), .B2(n10033), 
        .ZN(n10032) );
  OAI221_X1 U11114 ( .B1(n10034), .B2(keyinput3), .C1(n10033), .C2(keyinput41), 
        .A(n10032), .ZN(n10042) );
  AOI22_X1 U11115 ( .A1(n10037), .A2(keyinput19), .B1(keyinput6), .B2(n10036), 
        .ZN(n10035) );
  OAI221_X1 U11116 ( .B1(n10037), .B2(keyinput19), .C1(n10036), .C2(keyinput6), 
        .A(n10035), .ZN(n10041) );
  XNOR2_X1 U11117 ( .A(P2_REG1_REG_30__SCAN_IN), .B(keyinput116), .ZN(n10039)
         );
  XNOR2_X1 U11118 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput52), .ZN(n10038) );
  NAND2_X1 U11119 ( .A1(n10039), .A2(n10038), .ZN(n10040) );
  NOR4_X1 U11120 ( .A1(n10043), .A2(n10042), .A3(n10041), .A4(n10040), .ZN(
        n10086) );
  AOI22_X1 U11121 ( .A1(n5440), .A2(keyinput55), .B1(keyinput85), .B2(n10045), 
        .ZN(n10044) );
  OAI221_X1 U11122 ( .B1(n5440), .B2(keyinput55), .C1(n10045), .C2(keyinput85), 
        .A(n10044), .ZN(n10057) );
  AOI22_X1 U11123 ( .A1(n10048), .A2(keyinput74), .B1(keyinput17), .B2(n10047), 
        .ZN(n10046) );
  OAI221_X1 U11124 ( .B1(n10048), .B2(keyinput74), .C1(n10047), .C2(keyinput17), .A(n10046), .ZN(n10056) );
  AOI22_X1 U11125 ( .A1(n10051), .A2(keyinput99), .B1(n10050), .B2(keyinput37), 
        .ZN(n10049) );
  OAI221_X1 U11126 ( .B1(n10051), .B2(keyinput99), .C1(n10050), .C2(keyinput37), .A(n10049), .ZN(n10055) );
  XOR2_X1 U11127 ( .A(n4975), .B(keyinput101), .Z(n10053) );
  XNOR2_X1 U11128 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput115), .ZN(n10052) );
  NAND2_X1 U11129 ( .A1(n10053), .A2(n10052), .ZN(n10054) );
  NOR4_X1 U11130 ( .A1(n10057), .A2(n10056), .A3(n10055), .A4(n10054), .ZN(
        n10085) );
  INV_X1 U11131 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10059) );
  AOI22_X1 U11132 ( .A1(n6724), .A2(keyinput35), .B1(n10059), .B2(keyinput36), 
        .ZN(n10058) );
  OAI221_X1 U11133 ( .B1(n6724), .B2(keyinput35), .C1(n10059), .C2(keyinput36), 
        .A(n10058), .ZN(n10071) );
  AOI22_X1 U11134 ( .A1(n10062), .A2(keyinput106), .B1(n10061), .B2(keyinput24), .ZN(n10060) );
  OAI221_X1 U11135 ( .B1(n10062), .B2(keyinput106), .C1(n10061), .C2(
        keyinput24), .A(n10060), .ZN(n10070) );
  AOI22_X1 U11136 ( .A1(n10065), .A2(keyinput39), .B1(n10064), .B2(keyinput107), .ZN(n10063) );
  OAI221_X1 U11137 ( .B1(n10065), .B2(keyinput39), .C1(n10064), .C2(
        keyinput107), .A(n10063), .ZN(n10069) );
  XNOR2_X1 U11138 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput62), .ZN(n10067) );
  XNOR2_X1 U11139 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput25), .ZN(n10066)
         );
  NAND2_X1 U11140 ( .A1(n10067), .A2(n10066), .ZN(n10068) );
  NOR4_X1 U11141 ( .A1(n10071), .A2(n10070), .A3(n10069), .A4(n10068), .ZN(
        n10084) );
  AOI22_X1 U11142 ( .A1(n9659), .A2(keyinput77), .B1(keyinput83), .B2(P2_U3152), .ZN(n10072) );
  OAI221_X1 U11143 ( .B1(n9659), .B2(keyinput77), .C1(P2_U3152), .C2(
        keyinput83), .A(n10072), .ZN(n10082) );
  AOI22_X1 U11144 ( .A1(n10074), .A2(keyinput111), .B1(keyinput98), .B2(n6535), 
        .ZN(n10073) );
  OAI221_X1 U11145 ( .B1(n10074), .B2(keyinput111), .C1(n6535), .C2(keyinput98), .A(n10073), .ZN(n10081) );
  AOI22_X1 U11146 ( .A1(n6518), .A2(keyinput40), .B1(keyinput51), .B2(n10076), 
        .ZN(n10075) );
  OAI221_X1 U11147 ( .B1(n6518), .B2(keyinput40), .C1(n10076), .C2(keyinput51), 
        .A(n10075), .ZN(n10080) );
  AOI22_X1 U11148 ( .A1(n5551), .A2(keyinput86), .B1(keyinput97), .B2(n10078), 
        .ZN(n10077) );
  OAI221_X1 U11149 ( .B1(n5551), .B2(keyinput86), .C1(n10078), .C2(keyinput97), 
        .A(n10077), .ZN(n10079) );
  NOR4_X1 U11150 ( .A1(n10082), .A2(n10081), .A3(n10080), .A4(n10079), .ZN(
        n10083) );
  NAND4_X1 U11151 ( .A1(n10086), .A2(n10085), .A3(n10084), .A4(n10083), .ZN(
        n10204) );
  AOI22_X1 U11152 ( .A1(n7456), .A2(keyinput120), .B1(n10088), .B2(keyinput31), 
        .ZN(n10087) );
  OAI221_X1 U11153 ( .B1(n7456), .B2(keyinput120), .C1(n10088), .C2(keyinput31), .A(n10087), .ZN(n10099) );
  AOI22_X1 U11154 ( .A1(n7499), .A2(keyinput117), .B1(n5163), .B2(keyinput100), 
        .ZN(n10089) );
  OAI221_X1 U11155 ( .B1(n7499), .B2(keyinput117), .C1(n5163), .C2(keyinput100), .A(n10089), .ZN(n10098) );
  AOI22_X1 U11156 ( .A1(n10092), .A2(keyinput73), .B1(keyinput43), .B2(n10091), 
        .ZN(n10090) );
  OAI221_X1 U11157 ( .B1(n10092), .B2(keyinput73), .C1(n10091), .C2(keyinput43), .A(n10090), .ZN(n10097) );
  AOI22_X1 U11158 ( .A1(n10095), .A2(keyinput28), .B1(n10094), .B2(keyinput14), 
        .ZN(n10093) );
  OAI221_X1 U11159 ( .B1(n10095), .B2(keyinput28), .C1(n10094), .C2(keyinput14), .A(n10093), .ZN(n10096) );
  NOR4_X1 U11160 ( .A1(n10099), .A2(n10098), .A3(n10097), .A4(n10096), .ZN(
        n10140) );
  AOI22_X1 U11161 ( .A1(n10101), .A2(keyinput121), .B1(keyinput42), .B2(n8927), 
        .ZN(n10100) );
  OAI221_X1 U11162 ( .B1(n10101), .B2(keyinput121), .C1(n8927), .C2(keyinput42), .A(n10100), .ZN(n10110) );
  AOI22_X1 U11163 ( .A1(n9247), .A2(keyinput89), .B1(n10103), .B2(keyinput93), 
        .ZN(n10102) );
  OAI221_X1 U11164 ( .B1(n9247), .B2(keyinput89), .C1(n10103), .C2(keyinput93), 
        .A(n10102), .ZN(n10109) );
  AOI22_X1 U11165 ( .A1(n6605), .A2(keyinput50), .B1(n6079), .B2(keyinput23), 
        .ZN(n10104) );
  OAI221_X1 U11166 ( .B1(n6605), .B2(keyinput50), .C1(n6079), .C2(keyinput23), 
        .A(n10104), .ZN(n10108) );
  XNOR2_X1 U11167 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput127), .ZN(n10106)
         );
  XNOR2_X1 U11168 ( .A(SI_0_), .B(keyinput0), .ZN(n10105) );
  NAND2_X1 U11169 ( .A1(n10106), .A2(n10105), .ZN(n10107) );
  NOR4_X1 U11170 ( .A1(n10110), .A2(n10109), .A3(n10108), .A4(n10107), .ZN(
        n10139) );
  INV_X1 U11171 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10112) );
  AOI22_X1 U11172 ( .A1(n10112), .A2(keyinput57), .B1(keyinput59), .B2(n7572), 
        .ZN(n10111) );
  OAI221_X1 U11173 ( .B1(n10112), .B2(keyinput57), .C1(n7572), .C2(keyinput59), 
        .A(n10111), .ZN(n10122) );
  AOI22_X1 U11174 ( .A1(n6156), .A2(keyinput34), .B1(n5094), .B2(keyinput18), 
        .ZN(n10113) );
  OAI221_X1 U11175 ( .B1(n6156), .B2(keyinput34), .C1(n5094), .C2(keyinput18), 
        .A(n10113), .ZN(n10121) );
  AOI22_X1 U11176 ( .A1(n10116), .A2(keyinput11), .B1(keyinput29), .B2(n10115), 
        .ZN(n10114) );
  OAI221_X1 U11177 ( .B1(n10116), .B2(keyinput11), .C1(n10115), .C2(keyinput29), .A(n10114), .ZN(n10120) );
  AOI22_X1 U11178 ( .A1(n9134), .A2(keyinput126), .B1(keyinput102), .B2(n10118), .ZN(n10117) );
  OAI221_X1 U11179 ( .B1(n9134), .B2(keyinput126), .C1(n10118), .C2(
        keyinput102), .A(n10117), .ZN(n10119) );
  NOR4_X1 U11180 ( .A1(n10122), .A2(n10121), .A3(n10120), .A4(n10119), .ZN(
        n10138) );
  INV_X1 U11181 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10124) );
  AOI22_X1 U11182 ( .A1(n10125), .A2(keyinput71), .B1(keyinput108), .B2(n10124), .ZN(n10123) );
  OAI221_X1 U11183 ( .B1(n10125), .B2(keyinput71), .C1(n10124), .C2(
        keyinput108), .A(n10123), .ZN(n10136) );
  AOI22_X1 U11184 ( .A1(n10128), .A2(keyinput64), .B1(n10127), .B2(keyinput26), 
        .ZN(n10126) );
  OAI221_X1 U11185 ( .B1(n10128), .B2(keyinput64), .C1(n10127), .C2(keyinput26), .A(n10126), .ZN(n10135) );
  AOI22_X1 U11186 ( .A1(n10221), .A2(keyinput5), .B1(n10130), .B2(keyinput110), 
        .ZN(n10129) );
  OAI221_X1 U11187 ( .B1(n10221), .B2(keyinput5), .C1(n10130), .C2(keyinput110), .A(n10129), .ZN(n10134) );
  AOI22_X1 U11188 ( .A1(n10132), .A2(keyinput125), .B1(keyinput2), .B2(n10211), 
        .ZN(n10131) );
  OAI221_X1 U11189 ( .B1(n10132), .B2(keyinput125), .C1(n10211), .C2(keyinput2), .A(n10131), .ZN(n10133) );
  NOR4_X1 U11190 ( .A1(n10136), .A2(n10135), .A3(n10134), .A4(n10133), .ZN(
        n10137) );
  NAND4_X1 U11191 ( .A1(n10140), .A2(n10139), .A3(n10138), .A4(n10137), .ZN(
        n10203) );
  INV_X1 U11192 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10143) );
  AOI22_X1 U11193 ( .A1(n10143), .A2(keyinput75), .B1(keyinput49), .B2(n10142), 
        .ZN(n10141) );
  OAI221_X1 U11194 ( .B1(n10143), .B2(keyinput75), .C1(n10142), .C2(keyinput49), .A(n10141), .ZN(n10148) );
  AOI22_X1 U11195 ( .A1(n10146), .A2(keyinput94), .B1(n10145), .B2(keyinput58), 
        .ZN(n10144) );
  OAI221_X1 U11196 ( .B1(n10146), .B2(keyinput94), .C1(n10145), .C2(keyinput58), .A(n10144), .ZN(n10147) );
  NOR2_X1 U11197 ( .A1(n10148), .A2(n10147), .ZN(n10158) );
  INV_X1 U11198 ( .A(keyinput72), .ZN(n10149) );
  XNOR2_X1 U11199 ( .A(n10150), .B(n10149), .ZN(n10157) );
  XNOR2_X1 U11200 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput92), .ZN(n10156) );
  INV_X1 U11201 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10152) );
  AOI22_X1 U11202 ( .A1(n10153), .A2(keyinput47), .B1(n10152), .B2(keyinput32), 
        .ZN(n10151) );
  OAI221_X1 U11203 ( .B1(n10153), .B2(keyinput47), .C1(n10152), .C2(keyinput32), .A(n10151), .ZN(n10154) );
  INV_X1 U11204 ( .A(n10154), .ZN(n10155) );
  AND4_X1 U11205 ( .A1(n10158), .A2(n10157), .A3(n10156), .A4(n10155), .ZN(
        n10201) );
  AOI22_X1 U11206 ( .A1(n10160), .A2(keyinput66), .B1(keyinput33), .B2(n6725), 
        .ZN(n10159) );
  OAI221_X1 U11207 ( .B1(n10160), .B2(keyinput66), .C1(n6725), .C2(keyinput33), 
        .A(n10159), .ZN(n10170) );
  AOI22_X1 U11208 ( .A1(n5935), .A2(keyinput10), .B1(n10162), .B2(keyinput1), 
        .ZN(n10161) );
  OAI221_X1 U11209 ( .B1(n5935), .B2(keyinput10), .C1(n10162), .C2(keyinput1), 
        .A(n10161), .ZN(n10169) );
  INV_X1 U11210 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10238) );
  XOR2_X1 U11211 ( .A(n10238), .B(keyinput119), .Z(n10167) );
  INV_X1 U11212 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10163) );
  XOR2_X1 U11213 ( .A(n10163), .B(keyinput44), .Z(n10166) );
  XNOR2_X1 U11214 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput84), .ZN(n10165)
         );
  XNOR2_X1 U11215 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput12), .ZN(n10164) );
  NAND4_X1 U11216 ( .A1(n10167), .A2(n10166), .A3(n10165), .A4(n10164), .ZN(
        n10168) );
  NOR3_X1 U11217 ( .A1(n10170), .A2(n10169), .A3(n10168), .ZN(n10200) );
  AOI22_X1 U11218 ( .A1(n10172), .A2(keyinput27), .B1(keyinput56), .B2(n7541), 
        .ZN(n10171) );
  OAI221_X1 U11219 ( .B1(n10172), .B2(keyinput27), .C1(n7541), .C2(keyinput56), 
        .A(n10171), .ZN(n10182) );
  INV_X1 U11220 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U11221 ( .A1(n5873), .A2(keyinput122), .B1(keyinput81), .B2(n10174), 
        .ZN(n10173) );
  OAI221_X1 U11222 ( .B1(n5873), .B2(keyinput122), .C1(n10174), .C2(keyinput81), .A(n10173), .ZN(n10181) );
  XNOR2_X1 U11223 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput13), .ZN(n10177) );
  XNOR2_X1 U11224 ( .A(P1_REG2_REG_20__SCAN_IN), .B(keyinput78), .ZN(n10176)
         );
  XNOR2_X1 U11225 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput15), .ZN(n10175) );
  NAND3_X1 U11226 ( .A1(n10177), .A2(n10176), .A3(n10175), .ZN(n10180) );
  XNOR2_X1 U11227 ( .A(n10178), .B(keyinput104), .ZN(n10179) );
  NOR4_X1 U11228 ( .A1(n10182), .A2(n10181), .A3(n10180), .A4(n10179), .ZN(
        n10199) );
  AOI22_X1 U11229 ( .A1(n10185), .A2(keyinput82), .B1(n10184), .B2(keyinput8), 
        .ZN(n10183) );
  OAI221_X1 U11230 ( .B1(n10185), .B2(keyinput82), .C1(n10184), .C2(keyinput8), 
        .A(n10183), .ZN(n10197) );
  AOI22_X1 U11231 ( .A1(n10188), .A2(keyinput21), .B1(keyinput96), .B2(n10187), 
        .ZN(n10186) );
  OAI221_X1 U11232 ( .B1(n10188), .B2(keyinput21), .C1(n10187), .C2(keyinput96), .A(n10186), .ZN(n10196) );
  AOI22_X1 U11233 ( .A1(n10191), .A2(keyinput109), .B1(n10190), .B2(keyinput16), .ZN(n10189) );
  OAI221_X1 U11234 ( .B1(n10191), .B2(keyinput109), .C1(n10190), .C2(
        keyinput16), .A(n10189), .ZN(n10195) );
  XOR2_X1 U11235 ( .A(n6765), .B(keyinput54), .Z(n10193) );
  XNOR2_X1 U11236 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput20), .ZN(n10192) );
  NAND2_X1 U11237 ( .A1(n10193), .A2(n10192), .ZN(n10194) );
  NOR4_X1 U11238 ( .A1(n10197), .A2(n10196), .A3(n10195), .A4(n10194), .ZN(
        n10198) );
  NAND4_X1 U11239 ( .A1(n10201), .A2(n10200), .A3(n10199), .A4(n10198), .ZN(
        n10202) );
  NOR4_X1 U11240 ( .A1(n10205), .A2(n10204), .A3(n10203), .A4(n10202), .ZN(
        n10262) );
  NAND4_X1 U11241 ( .A1(SI_5_), .A2(P2_IR_REG_8__SCAN_IN), .A3(
        P2_REG3_REG_11__SCAN_IN), .A4(P2_REG0_REG_9__SCAN_IN), .ZN(n10209) );
  NAND4_X1 U11242 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_REG0_REG_21__SCAN_IN), .ZN(n10208) );
  NAND4_X1 U11243 ( .A1(P1_REG1_REG_22__SCAN_IN), .A2(P2_REG1_REG_13__SCAN_IN), 
        .A3(P2_REG1_REG_2__SCAN_IN), .A4(P2_REG1_REG_1__SCAN_IN), .ZN(n10207)
         );
  NAND4_X1 U11244 ( .A1(SI_19_), .A2(P2_IR_REG_16__SCAN_IN), .A3(
        P2_REG1_REG_12__SCAN_IN), .A4(P2_REG2_REG_9__SCAN_IN), .ZN(n10206) );
  NOR4_X1 U11245 ( .A1(n10209), .A2(n10208), .A3(n10207), .A4(n10206), .ZN(
        n10229) );
  NAND4_X1 U11246 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(SI_20_), .A3(SI_12_), .A4(
        P2_D_REG_0__SCAN_IN), .ZN(n10216) );
  NAND4_X1 U11247 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_U3084), .A3(n10211), 
        .A4(n10210), .ZN(n10215) );
  NAND4_X1 U11248 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), 
        .A3(P2_REG0_REG_23__SCAN_IN), .A4(P2_REG1_REG_31__SCAN_IN), .ZN(n10214) );
  NAND4_X1 U11249 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(SI_16_), .A3(
        P1_DATAO_REG_13__SCAN_IN), .A4(P2_REG3_REG_13__SCAN_IN), .ZN(n10213)
         );
  NOR4_X1 U11250 ( .A1(n10216), .A2(n10215), .A3(n10214), .A4(n10213), .ZN(
        n10228) );
  NAND4_X1 U11251 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), .A3(P1_REG2_REG_27__SCAN_IN), .A4(P1_REG2_REG_20__SCAN_IN), .ZN(n10220) );
  NAND4_X1 U11252 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(P1_REG2_REG_10__SCAN_IN), 
        .A3(P2_REG2_REG_29__SCAN_IN), .A4(P2_REG2_REG_30__SCAN_IN), .ZN(n10219) );
  NAND4_X1 U11253 ( .A1(n10217), .A2(P2_REG3_REG_17__SCAN_IN), .A3(
        P2_REG2_REG_21__SCAN_IN), .A4(P2_REG2_REG_18__SCAN_IN), .ZN(n10218) );
  NOR4_X1 U11254 ( .A1(n10221), .A2(n10220), .A3(n10219), .A4(n10218), .ZN(
        n10227) );
  NAND4_X1 U11255 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n10225) );
  NAND4_X1 U11256 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_REG0_REG_28__SCAN_IN), 
        .A3(P1_REG0_REG_22__SCAN_IN), .A4(P1_REG0_REG_29__SCAN_IN), .ZN(n10224) );
  NAND4_X1 U11257 ( .A1(P1_REG2_REG_23__SCAN_IN), .A2(P1_REG0_REG_16__SCAN_IN), 
        .A3(P1_REG1_REG_3__SCAN_IN), .A4(P1_DATAO_REG_30__SCAN_IN), .ZN(n10223) );
  NAND4_X1 U11258 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_REG3_REG_5__SCAN_IN), .A4(P1_REG0_REG_6__SCAN_IN), .ZN(n10222) );
  NOR4_X1 U11259 ( .A1(n10225), .A2(n10224), .A3(n10223), .A4(n10222), .ZN(
        n10226) );
  AND4_X1 U11260 ( .A1(n10229), .A2(n10228), .A3(n10227), .A4(n10226), .ZN(
        n10253) );
  NOR4_X1 U11261 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(P2_DATAO_REG_2__SCAN_IN), 
        .A3(SI_0_), .A4(P2_DATAO_REG_1__SCAN_IN), .ZN(n10230) );
  NAND3_X1 U11262 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n10230), .A3(n10270), 
        .ZN(n10236) );
  NOR4_X1 U11263 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .A3(
        P2_REG3_REG_10__SCAN_IN), .A4(P2_REG3_REG_5__SCAN_IN), .ZN(n10234) );
  NOR4_X1 U11264 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(P2_DATAO_REG_8__SCAN_IN), 
        .A3(P2_IR_REG_21__SCAN_IN), .A4(n10257), .ZN(n10233) );
  NOR4_X1 U11265 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(P2_REG0_REG_26__SCAN_IN), 
        .A3(P2_REG0_REG_20__SCAN_IN), .A4(P2_REG1_REG_30__SCAN_IN), .ZN(n10232) );
  NOR4_X1 U11266 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_D_REG_1__SCAN_IN), .A3(
        P2_IR_REG_17__SCAN_IN), .A4(P2_REG3_REG_8__SCAN_IN), .ZN(n10231) );
  NAND4_X1 U11267 ( .A1(n10234), .A2(n10233), .A3(n10232), .A4(n10231), .ZN(
        n10235) );
  NOR4_X1 U11268 ( .A1(P1_RD_REG_SCAN_IN), .A2(P2_U3152), .A3(n10236), .A4(
        n10235), .ZN(n10252) );
  NOR4_X1 U11269 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(n10238), .A4(n10237), .ZN(n10251) );
  NOR4_X1 U11270 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P2_DATAO_REG_11__SCAN_IN), 
        .A3(P1_REG0_REG_11__SCAN_IN), .A4(P1_REG1_REG_0__SCAN_IN), .ZN(n10242)
         );
  NOR4_X1 U11271 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_REG2_REG_8__SCAN_IN), 
        .A3(P1_REG2_REG_5__SCAN_IN), .A4(P1_REG2_REG_4__SCAN_IN), .ZN(n10241)
         );
  NOR4_X1 U11272 ( .A1(P2_REG2_REG_27__SCAN_IN), .A2(P2_REG2_REG_14__SCAN_IN), 
        .A3(P2_REG2_REG_13__SCAN_IN), .A4(P2_REG2_REG_22__SCAN_IN), .ZN(n10240) );
  NOR4_X1 U11273 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG0_REG_21__SCAN_IN), 
        .A3(P1_REG2_REG_18__SCAN_IN), .A4(P2_B_REG_SCAN_IN), .ZN(n10239) );
  AND4_X1 U11274 ( .A1(n10242), .A2(n10241), .A3(n10240), .A4(n10239), .ZN(
        n10249) );
  NOR4_X1 U11275 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(P2_REG2_REG_8__SCAN_IN), 
        .A3(P2_REG2_REG_6__SCAN_IN), .A4(P2_REG1_REG_3__SCAN_IN), .ZN(n10246)
         );
  NOR4_X1 U11276 ( .A1(SI_9_), .A2(P2_DATAO_REG_9__SCAN_IN), .A3(
        P2_IR_REG_12__SCAN_IN), .A4(P2_REG0_REG_8__SCAN_IN), .ZN(n10245) );
  NOR4_X1 U11277 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_REG1_REG_10__SCAN_IN), 
        .A3(P1_REG0_REG_8__SCAN_IN), .A4(P1_REG0_REG_3__SCAN_IN), .ZN(n10244)
         );
  NOR4_X1 U11278 ( .A1(P1_REG0_REG_27__SCAN_IN), .A2(P1_REG1_REG_26__SCAN_IN), 
        .A3(P1_REG2_REG_24__SCAN_IN), .A4(P1_REG0_REG_24__SCAN_IN), .ZN(n10243) );
  AND4_X1 U11279 ( .A1(n10246), .A2(n10245), .A3(n10244), .A4(n10243), .ZN(
        n10248) );
  AND4_X1 U11280 ( .A1(n10249), .A2(n10248), .A3(P2_REG3_REG_26__SCAN_IN), 
        .A4(n10247), .ZN(n10250) );
  NAND4_X1 U11281 ( .A1(n10253), .A2(n10252), .A3(n10251), .A4(n10250), .ZN(
        n10260) );
  OAI222_X1 U11282 ( .A1(n10258), .A2(n10257), .B1(n10256), .B2(n10255), .C1(
        P2_U3152), .C2(n10254), .ZN(n10259) );
  XOR2_X1 U11283 ( .A(n10260), .B(n10259), .Z(n10261) );
  XNOR2_X1 U11284 ( .A(n10262), .B(n10261), .ZN(P2_U3354) );
  XOR2_X1 U11285 ( .A(n10263), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11286 ( .A(n10264), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11287 ( .A1(n10266), .A2(n10265), .ZN(n10267) );
  XOR2_X1 U11288 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10267), .Z(ADD_1071_U51) );
  OAI21_X1 U11289 ( .B1(n10270), .B2(n10269), .A(n10268), .ZN(n10271) );
  XNOR2_X1 U11290 ( .A(n10271), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11291 ( .B1(n10274), .B2(n10273), .A(n10272), .ZN(ADD_1071_U47) );
  XOR2_X1 U11292 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10275), .Z(ADD_1071_U48) );
  XOR2_X1 U11293 ( .A(n10277), .B(n10276), .Z(ADD_1071_U54) );
  XOR2_X1 U11294 ( .A(n10279), .B(n10278), .Z(ADD_1071_U53) );
  XNOR2_X1 U11295 ( .A(n10281), .B(n10280), .ZN(ADD_1071_U52) );
  INV_X1 U4890 ( .A(n6177), .ZN(n6155) );
  CLKBUF_X1 U4898 ( .A(n7964), .Z(n4381) );
  CLKBUF_X1 U5047 ( .A(n5773), .Z(n6713) );
  CLKBUF_X1 U5061 ( .A(n5767), .Z(n6606) );
endmodule

