

module b20_C_AntiSAT_k_256_5 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, ADD_1068_U4, ADD_1068_U55, 
        ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, 
        ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, 
        ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, 
        ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, 
        P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, 
        P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, 
        P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, 
        P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, 
        P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, 
        P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, 
        P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, 
        P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, 
        P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, 
        P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, 
        P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, 
        P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492;

  NAND2_X1 U5013 ( .A1(n7921), .A2(n6712), .ZN(n6713) );
  CLKBUF_X2 U5014 ( .A(n6309), .Z(n6483) );
  NAND2_X1 U5015 ( .A1(n5294), .A2(n5295), .ZN(n5741) );
  INV_X1 U5016 ( .A(n5743), .ZN(n5618) );
  CLKBUF_X1 U5017 ( .A(n8790), .Z(n4507) );
  NOR2_X1 U5018 ( .A1(n7368), .A2(n8676), .ZN(n8790) );
  INV_X1 U5019 ( .A(n9696), .ZN(n4508) );
  INV_X2 U5020 ( .A(n4508), .ZN(n4509) );
  NAND2_X1 U5021 ( .A1(n4813), .A2(n5960), .ZN(n6066) );
  INV_X1 U5022 ( .A(n8798), .ZN(n8262) );
  CLKBUF_X3 U5023 ( .A(n5993), .Z(n8971) );
  AND2_X1 U5024 ( .A1(n5960), .A2(n7467), .ZN(n6043) );
  AND2_X1 U5025 ( .A1(n5064), .A2(n5266), .ZN(n5063) );
  INV_X1 U5026 ( .A(n8435), .ZN(n8439) );
  INV_X1 U5027 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8955) );
  NAND2_X2 U5028 ( .A1(n5949), .A2(n4511), .ZN(n6845) );
  OAI21_X1 U5029 ( .B1(n6814), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n4677), .ZN(
        n5135) );
  OAI211_X1 U5030 ( .C1(n7014), .C2(n6266), .A(n6268), .B(n6267), .ZN(n6573)
         );
  OR2_X1 U5031 ( .A1(n4594), .A2(n5421), .ZN(n5291) );
  INV_X1 U5032 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7406) );
  AOI222_X1 U5033 ( .A1(n9789), .A2(n9788), .B1(n9787), .B2(n9786), .C1(
        P1_REG2_REG_4__SCAN_IN), .C2(n9785), .ZN(n9799) );
  INV_X2 U5034 ( .A(n9516), .ZN(n9785) );
  NAND3_X2 U5035 ( .A1(n9692), .A2(n7513), .A3(n4877), .ZN(n7512) );
  NAND2_X2 U5036 ( .A1(n4876), .A2(n6013), .ZN(n9692) );
  NAND2_X1 U5037 ( .A1(n6266), .A2(n6265), .ZN(n4510) );
  NAND2_X1 U5038 ( .A1(n6266), .A2(n6265), .ZN(n6274) );
  INV_X1 U5039 ( .A(n6274), .ZN(n8249) );
  OR2_X2 U5040 ( .A1(n7923), .A2(n7924), .ZN(n7921) );
  OAI222_X1 U5041 ( .A1(n8965), .A2(n8001), .B1(P2_U3151), .B2(n7993), .C1(
        n7992), .C2(n8102), .ZN(P2_U3270) );
  AND3_X4 U5042 ( .A1(n5425), .A2(n5424), .A3(n5423), .ZN(n5883) );
  NAND2_X2 U5043 ( .A1(n6285), .A2(n6284), .ZN(n8799) );
  XNOR2_X2 U5044 ( .A(n5630), .B(n5629), .ZN(n9214) );
  XNOR2_X2 U5045 ( .A(n5139), .B(SI_2_), .ZN(n5623) );
  OAI222_X1 U5046 ( .A1(n9633), .A2(n8095), .B1(P1_U3086), .B2(n5949), .C1(
        n8961), .C2(n9629), .ZN(P1_U3327) );
  AND2_X1 U5047 ( .A1(n5949), .A2(n6843), .ZN(n9696) );
  NAND2_X1 U5048 ( .A1(n5292), .A2(n5294), .ZN(n5617) );
  NAND2_X1 U5049 ( .A1(n6066), .A2(n5983), .ZN(n5993) );
  NAND4_X2 U5050 ( .A1(n6260), .A2(n6259), .A3(n6258), .A4(n6257), .ZN(n6572)
         );
  NAND4_X2 U5051 ( .A1(n6273), .A2(n6272), .A3(n6271), .A4(n6270), .ZN(n8481)
         );
  NAND2_X1 U5052 ( .A1(n6545), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6273) );
  NAND2_X2 U5053 ( .A1(n6125), .A2(n6124), .ZN(n9036) );
  XNOR2_X2 U5054 ( .A(n6713), .B(n7740), .ZN(n7928) );
  OAI21_X2 U5055 ( .B1(n9636), .B2(n4873), .A(n4872), .ZN(n9138) );
  BUF_X2 U5056 ( .A(n5950), .Z(n4511) );
  XNOR2_X1 U5057 ( .A(n5272), .B(P1_IR_REG_27__SCAN_IN), .ZN(n5950) );
  INV_X1 U5058 ( .A(n8279), .ZN(n4512) );
  NAND2_X1 U5059 ( .A1(n7256), .A2(n7257), .ZN(n7255) );
  NAND2_X1 U5060 ( .A1(n6571), .A2(n8296), .ZN(n7173) );
  INV_X1 U5061 ( .A(n7539), .ZN(n9873) );
  INV_X2 U5062 ( .A(n6701), .ZN(n4513) );
  INV_X1 U5063 ( .A(n6572), .ZN(n6574) );
  BUF_X1 U5064 ( .A(n5634), .Z(n4516) );
  INV_X2 U5065 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5930) );
  OR2_X1 U5066 ( .A1(n6802), .A2(n10049), .ZN(n4936) );
  NAND2_X1 U5067 ( .A1(n9054), .A2(n9055), .ZN(n6182) );
  AOI21_X1 U5068 ( .B1(n9036), .B2(n9037), .A(n6132), .ZN(n9130) );
  NAND2_X1 U5069 ( .A1(n4957), .A2(n4956), .ZN(n8694) );
  AOI22_X1 U5070 ( .A1(n5873), .A2(n4783), .B1(n5871), .B2(n5872), .ZN(n4751)
         );
  XNOR2_X1 U5071 ( .A(n5728), .B(n5727), .ZN(n9626) );
  OAI22_X1 U5072 ( .A1(n5736), .A2(n5735), .B1(SI_30_), .B2(n5725), .ZN(n5728)
         );
  NAND2_X1 U5073 ( .A1(n8235), .A2(n8234), .ZN(n8233) );
  AOI21_X1 U5074 ( .B1(n4944), .B2(n4947), .A(n8653), .ZN(n4942) );
  OAI21_X1 U5075 ( .B1(n9450), .B2(n4796), .A(n4531), .ZN(n4801) );
  NAND2_X1 U5076 ( .A1(n8015), .A2(n8014), .ZN(n8013) );
  OAI21_X1 U5077 ( .B1(n4888), .B2(n7988), .A(n4885), .ZN(n8762) );
  NAND2_X1 U5078 ( .A1(n6065), .A2(n6068), .ZN(n9636) );
  NAND2_X1 U5079 ( .A1(n9460), .A2(n9459), .ZN(n9458) );
  AOI21_X1 U5080 ( .B1(n9005), .B2(n4862), .A(n9080), .ZN(n4861) );
  NAND3_X1 U5081 ( .A1(n9647), .A2(n9505), .A3(n9506), .ZN(n9504) );
  AND2_X1 U5082 ( .A1(n6131), .A2(n6130), .ZN(n6132) );
  OR2_X1 U5083 ( .A1(n9470), .A2(n8053), .ZN(n5115) );
  AND2_X1 U5084 ( .A1(n8052), .A2(n4600), .ZN(n5045) );
  NAND2_X1 U5085 ( .A1(n5352), .A2(n5351), .ZN(n9176) );
  NAND2_X1 U5086 ( .A1(n7661), .A2(n8323), .ZN(n7663) );
  AND2_X1 U5087 ( .A1(n7834), .A2(n4538), .ZN(n9660) );
  NAND2_X1 U5088 ( .A1(n4939), .A2(n4938), .ZN(n7601) );
  AND2_X1 U5089 ( .A1(n7756), .A2(n9892), .ZN(n7791) );
  AOI21_X1 U5090 ( .B1(n5107), .B2(n7502), .A(n4556), .ZN(n5105) );
  NAND2_X1 U5091 ( .A1(n5028), .A2(n5027), .ZN(n5511) );
  NAND2_X1 U5092 ( .A1(n5665), .A2(n5664), .ZN(n9883) );
  INV_X2 U5093 ( .A(n6701), .ZN(n6753) );
  OR2_X1 U5094 ( .A1(n7646), .A2(n7650), .ZN(n9792) );
  XNOR2_X1 U5095 ( .A(n4810), .B(n4809), .ZN(n6836) );
  AOI21_X1 U5096 ( .B1(n5690), .B2(n5156), .A(n4572), .ZN(n4810) );
  NAND4_X1 U5097 ( .A1(n6248), .A2(n6247), .A3(n6246), .A4(n6245), .ZN(n8482)
         );
  NAND2_X1 U5098 ( .A1(n5155), .A2(n5154), .ZN(n5690) );
  INV_X2 U5099 ( .A(n6256), .ZN(n6565) );
  NAND2_X1 U5100 ( .A1(n6277), .A2(n4542), .ZN(n9996) );
  OR2_X1 U5101 ( .A1(n6653), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6652) );
  NAND3_X1 U5102 ( .A1(n5614), .A2(n5613), .A3(n5129), .ZN(n5980) );
  AND3_X1 U5103 ( .A1(n6291), .A2(n6290), .A3(n6289), .ZN(n10003) );
  CLKBUF_X2 U5104 ( .A(n5634), .Z(n4517) );
  NAND2_X1 U5105 ( .A1(n5128), .A2(n4657), .ZN(n7113) );
  NAND4_X1 U5106 ( .A1(n5622), .A2(n5621), .A3(n5620), .A4(n5619), .ZN(n9197)
         );
  MUX2_X1 U5107 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9634), .S(n6845), .Z(n7673) );
  NAND2_X1 U5108 ( .A1(n8954), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6239) );
  AND2_X1 U5109 ( .A1(n5956), .A2(n7778), .ZN(n7472) );
  XNOR2_X1 U5110 ( .A(n6241), .B(n6236), .ZN(n8028) );
  INV_X1 U5111 ( .A(n5956), .ZN(n6931) );
  NAND2_X1 U5112 ( .A1(n6614), .A2(n6215), .ZN(n8437) );
  OR2_X1 U5113 ( .A1(n6250), .A2(n8955), .ZN(n6252) );
  NAND2_X1 U5114 ( .A1(n5796), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U5115 ( .A1(n4869), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U5116 ( .A1(n5945), .A2(n5944), .ZN(n8002) );
  XNOR2_X1 U5117 ( .A(n5795), .B(n5794), .ZN(n7778) );
  XNOR2_X1 U5118 ( .A(n5947), .B(n5266), .ZN(n7965) );
  OAI21_X1 U5119 ( .B1(n6216), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6214) );
  XNOR2_X1 U5120 ( .A(n5289), .B(n9622), .ZN(n5292) );
  OR2_X1 U5121 ( .A1(n5588), .A2(n5421), .ZN(n5795) );
  XNOR2_X1 U5122 ( .A(n5886), .B(n5885), .ZN(n7471) );
  AND2_X1 U5123 ( .A1(n6368), .A2(n6209), .ZN(n6378) );
  NAND2_X2 U5124 ( .A1(n4917), .A2(n4547), .ZN(n7099) );
  NOR2_X1 U5125 ( .A1(n5264), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n4765) );
  AND2_X1 U5126 ( .A1(n5259), .A2(n5258), .ZN(n5055) );
  AND2_X1 U5127 ( .A1(n5265), .A2(n5885), .ZN(n5064) );
  NOR2_X1 U5128 ( .A1(n6227), .A2(n6226), .ZN(n6229) );
  NOR2_X1 U5129 ( .A1(n6208), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5111) );
  AND2_X1 U5130 ( .A1(n4554), .A2(n6262), .ZN(n6314) );
  AND2_X1 U5131 ( .A1(n5056), .A2(n5054), .ZN(n4523) );
  AND2_X1 U5132 ( .A1(n4727), .A2(n5057), .ZN(n5056) );
  OR2_X1 U5133 ( .A1(n5581), .A2(n5421), .ZN(n5626) );
  AND3_X1 U5134 ( .A1(n5930), .A2(n5794), .A3(n5933), .ZN(n5265) );
  AND3_X1 U5135 ( .A1(n5494), .A2(n4624), .A3(n4623), .ZN(n5263) );
  INV_X1 U5136 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5494) );
  NOR2_X1 U5137 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5257) );
  INV_X1 U5138 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5794) );
  NOR2_X1 U5139 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4727) );
  AND2_X1 U5140 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5269) );
  INV_X1 U5141 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5933) );
  INV_X1 U5142 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6207) );
  INV_X1 U5143 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5131) );
  INV_X4 U5144 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5145 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6424) );
  INV_X1 U5146 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6224) );
  INV_X1 U5147 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6225) );
  NOR2_X1 U5148 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5262) );
  NOR2_X1 U5149 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5261) );
  NOR2_X1 U5150 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5260) );
  INV_X1 U5151 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6203) );
  INV_X1 U5152 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5885) );
  OR2_X2 U5153 ( .A1(n5633), .A2(n6823), .ZN(n5587) );
  INV_X4 U5154 ( .A(n6528), .ZN(n8254) );
  BUF_X4 U5155 ( .A(n5983), .Z(n4514) );
  OAI21_X2 U5156 ( .B1(n7377), .B2(n5078), .A(n5076), .ZN(n7501) );
  OAI211_X2 U5157 ( .C1(n5789), .C2(n5788), .A(n5787), .B(n5875), .ZN(n5887)
         );
  OR2_X2 U5158 ( .A1(n5782), .A2(n5781), .ZN(n5788) );
  XNOR2_X2 U5159 ( .A(n5271), .B(n5270), .ZN(n5949) );
  INV_X2 U5160 ( .A(n6295), .ZN(n4515) );
  AND2_X1 U5161 ( .A1(n8101), .A2(n6244), .ZN(n6280) );
  XNOR2_X2 U5162 ( .A(n6252), .B(n6251), .ZN(n6625) );
  NAND2_X1 U5163 ( .A1(n6845), .A2(n6814), .ZN(n5634) );
  AOI21_X2 U5164 ( .B1(n8201), .B2(n8202), .A(n4543), .ZN(n8172) );
  NAND2_X2 U5165 ( .A1(n6743), .A2(n6742), .ZN(n8201) );
  NAND2_X1 U5166 ( .A1(n6066), .A2(n5983), .ZN(n4518) );
  INV_X2 U5167 ( .A(n8481), .ZN(n4878) );
  XNOR2_X2 U5168 ( .A(n6683), .B(n6573), .ZN(n6685) );
  OAI21_X4 U5169 ( .B1(n6682), .B2(n7362), .A(n6681), .ZN(n6683) );
  AOI21_X2 U5170 ( .B1(n9013), .B2(n9014), .A(n5113), .ZN(n9109) );
  INV_X1 U5171 ( .A(n9789), .ZN(n4839) );
  OAI211_X2 U5172 ( .C1(n6889), .C2(n6845), .A(n5587), .B(n5586), .ZN(n9789)
         );
  NAND2_X1 U5173 ( .A1(n4726), .A2(n8435), .ZN(n4725) );
  NAND2_X1 U5174 ( .A1(n8301), .A2(n8439), .ZN(n4724) );
  INV_X1 U5175 ( .A(n8293), .ZN(n4726) );
  NAND2_X1 U5176 ( .A1(n6750), .A2(n8224), .ZN(n5103) );
  AND2_X1 U5177 ( .A1(n5111), .A2(n6230), .ZN(n5110) );
  NAND2_X1 U5178 ( .A1(n6562), .A2(n6561), .ZN(n8251) );
  NAND2_X1 U5179 ( .A1(n4966), .A2(n4569), .ZN(n8003) );
  AOI21_X1 U5180 ( .B1(n4946), .B2(n4945), .A(n4576), .ZN(n4944) );
  INV_X1 U5181 ( .A(n4950), .ZN(n4945) );
  INV_X1 U5182 ( .A(n5618), .ZN(n5591) );
  INV_X1 U5183 ( .A(n5741), .ZN(n5673) );
  INV_X1 U5184 ( .A(n5633), .ZN(n5737) );
  INV_X1 U5185 ( .A(n4516), .ZN(n5686) );
  INV_X1 U5186 ( .A(n6845), .ZN(n5692) );
  NAND2_X1 U5187 ( .A1(n4625), .A2(n4553), .ZN(n9763) );
  NAND2_X1 U5188 ( .A1(n6845), .A2(n6265), .ZN(n5633) );
  NAND3_X1 U5189 ( .A1(n5132), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4678) );
  INV_X1 U5190 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5132) );
  NAND2_X1 U5191 ( .A1(n4879), .A2(n8481), .ZN(n8298) );
  INV_X1 U5192 ( .A(n4710), .ZN(n4709) );
  OAI21_X1 U5193 ( .B1(n8320), .B2(n8435), .A(n4711), .ZN(n4710) );
  AND2_X1 U5194 ( .A1(n8333), .A2(n8323), .ZN(n4711) );
  AOI21_X1 U5195 ( .B1(n4740), .B2(n4741), .A(n4739), .ZN(n4738) );
  INV_X1 U5196 ( .A(n4742), .ZN(n4741) );
  INV_X1 U5197 ( .A(n5818), .ZN(n4739) );
  AND2_X1 U5198 ( .A1(n6210), .A2(n6211), .ZN(n5109) );
  INV_X1 U5199 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6211) );
  INV_X1 U5200 ( .A(n5451), .ZN(n5012) );
  INV_X1 U5201 ( .A(n5491), .ZN(n5189) );
  INV_X1 U5202 ( .A(SI_15_), .ZN(n5188) );
  INV_X1 U5203 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U5204 ( .A1(n4687), .A2(n4686), .ZN(n7192) );
  INV_X1 U5205 ( .A(n4683), .ZN(n4687) );
  AOI21_X1 U5206 ( .B1(n7288), .B2(n4520), .A(n4684), .ZN(n4683) );
  OR2_X1 U5207 ( .A1(n8722), .A2(n8705), .ZN(n8382) );
  AND2_X1 U5208 ( .A1(n6665), .A2(n6858), .ZN(n7361) );
  OR2_X1 U5209 ( .A1(n8902), .A2(n8174), .ZN(n8415) );
  INV_X1 U5210 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6670) );
  NOR2_X1 U5211 ( .A1(n6097), .A2(n4835), .ZN(n4834) );
  OR2_X1 U5212 ( .A1(n9532), .A2(n5302), .ZN(n5875) );
  OAI22_X1 U5213 ( .A1(n4521), .A2(n5073), .B1(n8067), .B2(n9375), .ZN(n5066)
         );
  INV_X1 U5214 ( .A(n9416), .ZN(n4797) );
  NOR2_X1 U5215 ( .A1(n9563), .A2(n9567), .ZN(n4757) );
  OR2_X1 U5216 ( .A1(n9563), .A2(n9178), .ZN(n8059) );
  NAND2_X1 U5217 ( .A1(n4667), .A2(n7955), .ZN(n4663) );
  INV_X1 U5218 ( .A(n4665), .ZN(n4664) );
  OAI21_X1 U5219 ( .B1(n7954), .B2(n4666), .A(n8043), .ZN(n4665) );
  NAND2_X1 U5220 ( .A1(n5252), .A2(n5251), .ZN(n5722) );
  INV_X1 U5221 ( .A(n5025), .ZN(n5024) );
  AND2_X1 U5222 ( .A1(n5233), .A2(n5232), .ZN(n5341) );
  AND2_X1 U5223 ( .A1(n5228), .A2(n5227), .ZN(n5354) );
  AOI21_X1 U5224 ( .B1(n5001), .B2(n4997), .A(n4610), .ZN(n4996) );
  NAND2_X1 U5225 ( .A1(n5660), .A2(n5119), .ZN(n5169) );
  OAI21_X1 U5226 ( .B1(n5690), .B2(n4993), .A(n4991), .ZN(n5660) );
  AOI21_X1 U5227 ( .B1(n5689), .B2(n4994), .A(n4992), .ZN(n4991) );
  INV_X1 U5228 ( .A(n4994), .ZN(n4993) );
  INV_X1 U5229 ( .A(n5162), .ZN(n4992) );
  AND2_X1 U5230 ( .A1(n7697), .A2(n6705), .ZN(n5107) );
  AND2_X1 U5231 ( .A1(n8449), .A2(n6680), .ZN(n6681) );
  AOI21_X1 U5232 ( .B1(n5100), .B2(n4543), .A(n5099), .ZN(n5098) );
  INV_X1 U5233 ( .A(n6748), .ZN(n5099) );
  NAND2_X1 U5234 ( .A1(n8233), .A2(n4570), .ZN(n8149) );
  INV_X1 U5235 ( .A(n8151), .ZN(n6728) );
  NAND2_X1 U5236 ( .A1(n8445), .A2(n8446), .ZN(n4720) );
  AND2_X1 U5237 ( .A1(n4895), .A2(n4894), .ZN(n8448) );
  AOI21_X1 U5238 ( .B1(n8659), .B2(n6565), .A(n6529), .ZN(n8224) );
  INV_X1 U5239 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6209) );
  XNOR2_X1 U5240 ( .A(n8485), .B(n9938), .ZN(n9947) );
  NAND2_X1 U5241 ( .A1(n4934), .A2(n4935), .ZN(n4933) );
  INV_X1 U5242 ( .A(n8561), .ZN(n4934) );
  INV_X1 U5243 ( .A(n8530), .ZN(n8528) );
  NAND2_X1 U5244 ( .A1(n4582), .A2(n4524), .ZN(n4983) );
  INV_X1 U5245 ( .A(n8657), .ZN(n8635) );
  INV_X1 U5246 ( .A(n6607), .ZN(n4948) );
  NOR2_X1 U5247 ( .A1(n6608), .A2(n4951), .ZN(n4950) );
  INV_X1 U5248 ( .A(n6605), .ZN(n4951) );
  NAND2_X1 U5249 ( .A1(n8405), .A2(n8406), .ZN(n8695) );
  AOI21_X1 U5250 ( .B1(n4958), .B2(n4960), .A(n4606), .ZN(n4956) );
  NAND2_X1 U5251 ( .A1(n8716), .A2(n4958), .ZN(n4957) );
  AND2_X1 U5252 ( .A1(n8354), .A2(n5126), .ZN(n4897) );
  AOI21_X1 U5253 ( .B1(n4969), .B2(n4968), .A(n4598), .ZN(n4967) );
  INV_X1 U5254 ( .A(n4975), .ZN(n4968) );
  INV_X1 U5255 ( .A(n6266), .ZN(n6470) );
  AND2_X1 U5256 ( .A1(n8439), .A2(n6782), .ZN(n8800) );
  INV_X1 U5257 ( .A(n8779), .ZN(n8801) );
  OR2_X1 U5258 ( .A1(n6635), .A2(n8463), .ZN(n10041) );
  NAND2_X1 U5259 ( .A1(n4651), .A2(n4647), .ZN(n5881) );
  AND2_X1 U5260 ( .A1(n4650), .A2(n4648), .ZN(n4647) );
  OR3_X1 U5261 ( .A1(n4751), .A2(n8070), .A3(n4652), .ZN(n4651) );
  AOI21_X1 U5262 ( .B1(n4654), .B2(n4529), .A(n4649), .ZN(n4648) );
  OR2_X1 U5263 ( .A1(n5294), .A2(n7679), .ZN(n4728) );
  INV_X1 U5264 ( .A(n9173), .ZN(n8068) );
  NAND2_X1 U5265 ( .A1(n5875), .A2(n5874), .ZN(n8070) );
  AND2_X1 U5266 ( .A1(n5801), .A2(n8035), .ZN(n8088) );
  OR2_X1 U5267 ( .A1(n9387), .A2(n8064), .ZN(n5071) );
  NAND2_X1 U5268 ( .A1(n9474), .A2(n9470), .ZN(n9463) );
  NOR2_X1 U5269 ( .A1(n4597), .A2(n5048), .ZN(n5047) );
  INV_X1 U5270 ( .A(n5112), .ZN(n5048) );
  NAND2_X1 U5271 ( .A1(n5060), .A2(n5058), .ZN(n9592) );
  NOR2_X1 U5272 ( .A1(n7952), .A2(n5059), .ZN(n5058) );
  INV_X1 U5273 ( .A(n5061), .ZN(n5059) );
  OR2_X1 U5274 ( .A1(n4732), .A2(n9779), .ZN(n4625) );
  AND2_X1 U5275 ( .A1(n6933), .A2(n6932), .ZN(n9765) );
  NAND2_X1 U5276 ( .A1(n5443), .A2(n5442), .ZN(n9588) );
  AND2_X1 U5277 ( .A1(n6162), .A2(n6161), .ZN(n9800) );
  INV_X1 U5278 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5054) );
  INV_X1 U5279 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5290) );
  XNOR2_X1 U5280 ( .A(n5303), .B(n5304), .ZN(n8094) );
  XNOR2_X1 U5281 ( .A(n5329), .B(n5330), .ZN(n8022) );
  NAND2_X1 U5282 ( .A1(n6631), .A2(n6630), .ZN(n8612) );
  OAI21_X1 U5283 ( .B1(n9631), .B2(n6563), .A(n6564), .ZN(n8616) );
  AOI21_X1 U5284 ( .B1(n4738), .B2(n4736), .A(n4807), .ZN(n4735) );
  INV_X1 U5285 ( .A(n4740), .ZN(n4736) );
  INV_X1 U5286 ( .A(n4738), .ZN(n4737) );
  NOR2_X1 U5287 ( .A1(n4632), .A2(n4630), .ZN(n4629) );
  NAND2_X1 U5288 ( .A1(n4805), .A2(n4631), .ZN(n4630) );
  NOR2_X1 U5289 ( .A1(n4599), .A2(n4633), .ZN(n4632) );
  NAND2_X1 U5290 ( .A1(n5906), .A2(n4635), .ZN(n4631) );
  INV_X1 U5291 ( .A(n4629), .ZN(n4628) );
  AND2_X1 U5292 ( .A1(n5879), .A2(n4750), .ZN(n4749) );
  NAND2_X1 U5293 ( .A1(n9357), .A2(n5872), .ZN(n4750) );
  NAND2_X1 U5294 ( .A1(n5074), .A2(n4545), .ZN(n5073) );
  AND2_X1 U5295 ( .A1(n5001), .A2(n5000), .ZN(n4999) );
  INV_X1 U5296 ( .A(n5213), .ZN(n5000) );
  INV_X1 U5297 ( .A(n5463), .ZN(n5192) );
  AND2_X1 U5298 ( .A1(n5032), .A2(n5524), .ZN(n5029) );
  INV_X1 U5299 ( .A(n8451), .ZN(n4896) );
  NAND2_X1 U5300 ( .A1(n7084), .A2(n6998), .ZN(n6999) );
  INV_X1 U5301 ( .A(n7193), .ZN(n4910) );
  AOI21_X1 U5302 ( .B1(n4985), .B2(n4983), .A(n4981), .ZN(n4980) );
  INV_X1 U5303 ( .A(n8430), .ZN(n4981) );
  INV_X1 U5304 ( .A(n4983), .ZN(n4982) );
  INV_X1 U5305 ( .A(n4955), .ZN(n4954) );
  OAI21_X1 U5306 ( .B1(n6584), .B2(n8476), .A(n7770), .ZN(n4955) );
  AND2_X1 U5307 ( .A1(n10030), .A2(n8476), .ZN(n8335) );
  INV_X1 U5308 ( .A(n8437), .ZN(n8432) );
  OR2_X1 U5309 ( .A1(n8908), .A2(n8205), .ZN(n8411) );
  OR2_X1 U5310 ( .A1(n8708), .A2(n6740), .ZN(n8399) );
  AND2_X1 U5311 ( .A1(n8344), .A2(n8328), .ZN(n7801) );
  OR2_X1 U5312 ( .A1(n7973), .A2(n7802), .ZN(n8345) );
  NAND2_X1 U5313 ( .A1(n6235), .A2(n4964), .ZN(n4963) );
  INV_X1 U5314 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6235) );
  INV_X1 U5315 ( .A(n6356), .ZN(n4714) );
  OR2_X1 U5316 ( .A1(n6439), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U5317 ( .A1(n6378), .A2(n5109), .ZN(n6415) );
  NAND2_X1 U5318 ( .A1(n9128), .A2(n4596), .ZN(n4867) );
  NAND2_X1 U5319 ( .A1(n4868), .A2(n4865), .ZN(n4864) );
  INV_X1 U5320 ( .A(n9128), .ZN(n4865) );
  INV_X1 U5321 ( .A(n4596), .ZN(n4868) );
  NOR2_X1 U5322 ( .A1(n4857), .A2(n6054), .ZN(n4856) );
  INV_X1 U5323 ( .A(n7729), .ZN(n4857) );
  CLKBUF_X1 U5324 ( .A(n6066), .Z(n6135) );
  NOR2_X1 U5325 ( .A1(n5750), .A2(n5749), .ZN(n5924) );
  INV_X1 U5326 ( .A(n8070), .ZN(n4776) );
  AOI21_X1 U5327 ( .B1(n4781), .B2(n4784), .A(n5314), .ZN(n4780) );
  NOR2_X1 U5328 ( .A1(n8038), .A2(n4549), .ZN(n4781) );
  INV_X1 U5329 ( .A(n5073), .ZN(n5068) );
  OR2_X1 U5330 ( .A1(n9543), .A2(n5328), .ZN(n5870) );
  INV_X1 U5331 ( .A(n4792), .ZN(n4791) );
  NOR2_X1 U5332 ( .A1(n4794), .A2(n4793), .ZN(n4792) );
  INV_X1 U5333 ( .A(n8032), .ZN(n4793) );
  INV_X1 U5334 ( .A(n4585), .ZN(n4794) );
  NOR2_X1 U5335 ( .A1(n9659), .A2(n9521), .ZN(n9494) );
  INV_X1 U5336 ( .A(n9735), .ZN(n4763) );
  INV_X1 U5337 ( .A(n7713), .ZN(n5043) );
  NOR2_X1 U5338 ( .A1(n5644), .A2(n5043), .ZN(n5040) );
  INV_X1 U5339 ( .A(n7778), .ZN(n6186) );
  OAI22_X1 U5340 ( .A1(n9592), .A2(n4661), .B1(n4660), .B2(n4664), .ZN(n9658)
         );
  NAND2_X1 U5341 ( .A1(n9655), .A2(n4662), .ZN(n4661) );
  INV_X1 U5342 ( .A(n4663), .ZN(n4662) );
  NAND2_X1 U5343 ( .A1(n5007), .A2(n5005), .ZN(n5413) );
  AND2_X1 U5344 ( .A1(n5006), .A2(n5203), .ZN(n5005) );
  INV_X1 U5345 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4870) );
  INV_X1 U5346 ( .A(n5033), .ZN(n5032) );
  OAI21_X1 U5347 ( .B1(n5036), .B2(n5034), .A(n5177), .ZN(n5033) );
  NAND2_X1 U5348 ( .A1(n5035), .A2(n5171), .ZN(n5034) );
  INV_X1 U5349 ( .A(n5539), .ZN(n5035) );
  NAND2_X1 U5350 ( .A1(n4986), .A2(n4988), .ZN(n5602) );
  AOI21_X1 U5351 ( .B1(n5648), .B2(n4989), .A(n4580), .ZN(n4988) );
  INV_X1 U5352 ( .A(n5149), .ZN(n4989) );
  OAI21_X1 U5353 ( .B1(n6265), .B2(P1_DATAO_REG_5__SCAN_IN), .A(n4622), .ZN(
        n5150) );
  NAND2_X1 U5354 ( .A1(n6265), .A2(n6826), .ZN(n4622) );
  OAI21_X1 U5355 ( .B1(n6814), .B2(P2_DATAO_REG_4__SCAN_IN), .A(n4811), .ZN(
        n5147) );
  NAND2_X1 U5356 ( .A1(n5089), .A2(n5088), .ZN(n5087) );
  INV_X1 U5357 ( .A(n8219), .ZN(n5088) );
  INV_X1 U5358 ( .A(n5087), .ZN(n5086) );
  NAND2_X1 U5359 ( .A1(n6254), .A2(n7369), .ZN(n6980) );
  INV_X1 U5360 ( .A(n8482), .ZN(n6254) );
  AOI21_X1 U5361 ( .B1(n5077), .B2(n7410), .A(n4558), .ZN(n5076) );
  INV_X1 U5362 ( .A(n7410), .ZN(n5078) );
  NAND2_X1 U5363 ( .A1(n5090), .A2(n5103), .ZN(n5089) );
  INV_X1 U5364 ( .A(n5095), .ZN(n5090) );
  AOI21_X1 U5365 ( .B1(n5098), .B2(n5101), .A(n5096), .ZN(n5095) );
  INV_X1 U5366 ( .A(n8142), .ZN(n5096) );
  INV_X1 U5367 ( .A(n5103), .ZN(n5093) );
  INV_X1 U5368 ( .A(n5098), .ZN(n5097) );
  AND2_X1 U5369 ( .A1(n4909), .A2(n7212), .ZN(n7317) );
  OR2_X1 U5370 ( .A1(n7324), .A2(n7323), .ZN(n7433) );
  XNOR2_X1 U5371 ( .A(n8491), .B(n9938), .ZN(n9940) );
  NAND2_X1 U5372 ( .A1(n4921), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4920) );
  NAND2_X1 U5373 ( .A1(n8486), .A2(n4921), .ZN(n4919) );
  INV_X1 U5374 ( .A(n9964), .ZN(n4921) );
  NAND2_X1 U5375 ( .A1(n6668), .A2(n6667), .ZN(n6947) );
  OAI21_X1 U5376 ( .B1(n8487), .B2(n4923), .A(n4922), .ZN(n9984) );
  NAND2_X1 U5377 ( .A1(n4924), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4923) );
  NAND2_X1 U5378 ( .A1(n8524), .A2(n4924), .ZN(n4922) );
  INV_X1 U5379 ( .A(n9985), .ZN(n4924) );
  OR2_X1 U5380 ( .A1(n8526), .A2(n8566), .ZN(n8561) );
  OR2_X1 U5381 ( .A1(n6554), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8614) );
  OR2_X1 U5382 ( .A1(n6505), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6514) );
  AND3_X1 U5383 ( .A1(n6486), .A2(n6485), .A3(n6484), .ZN(n8705) );
  AND2_X1 U5384 ( .A1(n8731), .A2(n6603), .ZN(n8716) );
  NAND2_X1 U5385 ( .A1(n8716), .A2(n8715), .ZN(n8714) );
  AOI21_X1 U5386 ( .B1(n8750), .B2(n8379), .A(n4907), .ZN(n4906) );
  INV_X1 U5387 ( .A(n8393), .ZN(n4907) );
  INV_X1 U5388 ( .A(n8474), .ZN(n7740) );
  NAND2_X1 U5389 ( .A1(n7605), .A2(n10008), .ZN(n4938) );
  NAND2_X1 U5390 ( .A1(n7592), .A2(n4564), .ZN(n4939) );
  OR2_X1 U5391 ( .A1(n7367), .A2(n7366), .ZN(n7368) );
  XNOR2_X1 U5392 ( .A(n8879), .B(n8468), .ZN(n8622) );
  INV_X1 U5393 ( .A(n8800), .ZN(n8748) );
  NOR2_X1 U5394 ( .A1(n4900), .A2(n8288), .ZN(n4899) );
  INV_X1 U5395 ( .A(n8420), .ZN(n4900) );
  XNOR2_X1 U5396 ( .A(n8884), .B(n8624), .ZN(n8633) );
  OR2_X1 U5397 ( .A1(n8288), .A2(n8289), .ZN(n8646) );
  OR2_X1 U5398 ( .A1(n8896), .A2(n8224), .ZN(n8420) );
  INV_X1 U5399 ( .A(n8646), .ZN(n8643) );
  NAND2_X1 U5400 ( .A1(n8742), .A2(n4940), .ZN(n8731) );
  NOR2_X1 U5401 ( .A1(n8736), .A2(n4941), .ZN(n4940) );
  INV_X1 U5402 ( .A(n6602), .ZN(n4941) );
  OR2_X1 U5403 ( .A1(n8854), .A2(n8164), .ZN(n8735) );
  AOI21_X1 U5404 ( .B1(n4889), .B2(n4887), .A(n4886), .ZN(n4885) );
  AND2_X1 U5405 ( .A1(n4891), .A2(n8373), .ZN(n4889) );
  OR2_X1 U5406 ( .A1(n8435), .A2(n6782), .ZN(n8779) );
  AND2_X1 U5407 ( .A1(n8386), .A2(n8373), .ZN(n8784) );
  AOI21_X1 U5408 ( .B1(n4541), .B2(n7984), .A(n4892), .ZN(n4891) );
  INV_X1 U5409 ( .A(n8387), .ZN(n4892) );
  NAND2_X1 U5410 ( .A1(n6428), .A2(n6427), .ZN(n8007) );
  INV_X1 U5411 ( .A(n8362), .ZN(n4971) );
  OR2_X1 U5412 ( .A1(n8012), .A2(n8197), .ZN(n8354) );
  NAND2_X1 U5413 ( .A1(n7897), .A2(n8352), .ZN(n4898) );
  NOR2_X1 U5414 ( .A1(n6594), .A2(n4976), .ZN(n4975) );
  INV_X1 U5415 ( .A(n6592), .ZN(n4976) );
  NAND2_X1 U5416 ( .A1(n4974), .A2(n8197), .ZN(n4973) );
  NAND2_X1 U5417 ( .A1(n4884), .A2(n6367), .ZN(n4883) );
  INV_X1 U5418 ( .A(n7738), .ZN(n4884) );
  AND3_X1 U5419 ( .A1(n6320), .A2(n6319), .A3(n6318), .ZN(n10012) );
  INV_X1 U5420 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6641) );
  XNOR2_X1 U5421 ( .A(n6671), .B(n6670), .ZN(n6945) );
  NAND2_X1 U5422 ( .A1(n6614), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6615) );
  NAND2_X1 U5423 ( .A1(n8955), .A2(n6203), .ZN(n4916) );
  NAND2_X1 U5424 ( .A1(n6113), .A2(n4826), .ZN(n4824) );
  AOI21_X1 U5425 ( .B1(n4823), .B2(n4822), .A(n4821), .ZN(n4820) );
  INV_X1 U5426 ( .A(n9149), .ZN(n4821) );
  INV_X1 U5427 ( .A(n9072), .ZN(n4822) );
  INV_X1 U5428 ( .A(n4824), .ZN(n4823) );
  NAND2_X1 U5429 ( .A1(n4817), .A2(n4819), .ZN(n4816) );
  INV_X1 U5430 ( .A(n4820), .ZN(n4817) );
  INV_X1 U5431 ( .A(n4834), .ZN(n4832) );
  AOI21_X1 U5432 ( .B1(n4834), .B2(n4831), .A(n4578), .ZN(n4830) );
  INV_X1 U5433 ( .A(n4544), .ZN(n4831) );
  NAND2_X1 U5434 ( .A1(n5279), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5430) );
  INV_X1 U5435 ( .A(n5445), .ZN(n5279) );
  INV_X1 U5436 ( .A(n9140), .ZN(n4875) );
  NOR2_X1 U5437 ( .A1(n4836), .A2(n8993), .ZN(n4835) );
  INV_X1 U5438 ( .A(n8994), .ZN(n4836) );
  NAND2_X1 U5439 ( .A1(n8097), .A2(n7471), .ZN(n6929) );
  NOR2_X1 U5440 ( .A1(n9286), .A2(n9285), .ZN(n9291) );
  NAND2_X1 U5441 ( .A1(n9375), .A2(n8036), .ZN(n4784) );
  OR2_X1 U5442 ( .A1(n8038), .A2(n5314), .ZN(n9361) );
  INV_X1 U5443 ( .A(n8063), .ZN(n5070) );
  OR2_X1 U5444 ( .A1(n9557), .A2(n8061), .ZN(n9392) );
  NAND2_X1 U5445 ( .A1(n4668), .A2(n4669), .ZN(n9387) );
  AOI21_X1 U5446 ( .B1(n4675), .B2(n4670), .A(n4532), .ZN(n4669) );
  AOI21_X1 U5447 ( .B1(n5051), .B2(n5050), .A(n4574), .ZN(n5049) );
  INV_X1 U5448 ( .A(n8058), .ZN(n5050) );
  NAND2_X1 U5449 ( .A1(n4535), .A2(n4585), .ZN(n4799) );
  NAND2_X1 U5450 ( .A1(n9450), .A2(n4792), .ZN(n4798) );
  AND2_X1 U5451 ( .A1(n8031), .A2(n5834), .ZN(n9459) );
  OAI22_X1 U5452 ( .A1(n9504), .A2(n4785), .B1(n4786), .B2(n5771), .ZN(n9460)
         );
  NAND2_X1 U5453 ( .A1(n5838), .A2(n5915), .ZN(n4785) );
  INV_X1 U5454 ( .A(n4787), .ZN(n4786) );
  INV_X1 U5455 ( .A(n9459), .ZN(n9456) );
  NAND2_X1 U5456 ( .A1(n9494), .A2(n9501), .ZN(n9495) );
  OR2_X1 U5457 ( .A1(n9501), .A2(n8049), .ZN(n5112) );
  AND2_X1 U5458 ( .A1(n5833), .A2(n5915), .ZN(n9479) );
  OR2_X1 U5459 ( .A1(n9588), .A2(n9183), .ZN(n8048) );
  OR2_X1 U5460 ( .A1(n9521), .A2(n8047), .ZN(n9489) );
  NAND2_X1 U5461 ( .A1(n9504), .A2(n4789), .ZN(n9487) );
  NAND2_X1 U5462 ( .A1(n5277), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5504) );
  OR2_X1 U5463 ( .A1(n9735), .A2(n5490), .ZN(n7947) );
  NAND2_X1 U5464 ( .A1(n5062), .A2(n5710), .ZN(n5061) );
  NAND2_X1 U5465 ( .A1(n7831), .A2(n4571), .ZN(n5060) );
  OR2_X1 U5466 ( .A1(n9897), .A2(n5711), .ZN(n7812) );
  NAND2_X1 U5467 ( .A1(n7827), .A2(n4659), .ZN(n7830) );
  NAND2_X1 U5468 ( .A1(n7829), .A2(n7828), .ZN(n4659) );
  AND2_X1 U5469 ( .A1(n5818), .A2(n5904), .ZN(n7832) );
  AOI21_X1 U5470 ( .B1(n5895), .B2(n4731), .A(n4550), .ZN(n4730) );
  INV_X1 U5471 ( .A(n5757), .ZN(n4731) );
  OAI21_X1 U5472 ( .B1(n7641), .B2(n5755), .A(n5891), .ZN(n9779) );
  OR2_X1 U5473 ( .A1(n9901), .A2(n6186), .ZN(n6926) );
  OR2_X1 U5474 ( .A1(n4768), .A2(n9353), .ZN(n4767) );
  INV_X1 U5475 ( .A(n4769), .ZN(n4768) );
  AOI21_X1 U5476 ( .B1(n9364), .B2(n9532), .A(n9600), .ZN(n4769) );
  INV_X1 U5477 ( .A(n7113), .ZN(n9844) );
  INV_X1 U5478 ( .A(n7472), .ZN(n7674) );
  INV_X1 U5479 ( .A(n9765), .ZN(n9782) );
  NOR2_X1 U5480 ( .A1(n8002), .A2(n7965), .ZN(n5948) );
  NAND2_X1 U5481 ( .A1(n5724), .A2(n5723), .ZN(n5736) );
  XNOR2_X1 U5482 ( .A(n5736), .B(n5735), .ZN(n8248) );
  XNOR2_X1 U5483 ( .A(n5315), .B(n5316), .ZN(n8096) );
  INV_X1 U5484 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U5485 ( .A1(n5884), .A2(n5063), .ZN(n5288) );
  NAND2_X1 U5486 ( .A1(n5941), .A2(n5943), .ZN(n5944) );
  NAND2_X1 U5487 ( .A1(n5023), .A2(n5228), .ZN(n5342) );
  NAND2_X1 U5488 ( .A1(n5355), .A2(n5354), .ZN(n5023) );
  OAI21_X1 U5489 ( .B1(n5377), .B2(n5376), .A(n5218), .ZN(n5366) );
  AND2_X1 U5490 ( .A1(n5222), .A2(n5221), .ZN(n5365) );
  XNOR2_X1 U5491 ( .A(n5934), .B(n5933), .ZN(n6842) );
  OAI21_X1 U5492 ( .B1(n5210), .B2(n5003), .A(n5001), .ZN(n5399) );
  NAND2_X1 U5493 ( .A1(n5004), .A2(n5008), .ZN(n5439) );
  OR2_X1 U5494 ( .A1(n5493), .A2(n5011), .ZN(n5004) );
  NAND2_X1 U5495 ( .A1(n5013), .A2(n5015), .ZN(n5452) );
  NAND2_X1 U5496 ( .A1(n5493), .A2(n5018), .ZN(n5013) );
  NAND2_X1 U5497 ( .A1(n5512), .A2(n4871), .ZN(n5466) );
  NAND2_X1 U5498 ( .A1(n5014), .A2(n5190), .ZN(n5465) );
  NAND2_X1 U5499 ( .A1(n5031), .A2(n5171), .ZN(n5540) );
  NAND2_X1 U5500 ( .A1(n5169), .A2(n5036), .ZN(n5031) );
  XNOR2_X1 U5501 ( .A(n5147), .B(SI_4_), .ZN(n5585) );
  NAND2_X1 U5502 ( .A1(n7503), .A2(n5107), .ZN(n7696) );
  NAND2_X1 U5503 ( .A1(n5075), .A2(n6691), .ZN(n7248) );
  INV_X1 U5504 ( .A(n7247), .ZN(n6692) );
  AOI21_X1 U5505 ( .B1(n4525), .B2(n5082), .A(n4602), .ZN(n5080) );
  AND2_X1 U5506 ( .A1(n6553), .A2(n6552), .ZN(n6788) );
  AND4_X1 U5507 ( .A1(n6435), .A2(n6434), .A3(n6433), .A4(n6432), .ZN(n8778)
         );
  NAND2_X1 U5508 ( .A1(n6480), .A2(n6479), .ZN(n8722) );
  INV_X1 U5509 ( .A(n8696), .ZN(n8205) );
  AND4_X1 U5510 ( .A1(n6458), .A2(n6457), .A3(n6456), .A4(n6455), .ZN(n8749)
         );
  AND2_X1 U5511 ( .A1(n6764), .A2(n8674), .ZN(n8245) );
  NAND2_X1 U5512 ( .A1(n6760), .A2(n6759), .ZN(n8232) );
  XNOR2_X1 U5513 ( .A(n6228), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8463) );
  INV_X1 U5514 ( .A(n8636), .ZN(n8468) );
  NAND2_X1 U5515 ( .A1(n6550), .A2(n6549), .ZN(n8647) );
  NAND2_X1 U5516 ( .A1(n6520), .A2(n6519), .ZN(n8685) );
  INV_X1 U5517 ( .A(n8705), .ZN(n8732) );
  INV_X1 U5518 ( .A(n8749), .ZN(n8787) );
  INV_X1 U5519 ( .A(n7802), .ZN(n8473) );
  XNOR2_X1 U5520 ( .A(n7099), .B(n6995), .ZN(n7086) );
  OR2_X1 U5521 ( .A1(n6994), .A2(n8540), .ZN(n9986) );
  NAND2_X1 U5522 ( .A1(n4933), .A2(n8583), .ZN(n4928) );
  AND2_X1 U5523 ( .A1(n4933), .A2(n4621), .ZN(n4926) );
  INV_X1 U5524 ( .A(n8592), .ZN(n4931) );
  NAND2_X1 U5525 ( .A1(n8528), .A2(n4617), .ZN(n4930) );
  AND2_X1 U5526 ( .A1(n8611), .A2(n9997), .ZN(n4937) );
  INV_X1 U5527 ( .A(n6788), .ZN(n8879) );
  NAND2_X1 U5528 ( .A1(n4949), .A2(n6607), .ZN(n8670) );
  NAND2_X1 U5529 ( .A1(n6606), .A2(n4950), .ZN(n4949) );
  NAND2_X1 U5530 ( .A1(n6405), .A2(n6404), .ZN(n8358) );
  INV_X1 U5531 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6217) );
  INV_X1 U5532 ( .A(n9153), .ZN(n9702) );
  NAND2_X1 U5533 ( .A1(n5393), .A2(n5392), .ZN(n9578) );
  NAND2_X1 U5534 ( .A1(n5379), .A2(n5378), .ZN(n9567) );
  AND2_X1 U5535 ( .A1(n6182), .A2(n6180), .ZN(n6184) );
  NAND2_X1 U5536 ( .A1(n5332), .A2(n5331), .ZN(n9546) );
  NOR2_X2 U5537 ( .A1(n6189), .A2(n6179), .ZN(n9096) );
  OAI21_X1 U5538 ( .B1(n4748), .B2(n4746), .A(n4620), .ZN(n4745) );
  NAND2_X1 U5539 ( .A1(n4747), .A2(n5872), .ZN(n4746) );
  NOR2_X1 U5540 ( .A1(n5881), .A2(n8097), .ZN(n4748) );
  NAND2_X1 U5541 ( .A1(n5340), .A2(n5339), .ZN(n9175) );
  OR2_X1 U5542 ( .A1(n5741), .A2(n5605), .ZN(n5606) );
  OR2_X1 U5543 ( .A1(n5743), .A2(n9920), .ZN(n5607) );
  OR2_X1 U5544 ( .A1(n5743), .A2(n9710), .ZN(n5567) );
  NOR2_X1 U5545 ( .A1(n7621), .A2(n7620), .ZN(n7854) );
  OR2_X1 U5546 ( .A1(n9340), .A2(n9727), .ZN(n4701) );
  AOI21_X1 U5547 ( .B1(n9341), .B2(n9720), .A(n9724), .ZN(n4700) );
  OAI21_X1 U5548 ( .B1(n9344), .B2(n5131), .A(n9343), .ZN(n4698) );
  NAND2_X1 U5549 ( .A1(n4778), .A2(n8070), .ZN(n4777) );
  NAND2_X1 U5550 ( .A1(n5516), .A2(n5515), .ZN(n9125) );
  AOI21_X1 U5551 ( .B1(n9800), .B2(n6165), .A(n6164), .ZN(n9620) );
  NAND2_X1 U5552 ( .A1(n5960), .A2(n6808), .ZN(n9833) );
  INV_X1 U5553 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9622) );
  AND3_X1 U5554 ( .A1(n4528), .A2(n5290), .A3(n5259), .ZN(n4752) );
  NAND2_X1 U5555 ( .A1(n5256), .A2(n5724), .ZN(n9631) );
  CLKBUF_X1 U5556 ( .A(n5959), .Z(n8097) );
  AND2_X1 U5557 ( .A1(n4744), .A2(n4743), .ZN(n4742) );
  NAND2_X1 U5558 ( .A1(n7779), .A2(n5816), .ZN(n4743) );
  AND2_X1 U5559 ( .A1(n7812), .A2(n5900), .ZN(n4744) );
  AOI21_X1 U5560 ( .B1(n4742), .B2(n5765), .A(n4575), .ZN(n4740) );
  INV_X1 U5561 ( .A(n5904), .ZN(n4635) );
  NAND2_X1 U5562 ( .A1(n8341), .A2(n4708), .ZN(n8349) );
  NAND2_X1 U5563 ( .A1(n4712), .A2(n4709), .ZN(n4708) );
  AOI21_X1 U5564 ( .B1(n4735), .B2(n4737), .A(n4583), .ZN(n4734) );
  OAI21_X1 U5565 ( .B1(n4628), .B2(n4634), .A(n5907), .ZN(n4627) );
  AND2_X1 U5566 ( .A1(n5837), .A2(n9489), .ZN(n5840) );
  AOI21_X1 U5567 ( .B1(n4645), .B2(n4646), .A(n4642), .ZN(n4641) );
  INV_X1 U5568 ( .A(n5848), .ZN(n4642) );
  NOR2_X1 U5569 ( .A1(n4522), .A2(n5872), .ZN(n4646) );
  INV_X1 U5570 ( .A(n5038), .ZN(n5627) );
  AOI21_X1 U5571 ( .B1(n4641), .B2(n5849), .A(n9427), .ZN(n4639) );
  INV_X1 U5572 ( .A(n4641), .ZN(n4640) );
  INV_X1 U5573 ( .A(n5228), .ZN(n5026) );
  NAND2_X1 U5574 ( .A1(n4685), .A2(n4688), .ZN(n4684) );
  NAND2_X1 U5575 ( .A1(n7289), .A2(n4520), .ZN(n4685) );
  AND2_X1 U5576 ( .A1(n8437), .A2(n8599), .ZN(n6768) );
  NAND2_X1 U5577 ( .A1(n6207), .A2(n6206), .ZN(n6208) );
  INV_X1 U5578 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6206) );
  NOR2_X1 U5579 ( .A1(n5022), .A2(n5026), .ZN(n5021) );
  INV_X1 U5580 ( .A(n5222), .ZN(n5022) );
  OAI21_X1 U5581 ( .B1(n5354), .B2(n5026), .A(n5341), .ZN(n5025) );
  NOR2_X1 U5582 ( .A1(n5213), .A2(n4998), .ZN(n4997) );
  INV_X1 U5583 ( .A(n5003), .ZN(n4998) );
  INV_X1 U5584 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5200) );
  INV_X1 U5585 ( .A(SI_17_), .ZN(n5195) );
  NOR2_X1 U5586 ( .A1(n5681), .A2(n4572), .ZN(n4994) );
  AND2_X1 U5587 ( .A1(n5648), .A2(n5585), .ZN(n4987) );
  INV_X1 U5588 ( .A(n6683), .ZN(n6701) );
  INV_X1 U5589 ( .A(n6699), .ZN(n5077) );
  NOR2_X1 U5590 ( .A1(n4543), .A2(n8202), .ZN(n5102) );
  NAND2_X1 U5591 ( .A1(n8869), .A2(n8285), .ZN(n4894) );
  AOI21_X1 U5592 ( .B1(n4723), .B2(n4563), .A(n4721), .ZN(n8453) );
  NAND2_X1 U5593 ( .A1(n4722), .A2(n8428), .ZN(n4721) );
  OAI21_X1 U5594 ( .B1(n7049), .B2(n10464), .A(n7157), .ZN(n7033) );
  AOI21_X1 U5595 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n8484), .A(n8483), .ZN(
        n8485) );
  OAI21_X1 U5596 ( .B1(n8537), .B2(n10226), .A(n9974), .ZN(n8553) );
  INV_X1 U5597 ( .A(n8559), .ZN(n4935) );
  OR2_X1 U5598 ( .A1(n8616), .A2(n8625), .ZN(n8451) );
  INV_X1 U5599 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6360) );
  INV_X1 U5600 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7195) );
  AND2_X1 U5601 ( .A1(n6348), .A2(n7195), .ZN(n6361) );
  NOR2_X1 U5602 ( .A1(n6335), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6348) );
  INV_X1 U5603 ( .A(n4959), .ZN(n4958) );
  OAI21_X1 U5604 ( .B1(n8715), .B2(n4960), .A(n8706), .ZN(n4959) );
  INV_X1 U5605 ( .A(n6604), .ZN(n4960) );
  INV_X1 U5606 ( .A(n4541), .ZN(n4887) );
  INV_X1 U5607 ( .A(n8343), .ZN(n4882) );
  NAND2_X1 U5608 ( .A1(n6355), .A2(n8327), .ZN(n7738) );
  AND2_X1 U5609 ( .A1(n6354), .A2(n8332), .ZN(n4908) );
  NOR2_X1 U5610 ( .A1(n6666), .A2(n7361), .ZN(n6775) );
  INV_X1 U5611 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6637) );
  NOR2_X1 U5612 ( .A1(n4863), .A2(n4860), .ZN(n4859) );
  INV_X1 U5613 ( .A(n4867), .ZN(n4860) );
  INV_X1 U5614 ( .A(n9005), .ZN(n4863) );
  INV_X1 U5615 ( .A(n4864), .ZN(n4862) );
  NAND2_X1 U5616 ( .A1(n4842), .A2(n4514), .ZN(n4841) );
  NAND2_X1 U5617 ( .A1(n5999), .A2(n5963), .ZN(n4847) );
  INV_X1 U5618 ( .A(n8971), .ZN(n4846) );
  AND2_X1 U5619 ( .A1(n5963), .A2(n9789), .ZN(n4840) );
  INV_X1 U5620 ( .A(n6066), .ZN(n5985) );
  NOR2_X1 U5621 ( .A1(n4855), .A2(n4850), .ZN(n4849) );
  INV_X1 U5622 ( .A(n6029), .ZN(n4850) );
  INV_X1 U5623 ( .A(n6053), .ZN(n4855) );
  AOI21_X1 U5624 ( .B1(n4854), .B2(n6053), .A(n4853), .ZN(n4852) );
  INV_X1 U5625 ( .A(n6061), .ZN(n4853) );
  INV_X1 U5626 ( .A(n4856), .ZN(n4854) );
  NOR2_X1 U5627 ( .A1(n5880), .A2(n4655), .ZN(n4654) );
  NOR2_X1 U5628 ( .A1(n9357), .A2(n5872), .ZN(n4655) );
  NAND2_X1 U5629 ( .A1(n9524), .A2(n5878), .ZN(n5880) );
  INV_X1 U5630 ( .A(n4581), .ZN(n4649) );
  NOR2_X1 U5631 ( .A1(n4749), .A2(n4654), .ZN(n4652) );
  NAND2_X1 U5632 ( .A1(n4749), .A2(n4557), .ZN(n4650) );
  NAND2_X1 U5633 ( .A1(n4784), .A2(n4783), .ZN(n4782) );
  INV_X1 U5634 ( .A(n9175), .ZN(n8065) );
  INV_X1 U5635 ( .A(n5049), .ZN(n4671) );
  NOR2_X1 U5636 ( .A1(n9557), .A2(n4756), .ZN(n4755) );
  INV_X1 U5637 ( .A(n4757), .ZN(n4756) );
  OR2_X1 U5638 ( .A1(n5382), .A2(n9009), .ZN(n5370) );
  OR2_X1 U5639 ( .A1(n9578), .A2(n9181), .ZN(n8052) );
  OAI21_X1 U5640 ( .B1(n4789), .B2(n4788), .A(n9479), .ZN(n4787) );
  NOR2_X1 U5641 ( .A1(n9051), .A2(n9125), .ZN(n4764) );
  AND2_X1 U5642 ( .A1(n7947), .A2(n5821), .ZN(n5819) );
  AND2_X1 U5643 ( .A1(n6931), .A2(n6186), .ZN(n6843) );
  NAND2_X1 U5644 ( .A1(n7834), .A2(n5062), .ZN(n7876) );
  NAND2_X1 U5645 ( .A1(n5959), .A2(n6931), .ZN(n6928) );
  INV_X1 U5646 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n4624) );
  INV_X1 U5647 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4623) );
  AND2_X1 U5648 ( .A1(n5251), .A2(n5250), .ZN(n5304) );
  AND2_X1 U5649 ( .A1(n5239), .A2(n5238), .ZN(n5330) );
  NOR2_X1 U5650 ( .A1(n5211), .A2(n10270), .ZN(n5003) );
  AOI21_X1 U5651 ( .B1(n4611), .B2(n5211), .A(n5002), .ZN(n5001) );
  NOR2_X1 U5652 ( .A1(n5209), .A2(SI_20_), .ZN(n5002) );
  AOI21_X1 U5653 ( .B1(n4546), .B2(n5010), .A(n5009), .ZN(n5008) );
  INV_X1 U5654 ( .A(n5199), .ZN(n5009) );
  INV_X1 U5655 ( .A(n5018), .ZN(n5010) );
  INV_X1 U5656 ( .A(n4546), .ZN(n5011) );
  NOR2_X1 U5657 ( .A1(n5194), .A2(n5019), .ZN(n5018) );
  INV_X1 U5658 ( .A(n5190), .ZN(n5019) );
  INV_X1 U5659 ( .A(n5016), .ZN(n5015) );
  OAI21_X1 U5660 ( .B1(n5017), .B2(n5194), .A(n5193), .ZN(n5016) );
  NAND2_X1 U5661 ( .A1(n5191), .A2(n5190), .ZN(n5017) );
  NOR2_X1 U5662 ( .A1(n4530), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n4871) );
  AOI21_X1 U5663 ( .B1(n5029), .B2(n5034), .A(n4579), .ZN(n5027) );
  NOR2_X1 U5664 ( .A1(n5172), .A2(n5037), .ZN(n5036) );
  INV_X1 U5665 ( .A(n5168), .ZN(n5037) );
  NOR2_X1 U5666 ( .A1(n5597), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5661) );
  NOR2_X2 U5667 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5582) );
  NAND2_X1 U5668 ( .A1(n6814), .A2(n6816), .ZN(n4677) );
  INV_X1 U5669 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5130) );
  XNOR2_X1 U5670 ( .A(n6253), .B(n4964), .ZN(n6626) );
  NAND2_X1 U5671 ( .A1(n6648), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6253) );
  OR2_X1 U5672 ( .A1(n8158), .A2(n5082), .ZN(n5081) );
  INV_X1 U5673 ( .A(n6732), .ZN(n5082) );
  INV_X1 U5674 ( .A(n8193), .ZN(n6720) );
  XNOR2_X1 U5675 ( .A(n6683), .B(n4879), .ZN(n6688) );
  NAND2_X1 U5676 ( .A1(n6730), .A2(n8158), .ZN(n8161) );
  AND4_X1 U5677 ( .A1(n6469), .A2(n6468), .A3(n6467), .A4(n6466), .ZN(n8164)
         );
  NAND2_X1 U5678 ( .A1(n8253), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6282) );
  NAND2_X1 U5679 ( .A1(n4682), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7127) );
  INV_X1 U5680 ( .A(n7125), .ZN(n4682) );
  NAND2_X1 U5681 ( .A1(n4914), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4913) );
  NAND2_X1 U5682 ( .A1(n4915), .A2(n7051), .ZN(n4914) );
  INV_X1 U5683 ( .A(n6999), .ZN(n4915) );
  NAND2_X1 U5684 ( .A1(n6999), .A2(n7029), .ZN(n7151) );
  NAND2_X1 U5685 ( .A1(n7271), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7290) );
  INV_X1 U5686 ( .A(n7192), .ZN(n7042) );
  AND2_X1 U5687 ( .A1(n4540), .A2(n4689), .ZN(n7040) );
  NOR2_X1 U5688 ( .A1(n7044), .A2(n7043), .ZN(n7191) );
  NAND2_X1 U5689 ( .A1(n7202), .A2(n7203), .ZN(n7207) );
  NAND2_X1 U5690 ( .A1(n7327), .A2(n7328), .ZN(n7330) );
  AND2_X1 U5691 ( .A1(n7433), .A2(n7432), .ZN(n7557) );
  NAND2_X1 U5692 ( .A1(n9940), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9939) );
  NOR2_X1 U5693 ( .A1(n9947), .A2(n10217), .ZN(n9946) );
  XNOR2_X1 U5694 ( .A(n8531), .B(n8522), .ZN(n8493) );
  NAND2_X1 U5695 ( .A1(n8493), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8533) );
  NOR2_X1 U5696 ( .A1(n9984), .A2(n4693), .ZN(n8526) );
  AND2_X1 U5697 ( .A1(n9994), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4693) );
  INV_X1 U5698 ( .A(n6626), .ZN(n8591) );
  AND2_X1 U5699 ( .A1(n8259), .A2(n6624), .ZN(n8436) );
  AOI21_X1 U5700 ( .B1(n4980), .B2(n4982), .A(n4577), .ZN(n4978) );
  AND2_X1 U5701 ( .A1(n6524), .A2(n8143), .ZN(n6532) );
  OR2_X1 U5702 ( .A1(n6497), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6505) );
  AND2_X1 U5703 ( .A1(n8382), .A2(n8379), .ZN(n4905) );
  OAI21_X1 U5704 ( .B1(n4906), .B2(n4904), .A(n8397), .ZN(n4903) );
  INV_X1 U5705 ( .A(n8382), .ZN(n4904) );
  NOR2_X1 U5706 ( .A1(n6481), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6489) );
  NAND2_X1 U5707 ( .A1(n6464), .A2(n6463), .ZN(n6473) );
  AND2_X1 U5708 ( .A1(n8735), .A2(n8392), .ZN(n8745) );
  NOR2_X1 U5709 ( .A1(n6429), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6444) );
  OR2_X1 U5710 ( .A1(n6418), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6429) );
  NOR2_X1 U5711 ( .A1(n6396), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6407) );
  AND2_X1 U5712 ( .A1(n4883), .A2(n8336), .ZN(n7799) );
  NAND2_X1 U5713 ( .A1(n4954), .A2(n8476), .ZN(n4953) );
  OR2_X1 U5714 ( .A1(n6321), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U5715 ( .A1(n6580), .A2(n6579), .ZN(n7592) );
  NAND2_X1 U5716 ( .A1(n8794), .A2(n6279), .ZN(n8294) );
  AND2_X1 U5717 ( .A1(n6618), .A2(n6780), .ZN(n7804) );
  INV_X1 U5718 ( .A(SI_10_), .ZN(n10097) );
  NAND2_X1 U5719 ( .A1(n6795), .A2(n6794), .ZN(n7366) );
  AND2_X1 U5720 ( .A1(n6560), .A2(n6559), .ZN(n8636) );
  AND2_X1 U5721 ( .A1(n8415), .A2(n8416), .ZN(n8669) );
  NAND2_X1 U5722 ( .A1(n8742), .A2(n6602), .ZN(n8729) );
  AND2_X1 U5723 ( .A1(n8395), .A2(n8393), .ZN(n8736) );
  OR2_X1 U5724 ( .A1(n8751), .A2(n8750), .ZN(n8753) );
  AND2_X1 U5725 ( .A1(n6333), .A2(n6332), .ZN(n10019) );
  NAND2_X1 U5726 ( .A1(n8446), .A2(n6633), .ZN(n6769) );
  OR2_X1 U5727 ( .A1(n8435), .A2(n6680), .ZN(n6780) );
  AND2_X1 U5728 ( .A1(n6775), .A2(n6857), .ZN(n6781) );
  AND2_X1 U5729 ( .A1(n6765), .A2(n6857), .ZN(n6762) );
  NAND2_X1 U5730 ( .A1(n7775), .A2(n7866), .ZN(n10029) );
  INV_X1 U5731 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n6238) );
  NOR2_X1 U5732 ( .A1(n4963), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4961) );
  INV_X1 U5733 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6236) );
  INV_X1 U5734 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5108) );
  XNOR2_X1 U5735 ( .A(n6393), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8490) );
  INV_X1 U5736 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U5737 ( .A1(n9130), .A2(n4867), .ZN(n4866) );
  NAND2_X1 U5738 ( .A1(n5993), .A2(n7673), .ZN(n5977) );
  OR2_X1 U5739 ( .A1(n5370), .A2(n9087), .ZN(n5359) );
  NAND2_X1 U5740 ( .A1(n6101), .A2(n4829), .ZN(n4828) );
  NAND2_X1 U5741 ( .A1(n4830), .A2(n4832), .ZN(n4829) );
  NAND2_X1 U5742 ( .A1(n7727), .A2(n4856), .ZN(n4851) );
  INV_X1 U5743 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9114) );
  NAND2_X1 U5744 ( .A1(n5280), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5405) );
  NOR2_X1 U5745 ( .A1(n9636), .A2(n9637), .ZN(n9635) );
  INV_X1 U5746 ( .A(n6014), .ZN(n6013) );
  NAND2_X1 U5747 ( .A1(n5882), .A2(n8097), .ZN(n4747) );
  NAND2_X1 U5748 ( .A1(n5883), .A2(n7778), .ZN(n5958) );
  NAND2_X1 U5749 ( .A1(n5924), .A2(n5957), .ZN(n5925) );
  INV_X1 U5750 ( .A(n5929), .ZN(n5926) );
  AND3_X1 U5751 ( .A1(n5734), .A2(n5733), .A3(n5732), .ZN(n9347) );
  OR2_X1 U5753 ( .A1(n6906), .A2(n6905), .ZN(n4706) );
  NOR2_X1 U5754 ( .A1(n6967), .A2(n4702), .ZN(n9266) );
  AND2_X1 U5755 ( .A1(n6968), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n4702) );
  AOI21_X1 U5756 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6968), .A(n6961), .ZN(
        n9261) );
  NAND2_X1 U5757 ( .A1(n9266), .A2(n9267), .ZN(n9265) );
  AOI21_X1 U5758 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7308), .A(n7303), .ZN(
        n7304) );
  NOR2_X1 U5759 ( .A1(n4696), .A2(n7307), .ZN(n7310) );
  AND2_X1 U5760 ( .A1(n7308), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4696) );
  NAND2_X1 U5761 ( .A1(n7310), .A2(n7309), .ZN(n7422) );
  AOI21_X1 U5762 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n7855), .A(n7850), .ZN(
        n9284) );
  NOR2_X1 U5763 ( .A1(n7854), .A2(n4704), .ZN(n9274) );
  AND2_X1 U5764 ( .A1(n7855), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4704) );
  AND2_X1 U5765 ( .A1(n9298), .A2(n9297), .ZN(n9299) );
  AND2_X1 U5766 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5420) );
  INV_X1 U5767 ( .A(n4782), .ZN(n4778) );
  AND2_X1 U5768 ( .A1(n4780), .A2(n4776), .ZN(n4775) );
  NAND2_X1 U5769 ( .A1(n4773), .A2(n4772), .ZN(n4771) );
  OR2_X1 U5770 ( .A1(n8070), .A2(n4780), .ZN(n4772) );
  NAND2_X1 U5771 ( .A1(n4774), .A2(n4780), .ZN(n4773) );
  NAND2_X1 U5772 ( .A1(n4776), .A2(n4782), .ZN(n4774) );
  OAI21_X1 U5773 ( .B1(n9387), .B2(n5067), .A(n5065), .ZN(n9359) );
  INV_X1 U5774 ( .A(n5066), .ZN(n5065) );
  INV_X1 U5775 ( .A(n8064), .ZN(n5072) );
  AND2_X1 U5776 ( .A1(n5800), .A2(n8033), .ZN(n9394) );
  INV_X1 U5777 ( .A(n4801), .ZN(n9407) );
  NAND2_X1 U5778 ( .A1(n4795), .A2(n4791), .ZN(n4790) );
  NAND2_X1 U5779 ( .A1(n9444), .A2(n4755), .ZN(n9402) );
  NAND2_X1 U5780 ( .A1(n9444), .A2(n9435), .ZN(n9429) );
  AND2_X1 U5781 ( .A1(n5837), .A2(n5838), .ZN(n9488) );
  INV_X1 U5782 ( .A(n5472), .ZN(n5278) );
  AND2_X1 U5783 ( .A1(n9489), .A2(n5832), .ZN(n9505) );
  INV_X1 U5784 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5470) );
  OR2_X1 U5785 ( .A1(n5504), .A2(n5470), .ZN(n5472) );
  NAND2_X1 U5786 ( .A1(n5276), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U5787 ( .A1(n9592), .A2(n7954), .ZN(n9593) );
  NAND2_X1 U5788 ( .A1(n7834), .A2(n4764), .ZN(n9601) );
  NAND2_X1 U5789 ( .A1(n7819), .A2(n4561), .ZN(n4806) );
  INV_X1 U5790 ( .A(n7874), .ZN(n4808) );
  INV_X1 U5791 ( .A(n5819), .ZN(n9597) );
  INV_X1 U5792 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10363) );
  OR2_X1 U5793 ( .A1(n5533), .A2(n10363), .ZN(n5519) );
  INV_X1 U5794 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5531) );
  OR2_X1 U5795 ( .A1(n5546), .A2(n5531), .ZN(n5533) );
  NAND2_X1 U5796 ( .A1(n5275), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5546) );
  INV_X1 U5797 ( .A(n5560), .ZN(n5275) );
  NAND2_X1 U5798 ( .A1(n5676), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5668) );
  OR2_X1 U5799 ( .A1(n5668), .A2(n5558), .ZN(n5560) );
  NAND2_X1 U5800 ( .A1(n5900), .A2(n7779), .ZN(n7829) );
  NAND2_X1 U5801 ( .A1(n4760), .A2(n4759), .ZN(n9756) );
  AND2_X1 U5802 ( .A1(n5698), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5676) );
  INV_X1 U5803 ( .A(n5042), .ZN(n5041) );
  OAI21_X1 U5804 ( .B1(n7533), .B2(n5043), .A(n7716), .ZN(n5042) );
  NAND2_X1 U5805 ( .A1(n9763), .A2(n9761), .ZN(n7534) );
  INV_X1 U5806 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5589) );
  NOR2_X1 U5807 ( .A1(n5653), .A2(n5589), .ZN(n5696) );
  AND2_X1 U5808 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5654) );
  XNOR2_X1 U5809 ( .A(n9197), .B(n9844), .ZN(n7518) );
  NAND2_X1 U5810 ( .A1(n7472), .A2(n7471), .ZN(n9600) );
  NAND2_X1 U5811 ( .A1(n5274), .A2(n5273), .ZN(n9532) );
  OR2_X1 U5812 ( .A1(n9631), .A2(n5633), .ZN(n5274) );
  INV_X1 U5813 ( .A(n9600), .ZN(n9793) );
  NAND2_X1 U5814 ( .A1(n5368), .A2(n5367), .ZN(n9563) );
  OAI22_X1 U5815 ( .A1(n9592), .A2(n4663), .B1(n4664), .B2(n8042), .ZN(n9656)
         );
  INV_X1 U5816 ( .A(n9898), .ZN(n9913) );
  AND2_X1 U5817 ( .A1(n6929), .A2(n7472), .ZN(n9898) );
  AND2_X1 U5818 ( .A1(n9831), .A2(n6927), .ZN(n9527) );
  XNOR2_X1 U5819 ( .A(n5722), .B(n5720), .ZN(n5253) );
  NAND2_X1 U5820 ( .A1(n5941), .A2(n5268), .ZN(n5272) );
  INV_X1 U5821 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5415) );
  INV_X1 U5822 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5414) );
  NAND2_X1 U5823 ( .A1(n5030), .A2(n5032), .ZN(n5525) );
  OR2_X1 U5824 ( .A1(n5169), .A2(n5034), .ZN(n5030) );
  INV_X1 U5825 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5057) );
  INV_X1 U5826 ( .A(n5084), .ZN(n5083) );
  OAI21_X1 U5827 ( .B1(n5087), .B2(n5092), .A(n8217), .ZN(n5084) );
  INV_X1 U5828 ( .A(n8685), .ZN(n8174) );
  INV_X1 U5829 ( .A(n5107), .ZN(n5106) );
  NAND2_X1 U5830 ( .A1(n6488), .A2(n6487), .ZN(n8708) );
  INV_X1 U5831 ( .A(n8471), .ZN(n8116) );
  NAND2_X1 U5832 ( .A1(n5094), .A2(n5098), .ZN(n8141) );
  NAND2_X1 U5833 ( .A1(n8201), .A2(n5100), .ZN(n5094) );
  NAND2_X1 U5834 ( .A1(n8233), .A2(n6727), .ZN(n8150) );
  NAND2_X1 U5835 ( .A1(n7377), .A2(n6699), .ZN(n7411) );
  NAND2_X1 U5836 ( .A1(n7248), .A2(n6694), .ZN(n7379) );
  AND4_X1 U5837 ( .A1(n6478), .A2(n6477), .A3(n6476), .A4(n6475), .ZN(n8747)
         );
  NAND2_X1 U5838 ( .A1(n8013), .A2(n6719), .ZN(n8192) );
  OR2_X1 U5839 ( .A1(n6784), .A2(n6782), .ZN(n8223) );
  NAND2_X1 U5840 ( .A1(n8161), .A2(n6732), .ZN(n8209) );
  NAND2_X1 U5841 ( .A1(n6461), .A2(n6460), .ZN(n8854) );
  NAND2_X1 U5842 ( .A1(n6703), .A2(n6702), .ZN(n7503) );
  INV_X1 U5843 ( .A(n8238), .ZN(n8211) );
  OAI21_X1 U5844 ( .B1(n8201), .B2(n5091), .A(n5089), .ZN(n8221) );
  INV_X1 U5845 ( .A(n8232), .ZN(n8230) );
  AND4_X1 U5846 ( .A1(n6449), .A2(n6448), .A3(n6447), .A4(n6446), .ZN(n8239)
         );
  OR2_X1 U5847 ( .A1(n6982), .A2(n6779), .ZN(n8241) );
  NAND2_X1 U5848 ( .A1(n8869), .A2(n8457), .ZN(n4716) );
  INV_X1 U5849 ( .A(n8458), .ZN(n4717) );
  INV_X1 U5850 ( .A(n8224), .ZN(n8671) );
  NAND2_X1 U5851 ( .A1(n6511), .A2(n6510), .ZN(n8696) );
  INV_X1 U5852 ( .A(n6740), .ZN(n8717) );
  INV_X1 U5853 ( .A(n8747), .ZN(n8718) );
  INV_X1 U5854 ( .A(n8164), .ZN(n8767) );
  NAND2_X1 U5855 ( .A1(n6309), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6260) );
  OR2_X2 U5856 ( .A1(n6947), .A2(n6981), .ZN(n8573) );
  OR2_X1 U5857 ( .A1(n6295), .A2(n6242), .ZN(n6248) );
  NAND2_X1 U5858 ( .A1(n7085), .A2(n7086), .ZN(n7084) );
  NAND2_X1 U5859 ( .A1(n7127), .A2(n6997), .ZN(n7085) );
  NAND2_X1 U5860 ( .A1(n4912), .A2(n7151), .ZN(n7153) );
  INV_X1 U5861 ( .A(n4913), .ZN(n4912) );
  NOR2_X1 U5862 ( .A1(n7320), .A2(n7319), .ZN(n7324) );
  XNOR2_X1 U5863 ( .A(n7557), .B(n7558), .ZN(n7434) );
  AND2_X1 U5864 ( .A1(n6378), .A2(n6210), .ZN(n6402) );
  XNOR2_X1 U5865 ( .A(n4925), .B(n8532), .ZN(n8487) );
  NOR2_X1 U5866 ( .A1(n8487), .A2(n8505), .ZN(n8523) );
  OR2_X1 U5867 ( .A1(P2_U3150), .A2(n6948), .ZN(n8515) );
  OR2_X1 U5868 ( .A1(n10029), .A2(n7455), .ZN(n8676) );
  NAND2_X1 U5869 ( .A1(n8714), .A2(n6604), .ZN(n8702) );
  NAND2_X1 U5870 ( .A1(n4902), .A2(n4906), .ZN(n8721) );
  NAND2_X1 U5871 ( .A1(n8751), .A2(n8379), .ZN(n4902) );
  NAND2_X1 U5872 ( .A1(n6472), .A2(n6471), .ZN(n8850) );
  NAND2_X1 U5873 ( .A1(n4541), .A2(n4893), .ZN(n8006) );
  OR2_X1 U5874 ( .A1(n7988), .A2(n7984), .ZN(n4893) );
  NAND2_X1 U5875 ( .A1(n7663), .A2(n8332), .ZN(n7633) );
  NAND2_X1 U5876 ( .A1(n6585), .A2(n6584), .ZN(n7634) );
  NAND2_X1 U5877 ( .A1(n6763), .A2(n7775), .ZN(n8674) );
  AND2_X1 U5878 ( .A1(n7368), .A2(n8674), .ZN(n8771) );
  INV_X1 U5879 ( .A(n10029), .ZN(n10046) );
  INV_X2 U5880 ( .A(n8771), .ZN(n8812) );
  INV_X1 U5881 ( .A(n8674), .ZN(n8808) );
  AOI21_X1 U5882 ( .B1(n8248), .B2(n8250), .A(n8247), .ZN(n8876) );
  NAND2_X1 U5883 ( .A1(n4979), .A2(n4983), .ZN(n8623) );
  NAND2_X1 U5884 ( .A1(n6542), .A2(n6541), .ZN(n8884) );
  NAND2_X1 U5885 ( .A1(n6531), .A2(n6530), .ZN(n8890) );
  NAND2_X1 U5886 ( .A1(n4901), .A2(n8420), .ZN(n8644) );
  NAND2_X1 U5887 ( .A1(n6523), .A2(n6522), .ZN(n8896) );
  NAND2_X1 U5888 ( .A1(n6513), .A2(n6512), .ZN(n8902) );
  NAND2_X1 U5889 ( .A1(n6504), .A2(n6503), .ZN(n8908) );
  NAND2_X1 U5890 ( .A1(n6606), .A2(n6605), .ZN(n8683) );
  NAND2_X1 U5891 ( .A1(n6496), .A2(n6495), .ZN(n8914) );
  NAND2_X1 U5892 ( .A1(n6454), .A2(n6453), .ZN(n8937) );
  NAND2_X1 U5893 ( .A1(n6442), .A2(n6441), .ZN(n8944) );
  NAND2_X1 U5894 ( .A1(n6597), .A2(n6596), .ZN(n8783) );
  NAND2_X1 U5895 ( .A1(n4890), .A2(n4891), .ZN(n8777) );
  NAND2_X1 U5896 ( .A1(n7988), .A2(n4541), .ZN(n4890) );
  NAND2_X1 U5897 ( .A1(n6417), .A2(n6416), .ZN(n8118) );
  OAI21_X1 U5898 ( .B1(n6593), .B2(n4970), .A(n4967), .ZN(n7985) );
  NAND2_X1 U5899 ( .A1(n4898), .A2(n8354), .ZN(n7944) );
  NAND2_X1 U5900 ( .A1(n4972), .A2(n4973), .ZN(n7941) );
  NAND2_X1 U5901 ( .A1(n6593), .A2(n4975), .ZN(n4972) );
  NAND2_X1 U5902 ( .A1(n6593), .A2(n6592), .ZN(n7898) );
  NAND2_X1 U5903 ( .A1(n4883), .A2(n4519), .ZN(n7882) );
  NAND2_X1 U5904 ( .A1(n6653), .A2(n6857), .ZN(n6865) );
  INV_X1 U5905 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6639) );
  NAND2_X1 U5906 ( .A1(n6643), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6640) );
  INV_X1 U5907 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7868) );
  INV_X1 U5908 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7774) );
  INV_X1 U5909 ( .A(n6679), .ZN(n7775) );
  INV_X1 U5910 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7617) );
  INV_X1 U5911 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10233) );
  INV_X1 U5912 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10284) );
  INV_X1 U5913 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7149) );
  INV_X1 U5914 ( .A(n8537), .ZN(n9994) );
  INV_X1 U5915 ( .A(n8502), .ZN(n9971) );
  INV_X1 U5916 ( .A(n8490), .ZN(n8484) );
  INV_X1 U5917 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10343) );
  INV_X1 U5918 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6870) );
  INV_X1 U5919 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6851) );
  OR2_X1 U5920 ( .A1(n6262), .A2(n4918), .ZN(n4917) );
  NAND2_X1 U5921 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4918) );
  NAND2_X1 U5922 ( .A1(n5318), .A2(n5317), .ZN(n9543) );
  AOI22_X1 U5923 ( .A1(n4820), .A2(n4824), .B1(n4818), .B2(n4825), .ZN(n4815)
         );
  NAND2_X1 U5924 ( .A1(n5427), .A2(n5426), .ZN(n9582) );
  AND2_X1 U5925 ( .A1(n8978), .A2(n8977), .ZN(n9030) );
  NAND2_X1 U5926 ( .A1(n5306), .A2(n5305), .ZN(n9538) );
  NAND2_X1 U5927 ( .A1(n5401), .A2(n5400), .ZN(n9572) );
  OAI21_X1 U5928 ( .B1(n8996), .B2(n4832), .A(n4830), .ZN(n9062) );
  NAND2_X1 U5929 ( .A1(n4875), .A2(n4874), .ZN(n4873) );
  NAND2_X1 U5930 ( .A1(n6069), .A2(n4875), .ZN(n4872) );
  INV_X1 U5931 ( .A(n9637), .ZN(n4874) );
  NAND2_X1 U5932 ( .A1(n5544), .A2(n5543), .ZN(n9897) );
  OAI22_X1 U5933 ( .A1(n6818), .A2(n6814), .B1(n6265), .B2(n6812), .ZN(n4658)
         );
  NAND2_X1 U5934 ( .A1(n6191), .A2(n6190), .ZN(n9153) );
  AOI21_X1 U5935 ( .B1(n9071), .B2(n9072), .A(n4825), .ZN(n9151) );
  INV_X1 U5936 ( .A(n4835), .ZN(n4833) );
  NAND2_X1 U5937 ( .A1(n8996), .A2(n4544), .ZN(n4837) );
  INV_X1 U5938 ( .A(n9096), .ZN(n9693) );
  NAND2_X1 U5939 ( .A1(n5313), .A2(n5312), .ZN(n9173) );
  OR2_X2 U5940 ( .A1(n5960), .A2(n6809), .ZN(n9198) );
  NAND2_X1 U5941 ( .A1(n9205), .A2(n9204), .ZN(n9203) );
  AOI21_X1 U5942 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n9252), .A(n9253), .ZN(
        n6903) );
  AND2_X1 U5943 ( .A1(n9246), .A2(n4707), .ZN(n6906) );
  NAND2_X1 U5944 ( .A1(n9252), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4707) );
  INV_X1 U5945 ( .A(n4706), .ZN(n6904) );
  AOI21_X1 U5946 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6907), .A(n6901), .ZN(
        n6915) );
  AND2_X1 U5947 ( .A1(n4706), .A2(n4705), .ZN(n6918) );
  NAND2_X1 U5948 ( .A1(n6907), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n4705) );
  AOI21_X1 U5949 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6919), .A(n6913), .ZN(
        n6882) );
  NOR2_X1 U5950 ( .A1(n6916), .A2(n4703), .ZN(n6895) );
  NOR2_X1 U5951 ( .A1(n6876), .A2(n6891), .ZN(n4703) );
  NOR2_X1 U5952 ( .A1(n6895), .A2(n6894), .ZN(n6967) );
  AOI21_X1 U5953 ( .B1(n7139), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7138), .ZN(
        n7142) );
  NOR2_X1 U5954 ( .A1(n7136), .A2(n7137), .ZN(n7307) );
  NOR2_X1 U5955 ( .A1(n7134), .A2(n4695), .ZN(n7137) );
  AND2_X1 U5956 ( .A1(n7139), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4695) );
  AOI21_X1 U5957 ( .B1(n7623), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7622), .ZN(
        n7626) );
  NOR2_X1 U5958 ( .A1(n7618), .A2(n4613), .ZN(n7621) );
  XNOR2_X1 U5959 ( .A(n9274), .B(n9283), .ZN(n7856) );
  INV_X1 U5960 ( .A(n4767), .ZN(n9534) );
  NAND2_X1 U5961 ( .A1(n4779), .A2(n4784), .ZN(n9360) );
  XNOR2_X1 U5962 ( .A(n4680), .B(n9374), .ZN(n9545) );
  NAND2_X1 U5963 ( .A1(n5069), .A2(n4545), .ZN(n4680) );
  NAND2_X1 U5964 ( .A1(n5071), .A2(n4521), .ZN(n5069) );
  NAND2_X1 U5965 ( .A1(n5071), .A2(n8063), .ZN(n8079) );
  NAND2_X1 U5966 ( .A1(n4672), .A2(n5049), .ZN(n9401) );
  NAND2_X1 U5967 ( .A1(n4674), .A2(n4673), .ZN(n4672) );
  INV_X1 U5968 ( .A(n9563), .ZN(n9424) );
  NAND2_X1 U5969 ( .A1(n4798), .A2(n4799), .ZN(n9417) );
  NAND2_X1 U5970 ( .A1(n5053), .A2(n8058), .ZN(n5052) );
  INV_X1 U5971 ( .A(n9578), .ZN(n9470) );
  AND2_X1 U5972 ( .A1(n5046), .A2(n4600), .ZN(n9457) );
  NAND2_X1 U5973 ( .A1(n9487), .A2(n5838), .ZN(n9480) );
  NAND2_X1 U5974 ( .A1(n8050), .A2(n5112), .ZN(n9473) );
  NAND2_X1 U5975 ( .A1(n5455), .A2(n5454), .ZN(n9521) );
  NAND2_X1 U5976 ( .A1(n5469), .A2(n5468), .ZN(n9654) );
  NAND2_X1 U5977 ( .A1(n5482), .A2(n5481), .ZN(n9735) );
  NAND2_X1 U5978 ( .A1(n7819), .A2(n5818), .ZN(n7869) );
  NAND2_X1 U5979 ( .A1(n5060), .A2(n5061), .ZN(n7953) );
  NAND2_X1 U5980 ( .A1(n7831), .A2(n7830), .ZN(n7873) );
  NAND2_X1 U5981 ( .A1(n9773), .A2(n9772), .ZN(n5044) );
  NAND2_X1 U5982 ( .A1(n4625), .A2(n4730), .ZN(n9766) );
  OAI21_X1 U5983 ( .B1(n9779), .B2(n5897), .A(n5757), .ZN(n7685) );
  INV_X1 U5984 ( .A(n9757), .ZN(n9661) );
  INV_X1 U5985 ( .A(n9797), .ZN(n9662) );
  NAND2_X1 U5986 ( .A1(n9516), .A2(n7475), .ZN(n9500) );
  OR2_X1 U5987 ( .A1(n6926), .A2(n9833), .ZN(n9513) );
  INV_X1 U5988 ( .A(n9500), .ZN(n9788) );
  INV_X1 U5989 ( .A(n9936), .ZN(n9934) );
  AND2_X2 U5990 ( .A1(n9527), .A2(n7465), .ZN(n9919) );
  NOR2_X1 U5991 ( .A1(n9800), .A2(n9833), .ZN(n9830) );
  NAND2_X1 U5992 ( .A1(n9621), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5289) );
  AND2_X1 U5993 ( .A1(n5063), .A2(n4528), .ZN(n4753) );
  NAND2_X1 U5994 ( .A1(n5944), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5942) );
  OR2_X1 U5995 ( .A1(n5941), .A2(n5943), .ZN(n5945) );
  INV_X1 U5996 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7865) );
  INV_X1 U5997 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7776) );
  NAND2_X1 U5998 ( .A1(n5210), .A2(n5209), .ZN(n5391) );
  INV_X1 U5999 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8100) );
  INV_X1 U6000 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7180) );
  INV_X1 U6001 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10331) );
  NAND2_X1 U6002 ( .A1(n4990), .A2(n5149), .ZN(n5649) );
  INV_X1 U6003 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6826) );
  XNOR2_X1 U6004 ( .A(n4694), .B(n5612), .ZN(n6883) );
  NAND2_X1 U6005 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4694) );
  OAI21_X1 U6006 ( .B1(n6788), .B2(n8245), .A(n6787), .ZN(n6789) );
  NAND2_X1 U6007 ( .A1(n4527), .A2(n9991), .ZN(n4681) );
  AOI211_X1 U6008 ( .C1(n8602), .C2(n9991), .A(n8601), .B(n8600), .ZN(n8603)
         );
  NAND2_X1 U6009 ( .A1(n4928), .A2(n8592), .ZN(n4927) );
  OAI22_X1 U6010 ( .A1(n6804), .A2(n8867), .B1(n10466), .B2(n6803), .ZN(n6805)
         );
  AOI21_X1 U6011 ( .B1(n8616), .B2(n8943), .A(n6677), .ZN(n6678) );
  OAI211_X1 U6012 ( .C1(n6184), .C2(n6183), .A(n9096), .B(n8986), .ZN(n6202)
         );
  NAND2_X1 U6013 ( .A1(n4745), .A2(n5937), .ZN(n5955) );
  AOI21_X1 U6014 ( .B1(n4699), .B2(n5883), .A(n4698), .ZN(n4697) );
  NAND2_X1 U6015 ( .A1(n4804), .A2(n4614), .ZN(P1_U3519) );
  NAND2_X1 U6016 ( .A1(n9607), .A2(n9919), .ZN(n4804) );
  INV_X1 U6017 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n4803) );
  AND2_X1 U6018 ( .A1(n7801), .A2(n8336), .ZN(n4519) );
  OR2_X1 U6019 ( .A1(n4691), .A2(n4690), .ZN(n4520) );
  OAI211_X1 U6020 ( .C1(n6266), .C2(n7172), .A(n6304), .B(n6303), .ZN(n7596)
         );
  NAND2_X1 U6021 ( .A1(n9003), .A2(n9005), .ZN(n9004) );
  INV_X1 U6022 ( .A(n9533), .ZN(n4766) );
  NOR2_X1 U6023 ( .A1(n8066), .A2(n5070), .ZN(n4521) );
  AND2_X1 U6024 ( .A1(n8031), .A2(n5833), .ZN(n4522) );
  OR2_X1 U6025 ( .A1(n8884), .A2(n8647), .ZN(n4524) );
  AND2_X1 U6026 ( .A1(n8210), .A2(n5081), .ZN(n4525) );
  INV_X1 U6027 ( .A(n4947), .ZN(n4946) );
  OR2_X1 U6028 ( .A1(n6609), .A2(n4948), .ZN(n4947) );
  AND2_X1 U6029 ( .A1(n4692), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4526) );
  NAND2_X1 U6030 ( .A1(n5739), .A2(n5738), .ZN(n9357) );
  INV_X1 U6031 ( .A(n9357), .ZN(n4656) );
  NAND2_X1 U6032 ( .A1(n5357), .A2(n5356), .ZN(n9557) );
  XNOR2_X1 U6033 ( .A(n8585), .B(n8586), .ZN(n4527) );
  AND2_X1 U6034 ( .A1(n5287), .A2(n5286), .ZN(n4528) );
  OR2_X1 U6035 ( .A1(n4653), .A2(n4656), .ZN(n4529) );
  OR2_X1 U6036 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4530) );
  AND2_X1 U6037 ( .A1(n4790), .A2(n4573), .ZN(n4531) );
  AND2_X1 U6038 ( .A1(n9406), .A2(n8061), .ZN(n4532) );
  NAND2_X1 U6039 ( .A1(n8118), .A2(n8470), .ZN(n4533) );
  AND2_X1 U6040 ( .A1(n5109), .A2(n4565), .ZN(n4534) );
  NAND2_X1 U6041 ( .A1(n4800), .A2(n9436), .ZN(n4535) );
  AND2_X1 U6042 ( .A1(n5008), .A2(n5438), .ZN(n4536) );
  NAND2_X1 U6043 ( .A1(n5499), .A2(n5498), .ZN(n9168) );
  AND2_X1 U6044 ( .A1(n4755), .A2(n4754), .ZN(n4537) );
  NOR2_X1 U6045 ( .A1(n4762), .A2(n9168), .ZN(n4538) );
  AND2_X1 U6046 ( .A1(n4526), .A2(n4688), .ZN(n4539) );
  AND2_X1 U6047 ( .A1(n4618), .A2(n4520), .ZN(n4540) );
  NAND2_X1 U6048 ( .A1(n7727), .A2(n7729), .ZN(n7728) );
  NAND2_X1 U6049 ( .A1(n8013), .A2(n4605), .ZN(n8190) );
  INV_X1 U6050 ( .A(n6115), .ZN(n4826) );
  INV_X1 U6051 ( .A(n6280), .ZN(n6528) );
  XNOR2_X1 U6052 ( .A(n5979), .B(n5980), .ZN(n5038) );
  INV_X2 U6053 ( .A(n5983), .ZN(n5963) );
  AND2_X1 U6054 ( .A1(n4512), .A2(n8368), .ZN(n4541) );
  AND2_X1 U6055 ( .A1(n6276), .A2(n6278), .ZN(n4542) );
  XNOR2_X1 U6056 ( .A(n6615), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6679) );
  INV_X1 U6057 ( .A(n8038), .ZN(n4783) );
  AND2_X1 U6058 ( .A1(n6744), .A2(n8704), .ZN(n4543) );
  NAND2_X1 U6059 ( .A1(n6161), .A2(n5948), .ZN(n5960) );
  INV_X1 U6060 ( .A(n6256), .ZN(n6545) );
  OR2_X1 U6061 ( .A1(n8101), .A2(n8028), .ZN(n6256) );
  NAND2_X1 U6062 ( .A1(n5187), .A2(n5186), .ZN(n5493) );
  NAND2_X1 U6063 ( .A1(n6574), .A2(n6573), .ZN(n6571) );
  NAND2_X1 U6064 ( .A1(n6316), .A2(n6205), .ZN(n6328) );
  OR2_X1 U6065 ( .A1(n8994), .A2(n4838), .ZN(n4544) );
  OR2_X1 U6066 ( .A1(n9546), .A2(n9175), .ZN(n4545) );
  AND2_X1 U6067 ( .A1(n5015), .A2(n5012), .ZN(n4546) );
  INV_X1 U6068 ( .A(n7289), .ZN(n4692) );
  AND2_X1 U6069 ( .A1(n6275), .A2(n4916), .ZN(n4547) );
  INV_X1 U6070 ( .A(n5055), .ZN(n5597) );
  AND2_X1 U6071 ( .A1(n5819), .A2(n5905), .ZN(n4805) );
  OR2_X1 U6072 ( .A1(n9567), .A2(n9179), .ZN(n4548) );
  OR2_X1 U6073 ( .A1(n10039), .A2(n7934), .ZN(n8336) );
  AND2_X1 U6074 ( .A1(n8036), .A2(n8035), .ZN(n4549) );
  NAND2_X1 U6075 ( .A1(n5085), .A2(n5083), .ZN(n8103) );
  INV_X1 U6076 ( .A(n4970), .ZN(n4969) );
  NAND2_X1 U6077 ( .A1(n4973), .A2(n4971), .ZN(n4970) );
  NAND2_X1 U6078 ( .A1(n6679), .A2(n8463), .ZN(n8435) );
  AND2_X1 U6079 ( .A1(n7529), .A2(n9859), .ZN(n4550) );
  NAND2_X1 U6080 ( .A1(n5292), .A2(n5293), .ZN(n5743) );
  AND2_X1 U6081 ( .A1(n5850), .A2(n6185), .ZN(n4551) );
  XNOR2_X1 U6082 ( .A(n5931), .B(n5930), .ZN(n5956) );
  INV_X4 U6083 ( .A(n6295), .ZN(n8253) );
  INV_X1 U6084 ( .A(n9408), .ZN(n4802) );
  NAND2_X1 U6085 ( .A1(n5288), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5941) );
  INV_X1 U6086 ( .A(n5876), .ZN(n4653) );
  AND2_X1 U6087 ( .A1(n8884), .A2(n8647), .ZN(n4552) );
  AND4_X1 U6088 ( .A1(n6353), .A2(n6352), .A3(n6351), .A4(n6350), .ZN(n7920)
         );
  NAND2_X1 U6089 ( .A1(n5530), .A2(n5529), .ZN(n9051) );
  AND2_X1 U6090 ( .A1(n4730), .A2(n5758), .ZN(n4553) );
  AND3_X1 U6091 ( .A1(n5104), .A2(n6203), .A3(n6301), .ZN(n4554) );
  AND2_X1 U6092 ( .A1(n4798), .A2(n4795), .ZN(n4555) );
  NAND2_X1 U6093 ( .A1(n6262), .A2(n6203), .ZN(n6275) );
  NAND2_X1 U6094 ( .A1(n5884), .A2(n5064), .ZN(n5946) );
  INV_X1 U6095 ( .A(n9557), .ZN(n9406) );
  AND2_X1 U6096 ( .A1(n6706), .A2(n8325), .ZN(n4556) );
  OR2_X1 U6097 ( .A1(n4653), .A2(n9357), .ZN(n4557) );
  AND2_X1 U6098 ( .A1(n6700), .A2(n7505), .ZN(n4558) );
  NOR2_X1 U6099 ( .A1(n9946), .A2(n8486), .ZN(n4559) );
  NOR2_X1 U6100 ( .A1(n8523), .A2(n8524), .ZN(n4560) );
  NAND2_X1 U6101 ( .A1(n4866), .A2(n4864), .ZN(n9003) );
  AND2_X1 U6102 ( .A1(n4808), .A2(n5818), .ZN(n4561) );
  NAND2_X1 U6103 ( .A1(n5759), .A2(n7707), .ZN(n4562) );
  AND2_X1 U6104 ( .A1(n8425), .A2(n8424), .ZN(n4563) );
  OR2_X1 U6105 ( .A1(n7605), .A2(n10008), .ZN(n4564) );
  NAND2_X1 U6106 ( .A1(n9444), .A2(n4757), .ZN(n4758) );
  AND2_X1 U6107 ( .A1(n6213), .A2(n6212), .ZN(n4565) );
  AND2_X1 U6108 ( .A1(n6584), .A2(n8476), .ZN(n4566) );
  NAND2_X1 U6109 ( .A1(n9051), .A2(n9189), .ZN(n4567) );
  INV_X1 U6110 ( .A(n5849), .ZN(n4645) );
  INV_X1 U6111 ( .A(n7955), .ZN(n4666) );
  INV_X1 U6112 ( .A(n5101), .ZN(n5100) );
  OR2_X1 U6113 ( .A1(n6749), .A2(n5102), .ZN(n5101) );
  INV_X1 U6114 ( .A(n4819), .ZN(n4818) );
  OAI21_X1 U6115 ( .B1(n9072), .B2(n4825), .A(n6115), .ZN(n4819) );
  NAND2_X1 U6116 ( .A1(n9532), .A2(n9898), .ZN(n4568) );
  AND2_X1 U6117 ( .A1(n4965), .A2(n6595), .ZN(n4569) );
  AND2_X1 U6118 ( .A1(n6728), .A2(n6727), .ZN(n4570) );
  AND2_X1 U6119 ( .A1(n7830), .A2(n4567), .ZN(n4571) );
  AND2_X1 U6120 ( .A1(n5157), .A2(SI_7_), .ZN(n4572) );
  AND2_X1 U6121 ( .A1(n8354), .A2(n8355), .ZN(n8352) );
  AND2_X1 U6122 ( .A1(n4802), .A2(n5851), .ZN(n4573) );
  INV_X1 U6123 ( .A(n8067), .ZN(n5074) );
  OR2_X1 U6124 ( .A1(n8944), .A2(n8239), .ZN(n8386) );
  INV_X1 U6125 ( .A(n8386), .ZN(n4886) );
  INV_X1 U6126 ( .A(n5838), .ZN(n4788) );
  NOR2_X1 U6127 ( .A1(n9424), .A2(n8060), .ZN(n4574) );
  NAND2_X1 U6128 ( .A1(n8451), .A2(n8252), .ZN(n8429) );
  INV_X1 U6129 ( .A(n8429), .ZN(n4722) );
  INV_X1 U6130 ( .A(n5092), .ZN(n5091) );
  NOR2_X1 U6131 ( .A1(n5097), .A2(n5093), .ZN(n5092) );
  INV_X1 U6132 ( .A(n4634), .ZN(n4633) );
  NOR2_X1 U6133 ( .A1(n4636), .A2(n5814), .ZN(n4634) );
  NAND2_X1 U6134 ( .A1(n5904), .A2(n5813), .ZN(n4575) );
  NOR2_X1 U6135 ( .A1(n8902), .A2(n8685), .ZN(n4576) );
  INV_X1 U6136 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5258) );
  INV_X1 U6137 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5513) );
  AND2_X1 U6138 ( .A1(n8879), .A2(n8468), .ZN(n4577) );
  INV_X1 U6139 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6205) );
  INV_X1 U6140 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6251) );
  AND4_X1 U6141 ( .A1(n6300), .A2(n6299), .A3(n6298), .A4(n6297), .ZN(n7605)
         );
  INV_X1 U6142 ( .A(n7605), .ZN(n8480) );
  INV_X1 U6143 ( .A(n4796), .ZN(n4795) );
  NAND2_X1 U6144 ( .A1(n4799), .A2(n4797), .ZN(n4796) );
  AND2_X1 U6145 ( .A1(n6096), .A2(n9160), .ZN(n4578) );
  AND2_X1 U6146 ( .A1(n5179), .A2(SI_12_), .ZN(n4579) );
  AND2_X1 U6147 ( .A1(n5151), .A2(SI_5_), .ZN(n4580) );
  INV_X1 U6148 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6828) );
  INV_X1 U6149 ( .A(n4675), .ZN(n4673) );
  NAND2_X1 U6150 ( .A1(n5051), .A2(n4676), .ZN(n4675) );
  INV_X1 U6151 ( .A(n9375), .ZN(n9374) );
  NAND2_X1 U6152 ( .A1(n5870), .A2(n8036), .ZN(n9375) );
  NAND2_X1 U6153 ( .A1(n9524), .A2(n9347), .ZN(n4581) );
  INV_X1 U6154 ( .A(n9524), .ZN(n5877) );
  NAND2_X1 U6155 ( .A1(n5730), .A2(n5729), .ZN(n9524) );
  INV_X1 U6156 ( .A(n4985), .ZN(n4984) );
  NAND2_X1 U6157 ( .A1(n4524), .A2(n5122), .ZN(n4985) );
  OR2_X1 U6158 ( .A1(n4552), .A2(n5121), .ZN(n4582) );
  NAND2_X1 U6159 ( .A1(n5819), .A2(n5906), .ZN(n4583) );
  INV_X1 U6160 ( .A(n5905), .ZN(n4807) );
  INV_X1 U6161 ( .A(n6113), .ZN(n4825) );
  NAND2_X1 U6162 ( .A1(n6112), .A2(n6111), .ZN(n6113) );
  AND2_X1 U6163 ( .A1(n8059), .A2(n4548), .ZN(n5051) );
  OR2_X1 U6164 ( .A1(n7823), .A2(n7822), .ZN(n7827) );
  AND2_X1 U6165 ( .A1(n4967), .A2(n4533), .ZN(n4584) );
  NAND2_X1 U6166 ( .A1(n8057), .A2(n9567), .ZN(n4585) );
  AND2_X1 U6167 ( .A1(n5052), .A2(n4548), .ZN(n4586) );
  OR2_X1 U6168 ( .A1(n4728), .A2(n5292), .ZN(n4587) );
  AND2_X1 U6169 ( .A1(n4871), .A2(n4870), .ZN(n4588) );
  NOR2_X1 U6170 ( .A1(n8260), .A2(n8431), .ZN(n4589) );
  AND2_X1 U6171 ( .A1(n6598), .A2(n6596), .ZN(n4590) );
  NOR2_X1 U6172 ( .A1(n8062), .A2(n4671), .ZN(n4670) );
  AND2_X1 U6173 ( .A1(n9535), .A2(n4568), .ZN(n4591) );
  INV_X1 U6174 ( .A(n4762), .ZN(n4761) );
  NAND2_X1 U6175 ( .A1(n4764), .A2(n4763), .ZN(n4762) );
  AND2_X1 U6176 ( .A1(n4534), .A2(n5108), .ZN(n4592) );
  OR2_X1 U6177 ( .A1(n4954), .A2(n4566), .ZN(n4593) );
  AND2_X1 U6178 ( .A1(n4753), .A2(n5884), .ZN(n4594) );
  INV_X1 U6179 ( .A(n7065), .ZN(n4688) );
  OR2_X1 U6180 ( .A1(n6330), .A2(n6329), .ZN(n7061) );
  INV_X1 U6181 ( .A(n7061), .ZN(n4691) );
  INV_X1 U6182 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4964) );
  NAND2_X1 U6183 ( .A1(n5344), .A2(n5343), .ZN(n9552) );
  INV_X1 U6184 ( .A(n9552), .ZN(n4754) );
  AND2_X1 U6185 ( .A1(n7834), .A2(n4761), .ZN(n4595) );
  NAND2_X1 U6186 ( .A1(n5055), .A2(n4523), .ZN(n5541) );
  NAND2_X1 U6187 ( .A1(n5364), .A2(n5363), .ZN(n9177) );
  NAND2_X1 U6188 ( .A1(n4837), .A2(n4833), .ZN(n9159) );
  NAND2_X1 U6189 ( .A1(n9593), .A2(n7955), .ZN(n8044) );
  XOR2_X1 U6190 ( .A(n6133), .B(n4514), .Z(n4596) );
  AND2_X1 U6191 ( .A1(n9582), .A2(n9182), .ZN(n4597) );
  AND2_X1 U6192 ( .A1(n8358), .A2(n8471), .ZN(n4598) );
  AND2_X1 U6193 ( .A1(n5813), .A2(n7779), .ZN(n4599) );
  NAND2_X1 U6194 ( .A1(n9478), .A2(n8051), .ZN(n4600) );
  INV_X1 U6195 ( .A(n6043), .ZN(n6076) );
  AND2_X1 U6196 ( .A1(n9448), .A2(n8056), .ZN(n4601) );
  NAND2_X1 U6197 ( .A1(n5055), .A2(n5056), .ZN(n5553) );
  NAND2_X1 U6198 ( .A1(n5512), .A2(n5513), .ZN(n5480) );
  AND2_X1 U6199 ( .A1(n6733), .A2(n8164), .ZN(n4602) );
  NAND2_X1 U6200 ( .A1(n4806), .A2(n5905), .ZN(n4603) );
  INV_X1 U6201 ( .A(n5902), .ZN(n4636) );
  AND2_X1 U6202 ( .A1(n4893), .A2(n8368), .ZN(n4604) );
  AND2_X1 U6203 ( .A1(n6720), .A2(n6719), .ZN(n4605) );
  NOR2_X1 U6204 ( .A1(n8708), .A2(n8717), .ZN(n4606) );
  NOR2_X1 U6205 ( .A1(n9635), .A2(n6069), .ZN(n4607) );
  OR2_X1 U6206 ( .A1(n5852), .A2(n6185), .ZN(n4608) );
  NAND2_X1 U6207 ( .A1(n5421), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n4609) );
  AND2_X1 U6208 ( .A1(n5212), .A2(SI_21_), .ZN(n4610) );
  NAND2_X1 U6209 ( .A1(n5209), .A2(SI_20_), .ZN(n4611) );
  NAND2_X1 U6210 ( .A1(n6378), .A2(n4534), .ZN(n4612) );
  XNOR2_X1 U6211 ( .A(n5942), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U6212 ( .A1(n7601), .A2(n8268), .ZN(n7491) );
  NOR2_X1 U6213 ( .A1(n9774), .A2(n7539), .ZN(n4760) );
  AND2_X1 U6214 ( .A1(n7623), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4613) );
  NAND2_X1 U6215 ( .A1(n5044), .A2(n7533), .ZN(n7714) );
  INV_X1 U6216 ( .A(n7558), .ZN(n7564) );
  AND2_X1 U6217 ( .A1(n6382), .A2(n6392), .ZN(n7558) );
  INV_X1 U6218 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n4690) );
  NAND2_X1 U6219 ( .A1(n6651), .A2(n6650), .ZN(n6653) );
  NAND2_X1 U6220 ( .A1(n4851), .A2(n6053), .ZN(n9095) );
  OR2_X1 U6221 ( .A1(n9919), .A2(n4803), .ZN(n4614) );
  INV_X1 U6222 ( .A(SI_20_), .ZN(n10270) );
  AND2_X1 U6223 ( .A1(n7503), .A2(n6705), .ZN(n4615) );
  NOR2_X2 U6224 ( .A1(n8097), .A2(n6931), .ZN(n6185) );
  INV_X1 U6225 ( .A(n9755), .ZN(n4759) );
  AND3_X2 U6226 ( .A1(n7366), .A2(n7365), .A3(n6801), .ZN(n10466) );
  INV_X1 U6227 ( .A(n10466), .ZN(n10463) );
  AND2_X1 U6228 ( .A1(n4935), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4616) );
  NAND2_X1 U6229 ( .A1(n6395), .A2(n6394), .ZN(n8012) );
  INV_X1 U6230 ( .A(n8012), .ZN(n4974) );
  AND2_X1 U6231 ( .A1(n8447), .A2(n6632), .ZN(n8782) );
  INV_X1 U6232 ( .A(n8782), .ZN(n8805) );
  AND2_X1 U6233 ( .A1(n4616), .A2(n8592), .ZN(n4617) );
  NAND2_X1 U6234 ( .A1(n6691), .A2(n6690), .ZN(n7246) );
  INV_X1 U6235 ( .A(n8799), .ZN(n6293) );
  OR2_X1 U6236 ( .A1(n7288), .A2(n7289), .ZN(n4618) );
  XNOR2_X1 U6237 ( .A(n6218), .B(n6217), .ZN(n8599) );
  AND2_X1 U6238 ( .A1(n4914), .A2(n7151), .ZN(n4619) );
  AND2_X1 U6239 ( .A1(n5958), .A2(n5957), .ZN(n4620) );
  AND2_X1 U6240 ( .A1(n8583), .A2(n4931), .ZN(n4621) );
  NAND2_X1 U6241 ( .A1(n4701), .A2(n4700), .ZN(n4699) );
  OAI21_X1 U6242 ( .B1(n9342), .B2(n5883), .A(n4697), .ZN(P1_U3262) );
  NAND2_X1 U6243 ( .A1(n4962), .A2(n4961), .ZN(n6240) );
  NAND2_X1 U6244 ( .A1(n7608), .A2(n7607), .ZN(n7606) );
  OAI21_X2 U6245 ( .B1(n8693), .B2(n6502), .A(n8406), .ZN(n8682) );
  NAND2_X2 U6246 ( .A1(n8759), .A2(n8376), .ZN(n8751) );
  OAI21_X1 U6247 ( .B1(n8448), .B2(n8447), .A(n4720), .ZN(n4719) );
  OAI21_X1 U6248 ( .B1(n4718), .B2(n4717), .A(n4716), .ZN(n4715) );
  AOI21_X2 U6249 ( .B1(n8751), .B2(n4905), .A(n4903), .ZN(n8707) );
  NAND3_X1 U6250 ( .A1(n5130), .A2(n7406), .A3(n5131), .ZN(n4679) );
  NAND2_X1 U6251 ( .A1(n8654), .A2(n8421), .ZN(n4901) );
  INV_X1 U6252 ( .A(n4889), .ZN(n4888) );
  OAI21_X1 U6253 ( .B1(n8251), .B2(n4896), .A(n4589), .ZN(n4895) );
  NOR2_X1 U6254 ( .A1(n8444), .A2(n4719), .ZN(n4718) );
  XNOR2_X1 U6255 ( .A(n4715), .B(n8599), .ZN(n8466) );
  NAND2_X1 U6256 ( .A1(n7219), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7327) );
  NAND2_X1 U6257 ( .A1(n7035), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7202) );
  INV_X1 U6258 ( .A(n4626), .ZN(n5827) );
  AOI21_X1 U6259 ( .B1(n5812), .B2(n4629), .A(n4627), .ZN(n4626) );
  NAND2_X1 U6260 ( .A1(n4638), .A2(n4637), .ZN(n4644) );
  AOI21_X1 U6261 ( .B1(n4639), .B2(n4640), .A(n4551), .ZN(n4637) );
  NAND2_X1 U6262 ( .A1(n5844), .A2(n4639), .ZN(n4638) );
  NAND2_X1 U6263 ( .A1(n4643), .A2(n4608), .ZN(n5853) );
  NAND2_X1 U6264 ( .A1(n4644), .A2(n5851), .ZN(n4643) );
  NAND2_X1 U6265 ( .A1(n6845), .A2(n4658), .ZN(n4657) );
  NAND2_X1 U6266 ( .A1(n9655), .A2(n4667), .ZN(n4660) );
  INV_X1 U6267 ( .A(n8042), .ZN(n4667) );
  INV_X1 U6268 ( .A(n8055), .ZN(n4674) );
  NAND2_X1 U6269 ( .A1(n8055), .A2(n4670), .ZN(n4668) );
  NOR2_X1 U6270 ( .A1(n8055), .A2(n4601), .ZN(n9428) );
  INV_X1 U6271 ( .A(n4601), .ZN(n4676) );
  AND2_X4 U6272 ( .A1(n4679), .A2(n4678), .ZN(n6814) );
  NOR2_X4 U6273 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6262) );
  NAND3_X1 U6274 ( .A1(n8581), .A2(n8580), .A3(n4681), .ZN(P2_U3200) );
  NAND2_X1 U6275 ( .A1(n7271), .A2(n4526), .ZN(n4689) );
  NAND2_X1 U6276 ( .A1(n7271), .A2(n4539), .ZN(n4686) );
  NAND2_X1 U6277 ( .A1(n4689), .A2(n4618), .ZN(n7291) );
  MUX2_X1 U6278 ( .A(n9920), .B(P1_REG1_REG_1__SCAN_IN), .S(n6883), .Z(n9205)
         );
  INV_X1 U6279 ( .A(n6573), .ZN(n7265) );
  NAND3_X1 U6280 ( .A1(n8319), .A2(n8435), .A3(n8318), .ZN(n4712) );
  AND2_X1 U6281 ( .A1(n6234), .A2(n6235), .ZN(n4713) );
  NAND2_X1 U6282 ( .A1(n4714), .A2(n6234), .ZN(n6646) );
  NAND2_X1 U6283 ( .A1(n4714), .A2(n4713), .ZN(n6648) );
  NAND3_X1 U6284 ( .A1(n8423), .A2(n8643), .A3(n8422), .ZN(n4723) );
  OAI211_X1 U6285 ( .C1(n8294), .C2(n4725), .A(n8302), .B(n4724), .ZN(n8313)
         );
  AND2_X1 U6286 ( .A1(n5566), .A2(n4587), .ZN(n4729) );
  OR2_X2 U6287 ( .A1(n5292), .A2(n5294), .ZN(n5637) );
  INV_X1 U6288 ( .A(n5294), .ZN(n5293) );
  INV_X1 U6289 ( .A(n5292), .ZN(n5295) );
  NAND3_X1 U6290 ( .A1(n4729), .A2(n5568), .A3(n5567), .ZN(n5974) );
  NAND2_X1 U6291 ( .A1(n5756), .A2(n5895), .ZN(n4732) );
  NAND2_X1 U6292 ( .A1(n4733), .A2(n4734), .ZN(n5825) );
  NAND2_X1 U6293 ( .A1(n5817), .A2(n4735), .ZN(n4733) );
  NAND4_X1 U6294 ( .A1(n5063), .A2(n4523), .A3(n4752), .A4(n4765), .ZN(n9621)
         );
  AND3_X2 U6295 ( .A1(n4765), .A2(n5259), .A3(n4523), .ZN(n5884) );
  NOR2_X2 U6296 ( .A1(n9495), .A2(n9582), .ZN(n9474) );
  AND2_X2 U6297 ( .A1(n9444), .A2(n4537), .ZN(n9388) );
  INV_X1 U6298 ( .A(n4758), .ZN(n9420) );
  NOR2_X2 U6299 ( .A1(n9756), .A2(n9883), .ZN(n7756) );
  NAND3_X1 U6300 ( .A1(n4591), .A2(n4767), .A3(n4766), .ZN(n9607) );
  NAND2_X1 U6301 ( .A1(n8086), .A2(n4775), .ZN(n4770) );
  OAI211_X1 U6302 ( .C1(n8086), .C2(n4777), .A(n4770), .B(n4771), .ZN(n8039)
         );
  NAND2_X1 U6303 ( .A1(n8086), .A2(n4549), .ZN(n4779) );
  NAND2_X1 U6304 ( .A1(n8086), .A2(n8035), .ZN(n9376) );
  AND2_X1 U6305 ( .A1(n9488), .A2(n9489), .ZN(n4789) );
  OAI21_X1 U6306 ( .B1(n9450), .B2(n9449), .A(n8032), .ZN(n9437) );
  NAND2_X1 U6307 ( .A1(n9449), .A2(n8032), .ZN(n4800) );
  NAND2_X1 U6308 ( .A1(n4806), .A2(n4805), .ZN(n9595) );
  INV_X1 U6309 ( .A(n5681), .ZN(n4809) );
  INV_X8 U6310 ( .A(n6814), .ZN(n6265) );
  NAND2_X1 U6311 ( .A1(n6814), .A2(n6822), .ZN(n4811) );
  NAND2_X2 U6312 ( .A1(n4812), .A2(n5960), .ZN(n5983) );
  NAND3_X1 U6313 ( .A1(n5958), .A2(n6932), .A3(n7674), .ZN(n4812) );
  NAND3_X1 U6314 ( .A1(n6928), .A2(n5958), .A3(n7471), .ZN(n4813) );
  NAND2_X1 U6315 ( .A1(n9071), .A2(n4816), .ZN(n4814) );
  NAND2_X1 U6316 ( .A1(n4814), .A2(n4815), .ZN(n9013) );
  AOI21_X1 U6317 ( .B1(n8996), .B2(n4830), .A(n4828), .ZN(n4827) );
  INV_X1 U6318 ( .A(n4827), .ZN(n6106) );
  INV_X1 U6319 ( .A(n8993), .ZN(n4838) );
  NAND2_X1 U6320 ( .A1(n5999), .A2(n4839), .ZN(n4842) );
  NAND2_X1 U6321 ( .A1(n4840), .A2(n8971), .ZN(n4843) );
  NAND2_X1 U6322 ( .A1(n4841), .A2(n4847), .ZN(n4844) );
  XNOR2_X1 U6323 ( .A(n6006), .B(n6007), .ZN(n7356) );
  NAND3_X1 U6324 ( .A1(n4844), .A2(n4845), .A3(n4843), .ZN(n6006) );
  NAND3_X1 U6325 ( .A1(n4846), .A2(n5999), .A3(n4514), .ZN(n4845) );
  NAND2_X1 U6326 ( .A1(n9689), .A2(n6029), .ZN(n7727) );
  NAND2_X1 U6327 ( .A1(n4848), .A2(n4852), .ZN(n6064) );
  NAND2_X1 U6328 ( .A1(n9689), .A2(n4849), .ZN(n4848) );
  NAND2_X1 U6329 ( .A1(n9130), .A2(n4859), .ZN(n4858) );
  NAND2_X1 U6330 ( .A1(n4858), .A2(n4861), .ZN(n6147) );
  NAND2_X1 U6331 ( .A1(n5512), .A2(n4588), .ZN(n4869) );
  NOR2_X2 U6332 ( .A1(n5541), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U6333 ( .A1(n6015), .A2(n6014), .ZN(n4877) );
  INV_X1 U6334 ( .A(n6015), .ZN(n4876) );
  AND2_X1 U6335 ( .A1(n9692), .A2(n4877), .ZN(n7511) );
  XNOR2_X2 U6336 ( .A(n9996), .B(n4878), .ZN(n8798) );
  INV_X1 U6337 ( .A(n9996), .ZN(n4879) );
  NAND2_X1 U6338 ( .A1(n7738), .A2(n4519), .ZN(n4880) );
  NAND2_X1 U6339 ( .A1(n4880), .A2(n4881), .ZN(n6391) );
  AOI21_X1 U6340 ( .B1(n4519), .B2(n8272), .A(n4882), .ZN(n4881) );
  NAND2_X1 U6341 ( .A1(n4898), .A2(n4897), .ZN(n6414) );
  NAND2_X1 U6342 ( .A1(n4901), .A2(n4899), .ZN(n6539) );
  INV_X1 U6343 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5104) );
  NAND2_X1 U6344 ( .A1(n7663), .A2(n4908), .ZN(n6355) );
  INV_X1 U6345 ( .A(n4911), .ZN(n7194) );
  INV_X1 U6346 ( .A(n4909), .ZN(n7213) );
  NAND2_X1 U6347 ( .A1(n4911), .A2(n4910), .ZN(n4909) );
  OR2_X1 U6348 ( .A1(n7191), .A2(n7192), .ZN(n4911) );
  NAND2_X1 U6349 ( .A1(n4913), .A2(n7151), .ZN(n7036) );
  OAI21_X1 U6350 ( .B1(n9947), .B2(n4920), .A(n4919), .ZN(n9963) );
  INV_X1 U6351 ( .A(n8521), .ZN(n4925) );
  NAND2_X1 U6352 ( .A1(n8528), .A2(n4616), .ZN(n4932) );
  NAND2_X1 U6353 ( .A1(n4932), .A2(n4926), .ZN(n4929) );
  NAND3_X1 U6354 ( .A1(n4929), .A2(n4930), .A3(n4927), .ZN(n8604) );
  NAND2_X1 U6355 ( .A1(n4932), .A2(n4933), .ZN(n8584) );
  NAND2_X1 U6356 ( .A1(n8528), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8560) );
  NAND2_X1 U6357 ( .A1(n4936), .A2(n6678), .ZN(P2_U3456) );
  NOR2_X1 U6358 ( .A1(n8612), .A2(n4937), .ZN(n6802) );
  NAND2_X1 U6359 ( .A1(n6597), .A2(n4590), .ZN(n8780) );
  NAND2_X1 U6360 ( .A1(n8780), .A2(n8763), .ZN(n6599) );
  NAND2_X1 U6361 ( .A1(n6601), .A2(n8750), .ZN(n8742) );
  OAI21_X1 U6362 ( .B1(n6606), .B2(n4947), .A(n4944), .ZN(n8656) );
  NAND2_X1 U6363 ( .A1(n4943), .A2(n4942), .ZN(n6611) );
  NAND2_X1 U6364 ( .A1(n6606), .A2(n4944), .ZN(n4943) );
  NAND2_X1 U6365 ( .A1(n6585), .A2(n4593), .ZN(n4952) );
  NAND2_X1 U6366 ( .A1(n4952), .A2(n4953), .ZN(n7739) );
  NOR2_X1 U6367 ( .A1(n6646), .A2(n4963), .ZN(n6250) );
  INV_X1 U6368 ( .A(n6646), .ZN(n4962) );
  NAND2_X1 U6369 ( .A1(n6593), .A2(n4584), .ZN(n4966) );
  NAND3_X1 U6370 ( .A1(n4967), .A2(n4970), .A3(n4533), .ZN(n4965) );
  NAND2_X1 U6371 ( .A1(n6612), .A2(n4980), .ZN(n4977) );
  NAND2_X1 U6372 ( .A1(n4977), .A2(n4978), .ZN(n6613) );
  NAND2_X1 U6373 ( .A1(n6612), .A2(n4984), .ZN(n4979) );
  AOI21_X1 U6374 ( .B1(n6612), .B2(n5122), .A(n5121), .ZN(n8634) );
  NAND2_X1 U6375 ( .A1(n5584), .A2(n5585), .ZN(n4990) );
  NAND2_X1 U6376 ( .A1(n5584), .A2(n4987), .ZN(n4986) );
  NAND2_X1 U6377 ( .A1(n5210), .A2(n4999), .ZN(n4995) );
  NAND2_X1 U6378 ( .A1(n4995), .A2(n4996), .ZN(n5377) );
  NAND2_X1 U6379 ( .A1(n5493), .A2(n4536), .ZN(n5007) );
  OR2_X1 U6380 ( .A1(n5493), .A2(n5191), .ZN(n5014) );
  NAND3_X1 U6381 ( .A1(n5008), .A2(n5011), .A3(n5438), .ZN(n5006) );
  NAND2_X1 U6382 ( .A1(n5223), .A2(n5021), .ZN(n5020) );
  NAND2_X1 U6383 ( .A1(n5223), .A2(n5222), .ZN(n5355) );
  NAND2_X1 U6384 ( .A1(n5020), .A2(n5024), .ZN(n5234) );
  NAND2_X1 U6385 ( .A1(n5169), .A2(n5029), .ZN(n5028) );
  NAND2_X1 U6386 ( .A1(n5169), .A2(n5168), .ZN(n5552) );
  OAI22_X1 U6387 ( .A1(n7549), .A2(n5038), .B1(n5979), .B2(n9835), .ZN(n7519)
         );
  NAND2_X1 U6388 ( .A1(n7545), .A2(n5038), .ZN(n5752) );
  XNOR2_X1 U6389 ( .A(n7549), .B(n5038), .ZN(n9836) );
  XNOR2_X1 U6390 ( .A(n7545), .B(n5038), .ZN(n7548) );
  NAND2_X1 U6391 ( .A1(n9773), .A2(n5040), .ZN(n5039) );
  NAND2_X1 U6392 ( .A1(n5039), .A2(n5041), .ZN(n9753) );
  NAND2_X1 U6393 ( .A1(n5046), .A2(n5045), .ZN(n8054) );
  NAND2_X1 U6394 ( .A1(n8050), .A2(n5047), .ZN(n5046) );
  INV_X1 U6395 ( .A(n9428), .ZN(n5053) );
  INV_X1 U6396 ( .A(n9051), .ZN(n5062) );
  AND2_X1 U6397 ( .A1(n5884), .A2(n5885), .ZN(n5588) );
  NAND2_X1 U6398 ( .A1(n5068), .A2(n5072), .ZN(n5067) );
  AND2_X1 U6399 ( .A1(n6692), .A2(n6690), .ZN(n5075) );
  NAND2_X1 U6400 ( .A1(n6696), .A2(n6695), .ZN(n7377) );
  NAND2_X1 U6401 ( .A1(n6730), .A2(n4525), .ZN(n5079) );
  NAND2_X1 U6402 ( .A1(n5079), .A2(n5080), .ZN(n8126) );
  NAND2_X1 U6403 ( .A1(n8201), .A2(n5086), .ZN(n5085) );
  NAND3_X1 U6404 ( .A1(n5104), .A2(n6262), .A3(n6203), .ZN(n6287) );
  OAI21_X2 U6405 ( .B1(n6703), .B2(n5106), .A(n5105), .ZN(n7764) );
  NAND2_X1 U6406 ( .A1(n6378), .A2(n4592), .ZN(n6216) );
  NAND2_X1 U6407 ( .A1(n6316), .A2(n5111), .ZN(n6356) );
  AND2_X2 U6408 ( .A1(n6316), .A2(n5110), .ZN(n6368) );
  OAI21_X1 U6409 ( .B1(n8987), .B2(n9026), .A(n9096), .ZN(n8992) );
  NAND2_X1 U6410 ( .A1(n5253), .A2(SI_29_), .ZN(n5724) );
  NAND2_X1 U6411 ( .A1(n5366), .A2(n5365), .ZN(n5223) );
  CLKBUF_X2 U6412 ( .A(n5980), .Z(n9835) );
  NAND2_X2 U6413 ( .A1(n6625), .A2(n6626), .ZN(n6266) );
  NAND2_X1 U6414 ( .A1(n6638), .A2(n6637), .ZN(n6669) );
  INV_X1 U6415 ( .A(n6636), .ZN(n6638) );
  OR2_X1 U6416 ( .A1(n5634), .A2(n6813), .ZN(n5614) );
  OAI21_X2 U6417 ( .B1(n8632), .B2(n8633), .A(n8426), .ZN(n8621) );
  OR2_X1 U6418 ( .A1(n5637), .A2(n9199), .ZN(n5608) );
  OR2_X1 U6419 ( .A1(n9389), .A2(n5637), .ZN(n5352) );
  OR2_X1 U6420 ( .A1(n8082), .A2(n5637), .ZN(n5340) );
  INV_X1 U6421 ( .A(n7650), .ZN(n5754) );
  OR2_X1 U6422 ( .A1(n6214), .A2(n6224), .ZN(n6215) );
  OAI22_X1 U6423 ( .A1(n8103), .A2(n8104), .B1(n8624), .B2(n6752), .ZN(n6755)
         );
  AOI21_X2 U6424 ( .B1(n9119), .B2(n9120), .A(n5117), .ZN(n8996) );
  INV_X2 U6425 ( .A(n10049), .ZN(n10047) );
  NAND2_X2 U6426 ( .A1(n7466), .A2(n9513), .ZN(n9516) );
  INV_X1 U6427 ( .A(n9704), .ZN(n6200) );
  AND2_X1 U6428 ( .A1(n6122), .A2(n6121), .ZN(n5113) );
  AND3_X1 U6429 ( .A1(n5746), .A2(n5745), .A3(n5744), .ZN(n8041) );
  INV_X1 U6430 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5558) );
  OR2_X1 U6431 ( .A1(n9110), .A2(n9111), .ZN(n5114) );
  AND2_X1 U6432 ( .A1(n6714), .A2(n7740), .ZN(n5116) );
  AND2_X1 U6433 ( .A1(n6088), .A2(n6087), .ZN(n5117) );
  NAND2_X1 U6434 ( .A1(n5422), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5118) );
  AND2_X1 U6435 ( .A1(n5168), .A2(n5167), .ZN(n5119) );
  INV_X1 U6436 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5421) );
  AND2_X1 U6437 ( .A1(n6061), .A2(n6062), .ZN(n5120) );
  INV_X1 U6438 ( .A(n9567), .ZN(n9435) );
  AND2_X1 U6439 ( .A1(n8890), .A2(n8657), .ZN(n5121) );
  OR2_X1 U6440 ( .A1(n8890), .A2(n8657), .ZN(n5122) );
  INV_X1 U6441 ( .A(n9546), .ZN(n8085) );
  OR2_X1 U6442 ( .A1(n8930), .A2(n8929), .ZN(P2_U3446) );
  OR2_X1 U6443 ( .A1(n8852), .A2(n8851), .ZN(P2_U3478) );
  OR2_X1 U6444 ( .A1(n8741), .A2(n8740), .ZN(P2_U3214) );
  NAND2_X1 U6445 ( .A1(n5240), .A2(n5239), .ZN(n5315) );
  OR2_X1 U6446 ( .A1(n8358), .A2(n8116), .ZN(n5126) );
  OR2_X1 U6447 ( .A1(n5935), .A2(n7910), .ZN(n5127) );
  INV_X1 U6448 ( .A(n10003), .ZN(n6292) );
  OR2_X1 U6449 ( .A1(n6845), .A2(n6885), .ZN(n5128) );
  NAND2_X1 U6450 ( .A1(n5234), .A2(n5233), .ZN(n5329) );
  OR2_X1 U6451 ( .A1(n6845), .A2(n6883), .ZN(n5129) );
  NAND2_X1 U6452 ( .A1(n5915), .A2(n5838), .ZN(n5839) );
  AOI21_X1 U6453 ( .B1(n5841), .B2(n5840), .A(n5839), .ZN(n5842) );
  INV_X1 U6454 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6230) );
  INV_X1 U6455 ( .A(n8041), .ZN(n5878) );
  INV_X1 U6456 ( .A(n8784), .ZN(n6598) );
  INV_X1 U6457 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U6458 ( .A1(n7040), .A2(n7065), .ZN(n7041) );
  INV_X1 U6459 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6406) );
  OR2_X1 U6460 ( .A1(n6653), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6665) );
  NAND2_X1 U6461 ( .A1(n6572), .A2(n7265), .ZN(n8296) );
  OR2_X1 U6462 ( .A1(n6104), .A2(n6103), .ZN(n6105) );
  INV_X1 U6463 ( .A(n5403), .ZN(n5280) );
  INV_X1 U6464 ( .A(n5519), .ZN(n5276) );
  INV_X1 U6465 ( .A(SI_23_), .ZN(n10219) );
  INV_X1 U6466 ( .A(n5397), .ZN(n5212) );
  INV_X1 U6467 ( .A(SI_19_), .ZN(n10294) );
  INV_X1 U6468 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U6469 ( .A1(n6361), .A2(n6360), .ZN(n6372) );
  NAND2_X1 U6470 ( .A1(n7042), .A2(n7041), .ZN(n7044) );
  OR2_X1 U6471 ( .A1(n6372), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6385) );
  OR2_X1 U6472 ( .A1(n6653), .A2(n6664), .ZN(n6796) );
  AND2_X1 U6473 ( .A1(n6183), .A2(n6180), .ZN(n6181) );
  INV_X1 U6474 ( .A(n6843), .ZN(n6178) );
  OR2_X1 U6475 ( .A1(n5334), .A2(n5319), .ZN(n5321) );
  NAND2_X1 U6476 ( .A1(n5282), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6477 ( .A1(n5281), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5382) );
  INV_X1 U6478 ( .A(n9178), .ZN(n8060) );
  NAND2_X1 U6479 ( .A1(n5278), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5458) );
  AND2_X1 U6480 ( .A1(n5696), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5698) );
  NOR2_X1 U6481 ( .A1(n7534), .A2(n7713), .ZN(n7708) );
  OR2_X1 U6482 ( .A1(n5722), .A2(n5721), .ZN(n5723) );
  INV_X1 U6483 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5270) );
  OR2_X1 U6484 ( .A1(n6473), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6481) );
  NAND2_X1 U6485 ( .A1(n6489), .A2(n8135), .ZN(n6497) );
  NOR2_X1 U6486 ( .A1(n6514), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6524) );
  INV_X1 U6487 ( .A(n7974), .ZN(n6715) );
  INV_X1 U6488 ( .A(n7502), .ZN(n6702) );
  AOI21_X1 U6489 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n9971), .A(n9963), .ZN(
        n8521) );
  AND2_X1 U6490 ( .A1(n6955), .A2(n8959), .ZN(n7012) );
  AND2_X1 U6491 ( .A1(n6532), .A2(n8222), .ZN(n6543) );
  AND2_X1 U6492 ( .A1(n6444), .A2(n6443), .ZN(n6464) );
  OR2_X1 U6493 ( .A1(n6385), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6396) );
  OR2_X1 U6494 ( .A1(n8435), .A2(n6768), .ZN(n6798) );
  OR2_X1 U6495 ( .A1(n6793), .A2(n7362), .ZN(n6795) );
  INV_X1 U6496 ( .A(n8647), .ZN(n8624) );
  INV_X1 U6497 ( .A(n8745), .ZN(n8750) );
  INV_X1 U6498 ( .A(n8475), .ZN(n7934) );
  AND2_X1 U6499 ( .A1(n6148), .A2(n6146), .ZN(n9079) );
  INV_X1 U6500 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9152) );
  AND2_X1 U6501 ( .A1(n5321), .A2(n5320), .ZN(n9381) );
  OR2_X1 U6502 ( .A1(n5430), .A2(n9114), .ZN(n5403) );
  NAND2_X1 U6503 ( .A1(n9379), .A2(n9371), .ZN(n9364) );
  NAND2_X1 U6504 ( .A1(n9567), .A2(n9179), .ZN(n8058) );
  INV_X1 U6505 ( .A(n9588), .ZN(n9501) );
  NAND2_X1 U6506 ( .A1(n7780), .A2(n5766), .ZN(n7815) );
  INV_X1 U6507 ( .A(n9505), .ZN(n9511) );
  AND2_X1 U6508 ( .A1(n5245), .A2(n5244), .ZN(n5316) );
  INV_X1 U6509 ( .A(n8223), .ZN(n8236) );
  INV_X1 U6510 ( .A(n8245), .ZN(n8227) );
  INV_X1 U6511 ( .A(n8599), .ZN(n8459) );
  AND3_X1 U6512 ( .A1(n6493), .A2(n6492), .A3(n6491), .ZN(n6740) );
  AND4_X1 U6513 ( .A1(n6390), .A2(n6389), .A3(n6388), .A4(n6387), .ZN(n7802)
         );
  NOR2_X1 U6514 ( .A1(n7560), .A2(n7559), .ZN(n7562) );
  INV_X1 U6515 ( .A(n8560), .ZN(n8529) );
  AND2_X1 U6516 ( .A1(n7012), .A2(n8540), .ZN(n9991) );
  OR2_X1 U6517 ( .A1(n6543), .A2(n6533), .ZN(n8650) );
  INV_X1 U6518 ( .A(n8793), .ZN(n8727) );
  OR2_X1 U6519 ( .A1(n7804), .A2(n8796), .ZN(n7456) );
  INV_X1 U6520 ( .A(n8867), .ZN(n8859) );
  AND2_X1 U6521 ( .A1(n6798), .A2(n6797), .ZN(n7365) );
  INV_X2 U6522 ( .A(n6563), .ZN(n8250) );
  AND2_X1 U6523 ( .A1(n8770), .A2(n8769), .ZN(n8936) );
  AND2_X1 U6524 ( .A1(n8367), .A2(n8368), .ZN(n8364) );
  INV_X1 U6525 ( .A(n8952), .ZN(n8943) );
  OR2_X1 U6526 ( .A1(n7804), .A2(n9997), .ZN(n10021) );
  AND2_X1 U6527 ( .A1(n6947), .A2(n6863), .ZN(n6857) );
  AND2_X1 U6528 ( .A1(n6450), .A2(n6440), .ZN(n8537) );
  INV_X1 U6529 ( .A(n9062), .ZN(n9063) );
  OR2_X1 U6530 ( .A1(n7081), .A2(n6195), .ZN(n6196) );
  OAI21_X1 U6531 ( .B1(n6189), .B2(n7474), .A(n9513), .ZN(n9167) );
  OR2_X1 U6532 ( .A1(n9367), .A2(n5637), .ZN(n5313) );
  OR2_X1 U6533 ( .A1(n5637), .A2(n7476), .ZN(n5620) );
  INV_X1 U6534 ( .A(n9720), .ZN(n9289) );
  INV_X1 U6535 ( .A(n9727), .ZN(n9338) );
  NAND2_X1 U6536 ( .A1(n9736), .A2(n7470), .ZN(n9797) );
  INV_X1 U6537 ( .A(n9916), .ZN(n9862) );
  NAND2_X1 U6538 ( .A1(n6185), .A2(n7471), .ZN(n9901) );
  NAND2_X1 U6539 ( .A1(n9872), .A2(n9901), .ZN(n9916) );
  AOI21_X1 U6540 ( .B1(n9800), .B2(n9832), .A(n6167), .ZN(n7463) );
  AND2_X1 U6541 ( .A1(n6842), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6808) );
  AND2_X1 U6542 ( .A1(n5685), .A2(n5684), .ZN(n6968) );
  INV_X1 U6543 ( .A(n6789), .ZN(n6790) );
  OR2_X1 U6544 ( .A1(n6784), .A2(n6783), .ZN(n8238) );
  INV_X1 U6545 ( .A(n8241), .ZN(n8165) );
  AND2_X1 U6546 ( .A1(n8259), .A2(n6570), .ZN(n8625) );
  INV_X1 U6547 ( .A(n8778), .ZN(n8469) );
  OR2_X1 U6548 ( .A1(n8573), .A2(n8460), .ZN(n9981) );
  INV_X1 U6549 ( .A(n9937), .ZN(n9995) );
  NAND2_X1 U6550 ( .A1(n8812), .A2(n7456), .ZN(n8793) );
  NAND2_X1 U6551 ( .A1(n10466), .A2(n10046), .ZN(n8867) );
  NAND2_X1 U6552 ( .A1(n10466), .A2(n10021), .ZN(n8862) );
  OR2_X1 U6553 ( .A1(n10049), .A2(n10029), .ZN(n8952) );
  OR2_X1 U6554 ( .A1(n10031), .A2(n10049), .ZN(n8947) );
  AND2_X1 U6555 ( .A1(n6676), .A2(n6675), .ZN(n10049) );
  AND2_X1 U6556 ( .A1(n6945), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6863) );
  INV_X1 U6557 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n10214) );
  INV_X1 U6558 ( .A(n7204), .ZN(n7216) );
  INV_X1 U6559 ( .A(n9167), .ZN(n9704) );
  NAND2_X1 U6560 ( .A1(n6196), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9708) );
  NAND2_X1 U6561 ( .A1(n5327), .A2(n5326), .ZN(n9174) );
  OR2_X1 U6562 ( .A1(n6880), .A2(n6846), .ZN(n9344) );
  AND2_X2 U6563 ( .A1(n9527), .A2(n9620), .ZN(n9936) );
  INV_X1 U6564 ( .A(n9919), .ZN(n9918) );
  CLKBUF_X1 U6565 ( .A(n9830), .Z(n9822) );
  INV_X1 U6566 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8095) );
  INV_X1 U6567 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7912) );
  INV_X1 U6568 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10364) );
  INV_X1 U6569 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6940) );
  INV_X1 U6570 ( .A(n8573), .ZN(P2_U3893) );
  INV_X1 U6571 ( .A(n9198), .ZN(P1_U3973) );
  NAND2_X1 U6572 ( .A1(n6202), .A2(n6201), .ZN(P1_U3240) );
  INV_X1 U6573 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6816) );
  INV_X1 U6574 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6813) );
  XNOR2_X1 U6575 ( .A(n5135), .B(SI_1_), .ZN(n5611) );
  AND2_X1 U6576 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5133) );
  NAND2_X1 U6577 ( .A1(n6265), .A2(n5133), .ZN(n5571) );
  NAND3_X1 U6578 ( .A1(n6814), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n5134) );
  NAND2_X1 U6579 ( .A1(n5571), .A2(n5134), .ZN(n5610) );
  NAND2_X1 U6580 ( .A1(n5611), .A2(n5610), .ZN(n5138) );
  INV_X1 U6581 ( .A(n5135), .ZN(n5136) );
  NAND2_X1 U6582 ( .A1(n5136), .A2(SI_1_), .ZN(n5137) );
  NAND2_X1 U6583 ( .A1(n5138), .A2(n5137), .ZN(n5624) );
  INV_X1 U6584 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6819) );
  INV_X1 U6585 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6812) );
  MUX2_X1 U6586 ( .A(n6819), .B(n6812), .S(n6265), .Z(n5139) );
  NAND2_X1 U6587 ( .A1(n5624), .A2(n5623), .ZN(n5142) );
  INV_X1 U6588 ( .A(n5139), .ZN(n5140) );
  NAND2_X1 U6589 ( .A1(n5140), .A2(SI_2_), .ZN(n5141) );
  NAND2_X1 U6590 ( .A1(n5142), .A2(n5141), .ZN(n5632) );
  INV_X1 U6591 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6817) );
  INV_X1 U6592 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6821) );
  MUX2_X1 U6593 ( .A(n6817), .B(n6821), .S(n6265), .Z(n5143) );
  XNOR2_X1 U6594 ( .A(n5143), .B(SI_3_), .ZN(n5631) );
  NAND2_X1 U6595 ( .A1(n5632), .A2(n5631), .ZN(n5146) );
  INV_X1 U6596 ( .A(n5143), .ZN(n5144) );
  NAND2_X1 U6597 ( .A1(n5144), .A2(SI_3_), .ZN(n5145) );
  NAND2_X1 U6598 ( .A1(n5146), .A2(n5145), .ZN(n5584) );
  INV_X1 U6599 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6822) );
  INV_X1 U6600 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6824) );
  INV_X1 U6601 ( .A(n5147), .ZN(n5148) );
  NAND2_X1 U6602 ( .A1(n5148), .A2(SI_4_), .ZN(n5149) );
  XNOR2_X1 U6603 ( .A(n5150), .B(SI_5_), .ZN(n5648) );
  INV_X1 U6604 ( .A(n5150), .ZN(n5151) );
  MUX2_X1 U6605 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6265), .Z(n5153) );
  XNOR2_X1 U6606 ( .A(n5153), .B(SI_6_), .ZN(n5601) );
  INV_X1 U6607 ( .A(n5601), .ZN(n5152) );
  NAND2_X1 U6608 ( .A1(n5602), .A2(n5152), .ZN(n5155) );
  NAND2_X1 U6609 ( .A1(n5153), .A2(SI_6_), .ZN(n5154) );
  MUX2_X1 U6610 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6265), .Z(n5157) );
  XNOR2_X1 U6611 ( .A(n5157), .B(SI_7_), .ZN(n5689) );
  INV_X1 U6612 ( .A(n5689), .ZN(n5156) );
  INV_X1 U6613 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6839) );
  INV_X1 U6614 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6837) );
  MUX2_X1 U6615 ( .A(n6839), .B(n6837), .S(n6265), .Z(n5159) );
  INV_X1 U6616 ( .A(SI_8_), .ZN(n5158) );
  NAND2_X1 U6617 ( .A1(n5159), .A2(n5158), .ZN(n5162) );
  INV_X1 U6618 ( .A(n5159), .ZN(n5160) );
  NAND2_X1 U6619 ( .A1(n5160), .A2(SI_8_), .ZN(n5161) );
  NAND2_X1 U6620 ( .A1(n5162), .A2(n5161), .ZN(n5681) );
  INV_X1 U6621 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5163) );
  MUX2_X1 U6622 ( .A(n6851), .B(n5163), .S(n6265), .Z(n5165) );
  INV_X1 U6623 ( .A(SI_9_), .ZN(n5164) );
  NAND2_X1 U6624 ( .A1(n5165), .A2(n5164), .ZN(n5168) );
  INV_X1 U6625 ( .A(n5165), .ZN(n5166) );
  NAND2_X1 U6626 ( .A1(n5166), .A2(SI_9_), .ZN(n5167) );
  MUX2_X1 U6627 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6265), .Z(n5170) );
  XNOR2_X1 U6628 ( .A(n5170), .B(n10097), .ZN(n5551) );
  INV_X1 U6629 ( .A(n5551), .ZN(n5172) );
  NAND2_X1 U6630 ( .A1(n5170), .A2(SI_10_), .ZN(n5171) );
  MUX2_X1 U6631 ( .A(n6870), .B(n10331), .S(n6265), .Z(n5174) );
  INV_X1 U6632 ( .A(SI_11_), .ZN(n5173) );
  NAND2_X1 U6633 ( .A1(n5174), .A2(n5173), .ZN(n5177) );
  INV_X1 U6634 ( .A(n5174), .ZN(n5175) );
  NAND2_X1 U6635 ( .A1(n5175), .A2(SI_11_), .ZN(n5176) );
  NAND2_X1 U6636 ( .A1(n5177), .A2(n5176), .ZN(n5539) );
  MUX2_X1 U6637 ( .A(n10343), .B(n6940), .S(n6265), .Z(n5178) );
  XNOR2_X1 U6638 ( .A(n5178), .B(SI_12_), .ZN(n5524) );
  INV_X1 U6639 ( .A(n5178), .ZN(n5179) );
  MUX2_X1 U6640 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6265), .Z(n5181) );
  XNOR2_X1 U6641 ( .A(n5181), .B(SI_13_), .ZN(n5510) );
  INV_X1 U6642 ( .A(n5510), .ZN(n5180) );
  NAND2_X1 U6643 ( .A1(n5511), .A2(n5180), .ZN(n5183) );
  NAND2_X1 U6644 ( .A1(n5181), .A2(SI_13_), .ZN(n5182) );
  NAND2_X1 U6645 ( .A1(n5183), .A2(n5182), .ZN(n5479) );
  MUX2_X1 U6646 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6265), .Z(n5185) );
  XNOR2_X1 U6647 ( .A(n5185), .B(SI_14_), .ZN(n5478) );
  INV_X1 U6648 ( .A(n5478), .ZN(n5184) );
  NAND2_X1 U6649 ( .A1(n5479), .A2(n5184), .ZN(n5187) );
  NAND2_X1 U6650 ( .A1(n5185), .A2(SI_14_), .ZN(n5186) );
  MUX2_X1 U6651 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6265), .Z(n5491) );
  NOR2_X1 U6652 ( .A1(n5189), .A2(n5188), .ZN(n5191) );
  NAND2_X1 U6653 ( .A1(n5189), .A2(n5188), .ZN(n5190) );
  MUX2_X1 U6654 ( .A(n7149), .B(n7180), .S(n6265), .Z(n5463) );
  NOR2_X1 U6655 ( .A1(n5192), .A2(SI_16_), .ZN(n5194) );
  NAND2_X1 U6656 ( .A1(n5192), .A2(SI_16_), .ZN(n5193) );
  MUX2_X1 U6657 ( .A(n10284), .B(n10364), .S(n6265), .Z(n5196) );
  NAND2_X1 U6658 ( .A1(n5196), .A2(n5195), .ZN(n5199) );
  INV_X1 U6659 ( .A(n5196), .ZN(n5197) );
  NAND2_X1 U6660 ( .A1(n5197), .A2(SI_17_), .ZN(n5198) );
  NAND2_X1 U6661 ( .A1(n5199), .A2(n5198), .ZN(n5451) );
  MUX2_X1 U6662 ( .A(n10233), .B(n5200), .S(n6265), .Z(n5201) );
  XNOR2_X1 U6663 ( .A(n5201), .B(SI_18_), .ZN(n5438) );
  INV_X1 U6664 ( .A(n5201), .ZN(n5202) );
  NAND2_X1 U6665 ( .A1(n5202), .A2(SI_18_), .ZN(n5203) );
  INV_X1 U6666 ( .A(n5413), .ZN(n5208) );
  MUX2_X1 U6667 ( .A(n7617), .B(n8100), .S(n6265), .Z(n5204) );
  NAND2_X1 U6668 ( .A1(n5204), .A2(n10294), .ZN(n5209) );
  INV_X1 U6669 ( .A(n5204), .ZN(n5205) );
  NAND2_X1 U6670 ( .A1(n5205), .A2(SI_19_), .ZN(n5206) );
  NAND2_X1 U6671 ( .A1(n5209), .A2(n5206), .ZN(n5412) );
  INV_X1 U6672 ( .A(n5412), .ZN(n5207) );
  NAND2_X1 U6673 ( .A1(n5208), .A2(n5207), .ZN(n5210) );
  MUX2_X1 U6674 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6265), .Z(n5389) );
  INV_X1 U6675 ( .A(n5389), .ZN(n5211) );
  MUX2_X1 U6676 ( .A(n7774), .B(n7776), .S(n6265), .Z(n5397) );
  NOR2_X1 U6677 ( .A1(n5212), .A2(SI_21_), .ZN(n5213) );
  MUX2_X1 U6678 ( .A(n7868), .B(n7865), .S(n6265), .Z(n5215) );
  INV_X1 U6679 ( .A(SI_22_), .ZN(n5214) );
  NAND2_X1 U6680 ( .A1(n5215), .A2(n5214), .ZN(n5218) );
  INV_X1 U6681 ( .A(n5215), .ZN(n5216) );
  NAND2_X1 U6682 ( .A1(n5216), .A2(SI_22_), .ZN(n5217) );
  NAND2_X1 U6683 ( .A1(n5218), .A2(n5217), .ZN(n5376) );
  MUX2_X1 U6684 ( .A(n10214), .B(n7912), .S(n6265), .Z(n5219) );
  NAND2_X1 U6685 ( .A1(n5219), .A2(n10219), .ZN(n5222) );
  INV_X1 U6686 ( .A(n5219), .ZN(n5220) );
  NAND2_X1 U6687 ( .A1(n5220), .A2(SI_23_), .ZN(n5221) );
  INV_X1 U6688 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7939) );
  INV_X1 U6689 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7963) );
  MUX2_X1 U6690 ( .A(n7939), .B(n7963), .S(n6265), .Z(n5225) );
  INV_X1 U6691 ( .A(SI_24_), .ZN(n5224) );
  NAND2_X1 U6692 ( .A1(n5225), .A2(n5224), .ZN(n5228) );
  INV_X1 U6693 ( .A(n5225), .ZN(n5226) );
  NAND2_X1 U6694 ( .A1(n5226), .A2(SI_24_), .ZN(n5227) );
  INV_X1 U6695 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7992) );
  INV_X1 U6696 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8000) );
  MUX2_X1 U6697 ( .A(n7992), .B(n8000), .S(n6265), .Z(n5230) );
  INV_X1 U6698 ( .A(SI_25_), .ZN(n5229) );
  NAND2_X1 U6699 ( .A1(n5230), .A2(n5229), .ZN(n5233) );
  INV_X1 U6700 ( .A(n5230), .ZN(n5231) );
  NAND2_X1 U6701 ( .A1(n5231), .A2(SI_25_), .ZN(n5232) );
  INV_X1 U6702 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8023) );
  INV_X1 U6703 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8025) );
  MUX2_X1 U6704 ( .A(n8023), .B(n8025), .S(n6265), .Z(n5236) );
  INV_X1 U6705 ( .A(SI_26_), .ZN(n5235) );
  NAND2_X1 U6706 ( .A1(n5236), .A2(n5235), .ZN(n5239) );
  INV_X1 U6707 ( .A(n5236), .ZN(n5237) );
  NAND2_X1 U6708 ( .A1(n5237), .A2(SI_26_), .ZN(n5238) );
  NAND2_X1 U6709 ( .A1(n5329), .A2(n5330), .ZN(n5240) );
  INV_X1 U6710 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6540) );
  INV_X1 U6711 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10342) );
  MUX2_X1 U6712 ( .A(n6540), .B(n10342), .S(n6265), .Z(n5242) );
  INV_X1 U6713 ( .A(SI_27_), .ZN(n5241) );
  NAND2_X1 U6714 ( .A1(n5242), .A2(n5241), .ZN(n5245) );
  INV_X1 U6715 ( .A(n5242), .ZN(n5243) );
  NAND2_X1 U6716 ( .A1(n5243), .A2(SI_27_), .ZN(n5244) );
  NAND2_X1 U6717 ( .A1(n5315), .A2(n5316), .ZN(n5246) );
  NAND2_X1 U6718 ( .A1(n5246), .A2(n5245), .ZN(n5303) );
  INV_X1 U6719 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6551) );
  MUX2_X1 U6720 ( .A(n6551), .B(n8095), .S(n6265), .Z(n5248) );
  INV_X1 U6721 ( .A(SI_28_), .ZN(n5247) );
  NAND2_X1 U6722 ( .A1(n5248), .A2(n5247), .ZN(n5251) );
  INV_X1 U6723 ( .A(n5248), .ZN(n5249) );
  NAND2_X1 U6724 ( .A1(n5249), .A2(SI_28_), .ZN(n5250) );
  NAND2_X1 U6725 ( .A1(n5303), .A2(n5304), .ZN(n5252) );
  MUX2_X1 U6726 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6265), .Z(n5720) );
  INV_X1 U6727 ( .A(n5253), .ZN(n5255) );
  INV_X1 U6728 ( .A(SI_29_), .ZN(n5254) );
  NAND2_X1 U6729 ( .A1(n5255), .A2(n5254), .ZN(n5256) );
  NOR2_X2 U6730 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5581) );
  NAND3_X1 U6731 ( .A1(n5581), .A2(n5582), .A3(n5257), .ZN(n5598) );
  INV_X1 U6732 ( .A(n5598), .ZN(n5259) );
  NAND4_X1 U6733 ( .A1(n5263), .A2(n5262), .A3(n5261), .A4(n5260), .ZN(n5264)
         );
  INV_X1 U6734 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5266) );
  NAND2_X1 U6735 ( .A1(n5943), .A2(n5267), .ZN(n5285) );
  NAND2_X1 U6736 ( .A1(n5285), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5268) );
  NOR2_X2 U6737 ( .A1(n5272), .A2(n5269), .ZN(n5271) );
  INV_X1 U6738 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9632) );
  OR2_X1 U6739 ( .A1(n4516), .A2(n9632), .ZN(n5273) );
  NAND2_X1 U6740 ( .A1(n5654), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5653) );
  INV_X1 U6741 ( .A(n5502), .ZN(n5277) );
  OR2_X2 U6742 ( .A1(n5458), .A2(n9152), .ZN(n5445) );
  INV_X1 U6743 ( .A(n5405), .ZN(n5281) );
  INV_X1 U6744 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9009) );
  INV_X1 U6745 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9087) );
  INV_X1 U6746 ( .A(n5359), .ZN(n5282) );
  INV_X1 U6747 ( .A(n5346), .ZN(n5283) );
  NAND2_X1 U6748 ( .A1(n5283), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5334) );
  INV_X1 U6749 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5319) );
  INV_X1 U6750 ( .A(n5321), .ZN(n5284) );
  NAND2_X1 U6751 ( .A1(n5284), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8074) );
  INV_X1 U6752 ( .A(n5285), .ZN(n5287) );
  NOR2_X1 U6753 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5286) );
  XNOR2_X2 U6754 ( .A(n5291), .B(n5290), .ZN(n5294) );
  OR2_X1 U6755 ( .A1(n8074), .A2(n5637), .ZN(n5301) );
  INV_X1 U6756 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5298) );
  INV_X2 U6757 ( .A(n5617), .ZN(n5740) );
  NAND2_X1 U6758 ( .A1(n5695), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5297) );
  INV_X1 U6759 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n8073) );
  OR2_X1 U6760 ( .A1(n5741), .A2(n8073), .ZN(n5296) );
  OAI211_X1 U6761 ( .C1(n5298), .C2(n5591), .A(n5297), .B(n5296), .ZN(n5299)
         );
  INV_X1 U6762 ( .A(n5299), .ZN(n5300) );
  NAND2_X1 U6763 ( .A1(n5301), .A2(n5300), .ZN(n9172) );
  INV_X1 U6764 ( .A(n9172), .ZN(n5302) );
  NAND2_X1 U6765 ( .A1(n9532), .A2(n5302), .ZN(n5874) );
  NAND2_X1 U6766 ( .A1(n8094), .A2(n5737), .ZN(n5306) );
  OR2_X1 U6767 ( .A1(n4517), .A2(n8095), .ZN(n5305) );
  INV_X1 U6768 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9027) );
  NAND2_X1 U6769 ( .A1(n5321), .A2(n9027), .ZN(n5307) );
  NAND2_X1 U6770 ( .A1(n8074), .A2(n5307), .ZN(n9367) );
  INV_X1 U6771 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10237) );
  NAND2_X1 U6772 ( .A1(n5673), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5310) );
  INV_X1 U6773 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5308) );
  OR2_X1 U6774 ( .A1(n5617), .A2(n5308), .ZN(n5309) );
  OAI211_X1 U6775 ( .C1(n5591), .C2(n10237), .A(n5310), .B(n5309), .ZN(n5311)
         );
  INV_X1 U6776 ( .A(n5311), .ZN(n5312) );
  NOR2_X1 U6777 ( .A1(n9538), .A2(n8068), .ZN(n8038) );
  NAND2_X1 U6778 ( .A1(n9538), .A2(n8068), .ZN(n8037) );
  INV_X1 U6779 ( .A(n8037), .ZN(n5314) );
  NAND2_X1 U6780 ( .A1(n8096), .A2(n5737), .ZN(n5318) );
  OR2_X1 U6781 ( .A1(n4516), .A2(n10342), .ZN(n5317) );
  NAND2_X1 U6782 ( .A1(n5334), .A2(n5319), .ZN(n5320) );
  INV_X1 U6783 ( .A(n5637), .ZN(n5446) );
  NAND2_X1 U6784 ( .A1(n9381), .A2(n5446), .ZN(n5327) );
  INV_X1 U6785 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10107) );
  NAND2_X1 U6786 ( .A1(n5673), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5324) );
  INV_X1 U6787 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n5322) );
  OR2_X1 U6788 ( .A1(n5617), .A2(n5322), .ZN(n5323) );
  OAI211_X1 U6789 ( .C1(n5591), .C2(n10107), .A(n5324), .B(n5323), .ZN(n5325)
         );
  INV_X1 U6790 ( .A(n5325), .ZN(n5326) );
  INV_X1 U6791 ( .A(n9174), .ZN(n5328) );
  NAND2_X1 U6792 ( .A1(n9543), .A2(n5328), .ZN(n8036) );
  NAND2_X1 U6793 ( .A1(n8022), .A2(n5737), .ZN(n5332) );
  OR2_X1 U6794 ( .A1(n4517), .A2(n8025), .ZN(n5331) );
  INV_X1 U6795 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n10122) );
  NAND2_X1 U6796 ( .A1(n5346), .A2(n10122), .ZN(n5333) );
  NAND2_X1 U6797 ( .A1(n5334), .A2(n5333), .ZN(n8082) );
  INV_X1 U6798 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5337) );
  NAND2_X1 U6799 ( .A1(n5673), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U6800 ( .A1(n5695), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5335) );
  OAI211_X1 U6801 ( .C1(n5337), .C2(n5591), .A(n5336), .B(n5335), .ZN(n5338)
         );
  INV_X1 U6802 ( .A(n5338), .ZN(n5339) );
  OR2_X1 U6803 ( .A1(n9546), .A2(n8065), .ZN(n5801) );
  NAND2_X1 U6804 ( .A1(n9546), .A2(n8065), .ZN(n8035) );
  XNOR2_X1 U6805 ( .A(n5342), .B(n5341), .ZN(n7991) );
  NAND2_X1 U6806 ( .A1(n7991), .A2(n5737), .ZN(n5344) );
  OR2_X1 U6807 ( .A1(n4516), .A2(n8000), .ZN(n5343) );
  INV_X1 U6808 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10359) );
  NAND2_X1 U6809 ( .A1(n5359), .A2(n10359), .ZN(n5345) );
  NAND2_X1 U6810 ( .A1(n5346), .A2(n5345), .ZN(n9389) );
  INV_X1 U6811 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U6812 ( .A1(n5673), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U6813 ( .A1(n5695), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5347) );
  OAI211_X1 U6814 ( .C1(n5349), .C2(n5591), .A(n5348), .B(n5347), .ZN(n5350)
         );
  INV_X1 U6815 ( .A(n5350), .ZN(n5351) );
  INV_X1 U6816 ( .A(n9176), .ZN(n5353) );
  OR2_X1 U6817 ( .A1(n9552), .A2(n5353), .ZN(n5800) );
  NAND2_X1 U6818 ( .A1(n9552), .A2(n5353), .ZN(n8033) );
  XNOR2_X1 U6819 ( .A(n5355), .B(n5354), .ZN(n7938) );
  NAND2_X1 U6820 ( .A1(n7938), .A2(n5737), .ZN(n5357) );
  OR2_X1 U6821 ( .A1(n4517), .A2(n7963), .ZN(n5356) );
  NAND2_X1 U6822 ( .A1(n5370), .A2(n9087), .ZN(n5358) );
  AND2_X1 U6823 ( .A1(n5359), .A2(n5358), .ZN(n9404) );
  NAND2_X1 U6824 ( .A1(n9404), .A2(n5446), .ZN(n5364) );
  INV_X1 U6825 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10268) );
  NAND2_X1 U6826 ( .A1(n5673), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6827 ( .A1(n5695), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5360) );
  OAI211_X1 U6828 ( .C1(n10268), .C2(n5591), .A(n5361), .B(n5360), .ZN(n5362)
         );
  INV_X1 U6829 ( .A(n5362), .ZN(n5363) );
  INV_X1 U6830 ( .A(n9177), .ZN(n8061) );
  NAND2_X1 U6831 ( .A1(n9557), .A2(n8061), .ZN(n5855) );
  NAND2_X1 U6832 ( .A1(n9392), .A2(n5855), .ZN(n9408) );
  XNOR2_X1 U6833 ( .A(n5366), .B(n5365), .ZN(n7914) );
  NAND2_X1 U6834 ( .A1(n7914), .A2(n5737), .ZN(n5368) );
  OR2_X1 U6835 ( .A1(n4516), .A2(n7912), .ZN(n5367) );
  NAND2_X1 U6836 ( .A1(n5382), .A2(n9009), .ZN(n5369) );
  NAND2_X1 U6837 ( .A1(n5370), .A2(n5369), .ZN(n9007) );
  OR2_X1 U6838 ( .A1(n9007), .A2(n5637), .ZN(n5375) );
  INV_X1 U6839 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10278) );
  NAND2_X1 U6840 ( .A1(n5673), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5372) );
  NAND2_X1 U6841 ( .A1(n5695), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5371) );
  OAI211_X1 U6842 ( .C1(n10278), .C2(n5591), .A(n5372), .B(n5371), .ZN(n5373)
         );
  INV_X1 U6843 ( .A(n5373), .ZN(n5374) );
  NAND2_X1 U6844 ( .A1(n5375), .A2(n5374), .ZN(n9178) );
  OR2_X1 U6845 ( .A1(n9563), .A2(n8060), .ZN(n5854) );
  NAND2_X1 U6846 ( .A1(n9563), .A2(n8060), .ZN(n5851) );
  NAND2_X1 U6847 ( .A1(n5854), .A2(n5851), .ZN(n9416) );
  XNOR2_X1 U6848 ( .A(n5377), .B(n5376), .ZN(n7864) );
  NAND2_X1 U6849 ( .A1(n7864), .A2(n5737), .ZN(n5379) );
  OR2_X1 U6850 ( .A1(n4516), .A2(n7865), .ZN(n5378) );
  INV_X1 U6851 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U6852 ( .A1(n5405), .A2(n5380), .ZN(n5381) );
  NAND2_X1 U6853 ( .A1(n5382), .A2(n5381), .ZN(n9432) );
  OR2_X1 U6854 ( .A1(n9432), .A2(n5637), .ZN(n5388) );
  INV_X1 U6855 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U6856 ( .A1(n5695), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U6857 ( .A1(n5673), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5383) );
  OAI211_X1 U6858 ( .C1(n5591), .C2(n5385), .A(n5384), .B(n5383), .ZN(n5386)
         );
  INV_X1 U6859 ( .A(n5386), .ZN(n5387) );
  NAND2_X1 U6860 ( .A1(n5388), .A2(n5387), .ZN(n9179) );
  XNOR2_X1 U6861 ( .A(n9567), .B(n9179), .ZN(n9436) );
  INV_X1 U6862 ( .A(n9436), .ZN(n9427) );
  XNOR2_X1 U6863 ( .A(n5389), .B(n10270), .ZN(n5390) );
  XNOR2_X1 U6864 ( .A(n5391), .B(n5390), .ZN(n7658) );
  NAND2_X1 U6865 ( .A1(n7658), .A2(n5737), .ZN(n5393) );
  INV_X1 U6866 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7657) );
  OR2_X1 U6867 ( .A1(n4517), .A2(n7657), .ZN(n5392) );
  NAND2_X1 U6868 ( .A1(n5430), .A2(n9114), .ZN(n5394) );
  NAND2_X1 U6869 ( .A1(n5403), .A2(n5394), .ZN(n9466) );
  AOI22_X1 U6870 ( .A1(n5618), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n5695), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U6871 ( .A1(n5673), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5395) );
  OAI211_X1 U6872 ( .C1(n9466), .C2(n5637), .A(n5396), .B(n5395), .ZN(n9181)
         );
  INV_X1 U6873 ( .A(n9181), .ZN(n8053) );
  OR2_X1 U6874 ( .A1(n9578), .A2(n8053), .ZN(n8031) );
  NAND2_X1 U6875 ( .A1(n9578), .A2(n8053), .ZN(n5834) );
  XNOR2_X1 U6876 ( .A(n5397), .B(SI_21_), .ZN(n5398) );
  XNOR2_X1 U6877 ( .A(n5399), .B(n5398), .ZN(n7773) );
  NAND2_X1 U6878 ( .A1(n7773), .A2(n5737), .ZN(n5401) );
  OR2_X1 U6879 ( .A1(n4517), .A2(n7776), .ZN(n5400) );
  INV_X1 U6880 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U6881 ( .A1(n5403), .A2(n5402), .ZN(n5404) );
  NAND2_X1 U6882 ( .A1(n5405), .A2(n5404), .ZN(n9445) );
  OR2_X1 U6883 ( .A1(n9445), .A2(n5637), .ZN(n5411) );
  INV_X1 U6884 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5408) );
  NAND2_X1 U6885 ( .A1(n5695), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U6886 ( .A1(n5673), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5406) );
  OAI211_X1 U6887 ( .C1(n5591), .C2(n5408), .A(n5407), .B(n5406), .ZN(n5409)
         );
  INV_X1 U6888 ( .A(n5409), .ZN(n5410) );
  NAND2_X1 U6889 ( .A1(n5411), .A2(n5410), .ZN(n9180) );
  INV_X1 U6890 ( .A(n9180), .ZN(n8056) );
  OR2_X1 U6891 ( .A1(n9572), .A2(n8056), .ZN(n5847) );
  NAND2_X1 U6892 ( .A1(n9572), .A2(n8056), .ZN(n8032) );
  NAND2_X1 U6893 ( .A1(n5847), .A2(n8032), .ZN(n9449) );
  XNOR2_X1 U6894 ( .A(n5413), .B(n5412), .ZN(n7616) );
  NAND2_X1 U6895 ( .A1(n7616), .A2(n5737), .ZN(n5427) );
  AND2_X2 U6896 ( .A1(n5526), .A2(n5414), .ZN(n5512) );
  NAND2_X1 U6897 ( .A1(n5453), .A2(n5415), .ZN(n5440) );
  INV_X1 U6898 ( .A(n5440), .ZN(n5419) );
  INV_X1 U6899 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5417) );
  INV_X1 U6900 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5416) );
  AND2_X1 U6901 ( .A1(n5417), .A2(n5416), .ZN(n5418) );
  NAND2_X1 U6902 ( .A1(n5419), .A2(n5418), .ZN(n5425) );
  NAND2_X1 U6903 ( .A1(n5440), .A2(n5420), .ZN(n5424) );
  NAND2_X1 U6904 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n5422) );
  NAND2_X1 U6905 ( .A1(n4609), .A2(n5118), .ZN(n5423) );
  AOI22_X1 U6906 ( .A1(n5686), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5883), .B2(
        n5692), .ZN(n5426) );
  INV_X1 U6907 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n5437) );
  INV_X1 U6908 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5428) );
  NAND2_X1 U6909 ( .A1(n5445), .A2(n5428), .ZN(n5429) );
  NAND2_X1 U6910 ( .A1(n5430), .A2(n5429), .ZN(n9475) );
  OR2_X1 U6911 ( .A1(n9475), .A2(n5637), .ZN(n5436) );
  INV_X1 U6912 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n5431) );
  OR2_X1 U6913 ( .A1(n5741), .A2(n5431), .ZN(n5434) );
  INV_X1 U6914 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n5432) );
  OR2_X1 U6915 ( .A1(n5617), .A2(n5432), .ZN(n5433) );
  AND2_X1 U6916 ( .A1(n5434), .A2(n5433), .ZN(n5435) );
  OAI211_X1 U6917 ( .C1(n5591), .C2(n5437), .A(n5436), .B(n5435), .ZN(n9182)
         );
  INV_X1 U6918 ( .A(n9182), .ZN(n8051) );
  OR2_X1 U6919 ( .A1(n9582), .A2(n8051), .ZN(n5833) );
  NAND2_X1 U6920 ( .A1(n9582), .A2(n8051), .ZN(n5915) );
  XNOR2_X1 U6921 ( .A(n5439), .B(n5438), .ZN(n7388) );
  NAND2_X1 U6922 ( .A1(n7388), .A2(n5737), .ZN(n5443) );
  NAND2_X1 U6923 ( .A1(n5440), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5441) );
  XNOR2_X1 U6924 ( .A(n5441), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9325) );
  AOI22_X1 U6925 ( .A1(n5686), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5692), .B2(
        n9325), .ZN(n5442) );
  NAND2_X1 U6926 ( .A1(n5458), .A2(n9152), .ZN(n5444) );
  AND2_X1 U6927 ( .A1(n5445), .A2(n5444), .ZN(n9497) );
  NAND2_X1 U6928 ( .A1(n9497), .A2(n5446), .ZN(n5450) );
  NAND2_X1 U6929 ( .A1(n5695), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U6930 ( .A1(n5673), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5448) );
  INV_X1 U6931 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10109) );
  OR2_X1 U6932 ( .A1(n5743), .A2(n10109), .ZN(n5447) );
  NAND4_X1 U6933 ( .A1(n5450), .A2(n5449), .A3(n5448), .A4(n5447), .ZN(n9183)
         );
  INV_X1 U6934 ( .A(n9183), .ZN(n8049) );
  OR2_X1 U6935 ( .A1(n9588), .A2(n8049), .ZN(n5837) );
  NAND2_X1 U6936 ( .A1(n9588), .A2(n8049), .ZN(n5838) );
  XNOR2_X1 U6937 ( .A(n5452), .B(n5451), .ZN(n7375) );
  NAND2_X1 U6938 ( .A1(n7375), .A2(n5737), .ZN(n5455) );
  XNOR2_X1 U6939 ( .A(n5453), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9318) );
  AOI22_X1 U6940 ( .A1(n5686), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5692), .B2(
        n9318), .ZN(n5454) );
  NAND2_X1 U6941 ( .A1(n5695), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5462) );
  INV_X1 U6942 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9515) );
  OR2_X1 U6943 ( .A1(n5741), .A2(n9515), .ZN(n5461) );
  INV_X1 U6944 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U6945 ( .A1(n5472), .A2(n5456), .ZN(n5457) );
  NAND2_X1 U6946 ( .A1(n5458), .A2(n5457), .ZN(n9514) );
  OR2_X1 U6947 ( .A1(n5637), .A2(n9514), .ZN(n5460) );
  INV_X1 U6948 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9302) );
  OR2_X1 U6949 ( .A1(n5591), .A2(n9302), .ZN(n5459) );
  NAND4_X1 U6950 ( .A1(n5462), .A2(n5461), .A3(n5460), .A4(n5459), .ZN(n9184)
         );
  INV_X1 U6951 ( .A(n9184), .ZN(n8047) );
  NAND2_X1 U6952 ( .A1(n9521), .A2(n8047), .ZN(n5832) );
  XNOR2_X1 U6953 ( .A(n5463), .B(SI_16_), .ZN(n5464) );
  XNOR2_X1 U6954 ( .A(n5465), .B(n5464), .ZN(n7148) );
  NAND2_X1 U6955 ( .A1(n7148), .A2(n5737), .ZN(n5469) );
  NAND2_X1 U6956 ( .A1(n5466), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5467) );
  XNOR2_X1 U6957 ( .A(n5467), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9305) );
  AOI22_X1 U6958 ( .A1(n5686), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5692), .B2(
        n9305), .ZN(n5468) );
  NAND2_X1 U6959 ( .A1(n5740), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5476) );
  INV_X1 U6960 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9287) );
  OR2_X1 U6961 ( .A1(n5741), .A2(n9287), .ZN(n5475) );
  NAND2_X1 U6962 ( .A1(n5504), .A2(n5470), .ZN(n5471) );
  NAND2_X1 U6963 ( .A1(n5472), .A2(n5471), .ZN(n9652) );
  OR2_X1 U6964 ( .A1(n5637), .A2(n9652), .ZN(n5474) );
  INV_X1 U6965 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9277) );
  OR2_X1 U6966 ( .A1(n5591), .A2(n9277), .ZN(n5473) );
  NAND4_X1 U6967 ( .A1(n5476), .A2(n5475), .A3(n5474), .A4(n5473), .ZN(n9185)
         );
  INV_X1 U6968 ( .A(n9185), .ZN(n5477) );
  OR2_X1 U6969 ( .A1(n9654), .A2(n5477), .ZN(n5828) );
  NAND2_X1 U6970 ( .A1(n9654), .A2(n5477), .ZN(n9506) );
  NAND2_X1 U6971 ( .A1(n5828), .A2(n9506), .ZN(n9655) );
  XNOR2_X1 U6972 ( .A(n5479), .B(n5478), .ZN(n6976) );
  NAND2_X1 U6973 ( .A1(n6976), .A2(n5737), .ZN(n5482) );
  NAND2_X1 U6974 ( .A1(n5480), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5495) );
  XNOR2_X1 U6975 ( .A(n5495), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7855) );
  AOI22_X1 U6976 ( .A1(n5686), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5692), .B2(
        n7855), .ZN(n5481) );
  NAND2_X1 U6977 ( .A1(n5673), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5489) );
  INV_X1 U6978 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5483) );
  OR2_X1 U6979 ( .A1(n5617), .A2(n5483), .ZN(n5488) );
  INV_X1 U6980 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U6981 ( .A1(n5519), .A2(n5484), .ZN(n5485) );
  NAND2_X1 U6982 ( .A1(n5502), .A2(n5485), .ZN(n9733) );
  OR2_X1 U6983 ( .A1(n5637), .A2(n9733), .ZN(n5487) );
  INV_X1 U6984 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7619) );
  OR2_X1 U6985 ( .A1(n5591), .A2(n7619), .ZN(n5486) );
  NAND4_X1 U6986 ( .A1(n5489), .A2(n5488), .A3(n5487), .A4(n5486), .ZN(n9187)
         );
  INV_X1 U6987 ( .A(n9187), .ZN(n5490) );
  NAND2_X1 U6988 ( .A1(n9735), .A2(n5490), .ZN(n5821) );
  XNOR2_X1 U6989 ( .A(n5491), .B(SI_15_), .ZN(n5492) );
  XNOR2_X1 U6990 ( .A(n5493), .B(n5492), .ZN(n6985) );
  NAND2_X1 U6991 ( .A1(n6985), .A2(n5737), .ZN(n5499) );
  NAND2_X1 U6992 ( .A1(n5495), .A2(n5494), .ZN(n5496) );
  NAND2_X1 U6993 ( .A1(n5496), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5497) );
  XNOR2_X1 U6994 ( .A(n5497), .B(P1_IR_REG_15__SCAN_IN), .ZN(n7857) );
  AOI22_X1 U6995 ( .A1(n5686), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5692), .B2(
        n7857), .ZN(n5498) );
  NAND2_X1 U6996 ( .A1(n5618), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5508) );
  INV_X1 U6997 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5500) );
  OR2_X1 U6998 ( .A1(n5617), .A2(n5500), .ZN(n5507) );
  INV_X1 U6999 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7957) );
  OR2_X1 U7000 ( .A1(n5741), .A2(n7957), .ZN(n5506) );
  INV_X1 U7001 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U7002 ( .A1(n5502), .A2(n5501), .ZN(n5503) );
  NAND2_X1 U7003 ( .A1(n5504), .A2(n5503), .ZN(n9165) );
  OR2_X1 U7004 ( .A1(n5637), .A2(n9165), .ZN(n5505) );
  NAND4_X1 U7005 ( .A1(n5508), .A2(n5507), .A3(n5506), .A4(n5505), .ZN(n9186)
         );
  INV_X1 U7006 ( .A(n9186), .ZN(n5509) );
  OR2_X1 U7007 ( .A1(n9168), .A2(n5509), .ZN(n5823) );
  NAND2_X1 U7008 ( .A1(n9168), .A2(n5509), .ZN(n5820) );
  NAND2_X1 U7009 ( .A1(n5823), .A2(n5820), .ZN(n7956) );
  XNOR2_X1 U7010 ( .A(n5511), .B(n5510), .ZN(n6941) );
  NAND2_X1 U7011 ( .A1(n6941), .A2(n5737), .ZN(n5516) );
  NOR2_X1 U7012 ( .A1(n5512), .A2(n5421), .ZN(n5514) );
  XNOR2_X1 U7013 ( .A(n5514), .B(n5513), .ZN(n7623) );
  AOI22_X1 U7014 ( .A1(n5686), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5692), .B2(
        n7623), .ZN(n5515) );
  NAND2_X1 U7015 ( .A1(n5673), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5523) );
  INV_X1 U7016 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5517) );
  OR2_X1 U7017 ( .A1(n5617), .A2(n5517), .ZN(n5522) );
  NAND2_X1 U7018 ( .A1(n5533), .A2(n10363), .ZN(n5518) );
  NAND2_X1 U7019 ( .A1(n5519), .A2(n5518), .ZN(n9123) );
  OR2_X1 U7020 ( .A1(n5637), .A2(n9123), .ZN(n5521) );
  INV_X1 U7021 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7421) );
  OR2_X1 U7022 ( .A1(n5591), .A2(n7421), .ZN(n5520) );
  NAND4_X1 U7023 ( .A1(n5523), .A2(n5522), .A3(n5521), .A4(n5520), .ZN(n9188)
         );
  INV_X1 U7024 ( .A(n9188), .ZN(n5768) );
  OR2_X1 U7025 ( .A1(n9125), .A2(n5768), .ZN(n5906) );
  NAND2_X1 U7026 ( .A1(n9125), .A2(n5768), .ZN(n5905) );
  XNOR2_X1 U7027 ( .A(n5525), .B(n5524), .ZN(n6938) );
  NAND2_X1 U7028 ( .A1(n6938), .A2(n5737), .ZN(n5530) );
  INV_X1 U7029 ( .A(n5526), .ZN(n5527) );
  NAND2_X1 U7030 ( .A1(n5527), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5528) );
  XNOR2_X1 U7031 ( .A(n5528), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7423) );
  AOI22_X1 U7032 ( .A1(n5686), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5692), .B2(
        n7423), .ZN(n5529) );
  NAND2_X1 U7033 ( .A1(n5740), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5538) );
  INV_X1 U7034 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7833) );
  OR2_X1 U7035 ( .A1(n5741), .A2(n7833), .ZN(n5537) );
  NAND2_X1 U7036 ( .A1(n5546), .A2(n5531), .ZN(n5532) );
  NAND2_X1 U7037 ( .A1(n5533), .A2(n5532), .ZN(n9049) );
  OR2_X1 U7038 ( .A1(n5637), .A2(n9049), .ZN(n5536) );
  INV_X1 U7039 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5534) );
  OR2_X1 U7040 ( .A1(n5743), .A2(n5534), .ZN(n5535) );
  NAND4_X1 U7041 ( .A1(n5538), .A2(n5537), .A3(n5536), .A4(n5535), .ZN(n9189)
         );
  INV_X1 U7042 ( .A(n9189), .ZN(n5710) );
  NAND2_X1 U7043 ( .A1(n9051), .A2(n5710), .ZN(n5904) );
  XNOR2_X1 U7044 ( .A(n5540), .B(n5539), .ZN(n6868) );
  NAND2_X1 U7045 ( .A1(n6868), .A2(n5737), .ZN(n5544) );
  NAND2_X1 U7046 ( .A1(n5541), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5542) );
  XNOR2_X1 U7047 ( .A(n5542), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7308) );
  AOI22_X1 U7048 ( .A1(n5686), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5692), .B2(
        n7308), .ZN(n5543) );
  NAND2_X1 U7049 ( .A1(n5740), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5550) );
  INV_X1 U7050 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10361) );
  NAND2_X1 U7051 ( .A1(n5560), .A2(n10361), .ZN(n5545) );
  NAND2_X1 U7052 ( .A1(n5546), .A2(n5545), .ZN(n9145) );
  OR2_X1 U7053 ( .A1(n5637), .A2(n9145), .ZN(n5549) );
  INV_X1 U7054 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7135) );
  OR2_X1 U7055 ( .A1(n5591), .A2(n7135), .ZN(n5548) );
  INV_X1 U7056 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7794) );
  OR2_X1 U7057 ( .A1(n5741), .A2(n7794), .ZN(n5547) );
  NAND4_X1 U7058 ( .A1(n5550), .A2(n5549), .A3(n5548), .A4(n5547), .ZN(n9190)
         );
  INV_X1 U7059 ( .A(n9190), .ZN(n5711) );
  NAND2_X1 U7060 ( .A1(n9897), .A2(n5711), .ZN(n5813) );
  XNOR2_X1 U7061 ( .A(n5552), .B(n5551), .ZN(n6853) );
  NAND2_X1 U7062 ( .A1(n6853), .A2(n5737), .ZN(n5557) );
  NAND2_X1 U7063 ( .A1(n5553), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5554) );
  MUX2_X1 U7064 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5554), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5555) );
  AND2_X1 U7065 ( .A1(n5555), .A2(n5541), .ZN(n7139) );
  AOI22_X1 U7066 ( .A1(n5686), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5692), .B2(
        n7139), .ZN(n5556) );
  NAND2_X1 U7067 ( .A1(n5557), .A2(n5556), .ZN(n7787) );
  NAND2_X1 U7068 ( .A1(n5740), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7069 ( .A1(n5668), .A2(n5558), .ZN(n5559) );
  NAND2_X1 U7070 ( .A1(n5560), .A2(n5559), .ZN(n9646) );
  OR2_X1 U7071 ( .A1(n5637), .A2(n9646), .ZN(n5563) );
  INV_X1 U7072 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6965) );
  OR2_X1 U7073 ( .A1(n5743), .A2(n6965), .ZN(n5562) );
  INV_X1 U7074 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6962) );
  OR2_X1 U7075 ( .A1(n5741), .A2(n6962), .ZN(n5561) );
  NAND4_X1 U7076 ( .A1(n5564), .A2(n5563), .A3(n5562), .A4(n5561), .ZN(n9191)
         );
  INV_X1 U7077 ( .A(n9191), .ZN(n6067) );
  OR2_X1 U7078 ( .A1(n7787), .A2(n6067), .ZN(n5900) );
  NAND2_X1 U7079 ( .A1(n7787), .A2(n6067), .ZN(n7779) );
  INV_X1 U7080 ( .A(n7829), .ZN(n5763) );
  INV_X1 U7081 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5565) );
  OR2_X1 U7082 ( .A1(n5741), .A2(n5565), .ZN(n5568) );
  INV_X1 U7083 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9710) );
  INV_X1 U7084 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7679) );
  NAND2_X1 U7085 ( .A1(n5740), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5566) );
  INV_X1 U7086 ( .A(n5974), .ZN(n5573) );
  INV_X1 U7087 ( .A(SI_0_), .ZN(n5570) );
  INV_X1 U7088 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5569) );
  OAI21_X1 U7089 ( .B1(n6814), .B2(n5570), .A(n5569), .ZN(n5572) );
  AND2_X1 U7090 ( .A1(n5572), .A2(n5571), .ZN(n9634) );
  AND2_X1 U7091 ( .A1(n5573), .A2(n7673), .ZN(n7545) );
  INV_X1 U7092 ( .A(n7673), .ZN(n6935) );
  AND2_X1 U7093 ( .A1(n6935), .A2(n5974), .ZN(n5893) );
  OR2_X1 U7094 ( .A1(n7545), .A2(n5893), .ZN(n7676) );
  NAND2_X1 U7095 ( .A1(n5740), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5580) );
  INV_X1 U7096 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5574) );
  OR2_X1 U7097 ( .A1(n5741), .A2(n5574), .ZN(n5579) );
  INV_X1 U7098 ( .A(n5654), .ZN(n5576) );
  INV_X1 U7099 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7259) );
  INV_X1 U7100 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9233) );
  NAND2_X1 U7101 ( .A1(n7259), .A2(n9233), .ZN(n5575) );
  NAND2_X1 U7102 ( .A1(n5576), .A2(n5575), .ZN(n9784) );
  OR2_X1 U7103 ( .A1(n5637), .A2(n9784), .ZN(n5578) );
  INV_X1 U7104 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6888) );
  OR2_X1 U7105 ( .A1(n5743), .A2(n6888), .ZN(n5577) );
  NAND4_X1 U7106 ( .A1(n5580), .A2(n5579), .A3(n5578), .A4(n5577), .ZN(n9195)
         );
  INV_X1 U7107 ( .A(n9195), .ZN(n7526) );
  OR2_X1 U7108 ( .A1(n5582), .A2(n5421), .ZN(n5583) );
  NAND2_X1 U7109 ( .A1(n5626), .A2(n5583), .ZN(n5646) );
  XNOR2_X1 U7110 ( .A(n5646), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6889) );
  XNOR2_X1 U7111 ( .A(n5584), .B(n5585), .ZN(n6823) );
  OR2_X1 U7112 ( .A1(n4517), .A2(n6824), .ZN(n5586) );
  NAND2_X1 U7113 ( .A1(n7526), .A2(n9789), .ZN(n5757) );
  NAND2_X1 U7114 ( .A1(n4839), .A2(n9195), .ZN(n5756) );
  NAND2_X1 U7115 ( .A1(n5757), .A2(n5756), .ZN(n9791) );
  NOR3_X1 U7116 ( .A1(n7676), .A2(n9791), .A3(n6186), .ZN(n5645) );
  NAND2_X1 U7117 ( .A1(n5740), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5596) );
  AND2_X1 U7118 ( .A1(n5653), .A2(n5589), .ZN(n5590) );
  OR2_X1 U7119 ( .A1(n5590), .A2(n5696), .ZN(n9769) );
  OR2_X1 U7120 ( .A1(n5637), .A2(n9769), .ZN(n5595) );
  INV_X1 U7121 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6890) );
  OR2_X1 U7122 ( .A1(n5591), .A2(n6890), .ZN(n5594) );
  INV_X1 U7123 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5592) );
  OR2_X1 U7124 ( .A1(n5741), .A2(n5592), .ZN(n5593) );
  NAND4_X1 U7125 ( .A1(n5596), .A2(n5595), .A3(n5594), .A4(n5593), .ZN(n9194)
         );
  INV_X1 U7126 ( .A(n9194), .ZN(n7532) );
  NAND2_X1 U7127 ( .A1(n5598), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5599) );
  MUX2_X1 U7128 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5599), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5600) );
  AND2_X1 U7129 ( .A1(n5597), .A2(n5600), .ZN(n6907) );
  INV_X1 U7130 ( .A(n6907), .ZN(n6875) );
  XNOR2_X1 U7131 ( .A(n5602), .B(n5601), .ZN(n6331) );
  INV_X1 U7132 ( .A(n6331), .ZN(n6830) );
  OR2_X1 U7133 ( .A1(n5633), .A2(n6830), .ZN(n5604) );
  INV_X1 U7134 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6831) );
  OR2_X1 U7135 ( .A1(n4517), .A2(n6831), .ZN(n5603) );
  OAI211_X1 U7136 ( .C1(n6845), .C2(n6875), .A(n5604), .B(n5603), .ZN(n9771)
         );
  NAND2_X1 U7137 ( .A1(n7532), .A2(n9771), .ZN(n5758) );
  INV_X1 U7138 ( .A(n9771), .ZN(n9867) );
  NAND2_X1 U7139 ( .A1(n9867), .A2(n9194), .ZN(n9761) );
  NAND2_X1 U7140 ( .A1(n5758), .A2(n9761), .ZN(n9772) );
  INV_X1 U7141 ( .A(n9772), .ZN(n5644) );
  NAND2_X1 U7142 ( .A1(n5740), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5609) );
  INV_X1 U7143 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9199) );
  INV_X1 U7144 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5605) );
  NAND4_X2 U7145 ( .A1(n5609), .A2(n5608), .A3(n5607), .A4(n5606), .ZN(n5979)
         );
  XNOR2_X1 U7146 ( .A(n5611), .B(n5610), .ZN(n6815) );
  OR2_X1 U7147 ( .A1(n5633), .A2(n6815), .ZN(n5613) );
  INV_X1 U7148 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5612) );
  INV_X1 U7149 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5615) );
  OR2_X1 U7150 ( .A1(n5741), .A2(n5615), .ZN(n5622) );
  INV_X1 U7151 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5616) );
  OR2_X1 U7152 ( .A1(n5617), .A2(n5616), .ZN(n5621) );
  INV_X1 U7153 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7476) );
  NAND2_X1 U7154 ( .A1(n5618), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5619) );
  XNOR2_X1 U7155 ( .A(n5624), .B(n5623), .ZN(n6818) );
  INV_X1 U7156 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7157 ( .A1(n5626), .A2(n5625), .ZN(n5628) );
  OAI21_X1 U7158 ( .B1(n5626), .B2(n5625), .A(n5628), .ZN(n6885) );
  NOR2_X1 U7159 ( .A1(n5627), .A2(n7518), .ZN(n5643) );
  NAND2_X1 U7160 ( .A1(n5628), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5630) );
  INV_X1 U7161 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5629) );
  XNOR2_X1 U7162 ( .A(n5632), .B(n5631), .ZN(n6820) );
  OR2_X1 U7163 ( .A1(n5633), .A2(n6820), .ZN(n5636) );
  OR2_X1 U7164 ( .A1(n4516), .A2(n6821), .ZN(n5635) );
  OAI211_X1 U7165 ( .C1(n6845), .C2(n9214), .A(n5636), .B(n5635), .ZN(n7650)
         );
  NAND2_X1 U7166 ( .A1(n5740), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5641) );
  OR2_X1 U7167 ( .A1(n5637), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5640) );
  INV_X1 U7168 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6887) );
  OR2_X1 U7169 ( .A1(n5743), .A2(n6887), .ZN(n5639) );
  OR2_X1 U7170 ( .A1(n5741), .A2(n7648), .ZN(n5638) );
  NAND4_X1 U7171 ( .A1(n5641), .A2(n5640), .A3(n5639), .A4(n5638), .ZN(n9196)
         );
  XNOR2_X1 U7172 ( .A(n5754), .B(n9196), .ZN(n7645) );
  INV_X1 U7173 ( .A(n7645), .ZN(n5642) );
  NAND4_X1 U7174 ( .A1(n5645), .A2(n5644), .A3(n5643), .A4(n5642), .ZN(n5659)
         );
  OAI21_X1 U7175 ( .B1(n5646), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5647) );
  XNOR2_X1 U7176 ( .A(n5647), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9252) );
  INV_X1 U7177 ( .A(n9252), .ZN(n6825) );
  XNOR2_X1 U7178 ( .A(n5649), .B(n5648), .ZN(n6827) );
  OR2_X1 U7179 ( .A1(n5633), .A2(n6827), .ZN(n5651) );
  OR2_X1 U7180 ( .A1(n4517), .A2(n6826), .ZN(n5650) );
  OAI211_X1 U7181 ( .C1(n6845), .C2(n6825), .A(n5651), .B(n5650), .ZN(n9859)
         );
  INV_X1 U7182 ( .A(n9859), .ZN(n7692) );
  NAND2_X1 U7183 ( .A1(n5618), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5658) );
  INV_X1 U7184 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7689) );
  OR2_X1 U7185 ( .A1(n5741), .A2(n7689), .ZN(n5657) );
  INV_X1 U7186 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5652) );
  OR2_X1 U7187 ( .A1(n5617), .A2(n5652), .ZN(n5656) );
  OAI21_X1 U7188 ( .B1(n5654), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5653), .ZN(
        n7691) );
  OR2_X1 U7189 ( .A1(n5637), .A2(n7691), .ZN(n5655) );
  NAND4_X1 U7190 ( .A1(n5658), .A2(n5657), .A3(n5656), .A4(n5655), .ZN(n9695)
         );
  XNOR2_X1 U7191 ( .A(n7692), .B(n9695), .ZN(n7684) );
  NOR2_X1 U7192 ( .A1(n5659), .A2(n7684), .ZN(n5708) );
  XNOR2_X1 U7193 ( .A(n5660), .B(n5119), .ZN(n6849) );
  NAND2_X1 U7194 ( .A1(n6849), .A2(n5737), .ZN(n5665) );
  OR2_X1 U7195 ( .A1(n5661), .A2(n5421), .ZN(n5682) );
  INV_X1 U7196 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7197 ( .A1(n5682), .A2(n5662), .ZN(n5684) );
  NAND2_X1 U7198 ( .A1(n5684), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5663) );
  XNOR2_X1 U7199 ( .A(n5663), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9269) );
  AOI22_X1 U7200 ( .A1(n5686), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5692), .B2(
        n9269), .ZN(n5664) );
  NAND2_X1 U7201 ( .A1(n5740), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5672) );
  INV_X1 U7202 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5666) );
  OR2_X1 U7203 ( .A1(n5743), .A2(n5666), .ZN(n5671) );
  OR2_X1 U7204 ( .A1(n5676), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5667) );
  NAND2_X1 U7205 ( .A1(n5668), .A2(n5667), .ZN(n9103) );
  OR2_X1 U7206 ( .A1(n5637), .A2(n9103), .ZN(n5670) );
  INV_X1 U7207 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7721) );
  OR2_X1 U7208 ( .A1(n5741), .A2(n7721), .ZN(n5669) );
  NAND4_X1 U7209 ( .A1(n5672), .A2(n5671), .A3(n5670), .A4(n5669), .ZN(n9192)
         );
  INV_X1 U7210 ( .A(n9192), .ZN(n5704) );
  OR2_X1 U7211 ( .A1(n9883), .A2(n5704), .ZN(n7707) );
  NAND2_X1 U7212 ( .A1(n5673), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5680) );
  INV_X1 U7213 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5674) );
  OR2_X1 U7214 ( .A1(n5617), .A2(n5674), .ZN(n5679) );
  NOR2_X1 U7215 ( .A1(n5698), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5675) );
  OR2_X1 U7216 ( .A1(n5676), .A2(n5675), .ZN(n9751) );
  OR2_X1 U7217 ( .A1(n5637), .A2(n9751), .ZN(n5678) );
  INV_X1 U7218 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6892) );
  OR2_X1 U7219 ( .A1(n5743), .A2(n6892), .ZN(n5677) );
  NAND4_X1 U7220 ( .A1(n5680), .A2(n5679), .A3(n5678), .A4(n5677), .ZN(n9193)
         );
  INV_X1 U7221 ( .A(n9193), .ZN(n5705) );
  NAND2_X1 U7222 ( .A1(n6836), .A2(n5737), .ZN(n5688) );
  INV_X1 U7223 ( .A(n5682), .ZN(n5683) );
  NAND2_X1 U7224 ( .A1(n5683), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5685) );
  AOI22_X1 U7225 ( .A1(n5686), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5692), .B2(
        n6968), .ZN(n5687) );
  NAND2_X1 U7226 ( .A1(n5688), .A2(n5687), .ZN(n9755) );
  OR2_X1 U7227 ( .A1(n5705), .A2(n9755), .ZN(n7710) );
  INV_X1 U7228 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6833) );
  XNOR2_X1 U7229 ( .A(n5690), .B(n5689), .ZN(n6832) );
  NAND2_X1 U7230 ( .A1(n6832), .A2(n5737), .ZN(n5694) );
  NAND2_X1 U7231 ( .A1(n5597), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5691) );
  XNOR2_X1 U7232 ( .A(n5691), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6919) );
  NAND2_X1 U7233 ( .A1(n5692), .A2(n6919), .ZN(n5693) );
  OAI211_X1 U7234 ( .C1(n4516), .C2(n6833), .A(n5694), .B(n5693), .ZN(n7539)
         );
  NAND2_X1 U7235 ( .A1(n5740), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5702) );
  INV_X1 U7236 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7540) );
  OR2_X1 U7237 ( .A1(n5741), .A2(n7540), .ZN(n5701) );
  NOR2_X1 U7238 ( .A1(n5696), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5697) );
  OR2_X1 U7239 ( .A1(n5698), .A2(n5697), .ZN(n7733) );
  OR2_X1 U7240 ( .A1(n5637), .A2(n7733), .ZN(n5700) );
  INV_X1 U7241 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6891) );
  OR2_X1 U7242 ( .A1(n5743), .A2(n6891), .ZN(n5699) );
  NAND4_X1 U7243 ( .A1(n5702), .A2(n5701), .A3(n5700), .A4(n5699), .ZN(n9697)
         );
  NAND2_X1 U7244 ( .A1(n9873), .A2(n9697), .ZN(n5703) );
  AND2_X1 U7245 ( .A1(n7710), .A2(n5703), .ZN(n5805) );
  AND2_X1 U7246 ( .A1(n7707), .A2(n5805), .ZN(n5761) );
  NAND2_X1 U7247 ( .A1(n9883), .A2(n5704), .ZN(n7706) );
  NAND2_X1 U7248 ( .A1(n9755), .A2(n5705), .ZN(n7709) );
  INV_X1 U7249 ( .A(n9697), .ZN(n7715) );
  NAND2_X1 U7250 ( .A1(n7715), .A2(n7539), .ZN(n9745) );
  NAND2_X1 U7251 ( .A1(n7709), .A2(n9745), .ZN(n5804) );
  NAND2_X1 U7252 ( .A1(n5804), .A2(n7710), .ZN(n5706) );
  NAND2_X1 U7253 ( .A1(n7706), .A2(n5706), .ZN(n5759) );
  INV_X1 U7254 ( .A(n5759), .ZN(n5707) );
  NAND4_X1 U7255 ( .A1(n5763), .A2(n5708), .A3(n5761), .A4(n5707), .ZN(n5709)
         );
  NOR2_X1 U7256 ( .A1(n4575), .A2(n5709), .ZN(n5712) );
  OR2_X1 U7257 ( .A1(n9051), .A2(n5710), .ZN(n5818) );
  AND2_X1 U7258 ( .A1(n5818), .A2(n7812), .ZN(n5902) );
  NAND4_X1 U7259 ( .A1(n5906), .A2(n5905), .A3(n5712), .A4(n5902), .ZN(n5713)
         );
  OR3_X1 U7260 ( .A1(n9597), .A2(n7956), .A3(n5713), .ZN(n5714) );
  NOR2_X1 U7261 ( .A1(n9655), .A2(n5714), .ZN(n5715) );
  NAND4_X1 U7262 ( .A1(n9479), .A2(n9488), .A3(n9505), .A4(n5715), .ZN(n5716)
         );
  OR3_X1 U7263 ( .A1(n9456), .A2(n9449), .A3(n5716), .ZN(n5717) );
  NOR3_X1 U7264 ( .A1(n9416), .A2(n9427), .A3(n5717), .ZN(n5718) );
  NAND4_X1 U7265 ( .A1(n8088), .A2(n9394), .A3(n4802), .A4(n5718), .ZN(n5719)
         );
  OR4_X1 U7266 ( .A1(n8070), .A2(n9361), .A3(n9375), .A4(n5719), .ZN(n5750) );
  INV_X1 U7267 ( .A(n5720), .ZN(n5721) );
  MUX2_X1 U7268 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6814), .Z(n5725) );
  XNOR2_X1 U7269 ( .A(n5725), .B(SI_30_), .ZN(n5735) );
  INV_X1 U7270 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10265) );
  INV_X1 U7271 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n10100) );
  MUX2_X1 U7272 ( .A(n10265), .B(n10100), .S(n6814), .Z(n5726) );
  XNOR2_X1 U7273 ( .A(n5726), .B(SI_31_), .ZN(n5727) );
  NAND2_X1 U7274 ( .A1(n9626), .A2(n5737), .ZN(n5730) );
  OR2_X1 U7275 ( .A1(n4517), .A2(n10265), .ZN(n5729) );
  NAND2_X1 U7276 ( .A1(n5695), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5734) );
  INV_X1 U7277 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n5731) );
  OR2_X1 U7278 ( .A1(n5743), .A2(n5731), .ZN(n5733) );
  INV_X1 U7279 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9348) );
  OR2_X1 U7280 ( .A1(n5741), .A2(n9348), .ZN(n5732) );
  NOR2_X1 U7281 ( .A1(n9524), .A2(n9347), .ZN(n5938) );
  INV_X1 U7282 ( .A(n5938), .ZN(n5748) );
  NAND2_X1 U7283 ( .A1(n8248), .A2(n5737), .ZN(n5739) );
  INV_X1 U7284 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9630) );
  OR2_X1 U7285 ( .A1(n4516), .A2(n9630), .ZN(n5738) );
  NAND2_X1 U7286 ( .A1(n5695), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5746) );
  INV_X1 U7287 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9355) );
  OR2_X1 U7288 ( .A1(n5741), .A2(n9355), .ZN(n5745) );
  INV_X1 U7289 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n5742) );
  OR2_X1 U7290 ( .A1(n5743), .A2(n5742), .ZN(n5744) );
  AND2_X1 U7291 ( .A1(n9357), .A2(n8041), .ZN(n5790) );
  NOR2_X1 U7292 ( .A1(n9357), .A2(n8041), .ZN(n5922) );
  NOR2_X1 U7293 ( .A1(n5790), .A2(n5922), .ZN(n5747) );
  NAND2_X1 U7294 ( .A1(n5748), .A2(n5747), .ZN(n5749) );
  INV_X1 U7295 ( .A(n5979), .ZN(n5892) );
  NAND2_X1 U7296 ( .A1(n5892), .A2(n9835), .ZN(n5751) );
  NAND2_X1 U7297 ( .A1(n5752), .A2(n5751), .ZN(n7479) );
  INV_X1 U7298 ( .A(n7518), .ZN(n7481) );
  NAND2_X1 U7299 ( .A1(n7479), .A2(n7481), .ZN(n7480) );
  INV_X1 U7300 ( .A(n9197), .ZN(n7520) );
  NAND2_X1 U7301 ( .A1(n7520), .A2(n7113), .ZN(n5753) );
  NAND2_X1 U7302 ( .A1(n7480), .A2(n5753), .ZN(n7641) );
  NOR2_X1 U7303 ( .A1(n5754), .A2(n9196), .ZN(n5755) );
  NAND2_X1 U7304 ( .A1(n5754), .A2(n9196), .ZN(n5891) );
  INV_X1 U7305 ( .A(n5756), .ZN(n5897) );
  NAND2_X1 U7306 ( .A1(n7692), .A2(n9695), .ZN(n5895) );
  INV_X1 U7307 ( .A(n9695), .ZN(n7529) );
  INV_X1 U7308 ( .A(n9763), .ZN(n5760) );
  NAND2_X1 U7309 ( .A1(n5760), .A2(n4562), .ZN(n7750) );
  NAND2_X1 U7310 ( .A1(n5761), .A2(n9761), .ZN(n5762) );
  NAND2_X1 U7311 ( .A1(n5762), .A2(n4562), .ZN(n7749) );
  AND2_X1 U7312 ( .A1(n5763), .A2(n7749), .ZN(n5764) );
  NAND2_X1 U7313 ( .A1(n7750), .A2(n5764), .ZN(n7780) );
  NAND2_X1 U7314 ( .A1(n7812), .A2(n5813), .ZN(n7790) );
  INV_X1 U7315 ( .A(n7779), .ZN(n5765) );
  NOR2_X1 U7316 ( .A1(n7790), .A2(n5765), .ZN(n5766) );
  NAND2_X1 U7317 ( .A1(n7815), .A2(n7812), .ZN(n5767) );
  NAND2_X1 U7318 ( .A1(n5767), .A2(n7832), .ZN(n7819) );
  XNOR2_X1 U7319 ( .A(n9125), .B(n5768), .ZN(n7874) );
  INV_X1 U7320 ( .A(n7947), .ZN(n5815) );
  NOR2_X1 U7321 ( .A1(n7956), .A2(n5815), .ZN(n5769) );
  NAND2_X1 U7322 ( .A1(n9595), .A2(n5769), .ZN(n5770) );
  NAND2_X1 U7323 ( .A1(n5770), .A2(n5820), .ZN(n9648) );
  INV_X1 U7324 ( .A(n9655), .ZN(n9649) );
  NAND2_X1 U7325 ( .A1(n9648), .A2(n9649), .ZN(n9647) );
  INV_X1 U7326 ( .A(n5915), .ZN(n5771) );
  NAND2_X1 U7327 ( .A1(n8037), .A2(n8036), .ZN(n5869) );
  NAND2_X1 U7328 ( .A1(n5870), .A2(n5801), .ZN(n5785) );
  INV_X1 U7329 ( .A(n9179), .ZN(n8057) );
  OR2_X1 U7330 ( .A1(n9567), .A2(n8057), .ZN(n5772) );
  NAND2_X1 U7331 ( .A1(n5854), .A2(n5772), .ZN(n5850) );
  NAND2_X1 U7332 ( .A1(n5850), .A2(n5851), .ZN(n5773) );
  NAND2_X1 U7333 ( .A1(n9392), .A2(n5773), .ZN(n5774) );
  NAND2_X1 U7334 ( .A1(n5774), .A2(n5855), .ZN(n5775) );
  AND2_X1 U7335 ( .A1(n5800), .A2(n5775), .ZN(n5783) );
  AND2_X1 U7336 ( .A1(n5851), .A2(n4585), .ZN(n5852) );
  NAND2_X1 U7337 ( .A1(n8032), .A2(n5834), .ZN(n5845) );
  NAND2_X1 U7338 ( .A1(n5845), .A2(n5847), .ZN(n5776) );
  NAND3_X1 U7339 ( .A1(n5855), .A2(n5852), .A3(n5776), .ZN(n5778) );
  INV_X1 U7340 ( .A(n8033), .ZN(n5777) );
  AOI21_X1 U7341 ( .B1(n5783), .B2(n5778), .A(n5777), .ZN(n5779) );
  NOR2_X1 U7342 ( .A1(n5785), .A2(n5779), .ZN(n5780) );
  NOR2_X1 U7343 ( .A1(n5869), .A2(n5780), .ZN(n5786) );
  INV_X1 U7344 ( .A(n5786), .ZN(n5782) );
  INV_X1 U7345 ( .A(n8035), .ZN(n5781) );
  INV_X1 U7346 ( .A(n5788), .ZN(n5916) );
  INV_X1 U7347 ( .A(n5783), .ZN(n5784) );
  NAND2_X1 U7348 ( .A1(n5847), .A2(n8031), .ZN(n5846) );
  NOR2_X1 U7349 ( .A1(n5784), .A2(n5846), .ZN(n5789) );
  AOI21_X1 U7350 ( .B1(n5786), .B2(n5785), .A(n8038), .ZN(n5787) );
  AOI21_X1 U7351 ( .B1(n9460), .B2(n5916), .A(n5887), .ZN(n5793) );
  INV_X1 U7352 ( .A(n5790), .ZN(n5791) );
  NAND2_X1 U7353 ( .A1(n5791), .A2(n5874), .ZN(n5919) );
  INV_X1 U7354 ( .A(n5922), .ZN(n5792) );
  OAI22_X1 U7355 ( .A1(n5793), .A2(n5919), .B1(n9347), .B2(n5792), .ZN(n5798)
         );
  INV_X1 U7356 ( .A(n9347), .ZN(n9171) );
  OAI21_X1 U7357 ( .B1(n9171), .B2(n9357), .A(n5877), .ZN(n5797) );
  NAND2_X1 U7358 ( .A1(n5795), .A2(n5794), .ZN(n5796) );
  AOI21_X1 U7359 ( .B1(n5798), .B2(n5797), .A(n6178), .ZN(n5799) );
  OAI21_X1 U7360 ( .B1(n5924), .B2(n5799), .A(n4581), .ZN(n5882) );
  INV_X1 U7361 ( .A(n5883), .ZN(n5959) );
  NAND2_X1 U7362 ( .A1(n8035), .A2(n8033), .ZN(n5863) );
  OR2_X1 U7363 ( .A1(n5863), .A2(n5800), .ZN(n5802) );
  NAND2_X1 U7364 ( .A1(n5802), .A2(n5801), .ZN(n5861) );
  INV_X1 U7365 ( .A(n5870), .ZN(n5803) );
  OR2_X1 U7366 ( .A1(n5861), .A2(n5803), .ZN(n5862) );
  INV_X1 U7367 ( .A(n6185), .ZN(n5872) );
  NOR2_X1 U7368 ( .A1(n5862), .A2(n5872), .ZN(n5859) );
  NOR3_X1 U7369 ( .A1(n5869), .A2(n6185), .A3(n5863), .ZN(n5858) );
  XNOR2_X1 U7370 ( .A(n7715), .B(n7539), .ZN(n7713) );
  OAI211_X1 U7371 ( .C1(n7708), .C2(n5804), .A(n7707), .B(n7710), .ZN(n5809)
         );
  INV_X1 U7372 ( .A(n7534), .ZN(n5806) );
  OAI21_X1 U7373 ( .B1(n5806), .B2(n7713), .A(n5805), .ZN(n5807) );
  NAND2_X1 U7374 ( .A1(n5807), .A2(n7709), .ZN(n5808) );
  MUX2_X1 U7375 ( .A(n5809), .B(n5808), .S(n6185), .Z(n5811) );
  INV_X1 U7376 ( .A(n7706), .ZN(n5810) );
  NOR2_X1 U7377 ( .A1(n5811), .A2(n5810), .ZN(n5817) );
  OAI21_X1 U7378 ( .B1(n5817), .B2(n5810), .A(n5900), .ZN(n5812) );
  INV_X1 U7379 ( .A(n5906), .ZN(n5814) );
  NAND2_X1 U7380 ( .A1(n5828), .A2(n5823), .ZN(n5888) );
  NOR2_X1 U7381 ( .A1(n5888), .A2(n5815), .ZN(n5907) );
  INV_X1 U7382 ( .A(n7707), .ZN(n5816) );
  NAND2_X1 U7383 ( .A1(n9506), .A2(n5820), .ZN(n5829) );
  INV_X1 U7384 ( .A(n5821), .ZN(n5822) );
  NOR2_X1 U7385 ( .A1(n5829), .A2(n5822), .ZN(n5912) );
  INV_X1 U7386 ( .A(n9506), .ZN(n5889) );
  OAI21_X1 U7387 ( .B1(n5889), .B2(n5823), .A(n5828), .ZN(n5824) );
  AOI21_X1 U7388 ( .B1(n5825), .B2(n5912), .A(n5824), .ZN(n5826) );
  MUX2_X1 U7389 ( .A(n5827), .B(n5826), .S(n6185), .Z(n5831) );
  NAND3_X1 U7390 ( .A1(n5829), .A2(n5872), .A3(n5828), .ZN(n5830) );
  AOI21_X1 U7391 ( .B1(n5831), .B2(n5830), .A(n9511), .ZN(n5836) );
  NAND2_X1 U7392 ( .A1(n5838), .A2(n5832), .ZN(n5913) );
  NOR2_X1 U7393 ( .A1(n5836), .A2(n5913), .ZN(n5835) );
  NAND2_X1 U7394 ( .A1(n5833), .A2(n5837), .ZN(n5917) );
  OAI211_X1 U7395 ( .C1(n5835), .C2(n5917), .A(n5834), .B(n5915), .ZN(n5843)
         );
  INV_X1 U7396 ( .A(n5836), .ZN(n5841) );
  MUX2_X1 U7397 ( .A(n5843), .B(n5842), .S(n6185), .Z(n5844) );
  MUX2_X1 U7398 ( .A(n5846), .B(n5845), .S(n6185), .Z(n5849) );
  MUX2_X1 U7399 ( .A(n8032), .B(n5847), .S(n6185), .Z(n5848) );
  INV_X1 U7400 ( .A(n5851), .ZN(n9409) );
  OAI211_X1 U7401 ( .C1(n6185), .C2(n5854), .A(n5853), .B(n4802), .ZN(n5857)
         );
  MUX2_X1 U7402 ( .A(n5855), .B(n9392), .S(n6185), .Z(n5856) );
  OAI211_X1 U7403 ( .C1(n5859), .C2(n5858), .A(n5857), .B(n5856), .ZN(n5868)
         );
  INV_X1 U7404 ( .A(n5869), .ZN(n5860) );
  NAND3_X1 U7405 ( .A1(n5861), .A2(n5860), .A3(n5872), .ZN(n5867) );
  INV_X1 U7406 ( .A(n5862), .ZN(n5864) );
  NAND3_X1 U7407 ( .A1(n5864), .A2(n6185), .A3(n5863), .ZN(n5866) );
  NAND2_X1 U7408 ( .A1(n5869), .A2(n6185), .ZN(n5865) );
  NAND4_X1 U7409 ( .A1(n5868), .A2(n5867), .A3(n5866), .A4(n5865), .ZN(n5873)
         );
  OAI21_X1 U7410 ( .B1(n5870), .B2(n5869), .A(n4783), .ZN(n5871) );
  MUX2_X1 U7411 ( .A(n5875), .B(n5874), .S(n6185), .Z(n5876) );
  AOI21_X1 U7412 ( .B1(n9171), .B2(n5878), .A(n5938), .ZN(n5879) );
  OR2_X1 U7413 ( .A1(n5884), .A2(n5421), .ZN(n5886) );
  INV_X1 U7414 ( .A(n7471), .ZN(n5957) );
  INV_X1 U7415 ( .A(n5887), .ZN(n5921) );
  INV_X1 U7416 ( .A(n5888), .ZN(n5890) );
  NOR2_X1 U7417 ( .A1(n5890), .A2(n5889), .ZN(n5911) );
  OAI21_X1 U7418 ( .B1(n5892), .B2(n9835), .A(n5891), .ZN(n5899) );
  INV_X1 U7419 ( .A(n5893), .ZN(n5894) );
  OAI211_X1 U7420 ( .C1(n7520), .C2(n7113), .A(n6186), .B(n5894), .ZN(n5898)
         );
  INV_X1 U7421 ( .A(n5895), .ZN(n5896) );
  NOR4_X1 U7422 ( .A1(n5899), .A2(n5898), .A3(n5897), .A4(n5896), .ZN(n5901)
         );
  OAI211_X1 U7423 ( .C1(n7750), .C2(n5901), .A(n5900), .B(n7749), .ZN(n5903)
         );
  AOI21_X1 U7424 ( .B1(n5903), .B2(n4599), .A(n4636), .ZN(n5909) );
  NAND2_X1 U7425 ( .A1(n5905), .A2(n5904), .ZN(n5908) );
  OAI211_X1 U7426 ( .C1(n5909), .C2(n5908), .A(n5907), .B(n5906), .ZN(n5910)
         );
  OAI21_X1 U7427 ( .B1(n5912), .B2(n5911), .A(n5910), .ZN(n5914) );
  AOI21_X1 U7428 ( .B1(n9489), .B2(n5914), .A(n5913), .ZN(n5918) );
  OAI211_X1 U7429 ( .C1(n5918), .C2(n5917), .A(n5916), .B(n5915), .ZN(n5920)
         );
  AOI21_X1 U7430 ( .B1(n5921), .B2(n5920), .A(n5919), .ZN(n5923) );
  NOR2_X1 U7431 ( .A1(n5923), .A2(n5922), .ZN(n5929) );
  OAI21_X1 U7432 ( .B1(n5926), .B2(n5957), .A(n5925), .ZN(n5927) );
  AOI22_X1 U7433 ( .A1(n5927), .A2(n4581), .B1(n5938), .B2(n7471), .ZN(n5928)
         );
  NOR2_X1 U7434 ( .A1(n5928), .A2(n8097), .ZN(n5936) );
  AOI211_X1 U7435 ( .C1(n5929), .C2(n4581), .A(n5938), .B(n6929), .ZN(n5935)
         );
  NAND2_X1 U7436 ( .A1(n5931), .A2(n5930), .ZN(n5932) );
  NAND2_X1 U7437 ( .A1(n5932), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5934) );
  OR2_X1 U7438 ( .A1(n6842), .A2(P1_U3086), .ZN(n7910) );
  NOR2_X1 U7439 ( .A1(n5936), .A2(n5127), .ZN(n5937) );
  OAI21_X1 U7440 ( .B1(n4581), .B2(n8097), .A(n5881), .ZN(n5940) );
  NAND2_X1 U7441 ( .A1(n5957), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7655) );
  NOR4_X1 U7442 ( .A1(n6842), .A2(n6931), .A3(n7778), .A4(n7655), .ZN(n5939)
         );
  OAI211_X1 U7443 ( .C1(n5748), .C2(n8097), .A(n5940), .B(n5939), .ZN(n5954)
         );
  OR2_X1 U7444 ( .A1(n6929), .A2(n6178), .ZN(n7675) );
  NAND2_X1 U7445 ( .A1(n5946), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5947) );
  OR2_X1 U7446 ( .A1(n5949), .A2(n4511), .ZN(n9227) );
  NOR3_X1 U7447 ( .A1(n7675), .A2(n9833), .A3(n9227), .ZN(n5952) );
  OAI21_X1 U7448 ( .B1(n7910), .B2(n6931), .A(P1_B_REG_SCAN_IN), .ZN(n5951) );
  OR2_X1 U7449 ( .A1(n5952), .A2(n5951), .ZN(n5953) );
  NAND3_X1 U7450 ( .A1(n5955), .A2(n5954), .A3(n5953), .ZN(P1_U3242) );
  NAND2_X1 U7451 ( .A1(n6186), .A2(n5957), .ZN(n6932) );
  NAND2_X1 U7452 ( .A1(n4518), .A2(n7113), .ZN(n5962) );
  AND2_X1 U7453 ( .A1(n6186), .A2(n7471), .ZN(n7467) );
  NAND2_X1 U7454 ( .A1(n9197), .A2(n6043), .ZN(n5961) );
  NAND2_X1 U7455 ( .A1(n5962), .A2(n5961), .ZN(n5964) );
  XNOR2_X1 U7456 ( .A(n5964), .B(n5963), .ZN(n5967) );
  NAND2_X1 U7458 ( .A1(n9197), .A2(n8975), .ZN(n5966) );
  NAND2_X1 U7459 ( .A1(n7113), .A2(n6043), .ZN(n5965) );
  AND2_X1 U7460 ( .A1(n5966), .A2(n5965), .ZN(n5968) );
  NAND2_X1 U7461 ( .A1(n5967), .A2(n5968), .ZN(n5992) );
  INV_X1 U7462 ( .A(n5967), .ZN(n5970) );
  INV_X1 U7463 ( .A(n5968), .ZN(n5969) );
  NAND2_X1 U7464 ( .A1(n5970), .A2(n5969), .ZN(n5971) );
  NAND2_X1 U7465 ( .A1(n5992), .A2(n5971), .ZN(n7107) );
  INV_X1 U7466 ( .A(n7107), .ZN(n5991) );
  NAND2_X1 U7467 ( .A1(n5974), .A2(n6043), .ZN(n5973) );
  OR2_X1 U7468 ( .A1(n5960), .A2(n9710), .ZN(n5972) );
  NAND3_X1 U7469 ( .A1(n5977), .A2(n5973), .A3(n5972), .ZN(n7080) );
  INV_X1 U7470 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9230) );
  NAND2_X1 U7471 ( .A1(n5974), .A2(n5985), .ZN(n5976) );
  NAND2_X1 U7472 ( .A1(n7673), .A2(n6043), .ZN(n5975) );
  OAI211_X1 U7473 ( .C1(n5960), .C2(n9230), .A(n5976), .B(n5975), .ZN(n7079)
         );
  NAND2_X1 U7474 ( .A1(n7080), .A2(n7079), .ZN(n7078) );
  NAND2_X1 U7475 ( .A1(n5977), .A2(n5963), .ZN(n5978) );
  NAND2_X1 U7476 ( .A1(n7078), .A2(n5978), .ZN(n7101) );
  NAND2_X1 U7477 ( .A1(n5979), .A2(n6043), .ZN(n5982) );
  NAND2_X1 U7478 ( .A1(n4518), .A2(n5980), .ZN(n5981) );
  NAND2_X1 U7479 ( .A1(n5982), .A2(n5981), .ZN(n5984) );
  XNOR2_X1 U7480 ( .A(n5984), .B(n5983), .ZN(n7100) );
  NAND2_X1 U7481 ( .A1(n5979), .A2(n8975), .ZN(n5987) );
  NAND2_X1 U7482 ( .A1(n9835), .A2(n6043), .ZN(n5986) );
  NAND2_X1 U7483 ( .A1(n5987), .A2(n5986), .ZN(n7102) );
  OAI21_X1 U7484 ( .B1(n7101), .B2(n7100), .A(n7102), .ZN(n5989) );
  NAND2_X1 U7485 ( .A1(n7101), .A2(n7100), .ZN(n5988) );
  NAND2_X1 U7486 ( .A1(n5989), .A2(n5988), .ZN(n7110) );
  INV_X1 U7487 ( .A(n7110), .ZN(n5990) );
  NAND2_X1 U7488 ( .A1(n5991), .A2(n5990), .ZN(n7108) );
  NAND2_X1 U7489 ( .A1(n7108), .A2(n5992), .ZN(n7256) );
  NAND2_X1 U7490 ( .A1(n4518), .A2(n7650), .ZN(n5995) );
  NAND2_X1 U7491 ( .A1(n9196), .A2(n6043), .ZN(n5994) );
  NAND2_X1 U7492 ( .A1(n5995), .A2(n5994), .ZN(n5996) );
  XNOR2_X1 U7493 ( .A(n5996), .B(n5963), .ZN(n6004) );
  NAND2_X1 U7494 ( .A1(n9196), .A2(n8975), .ZN(n5998) );
  NAND2_X1 U7495 ( .A1(n7650), .A2(n6043), .ZN(n5997) );
  NAND2_X1 U7496 ( .A1(n5998), .A2(n5997), .ZN(n6002) );
  XNOR2_X1 U7497 ( .A(n6004), .B(n6002), .ZN(n7257) );
  NAND2_X1 U7498 ( .A1(n9195), .A2(n6043), .ZN(n5999) );
  NAND2_X1 U7499 ( .A1(n9195), .A2(n8975), .ZN(n6001) );
  NAND2_X1 U7500 ( .A1(n9789), .A2(n6043), .ZN(n6000) );
  NAND2_X1 U7501 ( .A1(n6001), .A2(n6000), .ZN(n6007) );
  INV_X1 U7502 ( .A(n6002), .ZN(n6003) );
  NAND2_X1 U7503 ( .A1(n6004), .A2(n6003), .ZN(n7354) );
  AND2_X1 U7504 ( .A1(n7356), .A2(n7354), .ZN(n6005) );
  NAND2_X1 U7505 ( .A1(n7255), .A2(n6005), .ZN(n7355) );
  INV_X1 U7506 ( .A(n6006), .ZN(n6008) );
  NAND2_X1 U7507 ( .A1(n6008), .A2(n6007), .ZN(n6009) );
  NAND2_X1 U7508 ( .A1(n7355), .A2(n6009), .ZN(n6015) );
  NAND2_X1 U7509 ( .A1(n8971), .A2(n9859), .ZN(n6011) );
  NAND2_X1 U7510 ( .A1(n9695), .A2(n6152), .ZN(n6010) );
  NAND2_X1 U7511 ( .A1(n6011), .A2(n6010), .ZN(n6012) );
  XNOR2_X1 U7512 ( .A(n6012), .B(n4514), .ZN(n6014) );
  NAND2_X1 U7513 ( .A1(n9695), .A2(n8975), .ZN(n6017) );
  NAND2_X1 U7514 ( .A1(n9859), .A2(n6043), .ZN(n6016) );
  AND2_X1 U7515 ( .A1(n6017), .A2(n6016), .ZN(n7513) );
  NAND2_X1 U7516 ( .A1(n7512), .A2(n9692), .ZN(n6028) );
  NAND2_X1 U7517 ( .A1(n8971), .A2(n9771), .ZN(n6019) );
  NAND2_X1 U7518 ( .A1(n9194), .A2(n6152), .ZN(n6018) );
  NAND2_X1 U7519 ( .A1(n6019), .A2(n6018), .ZN(n6020) );
  XNOR2_X1 U7520 ( .A(n6020), .B(n5963), .ZN(n6023) );
  NAND2_X1 U7521 ( .A1(n9194), .A2(n8975), .ZN(n6022) );
  NAND2_X1 U7522 ( .A1(n9771), .A2(n6152), .ZN(n6021) );
  AND2_X1 U7523 ( .A1(n6022), .A2(n6021), .ZN(n6024) );
  NAND2_X1 U7524 ( .A1(n6023), .A2(n6024), .ZN(n6029) );
  INV_X1 U7525 ( .A(n6023), .ZN(n6026) );
  INV_X1 U7526 ( .A(n6024), .ZN(n6025) );
  NAND2_X1 U7527 ( .A1(n6026), .A2(n6025), .ZN(n6027) );
  AND2_X1 U7528 ( .A1(n6029), .A2(n6027), .ZN(n9690) );
  NAND2_X1 U7529 ( .A1(n6028), .A2(n9690), .ZN(n9689) );
  NAND2_X1 U7530 ( .A1(n7539), .A2(n8971), .ZN(n6031) );
  NAND2_X1 U7531 ( .A1(n9697), .A2(n6152), .ZN(n6030) );
  NAND2_X1 U7532 ( .A1(n6031), .A2(n6030), .ZN(n6032) );
  XNOR2_X1 U7533 ( .A(n6032), .B(n5963), .ZN(n6048) );
  NAND2_X1 U7534 ( .A1(n7539), .A2(n6152), .ZN(n6034) );
  NAND2_X1 U7535 ( .A1(n9697), .A2(n8975), .ZN(n6033) );
  NAND2_X1 U7536 ( .A1(n6034), .A2(n6033), .ZN(n6046) );
  XNOR2_X1 U7537 ( .A(n6048), .B(n6046), .ZN(n7729) );
  NAND2_X1 U7538 ( .A1(n9755), .A2(n8971), .ZN(n6036) );
  NAND2_X1 U7539 ( .A1(n9193), .A2(n6152), .ZN(n6035) );
  NAND2_X1 U7540 ( .A1(n6036), .A2(n6035), .ZN(n6037) );
  XNOR2_X1 U7541 ( .A(n6037), .B(n4514), .ZN(n6045) );
  NAND2_X1 U7542 ( .A1(n9755), .A2(n6152), .ZN(n6039) );
  NAND2_X1 U7543 ( .A1(n9193), .A2(n8975), .ZN(n6038) );
  NAND2_X1 U7544 ( .A1(n6039), .A2(n6038), .ZN(n7840) );
  AND2_X1 U7545 ( .A1(n6045), .A2(n7840), .ZN(n6054) );
  NAND2_X1 U7546 ( .A1(n9883), .A2(n8971), .ZN(n6041) );
  NAND2_X1 U7547 ( .A1(n9192), .A2(n6152), .ZN(n6040) );
  NAND2_X1 U7548 ( .A1(n6041), .A2(n6040), .ZN(n6042) );
  XNOR2_X1 U7549 ( .A(n6042), .B(n4514), .ZN(n6057) );
  AND2_X1 U7550 ( .A1(n9192), .A2(n8975), .ZN(n6044) );
  AOI21_X1 U7551 ( .B1(n9883), .B2(n6152), .A(n6044), .ZN(n6055) );
  XNOR2_X1 U7552 ( .A(n6057), .B(n6055), .ZN(n9097) );
  INV_X1 U7553 ( .A(n6045), .ZN(n9094) );
  INV_X1 U7554 ( .A(n6046), .ZN(n6047) );
  NAND2_X1 U7555 ( .A1(n6048), .A2(n6047), .ZN(n7839) );
  NAND2_X1 U7556 ( .A1(n7839), .A2(n7840), .ZN(n6051) );
  INV_X1 U7557 ( .A(n7839), .ZN(n6050) );
  INV_X1 U7558 ( .A(n7840), .ZN(n6049) );
  AOI22_X1 U7559 ( .A1(n9094), .A2(n6051), .B1(n6050), .B2(n6049), .ZN(n6052)
         );
  AND2_X1 U7560 ( .A1(n9097), .A2(n6052), .ZN(n6053) );
  INV_X1 U7561 ( .A(n6055), .ZN(n6056) );
  NAND2_X1 U7562 ( .A1(n6057), .A2(n6056), .ZN(n6061) );
  NAND2_X1 U7563 ( .A1(n7787), .A2(n8971), .ZN(n6059) );
  NAND2_X1 U7564 ( .A1(n9191), .A2(n6152), .ZN(n6058) );
  NAND2_X1 U7565 ( .A1(n6059), .A2(n6058), .ZN(n6060) );
  XNOR2_X1 U7566 ( .A(n6060), .B(n5963), .ZN(n6062) );
  NAND2_X1 U7567 ( .A1(n9095), .A2(n5120), .ZN(n6068) );
  INV_X1 U7568 ( .A(n6062), .ZN(n6063) );
  NAND2_X1 U7569 ( .A1(n6064), .A2(n6063), .ZN(n6065) );
  INV_X1 U7570 ( .A(n7787), .ZN(n9892) );
  OAI22_X1 U7571 ( .A1(n9892), .A2(n6076), .B1(n6067), .B2(n6135), .ZN(n9637)
         );
  INV_X1 U7572 ( .A(n6068), .ZN(n6069) );
  NAND2_X1 U7573 ( .A1(n9897), .A2(n8971), .ZN(n6071) );
  NAND2_X1 U7574 ( .A1(n9190), .A2(n6152), .ZN(n6070) );
  NAND2_X1 U7575 ( .A1(n6071), .A2(n6070), .ZN(n6072) );
  XNOR2_X1 U7576 ( .A(n6072), .B(n5963), .ZN(n6075) );
  AND2_X1 U7577 ( .A1(n9190), .A2(n8975), .ZN(n6073) );
  AOI21_X1 U7578 ( .B1(n9897), .B2(n6152), .A(n6073), .ZN(n6074) );
  NOR2_X1 U7579 ( .A1(n6075), .A2(n6074), .ZN(n9140) );
  AND2_X1 U7580 ( .A1(n6075), .A2(n6074), .ZN(n9139) );
  NOR2_X2 U7581 ( .A1(n9138), .A2(n9139), .ZN(n9045) );
  INV_X2 U7582 ( .A(n6076), .ZN(n6152) );
  AOI22_X1 U7583 ( .A1(n9051), .A2(n6152), .B1(n8975), .B2(n9189), .ZN(n6080)
         );
  NAND2_X1 U7584 ( .A1(n9051), .A2(n8971), .ZN(n6078) );
  NAND2_X1 U7585 ( .A1(n9189), .A2(n6152), .ZN(n6077) );
  NAND2_X1 U7586 ( .A1(n6078), .A2(n6077), .ZN(n6079) );
  XNOR2_X1 U7587 ( .A(n6079), .B(n4514), .ZN(n6082) );
  XOR2_X1 U7588 ( .A(n6080), .B(n6082), .Z(n9044) );
  INV_X1 U7589 ( .A(n6080), .ZN(n6081) );
  OAI22_X1 U7590 ( .A1(n9045), .A2(n9044), .B1(n6082), .B2(n6081), .ZN(n9119)
         );
  NAND2_X1 U7591 ( .A1(n9125), .A2(n8971), .ZN(n6084) );
  NAND2_X1 U7592 ( .A1(n9188), .A2(n6152), .ZN(n6083) );
  NAND2_X1 U7593 ( .A1(n6084), .A2(n6083), .ZN(n6085) );
  XNOR2_X1 U7594 ( .A(n6085), .B(n4514), .ZN(n6086) );
  AOI22_X1 U7595 ( .A1(n9125), .A2(n6152), .B1(n8975), .B2(n9188), .ZN(n6087)
         );
  XNOR2_X1 U7596 ( .A(n6086), .B(n6087), .ZN(n9120) );
  INV_X1 U7597 ( .A(n6086), .ZN(n6088) );
  AOI22_X1 U7598 ( .A1(n9735), .A2(n8971), .B1(n6152), .B2(n9187), .ZN(n6089)
         );
  XOR2_X1 U7599 ( .A(n4514), .B(n6089), .Z(n8994) );
  AOI22_X1 U7600 ( .A1(n9735), .A2(n6152), .B1(n8975), .B2(n9187), .ZN(n8993)
         );
  NAND2_X1 U7601 ( .A1(n9168), .A2(n8971), .ZN(n6091) );
  NAND2_X1 U7602 ( .A1(n9186), .A2(n6152), .ZN(n6090) );
  NAND2_X1 U7603 ( .A1(n6091), .A2(n6090), .ZN(n6092) );
  XNOR2_X1 U7604 ( .A(n6092), .B(n4514), .ZN(n9161) );
  NAND2_X1 U7605 ( .A1(n9168), .A2(n6152), .ZN(n6094) );
  NAND2_X1 U7606 ( .A1(n9186), .A2(n8975), .ZN(n6093) );
  NAND2_X1 U7607 ( .A1(n6094), .A2(n6093), .ZN(n6095) );
  AND2_X1 U7608 ( .A1(n9161), .A2(n6095), .ZN(n6097) );
  INV_X1 U7609 ( .A(n9161), .ZN(n6096) );
  INV_X1 U7610 ( .A(n6095), .ZN(n9160) );
  AOI22_X1 U7611 ( .A1(n9654), .A2(n6152), .B1(n8975), .B2(n9185), .ZN(n6102)
         );
  NAND2_X1 U7612 ( .A1(n9654), .A2(n8971), .ZN(n6099) );
  NAND2_X1 U7613 ( .A1(n9185), .A2(n6152), .ZN(n6098) );
  NAND2_X1 U7614 ( .A1(n6099), .A2(n6098), .ZN(n6100) );
  XNOR2_X1 U7615 ( .A(n6100), .B(n4514), .ZN(n6104) );
  XOR2_X1 U7616 ( .A(n6102), .B(n6104), .Z(n9064) );
  INV_X1 U7617 ( .A(n9064), .ZN(n6101) );
  INV_X1 U7618 ( .A(n6102), .ZN(n6103) );
  NAND2_X1 U7619 ( .A1(n6106), .A2(n6105), .ZN(n9071) );
  NAND2_X1 U7620 ( .A1(n9521), .A2(n8971), .ZN(n6108) );
  NAND2_X1 U7621 ( .A1(n9184), .A2(n6152), .ZN(n6107) );
  NAND2_X1 U7622 ( .A1(n6108), .A2(n6107), .ZN(n6109) );
  XNOR2_X1 U7623 ( .A(n6109), .B(n4514), .ZN(n6110) );
  AOI22_X1 U7624 ( .A1(n9521), .A2(n6152), .B1(n8975), .B2(n9184), .ZN(n6111)
         );
  XNOR2_X1 U7625 ( .A(n6110), .B(n6111), .ZN(n9072) );
  INV_X1 U7626 ( .A(n6110), .ZN(n6112) );
  AOI22_X1 U7627 ( .A1(n9588), .A2(n8971), .B1(n6152), .B2(n9183), .ZN(n6114)
         );
  XNOR2_X1 U7628 ( .A(n6114), .B(n4514), .ZN(n6115) );
  AOI22_X1 U7629 ( .A1(n9588), .A2(n6152), .B1(n8975), .B2(n9183), .ZN(n9149)
         );
  INV_X1 U7630 ( .A(n9582), .ZN(n9478) );
  OAI22_X1 U7631 ( .A1(n9478), .A2(n6076), .B1(n8051), .B2(n6135), .ZN(n6120)
         );
  NAND2_X1 U7632 ( .A1(n9582), .A2(n8971), .ZN(n6117) );
  NAND2_X1 U7633 ( .A1(n9182), .A2(n6152), .ZN(n6116) );
  NAND2_X1 U7634 ( .A1(n6117), .A2(n6116), .ZN(n6118) );
  XNOR2_X1 U7635 ( .A(n6118), .B(n4514), .ZN(n6119) );
  XOR2_X1 U7636 ( .A(n6120), .B(n6119), .Z(n9014) );
  INV_X1 U7637 ( .A(n6119), .ZN(n6122) );
  INV_X1 U7638 ( .A(n6120), .ZN(n6121) );
  AOI22_X1 U7639 ( .A1(n9578), .A2(n8971), .B1(n6152), .B2(n9181), .ZN(n6123)
         );
  XOR2_X1 U7640 ( .A(n4514), .B(n6123), .Z(n9110) );
  OAI22_X1 U7641 ( .A1(n9470), .A2(n6076), .B1(n8053), .B2(n6135), .ZN(n9111)
         );
  NAND2_X1 U7642 ( .A1(n9109), .A2(n5114), .ZN(n6125) );
  NAND2_X1 U7643 ( .A1(n9110), .A2(n9111), .ZN(n6124) );
  AND2_X1 U7644 ( .A1(n9180), .A2(n8975), .ZN(n6126) );
  AOI21_X1 U7645 ( .B1(n9572), .B2(n6152), .A(n6126), .ZN(n6129) );
  AOI22_X1 U7646 ( .A1(n9572), .A2(n8971), .B1(n6152), .B2(n9180), .ZN(n6127)
         );
  XNOR2_X1 U7647 ( .A(n6127), .B(n4514), .ZN(n6128) );
  XOR2_X1 U7648 ( .A(n6129), .B(n6128), .Z(n9037) );
  INV_X1 U7649 ( .A(n6128), .ZN(n6131) );
  INV_X1 U7650 ( .A(n6129), .ZN(n6130) );
  AOI22_X1 U7651 ( .A1(n9567), .A2(n8971), .B1(n6152), .B2(n9179), .ZN(n6133)
         );
  OAI22_X1 U7652 ( .A1(n9435), .A2(n6076), .B1(n8057), .B2(n6135), .ZN(n9128)
         );
  AOI22_X1 U7653 ( .A1(n9563), .A2(n8971), .B1(n6152), .B2(n9178), .ZN(n6134)
         );
  XOR2_X1 U7654 ( .A(n4514), .B(n6134), .Z(n6137) );
  OAI22_X1 U7655 ( .A1(n9424), .A2(n6076), .B1(n8060), .B2(n6135), .ZN(n6136)
         );
  NOR2_X1 U7656 ( .A1(n6137), .A2(n6136), .ZN(n9080) );
  AOI21_X1 U7657 ( .B1(n6137), .B2(n6136), .A(n9080), .ZN(n9005) );
  NAND2_X1 U7658 ( .A1(n9557), .A2(n8971), .ZN(n6139) );
  NAND2_X1 U7659 ( .A1(n9177), .A2(n6152), .ZN(n6138) );
  NAND2_X1 U7660 ( .A1(n6139), .A2(n6138), .ZN(n6140) );
  XNOR2_X1 U7661 ( .A(n6140), .B(n5963), .ZN(n6142) );
  AND2_X1 U7662 ( .A1(n9177), .A2(n8975), .ZN(n6141) );
  AOI21_X1 U7663 ( .B1(n9557), .B2(n6152), .A(n6141), .ZN(n6143) );
  NAND2_X1 U7664 ( .A1(n6142), .A2(n6143), .ZN(n6148) );
  INV_X1 U7665 ( .A(n6142), .ZN(n6145) );
  INV_X1 U7666 ( .A(n6143), .ZN(n6144) );
  NAND2_X1 U7667 ( .A1(n6145), .A2(n6144), .ZN(n6146) );
  NAND2_X1 U7668 ( .A1(n6147), .A2(n9079), .ZN(n9082) );
  NAND2_X1 U7669 ( .A1(n9082), .A2(n6148), .ZN(n9054) );
  NAND2_X1 U7670 ( .A1(n9552), .A2(n8971), .ZN(n6150) );
  NAND2_X1 U7671 ( .A1(n9176), .A2(n6152), .ZN(n6149) );
  NAND2_X1 U7672 ( .A1(n6150), .A2(n6149), .ZN(n6151) );
  XNOR2_X1 U7673 ( .A(n6151), .B(n5983), .ZN(n6153) );
  AOI22_X1 U7674 ( .A1(n9552), .A2(n6152), .B1(n8975), .B2(n9176), .ZN(n6154)
         );
  XNOR2_X1 U7675 ( .A(n6153), .B(n6154), .ZN(n9055) );
  INV_X1 U7676 ( .A(n6153), .ZN(n6155) );
  NAND2_X1 U7677 ( .A1(n6155), .A2(n6154), .ZN(n6180) );
  NAND2_X1 U7678 ( .A1(n9546), .A2(n8971), .ZN(n6157) );
  NAND2_X1 U7679 ( .A1(n9175), .A2(n6152), .ZN(n6156) );
  NAND2_X1 U7680 ( .A1(n6157), .A2(n6156), .ZN(n6158) );
  XNOR2_X1 U7681 ( .A(n6158), .B(n5983), .ZN(n8970) );
  AND2_X1 U7682 ( .A1(n9175), .A2(n8975), .ZN(n6159) );
  AOI21_X1 U7683 ( .B1(n9546), .B2(n6152), .A(n6159), .ZN(n8968) );
  XNOR2_X1 U7684 ( .A(n8970), .B(n8968), .ZN(n6183) );
  NAND2_X1 U7685 ( .A1(n8002), .A2(P1_B_REG_SCAN_IN), .ZN(n6160) );
  MUX2_X1 U7686 ( .A(P1_B_REG_SCAN_IN), .B(n6160), .S(n7965), .Z(n6162) );
  INV_X1 U7687 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6165) );
  INV_X1 U7688 ( .A(n7965), .ZN(n6163) );
  NOR2_X1 U7689 ( .A1(n6161), .A2(n6163), .ZN(n6164) );
  INV_X1 U7690 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9832) );
  INV_X1 U7691 ( .A(n8002), .ZN(n6166) );
  NOR2_X1 U7692 ( .A1(n6161), .A2(n6166), .ZN(n6167) );
  NOR2_X1 U7693 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .ZN(
        n6171) );
  NOR4_X1 U7694 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_31__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6170) );
  NOR4_X1 U7695 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6169) );
  NOR4_X1 U7696 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6168) );
  NAND4_X1 U7697 ( .A1(n6171), .A2(n6170), .A3(n6169), .A4(n6168), .ZN(n6177)
         );
  NOR4_X1 U7698 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6175) );
  NOR4_X1 U7699 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6174) );
  NOR4_X1 U7700 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n6173) );
  NOR4_X1 U7701 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6172) );
  NAND4_X1 U7702 ( .A1(n6175), .A2(n6174), .A3(n6173), .A4(n6172), .ZN(n6176)
         );
  OAI21_X1 U7703 ( .B1(n6177), .B2(n6176), .A(n9800), .ZN(n6925) );
  NAND3_X1 U7704 ( .A1(n9620), .A2(n7463), .A3(n6925), .ZN(n6193) );
  OR2_X1 U7705 ( .A1(n6193), .A2(n9833), .ZN(n6189) );
  NAND2_X1 U7706 ( .A1(n9913), .A2(n6178), .ZN(n6179) );
  NAND2_X1 U7707 ( .A1(n6182), .A2(n6181), .ZN(n8986) );
  OR2_X1 U7708 ( .A1(n7674), .A2(n7471), .ZN(n7474) );
  NAND2_X1 U7709 ( .A1(n9174), .A2(n4509), .ZN(n6188) );
  INV_X1 U7710 ( .A(n5949), .ZN(n9226) );
  NAND2_X1 U7711 ( .A1(n9226), .A2(n6843), .ZN(n8040) );
  INV_X2 U7712 ( .A(n8040), .ZN(n9131) );
  NAND2_X1 U7713 ( .A1(n9176), .A2(n9131), .ZN(n6187) );
  NAND2_X1 U7714 ( .A1(n6188), .A2(n6187), .ZN(n8089) );
  INV_X1 U7715 ( .A(n6189), .ZN(n6191) );
  INV_X1 U7716 ( .A(n6929), .ZN(n6190) );
  NAND2_X1 U7717 ( .A1(n9898), .A2(n7655), .ZN(n6192) );
  NAND2_X1 U7718 ( .A1(n6193), .A2(n6192), .ZN(n6194) );
  NAND2_X1 U7719 ( .A1(n6929), .A2(n6843), .ZN(n6924) );
  NAND2_X1 U7720 ( .A1(n6194), .A2(n6924), .ZN(n7081) );
  NAND2_X1 U7721 ( .A1(n5960), .A2(n6842), .ZN(n6195) );
  OAI22_X1 U7722 ( .A1(n8082), .A2(n9708), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10122), .ZN(n6197) );
  AOI21_X1 U7723 ( .B1(n8089), .B2(n9702), .A(n6197), .ZN(n6198) );
  INV_X1 U7724 ( .A(n6198), .ZN(n6199) );
  AOI21_X1 U7725 ( .B1(n9546), .B2(n6200), .A(n6199), .ZN(n6201) );
  AND2_X2 U7726 ( .A1(n6314), .A2(n6204), .ZN(n6316) );
  NOR2_X1 U7727 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n6210) );
  NAND2_X1 U7728 ( .A1(n6424), .A2(n6225), .ZN(n6436) );
  INV_X1 U7729 ( .A(n6436), .ZN(n6213) );
  NOR2_X1 U7730 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6212) );
  NAND2_X1 U7731 ( .A1(n6214), .A2(n6224), .ZN(n6614) );
  NAND2_X1 U7732 ( .A1(n6216), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U7733 ( .A1(n8437), .A2(n8459), .ZN(n6635) );
  NOR2_X1 U7734 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n6222) );
  NOR2_X1 U7735 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n6221) );
  NOR2_X1 U7736 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6220) );
  NOR2_X1 U7737 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n6219) );
  NAND4_X1 U7738 ( .A1(n6222), .A2(n6221), .A3(n6220), .A4(n6219), .ZN(n6227)
         );
  NAND4_X1 U7739 ( .A1(n6225), .A2(n6424), .A3(n6224), .A4(n6223), .ZN(n6226)
         );
  NAND2_X1 U7740 ( .A1(n6368), .A2(n6229), .ZN(n6636) );
  NAND2_X1 U7741 ( .A1(n6636), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6228) );
  INV_X1 U7742 ( .A(n10041), .ZN(n9997) );
  INV_X1 U7743 ( .A(n6229), .ZN(n6233) );
  NOR2_X1 U7744 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n6231) );
  NAND4_X1 U7745 ( .A1(n6231), .A2(n6230), .A3(n6641), .A4(n6670), .ZN(n6232)
         );
  NOR2_X1 U7746 ( .A1(n6233), .A2(n6232), .ZN(n6234) );
  INV_X1 U7747 ( .A(n6240), .ZN(n6237) );
  NAND2_X1 U7748 ( .A1(n6237), .A2(n6236), .ZN(n8954) );
  XNOR2_X2 U7749 ( .A(n6239), .B(n6238), .ZN(n8101) );
  NAND2_X1 U7750 ( .A1(n6240), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6241) );
  NAND2_X2 U7751 ( .A1(n8101), .A2(n8028), .ZN(n6295) );
  INV_X1 U7752 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U7753 ( .A1(n6545), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6247) );
  INV_X1 U7754 ( .A(n8101), .ZN(n6243) );
  AND2_X2 U7755 ( .A1(n6243), .A2(n8028), .ZN(n6309) );
  NAND2_X1 U7756 ( .A1(n6309), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6246) );
  INV_X1 U7757 ( .A(n8028), .ZN(n6244) );
  NAND2_X1 U7758 ( .A1(n6280), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7759 ( .A1(n6814), .A2(SI_0_), .ZN(n6249) );
  XNOR2_X1 U7760 ( .A(n6249), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8967) );
  MUX2_X1 U7761 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8967), .S(n6266), .Z(n7369) );
  INV_X1 U7762 ( .A(n7369), .ZN(n7119) );
  INV_X1 U7763 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6255) );
  OR2_X1 U7764 ( .A1(n6256), .A2(n6255), .ZN(n6259) );
  NAND2_X1 U7765 ( .A1(n8253), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6258) );
  NAND2_X1 U7766 ( .A1(n6280), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6257) );
  NAND2_X1 U7767 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6261) );
  MUX2_X1 U7768 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6261), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n6264) );
  INV_X1 U7769 ( .A(n6262), .ZN(n6263) );
  NAND2_X1 U7770 ( .A1(n6264), .A2(n6263), .ZN(n7014) );
  NAND2_X2 U7771 ( .A1(n6266), .A2(n6814), .ZN(n6563) );
  OR2_X1 U7772 ( .A1(n6563), .A2(n6815), .ZN(n6268) );
  OR2_X1 U7773 ( .A1(n4510), .A2(n6816), .ZN(n6267) );
  NAND2_X1 U7774 ( .A1(n6980), .A2(n6571), .ZN(n6269) );
  AND2_X1 U7775 ( .A1(n6269), .A2(n8296), .ZN(n8795) );
  NAND2_X1 U7776 ( .A1(n6280), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6272) );
  NAND2_X1 U7777 ( .A1(n6309), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U7778 ( .A1(n4515), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6270) );
  OR2_X1 U7779 ( .A1(n6563), .A2(n6818), .ZN(n6278) );
  OR2_X1 U7780 ( .A1(n6274), .A2(n6819), .ZN(n6277) );
  OR2_X1 U7781 ( .A1(n6266), .A2(n7099), .ZN(n6276) );
  NAND2_X1 U7782 ( .A1(n8795), .A2(n8262), .ZN(n8794) );
  NAND2_X1 U7783 ( .A1(n4878), .A2(n9996), .ZN(n6279) );
  NAND2_X1 U7784 ( .A1(n6280), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6283) );
  INV_X1 U7785 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7022) );
  NAND2_X1 U7786 ( .A1(n6545), .A2(n7022), .ZN(n6281) );
  AND3_X1 U7787 ( .A1(n6283), .A2(n6282), .A3(n6281), .ZN(n6285) );
  NAND2_X1 U7788 ( .A1(n6483), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6284) );
  OR2_X1 U7789 ( .A1(n6563), .A2(n6820), .ZN(n6291) );
  OR2_X1 U7790 ( .A1(n6274), .A2(n6817), .ZN(n6290) );
  NAND2_X1 U7791 ( .A1(n6275), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6286) );
  MUX2_X1 U7792 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6286), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n6288) );
  NAND2_X1 U7793 ( .A1(n6288), .A2(n6287), .ZN(n7029) );
  OR2_X1 U7794 ( .A1(n6266), .A2(n7029), .ZN(n6289) );
  NAND2_X1 U7795 ( .A1(n6293), .A2(n6292), .ZN(n8303) );
  NAND2_X1 U7796 ( .A1(n8799), .A2(n10003), .ZN(n8309) );
  NAND2_X1 U7797 ( .A1(n8303), .A2(n8309), .ZN(n7586) );
  INV_X1 U7798 ( .A(n7586), .ZN(n8264) );
  NAND2_X1 U7799 ( .A1(n8294), .A2(n8264), .ZN(n6294) );
  NAND2_X1 U7800 ( .A1(n6294), .A2(n8303), .ZN(n7594) );
  NAND2_X1 U7801 ( .A1(n8253), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U7802 ( .A1(n8254), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U7803 ( .A1(n6483), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6298) );
  NOR2_X1 U7804 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6307) );
  AND2_X1 U7805 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6296) );
  NOR2_X1 U7806 ( .A1(n6307), .A2(n6296), .ZN(n7381) );
  OR2_X1 U7807 ( .A1(n6256), .A2(n7381), .ZN(n6297) );
  NAND2_X1 U7808 ( .A1(n6287), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6302) );
  INV_X1 U7809 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6301) );
  XNOR2_X1 U7810 ( .A(n6302), .B(n6301), .ZN(n7172) );
  OR2_X1 U7811 ( .A1(n6563), .A2(n6823), .ZN(n6304) );
  OR2_X1 U7812 ( .A1(n6274), .A2(n6822), .ZN(n6303) );
  INV_X1 U7813 ( .A(n7596), .ZN(n10008) );
  NAND2_X1 U7814 ( .A1(n8480), .A2(n10008), .ZN(n8304) );
  NAND2_X1 U7815 ( .A1(n7594), .A2(n8304), .ZN(n6305) );
  NAND2_X1 U7816 ( .A1(n7605), .A2(n7596), .ZN(n8311) );
  NAND2_X1 U7817 ( .A1(n6305), .A2(n8311), .ZN(n7608) );
  NAND2_X1 U7818 ( .A1(n8253), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6313) );
  NAND2_X1 U7819 ( .A1(n8254), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U7820 ( .A1(n6307), .A2(n6306), .ZN(n6321) );
  OR2_X1 U7821 ( .A1(n6307), .A2(n6306), .ZN(n6308) );
  NAND2_X1 U7822 ( .A1(n6321), .A2(n6308), .ZN(n7609) );
  NAND2_X1 U7823 ( .A1(n6565), .A2(n7609), .ZN(n6311) );
  NAND2_X1 U7824 ( .A1(n6483), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6310) );
  NAND4_X1 U7825 ( .A1(n6313), .A2(n6312), .A3(n6311), .A4(n6310), .ZN(n8479)
         );
  OR2_X1 U7826 ( .A1(n6563), .A2(n6827), .ZN(n6320) );
  OR2_X1 U7827 ( .A1(n6274), .A2(n6828), .ZN(n6319) );
  NOR2_X1 U7828 ( .A1(n6314), .A2(n8955), .ZN(n6315) );
  MUX2_X1 U7829 ( .A(n8955), .B(n6315), .S(P2_IR_REG_5__SCAN_IN), .Z(n6317) );
  OR2_X1 U7830 ( .A1(n6317), .A2(n6316), .ZN(n7056) );
  OR2_X1 U7831 ( .A1(n6266), .A2(n7056), .ZN(n6318) );
  OR2_X1 U7832 ( .A1(n8479), .A2(n10012), .ZN(n8310) );
  NAND2_X1 U7833 ( .A1(n8479), .A2(n10012), .ZN(n8314) );
  NAND2_X1 U7834 ( .A1(n8310), .A2(n8314), .ZN(n8268) );
  INV_X1 U7835 ( .A(n8268), .ZN(n7607) );
  NAND2_X1 U7836 ( .A1(n8253), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U7837 ( .A1(n8254), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U7838 ( .A1(n6321), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6322) );
  NAND2_X1 U7839 ( .A1(n6335), .A2(n6322), .ZN(n7500) );
  NAND2_X1 U7840 ( .A1(n6565), .A2(n7500), .ZN(n6324) );
  NAND2_X1 U7841 ( .A1(n6483), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6323) );
  NAND4_X1 U7842 ( .A1(n6326), .A2(n6325), .A3(n6324), .A4(n6323), .ZN(n8478)
         );
  NOR2_X1 U7843 ( .A1(n6316), .A2(n8955), .ZN(n6327) );
  MUX2_X1 U7844 ( .A(n8955), .B(n6327), .S(P2_IR_REG_6__SCAN_IN), .Z(n6330) );
  INV_X1 U7845 ( .A(n6328), .ZN(n6329) );
  AOI22_X1 U7846 ( .A1(n8249), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6470), .B2(
        n4691), .ZN(n6333) );
  NAND2_X1 U7847 ( .A1(n6331), .A2(n8250), .ZN(n6332) );
  OR2_X1 U7848 ( .A1(n8478), .A2(n10019), .ZN(n8316) );
  AND2_X1 U7849 ( .A1(n8310), .A2(n8316), .ZN(n8307) );
  NAND2_X1 U7850 ( .A1(n7606), .A2(n8307), .ZN(n6334) );
  NAND2_X1 U7851 ( .A1(n8478), .A2(n10019), .ZN(n8318) );
  NAND2_X1 U7852 ( .A1(n6334), .A2(n8318), .ZN(n7661) );
  NAND2_X1 U7853 ( .A1(n8254), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6340) );
  NAND2_X1 U7854 ( .A1(n6483), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6339) );
  AND2_X1 U7855 ( .A1(n6335), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6336) );
  OR2_X1 U7856 ( .A1(n6336), .A2(n6348), .ZN(n7664) );
  NAND2_X1 U7857 ( .A1(n6565), .A2(n7664), .ZN(n6338) );
  NAND2_X1 U7858 ( .A1(n8253), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6337) );
  NAND4_X1 U7859 ( .A1(n6340), .A2(n6339), .A3(n6338), .A4(n6337), .ZN(n8477)
         );
  NAND2_X1 U7860 ( .A1(n6832), .A2(n8250), .ZN(n6342) );
  NAND2_X1 U7861 ( .A1(n6328), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6343) );
  XNOR2_X1 U7862 ( .A(n6343), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7065) );
  AOI22_X1 U7863 ( .A1(n8249), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6470), .B2(
        n7065), .ZN(n6341) );
  NAND2_X1 U7864 ( .A1(n6342), .A2(n6341), .ZN(n8324) );
  XNOR2_X1 U7865 ( .A(n8477), .B(n8324), .ZN(n8323) );
  INV_X1 U7866 ( .A(n8324), .ZN(n10024) );
  NAND2_X1 U7867 ( .A1(n10024), .A2(n8477), .ZN(n8332) );
  NAND2_X1 U7868 ( .A1(n6836), .A2(n8250), .ZN(n6347) );
  NAND2_X1 U7869 ( .A1(n6343), .A2(n6207), .ZN(n6344) );
  NAND2_X1 U7870 ( .A1(n6344), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6345) );
  XNOR2_X1 U7871 ( .A(n6345), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7204) );
  AOI22_X1 U7872 ( .A1(n8249), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6470), .B2(
        n7204), .ZN(n6346) );
  NAND2_X1 U7873 ( .A1(n6347), .A2(n6346), .ZN(n7770) );
  INV_X1 U7874 ( .A(n7770), .ZN(n10030) );
  NAND2_X1 U7875 ( .A1(n8254), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6353) );
  NAND2_X1 U7876 ( .A1(n8253), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6352) );
  NOR2_X1 U7877 ( .A1(n6348), .A2(n7195), .ZN(n6349) );
  OR2_X1 U7878 ( .A1(n6361), .A2(n6349), .ZN(n7765) );
  NAND2_X1 U7879 ( .A1(n6565), .A2(n7765), .ZN(n6351) );
  NAND2_X1 U7880 ( .A1(n6483), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6350) );
  INV_X1 U7881 ( .A(n7920), .ZN(n8476) );
  INV_X1 U7882 ( .A(n8335), .ZN(n6354) );
  NAND2_X1 U7883 ( .A1(n7770), .A2(n7920), .ZN(n8327) );
  NAND2_X1 U7884 ( .A1(n6849), .A2(n8250), .ZN(n6359) );
  NAND2_X1 U7885 ( .A1(n6356), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6357) );
  XNOR2_X1 U7886 ( .A(n6357), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7318) );
  AOI22_X1 U7887 ( .A1(n8249), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6470), .B2(
        n7318), .ZN(n6358) );
  NAND2_X1 U7888 ( .A1(n6359), .A2(n6358), .ZN(n10039) );
  NAND2_X1 U7889 ( .A1(n8253), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6366) );
  NAND2_X1 U7890 ( .A1(n8254), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6365) );
  OR2_X1 U7891 ( .A1(n6361), .A2(n6360), .ZN(n6362) );
  NAND2_X1 U7892 ( .A1(n6372), .A2(n6362), .ZN(n7916) );
  NAND2_X1 U7893 ( .A1(n6565), .A2(n7916), .ZN(n6364) );
  NAND2_X1 U7894 ( .A1(n6483), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6363) );
  NAND4_X1 U7895 ( .A1(n6366), .A2(n6365), .A3(n6364), .A4(n6363), .ZN(n8475)
         );
  NAND2_X1 U7896 ( .A1(n10039), .A2(n7934), .ZN(n8329) );
  NAND2_X1 U7897 ( .A1(n8336), .A2(n8329), .ZN(n8272) );
  INV_X1 U7898 ( .A(n8272), .ZN(n6367) );
  NAND2_X1 U7899 ( .A1(n6853), .A2(n8250), .ZN(n6371) );
  OR2_X1 U7900 ( .A1(n6368), .A2(n8955), .ZN(n6369) );
  XNOR2_X1 U7901 ( .A(n6369), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7338) );
  AOI22_X1 U7902 ( .A1(n8249), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6470), .B2(
        n7338), .ZN(n6370) );
  NAND2_X1 U7903 ( .A1(n6371), .A2(n6370), .ZN(n10045) );
  NAND2_X1 U7904 ( .A1(n8254), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6377) );
  NAND2_X1 U7905 ( .A1(n6483), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U7906 ( .A1(n6372), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U7907 ( .A1(n6385), .A2(n6373), .ZN(n7930) );
  NAND2_X1 U7908 ( .A1(n6565), .A2(n7930), .ZN(n6375) );
  NAND2_X1 U7909 ( .A1(n8253), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6374) );
  NAND4_X1 U7910 ( .A1(n6377), .A2(n6376), .A3(n6375), .A4(n6374), .ZN(n8474)
         );
  OR2_X1 U7911 ( .A1(n10045), .A2(n7740), .ZN(n8344) );
  NAND2_X1 U7912 ( .A1(n10045), .A2(n7740), .ZN(n8328) );
  NAND2_X1 U7913 ( .A1(n6868), .A2(n8250), .ZN(n6384) );
  OR2_X1 U7914 ( .A1(n6378), .A2(n8955), .ZN(n6381) );
  INV_X1 U7915 ( .A(n6381), .ZN(n6379) );
  NAND2_X1 U7916 ( .A1(n6379), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n6382) );
  INV_X1 U7917 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6380) );
  NAND2_X1 U7918 ( .A1(n6381), .A2(n6380), .ZN(n6392) );
  AOI22_X1 U7919 ( .A1(n8249), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6470), .B2(
        n7558), .ZN(n6383) );
  NAND2_X1 U7920 ( .A1(n6384), .A2(n6383), .ZN(n7973) );
  NAND2_X1 U7921 ( .A1(n8254), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6390) );
  NAND2_X1 U7922 ( .A1(n8253), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U7923 ( .A1(n6385), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U7924 ( .A1(n6396), .A2(n6386), .ZN(n7980) );
  NAND2_X1 U7925 ( .A1(n6565), .A2(n7980), .ZN(n6388) );
  NAND2_X1 U7926 ( .A1(n6483), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6387) );
  NAND2_X1 U7927 ( .A1(n7973), .A2(n7802), .ZN(n8346) );
  AND2_X1 U7928 ( .A1(n8346), .A2(n8328), .ZN(n8343) );
  NAND2_X1 U7929 ( .A1(n6391), .A2(n8345), .ZN(n7897) );
  NAND2_X1 U7930 ( .A1(n6938), .A2(n8250), .ZN(n6395) );
  NAND2_X1 U7931 ( .A1(n6392), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6393) );
  AOI22_X1 U7932 ( .A1(n8249), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8490), .B2(
        n6470), .ZN(n6394) );
  NAND2_X1 U7933 ( .A1(n8253), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6401) );
  NAND2_X1 U7934 ( .A1(n8254), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6400) );
  AND2_X1 U7935 ( .A1(n6396), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6397) );
  OR2_X1 U7936 ( .A1(n6397), .A2(n6407), .ZN(n8019) );
  NAND2_X1 U7937 ( .A1(n6565), .A2(n8019), .ZN(n6399) );
  NAND2_X1 U7938 ( .A1(n6483), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6398) );
  NAND4_X1 U7939 ( .A1(n6401), .A2(n6400), .A3(n6399), .A4(n6398), .ZN(n8472)
         );
  INV_X1 U7940 ( .A(n8472), .ZN(n8197) );
  NAND2_X1 U7941 ( .A1(n8012), .A2(n8197), .ZN(n8355) );
  NAND2_X1 U7942 ( .A1(n6941), .A2(n8250), .ZN(n6405) );
  OR2_X1 U7943 ( .A1(n6402), .A2(n8955), .ZN(n6403) );
  XNOR2_X1 U7944 ( .A(n6403), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9938) );
  AOI22_X1 U7945 ( .A1(n8249), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6470), .B2(
        n9938), .ZN(n6404) );
  NAND2_X1 U7946 ( .A1(n8253), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6412) );
  NAND2_X1 U7947 ( .A1(n8254), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6411) );
  NAND2_X1 U7948 ( .A1(n6407), .A2(n6406), .ZN(n6418) );
  OR2_X1 U7949 ( .A1(n6407), .A2(n6406), .ZN(n6408) );
  NAND2_X1 U7950 ( .A1(n6418), .A2(n6408), .ZN(n8194) );
  NAND2_X1 U7951 ( .A1(n6565), .A2(n8194), .ZN(n6410) );
  NAND2_X1 U7952 ( .A1(n6309), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6409) );
  NAND4_X1 U7953 ( .A1(n6412), .A2(n6411), .A3(n6410), .A4(n6409), .ZN(n8471)
         );
  NAND2_X1 U7954 ( .A1(n8358), .A2(n8116), .ZN(n6413) );
  NAND2_X1 U7955 ( .A1(n6414), .A2(n6413), .ZN(n7988) );
  NAND2_X1 U7956 ( .A1(n6976), .A2(n8250), .ZN(n6417) );
  NAND2_X1 U7957 ( .A1(n6415), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6438) );
  XNOR2_X1 U7958 ( .A(n6438), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8502) );
  AOI22_X1 U7959 ( .A1(n8249), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8502), .B2(
        n6470), .ZN(n6416) );
  NAND2_X1 U7960 ( .A1(n4515), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6423) );
  NAND2_X1 U7961 ( .A1(n8254), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6422) );
  NAND2_X1 U7962 ( .A1(n6418), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6419) );
  NAND2_X1 U7963 ( .A1(n6429), .A2(n6419), .ZN(n8113) );
  NAND2_X1 U7964 ( .A1(n6565), .A2(n8113), .ZN(n6421) );
  NAND2_X1 U7965 ( .A1(n6309), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6420) );
  NAND4_X1 U7966 ( .A1(n6423), .A2(n6422), .A3(n6421), .A4(n6420), .ZN(n8470)
         );
  INV_X1 U7967 ( .A(n8470), .ZN(n8005) );
  AND2_X1 U7968 ( .A1(n8118), .A2(n8005), .ZN(n7984) );
  OR2_X1 U7969 ( .A1(n8118), .A2(n8005), .ZN(n8368) );
  NAND2_X1 U7970 ( .A1(n6985), .A2(n8250), .ZN(n6428) );
  NAND2_X1 U7971 ( .A1(n6438), .A2(n6424), .ZN(n6425) );
  NAND2_X1 U7972 ( .A1(n6425), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6426) );
  XNOR2_X1 U7973 ( .A(n6426), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8522) );
  AOI22_X1 U7974 ( .A1(n8522), .A2(n6470), .B1(n8249), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6427) );
  NAND2_X1 U7975 ( .A1(n8253), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6435) );
  NAND2_X1 U7976 ( .A1(n8254), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6434) );
  INV_X1 U7977 ( .A(n6444), .ZN(n6431) );
  NAND2_X1 U7978 ( .A1(n6429), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6430) );
  NAND2_X1 U7979 ( .A1(n6431), .A2(n6430), .ZN(n8242) );
  NAND2_X1 U7980 ( .A1(n6565), .A2(n8242), .ZN(n6433) );
  NAND2_X1 U7981 ( .A1(n6309), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6432) );
  OR2_X1 U7982 ( .A1(n8007), .A2(n8778), .ZN(n8372) );
  NAND2_X1 U7983 ( .A1(n8007), .A2(n8778), .ZN(n8387) );
  NAND2_X1 U7984 ( .A1(n8372), .A2(n8387), .ZN(n8279) );
  NAND2_X1 U7985 ( .A1(n7148), .A2(n8250), .ZN(n6442) );
  NAND2_X1 U7986 ( .A1(n6436), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6437) );
  NAND2_X1 U7987 ( .A1(n6438), .A2(n6437), .ZN(n6439) );
  NAND2_X1 U7988 ( .A1(n6439), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n6440) );
  AOI22_X1 U7989 ( .A1(n8537), .A2(n6470), .B1(n8249), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n6441) );
  NAND2_X1 U7990 ( .A1(n8254), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6449) );
  NAND2_X1 U7991 ( .A1(n6483), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6448) );
  INV_X1 U7992 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6443) );
  NOR2_X1 U7993 ( .A1(n6444), .A2(n6443), .ZN(n6445) );
  OR2_X1 U7994 ( .A1(n6464), .A2(n6445), .ZN(n8789) );
  NAND2_X1 U7995 ( .A1(n6565), .A2(n8789), .ZN(n6447) );
  NAND2_X1 U7996 ( .A1(n4515), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6446) );
  NAND2_X1 U7997 ( .A1(n8944), .A2(n8239), .ZN(n8373) );
  NAND2_X1 U7998 ( .A1(n7375), .A2(n8250), .ZN(n6454) );
  NAND2_X1 U7999 ( .A1(n6450), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6451) );
  XNOR2_X1 U8000 ( .A(n6451), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8566) );
  NOR2_X1 U8001 ( .A1(n6274), .A2(n10284), .ZN(n6452) );
  AOI21_X1 U8002 ( .B1(n8566), .B2(n6470), .A(n6452), .ZN(n6453) );
  NAND2_X1 U8003 ( .A1(n8254), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U8004 ( .A1(n4515), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6457) );
  NAND2_X1 U8005 ( .A1(n6309), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6456) );
  XNOR2_X1 U8006 ( .A(n6464), .B(P2_REG3_REG_17__SCAN_IN), .ZN(n8773) );
  OR2_X1 U8007 ( .A1(n6256), .A2(n8773), .ZN(n6455) );
  OR2_X1 U8008 ( .A1(n8937), .A2(n8749), .ZN(n8389) );
  NAND2_X1 U8009 ( .A1(n8937), .A2(n8749), .ZN(n8376) );
  NAND2_X1 U8010 ( .A1(n8389), .A2(n8376), .ZN(n8761) );
  OR2_X2 U8011 ( .A1(n8762), .A2(n8761), .ZN(n8759) );
  NAND2_X1 U8012 ( .A1(n7388), .A2(n8250), .ZN(n6461) );
  NAND2_X1 U8013 ( .A1(n4612), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6459) );
  XNOR2_X1 U8014 ( .A(n6459), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8557) );
  AOI22_X1 U8015 ( .A1(n8557), .A2(n6470), .B1(n8249), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n6460) );
  NAND2_X1 U8016 ( .A1(n8253), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6469) );
  NAND2_X1 U8017 ( .A1(n8254), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6468) );
  INV_X1 U8018 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10348) );
  NAND2_X1 U8019 ( .A1(n6464), .A2(n10348), .ZN(n6462) );
  NAND2_X1 U8020 ( .A1(n6462), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6465) );
  NOR2_X1 U8021 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_17__SCAN_IN), 
        .ZN(n6463) );
  NAND2_X1 U8022 ( .A1(n6465), .A2(n6473), .ZN(n8754) );
  NAND2_X1 U8023 ( .A1(n6565), .A2(n8754), .ZN(n6467) );
  NAND2_X1 U8024 ( .A1(n6483), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U8025 ( .A1(n8854), .A2(n8164), .ZN(n8392) );
  NAND2_X1 U8026 ( .A1(n7616), .A2(n8250), .ZN(n6472) );
  AOI22_X1 U8027 ( .A1(n8459), .A2(n6470), .B1(n8249), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U8028 ( .A1(n6473), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6474) );
  NAND2_X1 U8029 ( .A1(n6481), .A2(n6474), .ZN(n8738) );
  NAND2_X1 U8030 ( .A1(n8738), .A2(n6565), .ZN(n6478) );
  NAND2_X1 U8031 ( .A1(n8253), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U8032 ( .A1(n8254), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6476) );
  NAND2_X1 U8033 ( .A1(n6309), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6475) );
  OR2_X1 U8034 ( .A1(n8850), .A2(n8747), .ZN(n8395) );
  AND2_X1 U8035 ( .A1(n8395), .A2(n8735), .ZN(n8379) );
  NAND2_X1 U8036 ( .A1(n8850), .A2(n8747), .ZN(n8393) );
  NAND2_X1 U8037 ( .A1(n7658), .A2(n8250), .ZN(n6480) );
  INV_X1 U8038 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7659) );
  OR2_X1 U8039 ( .A1(n6274), .A2(n7659), .ZN(n6479) );
  AND2_X1 U8040 ( .A1(n6481), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6482) );
  OR2_X1 U8041 ( .A1(n6482), .A2(n6489), .ZN(n8723) );
  NAND2_X1 U8042 ( .A1(n8723), .A2(n6565), .ZN(n6486) );
  AOI22_X1 U8043 ( .A1(n8253), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n8254), .B2(
        P2_REG1_REG_20__SCAN_IN), .ZN(n6485) );
  NAND2_X1 U8044 ( .A1(n6483), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6484) );
  NAND2_X1 U8045 ( .A1(n8722), .A2(n8705), .ZN(n8397) );
  NAND2_X1 U8046 ( .A1(n7773), .A2(n8250), .ZN(n6488) );
  OR2_X1 U8047 ( .A1(n6274), .A2(n7774), .ZN(n6487) );
  INV_X1 U8048 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8135) );
  OR2_X1 U8049 ( .A1(n6489), .A2(n8135), .ZN(n6490) );
  NAND2_X1 U8050 ( .A1(n6497), .A2(n6490), .ZN(n8709) );
  NAND2_X1 U8051 ( .A1(n8709), .A2(n6565), .ZN(n6493) );
  AOI22_X1 U8052 ( .A1(n4515), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n8254), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n6492) );
  NAND2_X1 U8053 ( .A1(n6309), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6491) );
  NAND2_X1 U8054 ( .A1(n8708), .A2(n6740), .ZN(n8398) );
  NAND2_X1 U8055 ( .A1(n8707), .A2(n8398), .ZN(n6494) );
  NAND2_X1 U8056 ( .A1(n6494), .A2(n8399), .ZN(n8693) );
  NAND2_X1 U8057 ( .A1(n7864), .A2(n8250), .ZN(n6496) );
  OR2_X1 U8058 ( .A1(n6274), .A2(n7868), .ZN(n6495) );
  NAND2_X1 U8059 ( .A1(n6497), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6498) );
  NAND2_X1 U8060 ( .A1(n6505), .A2(n6498), .ZN(n8699) );
  INV_X1 U8061 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8698) );
  INV_X1 U8062 ( .A(n6309), .ZN(n6621) );
  NAND2_X1 U8063 ( .A1(n8253), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6500) );
  NAND2_X1 U8064 ( .A1(n8254), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6499) );
  OAI211_X1 U8065 ( .C1(n8698), .C2(n6621), .A(n6500), .B(n6499), .ZN(n6501)
         );
  AOI21_X1 U8066 ( .B1(n8699), .B2(n6565), .A(n6501), .ZN(n8704) );
  OR2_X1 U8067 ( .A1(n8914), .A2(n8704), .ZN(n8405) );
  INV_X1 U8068 ( .A(n8405), .ZN(n6502) );
  NAND2_X1 U8069 ( .A1(n8914), .A2(n8704), .ZN(n8406) );
  NAND2_X1 U8070 ( .A1(n7914), .A2(n8250), .ZN(n6504) );
  OR2_X1 U8071 ( .A1(n6274), .A2(n10214), .ZN(n6503) );
  NAND2_X1 U8072 ( .A1(n6505), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U8073 ( .A1(n6514), .A2(n6506), .ZN(n8689) );
  NAND2_X1 U8074 ( .A1(n8689), .A2(n6565), .ZN(n6511) );
  INV_X1 U8075 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8688) );
  NAND2_X1 U8076 ( .A1(n8254), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6508) );
  NAND2_X1 U8077 ( .A1(n4515), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6507) );
  OAI211_X1 U8078 ( .C1(n6621), .C2(n8688), .A(n6508), .B(n6507), .ZN(n6509)
         );
  INV_X1 U8079 ( .A(n6509), .ZN(n6510) );
  NAND2_X1 U8080 ( .A1(n8682), .A2(n8411), .ZN(n8667) );
  NAND2_X1 U8081 ( .A1(n7938), .A2(n8250), .ZN(n6513) );
  OR2_X1 U8082 ( .A1(n6274), .A2(n7939), .ZN(n6512) );
  AND2_X1 U8083 ( .A1(n6514), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6515) );
  OR2_X1 U8084 ( .A1(n6515), .A2(n6524), .ZN(n8673) );
  NAND2_X1 U8085 ( .A1(n8673), .A2(n6565), .ZN(n6520) );
  INV_X1 U8086 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8901) );
  NAND2_X1 U8087 ( .A1(n8254), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U8088 ( .A1(n6483), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6516) );
  OAI211_X1 U8089 ( .C1(n8901), .C2(n6295), .A(n6517), .B(n6516), .ZN(n6518)
         );
  INV_X1 U8090 ( .A(n6518), .ZN(n6519) );
  NAND2_X1 U8091 ( .A1(n8902), .A2(n8174), .ZN(n8416) );
  NAND2_X1 U8092 ( .A1(n8908), .A2(n8205), .ZN(n8666) );
  AND2_X1 U8093 ( .A1(n8416), .A2(n8666), .ZN(n8412) );
  NAND2_X1 U8094 ( .A1(n8667), .A2(n8412), .ZN(n6521) );
  NAND2_X1 U8095 ( .A1(n6521), .A2(n8415), .ZN(n8654) );
  NAND2_X1 U8096 ( .A1(n7991), .A2(n8250), .ZN(n6523) );
  OR2_X1 U8097 ( .A1(n4510), .A2(n7992), .ZN(n6522) );
  INV_X1 U8098 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8143) );
  NOR2_X1 U8099 ( .A1(n6524), .A2(n8143), .ZN(n6525) );
  OR2_X1 U8100 ( .A1(n6532), .A2(n6525), .ZN(n8659) );
  INV_X1 U8101 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n10293) );
  NAND2_X1 U8102 ( .A1(n8253), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6527) );
  NAND2_X1 U8103 ( .A1(n6309), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6526) );
  OAI211_X1 U8104 ( .C1(n6528), .C2(n10293), .A(n6527), .B(n6526), .ZN(n6529)
         );
  NAND2_X1 U8105 ( .A1(n8896), .A2(n8224), .ZN(n8421) );
  NAND2_X1 U8106 ( .A1(n8022), .A2(n8250), .ZN(n6531) );
  OR2_X1 U8107 ( .A1(n6274), .A2(n8023), .ZN(n6530) );
  INV_X1 U8108 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8222) );
  NOR2_X1 U8109 ( .A1(n6532), .A2(n8222), .ZN(n6533) );
  NAND2_X1 U8110 ( .A1(n8650), .A2(n6565), .ZN(n6538) );
  INV_X1 U8111 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8649) );
  NAND2_X1 U8112 ( .A1(n8253), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6535) );
  NAND2_X1 U8113 ( .A1(n8254), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6534) );
  OAI211_X1 U8114 ( .C1(n8649), .C2(n6621), .A(n6535), .B(n6534), .ZN(n6536)
         );
  INV_X1 U8115 ( .A(n6536), .ZN(n6537) );
  NAND2_X1 U8116 ( .A1(n6538), .A2(n6537), .ZN(n8657) );
  NOR2_X1 U8117 ( .A1(n8890), .A2(n8635), .ZN(n8288) );
  NAND2_X1 U8118 ( .A1(n8890), .A2(n8635), .ZN(n8261) );
  NAND2_X1 U8119 ( .A1(n6539), .A2(n8261), .ZN(n8632) );
  NAND2_X1 U8120 ( .A1(n8096), .A2(n8250), .ZN(n6542) );
  OR2_X1 U8121 ( .A1(n4510), .A2(n6540), .ZN(n6541) );
  INV_X1 U8122 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8105) );
  NAND2_X1 U8123 ( .A1(n6543), .A2(n8105), .ZN(n6554) );
  OR2_X1 U8124 ( .A1(n6543), .A2(n8105), .ZN(n6544) );
  NAND2_X1 U8125 ( .A1(n6554), .A2(n6544), .ZN(n8640) );
  NAND2_X1 U8126 ( .A1(n8640), .A2(n6545), .ZN(n6550) );
  INV_X1 U8127 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n10311) );
  NAND2_X1 U8128 ( .A1(n6309), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6547) );
  NAND2_X1 U8129 ( .A1(n8254), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6546) );
  OAI211_X1 U8130 ( .C1(n6295), .C2(n10311), .A(n6547), .B(n6546), .ZN(n6548)
         );
  INV_X1 U8131 ( .A(n6548), .ZN(n6549) );
  OR2_X1 U8132 ( .A1(n8884), .A2(n8624), .ZN(n8426) );
  NAND2_X1 U8133 ( .A1(n8094), .A2(n8250), .ZN(n6553) );
  OR2_X1 U8134 ( .A1(n6274), .A2(n6551), .ZN(n6552) );
  NAND2_X1 U8135 ( .A1(n6554), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6555) );
  NAND2_X1 U8136 ( .A1(n8614), .A2(n6555), .ZN(n8629) );
  NAND2_X1 U8137 ( .A1(n8629), .A2(n6565), .ZN(n6560) );
  INV_X1 U8138 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U8139 ( .A1(n8253), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6557) );
  NAND2_X1 U8140 ( .A1(n8254), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6556) );
  OAI211_X1 U8141 ( .C1(n8628), .C2(n6621), .A(n6557), .B(n6556), .ZN(n6558)
         );
  INV_X1 U8142 ( .A(n6558), .ZN(n6559) );
  NAND2_X1 U8143 ( .A1(n8621), .A2(n8622), .ZN(n6562) );
  OR2_X1 U8144 ( .A1(n8879), .A2(n8636), .ZN(n6561) );
  INV_X1 U8145 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n10238) );
  OR2_X1 U8146 ( .A1(n6274), .A2(n10238), .ZN(n6564) );
  INV_X1 U8147 ( .A(n8614), .ZN(n6566) );
  NAND2_X1 U8148 ( .A1(n6566), .A2(n6565), .ZN(n8259) );
  INV_X1 U8149 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n10271) );
  NAND2_X1 U8150 ( .A1(n8254), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6568) );
  NAND2_X1 U8151 ( .A1(n6309), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6567) );
  OAI211_X1 U8152 ( .C1(n10271), .C2(n6295), .A(n6568), .B(n6567), .ZN(n6569)
         );
  INV_X1 U8153 ( .A(n6569), .ZN(n6570) );
  NAND2_X1 U8154 ( .A1(n8616), .A2(n8625), .ZN(n8252) );
  XNOR2_X1 U8155 ( .A(n8251), .B(n8429), .ZN(n8611) );
  NAND2_X1 U8156 ( .A1(n8482), .A2(n7369), .ZN(n7175) );
  NAND2_X1 U8157 ( .A1(n7173), .A2(n7175), .ZN(n6576) );
  NAND2_X1 U8158 ( .A1(n6574), .A2(n7265), .ZN(n6575) );
  NAND2_X1 U8159 ( .A1(n6576), .A2(n6575), .ZN(n8797) );
  NAND2_X1 U8160 ( .A1(n8797), .A2(n8798), .ZN(n6578) );
  OR2_X1 U8161 ( .A1(n8481), .A2(n9996), .ZN(n6577) );
  NAND2_X1 U8162 ( .A1(n6578), .A2(n6577), .ZN(n7585) );
  NAND2_X1 U8163 ( .A1(n7585), .A2(n7586), .ZN(n6580) );
  OR2_X1 U8164 ( .A1(n8799), .A2(n6292), .ZN(n6579) );
  INV_X1 U8165 ( .A(n10012), .ZN(n7610) );
  OR2_X1 U8166 ( .A1(n8479), .A2(n7610), .ZN(n7492) );
  NAND2_X1 U8167 ( .A1(n7491), .A2(n7492), .ZN(n6581) );
  NAND2_X1 U8168 ( .A1(n8316), .A2(n8318), .ZN(n8266) );
  NAND2_X1 U8169 ( .A1(n6581), .A2(n8266), .ZN(n7495) );
  INV_X1 U8170 ( .A(n10019), .ZN(n7497) );
  OR2_X1 U8171 ( .A1(n8478), .A2(n7497), .ZN(n6582) );
  NAND2_X1 U8172 ( .A1(n7495), .A2(n6582), .ZN(n7665) );
  NAND2_X1 U8173 ( .A1(n8477), .A2(n8324), .ZN(n6583) );
  NAND2_X1 U8174 ( .A1(n7665), .A2(n6583), .ZN(n6585) );
  OR2_X1 U8175 ( .A1(n8477), .A2(n8324), .ZN(n6584) );
  OR2_X1 U8176 ( .A1(n10039), .A2(n8475), .ZN(n6586) );
  NAND2_X1 U8177 ( .A1(n7739), .A2(n6586), .ZN(n6588) );
  NAND2_X1 U8178 ( .A1(n10039), .A2(n8475), .ZN(n6587) );
  NAND2_X1 U8179 ( .A1(n6588), .A2(n6587), .ZN(n7800) );
  OR2_X1 U8180 ( .A1(n10045), .A2(n8474), .ZN(n6589) );
  NAND2_X1 U8181 ( .A1(n7800), .A2(n6589), .ZN(n6591) );
  NAND2_X1 U8182 ( .A1(n10045), .A2(n8474), .ZN(n6590) );
  NAND2_X1 U8183 ( .A1(n6591), .A2(n6590), .ZN(n7884) );
  NAND2_X1 U8184 ( .A1(n8345), .A2(n8346), .ZN(n8275) );
  NAND2_X1 U8185 ( .A1(n7884), .A2(n8275), .ZN(n6593) );
  NAND2_X1 U8186 ( .A1(n7973), .A2(n8473), .ZN(n6592) );
  AND2_X1 U8187 ( .A1(n8012), .A2(n8472), .ZN(n6594) );
  NOR2_X1 U8188 ( .A1(n8358), .A2(n8471), .ZN(n8362) );
  OR2_X1 U8189 ( .A1(n8118), .A2(n8470), .ZN(n6595) );
  NAND2_X1 U8190 ( .A1(n8003), .A2(n8279), .ZN(n6597) );
  OR2_X1 U8191 ( .A1(n8007), .A2(n8469), .ZN(n6596) );
  INV_X1 U8192 ( .A(n8239), .ZN(n8768) );
  NAND2_X1 U8193 ( .A1(n8944), .A2(n8768), .ZN(n8763) );
  NAND2_X1 U8194 ( .A1(n6599), .A2(n8761), .ZN(n8766) );
  NAND2_X1 U8195 ( .A1(n8937), .A2(n8787), .ZN(n6600) );
  NAND2_X1 U8196 ( .A1(n8766), .A2(n6600), .ZN(n8744) );
  INV_X1 U8197 ( .A(n8744), .ZN(n6601) );
  OR2_X1 U8198 ( .A1(n8854), .A2(n8767), .ZN(n6602) );
  NAND2_X1 U8199 ( .A1(n8850), .A2(n8718), .ZN(n6603) );
  NAND2_X1 U8200 ( .A1(n8382), .A2(n8397), .ZN(n8715) );
  OR2_X1 U8201 ( .A1(n8722), .A2(n8732), .ZN(n6604) );
  NAND2_X1 U8202 ( .A1(n8399), .A2(n8398), .ZN(n8706) );
  NAND2_X1 U8203 ( .A1(n8694), .A2(n8695), .ZN(n6606) );
  INV_X1 U8204 ( .A(n8704), .ZN(n8686) );
  OR2_X1 U8205 ( .A1(n8686), .A2(n8914), .ZN(n6605) );
  NOR2_X1 U8206 ( .A1(n8908), .A2(n8696), .ZN(n6608) );
  NAND2_X1 U8207 ( .A1(n8908), .A2(n8696), .ZN(n6607) );
  AND2_X1 U8208 ( .A1(n8685), .A2(n8902), .ZN(n6609) );
  NAND2_X1 U8209 ( .A1(n8420), .A2(n8421), .ZN(n8655) );
  OR2_X1 U8210 ( .A1(n8896), .A2(n8671), .ZN(n6610) );
  NAND2_X1 U8211 ( .A1(n6611), .A2(n6610), .ZN(n8645) );
  INV_X1 U8212 ( .A(n8645), .ZN(n6612) );
  NAND2_X1 U8213 ( .A1(n6788), .A2(n8636), .ZN(n8430) );
  XNOR2_X1 U8214 ( .A(n6613), .B(n4722), .ZN(n6616) );
  NAND2_X1 U8215 ( .A1(n6679), .A2(n8432), .ZN(n8447) );
  NAND2_X1 U8216 ( .A1(n8459), .A2(n8463), .ZN(n6632) );
  NAND2_X1 U8217 ( .A1(n6616), .A2(n8805), .ZN(n6631) );
  INV_X1 U8218 ( .A(n8463), .ZN(n7866) );
  AOI21_X1 U8219 ( .B1(n8432), .B2(n7866), .A(n8459), .ZN(n6617) );
  AND2_X1 U8220 ( .A1(n10029), .A2(n6617), .ZN(n6618) );
  INV_X1 U8221 ( .A(n6768), .ZN(n6680) );
  INV_X1 U8222 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6622) );
  NAND2_X1 U8223 ( .A1(n8253), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6620) );
  NAND2_X1 U8224 ( .A1(n8254), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6619) );
  OAI211_X1 U8225 ( .C1(n6622), .C2(n6621), .A(n6620), .B(n6619), .ZN(n6623)
         );
  INV_X1 U8226 ( .A(n6623), .ZN(n6624) );
  INV_X1 U8227 ( .A(n6625), .ZN(n8460) );
  NAND2_X1 U8228 ( .A1(n8460), .A2(n8591), .ZN(n6627) );
  NAND2_X1 U8229 ( .A1(n6266), .A2(n6627), .ZN(n6782) );
  NAND2_X1 U8230 ( .A1(n6266), .A2(P2_B_REG_SCAN_IN), .ZN(n6628) );
  NAND2_X1 U8231 ( .A1(n8800), .A2(n6628), .ZN(n8605) );
  OAI22_X1 U8232 ( .A1(n8436), .A2(n8605), .B1(n8636), .B2(n8779), .ZN(n6629)
         );
  AOI21_X1 U8233 ( .B1(n8611), .B2(n7804), .A(n6629), .ZN(n6630) );
  OR2_X1 U8234 ( .A1(n6679), .A2(n8437), .ZN(n6682) );
  INV_X1 U8235 ( .A(n6682), .ZN(n8446) );
  INV_X1 U8236 ( .A(n6632), .ZN(n6633) );
  AND2_X1 U8237 ( .A1(n8435), .A2(n10029), .ZN(n6634) );
  NAND2_X1 U8238 ( .A1(n6769), .A2(n6634), .ZN(n6756) );
  INV_X1 U8239 ( .A(n6635), .ZN(n7455) );
  NAND2_X1 U8240 ( .A1(n6756), .A2(n8676), .ZN(n6767) );
  OAI21_X2 U8241 ( .B1(n6669), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6642) );
  NAND2_X1 U8242 ( .A1(n6642), .A2(n6641), .ZN(n6643) );
  XNOR2_X2 U8243 ( .A(n6640), .B(n6639), .ZN(n7993) );
  OR2_X1 U8244 ( .A1(n6642), .A2(n6641), .ZN(n6644) );
  NAND2_X2 U8245 ( .A1(n6644), .A2(n6643), .ZN(n7940) );
  XNOR2_X1 U8246 ( .A(n7940), .B(P2_B_REG_SCAN_IN), .ZN(n6645) );
  NAND2_X1 U8247 ( .A1(n7993), .A2(n6645), .ZN(n6651) );
  NAND2_X1 U8248 ( .A1(n6646), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6647) );
  MUX2_X1 U8249 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6647), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6649) );
  NAND2_X1 U8250 ( .A1(n6649), .A2(n6648), .ZN(n8024) );
  INV_X1 U8251 ( .A(n8024), .ZN(n6650) );
  NAND2_X1 U8252 ( .A1(n7940), .A2(n8024), .ZN(n6861) );
  NAND2_X2 U8253 ( .A1(n6652), .A2(n6861), .ZN(n7362) );
  NOR2_X1 U8254 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .ZN(
        n6657) );
  NOR4_X1 U8255 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6656) );
  NOR4_X1 U8256 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6655) );
  NOR4_X1 U8257 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6654) );
  NAND4_X1 U8258 ( .A1(n6657), .A2(n6656), .A3(n6655), .A4(n6654), .ZN(n6663)
         );
  NOR4_X1 U8259 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6661) );
  NOR4_X1 U8260 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6660) );
  NOR4_X1 U8261 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n6659) );
  NOR4_X1 U8262 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6658) );
  NAND4_X1 U8263 ( .A1(n6661), .A2(n6660), .A3(n6659), .A4(n6658), .ZN(n6662)
         );
  NOR2_X1 U8264 ( .A1(n6663), .A2(n6662), .ZN(n6664) );
  NAND2_X1 U8265 ( .A1(n7362), .A2(n6796), .ZN(n6666) );
  NAND2_X1 U8266 ( .A1(n7993), .A2(n8024), .ZN(n6858) );
  INV_X1 U8267 ( .A(n7993), .ZN(n6668) );
  NOR2_X1 U8268 ( .A1(n7940), .A2(n8024), .ZN(n6667) );
  NAND2_X1 U8269 ( .A1(n6669), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6671) );
  NAND2_X1 U8270 ( .A1(n6767), .A2(n6781), .ZN(n6676) );
  INV_X1 U8271 ( .A(n7362), .ZN(n6672) );
  NAND2_X1 U8272 ( .A1(n7361), .A2(n6672), .ZN(n6799) );
  INV_X1 U8273 ( .A(n6796), .ZN(n6673) );
  NOR2_X1 U8274 ( .A1(n6799), .A2(n6673), .ZN(n6765) );
  NAND2_X1 U8275 ( .A1(n6769), .A2(n6780), .ZN(n6674) );
  NAND2_X1 U8276 ( .A1(n6762), .A2(n6674), .ZN(n6675) );
  INV_X1 U8277 ( .A(n8616), .ZN(n6804) );
  NOR2_X1 U8278 ( .A1(n10047), .A2(n10271), .ZN(n6677) );
  INV_X2 U8279 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NAND2_X1 U8280 ( .A1(n6679), .A2(n8437), .ZN(n8449) );
  XNOR2_X1 U8281 ( .A(n6685), .B(n6572), .ZN(n6989) );
  OR2_X1 U8282 ( .A1(n6683), .A2(n7369), .ZN(n6684) );
  NAND2_X1 U8283 ( .A1(n6684), .A2(n6980), .ZN(n6988) );
  NAND2_X1 U8284 ( .A1(n6989), .A2(n6988), .ZN(n6687) );
  NAND2_X1 U8285 ( .A1(n6685), .A2(n6574), .ZN(n6686) );
  NAND2_X1 U8286 ( .A1(n6687), .A2(n6686), .ZN(n7240) );
  XNOR2_X1 U8287 ( .A(n6688), .B(n4878), .ZN(n7239) );
  NAND2_X1 U8288 ( .A1(n7240), .A2(n7239), .ZN(n6691) );
  INV_X1 U8289 ( .A(n6688), .ZN(n6689) );
  NAND2_X1 U8290 ( .A1(n6689), .A2(n4878), .ZN(n6690) );
  XNOR2_X1 U8291 ( .A(n6683), .B(n10003), .ZN(n6693) );
  XNOR2_X1 U8292 ( .A(n6693), .B(n8799), .ZN(n7247) );
  NAND2_X1 U8293 ( .A1(n6693), .A2(n8799), .ZN(n6694) );
  INV_X1 U8294 ( .A(n7379), .ZN(n6696) );
  XNOR2_X1 U8295 ( .A(n4513), .B(n10008), .ZN(n6697) );
  XNOR2_X1 U8296 ( .A(n6697), .B(n8480), .ZN(n7380) );
  INV_X1 U8297 ( .A(n7380), .ZN(n6695) );
  INV_X1 U8298 ( .A(n6697), .ZN(n6698) );
  NAND2_X1 U8299 ( .A1(n6698), .A2(n7605), .ZN(n6699) );
  XNOR2_X1 U8300 ( .A(n4513), .B(n7610), .ZN(n6700) );
  XNOR2_X1 U8301 ( .A(n6700), .B(n8479), .ZN(n7410) );
  INV_X1 U8302 ( .A(n8479), .ZN(n7505) );
  INV_X1 U8303 ( .A(n7501), .ZN(n6703) );
  XNOR2_X1 U8304 ( .A(n6753), .B(n10019), .ZN(n6704) );
  XNOR2_X1 U8305 ( .A(n6704), .B(n8478), .ZN(n7502) );
  NAND2_X1 U8306 ( .A1(n6704), .A2(n8478), .ZN(n6705) );
  XNOR2_X1 U8307 ( .A(n6753), .B(n8324), .ZN(n6706) );
  XNOR2_X1 U8308 ( .A(n6706), .B(n8477), .ZN(n7697) );
  INV_X1 U8309 ( .A(n8477), .ZN(n8325) );
  XNOR2_X1 U8310 ( .A(n6753), .B(n10030), .ZN(n6707) );
  XNOR2_X1 U8311 ( .A(n6707), .B(n7920), .ZN(n7763) );
  NAND2_X1 U8312 ( .A1(n7764), .A2(n7763), .ZN(n6710) );
  INV_X1 U8313 ( .A(n6707), .ZN(n6708) );
  NAND2_X1 U8314 ( .A1(n6708), .A2(n7920), .ZN(n6709) );
  NAND2_X1 U8315 ( .A1(n6710), .A2(n6709), .ZN(n7923) );
  XNOR2_X1 U8316 ( .A(n6753), .B(n10039), .ZN(n6711) );
  XNOR2_X1 U8317 ( .A(n6711), .B(n7934), .ZN(n7924) );
  OR2_X1 U8318 ( .A1(n6711), .A2(n7934), .ZN(n6712) );
  XNOR2_X1 U8319 ( .A(n10045), .B(n6753), .ZN(n7929) );
  INV_X1 U8320 ( .A(n6713), .ZN(n6714) );
  AOI21_X2 U8321 ( .B1(n7928), .B2(n7929), .A(n5116), .ZN(n7976) );
  XNOR2_X1 U8322 ( .A(n8275), .B(n6753), .ZN(n7974) );
  NAND2_X1 U8323 ( .A1(n7976), .A2(n6715), .ZN(n7975) );
  NAND2_X1 U8324 ( .A1(n7974), .A2(n8473), .ZN(n6716) );
  NAND2_X1 U8325 ( .A1(n7975), .A2(n6716), .ZN(n8015) );
  XNOR2_X1 U8326 ( .A(n8012), .B(n6753), .ZN(n6717) );
  XNOR2_X1 U8327 ( .A(n6717), .B(n8472), .ZN(n8014) );
  INV_X1 U8328 ( .A(n6717), .ZN(n6718) );
  NAND2_X1 U8329 ( .A1(n6718), .A2(n8472), .ZN(n6719) );
  XNOR2_X1 U8330 ( .A(n8358), .B(n6753), .ZN(n6721) );
  XNOR2_X1 U8331 ( .A(n6721), .B(n8116), .ZN(n8193) );
  NAND2_X1 U8332 ( .A1(n6721), .A2(n8116), .ZN(n6722) );
  NAND2_X1 U8333 ( .A1(n8190), .A2(n6722), .ZN(n8112) );
  XNOR2_X1 U8334 ( .A(n8118), .B(n6753), .ZN(n6723) );
  XNOR2_X1 U8335 ( .A(n6723), .B(n8470), .ZN(n8111) );
  AND2_X1 U8336 ( .A1(n6723), .A2(n8005), .ZN(n6724) );
  AOI21_X2 U8337 ( .B1(n8112), .B2(n8111), .A(n6724), .ZN(n8235) );
  XNOR2_X1 U8338 ( .A(n8007), .B(n6753), .ZN(n6725) );
  XNOR2_X1 U8339 ( .A(n6725), .B(n8469), .ZN(n8234) );
  INV_X1 U8340 ( .A(n6725), .ZN(n6726) );
  NAND2_X1 U8341 ( .A1(n6726), .A2(n8469), .ZN(n6727) );
  XNOR2_X1 U8342 ( .A(n8944), .B(n6753), .ZN(n6729) );
  XNOR2_X1 U8343 ( .A(n6729), .B(n8239), .ZN(n8151) );
  NAND2_X1 U8344 ( .A1(n6729), .A2(n8239), .ZN(n8157) );
  NAND2_X1 U8345 ( .A1(n8149), .A2(n8157), .ZN(n6730) );
  XNOR2_X1 U8346 ( .A(n8937), .B(n6753), .ZN(n6731) );
  XNOR2_X1 U8347 ( .A(n6731), .B(n8787), .ZN(n8158) );
  NAND2_X1 U8348 ( .A1(n6731), .A2(n8749), .ZN(n6732) );
  XNOR2_X1 U8349 ( .A(n8854), .B(n4513), .ZN(n6733) );
  XNOR2_X1 U8350 ( .A(n6733), .B(n8767), .ZN(n8210) );
  XNOR2_X1 U8351 ( .A(n8850), .B(n4513), .ZN(n6734) );
  XNOR2_X1 U8352 ( .A(n6734), .B(n8718), .ZN(n8127) );
  NAND2_X1 U8353 ( .A1(n8126), .A2(n8127), .ZN(n6736) );
  NAND2_X1 U8354 ( .A1(n6734), .A2(n8747), .ZN(n6735) );
  NAND2_X1 U8355 ( .A1(n6736), .A2(n6735), .ZN(n8183) );
  XNOR2_X1 U8356 ( .A(n8722), .B(n6753), .ZN(n6737) );
  XNOR2_X1 U8357 ( .A(n6737), .B(n8732), .ZN(n8184) );
  NAND2_X1 U8358 ( .A1(n8183), .A2(n8184), .ZN(n6739) );
  NAND2_X1 U8359 ( .A1(n6737), .A2(n8705), .ZN(n6738) );
  NAND2_X1 U8360 ( .A1(n6739), .A2(n6738), .ZN(n8133) );
  XNOR2_X1 U8361 ( .A(n8708), .B(n6753), .ZN(n6741) );
  XNOR2_X1 U8362 ( .A(n6741), .B(n8717), .ZN(n8134) );
  NAND2_X1 U8363 ( .A1(n8133), .A2(n8134), .ZN(n6743) );
  NAND2_X1 U8364 ( .A1(n6741), .A2(n6740), .ZN(n6742) );
  XNOR2_X1 U8365 ( .A(n8914), .B(n6753), .ZN(n6744) );
  XNOR2_X1 U8366 ( .A(n6744), .B(n8686), .ZN(n8202) );
  XNOR2_X1 U8367 ( .A(n8902), .B(n6753), .ZN(n8175) );
  XNOR2_X1 U8368 ( .A(n8908), .B(n6701), .ZN(n8171) );
  INV_X1 U8369 ( .A(n8171), .ZN(n6745) );
  OAI22_X1 U8370 ( .A1(n8175), .A2(n8174), .B1(n8205), .B2(n6745), .ZN(n6749)
         );
  OAI21_X1 U8371 ( .B1(n8171), .B2(n8696), .A(n8685), .ZN(n6747) );
  NOR2_X1 U8372 ( .A1(n8685), .A2(n8696), .ZN(n6746) );
  AOI22_X1 U8373 ( .A1(n6747), .A2(n8175), .B1(n6746), .B2(n6745), .ZN(n6748)
         );
  XNOR2_X1 U8374 ( .A(n8896), .B(n4513), .ZN(n6750) );
  XNOR2_X1 U8375 ( .A(n6750), .B(n8671), .ZN(n8142) );
  XNOR2_X1 U8376 ( .A(n8890), .B(n4513), .ZN(n6751) );
  NOR2_X1 U8377 ( .A1(n6751), .A2(n8635), .ZN(n8219) );
  NAND2_X1 U8378 ( .A1(n6751), .A2(n8635), .ZN(n8217) );
  XNOR2_X1 U8379 ( .A(n8884), .B(n6753), .ZN(n6752) );
  XNOR2_X1 U8380 ( .A(n6752), .B(n8624), .ZN(n8104) );
  XOR2_X1 U8381 ( .A(n4513), .B(n8622), .Z(n6754) );
  XNOR2_X1 U8382 ( .A(n6755), .B(n6754), .ZN(n6761) );
  INV_X1 U8383 ( .A(n6756), .ZN(n6757) );
  NAND2_X1 U8384 ( .A1(n6757), .A2(n6762), .ZN(n6760) );
  INV_X1 U8385 ( .A(n6769), .ZN(n6758) );
  NAND2_X1 U8386 ( .A1(n6781), .A2(n6758), .ZN(n6759) );
  NAND2_X1 U8387 ( .A1(n6761), .A2(n8232), .ZN(n6791) );
  NAND2_X1 U8388 ( .A1(n6762), .A2(n10046), .ZN(n6764) );
  INV_X1 U8389 ( .A(n6857), .ZN(n6774) );
  NOR2_X1 U8390 ( .A1(n10041), .A2(n6774), .ZN(n6763) );
  INV_X1 U8391 ( .A(n6765), .ZN(n6766) );
  NAND2_X1 U8392 ( .A1(n6767), .A2(n6766), .ZN(n6772) );
  OAI211_X1 U8393 ( .C1(n6769), .C2(n6775), .A(n6947), .B(n6798), .ZN(n6770)
         );
  INV_X1 U8394 ( .A(n6770), .ZN(n6771) );
  NAND2_X1 U8395 ( .A1(n6772), .A2(n6771), .ZN(n6773) );
  NAND2_X1 U8396 ( .A1(n6773), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6778) );
  NOR2_X1 U8397 ( .A1(n6780), .A2(n6774), .ZN(n8461) );
  INV_X1 U8398 ( .A(n6775), .ZN(n6776) );
  NAND2_X1 U8399 ( .A1(n8461), .A2(n6776), .ZN(n6777) );
  NAND2_X1 U8400 ( .A1(n6778), .A2(n6777), .ZN(n6982) );
  OR2_X1 U8401 ( .A1(n6945), .A2(P2_U3151), .ZN(n8465) );
  INV_X1 U8402 ( .A(n8465), .ZN(n6779) );
  INV_X1 U8403 ( .A(n6780), .ZN(n7370) );
  NAND2_X1 U8404 ( .A1(n6781), .A2(n7370), .ZN(n6784) );
  INV_X1 U8405 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10349) );
  OAI22_X1 U8406 ( .A1(n8624), .A2(n8223), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10349), .ZN(n6786) );
  INV_X1 U8407 ( .A(n6782), .ZN(n6783) );
  NOR2_X1 U8408 ( .A1(n8625), .A2(n8238), .ZN(n6785) );
  AOI211_X1 U8409 ( .C1(n8629), .C2(n8241), .A(n6786), .B(n6785), .ZN(n6787)
         );
  NAND2_X1 U8410 ( .A1(n6791), .A2(n6790), .ZN(P2_U3160) );
  NAND3_X1 U8411 ( .A1(n8432), .A2(n8463), .A3(n8599), .ZN(n6792) );
  NAND2_X1 U8412 ( .A1(n8435), .A2(n6792), .ZN(n6793) );
  NAND2_X1 U8413 ( .A1(n6793), .A2(n7361), .ZN(n6794) );
  AND2_X1 U8414 ( .A1(n6796), .A2(n6857), .ZN(n6797) );
  OAI21_X1 U8415 ( .B1(n6679), .B2(n10041), .A(n6799), .ZN(n6800) );
  INV_X1 U8416 ( .A(n6800), .ZN(n6801) );
  OR2_X1 U8417 ( .A1(n6802), .A2(n10463), .ZN(n6807) );
  INV_X1 U8418 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6803) );
  INV_X1 U8419 ( .A(n6805), .ZN(n6806) );
  NAND2_X1 U8420 ( .A1(n6807), .A2(n6806), .ZN(P2_U3488) );
  INV_X1 U8421 ( .A(n6808), .ZN(n6809) );
  INV_X1 U8422 ( .A(n6863), .ZN(n6981) );
  NAND2_X1 U8423 ( .A1(n8435), .A2(n6947), .ZN(n6810) );
  NAND2_X1 U8424 ( .A1(n6810), .A2(n6945), .ZN(n6955) );
  NAND2_X1 U8425 ( .A1(n6955), .A2(n6266), .ZN(n6811) );
  NAND2_X1 U8426 ( .A1(n6811), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  AND2_X1 U8427 ( .A1(n6814), .A2(P1_U3086), .ZN(n7389) );
  NOR2_X1 U8428 ( .A1(n6814), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9625) );
  INV_X2 U8429 ( .A(n9625), .ZN(n9629) );
  OAI222_X1 U8430 ( .A1(n9633), .A2(n6812), .B1(n9629), .B2(n6818), .C1(
        P1_U3086), .C2(n6885), .ZN(P1_U3353) );
  INV_X2 U8431 ( .A(n7389), .ZN(n9633) );
  OAI222_X1 U8432 ( .A1(n9633), .A2(n6813), .B1(n9629), .B2(n6815), .C1(
        P1_U3086), .C2(n6883), .ZN(P1_U3354) );
  NOR2_X1 U8433 ( .A1(n6814), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8963) );
  INV_X2 U8434 ( .A(n8963), .ZN(n8102) );
  AND2_X1 U8435 ( .A1(n6814), .A2(P2_U3151), .ZN(n7913) );
  INV_X2 U8436 ( .A(n7913), .ZN(n8965) );
  OAI222_X1 U8437 ( .A1(n8102), .A2(n6816), .B1(n8965), .B2(n6815), .C1(
        P2_U3151), .C2(n7014), .ZN(P2_U3294) );
  OAI222_X1 U8438 ( .A1(n8102), .A2(n6817), .B1(n8965), .B2(n6820), .C1(
        P2_U3151), .C2(n7029), .ZN(P2_U3292) );
  OAI222_X1 U8439 ( .A1(n8102), .A2(n6819), .B1(n8965), .B2(n6818), .C1(
        P2_U3151), .C2(n7099), .ZN(P2_U3293) );
  OAI222_X1 U8440 ( .A1(n9633), .A2(n6821), .B1(n9629), .B2(n6820), .C1(
        P1_U3086), .C2(n9214), .ZN(P1_U3352) );
  OAI222_X1 U8441 ( .A1(n8102), .A2(n6822), .B1(n8965), .B2(n6823), .C1(
        P2_U3151), .C2(n7172), .ZN(P2_U3291) );
  OAI222_X1 U8442 ( .A1(n6824), .A2(n9633), .B1(P1_U3086), .B2(n6889), .C1(
        n9629), .C2(n6823), .ZN(P1_U3351) );
  OAI222_X1 U8443 ( .A1(n9633), .A2(n6826), .B1(n9629), .B2(n6827), .C1(
        P1_U3086), .C2(n6825), .ZN(P1_U3350) );
  OAI222_X1 U8444 ( .A1(n8102), .A2(n6828), .B1(n8965), .B2(n6827), .C1(
        P2_U3151), .C2(n7056), .ZN(P2_U3290) );
  INV_X1 U8445 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6829) );
  OAI222_X1 U8446 ( .A1(n8102), .A2(n6829), .B1(n8965), .B2(n6830), .C1(
        P2_U3151), .C2(n7061), .ZN(P2_U3289) );
  OAI222_X1 U8447 ( .A1(n9633), .A2(n6831), .B1(n9629), .B2(n6830), .C1(
        P1_U3086), .C2(n6875), .ZN(P1_U3349) );
  INV_X1 U8448 ( .A(n6832), .ZN(n6834) );
  INV_X1 U8449 ( .A(n6919), .ZN(n6876) );
  OAI222_X1 U8450 ( .A1(n9633), .A2(n6833), .B1(n9629), .B2(n6834), .C1(
        P1_U3086), .C2(n6876), .ZN(P1_U3348) );
  INV_X1 U8451 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6835) );
  OAI222_X1 U8452 ( .A1(n8102), .A2(n6835), .B1(n8965), .B2(n6834), .C1(
        P2_U3151), .C2(n4688), .ZN(P2_U3288) );
  INV_X1 U8453 ( .A(n6836), .ZN(n6838) );
  INV_X1 U8454 ( .A(n6968), .ZN(n6877) );
  OAI222_X1 U8455 ( .A1(n9633), .A2(n6837), .B1(n9629), .B2(n6838), .C1(
        P1_U3086), .C2(n6877), .ZN(P1_U3347) );
  OAI222_X1 U8456 ( .A1(n8102), .A2(n6839), .B1(n8965), .B2(n6838), .C1(
        P2_U3151), .C2(n7216), .ZN(P2_U3287) );
  INV_X1 U8457 ( .A(n6842), .ZN(n6840) );
  OR2_X1 U8458 ( .A1(n5960), .A2(n6840), .ZN(n6841) );
  NAND2_X1 U8459 ( .A1(n6841), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6880) );
  NAND2_X1 U8460 ( .A1(n6843), .A2(n6842), .ZN(n6844) );
  NAND2_X1 U8461 ( .A1(n6845), .A2(n6844), .ZN(n6879) );
  INV_X1 U8462 ( .A(n6879), .ZN(n6846) );
  INV_X1 U8463 ( .A(n9344), .ZN(n9715) );
  NOR2_X1 U8464 ( .A1(n9715), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8465 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6848) );
  NAND2_X1 U8466 ( .A1(n5974), .A2(P1_U3973), .ZN(n6847) );
  OAI21_X1 U8467 ( .B1(P1_U3973), .B2(n6848), .A(n6847), .ZN(P1_U3554) );
  INV_X1 U8468 ( .A(n6849), .ZN(n6852) );
  AOI22_X1 U8469 ( .A1(n9269), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n7389), .ZN(n6850) );
  OAI21_X1 U8470 ( .B1(n6852), .B2(n9629), .A(n6850), .ZN(P1_U3346) );
  INV_X1 U8471 ( .A(n7318), .ZN(n7326) );
  OAI222_X1 U8472 ( .A1(n8965), .A2(n6852), .B1(n7326), .B2(P2_U3151), .C1(
        n6851), .C2(n8102), .ZN(P2_U3286) );
  INV_X1 U8473 ( .A(n6853), .ZN(n6856) );
  AOI22_X1 U8474 ( .A1(n7139), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n7389), .ZN(n6854) );
  OAI21_X1 U8475 ( .B1(n6856), .B2(n9629), .A(n6854), .ZN(P1_U3345) );
  INV_X1 U8476 ( .A(n7338), .ZN(n7435) );
  INV_X1 U8477 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6855) );
  OAI222_X1 U8478 ( .A1(n8965), .A2(n6856), .B1(n7435), .B2(P2_U3151), .C1(
        n6855), .C2(n8102), .ZN(P2_U3285) );
  INV_X1 U8479 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6860) );
  INV_X1 U8480 ( .A(n6858), .ZN(n6859) );
  AOI22_X1 U8481 ( .A1(n6865), .A2(n6860), .B1(n6863), .B2(n6859), .ZN(
        P2_U3377) );
  INV_X1 U8482 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6864) );
  INV_X1 U8483 ( .A(n6861), .ZN(n6862) );
  AOI22_X1 U8484 ( .A1(n6865), .A2(n6864), .B1(n6863), .B2(n6862), .ZN(
        P2_U3376) );
  AND2_X1 U8485 ( .A1(n6865), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8486 ( .A1(n6865), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8487 ( .A1(n6865), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8488 ( .A1(n6865), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8489 ( .A1(n6865), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8490 ( .A1(n6865), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8491 ( .A1(n6865), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8492 ( .A1(n6865), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8493 ( .A1(n6865), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8494 ( .A1(n6865), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8495 ( .A1(n6865), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8496 ( .A1(n6865), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8497 ( .A1(n6865), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8498 ( .A1(n6865), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8499 ( .A1(n6865), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8500 ( .A1(n6865), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8501 ( .A1(n6865), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8502 ( .A1(n6865), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8503 ( .A1(n6865), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8504 ( .A1(n6865), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8505 ( .A1(n6865), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8506 ( .A1(n6865), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8507 ( .A1(n6865), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8508 ( .A1(n6865), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8509 ( .A1(n6865), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  INV_X1 U8510 ( .A(n6865), .ZN(n6867) );
  INV_X1 U8511 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n10306) );
  NOR2_X1 U8512 ( .A1(n6867), .A2(n10306), .ZN(P2_U3235) );
  INV_X1 U8513 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10098) );
  NOR2_X1 U8514 ( .A1(n6867), .A2(n10098), .ZN(P2_U3263) );
  INV_X1 U8515 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n10308) );
  NOR2_X1 U8516 ( .A1(n6867), .A2(n10308), .ZN(P2_U3246) );
  INV_X1 U8517 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6866) );
  NOR2_X1 U8518 ( .A1(n6867), .A2(n6866), .ZN(P2_U3260) );
  INV_X1 U8519 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10328) );
  NOR2_X1 U8520 ( .A1(n6867), .A2(n10328), .ZN(P2_U3254) );
  INV_X1 U8521 ( .A(n6868), .ZN(n6869) );
  INV_X1 U8522 ( .A(n7308), .ZN(n7140) );
  OAI222_X1 U8523 ( .A1(n9633), .A2(n10331), .B1(n9629), .B2(n6869), .C1(
        P1_U3086), .C2(n7140), .ZN(P1_U3344) );
  OAI222_X1 U8524 ( .A1(n8102), .A2(n6870), .B1(n8965), .B2(n6869), .C1(
        P2_U3151), .C2(n7564), .ZN(P2_U3284) );
  MUX2_X1 U8525 ( .A(n5615), .B(P1_REG2_REG_2__SCAN_IN), .S(n6885), .Z(n9722)
         );
  MUX2_X1 U8526 ( .A(n5605), .B(P1_REG2_REG_1__SCAN_IN), .S(n6883), .Z(n9207)
         );
  AND2_X1 U8527 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9228) );
  NAND2_X1 U8528 ( .A1(n9207), .A2(n9228), .ZN(n9206) );
  INV_X1 U8529 ( .A(n6883), .ZN(n9202) );
  NAND2_X1 U8530 ( .A1(n9202), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6871) );
  NAND2_X1 U8531 ( .A1(n9206), .A2(n6871), .ZN(n9721) );
  NAND2_X1 U8532 ( .A1(n9722), .A2(n9721), .ZN(n9719) );
  INV_X1 U8533 ( .A(n6885), .ZN(n9723) );
  NAND2_X1 U8534 ( .A1(n9723), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6872) );
  NAND2_X1 U8535 ( .A1(n9719), .A2(n6872), .ZN(n9220) );
  INV_X1 U8536 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7648) );
  MUX2_X1 U8537 ( .A(n7648), .B(P1_REG2_REG_3__SCAN_IN), .S(n9214), .Z(n9221)
         );
  NAND2_X1 U8538 ( .A1(n9220), .A2(n9221), .ZN(n9219) );
  OR2_X1 U8539 ( .A1(n9214), .A2(n7648), .ZN(n6873) );
  NAND2_X1 U8540 ( .A1(n9219), .A2(n6873), .ZN(n9241) );
  XNOR2_X1 U8541 ( .A(n6889), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9242) );
  NAND2_X1 U8542 ( .A1(n9241), .A2(n9242), .ZN(n9240) );
  INV_X1 U8543 ( .A(n6889), .ZN(n9236) );
  NAND2_X1 U8544 ( .A1(n9236), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6874) );
  NAND2_X1 U8545 ( .A1(n9240), .A2(n6874), .ZN(n9255) );
  MUX2_X1 U8546 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7689), .S(n9252), .Z(n9256)
         );
  AND2_X1 U8547 ( .A1(n9255), .A2(n9256), .ZN(n9253) );
  AOI22_X1 U8548 ( .A1(n6907), .A2(n5592), .B1(P1_REG2_REG_6__SCAN_IN), .B2(
        n6875), .ZN(n6902) );
  NOR2_X1 U8549 ( .A1(n6903), .A2(n6902), .ZN(n6901) );
  AOI22_X1 U8550 ( .A1(n6919), .A2(n7540), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n6876), .ZN(n6914) );
  NOR2_X1 U8551 ( .A1(n6915), .A2(n6914), .ZN(n6913) );
  INV_X1 U8552 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6878) );
  AOI22_X1 U8553 ( .A1(n6968), .A2(n6878), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n6877), .ZN(n6881) );
  NOR2_X1 U8554 ( .A1(n6882), .A2(n6881), .ZN(n6961) );
  OR2_X1 U8555 ( .A1(n6880), .A2(n6879), .ZN(n9713) );
  NOR2_X2 U8556 ( .A1(n9713), .A2(n9227), .ZN(n9720) );
  AOI211_X1 U8557 ( .C1(n6882), .C2(n6881), .A(n6961), .B(n9289), .ZN(n6900)
         );
  INV_X1 U8558 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6886) );
  MUX2_X1 U8559 ( .A(n6886), .B(P1_REG1_REG_2__SCAN_IN), .S(n6885), .Z(n9718)
         );
  INV_X1 U8560 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9920) );
  AND2_X1 U8561 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9204) );
  NAND2_X1 U8562 ( .A1(n9202), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6884) );
  NAND2_X1 U8563 ( .A1(n9203), .A2(n6884), .ZN(n9717) );
  NAND2_X1 U8564 ( .A1(n9718), .A2(n9717), .ZN(n9716) );
  OAI21_X1 U8565 ( .B1(n6886), .B2(n6885), .A(n9716), .ZN(n9212) );
  MUX2_X1 U8566 ( .A(n6887), .B(P1_REG1_REG_3__SCAN_IN), .S(n9214), .Z(n9213)
         );
  NAND2_X1 U8567 ( .A1(n9212), .A2(n9213), .ZN(n9211) );
  OAI21_X1 U8568 ( .B1(n6887), .B2(n9214), .A(n9211), .ZN(n9238) );
  XNOR2_X1 U8569 ( .A(n6889), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9239) );
  NAND2_X1 U8570 ( .A1(n9238), .A2(n9239), .ZN(n9237) );
  OAI21_X1 U8571 ( .B1(n6889), .B2(n6888), .A(n9237), .ZN(n9247) );
  INV_X1 U8572 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9925) );
  MUX2_X1 U8573 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9925), .S(n9252), .Z(n9248)
         );
  NAND2_X1 U8574 ( .A1(n9247), .A2(n9248), .ZN(n9246) );
  MUX2_X1 U8575 ( .A(n6890), .B(P1_REG1_REG_6__SCAN_IN), .S(n6907), .Z(n6905)
         );
  MUX2_X1 U8576 ( .A(n6891), .B(P1_REG1_REG_7__SCAN_IN), .S(n6919), .Z(n6917)
         );
  NOR2_X1 U8577 ( .A1(n6918), .A2(n6917), .ZN(n6916) );
  MUX2_X1 U8578 ( .A(n6892), .B(P1_REG1_REG_8__SCAN_IN), .S(n6968), .Z(n6894)
         );
  INV_X1 U8579 ( .A(n9713), .ZN(n6893) );
  NAND2_X1 U8580 ( .A1(n6893), .A2(n4511), .ZN(n9727) );
  AOI211_X1 U8581 ( .C1(n6895), .C2(n6894), .A(n6967), .B(n9727), .ZN(n6899)
         );
  INV_X1 U8582 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6897) );
  NOR2_X2 U8583 ( .A1(n9713), .A2(n9226), .ZN(n9724) );
  NAND2_X1 U8584 ( .A1(n9724), .A2(n6968), .ZN(n6896) );
  NAND2_X1 U8585 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7844) );
  OAI211_X1 U8586 ( .C1(n6897), .C2(n9344), .A(n6896), .B(n7844), .ZN(n6898)
         );
  OR3_X1 U8587 ( .A1(n6900), .A2(n6899), .A3(n6898), .ZN(P1_U3251) );
  AOI211_X1 U8588 ( .C1(n6903), .C2(n6902), .A(n6901), .B(n9289), .ZN(n6912)
         );
  AOI211_X1 U8589 ( .C1(n6906), .C2(n6905), .A(n6904), .B(n9727), .ZN(n6911)
         );
  INV_X1 U8590 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6909) );
  NAND2_X1 U8591 ( .A1(n9724), .A2(n6907), .ZN(n6908) );
  NAND2_X1 U8592 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9700) );
  OAI211_X1 U8593 ( .C1(n6909), .C2(n9344), .A(n6908), .B(n9700), .ZN(n6910)
         );
  OR3_X1 U8594 ( .A1(n6912), .A2(n6911), .A3(n6910), .ZN(P1_U3249) );
  AOI211_X1 U8595 ( .C1(n6915), .C2(n6914), .A(n6913), .B(n9289), .ZN(n6923)
         );
  AOI211_X1 U8596 ( .C1(n6918), .C2(n6917), .A(n6916), .B(n9727), .ZN(n6922)
         );
  INV_X1 U8597 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10305) );
  NAND2_X1 U8598 ( .A1(n9724), .A2(n6919), .ZN(n6920) );
  NAND2_X1 U8599 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n7731) );
  OAI211_X1 U8600 ( .C1(n10305), .C2(n9344), .A(n6920), .B(n7731), .ZN(n6921)
         );
  OR3_X1 U8601 ( .A1(n6923), .A2(n6922), .A3(n6921), .ZN(P1_U3250) );
  NOR2_X1 U8602 ( .A1(n7463), .A2(n9833), .ZN(n9831) );
  AND2_X1 U8603 ( .A1(n6925), .A2(n6924), .ZN(n7462) );
  AND2_X1 U8604 ( .A1(n7462), .A2(n6926), .ZN(n6927) );
  INV_X1 U8605 ( .A(n9620), .ZN(n7465) );
  INV_X1 U8606 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6937) );
  AOI21_X1 U8607 ( .B1(n6929), .B2(n6928), .A(n7472), .ZN(n6930) );
  NAND2_X1 U8608 ( .A1(n6930), .A2(n7675), .ZN(n9872) );
  NAND2_X1 U8609 ( .A1(n5883), .A2(n6931), .ZN(n6933) );
  OAI21_X1 U8610 ( .B1(n9916), .B2(n9782), .A(n7676), .ZN(n6934) );
  NAND2_X1 U8611 ( .A1(n5979), .A2(n4509), .ZN(n7677) );
  OAI211_X1 U8612 ( .C1(n7674), .C2(n6935), .A(n6934), .B(n7677), .ZN(n9604)
         );
  NAND2_X1 U8613 ( .A1(n9604), .A2(n9919), .ZN(n6936) );
  OAI21_X1 U8614 ( .B1(n9919), .B2(n6937), .A(n6936), .ZN(P1_U3453) );
  INV_X1 U8615 ( .A(n6938), .ZN(n6939) );
  OAI222_X1 U8616 ( .A1(n8965), .A2(n6939), .B1(n8484), .B2(P2_U3151), .C1(
        n10343), .C2(n8102), .ZN(P2_U3283) );
  INV_X1 U8617 ( .A(n7423), .ZN(n7312) );
  OAI222_X1 U8618 ( .A1(n9633), .A2(n6940), .B1(n9629), .B2(n6939), .C1(n7312), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8619 ( .A(n6941), .ZN(n6943) );
  AOI22_X1 U8620 ( .A1(n7623), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n7389), .ZN(n6942) );
  OAI21_X1 U8621 ( .B1(n6943), .B2(n9629), .A(n6942), .ZN(P1_U3342) );
  INV_X1 U8622 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6944) );
  INV_X1 U8623 ( .A(n9938), .ZN(n8496) );
  OAI222_X1 U8624 ( .A1(n8102), .A2(n6944), .B1(n8965), .B2(n6943), .C1(
        P2_U3151), .C2(n8496), .ZN(P2_U3282) );
  INV_X1 U8625 ( .A(n6945), .ZN(n6946) );
  NOR2_X1 U8626 ( .A1(n6947), .A2(n6946), .ZN(n6948) );
  INV_X1 U8627 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6959) );
  NOR2_X1 U8628 ( .A1(n6625), .A2(P2_U3151), .ZN(n8959) );
  INV_X1 U8629 ( .A(n7012), .ZN(n6994) );
  INV_X1 U8630 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6950) );
  INV_X1 U8631 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6949) );
  INV_X2 U8632 ( .A(n8591), .ZN(n8540) );
  MUX2_X1 U8633 ( .A(n6950), .B(n6949), .S(n8540), .Z(n6951) );
  NAND2_X1 U8634 ( .A1(n6951), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7122) );
  INV_X1 U8635 ( .A(n6951), .ZN(n6952) );
  INV_X1 U8636 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7015) );
  NAND2_X1 U8637 ( .A1(n6952), .A2(n7015), .ZN(n6953) );
  AOI22_X1 U8638 ( .A1(n6994), .A2(n9981), .B1(n7122), .B2(n6953), .ZN(n6954)
         );
  AOI21_X1 U8639 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n6954), .ZN(
        n6958) );
  NOR2_X1 U8640 ( .A1(n8540), .A2(P2_U3151), .ZN(n8962) );
  AND2_X1 U8641 ( .A1(n6955), .A2(n8962), .ZN(n6956) );
  MUX2_X1 U8642 ( .A(P2_U3893), .B(n6956), .S(n6625), .Z(n9937) );
  NAND2_X1 U8643 ( .A1(n9937), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6957) );
  OAI211_X1 U8644 ( .C1(n8515), .C2(n6959), .A(n6958), .B(n6957), .ZN(P2_U3182) );
  NOR2_X1 U8645 ( .A1(n9269), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6960) );
  AOI21_X1 U8646 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n9269), .A(n6960), .ZN(
        n9262) );
  NAND2_X1 U8647 ( .A1(n9262), .A2(n9261), .ZN(n9260) );
  OAI21_X1 U8648 ( .B1(n9269), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9260), .ZN(
        n6964) );
  MUX2_X1 U8649 ( .A(n6962), .B(P1_REG2_REG_10__SCAN_IN), .S(n7139), .Z(n6963)
         );
  NOR2_X1 U8650 ( .A1(n6964), .A2(n6963), .ZN(n7138) );
  AOI211_X1 U8651 ( .C1(n6964), .C2(n6963), .A(n9289), .B(n7138), .ZN(n6975)
         );
  MUX2_X1 U8652 ( .A(n6965), .B(P1_REG1_REG_10__SCAN_IN), .S(n7139), .Z(n6970)
         );
  NOR2_X1 U8653 ( .A1(n9269), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6966) );
  AOI21_X1 U8654 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9269), .A(n6966), .ZN(
        n9267) );
  OAI21_X1 U8655 ( .B1(n9269), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9265), .ZN(
        n6969) );
  NOR2_X1 U8656 ( .A1(n6969), .A2(n6970), .ZN(n7134) );
  AOI211_X1 U8657 ( .C1(n6970), .C2(n6969), .A(n9727), .B(n7134), .ZN(n6974)
         );
  INV_X1 U8658 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6972) );
  NAND2_X1 U8659 ( .A1(n9724), .A2(n7139), .ZN(n6971) );
  NAND2_X1 U8660 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9638) );
  OAI211_X1 U8661 ( .C1(n6972), .C2(n9344), .A(n6971), .B(n9638), .ZN(n6973)
         );
  OR3_X1 U8662 ( .A1(n6975), .A2(n6974), .A3(n6973), .ZN(P1_U3253) );
  INV_X1 U8663 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6977) );
  INV_X1 U8664 ( .A(n6976), .ZN(n6979) );
  OAI222_X1 U8665 ( .A1(n8102), .A2(n6977), .B1(n8965), .B2(n6979), .C1(
        P2_U3151), .C2(n9971), .ZN(P2_U3281) );
  INV_X1 U8666 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10371) );
  INV_X1 U8667 ( .A(n7855), .ZN(n6978) );
  OAI222_X1 U8668 ( .A1(n9633), .A2(n10371), .B1(n9629), .B2(n6979), .C1(
        P1_U3086), .C2(n6978), .ZN(P1_U3341) );
  INV_X1 U8669 ( .A(n6980), .ZN(n7174) );
  NAND2_X1 U8670 ( .A1(n8482), .A2(n7119), .ZN(n8291) );
  INV_X1 U8671 ( .A(n8291), .ZN(n8295) );
  NOR2_X1 U8672 ( .A1(n7174), .A2(n8295), .ZN(n8265) );
  INV_X1 U8673 ( .A(n8265), .ZN(n7116) );
  AOI22_X1 U8674 ( .A1(n8227), .A2(n7369), .B1(n8232), .B2(n7116), .ZN(n6984)
         );
  OR2_X1 U8675 ( .A1(n6982), .A2(n6981), .ZN(n7243) );
  NAND2_X1 U8676 ( .A1(n7243), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6983) );
  OAI211_X1 U8677 ( .C1(n6574), .C2(n8238), .A(n6984), .B(n6983), .ZN(P2_U3172) );
  INV_X1 U8678 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6986) );
  INV_X1 U8679 ( .A(n6985), .ZN(n6987) );
  INV_X1 U8680 ( .A(n8522), .ZN(n8532) );
  OAI222_X1 U8681 ( .A1(n8102), .A2(n6986), .B1(n8965), .B2(n6987), .C1(
        P2_U3151), .C2(n8532), .ZN(P2_U3280) );
  INV_X1 U8682 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10326) );
  INV_X1 U8683 ( .A(n7857), .ZN(n9283) );
  OAI222_X1 U8684 ( .A1(n9633), .A2(n10326), .B1(n9629), .B2(n6987), .C1(
        P1_U3086), .C2(n9283), .ZN(P1_U3340) );
  XOR2_X1 U8685 ( .A(n6989), .B(n6988), .Z(n6993) );
  OAI22_X1 U8686 ( .A1(n8245), .A2(n7265), .B1(n8238), .B2(n4878), .ZN(n6990)
         );
  AOI21_X1 U8687 ( .B1(n8236), .B2(n8482), .A(n6990), .ZN(n6992) );
  NAND2_X1 U8688 ( .A1(n7243), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6991) );
  OAI211_X1 U8689 ( .C1(n6993), .C2(n8230), .A(n6992), .B(n6991), .ZN(P2_U3162) );
  INV_X1 U8690 ( .A(n9986), .ZN(n8562) );
  INV_X1 U8691 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6995) );
  AND2_X1 U8692 ( .A1(n7015), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6996) );
  NAND2_X1 U8693 ( .A1(n6262), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6997) );
  OAI21_X1 U8694 ( .B1(n7014), .B2(n6996), .A(n6997), .ZN(n7125) );
  INV_X1 U8695 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7457) );
  NAND2_X1 U8696 ( .A1(n7099), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6998) );
  INV_X1 U8697 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10339) );
  OAI21_X1 U8698 ( .B1(n4619), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7153), .ZN(
        n7026) );
  INV_X1 U8699 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7011) );
  MUX2_X1 U8700 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8540), .Z(n7000) );
  INV_X1 U8701 ( .A(n7014), .ZN(n7131) );
  XNOR2_X1 U8702 ( .A(n7000), .B(n7131), .ZN(n7123) );
  NAND2_X1 U8703 ( .A1(n7123), .A2(n7122), .ZN(n7002) );
  NAND2_X1 U8704 ( .A1(n7000), .A2(n7014), .ZN(n7001) );
  NAND2_X1 U8705 ( .A1(n7002), .A2(n7001), .ZN(n7088) );
  MUX2_X1 U8706 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8540), .Z(n7004) );
  INV_X1 U8707 ( .A(n7099), .ZN(n7003) );
  XNOR2_X1 U8708 ( .A(n7004), .B(n7003), .ZN(n7087) );
  NAND2_X1 U8709 ( .A1(n7088), .A2(n7087), .ZN(n7006) );
  NAND2_X1 U8710 ( .A1(n7004), .A2(n7099), .ZN(n7005) );
  NAND2_X1 U8711 ( .A1(n7006), .A2(n7005), .ZN(n7008) );
  MUX2_X1 U8712 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8540), .Z(n7050) );
  XNOR2_X1 U8713 ( .A(n7050), .B(n7029), .ZN(n7007) );
  OR2_X1 U8714 ( .A1(n7008), .A2(n7007), .ZN(n7166) );
  NAND2_X1 U8715 ( .A1(n7008), .A2(n7007), .ZN(n7009) );
  AND2_X1 U8716 ( .A1(n7166), .A2(n7009), .ZN(n7010) );
  OAI22_X1 U8717 ( .A1(n8515), .A2(n7011), .B1(n7010), .B2(n9981), .ZN(n7025)
         );
  INV_X1 U8718 ( .A(n9991), .ZN(n8582) );
  INV_X1 U8719 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7013) );
  MUX2_X1 U8720 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n7013), .S(n7099), .Z(n7092)
         );
  NAND2_X1 U8721 ( .A1(n6262), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7019) );
  NAND2_X1 U8722 ( .A1(n7014), .A2(n7019), .ZN(n7018) );
  NAND2_X1 U8723 ( .A1(n7015), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7016) );
  OR2_X1 U8724 ( .A1(n7016), .A2(n6262), .ZN(n7017) );
  NAND2_X1 U8725 ( .A1(n7018), .A2(n7017), .ZN(n7121) );
  NAND2_X1 U8726 ( .A1(n7121), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7020) );
  NAND2_X1 U8727 ( .A1(n7020), .A2(n7019), .ZN(n7091) );
  NAND2_X1 U8728 ( .A1(n7092), .A2(n7091), .ZN(n7090) );
  NAND2_X1 U8729 ( .A1(n7099), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7021) );
  NAND2_X1 U8730 ( .A1(n7090), .A2(n7021), .ZN(n7030) );
  INV_X1 U8731 ( .A(n7029), .ZN(n7051) );
  XNOR2_X1 U8732 ( .A(n7030), .B(n7051), .ZN(n7028) );
  XOR2_X1 U8733 ( .A(n7028), .B(P2_REG1_REG_3__SCAN_IN), .Z(n7023) );
  OR2_X1 U8734 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7022), .ZN(n7250) );
  OAI21_X1 U8735 ( .B1(n8582), .B2(n7023), .A(n7250), .ZN(n7024) );
  AOI211_X1 U8736 ( .C1(n8562), .C2(n7026), .A(n7025), .B(n7024), .ZN(n7027)
         );
  OAI21_X1 U8737 ( .B1(n7029), .B2(n9995), .A(n7027), .ZN(P2_U3185) );
  INV_X1 U8738 ( .A(n7172), .ZN(n7049) );
  INV_X1 U8739 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10464) );
  NAND2_X1 U8740 ( .A1(n7028), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7032) );
  NAND2_X1 U8741 ( .A1(n7030), .A2(n7029), .ZN(n7031) );
  NAND2_X1 U8742 ( .A1(n7032), .A2(n7031), .ZN(n7158) );
  MUX2_X1 U8743 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10464), .S(n7172), .Z(n7159)
         );
  NAND2_X1 U8744 ( .A1(n7158), .A2(n7159), .ZN(n7157) );
  INV_X1 U8745 ( .A(n7056), .ZN(n7279) );
  XNOR2_X1 U8746 ( .A(n7033), .B(n7279), .ZN(n7273) );
  AOI22_X1 U8747 ( .A1(n7273), .A2(P2_REG1_REG_5__SCAN_IN), .B1(n7056), .B2(
        n7033), .ZN(n7286) );
  INV_X1 U8748 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10055) );
  MUX2_X1 U8749 ( .A(n10055), .B(P2_REG1_REG_6__SCAN_IN), .S(n7061), .Z(n7287)
         );
  NOR2_X1 U8750 ( .A1(n7286), .A2(n7287), .ZN(n7285) );
  AOI21_X1 U8751 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n7061), .A(n7285), .ZN(
        n7034) );
  INV_X1 U8752 ( .A(n7034), .ZN(n7201) );
  XNOR2_X1 U8753 ( .A(n7201), .B(n7065), .ZN(n7035) );
  OAI21_X1 U8754 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n7035), .A(n7202), .ZN(
        n7048) );
  INV_X1 U8755 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7598) );
  MUX2_X1 U8756 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7598), .S(n7172), .Z(n7150)
         );
  NAND2_X1 U8757 ( .A1(n7036), .A2(n7150), .ZN(n7155) );
  NAND2_X1 U8758 ( .A1(n7172), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7037) );
  NAND2_X1 U8759 ( .A1(n7155), .A2(n7037), .ZN(n7038) );
  OR2_X1 U8760 ( .A1(n7038), .A2(n7056), .ZN(n7039) );
  NAND2_X1 U8761 ( .A1(n7038), .A2(n7056), .ZN(n7288) );
  AND2_X1 U8762 ( .A1(n7039), .A2(n7288), .ZN(n7271) );
  XNOR2_X1 U8763 ( .A(n7061), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n7289) );
  INV_X1 U8764 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7043) );
  AOI21_X1 U8765 ( .B1(n7044), .B2(n7043), .A(n7191), .ZN(n7046) );
  INV_X1 U8766 ( .A(n8515), .ZN(n9973) );
  AND2_X1 U8767 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7699) );
  AOI21_X1 U8768 ( .B1(n9973), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7699), .ZN(
        n7045) );
  OAI21_X1 U8769 ( .B1(n7046), .B2(n9986), .A(n7045), .ZN(n7047) );
  AOI21_X1 U8770 ( .B1(n9991), .B2(n7048), .A(n7047), .ZN(n7077) );
  MUX2_X1 U8771 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8540), .Z(n7054) );
  XNOR2_X1 U8772 ( .A(n7054), .B(n7049), .ZN(n7168) );
  INV_X1 U8773 ( .A(n7050), .ZN(n7052) );
  NAND2_X1 U8774 ( .A1(n7052), .A2(n7051), .ZN(n7165) );
  AND2_X1 U8775 ( .A1(n7168), .A2(n7165), .ZN(n7053) );
  NAND2_X1 U8776 ( .A1(n7166), .A2(n7053), .ZN(n7167) );
  NAND2_X1 U8777 ( .A1(n7054), .A2(n7172), .ZN(n7055) );
  NAND2_X1 U8778 ( .A1(n7167), .A2(n7055), .ZN(n7270) );
  MUX2_X1 U8779 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8540), .Z(n7057) );
  XNOR2_X1 U8780 ( .A(n7057), .B(n7279), .ZN(n7269) );
  NAND2_X1 U8781 ( .A1(n7270), .A2(n7269), .ZN(n7059) );
  NAND2_X1 U8782 ( .A1(n7057), .A2(n7056), .ZN(n7058) );
  NAND2_X1 U8783 ( .A1(n7059), .A2(n7058), .ZN(n7283) );
  MUX2_X1 U8784 ( .A(n4690), .B(n10055), .S(n8540), .Z(n7060) );
  NAND2_X1 U8785 ( .A1(n7060), .A2(n4691), .ZN(n7070) );
  INV_X1 U8786 ( .A(n7060), .ZN(n7062) );
  NAND2_X1 U8787 ( .A1(n7062), .A2(n7061), .ZN(n7063) );
  NAND2_X1 U8788 ( .A1(n7070), .A2(n7063), .ZN(n7284) );
  OR2_X1 U8789 ( .A1(n7283), .A2(n7284), .ZN(n7071) );
  INV_X1 U8790 ( .A(n7071), .ZN(n7282) );
  INV_X1 U8791 ( .A(n7070), .ZN(n7069) );
  INV_X1 U8792 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7064) );
  MUX2_X1 U8793 ( .A(n7043), .B(n7064), .S(n8540), .Z(n7066) );
  NAND2_X1 U8794 ( .A1(n7066), .A2(n7065), .ZN(n7186) );
  INV_X1 U8795 ( .A(n7066), .ZN(n7067) );
  NAND2_X1 U8796 ( .A1(n7067), .A2(n4688), .ZN(n7068) );
  AND2_X1 U8797 ( .A1(n7186), .A2(n7068), .ZN(n7072) );
  NOR3_X1 U8798 ( .A1(n7282), .A2(n7069), .A3(n7072), .ZN(n7075) );
  NAND2_X1 U8799 ( .A1(n7071), .A2(n7070), .ZN(n7073) );
  NAND2_X1 U8800 ( .A1(n7073), .A2(n7072), .ZN(n7189) );
  INV_X1 U8801 ( .A(n7189), .ZN(n7074) );
  INV_X1 U8802 ( .A(n9981), .ZN(n7348) );
  OAI21_X1 U8803 ( .B1(n7075), .B2(n7074), .A(n7348), .ZN(n7076) );
  OAI211_X1 U8804 ( .C1(n9995), .C2(n4688), .A(n7077), .B(n7076), .ZN(P2_U3189) );
  OAI21_X1 U8805 ( .B1(n7080), .B2(n7079), .A(n7078), .ZN(n9225) );
  NOR2_X1 U8806 ( .A1(n7081), .A2(n9833), .ZN(n7111) );
  OAI22_X1 U8807 ( .A1(n7111), .A2(n7679), .B1(n9153), .B2(n7677), .ZN(n7082)
         );
  AOI21_X1 U8808 ( .B1(n7673), .B2(n6200), .A(n7082), .ZN(n7083) );
  OAI21_X1 U8809 ( .B1(n9693), .B2(n9225), .A(n7083), .ZN(P1_U3232) );
  OAI21_X1 U8810 ( .B1(n7086), .B2(n7085), .A(n7084), .ZN(n7097) );
  INV_X1 U8811 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10314) );
  XNOR2_X1 U8812 ( .A(n7088), .B(n7087), .ZN(n7089) );
  OAI22_X1 U8813 ( .A1(n8515), .A2(n10314), .B1(n9981), .B2(n7089), .ZN(n7096)
         );
  OAI21_X1 U8814 ( .B1(n7092), .B2(n7091), .A(n7090), .ZN(n7093) );
  AOI22_X1 U8815 ( .A1(n9991), .A2(n7093), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n7094) );
  INV_X1 U8816 ( .A(n7094), .ZN(n7095) );
  AOI211_X1 U8817 ( .C1(n8562), .C2(n7097), .A(n7096), .B(n7095), .ZN(n7098)
         );
  OAI21_X1 U8818 ( .B1(n7099), .B2(n9995), .A(n7098), .ZN(P2_U3184) );
  XNOR2_X1 U8819 ( .A(n7101), .B(n7102), .ZN(n7103) );
  XOR2_X1 U8820 ( .A(n7100), .B(n7103), .Z(n7106) );
  AOI22_X1 U8821 ( .A1(n4509), .A2(n9197), .B1(n5974), .B2(n9131), .ZN(n7546)
         );
  OAI22_X1 U8822 ( .A1(n7111), .A2(n9199), .B1(n9153), .B2(n7546), .ZN(n7104)
         );
  AOI21_X1 U8823 ( .B1(n9835), .B2(n6200), .A(n7104), .ZN(n7105) );
  OAI21_X1 U8824 ( .B1(n7106), .B2(n9693), .A(n7105), .ZN(P1_U3222) );
  INV_X1 U8825 ( .A(n7108), .ZN(n7109) );
  AOI21_X1 U8826 ( .B1(n7107), .B2(n7110), .A(n7109), .ZN(n7115) );
  AOI22_X1 U8827 ( .A1(n9131), .A2(n5979), .B1(n9196), .B2(n4509), .ZN(n7482)
         );
  OAI22_X1 U8828 ( .A1(n7111), .A2(n7476), .B1(n9153), .B2(n7482), .ZN(n7112)
         );
  AOI21_X1 U8829 ( .B1(n7113), .B2(n6200), .A(n7112), .ZN(n7114) );
  OAI21_X1 U8830 ( .B1(n7115), .B2(n9693), .A(n7114), .ZN(P1_U3237) );
  OAI21_X1 U8831 ( .B1(n10021), .B2(n8805), .A(n7116), .ZN(n7118) );
  AND2_X1 U8832 ( .A1(n8800), .A2(n6572), .ZN(n7372) );
  INV_X1 U8833 ( .A(n7372), .ZN(n7117) );
  OAI211_X1 U8834 ( .C1(n7119), .C2(n10029), .A(n7118), .B(n7117), .ZN(n8868)
         );
  NAND2_X1 U8835 ( .A1(n10047), .A2(n8868), .ZN(n7120) );
  OAI21_X1 U8836 ( .B1(n10047), .B2(n6242), .A(n7120), .ZN(P2_U3390) );
  INV_X1 U8837 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10065) );
  XNOR2_X1 U8838 ( .A(n7121), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n7130) );
  XNOR2_X1 U8839 ( .A(n7123), .B(n7122), .ZN(n7124) );
  OAI22_X1 U8840 ( .A1(n9981), .A2(n7124), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6255), .ZN(n7129) );
  NAND2_X1 U8841 ( .A1(n7125), .A2(n7457), .ZN(n7126) );
  AOI21_X1 U8842 ( .B1(n7127), .B2(n7126), .A(n9986), .ZN(n7128) );
  AOI211_X1 U8843 ( .C1(n9991), .C2(n7130), .A(n7129), .B(n7128), .ZN(n7133)
         );
  NAND2_X1 U8844 ( .A1(n9937), .A2(n7131), .ZN(n7132) );
  OAI211_X1 U8845 ( .C1(n10065), .C2(n8515), .A(n7133), .B(n7132), .ZN(
        P2_U3183) );
  MUX2_X1 U8846 ( .A(n7135), .B(P1_REG1_REG_11__SCAN_IN), .S(n7308), .Z(n7136)
         );
  AOI211_X1 U8847 ( .C1(n7137), .C2(n7136), .A(n9727), .B(n7307), .ZN(n7147)
         );
  AOI22_X1 U8848 ( .A1(n7308), .A2(n7794), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n7140), .ZN(n7141) );
  NOR2_X1 U8849 ( .A1(n7142), .A2(n7141), .ZN(n7303) );
  AOI211_X1 U8850 ( .C1(n7142), .C2(n7141), .A(n7303), .B(n9289), .ZN(n7146)
         );
  INV_X1 U8851 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10350) );
  NAND2_X1 U8852 ( .A1(n9724), .A2(n7308), .ZN(n7144) );
  NAND2_X1 U8853 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n7143) );
  OAI211_X1 U8854 ( .C1(n10350), .C2(n9344), .A(n7144), .B(n7143), .ZN(n7145)
         );
  OR3_X1 U8855 ( .A1(n7147), .A2(n7146), .A3(n7145), .ZN(P1_U3254) );
  INV_X1 U8856 ( .A(n7148), .ZN(n7181) );
  OAI222_X1 U8857 ( .A1(n8965), .A2(n7181), .B1(n9994), .B2(P2_U3151), .C1(
        n7149), .C2(n8102), .ZN(P2_U3279) );
  INV_X1 U8858 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7163) );
  INV_X1 U8859 ( .A(n7150), .ZN(n7152) );
  NAND3_X1 U8860 ( .A1(n7153), .A2(n7152), .A3(n7151), .ZN(n7154) );
  NAND2_X1 U8861 ( .A1(n7155), .A2(n7154), .ZN(n7156) );
  INV_X1 U8862 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10235) );
  NOR2_X1 U8863 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10235), .ZN(n7382) );
  AOI21_X1 U8864 ( .B1(n8562), .B2(n7156), .A(n7382), .ZN(n7162) );
  OAI21_X1 U8865 ( .B1(n7159), .B2(n7158), .A(n7157), .ZN(n7160) );
  NAND2_X1 U8866 ( .A1(n9991), .A2(n7160), .ZN(n7161) );
  OAI211_X1 U8867 ( .C1(n7163), .C2(n8515), .A(n7162), .B(n7161), .ZN(n7164)
         );
  INV_X1 U8868 ( .A(n7164), .ZN(n7171) );
  AND2_X1 U8869 ( .A1(n7166), .A2(n7165), .ZN(n7169) );
  OAI211_X1 U8870 ( .C1(n7169), .C2(n7168), .A(n7348), .B(n7167), .ZN(n7170)
         );
  OAI211_X1 U8871 ( .C1(n9995), .C2(n7172), .A(n7171), .B(n7170), .ZN(P2_U3186) );
  INV_X1 U8872 ( .A(n10021), .ZN(n10031) );
  XNOR2_X1 U8873 ( .A(n7173), .B(n7174), .ZN(n7461) );
  XNOR2_X1 U8874 ( .A(n7175), .B(n7173), .ZN(n7176) );
  AOI222_X1 U8875 ( .A1(n8805), .A2(n7176), .B1(n8482), .B2(n8801), .C1(n8481), 
        .C2(n8800), .ZN(n7458) );
  OAI21_X1 U8876 ( .B1(n10031), .B2(n7461), .A(n7458), .ZN(n7267) );
  INV_X1 U8877 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7177) );
  OAI22_X1 U8878 ( .A1(n8867), .A2(n7265), .B1(n10466), .B2(n7177), .ZN(n7178)
         );
  AOI21_X1 U8879 ( .B1(n7267), .B2(n10466), .A(n7178), .ZN(n7179) );
  INV_X1 U8880 ( .A(n7179), .ZN(P2_U3460) );
  INV_X1 U8881 ( .A(n9305), .ZN(n9282) );
  OAI222_X1 U8882 ( .A1(P1_U3086), .A2(n9282), .B1(n9629), .B2(n7181), .C1(
        n7180), .C2(n9633), .ZN(P1_U3339) );
  INV_X1 U8883 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7637) );
  INV_X1 U8884 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7205) );
  MUX2_X1 U8885 ( .A(n7637), .B(n7205), .S(n8540), .Z(n7182) );
  NAND2_X1 U8886 ( .A1(n7182), .A2(n7204), .ZN(n7231) );
  INV_X1 U8887 ( .A(n7182), .ZN(n7183) );
  NAND2_X1 U8888 ( .A1(n7183), .A2(n7216), .ZN(n7184) );
  AND2_X1 U8889 ( .A1(n7231), .A2(n7184), .ZN(n7187) );
  INV_X1 U8890 ( .A(n7186), .ZN(n7185) );
  NOR2_X1 U8891 ( .A1(n7187), .A2(n7185), .ZN(n7190) );
  NAND2_X1 U8892 ( .A1(n7189), .A2(n7186), .ZN(n7188) );
  NAND2_X1 U8893 ( .A1(n7188), .A2(n7187), .ZN(n7232) );
  INV_X1 U8894 ( .A(n7232), .ZN(n7230) );
  AOI21_X1 U8895 ( .B1(n7190), .B2(n7189), .A(n7230), .ZN(n7211) );
  NAND2_X1 U8896 ( .A1(n7216), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7212) );
  OAI21_X1 U8897 ( .B1(n7216), .B2(P2_REG2_REG_8__SCAN_IN), .A(n7212), .ZN(
        n7193) );
  AOI21_X1 U8898 ( .B1(n7194), .B2(n7193), .A(n7213), .ZN(n7197) );
  NOR2_X1 U8899 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7195), .ZN(n7766) );
  INV_X1 U8900 ( .A(n7766), .ZN(n7196) );
  OAI21_X1 U8901 ( .B1(n9986), .B2(n7197), .A(n7196), .ZN(n7200) );
  INV_X1 U8902 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7198) );
  NOR2_X1 U8903 ( .A1(n8515), .A2(n7198), .ZN(n7199) );
  AOI211_X1 U8904 ( .C1(n9937), .C2(n7204), .A(n7200), .B(n7199), .ZN(n7210)
         );
  NAND2_X1 U8905 ( .A1(n4688), .A2(n7201), .ZN(n7203) );
  MUX2_X1 U8906 ( .A(n7205), .B(P2_REG1_REG_8__SCAN_IN), .S(n7204), .Z(n7206)
         );
  NAND2_X1 U8907 ( .A1(n7206), .A2(n7207), .ZN(n7217) );
  OAI21_X1 U8908 ( .B1(n7207), .B2(n7206), .A(n7217), .ZN(n7208) );
  NAND2_X1 U8909 ( .A1(n7208), .A2(n9991), .ZN(n7209) );
  OAI211_X1 U8910 ( .C1(n7211), .C2(n9981), .A(n7210), .B(n7209), .ZN(P2_U3190) );
  INV_X1 U8911 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7215) );
  XNOR2_X1 U8912 ( .A(n7318), .B(n7317), .ZN(n7214) );
  NOR2_X1 U8913 ( .A1(n7215), .A2(n7214), .ZN(n7320) );
  AOI21_X1 U8914 ( .B1(n7215), .B2(n7214), .A(n7320), .ZN(n7238) );
  NAND2_X1 U8915 ( .A1(n7216), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7218) );
  NAND2_X1 U8916 ( .A1(n7218), .A2(n7217), .ZN(n7325) );
  XOR2_X1 U8917 ( .A(n7326), .B(n7325), .Z(n7219) );
  OAI21_X1 U8918 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n7219), .A(n7327), .ZN(
        n7224) );
  INV_X1 U8919 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7222) );
  NAND2_X1 U8920 ( .A1(n9937), .A2(n7318), .ZN(n7221) );
  AND2_X1 U8921 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7917) );
  INV_X1 U8922 ( .A(n7917), .ZN(n7220) );
  OAI211_X1 U8923 ( .C1(n7222), .C2(n8515), .A(n7221), .B(n7220), .ZN(n7223)
         );
  AOI21_X1 U8924 ( .B1(n7224), .B2(n9991), .A(n7223), .ZN(n7237) );
  INV_X1 U8925 ( .A(n7231), .ZN(n7229) );
  INV_X1 U8926 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7225) );
  MUX2_X1 U8927 ( .A(n7215), .B(n7225), .S(n8540), .Z(n7226) );
  NAND2_X1 U8928 ( .A1(n7226), .A2(n7318), .ZN(n7344) );
  INV_X1 U8929 ( .A(n7226), .ZN(n7227) );
  NAND2_X1 U8930 ( .A1(n7227), .A2(n7326), .ZN(n7228) );
  AND2_X1 U8931 ( .A1(n7344), .A2(n7228), .ZN(n7233) );
  NOR3_X1 U8932 ( .A1(n7230), .A2(n7229), .A3(n7233), .ZN(n7235) );
  NAND2_X1 U8933 ( .A1(n7232), .A2(n7231), .ZN(n7234) );
  NAND2_X1 U8934 ( .A1(n7234), .A2(n7233), .ZN(n7345) );
  INV_X1 U8935 ( .A(n7345), .ZN(n7343) );
  OAI21_X1 U8936 ( .B1(n7235), .B2(n7343), .A(n7348), .ZN(n7236) );
  OAI211_X1 U8937 ( .C1(n7238), .C2(n9986), .A(n7237), .B(n7236), .ZN(P2_U3191) );
  XOR2_X1 U8938 ( .A(n7240), .B(n7239), .Z(n7245) );
  AOI22_X1 U8939 ( .A1(n8227), .A2(n9996), .B1(n8211), .B2(n8799), .ZN(n7241)
         );
  OAI21_X1 U8940 ( .B1(n6574), .B2(n8223), .A(n7241), .ZN(n7242) );
  AOI21_X1 U8941 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7243), .A(n7242), .ZN(
        n7244) );
  OAI21_X1 U8942 ( .B1(n7245), .B2(n8230), .A(n7244), .ZN(P2_U3177) );
  AOI21_X1 U8943 ( .B1(n7246), .B2(n7247), .A(n8230), .ZN(n7249) );
  NAND2_X1 U8944 ( .A1(n7249), .A2(n7248), .ZN(n7254) );
  OAI21_X1 U8945 ( .B1(n8245), .B2(n10003), .A(n7250), .ZN(n7252) );
  OAI22_X1 U8946 ( .A1(n4878), .A2(n8223), .B1(n8238), .B2(n7605), .ZN(n7251)
         );
  NOR2_X1 U8947 ( .A1(n7252), .A2(n7251), .ZN(n7253) );
  OAI211_X1 U8948 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8165), .A(n7254), .B(
        n7253), .ZN(P2_U3158) );
  OAI21_X1 U8949 ( .B1(n7257), .B2(n7256), .A(n7255), .ZN(n7258) );
  NAND2_X1 U8950 ( .A1(n7258), .A2(n9096), .ZN(n7262) );
  AOI22_X1 U8951 ( .A1(n9131), .A2(n9197), .B1(n9195), .B2(n4509), .ZN(n7642)
         );
  OAI22_X1 U8952 ( .A1(n9153), .A2(n7642), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7259), .ZN(n7260) );
  AOI21_X1 U8953 ( .B1(n7650), .B2(n6200), .A(n7260), .ZN(n7261) );
  OAI211_X1 U8954 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9708), .A(n7262), .B(
        n7261), .ZN(P1_U3218) );
  NAND2_X1 U8955 ( .A1(n8573), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7263) );
  OAI21_X1 U8956 ( .B1(n8625), .B2(n8573), .A(n7263), .ZN(P2_U3520) );
  INV_X1 U8957 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7264) );
  OAI22_X1 U8958 ( .A1(n7265), .A2(n8952), .B1(n10047), .B2(n7264), .ZN(n7266)
         );
  AOI21_X1 U8959 ( .B1(n7267), .B2(n10047), .A(n7266), .ZN(n7268) );
  INV_X1 U8960 ( .A(n7268), .ZN(P2_U3393) );
  XNOR2_X1 U8961 ( .A(n7270), .B(n7269), .ZN(n7281) );
  INV_X1 U8962 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7277) );
  OAI21_X1 U8963 ( .B1(n7271), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7290), .ZN(
        n7272) );
  AND2_X1 U8964 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7412) );
  AOI21_X1 U8965 ( .B1(n8562), .B2(n7272), .A(n7412), .ZN(n7276) );
  XNOR2_X1 U8966 ( .A(n7273), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n7274) );
  NAND2_X1 U8967 ( .A1(n9991), .A2(n7274), .ZN(n7275) );
  OAI211_X1 U8968 ( .C1(n8515), .C2(n7277), .A(n7276), .B(n7275), .ZN(n7278)
         );
  AOI21_X1 U8969 ( .B1(n7279), .B2(n9937), .A(n7278), .ZN(n7280) );
  OAI21_X1 U8970 ( .B1(n9981), .B2(n7281), .A(n7280), .ZN(P2_U3187) );
  AOI21_X1 U8971 ( .B1(n7284), .B2(n7283), .A(n7282), .ZN(n7301) );
  AOI21_X1 U8972 ( .B1(n7287), .B2(n7286), .A(n7285), .ZN(n7298) );
  AND3_X1 U8973 ( .A1(n7290), .A2(n7289), .A3(n7288), .ZN(n7292) );
  OR2_X1 U8974 ( .A1(n7292), .A2(n7291), .ZN(n7294) );
  INV_X1 U8975 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7293) );
  NOR2_X1 U8976 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7293), .ZN(n7507) );
  AOI21_X1 U8977 ( .B1(n8562), .B2(n7294), .A(n7507), .ZN(n7297) );
  INV_X1 U8978 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7295) );
  OR2_X1 U8979 ( .A1(n8515), .A2(n7295), .ZN(n7296) );
  OAI211_X1 U8980 ( .C1(n8582), .C2(n7298), .A(n7297), .B(n7296), .ZN(n7299)
         );
  AOI21_X1 U8981 ( .B1(n4691), .B2(n9937), .A(n7299), .ZN(n7300) );
  OAI21_X1 U8982 ( .B1(n7301), .B2(n9981), .A(n7300), .ZN(P2_U3188) );
  NOR2_X1 U8983 ( .A1(n7423), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7302) );
  AOI21_X1 U8984 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7423), .A(n7302), .ZN(
        n7305) );
  NAND2_X1 U8985 ( .A1(n7305), .A2(n7304), .ZN(n7418) );
  OAI21_X1 U8986 ( .B1(n7305), .B2(n7304), .A(n7418), .ZN(n7306) );
  NAND2_X1 U8987 ( .A1(n7306), .A2(n9720), .ZN(n7316) );
  AOI22_X1 U8988 ( .A1(n7423), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n5534), .B2(
        n7312), .ZN(n7309) );
  OAI21_X1 U8989 ( .B1(n7310), .B2(n7309), .A(n7422), .ZN(n7314) );
  INV_X1 U8990 ( .A(n9724), .ZN(n9311) );
  NAND2_X1 U8991 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U8992 ( .A1(n9715), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n7311) );
  OAI211_X1 U8993 ( .C1(n9311), .C2(n7312), .A(n9047), .B(n7311), .ZN(n7313)
         );
  AOI21_X1 U8994 ( .B1(n7314), .B2(n9338), .A(n7313), .ZN(n7315) );
  NAND2_X1 U8995 ( .A1(n7316), .A2(n7315), .ZN(P1_U3255) );
  NOR2_X1 U8996 ( .A1(n7318), .A2(n7317), .ZN(n7319) );
  NAND2_X1 U8997 ( .A1(n7435), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7432) );
  INV_X1 U8998 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7337) );
  NAND2_X1 U8999 ( .A1(n7338), .A2(n7337), .ZN(n7321) );
  NAND2_X1 U9000 ( .A1(n7432), .A2(n7321), .ZN(n7323) );
  INV_X1 U9001 ( .A(n7433), .ZN(n7322) );
  AOI21_X1 U9002 ( .B1(n7324), .B2(n7323), .A(n7322), .ZN(n7353) );
  NAND2_X1 U9003 ( .A1(n7326), .A2(n7325), .ZN(n7328) );
  INV_X1 U9004 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7336) );
  MUX2_X1 U9005 ( .A(n7336), .B(P2_REG1_REG_10__SCAN_IN), .S(n7338), .Z(n7329)
         );
  NAND2_X1 U9006 ( .A1(n7329), .A2(n7330), .ZN(n7436) );
  OAI21_X1 U9007 ( .B1(n7330), .B2(n7329), .A(n7436), .ZN(n7335) );
  INV_X1 U9008 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7333) );
  NAND2_X1 U9009 ( .A1(n9937), .A2(n7338), .ZN(n7332) );
  INV_X1 U9010 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10296) );
  NOR2_X1 U9011 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10296), .ZN(n7931) );
  INV_X1 U9012 ( .A(n7931), .ZN(n7331) );
  OAI211_X1 U9013 ( .C1(n7333), .C2(n8515), .A(n7332), .B(n7331), .ZN(n7334)
         );
  AOI21_X1 U9014 ( .B1(n7335), .B2(n9991), .A(n7334), .ZN(n7352) );
  INV_X1 U9015 ( .A(n7344), .ZN(n7342) );
  MUX2_X1 U9016 ( .A(n7337), .B(n7336), .S(n8540), .Z(n7339) );
  NAND2_X1 U9017 ( .A1(n7339), .A2(n7338), .ZN(n7445) );
  INV_X1 U9018 ( .A(n7339), .ZN(n7340) );
  NAND2_X1 U9019 ( .A1(n7340), .A2(n7435), .ZN(n7341) );
  AND2_X1 U9020 ( .A1(n7445), .A2(n7341), .ZN(n7346) );
  NOR3_X1 U9021 ( .A1(n7343), .A2(n7342), .A3(n7346), .ZN(n7350) );
  NAND2_X1 U9022 ( .A1(n7345), .A2(n7344), .ZN(n7347) );
  NAND2_X1 U9023 ( .A1(n7347), .A2(n7346), .ZN(n7446) );
  INV_X1 U9024 ( .A(n7446), .ZN(n7349) );
  OAI21_X1 U9025 ( .B1(n7350), .B2(n7349), .A(n7348), .ZN(n7351) );
  OAI211_X1 U9026 ( .C1(n7353), .C2(n9986), .A(n7352), .B(n7351), .ZN(P2_U3192) );
  AND2_X1 U9027 ( .A1(n7255), .A2(n7354), .ZN(n7357) );
  OAI211_X1 U9028 ( .C1(n7357), .C2(n7356), .A(n9096), .B(n7355), .ZN(n7360)
         );
  AOI22_X1 U9029 ( .A1(n9131), .A2(n9196), .B1(n9695), .B2(n4509), .ZN(n9780)
         );
  OAI22_X1 U9030 ( .A1(n9153), .A2(n9780), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9233), .ZN(n7358) );
  AOI21_X1 U9031 ( .B1(n9789), .B2(n6200), .A(n7358), .ZN(n7359) );
  OAI211_X1 U9032 ( .C1(n9708), .C2(n9784), .A(n7360), .B(n7359), .ZN(P1_U3230) );
  INV_X1 U9033 ( .A(n7361), .ZN(n7363) );
  NAND2_X1 U9034 ( .A1(n7363), .A2(n7362), .ZN(n7364) );
  NAND2_X1 U9035 ( .A1(n7365), .A2(n7364), .ZN(n7367) );
  AOI22_X1 U9036 ( .A1(n4507), .A2(n7369), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8808), .ZN(n7374) );
  NOR3_X1 U9037 ( .A1(n8265), .A2(n7370), .A3(n10046), .ZN(n7371) );
  OAI21_X1 U9038 ( .B1(n7372), .B2(n7371), .A(n8812), .ZN(n7373) );
  OAI211_X1 U9039 ( .C1(n6950), .C2(n8812), .A(n7374), .B(n7373), .ZN(P2_U3233) );
  INV_X1 U9040 ( .A(n7375), .ZN(n7376) );
  INV_X1 U9041 ( .A(n8566), .ZN(n8554) );
  OAI222_X1 U9042 ( .A1(n8102), .A2(n10284), .B1(n8965), .B2(n7376), .C1(
        P2_U3151), .C2(n8554), .ZN(P2_U3278) );
  INV_X1 U9043 ( .A(n9318), .ZN(n9310) );
  OAI222_X1 U9044 ( .A1(n9633), .A2(n10364), .B1(n9629), .B2(n7376), .C1(
        P1_U3086), .C2(n9310), .ZN(P1_U3338) );
  INV_X1 U9045 ( .A(n7377), .ZN(n7378) );
  AOI21_X1 U9046 ( .B1(n7380), .B2(n7379), .A(n7378), .ZN(n7387) );
  INV_X1 U9047 ( .A(n7381), .ZN(n7595) );
  OAI22_X1 U9048 ( .A1(n7505), .A2(n8238), .B1(n8223), .B2(n6293), .ZN(n7384)
         );
  NOR2_X1 U9049 ( .A1(n8245), .A2(n10008), .ZN(n7383) );
  OR3_X1 U9050 ( .A1(n7384), .A2(n7383), .A3(n7382), .ZN(n7385) );
  AOI21_X1 U9051 ( .B1(n7595), .B2(n8241), .A(n7385), .ZN(n7386) );
  OAI21_X1 U9052 ( .B1(n7387), .B2(n8230), .A(n7386), .ZN(P2_U3170) );
  INV_X1 U9053 ( .A(n7388), .ZN(n7409) );
  AOI22_X1 U9054 ( .A1(n9325), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n7389), .ZN(n7390) );
  OAI21_X1 U9055 ( .B1(n7409), .B2(n9629), .A(n7390), .ZN(P1_U3337) );
  INV_X1 U9056 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10067) );
  INV_X1 U9057 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10356) );
  INV_X1 U9058 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10277) );
  AOI22_X1 U9059 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n10356), .B2(n10277), .ZN(n10072) );
  NOR2_X1 U9060 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7391) );
  AOI21_X1 U9061 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7391), .ZN(n10075) );
  NOR2_X1 U9062 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7392) );
  AOI21_X1 U9063 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7392), .ZN(n10078) );
  INV_X1 U9064 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10312) );
  INV_X1 U9065 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10267) );
  AOI22_X1 U9066 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .B1(n10312), .B2(n10267), .ZN(n10081) );
  NOR2_X1 U9067 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7393) );
  AOI21_X1 U9068 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7393), .ZN(n10084) );
  NOR2_X1 U9069 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7394) );
  AOI21_X1 U9070 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7394), .ZN(n10087) );
  INV_X1 U9071 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7449) );
  AOI22_X1 U9072 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .B1(n10350), .B2(n7449), .ZN(n10090) );
  NOR2_X1 U9073 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7395) );
  AOI21_X1 U9074 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7395), .ZN(n10093) );
  NOR2_X1 U9075 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7396) );
  AOI21_X1 U9076 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7396), .ZN(n10477) );
  NOR2_X1 U9077 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7397) );
  AOI21_X1 U9078 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7397), .ZN(n10483) );
  INV_X1 U9079 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7398) );
  AOI22_X1 U9080 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(P2_ADDR_REG_7__SCAN_IN), 
        .B1(n7398), .B2(n10305), .ZN(n10480) );
  NOR2_X1 U9081 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7399) );
  AOI21_X1 U9082 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7399), .ZN(n10471) );
  NOR2_X1 U9083 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7400) );
  AOI21_X1 U9084 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7400), .ZN(n10474) );
  AND2_X1 U9085 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7401) );
  NOR2_X1 U9086 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7401), .ZN(n10062) );
  INV_X1 U9087 ( .A(n10062), .ZN(n10063) );
  NAND3_X1 U9088 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10064) );
  NAND2_X1 U9089 ( .A1(n10065), .A2(n10064), .ZN(n10061) );
  NAND2_X1 U9090 ( .A1(n10063), .A2(n10061), .ZN(n10486) );
  NAND2_X1 U9091 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7402) );
  OAI21_X1 U9092 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n7402), .ZN(n10485) );
  NOR2_X1 U9093 ( .A1(n10486), .A2(n10485), .ZN(n10484) );
  AOI21_X1 U9094 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10484), .ZN(n10489) );
  NAND2_X1 U9095 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7403) );
  OAI21_X1 U9096 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7403), .ZN(n10488) );
  NOR2_X1 U9097 ( .A1(n10489), .A2(n10488), .ZN(n10487) );
  AOI21_X1 U9098 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10487), .ZN(n10492) );
  NOR2_X1 U9099 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7404) );
  AOI21_X1 U9100 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7404), .ZN(n10491) );
  NAND2_X1 U9101 ( .A1(n10492), .A2(n10491), .ZN(n10490) );
  OAI21_X1 U9102 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10490), .ZN(n10473) );
  NAND2_X1 U9103 ( .A1(n10474), .A2(n10473), .ZN(n10472) );
  OAI21_X1 U9104 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10472), .ZN(n10470) );
  NAND2_X1 U9105 ( .A1(n10471), .A2(n10470), .ZN(n10469) );
  OAI21_X1 U9106 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10469), .ZN(n10479) );
  NAND2_X1 U9107 ( .A1(n10480), .A2(n10479), .ZN(n10478) );
  OAI21_X1 U9108 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n10478), .ZN(n10482) );
  NAND2_X1 U9109 ( .A1(n10483), .A2(n10482), .ZN(n10481) );
  OAI21_X1 U9110 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10481), .ZN(n10476) );
  NAND2_X1 U9111 ( .A1(n10477), .A2(n10476), .ZN(n10475) );
  OAI21_X1 U9112 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10475), .ZN(n10092) );
  NAND2_X1 U9113 ( .A1(n10093), .A2(n10092), .ZN(n10091) );
  OAI21_X1 U9114 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10091), .ZN(n10089) );
  NAND2_X1 U9115 ( .A1(n10090), .A2(n10089), .ZN(n10088) );
  OAI21_X1 U9116 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10088), .ZN(n10086) );
  NAND2_X1 U9117 ( .A1(n10087), .A2(n10086), .ZN(n10085) );
  OAI21_X1 U9118 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10085), .ZN(n10083) );
  NAND2_X1 U9119 ( .A1(n10084), .A2(n10083), .ZN(n10082) );
  OAI21_X1 U9120 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10082), .ZN(n10080) );
  NAND2_X1 U9121 ( .A1(n10081), .A2(n10080), .ZN(n10079) );
  OAI21_X1 U9122 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10079), .ZN(n10077) );
  NAND2_X1 U9123 ( .A1(n10078), .A2(n10077), .ZN(n10076) );
  OAI21_X1 U9124 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10076), .ZN(n10074) );
  NAND2_X1 U9125 ( .A1(n10075), .A2(n10074), .ZN(n10073) );
  OAI21_X1 U9126 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10073), .ZN(n10071) );
  NAND2_X1 U9127 ( .A1(n10072), .A2(n10071), .ZN(n10070) );
  OAI21_X1 U9128 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10070), .ZN(n10068) );
  NAND2_X1 U9129 ( .A1(n10067), .A2(n10068), .ZN(n7405) );
  NOR2_X1 U9130 ( .A1(n10067), .A2(n10068), .ZN(n10066) );
  AOI21_X1 U9131 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7405), .A(n10066), .ZN(
        n7408) );
  XNOR2_X1 U9132 ( .A(n7406), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7407) );
  XNOR2_X1 U9133 ( .A(n7408), .B(n7407), .ZN(ADD_1068_U4) );
  INV_X1 U9134 ( .A(n8557), .ZN(n8590) );
  OAI222_X1 U9135 ( .A1(n8102), .A2(n10233), .B1(n8590), .B2(P2_U3151), .C1(
        n8965), .C2(n7409), .ZN(P2_U3277) );
  XOR2_X1 U9136 ( .A(n7411), .B(n7410), .Z(n7417) );
  INV_X1 U9137 ( .A(n8478), .ZN(n7701) );
  OAI22_X1 U9138 ( .A1(n7605), .A2(n8223), .B1(n8238), .B2(n7701), .ZN(n7414)
         );
  NOR2_X1 U9139 ( .A1(n8245), .A2(n10012), .ZN(n7413) );
  OR3_X1 U9140 ( .A1(n7414), .A2(n7413), .A3(n7412), .ZN(n7415) );
  AOI21_X1 U9141 ( .B1(n7609), .B2(n8241), .A(n7415), .ZN(n7416) );
  OAI21_X1 U9142 ( .B1(n7417), .B2(n8230), .A(n7416), .ZN(P2_U3167) );
  OAI21_X1 U9143 ( .B1(n7423), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7418), .ZN(
        n7420) );
  XNOR2_X1 U9144 ( .A(n7623), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n7419) );
  NOR2_X1 U9145 ( .A1(n7420), .A2(n7419), .ZN(n7622) );
  AOI211_X1 U9146 ( .C1(n7420), .C2(n7419), .A(n9289), .B(n7622), .ZN(n7431)
         );
  MUX2_X1 U9147 ( .A(n7421), .B(P1_REG1_REG_13__SCAN_IN), .S(n7623), .Z(n7425)
         );
  OAI21_X1 U9148 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n7423), .A(n7422), .ZN(
        n7424) );
  NOR2_X1 U9149 ( .A1(n7424), .A2(n7425), .ZN(n7618) );
  AOI211_X1 U9150 ( .C1(n7425), .C2(n7424), .A(n9727), .B(n7618), .ZN(n7430)
         );
  INV_X1 U9151 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7428) );
  NAND2_X1 U9152 ( .A1(n9724), .A2(n7623), .ZN(n7427) );
  NAND2_X1 U9153 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n7426) );
  OAI211_X1 U9154 ( .C1(n7428), .C2(n9344), .A(n7427), .B(n7426), .ZN(n7429)
         );
  OR3_X1 U9155 ( .A1(n7431), .A2(n7430), .A3(n7429), .ZN(P1_U3256) );
  INV_X1 U9156 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7893) );
  NOR2_X1 U9157 ( .A1(n7893), .A2(n7434), .ZN(n7559) );
  AOI21_X1 U9158 ( .B1(n7893), .B2(n7434), .A(n7559), .ZN(n7454) );
  NAND2_X1 U9159 ( .A1(n7435), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7437) );
  NAND2_X1 U9160 ( .A1(n7437), .A2(n7436), .ZN(n7563) );
  XNOR2_X1 U9161 ( .A(n7563), .B(n7558), .ZN(n7438) );
  NAND2_X1 U9162 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n7438), .ZN(n7565) );
  OAI21_X1 U9163 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7438), .A(n7565), .ZN(
        n7452) );
  NAND2_X1 U9164 ( .A1(n7446), .A2(n7445), .ZN(n7442) );
  INV_X1 U9165 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7889) );
  MUX2_X1 U9166 ( .A(n7893), .B(n7889), .S(n8540), .Z(n7439) );
  NAND2_X1 U9167 ( .A1(n7439), .A2(n7558), .ZN(n7574) );
  INV_X1 U9168 ( .A(n7439), .ZN(n7440) );
  NAND2_X1 U9169 ( .A1(n7440), .A2(n7564), .ZN(n7441) );
  AND2_X1 U9170 ( .A1(n7574), .A2(n7441), .ZN(n7443) );
  NAND2_X1 U9171 ( .A1(n7442), .A2(n7443), .ZN(n7575) );
  INV_X1 U9172 ( .A(n7443), .ZN(n7444) );
  NAND3_X1 U9173 ( .A1(n7446), .A2(n7445), .A3(n7444), .ZN(n7447) );
  AOI21_X1 U9174 ( .B1(n7575), .B2(n7447), .A(n9981), .ZN(n7451) );
  NAND2_X1 U9175 ( .A1(n9937), .A2(n7558), .ZN(n7448) );
  NAND2_X1 U9176 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7977) );
  OAI211_X1 U9177 ( .C1(n7449), .C2(n8515), .A(n7448), .B(n7977), .ZN(n7450)
         );
  AOI211_X1 U9178 ( .C1(n7452), .C2(n9991), .A(n7451), .B(n7450), .ZN(n7453)
         );
  OAI21_X1 U9179 ( .B1(n7454), .B2(n9986), .A(n7453), .ZN(P2_U3193) );
  AND2_X1 U9180 ( .A1(n7455), .A2(n6679), .ZN(n8796) );
  MUX2_X1 U9181 ( .A(n7458), .B(n7457), .S(n8771), .Z(n7460) );
  AOI22_X1 U9182 ( .A1(n4507), .A2(n6573), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8808), .ZN(n7459) );
  OAI211_X1 U9183 ( .C1(n7461), .C2(n8793), .A(n7460), .B(n7459), .ZN(P2_U3232) );
  INV_X1 U9184 ( .A(n9833), .ZN(n7464) );
  NAND4_X1 U9185 ( .A1(n7465), .A2(n7464), .A3(n7463), .A4(n7462), .ZN(n7466)
         );
  INV_X1 U9186 ( .A(n7467), .ZN(n7468) );
  NOR2_X1 U9187 ( .A1(n8097), .A2(n7468), .ZN(n7469) );
  NAND2_X1 U9188 ( .A1(n9516), .A2(n7469), .ZN(n9736) );
  INV_X1 U9189 ( .A(n9872), .ZN(n9905) );
  NAND2_X1 U9190 ( .A1(n9516), .A2(n9905), .ZN(n7470) );
  AND2_X1 U9191 ( .A1(n5974), .A2(n7673), .ZN(n7549) );
  XNOR2_X1 U9192 ( .A(n7519), .B(n7518), .ZN(n9846) );
  INV_X1 U9193 ( .A(n9846), .ZN(n7489) );
  NOR2_X1 U9194 ( .A1(n9835), .A2(n7673), .ZN(n7473) );
  NAND2_X1 U9195 ( .A1(n7473), .A2(n9844), .ZN(n7646) );
  OAI211_X1 U9196 ( .C1(n7473), .C2(n9844), .A(n9793), .B(n7646), .ZN(n9842)
         );
  INV_X1 U9197 ( .A(n9842), .ZN(n7487) );
  NOR2_X2 U9198 ( .A1(n9785), .A2(n5883), .ZN(n9757) );
  INV_X1 U9199 ( .A(n7474), .ZN(n7475) );
  NOR2_X1 U9200 ( .A1(n9513), .A2(n7476), .ZN(n7477) );
  AOI21_X1 U9201 ( .B1(n9785), .B2(P1_REG2_REG_2__SCAN_IN), .A(n7477), .ZN(
        n7478) );
  OAI21_X1 U9202 ( .B1(n9500), .B2(n9844), .A(n7478), .ZN(n7486) );
  OAI21_X1 U9203 ( .B1(n7479), .B2(n7481), .A(n7480), .ZN(n7484) );
  INV_X1 U9204 ( .A(n7482), .ZN(n7483) );
  AOI21_X1 U9205 ( .B1(n7484), .B2(n9782), .A(n7483), .ZN(n9843) );
  NOR2_X1 U9206 ( .A1(n9843), .A2(n9785), .ZN(n7485) );
  AOI211_X1 U9207 ( .C1(n7487), .C2(n9757), .A(n7486), .B(n7485), .ZN(n7488)
         );
  OAI21_X1 U9208 ( .B1(n9662), .B2(n7489), .A(n7488), .ZN(P1_U3291) );
  NAND2_X1 U9209 ( .A1(n7606), .A2(n8310), .ZN(n7490) );
  XNOR2_X1 U9210 ( .A(n7490), .B(n8266), .ZN(n10017) );
  INV_X1 U9211 ( .A(n8266), .ZN(n7493) );
  NAND3_X1 U9212 ( .A1(n7491), .A2(n7493), .A3(n7492), .ZN(n7494) );
  NAND2_X1 U9213 ( .A1(n7495), .A2(n7494), .ZN(n7496) );
  AOI222_X1 U9214 ( .A1(n8805), .A2(n7496), .B1(n8477), .B2(n8800), .C1(n8479), 
        .C2(n8801), .ZN(n10018) );
  MUX2_X1 U9215 ( .A(n4690), .B(n10018), .S(n8812), .Z(n7499) );
  AOI22_X1 U9216 ( .A1(n4507), .A2(n7497), .B1(n8808), .B2(n7500), .ZN(n7498)
         );
  OAI211_X1 U9217 ( .C1(n8793), .C2(n10017), .A(n7499), .B(n7498), .ZN(
        P2_U3227) );
  INV_X1 U9218 ( .A(n7500), .ZN(n7510) );
  AOI21_X1 U9219 ( .B1(n7501), .B2(n7502), .A(n8230), .ZN(n7504) );
  NAND2_X1 U9220 ( .A1(n7504), .A2(n7503), .ZN(n7509) );
  OAI22_X1 U9221 ( .A1(n8245), .A2(n10019), .B1(n8223), .B2(n7505), .ZN(n7506)
         );
  AOI211_X1 U9222 ( .C1(n8211), .C2(n8477), .A(n7507), .B(n7506), .ZN(n7508)
         );
  OAI211_X1 U9223 ( .C1(n7510), .C2(n8165), .A(n7509), .B(n7508), .ZN(P2_U3179) );
  OAI21_X1 U9224 ( .B1(n7513), .B2(n7511), .A(n7512), .ZN(n7514) );
  NAND2_X1 U9225 ( .A1(n7514), .A2(n9096), .ZN(n7517) );
  AOI22_X1 U9226 ( .A1(n9131), .A2(n9195), .B1(n9194), .B2(n4509), .ZN(n7686)
         );
  NAND2_X1 U9227 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9249) );
  OAI21_X1 U9228 ( .B1(n9153), .B2(n7686), .A(n9249), .ZN(n7515) );
  AOI21_X1 U9229 ( .B1(n9859), .B2(n6200), .A(n7515), .ZN(n7516) );
  OAI211_X1 U9230 ( .C1(n9708), .C2(n7691), .A(n7517), .B(n7516), .ZN(P1_U3227) );
  NAND2_X1 U9231 ( .A1(n7519), .A2(n7518), .ZN(n7522) );
  NAND2_X1 U9232 ( .A1(n7520), .A2(n9844), .ZN(n7521) );
  NAND2_X1 U9233 ( .A1(n7522), .A2(n7521), .ZN(n7644) );
  NAND2_X1 U9234 ( .A1(n7644), .A2(n7645), .ZN(n7525) );
  INV_X1 U9235 ( .A(n9196), .ZN(n7523) );
  NAND2_X1 U9236 ( .A1(n7523), .A2(n5754), .ZN(n7524) );
  NAND2_X1 U9237 ( .A1(n7525), .A2(n7524), .ZN(n9790) );
  NAND2_X1 U9238 ( .A1(n9790), .A2(n9791), .ZN(n7528) );
  NAND2_X1 U9239 ( .A1(n7526), .A2(n4839), .ZN(n7527) );
  NAND2_X1 U9240 ( .A1(n7528), .A2(n7527), .ZN(n7683) );
  NAND2_X1 U9241 ( .A1(n7683), .A2(n7684), .ZN(n7531) );
  NAND2_X1 U9242 ( .A1(n7529), .A2(n7692), .ZN(n7530) );
  NAND2_X1 U9243 ( .A1(n7531), .A2(n7530), .ZN(n9773) );
  NAND2_X1 U9244 ( .A1(n7532), .A2(n9867), .ZN(n7533) );
  XOR2_X1 U9245 ( .A(n7714), .B(n7713), .Z(n9871) );
  AOI21_X1 U9246 ( .B1(n7713), .B2(n7534), .A(n7708), .ZN(n7538) );
  NAND2_X1 U9247 ( .A1(n9193), .A2(n4509), .ZN(n7536) );
  NAND2_X1 U9248 ( .A1(n9194), .A2(n9131), .ZN(n7535) );
  NAND2_X1 U9249 ( .A1(n7536), .A2(n7535), .ZN(n7730) );
  INV_X1 U9250 ( .A(n7730), .ZN(n7537) );
  OAI21_X1 U9251 ( .B1(n7538), .B2(n9765), .A(n7537), .ZN(n9877) );
  NAND2_X1 U9252 ( .A1(n9877), .A2(n9516), .ZN(n7544) );
  NOR2_X1 U9253 ( .A1(n9792), .A2(n9789), .ZN(n7690) );
  AND2_X1 U9254 ( .A1(n7690), .A2(n7692), .ZN(n9775) );
  NAND2_X1 U9255 ( .A1(n9775), .A2(n9867), .ZN(n9774) );
  AOI211_X1 U9256 ( .C1(n7539), .C2(n9774), .A(n9600), .B(n4760), .ZN(n9875)
         );
  NOR2_X1 U9257 ( .A1(n9500), .A2(n9873), .ZN(n7542) );
  OAI22_X1 U9258 ( .A1(n9516), .A2(n7540), .B1(n7733), .B2(n9513), .ZN(n7541)
         );
  AOI211_X1 U9259 ( .C1(n9875), .C2(n9757), .A(n7542), .B(n7541), .ZN(n7543)
         );
  OAI211_X1 U9260 ( .C1(n9662), .C2(n9871), .A(n7544), .B(n7543), .ZN(P1_U3286) );
  INV_X1 U9261 ( .A(n7546), .ZN(n7547) );
  AOI21_X1 U9262 ( .B1(n7548), .B2(n9782), .A(n7547), .ZN(n9840) );
  INV_X1 U9263 ( .A(n9835), .ZN(n7554) );
  NAND2_X1 U9264 ( .A1(n9835), .A2(n7673), .ZN(n7550) );
  NAND2_X1 U9265 ( .A1(n7550), .A2(n9793), .ZN(n7551) );
  NOR2_X1 U9266 ( .A1(n7473), .A2(n7551), .ZN(n9834) );
  NAND2_X1 U9267 ( .A1(n9757), .A2(n9834), .ZN(n7553) );
  INV_X1 U9268 ( .A(n9513), .ZN(n9786) );
  AOI22_X1 U9269 ( .A1(n9785), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9786), .ZN(n7552) );
  OAI211_X1 U9270 ( .C1(n9500), .C2(n7554), .A(n7553), .B(n7552), .ZN(n7555)
         );
  AOI21_X1 U9271 ( .B1(n9836), .B2(n9797), .A(n7555), .ZN(n7556) );
  OAI21_X1 U9272 ( .B1(n9785), .B2(n9840), .A(n7556), .ZN(P1_U3292) );
  NOR2_X1 U9273 ( .A1(n7558), .A2(n7557), .ZN(n7560) );
  INV_X1 U9274 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7906) );
  AOI22_X1 U9275 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8490), .B1(n8484), .B2(
        n7906), .ZN(n7561) );
  NOR2_X1 U9276 ( .A1(n7562), .A2(n7561), .ZN(n8483) );
  AOI21_X1 U9277 ( .B1(n7562), .B2(n7561), .A(n8483), .ZN(n7584) );
  INV_X1 U9278 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8489) );
  AOI22_X1 U9279 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8484), .B1(n8490), .B2(
        n8489), .ZN(n7568) );
  NAND2_X1 U9280 ( .A1(n7564), .A2(n7563), .ZN(n7566) );
  NAND2_X1 U9281 ( .A1(n7566), .A2(n7565), .ZN(n7567) );
  NAND2_X1 U9282 ( .A1(n7568), .A2(n7567), .ZN(n8488) );
  OAI21_X1 U9283 ( .B1(n7568), .B2(n7567), .A(n8488), .ZN(n7582) );
  NAND2_X1 U9284 ( .A1(n7575), .A2(n7574), .ZN(n7571) );
  MUX2_X1 U9285 ( .A(n7906), .B(n8489), .S(n8540), .Z(n7569) );
  OR2_X1 U9286 ( .A1(n8490), .A2(n7569), .ZN(n7570) );
  NAND2_X1 U9287 ( .A1(n7569), .A2(n8490), .ZN(n9943) );
  AND2_X1 U9288 ( .A1(n7570), .A2(n9943), .ZN(n7572) );
  NAND2_X1 U9289 ( .A1(n7571), .A2(n7572), .ZN(n9944) );
  INV_X1 U9290 ( .A(n7572), .ZN(n7573) );
  NAND3_X1 U9291 ( .A1(n7575), .A2(n7574), .A3(n7573), .ZN(n7576) );
  AOI21_X1 U9292 ( .B1(n9944), .B2(n7576), .A(n9981), .ZN(n7581) );
  INV_X1 U9293 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7579) );
  NAND2_X1 U9294 ( .A1(n9937), .A2(n8490), .ZN(n7578) );
  INV_X1 U9295 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7577) );
  OR2_X1 U9296 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7577), .ZN(n8016) );
  OAI211_X1 U9297 ( .C1(n7579), .C2(n8515), .A(n7578), .B(n8016), .ZN(n7580)
         );
  AOI211_X1 U9298 ( .C1(n7582), .C2(n9991), .A(n7581), .B(n7580), .ZN(n7583)
         );
  OAI21_X1 U9299 ( .B1(n7584), .B2(n9986), .A(n7583), .ZN(P2_U3194) );
  XNOR2_X1 U9300 ( .A(n7585), .B(n7586), .ZN(n7587) );
  AOI222_X1 U9301 ( .A1(n8805), .A2(n7587), .B1(n8480), .B2(n8800), .C1(n8481), 
        .C2(n8801), .ZN(n10002) );
  XNOR2_X1 U9302 ( .A(n8294), .B(n8264), .ZN(n10005) );
  NAND2_X1 U9303 ( .A1(n4507), .A2(n6292), .ZN(n7589) );
  NAND2_X1 U9304 ( .A1(n8771), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7588) );
  OAI211_X1 U9305 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8674), .A(n7589), .B(
        n7588), .ZN(n7590) );
  AOI21_X1 U9306 ( .B1(n8727), .B2(n10005), .A(n7590), .ZN(n7591) );
  OAI21_X1 U9307 ( .B1(n10002), .B2(n8771), .A(n7591), .ZN(P2_U3230) );
  AND2_X1 U9308 ( .A1(n8311), .A2(n8304), .ZN(n8302) );
  INV_X1 U9309 ( .A(n8302), .ZN(n8267) );
  XNOR2_X1 U9310 ( .A(n7592), .B(n8267), .ZN(n7593) );
  AOI222_X1 U9311 ( .A1(n8805), .A2(n7593), .B1(n8799), .B2(n8801), .C1(n8479), 
        .C2(n8800), .ZN(n10007) );
  XNOR2_X1 U9312 ( .A(n7594), .B(n8302), .ZN(n10010) );
  AOI22_X1 U9313 ( .A1(n4507), .A2(n7596), .B1(n8808), .B2(n7595), .ZN(n7597)
         );
  OAI21_X1 U9314 ( .B1(n7598), .B2(n8812), .A(n7597), .ZN(n7599) );
  AOI21_X1 U9315 ( .B1(n8727), .B2(n10010), .A(n7599), .ZN(n7600) );
  OAI21_X1 U9316 ( .B1(n10007), .B2(n8771), .A(n7600), .ZN(P2_U3229) );
  INV_X1 U9317 ( .A(n7601), .ZN(n7603) );
  INV_X1 U9318 ( .A(n7491), .ZN(n7602) );
  AOI21_X1 U9319 ( .B1(n7607), .B2(n7603), .A(n7602), .ZN(n7604) );
  OAI222_X1 U9320 ( .A1(n8748), .A2(n7701), .B1(n8779), .B2(n7605), .C1(n8782), 
        .C2(n7604), .ZN(n10013) );
  INV_X1 U9321 ( .A(n10013), .ZN(n7615) );
  OAI21_X1 U9322 ( .B1(n7608), .B2(n7607), .A(n7606), .ZN(n10015) );
  INV_X1 U9323 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7612) );
  AOI22_X1 U9324 ( .A1(n4507), .A2(n7610), .B1(n8808), .B2(n7609), .ZN(n7611)
         );
  OAI21_X1 U9325 ( .B1(n7612), .B2(n8812), .A(n7611), .ZN(n7613) );
  AOI21_X1 U9326 ( .B1(n8727), .B2(n10015), .A(n7613), .ZN(n7614) );
  OAI21_X1 U9327 ( .B1(n7615), .B2(n8771), .A(n7614), .ZN(P2_U3228) );
  INV_X1 U9328 ( .A(n7616), .ZN(n8099) );
  OAI222_X1 U9329 ( .A1(n8102), .A2(n7617), .B1(n8965), .B2(n8099), .C1(n8599), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  MUX2_X1 U9330 ( .A(n7619), .B(P1_REG1_REG_14__SCAN_IN), .S(n7855), .Z(n7620)
         );
  AOI211_X1 U9331 ( .C1(n7621), .C2(n7620), .A(n9727), .B(n7854), .ZN(n7631)
         );
  NAND2_X1 U9332 ( .A1(n7855), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7624) );
  OAI21_X1 U9333 ( .B1(n7855), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7624), .ZN(
        n7625) );
  NOR2_X1 U9334 ( .A1(n7626), .A2(n7625), .ZN(n7850) );
  AOI211_X1 U9335 ( .C1(n7626), .C2(n7625), .A(n7850), .B(n9289), .ZN(n7630)
         );
  NAND2_X1 U9336 ( .A1(n9724), .A2(n7855), .ZN(n7628) );
  NAND2_X1 U9337 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n7627) );
  OAI211_X1 U9338 ( .C1(n10312), .C2(n9344), .A(n7628), .B(n7627), .ZN(n7629)
         );
  OR3_X1 U9339 ( .A1(n7631), .A2(n7630), .A3(n7629), .ZN(P1_U3257) );
  INV_X1 U9340 ( .A(n8327), .ZN(n7632) );
  NOR2_X1 U9341 ( .A1(n8335), .A2(n7632), .ZN(n8270) );
  XNOR2_X1 U9342 ( .A(n7633), .B(n8270), .ZN(n10032) );
  XNOR2_X1 U9343 ( .A(n7634), .B(n8270), .ZN(n7635) );
  OAI222_X1 U9344 ( .A1(n8748), .A2(n7934), .B1(n8779), .B2(n8325), .C1(n8782), 
        .C2(n7635), .ZN(n10034) );
  NAND2_X1 U9345 ( .A1(n10034), .A2(n8812), .ZN(n7640) );
  INV_X1 U9346 ( .A(n7765), .ZN(n7636) );
  OAI22_X1 U9347 ( .A1(n8812), .A2(n7637), .B1(n7636), .B2(n8674), .ZN(n7638)
         );
  AOI21_X1 U9348 ( .B1(n4507), .B2(n7770), .A(n7638), .ZN(n7639) );
  OAI211_X1 U9349 ( .C1(n10032), .C2(n8793), .A(n7640), .B(n7639), .ZN(
        P2_U3225) );
  XNOR2_X1 U9350 ( .A(n7641), .B(n7645), .ZN(n7643) );
  OAI21_X1 U9351 ( .B1(n7643), .B2(n9765), .A(n7642), .ZN(n9848) );
  INV_X1 U9352 ( .A(n9848), .ZN(n7654) );
  XNOR2_X1 U9353 ( .A(n7644), .B(n7645), .ZN(n9850) );
  INV_X1 U9354 ( .A(n7646), .ZN(n7647) );
  OAI211_X1 U9355 ( .C1(n7647), .C2(n5754), .A(n9793), .B(n9792), .ZN(n9847)
         );
  OAI22_X1 U9356 ( .A1(n9516), .A2(n7648), .B1(n9513), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n7649) );
  AOI21_X1 U9357 ( .B1(n9788), .B2(n7650), .A(n7649), .ZN(n7651) );
  OAI21_X1 U9358 ( .B1(n9661), .B2(n9847), .A(n7651), .ZN(n7652) );
  AOI21_X1 U9359 ( .B1(n9850), .B2(n9797), .A(n7652), .ZN(n7653) );
  OAI21_X1 U9360 ( .B1(n7654), .B2(n9785), .A(n7653), .ZN(P1_U3290) );
  NAND2_X1 U9361 ( .A1(n7658), .A2(n9625), .ZN(n7656) );
  OAI211_X1 U9362 ( .C1(n7657), .C2(n9633), .A(n7656), .B(n7655), .ZN(P1_U3335) );
  INV_X1 U9363 ( .A(n7658), .ZN(n7660) );
  OAI222_X1 U9364 ( .A1(n8965), .A2(n7660), .B1(P2_U3151), .B2(n8437), .C1(
        n7659), .C2(n8102), .ZN(P2_U3275) );
  INV_X1 U9365 ( .A(n4507), .ZN(n8725) );
  OR2_X1 U9366 ( .A1(n7661), .A2(n8323), .ZN(n7662) );
  NAND2_X1 U9367 ( .A1(n7663), .A2(n7662), .ZN(n10025) );
  INV_X1 U9368 ( .A(n10025), .ZN(n7670) );
  INV_X1 U9369 ( .A(n7664), .ZN(n7705) );
  NOR2_X1 U9370 ( .A1(n8674), .A2(n7705), .ZN(n7669) );
  INV_X1 U9371 ( .A(n7804), .ZN(n8803) );
  XOR2_X1 U9372 ( .A(n7665), .B(n8323), .Z(n7666) );
  NAND2_X1 U9373 ( .A1(n7666), .A2(n8805), .ZN(n7668) );
  AOI22_X1 U9374 ( .A1(n8801), .A2(n8478), .B1(n8800), .B2(n8476), .ZN(n7667)
         );
  OAI211_X1 U9375 ( .C1(n8803), .C2(n10025), .A(n7668), .B(n7667), .ZN(n10027)
         );
  AOI211_X1 U9376 ( .C1(n7670), .C2(n8796), .A(n7669), .B(n10027), .ZN(n7671)
         );
  MUX2_X1 U9377 ( .A(n7043), .B(n7671), .S(n8812), .Z(n7672) );
  OAI21_X1 U9378 ( .B1(n10024), .B2(n8725), .A(n7672), .ZN(P2_U3226) );
  NOR2_X1 U9379 ( .A1(n9661), .A2(n9600), .ZN(n9345) );
  OAI21_X1 U9380 ( .B1(n9345), .B2(n9788), .A(n7673), .ZN(n7682) );
  NAND3_X1 U9381 ( .A1(n7676), .A2(n7675), .A3(n7674), .ZN(n7678) );
  OAI211_X1 U9382 ( .C1(n9513), .C2(n7679), .A(n7678), .B(n7677), .ZN(n7680)
         );
  NAND2_X1 U9383 ( .A1(n7680), .A2(n9516), .ZN(n7681) );
  OAI211_X1 U9384 ( .C1(n5565), .C2(n9516), .A(n7682), .B(n7681), .ZN(P1_U3293) );
  XOR2_X1 U9385 ( .A(n7683), .B(n7684), .Z(n9863) );
  XOR2_X1 U9386 ( .A(n7685), .B(n7684), .Z(n7688) );
  INV_X1 U9387 ( .A(n7686), .ZN(n7687) );
  AOI21_X1 U9388 ( .B1(n7688), .B2(n9782), .A(n7687), .ZN(n9861) );
  MUX2_X1 U9389 ( .A(n7689), .B(n9861), .S(n9516), .Z(n7695) );
  INV_X1 U9390 ( .A(n7690), .ZN(n9794) );
  AOI211_X1 U9391 ( .C1(n9859), .C2(n9794), .A(n9600), .B(n9775), .ZN(n9858)
         );
  OAI22_X1 U9392 ( .A1(n9500), .A2(n7692), .B1(n9513), .B2(n7691), .ZN(n7693)
         );
  AOI21_X1 U9393 ( .B1(n9858), .B2(n9757), .A(n7693), .ZN(n7694) );
  OAI211_X1 U9394 ( .C1(n9662), .C2(n9863), .A(n7695), .B(n7694), .ZN(P1_U3288) );
  OAI21_X1 U9395 ( .B1(n4615), .B2(n7697), .A(n7696), .ZN(n7698) );
  NAND2_X1 U9396 ( .A1(n7698), .A2(n8232), .ZN(n7704) );
  AOI21_X1 U9397 ( .B1(n8211), .B2(n8476), .A(n7699), .ZN(n7700) );
  OAI21_X1 U9398 ( .B1(n7701), .B2(n8223), .A(n7700), .ZN(n7702) );
  AOI21_X1 U9399 ( .B1(n8324), .B2(n8227), .A(n7702), .ZN(n7703) );
  OAI211_X1 U9400 ( .C1(n7705), .C2(n8165), .A(n7704), .B(n7703), .ZN(P2_U3153) );
  NAND2_X1 U9401 ( .A1(n7707), .A2(n7706), .ZN(n7759) );
  INV_X1 U9402 ( .A(n7708), .ZN(n9746) );
  NAND2_X1 U9403 ( .A1(n7710), .A2(n7709), .ZN(n9754) );
  INV_X1 U9404 ( .A(n9754), .ZN(n9744) );
  NAND3_X1 U9405 ( .A1(n9746), .A2(n9744), .A3(n9745), .ZN(n9743) );
  NAND2_X1 U9406 ( .A1(n9743), .A2(n7710), .ZN(n7711) );
  XOR2_X1 U9407 ( .A(n7759), .B(n7711), .Z(n7712) );
  NAND2_X1 U9408 ( .A1(n9193), .A2(n9131), .ZN(n9099) );
  OAI21_X1 U9409 ( .B1(n7712), .B2(n9765), .A(n9099), .ZN(n9886) );
  INV_X1 U9410 ( .A(n9886), .ZN(n7726) );
  NAND2_X1 U9411 ( .A1(n9873), .A2(n7715), .ZN(n7716) );
  NAND2_X1 U9412 ( .A1(n9753), .A2(n9754), .ZN(n7718) );
  OR2_X1 U9413 ( .A1(n9755), .A2(n9193), .ZN(n7717) );
  NAND2_X1 U9414 ( .A1(n7718), .A2(n7717), .ZN(n7760) );
  XNOR2_X1 U9415 ( .A(n7760), .B(n7759), .ZN(n9888) );
  AOI211_X1 U9416 ( .C1(n9883), .C2(n9756), .A(n9600), .B(n7756), .ZN(n7720)
         );
  NAND2_X1 U9417 ( .A1(n9191), .A2(n4509), .ZN(n9100) );
  INV_X1 U9418 ( .A(n9100), .ZN(n7719) );
  NOR2_X1 U9419 ( .A1(n7720), .A2(n7719), .ZN(n9884) );
  OAI22_X1 U9420 ( .A1(n9516), .A2(n7721), .B1(n9103), .B2(n9513), .ZN(n7722)
         );
  AOI21_X1 U9421 ( .B1(n9788), .B2(n9883), .A(n7722), .ZN(n7723) );
  OAI21_X1 U9422 ( .B1(n9884), .B2(n9661), .A(n7723), .ZN(n7724) );
  AOI21_X1 U9423 ( .B1(n9797), .B2(n9888), .A(n7724), .ZN(n7725) );
  OAI21_X1 U9424 ( .B1(n7726), .B2(n9785), .A(n7725), .ZN(P1_U3284) );
  OAI21_X1 U9425 ( .B1(n7729), .B2(n7727), .A(n7728), .ZN(n7736) );
  NOR2_X1 U9426 ( .A1(n9704), .A2(n9873), .ZN(n7735) );
  NAND2_X1 U9427 ( .A1(n9702), .A2(n7730), .ZN(n7732) );
  OAI211_X1 U9428 ( .C1(n9708), .C2(n7733), .A(n7732), .B(n7731), .ZN(n7734)
         );
  AOI211_X1 U9429 ( .C1(n7736), .C2(n9096), .A(n7735), .B(n7734), .ZN(n7737)
         );
  INV_X1 U9430 ( .A(n7737), .ZN(P1_U3213) );
  XOR2_X1 U9431 ( .A(n8272), .B(n7738), .Z(n7742) );
  INV_X1 U9432 ( .A(n7742), .ZN(n10036) );
  NAND2_X1 U9433 ( .A1(n8812), .A2(n8796), .ZN(n8619) );
  XNOR2_X1 U9434 ( .A(n7739), .B(n8272), .ZN(n7744) );
  OAI22_X1 U9435 ( .A1(n8748), .A2(n7740), .B1(n7920), .B2(n8779), .ZN(n7741)
         );
  AOI21_X1 U9436 ( .B1(n7742), .B2(n7804), .A(n7741), .ZN(n7743) );
  OAI21_X1 U9437 ( .B1(n8782), .B2(n7744), .A(n7743), .ZN(n10037) );
  NAND2_X1 U9438 ( .A1(n10037), .A2(n8812), .ZN(n7748) );
  INV_X1 U9439 ( .A(n7916), .ZN(n7745) );
  OAI22_X1 U9440 ( .A1(n8812), .A2(n7215), .B1(n7745), .B2(n8674), .ZN(n7746)
         );
  AOI21_X1 U9441 ( .B1(n4507), .B2(n10039), .A(n7746), .ZN(n7747) );
  OAI211_X1 U9442 ( .C1(n10036), .C2(n8619), .A(n7748), .B(n7747), .ZN(
        P2_U3224) );
  NAND2_X1 U9443 ( .A1(n7750), .A2(n7749), .ZN(n7751) );
  NAND2_X1 U9444 ( .A1(n7751), .A2(n7829), .ZN(n7752) );
  NAND2_X1 U9445 ( .A1(n7752), .A2(n7780), .ZN(n7755) );
  NAND2_X1 U9446 ( .A1(n9192), .A2(n9131), .ZN(n7754) );
  NAND2_X1 U9447 ( .A1(n9190), .A2(n4509), .ZN(n7753) );
  NAND2_X1 U9448 ( .A1(n7754), .A2(n7753), .ZN(n9641) );
  AOI21_X1 U9449 ( .B1(n7755), .B2(n9782), .A(n9641), .ZN(n9891) );
  OAI22_X1 U9450 ( .A1(n9516), .A2(n6962), .B1(n9646), .B2(n9513), .ZN(n7758)
         );
  INV_X1 U9451 ( .A(n7791), .ZN(n7792) );
  OAI211_X1 U9452 ( .C1(n9892), .C2(n7756), .A(n7792), .B(n9793), .ZN(n9890)
         );
  NOR2_X1 U9453 ( .A1(n9890), .A2(n9661), .ZN(n7757) );
  AOI211_X1 U9454 ( .C1(n9788), .C2(n7787), .A(n7758), .B(n7757), .ZN(n7762)
         );
  NAND2_X1 U9455 ( .A1(n7760), .A2(n7759), .ZN(n7826) );
  OR2_X1 U9456 ( .A1(n9883), .A2(n9192), .ZN(n7824) );
  NAND2_X1 U9457 ( .A1(n7826), .A2(n7824), .ZN(n7786) );
  XNOR2_X1 U9458 ( .A(n7786), .B(n7829), .ZN(n9894) );
  NAND2_X1 U9459 ( .A1(n9894), .A2(n9797), .ZN(n7761) );
  OAI211_X1 U9460 ( .C1(n9785), .C2(n9891), .A(n7762), .B(n7761), .ZN(P1_U3283) );
  XOR2_X1 U9461 ( .A(n7764), .B(n7763), .Z(n7772) );
  NAND2_X1 U9462 ( .A1(n8241), .A2(n7765), .ZN(n7768) );
  AOI21_X1 U9463 ( .B1(n8211), .B2(n8475), .A(n7766), .ZN(n7767) );
  OAI211_X1 U9464 ( .C1(n8325), .C2(n8223), .A(n7768), .B(n7767), .ZN(n7769)
         );
  AOI21_X1 U9465 ( .B1(n7770), .B2(n8227), .A(n7769), .ZN(n7771) );
  OAI21_X1 U9466 ( .B1(n7772), .B2(n8230), .A(n7771), .ZN(P2_U3161) );
  INV_X1 U9467 ( .A(n7773), .ZN(n7777) );
  OAI222_X1 U9468 ( .A1(n8965), .A2(n7777), .B1(P2_U3151), .B2(n7775), .C1(
        n7774), .C2(n8102), .ZN(P2_U3274) );
  OAI222_X1 U9469 ( .A1(P1_U3086), .A2(n7778), .B1(n9629), .B2(n7777), .C1(
        n7776), .C2(n9633), .ZN(P1_U3334) );
  NAND2_X1 U9470 ( .A1(n7780), .A2(n7779), .ZN(n7782) );
  INV_X1 U9471 ( .A(n7815), .ZN(n7781) );
  AOI211_X1 U9472 ( .C1(n7790), .C2(n7782), .A(n9765), .B(n7781), .ZN(n7785)
         );
  NAND2_X1 U9473 ( .A1(n9189), .A2(n4509), .ZN(n7784) );
  NAND2_X1 U9474 ( .A1(n9191), .A2(n9131), .ZN(n7783) );
  NAND2_X1 U9475 ( .A1(n7784), .A2(n7783), .ZN(n9143) );
  NOR2_X1 U9476 ( .A1(n7785), .A2(n9143), .ZN(n9900) );
  NAND2_X1 U9477 ( .A1(n7786), .A2(n7829), .ZN(n7788) );
  OR2_X1 U9478 ( .A1(n7787), .A2(n9191), .ZN(n7821) );
  NAND2_X1 U9479 ( .A1(n7788), .A2(n7821), .ZN(n7789) );
  XOR2_X1 U9480 ( .A(n7790), .B(n7789), .Z(n9902) );
  INV_X1 U9481 ( .A(n9902), .ZN(n9904) );
  NAND2_X1 U9482 ( .A1(n9904), .A2(n9797), .ZN(n7798) );
  INV_X1 U9483 ( .A(n9897), .ZN(n7793) );
  AND2_X2 U9484 ( .A1(n7791), .A2(n7793), .ZN(n7834) );
  AOI211_X1 U9485 ( .C1(n9897), .C2(n7792), .A(n9600), .B(n7834), .ZN(n9896)
         );
  NOR2_X1 U9486 ( .A1(n7793), .A2(n9500), .ZN(n7796) );
  OAI22_X1 U9487 ( .A1(n9516), .A2(n7794), .B1(n9145), .B2(n9513), .ZN(n7795)
         );
  AOI211_X1 U9488 ( .C1(n9896), .C2(n9757), .A(n7796), .B(n7795), .ZN(n7797)
         );
  OAI211_X1 U9489 ( .C1(n9785), .C2(n9900), .A(n7798), .B(n7797), .ZN(P1_U3282) );
  XNOR2_X1 U9490 ( .A(n7799), .B(n7801), .ZN(n7805) );
  INV_X1 U9491 ( .A(n7805), .ZN(n10042) );
  INV_X1 U9492 ( .A(n7801), .ZN(n8273) );
  XNOR2_X1 U9493 ( .A(n7800), .B(n8273), .ZN(n7807) );
  OAI22_X1 U9494 ( .A1(n8748), .A2(n7802), .B1(n7934), .B2(n8779), .ZN(n7803)
         );
  AOI21_X1 U9495 ( .B1(n7805), .B2(n7804), .A(n7803), .ZN(n7806) );
  OAI21_X1 U9496 ( .B1(n7807), .B2(n8782), .A(n7806), .ZN(n10043) );
  NAND2_X1 U9497 ( .A1(n10043), .A2(n8812), .ZN(n7811) );
  INV_X1 U9498 ( .A(n7930), .ZN(n7808) );
  OAI22_X1 U9499 ( .A1(n8812), .A2(n7337), .B1(n7808), .B2(n8674), .ZN(n7809)
         );
  AOI21_X1 U9500 ( .B1(n4507), .B2(n10045), .A(n7809), .ZN(n7810) );
  OAI211_X1 U9501 ( .C1(n10042), .C2(n8619), .A(n7811), .B(n7810), .ZN(
        P2_U3223) );
  INV_X1 U9502 ( .A(n7812), .ZN(n7813) );
  NOR2_X1 U9503 ( .A1(n7832), .A2(n7813), .ZN(n7814) );
  AOI21_X1 U9504 ( .B1(n7815), .B2(n7814), .A(n9765), .ZN(n7818) );
  NAND2_X1 U9505 ( .A1(n9188), .A2(n4509), .ZN(n7817) );
  NAND2_X1 U9506 ( .A1(n9190), .A2(n9131), .ZN(n7816) );
  NAND2_X1 U9507 ( .A1(n7817), .A2(n7816), .ZN(n9046) );
  AOI21_X1 U9508 ( .B1(n7819), .B2(n7818), .A(n9046), .ZN(n9907) );
  NAND2_X1 U9509 ( .A1(n9897), .A2(n9190), .ZN(n7828) );
  INV_X1 U9510 ( .A(n7828), .ZN(n7823) );
  OR2_X1 U9511 ( .A1(n9897), .A2(n9190), .ZN(n7820) );
  AND2_X1 U9512 ( .A1(n7821), .A2(n7820), .ZN(n7822) );
  AND2_X1 U9513 ( .A1(n7824), .A2(n7827), .ZN(n7825) );
  NAND2_X1 U9514 ( .A1(n7826), .A2(n7825), .ZN(n7831) );
  XNOR2_X1 U9515 ( .A(n7873), .B(n7832), .ZN(n9909) );
  NAND2_X1 U9516 ( .A1(n9909), .A2(n9797), .ZN(n7838) );
  OAI22_X1 U9517 ( .A1(n9516), .A2(n7833), .B1(n9049), .B2(n9513), .ZN(n7836)
         );
  OAI211_X1 U9518 ( .C1(n7834), .C2(n5062), .A(n9793), .B(n7876), .ZN(n9906)
         );
  NOR2_X1 U9519 ( .A1(n9906), .A2(n9661), .ZN(n7835) );
  AOI211_X1 U9520 ( .C1(n9788), .C2(n9051), .A(n7836), .B(n7835), .ZN(n7837)
         );
  OAI211_X1 U9521 ( .C1(n9785), .C2(n9907), .A(n7838), .B(n7837), .ZN(P1_U3281) );
  NAND2_X1 U9522 ( .A1(n7728), .A2(n7839), .ZN(n9093) );
  XNOR2_X1 U9523 ( .A(n9093), .B(n9094), .ZN(n7841) );
  NOR2_X1 U9524 ( .A1(n7841), .A2(n7840), .ZN(n9092) );
  AOI21_X1 U9525 ( .B1(n7841), .B2(n7840), .A(n9092), .ZN(n7849) );
  NAND2_X1 U9526 ( .A1(n9697), .A2(n9131), .ZN(n7843) );
  NAND2_X1 U9527 ( .A1(n9192), .A2(n4509), .ZN(n7842) );
  NAND2_X1 U9528 ( .A1(n7843), .A2(n7842), .ZN(n9749) );
  INV_X1 U9529 ( .A(n7844), .ZN(n7845) );
  AOI21_X1 U9530 ( .B1(n9702), .B2(n9749), .A(n7845), .ZN(n7846) );
  OAI21_X1 U9531 ( .B1(n9751), .B2(n9708), .A(n7846), .ZN(n7847) );
  AOI21_X1 U9532 ( .B1(n9755), .B2(n6200), .A(n7847), .ZN(n7848) );
  OAI21_X1 U9533 ( .B1(n7849), .B2(n9693), .A(n7848), .ZN(P1_U3221) );
  XOR2_X1 U9534 ( .A(n7857), .B(n9284), .Z(n7853) );
  NOR2_X1 U9535 ( .A1(n7957), .A2(n7853), .ZN(n9285) );
  INV_X1 U9536 ( .A(n9285), .ZN(n7851) );
  NAND2_X1 U9537 ( .A1(n9720), .A2(n7851), .ZN(n7852) );
  AOI21_X1 U9538 ( .B1(n7853), .B2(n7957), .A(n7852), .ZN(n7863) );
  INV_X1 U9539 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9683) );
  NOR2_X1 U9540 ( .A1(n9683), .A2(n7856), .ZN(n9275) );
  AOI211_X1 U9541 ( .C1(n7856), .C2(n9683), .A(n9275), .B(n9727), .ZN(n7862)
         );
  INV_X1 U9542 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7860) );
  NAND2_X1 U9543 ( .A1(n9724), .A2(n7857), .ZN(n7859) );
  NAND2_X1 U9544 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n7858) );
  OAI211_X1 U9545 ( .C1(n7860), .C2(n9344), .A(n7859), .B(n7858), .ZN(n7861)
         );
  OR3_X1 U9546 ( .A1(n7863), .A2(n7862), .A3(n7861), .ZN(P1_U3258) );
  INV_X1 U9547 ( .A(n7864), .ZN(n7867) );
  OAI222_X1 U9548 ( .A1(n9633), .A2(n7865), .B1(n9629), .B2(n7867), .C1(
        P1_U3086), .C2(n5956), .ZN(P1_U3333) );
  OAI222_X1 U9549 ( .A1(n8102), .A2(n7868), .B1(n8965), .B2(n7867), .C1(n7866), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  XNOR2_X1 U9550 ( .A(n7869), .B(n7874), .ZN(n7872) );
  NAND2_X1 U9551 ( .A1(n9189), .A2(n9131), .ZN(n7871) );
  NAND2_X1 U9552 ( .A1(n9187), .A2(n4509), .ZN(n7870) );
  NAND2_X1 U9553 ( .A1(n7871), .A2(n7870), .ZN(n9121) );
  AOI21_X1 U9554 ( .B1(n7872), .B2(n9782), .A(n9121), .ZN(n9912) );
  XNOR2_X1 U9555 ( .A(n7953), .B(n7874), .ZN(n9917) );
  NAND2_X1 U9556 ( .A1(n9917), .A2(n9797), .ZN(n7881) );
  INV_X1 U9557 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7875) );
  OAI22_X1 U9558 ( .A1(n9516), .A2(n7875), .B1(n9123), .B2(n9513), .ZN(n7879)
         );
  INV_X1 U9559 ( .A(n7876), .ZN(n7877) );
  INV_X1 U9560 ( .A(n9125), .ZN(n9914) );
  OAI211_X1 U9561 ( .C1(n7877), .C2(n9914), .A(n9793), .B(n9601), .ZN(n9911)
         );
  NOR2_X1 U9562 ( .A1(n9911), .A2(n9661), .ZN(n7878) );
  AOI211_X1 U9563 ( .C1(n9788), .C2(n9125), .A(n7879), .B(n7878), .ZN(n7880)
         );
  OAI211_X1 U9564 ( .C1(n9785), .C2(n9912), .A(n7881), .B(n7880), .ZN(P1_U3280) );
  NAND2_X1 U9565 ( .A1(n7882), .A2(n8328), .ZN(n7883) );
  XNOR2_X1 U9566 ( .A(n7883), .B(n8275), .ZN(n7896) );
  INV_X1 U9567 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7886) );
  XOR2_X1 U9568 ( .A(n7884), .B(n8275), .Z(n7885) );
  AOI222_X1 U9569 ( .A1(n8805), .A2(n7885), .B1(n8472), .B2(n8800), .C1(n8474), 
        .C2(n8801), .ZN(n7892) );
  MUX2_X1 U9570 ( .A(n7886), .B(n7892), .S(n10047), .Z(n7888) );
  NAND2_X1 U9571 ( .A1(n8943), .A2(n7973), .ZN(n7887) );
  OAI211_X1 U9572 ( .C1(n7896), .C2(n8947), .A(n7888), .B(n7887), .ZN(P2_U3423) );
  MUX2_X1 U9573 ( .A(n7889), .B(n7892), .S(n10466), .Z(n7891) );
  NAND2_X1 U9574 ( .A1(n8859), .A2(n7973), .ZN(n7890) );
  OAI211_X1 U9575 ( .C1(n8862), .C2(n7896), .A(n7891), .B(n7890), .ZN(P2_U3470) );
  MUX2_X1 U9576 ( .A(n7893), .B(n7892), .S(n8812), .Z(n7895) );
  AOI22_X1 U9577 ( .A1(n4507), .A2(n7973), .B1(n8808), .B2(n7980), .ZN(n7894)
         );
  OAI211_X1 U9578 ( .C1(n7896), .C2(n8793), .A(n7895), .B(n7894), .ZN(P2_U3222) );
  XNOR2_X1 U9579 ( .A(n7897), .B(n8352), .ZN(n7909) );
  INV_X1 U9580 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7900) );
  XNOR2_X1 U9581 ( .A(n7898), .B(n8352), .ZN(n7899) );
  AOI222_X1 U9582 ( .A1(n8805), .A2(n7899), .B1(n8471), .B2(n8800), .C1(n8473), 
        .C2(n8801), .ZN(n7905) );
  MUX2_X1 U9583 ( .A(n7900), .B(n7905), .S(n10047), .Z(n7902) );
  NAND2_X1 U9584 ( .A1(n8943), .A2(n8012), .ZN(n7901) );
  OAI211_X1 U9585 ( .C1(n7909), .C2(n8947), .A(n7902), .B(n7901), .ZN(P2_U3426) );
  MUX2_X1 U9586 ( .A(n8489), .B(n7905), .S(n10466), .Z(n7904) );
  NAND2_X1 U9587 ( .A1(n8012), .A2(n8859), .ZN(n7903) );
  OAI211_X1 U9588 ( .C1(n7909), .C2(n8862), .A(n7904), .B(n7903), .ZN(P2_U3471) );
  MUX2_X1 U9589 ( .A(n7906), .B(n7905), .S(n8812), .Z(n7908) );
  AOI22_X1 U9590 ( .A1(n8012), .A2(n4507), .B1(n8808), .B2(n8019), .ZN(n7907)
         );
  OAI211_X1 U9591 ( .C1(n7909), .C2(n8793), .A(n7908), .B(n7907), .ZN(P2_U3221) );
  NAND2_X1 U9592 ( .A1(n7914), .A2(n9625), .ZN(n7911) );
  OAI211_X1 U9593 ( .C1(n7912), .C2(n9633), .A(n7911), .B(n7910), .ZN(P1_U3332) );
  NAND2_X1 U9594 ( .A1(n7914), .A2(n7913), .ZN(n7915) );
  OAI211_X1 U9595 ( .C1(n10214), .C2(n8102), .A(n7915), .B(n8465), .ZN(
        P2_U3272) );
  NAND2_X1 U9596 ( .A1(n8241), .A2(n7916), .ZN(n7919) );
  AOI21_X1 U9597 ( .B1(n8211), .B2(n8474), .A(n7917), .ZN(n7918) );
  OAI211_X1 U9598 ( .C1(n7920), .C2(n8223), .A(n7919), .B(n7918), .ZN(n7926)
         );
  INV_X1 U9599 ( .A(n7921), .ZN(n7922) );
  AOI211_X1 U9600 ( .C1(n7924), .C2(n7923), .A(n8230), .B(n7922), .ZN(n7925)
         );
  AOI211_X1 U9601 ( .C1(n10039), .C2(n8227), .A(n7926), .B(n7925), .ZN(n7927)
         );
  INV_X1 U9602 ( .A(n7927), .ZN(P2_U3171) );
  XOR2_X1 U9603 ( .A(n7928), .B(n7929), .Z(n7937) );
  NAND2_X1 U9604 ( .A1(n8241), .A2(n7930), .ZN(n7933) );
  AOI21_X1 U9605 ( .B1(n8211), .B2(n8473), .A(n7931), .ZN(n7932) );
  OAI211_X1 U9606 ( .C1(n7934), .C2(n8223), .A(n7933), .B(n7932), .ZN(n7935)
         );
  AOI21_X1 U9607 ( .B1(n10045), .B2(n8227), .A(n7935), .ZN(n7936) );
  OAI21_X1 U9608 ( .B1(n7937), .B2(n8230), .A(n7936), .ZN(P2_U3157) );
  INV_X1 U9609 ( .A(n7938), .ZN(n7964) );
  OAI222_X1 U9610 ( .A1(n8965), .A2(n7964), .B1(P2_U3151), .B2(n7940), .C1(
        n7939), .C2(n8102), .ZN(P2_U3271) );
  XNOR2_X1 U9611 ( .A(n8358), .B(n8471), .ZN(n8276) );
  XOR2_X1 U9612 ( .A(n8276), .B(n7941), .Z(n7942) );
  AOI222_X1 U9613 ( .A1(n8805), .A2(n7942), .B1(n8472), .B2(n8801), .C1(n8470), 
        .C2(n8800), .ZN(n7969) );
  INV_X1 U9614 ( .A(n8676), .ZN(n8807) );
  AOI22_X1 U9615 ( .A1(n8358), .A2(n8807), .B1(n8808), .B2(n8194), .ZN(n7943)
         );
  AOI21_X1 U9616 ( .B1(n7969), .B2(n7943), .A(n8771), .ZN(n7946) );
  XNOR2_X1 U9617 ( .A(n7944), .B(n8276), .ZN(n7972) );
  INV_X1 U9618 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10217) );
  OAI22_X1 U9619 ( .A1(n7972), .A2(n8793), .B1(n10217), .B2(n8812), .ZN(n7945)
         );
  OR2_X1 U9620 ( .A1(n7946), .A2(n7945), .ZN(P2_U3220) );
  NAND2_X1 U9621 ( .A1(n9595), .A2(n7947), .ZN(n7948) );
  XNOR2_X1 U9622 ( .A(n7948), .B(n7956), .ZN(n7951) );
  NAND2_X1 U9623 ( .A1(n9187), .A2(n9131), .ZN(n7950) );
  NAND2_X1 U9624 ( .A1(n9185), .A2(n4509), .ZN(n7949) );
  NAND2_X1 U9625 ( .A1(n7950), .A2(n7949), .ZN(n9163) );
  AOI21_X1 U9626 ( .B1(n7951), .B2(n9782), .A(n9163), .ZN(n9679) );
  NOR2_X1 U9627 ( .A1(n9125), .A2(n9188), .ZN(n7952) );
  NAND2_X1 U9628 ( .A1(n9125), .A2(n9188), .ZN(n9591) );
  AND2_X1 U9629 ( .A1(n9597), .A2(n9591), .ZN(n7954) );
  OR2_X1 U9630 ( .A1(n9735), .A2(n9187), .ZN(n7955) );
  XNOR2_X1 U9631 ( .A(n8044), .B(n7956), .ZN(n9682) );
  NAND2_X1 U9632 ( .A1(n9682), .A2(n9797), .ZN(n7962) );
  OAI22_X1 U9633 ( .A1(n9516), .A2(n7957), .B1(n9165), .B2(n9513), .ZN(n7960)
         );
  INV_X1 U9634 ( .A(n9168), .ZN(n9680) );
  INV_X1 U9635 ( .A(n9660), .ZN(n7958) );
  OAI211_X1 U9636 ( .C1(n9680), .C2(n4595), .A(n7958), .B(n9793), .ZN(n9678)
         );
  NOR2_X1 U9637 ( .A1(n9678), .A2(n9661), .ZN(n7959) );
  AOI211_X1 U9638 ( .C1(n9788), .C2(n9168), .A(n7960), .B(n7959), .ZN(n7961)
         );
  OAI211_X1 U9639 ( .C1(n9785), .C2(n9679), .A(n7962), .B(n7961), .ZN(P1_U3278) );
  OAI222_X1 U9640 ( .A1(n7965), .A2(P1_U3086), .B1(n9629), .B2(n7964), .C1(
        n7963), .C2(n9633), .ZN(P1_U3331) );
  INV_X1 U9641 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7966) );
  MUX2_X1 U9642 ( .A(n7966), .B(n7969), .S(n10047), .Z(n7968) );
  NAND2_X1 U9643 ( .A1(n8358), .A2(n8943), .ZN(n7967) );
  OAI211_X1 U9644 ( .C1(n7972), .C2(n8947), .A(n7968), .B(n7967), .ZN(P2_U3429) );
  INV_X1 U9645 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10309) );
  MUX2_X1 U9646 ( .A(n10309), .B(n7969), .S(n10466), .Z(n7971) );
  NAND2_X1 U9647 ( .A1(n8358), .A2(n8859), .ZN(n7970) );
  OAI211_X1 U9648 ( .C1(n8862), .C2(n7972), .A(n7971), .B(n7970), .ZN(P2_U3472) );
  INV_X1 U9649 ( .A(n7973), .ZN(n7983) );
  OAI211_X1 U9650 ( .C1(n7976), .C2(n6715), .A(n8232), .B(n7975), .ZN(n7982)
         );
  NAND2_X1 U9651 ( .A1(n8236), .A2(n8474), .ZN(n7978) );
  OAI211_X1 U9652 ( .C1(n8197), .C2(n8238), .A(n7978), .B(n7977), .ZN(n7979)
         );
  AOI21_X1 U9653 ( .B1(n7980), .B2(n8241), .A(n7979), .ZN(n7981) );
  OAI211_X1 U9654 ( .C1(n7983), .C2(n8245), .A(n7982), .B(n7981), .ZN(P2_U3176) );
  INV_X1 U9655 ( .A(n7984), .ZN(n8367) );
  XNOR2_X1 U9656 ( .A(n7985), .B(n8364), .ZN(n7986) );
  AOI222_X1 U9657 ( .A1(n8805), .A2(n7986), .B1(n8469), .B2(n8800), .C1(n8471), 
        .C2(n8801), .ZN(n7996) );
  AOI22_X1 U9658 ( .A1(n8118), .A2(n8807), .B1(n8808), .B2(n8113), .ZN(n7987)
         );
  AOI21_X1 U9659 ( .B1(n7996), .B2(n7987), .A(n8771), .ZN(n7990) );
  XOR2_X1 U9660 ( .A(n8364), .B(n7988), .Z(n7999) );
  INV_X1 U9661 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8500) );
  OAI22_X1 U9662 ( .A1(n7999), .A2(n8793), .B1(n8500), .B2(n8812), .ZN(n7989)
         );
  OR2_X1 U9663 ( .A1(n7990), .A2(n7989), .ZN(P2_U3219) );
  INV_X1 U9664 ( .A(n7991), .ZN(n8001) );
  INV_X1 U9665 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10280) );
  MUX2_X1 U9666 ( .A(n10280), .B(n7996), .S(n10047), .Z(n7995) );
  NAND2_X1 U9667 ( .A1(n8118), .A2(n8943), .ZN(n7994) );
  OAI211_X1 U9668 ( .C1(n7999), .C2(n8947), .A(n7995), .B(n7994), .ZN(P2_U3432) );
  INV_X1 U9669 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8499) );
  MUX2_X1 U9670 ( .A(n8499), .B(n7996), .S(n10466), .Z(n7998) );
  NAND2_X1 U9671 ( .A1(n8118), .A2(n8859), .ZN(n7997) );
  OAI211_X1 U9672 ( .C1(n8862), .C2(n7999), .A(n7998), .B(n7997), .ZN(P2_U3473) );
  OAI222_X1 U9673 ( .A1(n8002), .A2(P1_U3086), .B1(n9629), .B2(n8001), .C1(
        n8000), .C2(n9633), .ZN(P1_U3330) );
  XNOR2_X1 U9674 ( .A(n8003), .B(n4512), .ZN(n8004) );
  OAI222_X1 U9675 ( .A1(n8748), .A2(n8239), .B1(n8779), .B2(n8005), .C1(n8782), 
        .C2(n8004), .ZN(n8863) );
  INV_X1 U9676 ( .A(n8863), .ZN(n8011) );
  OAI21_X1 U9677 ( .B1(n4604), .B2(n4512), .A(n8006), .ZN(n8864) );
  INV_X1 U9678 ( .A(n8007), .ZN(n8953) );
  AOI22_X1 U9679 ( .A1(n8771), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8808), .B2(
        n8242), .ZN(n8008) );
  OAI21_X1 U9680 ( .B1(n8953), .B2(n8725), .A(n8008), .ZN(n8009) );
  AOI21_X1 U9681 ( .B1(n8864), .B2(n8727), .A(n8009), .ZN(n8010) );
  OAI21_X1 U9682 ( .B1(n8011), .B2(n8771), .A(n8010), .ZN(P2_U3218) );
  OAI211_X1 U9683 ( .C1(n8015), .C2(n8014), .A(n8013), .B(n8232), .ZN(n8021)
         );
  NAND2_X1 U9684 ( .A1(n8236), .A2(n8473), .ZN(n8017) );
  OAI211_X1 U9685 ( .C1(n8116), .C2(n8238), .A(n8017), .B(n8016), .ZN(n8018)
         );
  AOI21_X1 U9686 ( .B1(n8019), .B2(n8241), .A(n8018), .ZN(n8020) );
  OAI211_X1 U9687 ( .C1(n4974), .C2(n8245), .A(n8021), .B(n8020), .ZN(P2_U3164) );
  INV_X1 U9688 ( .A(n8022), .ZN(n8026) );
  OAI222_X1 U9689 ( .A1(n8965), .A2(n8026), .B1(P2_U3151), .B2(n8024), .C1(
        n8023), .C2(n8102), .ZN(P2_U3269) );
  INV_X1 U9690 ( .A(n6161), .ZN(n8027) );
  OAI222_X1 U9691 ( .A1(n8027), .A2(P1_U3086), .B1(n9629), .B2(n8026), .C1(
        n8025), .C2(n9633), .ZN(P1_U3329) );
  OAI222_X1 U9692 ( .A1(n8965), .A2(n9631), .B1(n8028), .B2(P2_U3151), .C1(
        n10238), .C2(n8102), .ZN(P2_U3266) );
  INV_X1 U9693 ( .A(P1_B_REG_SCAN_IN), .ZN(n8029) );
  OR2_X1 U9694 ( .A1(n4511), .A2(n8029), .ZN(n8030) );
  NAND2_X1 U9695 ( .A1(n4509), .A2(n8030), .ZN(n9346) );
  NAND2_X1 U9696 ( .A1(n9458), .A2(n8031), .ZN(n9450) );
  NAND2_X1 U9697 ( .A1(n9394), .A2(n9392), .ZN(n8034) );
  OAI21_X1 U9698 ( .B1(n9407), .B2(n8034), .A(n8033), .ZN(n8087) );
  NAND2_X1 U9699 ( .A1(n8087), .A2(n8088), .ZN(n8086) );
  OAI222_X1 U9700 ( .A1(n9346), .A2(n8041), .B1(n8040), .B2(n8068), .C1(n8039), 
        .C2(n9765), .ZN(n9533) );
  INV_X1 U9701 ( .A(n9572), .ZN(n9448) );
  NAND2_X1 U9702 ( .A1(n9168), .A2(n9186), .ZN(n8043) );
  NOR2_X1 U9703 ( .A1(n9168), .A2(n9186), .ZN(n8042) );
  AOI21_X1 U9704 ( .B1(n9185), .B2(n9654), .A(n9658), .ZN(n9512) );
  INV_X1 U9705 ( .A(n9512), .ZN(n8045) );
  AOI21_X1 U9706 ( .B1(n8045), .B2(n9184), .A(n9521), .ZN(n8046) );
  AOI21_X1 U9707 ( .B1(n9512), .B2(n8047), .A(n8046), .ZN(n9486) );
  NAND2_X1 U9708 ( .A1(n9486), .A2(n8048), .ZN(n8050) );
  NAND2_X1 U9709 ( .A1(n8054), .A2(n5115), .ZN(n9443) );
  AOI21_X1 U9710 ( .B1(n9180), .B2(n9572), .A(n9443), .ZN(n8055) );
  NOR2_X1 U9711 ( .A1(n9406), .A2(n8061), .ZN(n8062) );
  NOR2_X1 U9712 ( .A1(n9552), .A2(n9176), .ZN(n8064) );
  NAND2_X1 U9713 ( .A1(n9552), .A2(n9176), .ZN(n8063) );
  NOR2_X1 U9714 ( .A1(n8085), .A2(n8065), .ZN(n8066) );
  NOR2_X1 U9715 ( .A1(n9543), .A2(n9174), .ZN(n8067) );
  INV_X1 U9716 ( .A(n9538), .ZN(n9371) );
  NAND2_X1 U9717 ( .A1(n9371), .A2(n8068), .ZN(n8069) );
  AOI22_X1 U9718 ( .A1(n9359), .A2(n8069), .B1(n9538), .B2(n9173), .ZN(n8071)
         );
  XNOR2_X1 U9719 ( .A(n8071), .B(n8070), .ZN(n9531) );
  NAND2_X1 U9720 ( .A1(n9531), .A2(n9797), .ZN(n8078) );
  INV_X1 U9721 ( .A(n9654), .ZN(n9674) );
  NAND2_X1 U9722 ( .A1(n9660), .A2(n9674), .ZN(n9659) );
  NOR2_X2 U9723 ( .A1(n9463), .A2(n9572), .ZN(n9444) );
  NAND2_X1 U9724 ( .A1(n9388), .A2(n8085), .ZN(n9380) );
  NOR2_X2 U9725 ( .A1(n9380), .A2(n9543), .ZN(n9379) );
  NOR2_X2 U9726 ( .A1(n9364), .A2(n9532), .ZN(n9353) );
  INV_X1 U9727 ( .A(n9532), .ZN(n8072) );
  NOR2_X1 U9728 ( .A1(n8072), .A2(n9500), .ZN(n8076) );
  OAI22_X1 U9729 ( .A1(n8074), .A2(n9513), .B1(n8073), .B2(n9516), .ZN(n8075)
         );
  AOI211_X1 U9730 ( .C1(n9534), .C2(n9757), .A(n8076), .B(n8075), .ZN(n8077)
         );
  OAI211_X1 U9731 ( .C1(n4766), .C2(n9785), .A(n8078), .B(n8077), .ZN(P1_U3356) );
  XOR2_X1 U9732 ( .A(n8088), .B(n8079), .Z(n9550) );
  INV_X1 U9733 ( .A(n9388), .ZN(n8081) );
  INV_X1 U9734 ( .A(n9380), .ZN(n8080) );
  AOI21_X1 U9735 ( .B1(n9546), .B2(n8081), .A(n8080), .ZN(n9547) );
  INV_X1 U9736 ( .A(n8082), .ZN(n8083) );
  AOI22_X1 U9737 ( .A1(n8083), .A2(n9786), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9785), .ZN(n8084) );
  OAI21_X1 U9738 ( .B1(n8085), .B2(n9500), .A(n8084), .ZN(n8092) );
  OAI21_X1 U9739 ( .B1(n8088), .B2(n8087), .A(n8086), .ZN(n8090) );
  AOI21_X1 U9740 ( .B1(n8090), .B2(n9782), .A(n8089), .ZN(n9549) );
  NOR2_X1 U9741 ( .A1(n9549), .A2(n9785), .ZN(n8091) );
  AOI211_X1 U9742 ( .C1(n9547), .C2(n9345), .A(n8092), .B(n8091), .ZN(n8093)
         );
  OAI21_X1 U9743 ( .B1(n9550), .B2(n9662), .A(n8093), .ZN(P1_U3267) );
  INV_X1 U9744 ( .A(n8094), .ZN(n8961) );
  INV_X1 U9745 ( .A(n8096), .ZN(n8966) );
  OAI222_X1 U9746 ( .A1(n9633), .A2(n10342), .B1(P1_U3086), .B2(n4511), .C1(
        n8966), .C2(n9629), .ZN(P1_U3328) );
  OAI222_X1 U9747 ( .A1(n9633), .A2(n8100), .B1(n9629), .B2(n8099), .C1(
        P1_U3086), .C2(n8097), .ZN(P1_U3336) );
  INV_X1 U9748 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8246) );
  INV_X1 U9749 ( .A(n8248), .ZN(n9628) );
  OAI222_X1 U9750 ( .A1(n8102), .A2(n8246), .B1(n8965), .B2(n9628), .C1(
        P2_U3151), .C2(n8101), .ZN(P2_U3265) );
  XNOR2_X1 U9751 ( .A(n8103), .B(n8104), .ZN(n8110) );
  OAI22_X1 U9752 ( .A1(n8635), .A2(n8223), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8105), .ZN(n8107) );
  NOR2_X1 U9753 ( .A1(n8636), .A2(n8238), .ZN(n8106) );
  AOI211_X1 U9754 ( .C1(n8640), .C2(n8241), .A(n8107), .B(n8106), .ZN(n8109)
         );
  NAND2_X1 U9755 ( .A1(n8884), .A2(n8227), .ZN(n8108) );
  OAI211_X1 U9756 ( .C1(n8110), .C2(n8230), .A(n8109), .B(n8108), .ZN(P2_U3154) );
  XOR2_X1 U9757 ( .A(n8112), .B(n8111), .Z(n8120) );
  NAND2_X1 U9758 ( .A1(n8241), .A2(n8113), .ZN(n8115) );
  AOI22_X1 U9759 ( .A1(n8211), .A2(n8469), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n8114) );
  OAI211_X1 U9760 ( .C1(n8116), .C2(n8223), .A(n8115), .B(n8114), .ZN(n8117)
         );
  AOI21_X1 U9761 ( .B1(n8118), .B2(n8227), .A(n8117), .ZN(n8119) );
  OAI21_X1 U9762 ( .B1(n8120), .B2(n8230), .A(n8119), .ZN(P2_U3155) );
  XNOR2_X1 U9763 ( .A(n8172), .B(n8171), .ZN(n8173) );
  XNOR2_X1 U9764 ( .A(n8173), .B(n8205), .ZN(n8125) );
  NAND2_X1 U9765 ( .A1(n8241), .A2(n8689), .ZN(n8122) );
  AOI22_X1 U9766 ( .A1(n8236), .A2(n8686), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8121) );
  OAI211_X1 U9767 ( .C1(n8174), .C2(n8238), .A(n8122), .B(n8121), .ZN(n8123)
         );
  AOI21_X1 U9768 ( .B1(n8908), .B2(n8227), .A(n8123), .ZN(n8124) );
  OAI21_X1 U9769 ( .B1(n8125), .B2(n8230), .A(n8124), .ZN(P2_U3156) );
  XOR2_X1 U9770 ( .A(n8127), .B(n8126), .Z(n8132) );
  NAND2_X1 U9771 ( .A1(n8211), .A2(n8732), .ZN(n8128) );
  NAND2_X1 U9772 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8598) );
  OAI211_X1 U9773 ( .C1(n8164), .C2(n8223), .A(n8128), .B(n8598), .ZN(n8129)
         );
  AOI21_X1 U9774 ( .B1(n8738), .B2(n8241), .A(n8129), .ZN(n8131) );
  NAND2_X1 U9775 ( .A1(n8850), .A2(n8227), .ZN(n8130) );
  OAI211_X1 U9776 ( .C1(n8132), .C2(n8230), .A(n8131), .B(n8130), .ZN(P2_U3159) );
  XOR2_X1 U9777 ( .A(n8134), .B(n8133), .Z(n8140) );
  NOR2_X1 U9778 ( .A1(n8223), .A2(n8705), .ZN(n8137) );
  OAI22_X1 U9779 ( .A1(n8238), .A2(n8704), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8135), .ZN(n8136) );
  AOI211_X1 U9780 ( .C1(n8241), .C2(n8709), .A(n8137), .B(n8136), .ZN(n8139)
         );
  NAND2_X1 U9781 ( .A1(n8708), .A2(n8227), .ZN(n8138) );
  OAI211_X1 U9782 ( .C1(n8140), .C2(n8230), .A(n8139), .B(n8138), .ZN(P2_U3163) );
  XOR2_X1 U9783 ( .A(n8142), .B(n8141), .Z(n8148) );
  NOR2_X1 U9784 ( .A1(n8174), .A2(n8223), .ZN(n8145) );
  OAI22_X1 U9785 ( .A1(n8635), .A2(n8238), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8143), .ZN(n8144) );
  AOI211_X1 U9786 ( .C1(n8659), .C2(n8241), .A(n8145), .B(n8144), .ZN(n8147)
         );
  NAND2_X1 U9787 ( .A1(n8896), .A2(n8227), .ZN(n8146) );
  OAI211_X1 U9788 ( .C1(n8148), .C2(n8230), .A(n8147), .B(n8146), .ZN(P2_U3165) );
  INV_X1 U9789 ( .A(n8149), .ZN(n8160) );
  AOI21_X1 U9790 ( .B1(n8151), .B2(n8150), .A(n8160), .ZN(n8156) );
  NAND2_X1 U9791 ( .A1(n8241), .A2(n8789), .ZN(n8153) );
  AOI22_X1 U9792 ( .A1(n8211), .A2(n8787), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3151), .ZN(n8152) );
  OAI211_X1 U9793 ( .C1(n8778), .C2(n8223), .A(n8153), .B(n8152), .ZN(n8154)
         );
  AOI21_X1 U9794 ( .B1(n8944), .B2(n8227), .A(n8154), .ZN(n8155) );
  OAI21_X1 U9795 ( .B1(n8156), .B2(n8230), .A(n8155), .ZN(P2_U3166) );
  INV_X1 U9796 ( .A(n8937), .ZN(n8170) );
  INV_X1 U9797 ( .A(n8157), .ZN(n8159) );
  NOR3_X1 U9798 ( .A1(n8160), .A2(n8159), .A3(n8158), .ZN(n8163) );
  INV_X1 U9799 ( .A(n8161), .ZN(n8162) );
  OAI21_X1 U9800 ( .B1(n8163), .B2(n8162), .A(n8232), .ZN(n8169) );
  OAI22_X1 U9801 ( .A1(n8238), .A2(n8164), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10348), .ZN(n8167) );
  NOR2_X1 U9802 ( .A1(n8165), .A2(n8773), .ZN(n8166) );
  AOI211_X1 U9803 ( .C1(n8236), .C2(n8768), .A(n8167), .B(n8166), .ZN(n8168)
         );
  OAI211_X1 U9804 ( .C1(n8170), .C2(n8245), .A(n8169), .B(n8168), .ZN(P2_U3168) );
  OAI22_X1 U9805 ( .A1(n8173), .A2(n8696), .B1(n8172), .B2(n8171), .ZN(n8177)
         );
  XNOR2_X1 U9806 ( .A(n8175), .B(n8174), .ZN(n8176) );
  XNOR2_X1 U9807 ( .A(n8177), .B(n8176), .ZN(n8182) );
  NOR2_X1 U9808 ( .A1(n8223), .A2(n8205), .ZN(n8179) );
  INV_X1 U9809 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10358) );
  OAI22_X1 U9810 ( .A1(n8224), .A2(n8238), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10358), .ZN(n8178) );
  AOI211_X1 U9811 ( .C1(n8673), .C2(n8241), .A(n8179), .B(n8178), .ZN(n8181)
         );
  NAND2_X1 U9812 ( .A1(n8902), .A2(n8227), .ZN(n8180) );
  OAI211_X1 U9813 ( .C1(n8182), .C2(n8230), .A(n8181), .B(n8180), .ZN(P2_U3169) );
  XOR2_X1 U9814 ( .A(n8184), .B(n8183), .Z(n8189) );
  NAND2_X1 U9815 ( .A1(n8241), .A2(n8723), .ZN(n8186) );
  AOI22_X1 U9816 ( .A1(n8211), .A2(n8717), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8185) );
  OAI211_X1 U9817 ( .C1(n8747), .C2(n8223), .A(n8186), .B(n8185), .ZN(n8187)
         );
  AOI21_X1 U9818 ( .B1(n8722), .B2(n8227), .A(n8187), .ZN(n8188) );
  OAI21_X1 U9819 ( .B1(n8189), .B2(n8230), .A(n8188), .ZN(P2_U3173) );
  INV_X1 U9820 ( .A(n8190), .ZN(n8191) );
  AOI21_X1 U9821 ( .B1(n8193), .B2(n8192), .A(n8191), .ZN(n8200) );
  NAND2_X1 U9822 ( .A1(n8241), .A2(n8194), .ZN(n8196) );
  AOI22_X1 U9823 ( .A1(n8211), .A2(n8470), .B1(P2_REG3_REG_13__SCAN_IN), .B2(
        P2_U3151), .ZN(n8195) );
  OAI211_X1 U9824 ( .C1(n8197), .C2(n8223), .A(n8196), .B(n8195), .ZN(n8198)
         );
  AOI21_X1 U9825 ( .B1(n8358), .B2(n8227), .A(n8198), .ZN(n8199) );
  OAI21_X1 U9826 ( .B1(n8200), .B2(n8230), .A(n8199), .ZN(P2_U3174) );
  XOR2_X1 U9827 ( .A(n8202), .B(n8201), .Z(n8208) );
  NAND2_X1 U9828 ( .A1(n8241), .A2(n8699), .ZN(n8204) );
  AOI22_X1 U9829 ( .A1(n8236), .A2(n8717), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8203) );
  OAI211_X1 U9830 ( .C1(n8205), .C2(n8238), .A(n8204), .B(n8203), .ZN(n8206)
         );
  AOI21_X1 U9831 ( .B1(n8914), .B2(n8227), .A(n8206), .ZN(n8207) );
  OAI21_X1 U9832 ( .B1(n8208), .B2(n8230), .A(n8207), .ZN(P2_U3175) );
  XOR2_X1 U9833 ( .A(n8210), .B(n8209), .Z(n8216) );
  NAND2_X1 U9834 ( .A1(n8241), .A2(n8754), .ZN(n8213) );
  INV_X1 U9835 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10281) );
  NOR2_X1 U9836 ( .A1(n10281), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8579) );
  AOI21_X1 U9837 ( .B1(n8211), .B2(n8718), .A(n8579), .ZN(n8212) );
  OAI211_X1 U9838 ( .C1(n8749), .C2(n8223), .A(n8213), .B(n8212), .ZN(n8214)
         );
  AOI21_X1 U9839 ( .B1(n8854), .B2(n8227), .A(n8214), .ZN(n8215) );
  OAI21_X1 U9840 ( .B1(n8216), .B2(n8230), .A(n8215), .ZN(P2_U3178) );
  INV_X1 U9841 ( .A(n8217), .ZN(n8218) );
  NOR2_X1 U9842 ( .A1(n8219), .A2(n8218), .ZN(n8220) );
  XNOR2_X1 U9843 ( .A(n8221), .B(n8220), .ZN(n8231) );
  OAI22_X1 U9844 ( .A1(n8224), .A2(n8223), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8222), .ZN(n8226) );
  NOR2_X1 U9845 ( .A1(n8624), .A2(n8238), .ZN(n8225) );
  AOI211_X1 U9846 ( .C1(n8650), .C2(n8241), .A(n8226), .B(n8225), .ZN(n8229)
         );
  NAND2_X1 U9847 ( .A1(n8890), .A2(n8227), .ZN(n8228) );
  OAI211_X1 U9848 ( .C1(n8231), .C2(n8230), .A(n8229), .B(n8228), .ZN(P2_U3180) );
  OAI211_X1 U9849 ( .C1(n8235), .C2(n8234), .A(n8233), .B(n8232), .ZN(n8244)
         );
  NAND2_X1 U9850 ( .A1(n8236), .A2(n8470), .ZN(n8237) );
  NAND2_X1 U9851 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8513) );
  OAI211_X1 U9852 ( .C1(n8239), .C2(n8238), .A(n8237), .B(n8513), .ZN(n8240)
         );
  AOI21_X1 U9853 ( .B1(n8242), .B2(n8241), .A(n8240), .ZN(n8243) );
  OAI211_X1 U9854 ( .C1(n8953), .C2(n8245), .A(n8244), .B(n8243), .ZN(P2_U3181) );
  NOR2_X1 U9855 ( .A1(n4510), .A2(n8246), .ZN(n8247) );
  INV_X1 U9856 ( .A(n8436), .ZN(n8467) );
  AND2_X1 U9857 ( .A1(n8876), .A2(n8467), .ZN(n8285) );
  AOI22_X1 U9858 ( .A1(n9626), .A2(n8250), .B1(n8249), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n8815) );
  INV_X1 U9859 ( .A(n8815), .ZN(n8869) );
  INV_X1 U9860 ( .A(n8876), .ZN(n8816) );
  NAND2_X1 U9861 ( .A1(n8816), .A2(n8436), .ZN(n8286) );
  NAND2_X1 U9862 ( .A1(n8286), .A2(n8252), .ZN(n8431) );
  NAND2_X1 U9863 ( .A1(n6483), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8257) );
  NAND2_X1 U9864 ( .A1(n4515), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8256) );
  NAND2_X1 U9865 ( .A1(n8254), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8255) );
  AND3_X1 U9866 ( .A1(n8257), .A2(n8256), .A3(n8255), .ZN(n8258) );
  NAND2_X1 U9867 ( .A1(n8259), .A2(n8258), .ZN(n8607) );
  NAND2_X1 U9868 ( .A1(n8815), .A2(n8607), .ZN(n8440) );
  OAI21_X1 U9869 ( .B1(n8876), .B2(n8869), .A(n8440), .ZN(n8260) );
  INV_X1 U9870 ( .A(n8622), .ZN(n8284) );
  INV_X1 U9871 ( .A(n8261), .ZN(n8289) );
  INV_X1 U9872 ( .A(n8655), .ZN(n8653) );
  NAND2_X1 U9873 ( .A1(n8411), .A2(n8666), .ZN(n8684) );
  INV_X1 U9874 ( .A(n8715), .ZN(n8720) );
  INV_X1 U9875 ( .A(n7173), .ZN(n8263) );
  NAND4_X1 U9876 ( .A1(n8265), .A2(n8264), .A3(n8263), .A4(n8262), .ZN(n8269)
         );
  NOR4_X1 U9877 ( .A1(n8269), .A2(n8268), .A3(n8267), .A4(n8266), .ZN(n8271)
         );
  NAND3_X1 U9878 ( .A1(n8271), .A2(n8270), .A3(n8323), .ZN(n8274) );
  NOR4_X1 U9879 ( .A1(n8275), .A2(n8274), .A3(n8273), .A4(n8272), .ZN(n8277)
         );
  NAND4_X1 U9880 ( .A1(n8364), .A2(n8352), .A3(n8277), .A4(n8276), .ZN(n8278)
         );
  NOR4_X1 U9881 ( .A1(n8761), .A2(n6598), .A3(n8279), .A4(n8278), .ZN(n8280)
         );
  NAND4_X1 U9882 ( .A1(n8720), .A2(n8745), .A3(n8736), .A4(n8280), .ZN(n8281)
         );
  NOR4_X1 U9883 ( .A1(n8684), .A2(n8695), .A3(n8706), .A4(n8281), .ZN(n8282)
         );
  NAND4_X1 U9884 ( .A1(n8643), .A2(n8653), .A3(n8669), .A4(n8282), .ZN(n8283)
         );
  NOR4_X1 U9885 ( .A1(n8429), .A2(n8284), .A3(n8633), .A4(n8283), .ZN(n8287)
         );
  INV_X1 U9886 ( .A(n8285), .ZN(n8454) );
  NAND4_X1 U9887 ( .A1(n8440), .A2(n8287), .A3(n8286), .A4(n8454), .ZN(n8445)
         );
  INV_X1 U9888 ( .A(n8633), .ZN(n8425) );
  MUX2_X1 U9889 ( .A(n8289), .B(n8288), .S(n8439), .Z(n8290) );
  INV_X1 U9890 ( .A(n8290), .ZN(n8424) );
  NAND3_X1 U9891 ( .A1(n8296), .A2(n8291), .A3(n6679), .ZN(n8292) );
  OAI21_X1 U9892 ( .B1(n8798), .B2(n8292), .A(n8303), .ZN(n8293) );
  NAND2_X1 U9893 ( .A1(n8295), .A2(n6571), .ZN(n8297) );
  NAND2_X1 U9894 ( .A1(n8297), .A2(n8296), .ZN(n8300) );
  NAND2_X1 U9895 ( .A1(n8309), .A2(n8298), .ZN(n8299) );
  AOI21_X1 U9896 ( .B1(n8262), .B2(n8300), .A(n8299), .ZN(n8301) );
  INV_X1 U9897 ( .A(n8303), .ZN(n8305) );
  OAI211_X1 U9898 ( .C1(n8313), .C2(n8305), .A(n8304), .B(n8314), .ZN(n8308)
         );
  INV_X1 U9899 ( .A(n8318), .ZN(n8306) );
  AOI21_X1 U9900 ( .B1(n8308), .B2(n8307), .A(n8306), .ZN(n8320) );
  INV_X1 U9901 ( .A(n8309), .ZN(n8312) );
  OAI211_X1 U9902 ( .C1(n8313), .C2(n8312), .A(n8311), .B(n8310), .ZN(n8315)
         );
  NAND2_X1 U9903 ( .A1(n8315), .A2(n8314), .ZN(n8317) );
  NAND2_X1 U9904 ( .A1(n8317), .A2(n8316), .ZN(n8319) );
  NOR2_X1 U9905 ( .A1(n8335), .A2(n8435), .ZN(n8321) );
  NAND2_X1 U9906 ( .A1(n8321), .A2(n8336), .ZN(n8331) );
  NAND3_X1 U9907 ( .A1(n8329), .A2(n8435), .A3(n8327), .ZN(n8322) );
  NAND2_X1 U9908 ( .A1(n8331), .A2(n8322), .ZN(n8333) );
  NAND2_X1 U9909 ( .A1(n8325), .A2(n8324), .ZN(n8326) );
  AND2_X1 U9910 ( .A1(n8327), .A2(n8326), .ZN(n8330) );
  OAI211_X1 U9911 ( .C1(n8331), .C2(n8330), .A(n8329), .B(n8328), .ZN(n8339)
         );
  INV_X1 U9912 ( .A(n8332), .ZN(n8334) );
  OAI21_X1 U9913 ( .B1(n8335), .B2(n8334), .A(n8333), .ZN(n8337) );
  NAND3_X1 U9914 ( .A1(n8337), .A2(n8336), .A3(n8344), .ZN(n8338) );
  MUX2_X1 U9915 ( .A(n8339), .B(n8338), .S(n8435), .Z(n8340) );
  INV_X1 U9916 ( .A(n8340), .ZN(n8341) );
  INV_X1 U9917 ( .A(n8345), .ZN(n8342) );
  AOI21_X1 U9918 ( .B1(n8349), .B2(n8343), .A(n8342), .ZN(n8351) );
  AND2_X1 U9919 ( .A1(n8345), .A2(n8344), .ZN(n8348) );
  INV_X1 U9920 ( .A(n8346), .ZN(n8347) );
  AOI21_X1 U9921 ( .B1(n8349), .B2(n8348), .A(n8347), .ZN(n8350) );
  MUX2_X1 U9922 ( .A(n8351), .B(n8350), .S(n8439), .Z(n8353) );
  NAND2_X1 U9923 ( .A1(n8353), .A2(n8352), .ZN(n8357) );
  MUX2_X1 U9924 ( .A(n8355), .B(n8354), .S(n8439), .Z(n8356) );
  NAND2_X1 U9925 ( .A1(n8357), .A2(n8356), .ZN(n8361) );
  NAND2_X1 U9926 ( .A1(n8361), .A2(n4598), .ZN(n8360) );
  MUX2_X1 U9927 ( .A(n8471), .B(n8358), .S(n8439), .Z(n8359) );
  NAND2_X1 U9928 ( .A1(n8360), .A2(n8359), .ZN(n8366) );
  INV_X1 U9929 ( .A(n8361), .ZN(n8363) );
  NAND2_X1 U9930 ( .A1(n8363), .A2(n8362), .ZN(n8365) );
  NAND3_X1 U9931 ( .A1(n8366), .A2(n8365), .A3(n8364), .ZN(n8370) );
  MUX2_X1 U9932 ( .A(n8368), .B(n8367), .S(n8435), .Z(n8369) );
  NAND2_X1 U9933 ( .A1(n8370), .A2(n8369), .ZN(n8371) );
  NAND2_X1 U9934 ( .A1(n8371), .A2(n4512), .ZN(n8388) );
  NAND3_X1 U9935 ( .A1(n8388), .A2(n8784), .A3(n8372), .ZN(n8375) );
  XNOR2_X1 U9936 ( .A(n8373), .B(n8439), .ZN(n8374) );
  NAND2_X1 U9937 ( .A1(n8375), .A2(n8374), .ZN(n8378) );
  INV_X1 U9938 ( .A(n8761), .ZN(n8764) );
  AOI21_X1 U9939 ( .B1(n8392), .B2(n8376), .A(n8435), .ZN(n8377) );
  AOI21_X1 U9940 ( .B1(n8378), .B2(n8764), .A(n8377), .ZN(n8391) );
  INV_X1 U9941 ( .A(n8391), .ZN(n8380) );
  NAND2_X1 U9942 ( .A1(n8380), .A2(n8379), .ZN(n8381) );
  NAND3_X1 U9943 ( .A1(n8381), .A2(n8397), .A3(n8393), .ZN(n8385) );
  AND2_X1 U9944 ( .A1(n8399), .A2(n8382), .ZN(n8384) );
  INV_X1 U9945 ( .A(n8398), .ZN(n8383) );
  AOI21_X1 U9946 ( .B1(n8385), .B2(n8384), .A(n8383), .ZN(n8404) );
  AOI21_X1 U9947 ( .B1(n8388), .B2(n8387), .A(n4886), .ZN(n8390) );
  OAI211_X1 U9948 ( .C1(n8391), .C2(n8390), .A(n8389), .B(n8735), .ZN(n8394)
         );
  NAND3_X1 U9949 ( .A1(n8394), .A2(n8393), .A3(n8392), .ZN(n8396) );
  NAND3_X1 U9950 ( .A1(n8396), .A2(n8720), .A3(n8395), .ZN(n8402) );
  AND2_X1 U9951 ( .A1(n8398), .A2(n8397), .ZN(n8401) );
  INV_X1 U9952 ( .A(n8399), .ZN(n8400) );
  AOI21_X1 U9953 ( .B1(n8402), .B2(n8401), .A(n8400), .ZN(n8403) );
  MUX2_X1 U9954 ( .A(n8404), .B(n8403), .S(n8435), .Z(n8410) );
  INV_X1 U9955 ( .A(n8695), .ZN(n8692) );
  NAND2_X1 U9956 ( .A1(n8411), .A2(n8405), .ZN(n8408) );
  NAND2_X1 U9957 ( .A1(n8666), .A2(n8406), .ZN(n8407) );
  MUX2_X1 U9958 ( .A(n8408), .B(n8407), .S(n8435), .Z(n8409) );
  AOI21_X1 U9959 ( .B1(n8410), .B2(n8692), .A(n8409), .ZN(n8419) );
  NAND2_X1 U9960 ( .A1(n8415), .A2(n8411), .ZN(n8414) );
  INV_X1 U9961 ( .A(n8412), .ZN(n8413) );
  MUX2_X1 U9962 ( .A(n8414), .B(n8413), .S(n8439), .Z(n8418) );
  MUX2_X1 U9963 ( .A(n8416), .B(n8415), .S(n8439), .Z(n8417) );
  OAI211_X1 U9964 ( .C1(n8419), .C2(n8418), .A(n8653), .B(n8417), .ZN(n8423)
         );
  MUX2_X1 U9965 ( .A(n8421), .B(n8420), .S(n8435), .Z(n8422) );
  NAND2_X1 U9966 ( .A1(n8884), .A2(n8624), .ZN(n8427) );
  MUX2_X1 U9967 ( .A(n8427), .B(n8426), .S(n8435), .Z(n8428) );
  AOI21_X1 U9968 ( .B1(n4722), .B2(n8430), .A(n8453), .ZN(n8456) );
  INV_X1 U9969 ( .A(n8431), .ZN(n8434) );
  AOI21_X1 U9970 ( .B1(n8453), .B2(n8879), .A(n8432), .ZN(n8433) );
  OAI211_X1 U9971 ( .C1(n8456), .C2(n8468), .A(n8434), .B(n8433), .ZN(n8443)
         );
  OAI21_X1 U9972 ( .B1(n8436), .B2(n8435), .A(n8816), .ZN(n8438) );
  OAI211_X1 U9973 ( .C1(n8439), .C2(n8467), .A(n8438), .B(n8437), .ZN(n8442)
         );
  INV_X1 U9974 ( .A(n8440), .ZN(n8441) );
  AOI21_X1 U9975 ( .B1(n8443), .B2(n8442), .A(n8441), .ZN(n8444) );
  INV_X1 U9976 ( .A(n8449), .ZN(n8450) );
  NAND3_X1 U9977 ( .A1(n8451), .A2(n8450), .A3(n8463), .ZN(n8452) );
  AOI21_X1 U9978 ( .B1(n8453), .B2(n8468), .A(n8452), .ZN(n8455) );
  OAI211_X1 U9979 ( .C1(n8456), .C2(n8879), .A(n8455), .B(n8454), .ZN(n8458)
         );
  INV_X1 U9980 ( .A(n8607), .ZN(n8457) );
  NAND3_X1 U9981 ( .A1(n8461), .A2(n8460), .A3(n8540), .ZN(n8462) );
  OAI211_X1 U9982 ( .C1(n8463), .C2(n8465), .A(n8462), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8464) );
  OAI21_X1 U9983 ( .B1(n8466), .B2(n8465), .A(n8464), .ZN(P2_U3296) );
  MUX2_X1 U9984 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8607), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9985 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8467), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9986 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8468), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9987 ( .A(n8647), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8573), .Z(
        P2_U3518) );
  MUX2_X1 U9988 ( .A(n8657), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8573), .Z(
        P2_U3517) );
  MUX2_X1 U9989 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8671), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9990 ( .A(n8685), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8573), .Z(
        P2_U3515) );
  MUX2_X1 U9991 ( .A(n8696), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8573), .Z(
        P2_U3514) );
  MUX2_X1 U9992 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8686), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9993 ( .A(n8717), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8573), .Z(
        P2_U3512) );
  MUX2_X1 U9994 ( .A(n8732), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8573), .Z(
        P2_U3511) );
  MUX2_X1 U9995 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8718), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9996 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8767), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9997 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8787), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9998 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8768), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9999 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8469), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10000 ( .A(n8470), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8573), .Z(
        P2_U3505) );
  MUX2_X1 U10001 ( .A(n8471), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8573), .Z(
        P2_U3504) );
  MUX2_X1 U10002 ( .A(n8472), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8573), .Z(
        P2_U3503) );
  MUX2_X1 U10003 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8473), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10004 ( .A(n8474), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8573), .Z(
        P2_U3501) );
  MUX2_X1 U10005 ( .A(n8475), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8573), .Z(
        P2_U3500) );
  MUX2_X1 U10006 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8476), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U10007 ( .A(n8477), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8573), .Z(
        P2_U3498) );
  MUX2_X1 U10008 ( .A(n8478), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8573), .Z(
        P2_U3497) );
  MUX2_X1 U10009 ( .A(n8479), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8573), .Z(
        P2_U3496) );
  MUX2_X1 U10010 ( .A(n8480), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8573), .Z(
        P2_U3495) );
  MUX2_X1 U10011 ( .A(n8799), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8573), .Z(
        P2_U3494) );
  MUX2_X1 U10012 ( .A(n8481), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8573), .Z(
        P2_U3493) );
  MUX2_X1 U10013 ( .A(n6572), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8573), .Z(
        P2_U3492) );
  MUX2_X1 U10014 ( .A(n8482), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8573), .Z(
        P2_U3491) );
  INV_X1 U10015 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8505) );
  NOR2_X1 U10016 ( .A1(n9938), .A2(n8485), .ZN(n8486) );
  AOI22_X1 U10017 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8502), .B1(n9971), .B2(
        n8500), .ZN(n9964) );
  AOI21_X1 U10018 ( .B1(n8505), .B2(n8487), .A(n8523), .ZN(n8520) );
  AOI22_X1 U10019 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n9971), .B1(n8502), .B2(
        n8499), .ZN(n9956) );
  OAI21_X1 U10020 ( .B1(n8490), .B2(n8489), .A(n8488), .ZN(n8491) );
  NAND2_X1 U10021 ( .A1(n8496), .A2(n8491), .ZN(n8492) );
  NAND2_X1 U10022 ( .A1(n8492), .A2(n9939), .ZN(n9955) );
  NAND2_X1 U10023 ( .A1(n9956), .A2(n9955), .ZN(n9954) );
  OAI21_X1 U10024 ( .B1(n8502), .B2(n8499), .A(n9954), .ZN(n8531) );
  OAI21_X1 U10025 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n8493), .A(n8533), .ZN(
        n8518) );
  NAND2_X1 U10026 ( .A1(n9944), .A2(n9943), .ZN(n8498) );
  MUX2_X1 U10027 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8540), .Z(n8495) );
  INV_X1 U10028 ( .A(n8495), .ZN(n8494) );
  NAND2_X1 U10029 ( .A1(n8494), .A2(n9938), .ZN(n9959) );
  NAND2_X1 U10030 ( .A1(n8496), .A2(n8495), .ZN(n8497) );
  AND2_X1 U10031 ( .A1(n9959), .A2(n8497), .ZN(n9941) );
  NAND2_X1 U10032 ( .A1(n8498), .A2(n9941), .ZN(n9960) );
  NAND2_X1 U10033 ( .A1(n9960), .A2(n9959), .ZN(n8504) );
  MUX2_X1 U10034 ( .A(n8500), .B(n8499), .S(n8540), .Z(n8501) );
  NAND2_X1 U10035 ( .A1(n8502), .A2(n8501), .ZN(n8511) );
  OR2_X1 U10036 ( .A1(n8502), .A2(n8501), .ZN(n8503) );
  AND2_X1 U10037 ( .A1(n8511), .A2(n8503), .ZN(n9957) );
  NAND2_X1 U10038 ( .A1(n8504), .A2(n9957), .ZN(n9962) );
  NAND2_X1 U10039 ( .A1(n9962), .A2(n8511), .ZN(n8508) );
  INV_X1 U10040 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8865) );
  MUX2_X1 U10041 ( .A(n8505), .B(n8865), .S(n8540), .Z(n8506) );
  NAND2_X1 U10042 ( .A1(n8522), .A2(n8506), .ZN(n9979) );
  OR2_X1 U10043 ( .A1(n8522), .A2(n8506), .ZN(n8507) );
  AND2_X1 U10044 ( .A1(n9979), .A2(n8507), .ZN(n8509) );
  NAND2_X1 U10045 ( .A1(n8508), .A2(n8509), .ZN(n9980) );
  INV_X1 U10046 ( .A(n8509), .ZN(n8510) );
  NAND3_X1 U10047 ( .A1(n9962), .A2(n8511), .A3(n8510), .ZN(n8512) );
  AOI21_X1 U10048 ( .B1(n9980), .B2(n8512), .A(n9981), .ZN(n8517) );
  INV_X1 U10049 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10291) );
  NAND2_X1 U10050 ( .A1(n9937), .A2(n8522), .ZN(n8514) );
  OAI211_X1 U10051 ( .C1(n10291), .C2(n8515), .A(n8514), .B(n8513), .ZN(n8516)
         );
  AOI211_X1 U10052 ( .C1(n8518), .C2(n9991), .A(n8517), .B(n8516), .ZN(n8519)
         );
  OAI21_X1 U10053 ( .B1(n8520), .B2(n9986), .A(n8519), .ZN(P2_U3197) );
  NOR2_X1 U10054 ( .A1(n8522), .A2(n8521), .ZN(n8524) );
  NAND2_X1 U10055 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n9994), .ZN(n8525) );
  OAI21_X1 U10056 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n9994), .A(n8525), .ZN(
        n9985) );
  INV_X1 U10057 ( .A(n8526), .ZN(n8527) );
  OAI21_X1 U10058 ( .B1(n8527), .B2(n8554), .A(n8561), .ZN(n8530) );
  INV_X1 U10059 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8772) );
  AOI21_X1 U10060 ( .B1(n8530), .B2(n8772), .A(n8529), .ZN(n8552) );
  INV_X1 U10061 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n10226) );
  AOI22_X1 U10062 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n9994), .B1(n8537), .B2(
        n10226), .ZN(n9976) );
  NAND2_X1 U10063 ( .A1(n8532), .A2(n8531), .ZN(n8534) );
  NAND2_X1 U10064 ( .A1(n8534), .A2(n8533), .ZN(n9975) );
  NAND2_X1 U10065 ( .A1(n9976), .A2(n9975), .ZN(n9974) );
  XNOR2_X1 U10066 ( .A(n8553), .B(n8566), .ZN(n8535) );
  NAND2_X1 U10067 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n8535), .ZN(n8555) );
  OAI21_X1 U10068 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8535), .A(n8555), .ZN(
        n8550) );
  NAND2_X1 U10069 ( .A1(n9980), .A2(n9979), .ZN(n8539) );
  INV_X1 U10070 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8788) );
  MUX2_X1 U10071 ( .A(n8788), .B(n10226), .S(n8540), .Z(n8536) );
  OR2_X1 U10072 ( .A1(n8537), .A2(n8536), .ZN(n8538) );
  NAND2_X1 U10073 ( .A1(n8537), .A2(n8536), .ZN(n8543) );
  AND2_X1 U10074 ( .A1(n8538), .A2(n8543), .ZN(n9977) );
  NAND2_X1 U10075 ( .A1(n8539), .A2(n9977), .ZN(n9983) );
  NAND2_X1 U10076 ( .A1(n9983), .A2(n8543), .ZN(n8541) );
  MUX2_X1 U10077 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8540), .Z(n8564) );
  XNOR2_X1 U10078 ( .A(n8566), .B(n8564), .ZN(n8542) );
  NAND2_X1 U10079 ( .A1(n8541), .A2(n8542), .ZN(n8568) );
  INV_X1 U10080 ( .A(n8542), .ZN(n8544) );
  NAND3_X1 U10081 ( .A1(n9983), .A2(n8544), .A3(n8543), .ZN(n8545) );
  AOI21_X1 U10082 ( .B1(n8568), .B2(n8545), .A(n9981), .ZN(n8549) );
  NOR2_X1 U10083 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10348), .ZN(n8546) );
  AOI21_X1 U10084 ( .B1(n9973), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8546), .ZN(
        n8547) );
  OAI21_X1 U10085 ( .B1(n9995), .B2(n8554), .A(n8547), .ZN(n8548) );
  AOI211_X1 U10086 ( .C1(n8550), .C2(n9991), .A(n8549), .B(n8548), .ZN(n8551)
         );
  OAI21_X1 U10087 ( .B1(n8552), .B2(n9986), .A(n8551), .ZN(P2_U3199) );
  XNOR2_X1 U10088 ( .A(n8557), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8585) );
  NAND2_X1 U10089 ( .A1(n8554), .A2(n8553), .ZN(n8556) );
  NAND2_X1 U10090 ( .A1(n8556), .A2(n8555), .ZN(n8586) );
  INV_X1 U10091 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8569) );
  OR2_X1 U10092 ( .A1(n8557), .A2(n8569), .ZN(n8583) );
  NAND2_X1 U10093 ( .A1(n8557), .A2(n8569), .ZN(n8558) );
  NAND2_X1 U10094 ( .A1(n8583), .A2(n8558), .ZN(n8559) );
  AND3_X1 U10095 ( .A1(n8561), .A2(n8560), .A3(n8559), .ZN(n8563) );
  OAI21_X1 U10096 ( .B1(n8584), .B2(n8563), .A(n8562), .ZN(n8581) );
  INV_X1 U10097 ( .A(n8564), .ZN(n8565) );
  NAND2_X1 U10098 ( .A1(n8566), .A2(n8565), .ZN(n8567) );
  NAND2_X1 U10099 ( .A1(n8568), .A2(n8567), .ZN(n8571) );
  INV_X1 U10100 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8855) );
  MUX2_X1 U10101 ( .A(n8569), .B(n8855), .S(n8540), .Z(n8570) );
  NOR2_X1 U10102 ( .A1(n8571), .A2(n8570), .ZN(n8588) );
  NAND2_X1 U10103 ( .A1(n8571), .A2(n8570), .ZN(n8589) );
  INV_X1 U10104 ( .A(n8589), .ZN(n8572) );
  OR2_X1 U10105 ( .A1(n8588), .A2(n8572), .ZN(n8574) );
  OAI21_X1 U10106 ( .B1(n8574), .B2(n8573), .A(n9995), .ZN(n8577) );
  INV_X1 U10107 ( .A(n8574), .ZN(n8575) );
  NOR2_X1 U10108 ( .A1(n8575), .A2(n9981), .ZN(n8576) );
  MUX2_X1 U10109 ( .A(n8577), .B(n8576), .S(n8590), .Z(n8578) );
  AOI211_X1 U10110 ( .C1(n9973), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8579), .B(
        n8578), .ZN(n8580) );
  XNOR2_X1 U10111 ( .A(n8599), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8592) );
  AOI22_X1 U10112 ( .A1(n8586), .A2(n8585), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8590), .ZN(n8587) );
  XNOR2_X1 U10113 ( .A(n8599), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8593) );
  XNOR2_X1 U10114 ( .A(n8587), .B(n8593), .ZN(n8602) );
  AOI21_X1 U10115 ( .B1(n8590), .B2(n8589), .A(n8588), .ZN(n8595) );
  MUX2_X1 U10116 ( .A(n8593), .B(n8592), .S(n8591), .Z(n8594) );
  XNOR2_X1 U10117 ( .A(n8595), .B(n8594), .ZN(n8596) );
  NOR2_X1 U10118 ( .A1(n8596), .A2(n9981), .ZN(n8601) );
  NAND2_X1 U10119 ( .A1(n9973), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8597) );
  OAI211_X1 U10120 ( .C1(n9995), .C2(n8599), .A(n8598), .B(n8597), .ZN(n8600)
         );
  OAI21_X1 U10121 ( .B1(n8604), .B2(n9986), .A(n8603), .ZN(P2_U3201) );
  INV_X1 U10122 ( .A(n8605), .ZN(n8606) );
  NAND2_X1 U10123 ( .A1(n8607), .A2(n8606), .ZN(n8870) );
  OAI22_X1 U10124 ( .A1(n8771), .A2(n8870), .B1(n8614), .B2(n8674), .ZN(n8609)
         );
  AOI21_X1 U10125 ( .B1(n8771), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8609), .ZN(
        n8608) );
  OAI21_X1 U10126 ( .B1(n8815), .B2(n8725), .A(n8608), .ZN(P2_U3202) );
  AOI21_X1 U10127 ( .B1(n8771), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8609), .ZN(
        n8610) );
  OAI21_X1 U10128 ( .B1(n8876), .B2(n8725), .A(n8610), .ZN(P2_U3203) );
  INV_X1 U10129 ( .A(n8611), .ZN(n8620) );
  NAND2_X1 U10130 ( .A1(n8612), .A2(n8812), .ZN(n8618) );
  INV_X1 U10131 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8613) );
  OAI22_X1 U10132 ( .A1(n8614), .A2(n8674), .B1(n8613), .B2(n8812), .ZN(n8615)
         );
  AOI21_X1 U10133 ( .B1(n8616), .B2(n4507), .A(n8615), .ZN(n8617) );
  OAI211_X1 U10134 ( .C1(n8620), .C2(n8619), .A(n8618), .B(n8617), .ZN(
        P2_U3204) );
  XNOR2_X1 U10135 ( .A(n8621), .B(n8622), .ZN(n8882) );
  XNOR2_X1 U10136 ( .A(n8623), .B(n8622), .ZN(n8627) );
  OAI22_X1 U10137 ( .A1(n8625), .A2(n8748), .B1(n8624), .B2(n8779), .ZN(n8626)
         );
  AOI21_X1 U10138 ( .B1(n8627), .B2(n8805), .A(n8626), .ZN(n8877) );
  MUX2_X1 U10139 ( .A(n8628), .B(n8877), .S(n8812), .Z(n8631) );
  AOI22_X1 U10140 ( .A1(n8879), .A2(n4507), .B1(n8808), .B2(n8629), .ZN(n8630)
         );
  OAI211_X1 U10141 ( .C1(n8882), .C2(n8793), .A(n8631), .B(n8630), .ZN(
        P2_U3205) );
  XNOR2_X1 U10142 ( .A(n8632), .B(n8633), .ZN(n8887) );
  INV_X1 U10143 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8639) );
  XNOR2_X1 U10144 ( .A(n8634), .B(n8633), .ZN(n8638) );
  OAI22_X1 U10145 ( .A1(n8636), .A2(n8748), .B1(n8635), .B2(n8779), .ZN(n8637)
         );
  AOI21_X1 U10146 ( .B1(n8638), .B2(n8805), .A(n8637), .ZN(n8883) );
  MUX2_X1 U10147 ( .A(n8639), .B(n8883), .S(n8812), .Z(n8642) );
  AOI22_X1 U10148 ( .A1(n8884), .A2(n4507), .B1(n8808), .B2(n8640), .ZN(n8641)
         );
  OAI211_X1 U10149 ( .C1(n8887), .C2(n8793), .A(n8642), .B(n8641), .ZN(
        P2_U3206) );
  XNOR2_X1 U10150 ( .A(n8644), .B(n8643), .ZN(n8893) );
  XNOR2_X1 U10151 ( .A(n8645), .B(n8646), .ZN(n8648) );
  AOI222_X1 U10152 ( .A1(n8805), .A2(n8648), .B1(n8647), .B2(n8800), .C1(n8671), .C2(n8801), .ZN(n8888) );
  MUX2_X1 U10153 ( .A(n8649), .B(n8888), .S(n8812), .Z(n8652) );
  AOI22_X1 U10154 ( .A1(n8890), .A2(n4507), .B1(n8808), .B2(n8650), .ZN(n8651)
         );
  OAI211_X1 U10155 ( .C1(n8893), .C2(n8793), .A(n8652), .B(n8651), .ZN(
        P2_U3207) );
  XNOR2_X1 U10156 ( .A(n8654), .B(n8653), .ZN(n8899) );
  XNOR2_X1 U10157 ( .A(n8656), .B(n8655), .ZN(n8658) );
  AOI222_X1 U10158 ( .A1(n8805), .A2(n8658), .B1(n8657), .B2(n8800), .C1(n8685), .C2(n8801), .ZN(n8894) );
  INV_X1 U10159 ( .A(n8894), .ZN(n8663) );
  INV_X1 U10160 ( .A(n8896), .ZN(n8661) );
  INV_X1 U10161 ( .A(n8659), .ZN(n8660) );
  OAI22_X1 U10162 ( .A1(n8661), .A2(n8676), .B1(n8660), .B2(n8674), .ZN(n8662)
         );
  OAI21_X1 U10163 ( .B1(n8663), .B2(n8662), .A(n8812), .ZN(n8665) );
  NAND2_X1 U10164 ( .A1(n8771), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8664) );
  OAI211_X1 U10165 ( .C1(n8899), .C2(n8793), .A(n8665), .B(n8664), .ZN(
        P2_U3208) );
  NAND2_X1 U10166 ( .A1(n8667), .A2(n8666), .ZN(n8668) );
  XOR2_X1 U10167 ( .A(n8669), .B(n8668), .Z(n8905) );
  XNOR2_X1 U10168 ( .A(n8670), .B(n8669), .ZN(n8672) );
  AOI222_X1 U10169 ( .A1(n8805), .A2(n8672), .B1(n8696), .B2(n8801), .C1(n8671), .C2(n8800), .ZN(n8900) );
  INV_X1 U10170 ( .A(n8900), .ZN(n8679) );
  INV_X1 U10171 ( .A(n8902), .ZN(n8677) );
  INV_X1 U10172 ( .A(n8673), .ZN(n8675) );
  OAI22_X1 U10173 ( .A1(n8677), .A2(n8676), .B1(n8675), .B2(n8674), .ZN(n8678)
         );
  OAI21_X1 U10174 ( .B1(n8679), .B2(n8678), .A(n8812), .ZN(n8681) );
  NAND2_X1 U10175 ( .A1(n8771), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8680) );
  OAI211_X1 U10176 ( .C1(n8905), .C2(n8793), .A(n8681), .B(n8680), .ZN(
        P2_U3209) );
  XNOR2_X1 U10177 ( .A(n8682), .B(n8684), .ZN(n8911) );
  XNOR2_X1 U10178 ( .A(n8683), .B(n8684), .ZN(n8687) );
  AOI222_X1 U10179 ( .A1(n8805), .A2(n8687), .B1(n8686), .B2(n8801), .C1(n8685), .C2(n8800), .ZN(n8906) );
  MUX2_X1 U10180 ( .A(n8688), .B(n8906), .S(n8812), .Z(n8691) );
  AOI22_X1 U10181 ( .A1(n8908), .A2(n4507), .B1(n8808), .B2(n8689), .ZN(n8690)
         );
  OAI211_X1 U10182 ( .C1(n8911), .C2(n8793), .A(n8691), .B(n8690), .ZN(
        P2_U3210) );
  XNOR2_X1 U10183 ( .A(n8693), .B(n8692), .ZN(n8917) );
  XNOR2_X1 U10184 ( .A(n8694), .B(n8695), .ZN(n8697) );
  AOI222_X1 U10185 ( .A1(n8805), .A2(n8697), .B1(n8717), .B2(n8801), .C1(n8696), .C2(n8800), .ZN(n8912) );
  MUX2_X1 U10186 ( .A(n8698), .B(n8912), .S(n8812), .Z(n8701) );
  AOI22_X1 U10187 ( .A1(n8914), .A2(n4507), .B1(n8808), .B2(n8699), .ZN(n8700)
         );
  OAI211_X1 U10188 ( .C1(n8917), .C2(n8793), .A(n8701), .B(n8700), .ZN(
        P2_U3211) );
  XOR2_X1 U10189 ( .A(n8702), .B(n8706), .Z(n8703) );
  OAI222_X1 U10190 ( .A1(n8779), .A2(n8705), .B1(n8748), .B2(n8704), .C1(n8782), .C2(n8703), .ZN(n8841) );
  INV_X1 U10191 ( .A(n8841), .ZN(n8713) );
  XNOR2_X1 U10192 ( .A(n8707), .B(n8706), .ZN(n8842) );
  INV_X1 U10193 ( .A(n8708), .ZN(n8921) );
  AOI22_X1 U10194 ( .A1(n8771), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8808), .B2(
        n8709), .ZN(n8710) );
  OAI21_X1 U10195 ( .B1(n8921), .B2(n8725), .A(n8710), .ZN(n8711) );
  AOI21_X1 U10196 ( .B1(n8842), .B2(n8727), .A(n8711), .ZN(n8712) );
  OAI21_X1 U10197 ( .B1(n8713), .B2(n8771), .A(n8712), .ZN(P2_U3212) );
  OAI21_X1 U10198 ( .B1(n8716), .B2(n8715), .A(n8714), .ZN(n8719) );
  AOI222_X1 U10199 ( .A1(n8805), .A2(n8719), .B1(n8718), .B2(n8801), .C1(n8717), .C2(n8800), .ZN(n8845) );
  XNOR2_X1 U10200 ( .A(n8721), .B(n8720), .ZN(n8847) );
  INV_X1 U10201 ( .A(n8722), .ZN(n8925) );
  AOI22_X1 U10202 ( .A1(n8771), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8808), .B2(
        n8723), .ZN(n8724) );
  OAI21_X1 U10203 ( .B1(n8925), .B2(n8725), .A(n8724), .ZN(n8726) );
  AOI21_X1 U10204 ( .B1(n8847), .B2(n8727), .A(n8726), .ZN(n8728) );
  OAI21_X1 U10205 ( .B1(n8845), .B2(n8771), .A(n8728), .ZN(P2_U3213) );
  NAND2_X1 U10206 ( .A1(n8729), .A2(n8736), .ZN(n8730) );
  NAND3_X1 U10207 ( .A1(n8731), .A2(n8805), .A3(n8730), .ZN(n8734) );
  AOI22_X1 U10208 ( .A1(n8732), .A2(n8800), .B1(n8801), .B2(n8767), .ZN(n8733)
         );
  NAND2_X1 U10209 ( .A1(n8734), .A2(n8733), .ZN(n8926) );
  MUX2_X1 U10210 ( .A(n8926), .B(P2_REG2_REG_19__SCAN_IN), .S(n8771), .Z(n8741) );
  NAND2_X1 U10211 ( .A1(n8753), .A2(n8735), .ZN(n8737) );
  XNOR2_X1 U10212 ( .A(n8737), .B(n8736), .ZN(n8928) );
  AOI22_X1 U10213 ( .A1(n8850), .A2(n4507), .B1(n8808), .B2(n8738), .ZN(n8739)
         );
  OAI21_X1 U10214 ( .B1(n8928), .B2(n8793), .A(n8739), .ZN(n8740) );
  INV_X1 U10215 ( .A(n8742), .ZN(n8743) );
  AOI21_X1 U10216 ( .B1(n8745), .B2(n8744), .A(n8743), .ZN(n8746) );
  OAI222_X1 U10217 ( .A1(n8779), .A2(n8749), .B1(n8748), .B2(n8747), .C1(n8782), .C2(n8746), .ZN(n8853) );
  NAND2_X1 U10218 ( .A1(n8751), .A2(n8750), .ZN(n8752) );
  NAND2_X1 U10219 ( .A1(n8753), .A2(n8752), .ZN(n8934) );
  AOI22_X1 U10220 ( .A1(n8771), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8808), .B2(
        n8754), .ZN(n8756) );
  NAND2_X1 U10221 ( .A1(n8854), .A2(n4507), .ZN(n8755) );
  OAI211_X1 U10222 ( .C1(n8934), .C2(n8793), .A(n8756), .B(n8755), .ZN(n8757)
         );
  AOI21_X1 U10223 ( .B1(n8853), .B2(n8812), .A(n8757), .ZN(n8758) );
  INV_X1 U10224 ( .A(n8758), .ZN(P2_U3215) );
  INV_X1 U10225 ( .A(n8759), .ZN(n8760) );
  AOI21_X1 U10226 ( .B1(n8762), .B2(n8761), .A(n8760), .ZN(n8940) );
  NAND3_X1 U10227 ( .A1(n8780), .A2(n8764), .A3(n8763), .ZN(n8765) );
  NAND3_X1 U10228 ( .A1(n8766), .A2(n8805), .A3(n8765), .ZN(n8770) );
  AOI22_X1 U10229 ( .A1(n8801), .A2(n8768), .B1(n8800), .B2(n8767), .ZN(n8769)
         );
  MUX2_X1 U10230 ( .A(n8936), .B(n8772), .S(n8771), .Z(n8776) );
  INV_X1 U10231 ( .A(n8773), .ZN(n8774) );
  AOI22_X1 U10232 ( .A1(n8937), .A2(n4507), .B1(n8774), .B2(n8808), .ZN(n8775)
         );
  OAI211_X1 U10233 ( .C1(n8940), .C2(n8793), .A(n8776), .B(n8775), .ZN(
        P2_U3216) );
  XNOR2_X1 U10234 ( .A(n8777), .B(n6598), .ZN(n8948) );
  NOR2_X1 U10235 ( .A1(n8779), .A2(n8778), .ZN(n8786) );
  INV_X1 U10236 ( .A(n8780), .ZN(n8781) );
  AOI211_X1 U10237 ( .C1(n8784), .C2(n8783), .A(n8782), .B(n8781), .ZN(n8785)
         );
  AOI211_X1 U10238 ( .C1(n8800), .C2(n8787), .A(n8786), .B(n8785), .ZN(n8941)
         );
  MUX2_X1 U10239 ( .A(n8788), .B(n8941), .S(n8812), .Z(n8792) );
  AOI22_X1 U10240 ( .A1(n8944), .A2(n4507), .B1(n8808), .B2(n8789), .ZN(n8791)
         );
  OAI211_X1 U10241 ( .C1(n8948), .C2(n8793), .A(n8792), .B(n8791), .ZN(
        P2_U3217) );
  OAI21_X1 U10242 ( .B1(n8262), .B2(n8795), .A(n8794), .ZN(n9998) );
  INV_X1 U10243 ( .A(n9998), .ZN(n8811) );
  INV_X1 U10244 ( .A(n8796), .ZN(n8810) );
  XNOR2_X1 U10245 ( .A(n8797), .B(n8798), .ZN(n8806) );
  AOI22_X1 U10246 ( .A1(n8801), .A2(n6572), .B1(n8800), .B2(n8799), .ZN(n8802)
         );
  OAI21_X1 U10247 ( .B1(n8811), .B2(n8803), .A(n8802), .ZN(n8804) );
  AOI21_X1 U10248 ( .B1(n8806), .B2(n8805), .A(n8804), .ZN(n10000) );
  AOI22_X1 U10249 ( .A1(n8808), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n8807), .B2(
        n9996), .ZN(n8809) );
  OAI211_X1 U10250 ( .C1(n8811), .C2(n8810), .A(n10000), .B(n8809), .ZN(n8813)
         );
  MUX2_X1 U10251 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n8813), .S(n8812), .Z(
        P2_U3231) );
  NOR2_X1 U10252 ( .A1(n8870), .A2(n10463), .ZN(n8817) );
  AOI21_X1 U10253 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10463), .A(n8817), .ZN(
        n8814) );
  OAI21_X1 U10254 ( .B1(n8815), .B2(n8867), .A(n8814), .ZN(P2_U3490) );
  INV_X1 U10255 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8820) );
  NAND2_X1 U10256 ( .A1(n8816), .A2(n8859), .ZN(n8819) );
  INV_X1 U10257 ( .A(n8817), .ZN(n8818) );
  OAI211_X1 U10258 ( .C1(n10466), .C2(n8820), .A(n8819), .B(n8818), .ZN(
        P2_U3489) );
  INV_X1 U10259 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8821) );
  MUX2_X1 U10260 ( .A(n8821), .B(n8877), .S(n10466), .Z(n8823) );
  NAND2_X1 U10261 ( .A1(n8879), .A2(n8859), .ZN(n8822) );
  OAI211_X1 U10262 ( .C1(n8882), .C2(n8862), .A(n8823), .B(n8822), .ZN(
        P2_U3487) );
  INV_X1 U10263 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8824) );
  MUX2_X1 U10264 ( .A(n8824), .B(n8883), .S(n10466), .Z(n8826) );
  NAND2_X1 U10265 ( .A1(n8884), .A2(n8859), .ZN(n8825) );
  OAI211_X1 U10266 ( .C1(n8887), .C2(n8862), .A(n8826), .B(n8825), .ZN(
        P2_U3486) );
  INV_X1 U10267 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8827) );
  MUX2_X1 U10268 ( .A(n8827), .B(n8888), .S(n10466), .Z(n8829) );
  NAND2_X1 U10269 ( .A1(n8890), .A2(n8859), .ZN(n8828) );
  OAI211_X1 U10270 ( .C1(n8893), .C2(n8862), .A(n8829), .B(n8828), .ZN(
        P2_U3485) );
  MUX2_X1 U10271 ( .A(n10293), .B(n8894), .S(n10466), .Z(n8831) );
  NAND2_X1 U10272 ( .A1(n8896), .A2(n8859), .ZN(n8830) );
  OAI211_X1 U10273 ( .C1(n8899), .C2(n8862), .A(n8831), .B(n8830), .ZN(
        P2_U3484) );
  INV_X1 U10274 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8832) );
  MUX2_X1 U10275 ( .A(n8832), .B(n8900), .S(n10466), .Z(n8834) );
  NAND2_X1 U10276 ( .A1(n8902), .A2(n8859), .ZN(n8833) );
  OAI211_X1 U10277 ( .C1(n8862), .C2(n8905), .A(n8834), .B(n8833), .ZN(
        P2_U3483) );
  INV_X1 U10278 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8835) );
  MUX2_X1 U10279 ( .A(n8835), .B(n8906), .S(n10466), .Z(n8837) );
  NAND2_X1 U10280 ( .A1(n8908), .A2(n8859), .ZN(n8836) );
  OAI211_X1 U10281 ( .C1(n8862), .C2(n8911), .A(n8837), .B(n8836), .ZN(
        P2_U3482) );
  INV_X1 U10282 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8838) );
  MUX2_X1 U10283 ( .A(n8838), .B(n8912), .S(n10466), .Z(n8840) );
  NAND2_X1 U10284 ( .A1(n8914), .A2(n8859), .ZN(n8839) );
  OAI211_X1 U10285 ( .C1(n8917), .C2(n8862), .A(n8840), .B(n8839), .ZN(
        P2_U3481) );
  INV_X1 U10286 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8843) );
  AOI21_X1 U10287 ( .B1(n8842), .B2(n10021), .A(n8841), .ZN(n8918) );
  MUX2_X1 U10288 ( .A(n8843), .B(n8918), .S(n10466), .Z(n8844) );
  OAI21_X1 U10289 ( .B1(n8921), .B2(n8867), .A(n8844), .ZN(P2_U3480) );
  INV_X1 U10290 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8848) );
  INV_X1 U10291 ( .A(n8845), .ZN(n8846) );
  AOI21_X1 U10292 ( .B1(n8847), .B2(n10021), .A(n8846), .ZN(n8922) );
  MUX2_X1 U10293 ( .A(n8848), .B(n8922), .S(n10466), .Z(n8849) );
  OAI21_X1 U10294 ( .B1(n8925), .B2(n8867), .A(n8849), .ZN(P2_U3479) );
  MUX2_X1 U10295 ( .A(n8926), .B(P2_REG1_REG_19__SCAN_IN), .S(n10463), .Z(
        n8852) );
  INV_X1 U10296 ( .A(n8850), .ZN(n8927) );
  OAI22_X1 U10297 ( .A1(n8928), .A2(n8862), .B1(n8927), .B2(n8867), .ZN(n8851)
         );
  AOI21_X1 U10298 ( .B1(n10046), .B2(n8854), .A(n8853), .ZN(n8931) );
  MUX2_X1 U10299 ( .A(n8855), .B(n8931), .S(n10466), .Z(n8856) );
  OAI21_X1 U10300 ( .B1(n8862), .B2(n8934), .A(n8856), .ZN(P2_U3477) );
  INV_X1 U10301 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n10297) );
  MUX2_X1 U10302 ( .A(n8936), .B(n10297), .S(n10463), .Z(n8858) );
  NAND2_X1 U10303 ( .A1(n8937), .A2(n8859), .ZN(n8857) );
  OAI211_X1 U10304 ( .C1(n8940), .C2(n8862), .A(n8858), .B(n8857), .ZN(
        P2_U3476) );
  MUX2_X1 U10305 ( .A(n10226), .B(n8941), .S(n10466), .Z(n8861) );
  NAND2_X1 U10306 ( .A1(n8944), .A2(n8859), .ZN(n8860) );
  OAI211_X1 U10307 ( .C1(n8862), .C2(n8948), .A(n8861), .B(n8860), .ZN(
        P2_U3475) );
  AOI21_X1 U10308 ( .B1(n10021), .B2(n8864), .A(n8863), .ZN(n8949) );
  MUX2_X1 U10309 ( .A(n8865), .B(n8949), .S(n10466), .Z(n8866) );
  OAI21_X1 U10310 ( .B1(n8953), .B2(n8867), .A(n8866), .ZN(P2_U3474) );
  MUX2_X1 U10311 ( .A(n8868), .B(P2_REG1_REG_0__SCAN_IN), .S(n10463), .Z(
        P2_U3459) );
  INV_X1 U10312 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8873) );
  NAND2_X1 U10313 ( .A1(n8869), .A2(n8943), .ZN(n8872) );
  INV_X1 U10314 ( .A(n8870), .ZN(n8871) );
  NAND2_X1 U10315 ( .A1(n8871), .A2(n10047), .ZN(n8874) );
  OAI211_X1 U10316 ( .C1(n8873), .C2(n10047), .A(n8872), .B(n8874), .ZN(
        P2_U3458) );
  NAND2_X1 U10317 ( .A1(n10049), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8875) );
  OAI211_X1 U10318 ( .C1(n8876), .C2(n8952), .A(n8875), .B(n8874), .ZN(
        P2_U3457) );
  INV_X1 U10319 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8878) );
  MUX2_X1 U10320 ( .A(n8878), .B(n8877), .S(n10047), .Z(n8881) );
  NAND2_X1 U10321 ( .A1(n8879), .A2(n8943), .ZN(n8880) );
  OAI211_X1 U10322 ( .C1(n8882), .C2(n8947), .A(n8881), .B(n8880), .ZN(
        P2_U3455) );
  MUX2_X1 U10323 ( .A(n10311), .B(n8883), .S(n10047), .Z(n8886) );
  NAND2_X1 U10324 ( .A1(n8884), .A2(n8943), .ZN(n8885) );
  OAI211_X1 U10325 ( .C1(n8887), .C2(n8947), .A(n8886), .B(n8885), .ZN(
        P2_U3454) );
  INV_X1 U10326 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8889) );
  MUX2_X1 U10327 ( .A(n8889), .B(n8888), .S(n10047), .Z(n8892) );
  NAND2_X1 U10328 ( .A1(n8890), .A2(n8943), .ZN(n8891) );
  OAI211_X1 U10329 ( .C1(n8893), .C2(n8947), .A(n8892), .B(n8891), .ZN(
        P2_U3453) );
  INV_X1 U10330 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8895) );
  MUX2_X1 U10331 ( .A(n8895), .B(n8894), .S(n10047), .Z(n8898) );
  NAND2_X1 U10332 ( .A1(n8896), .A2(n8943), .ZN(n8897) );
  OAI211_X1 U10333 ( .C1(n8899), .C2(n8947), .A(n8898), .B(n8897), .ZN(
        P2_U3452) );
  MUX2_X1 U10334 ( .A(n8901), .B(n8900), .S(n10047), .Z(n8904) );
  NAND2_X1 U10335 ( .A1(n8902), .A2(n8943), .ZN(n8903) );
  OAI211_X1 U10336 ( .C1(n8905), .C2(n8947), .A(n8904), .B(n8903), .ZN(
        P2_U3451) );
  INV_X1 U10337 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8907) );
  MUX2_X1 U10338 ( .A(n8907), .B(n8906), .S(n10047), .Z(n8910) );
  NAND2_X1 U10339 ( .A1(n8908), .A2(n8943), .ZN(n8909) );
  OAI211_X1 U10340 ( .C1(n8911), .C2(n8947), .A(n8910), .B(n8909), .ZN(
        P2_U3450) );
  INV_X1 U10341 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8913) );
  MUX2_X1 U10342 ( .A(n8913), .B(n8912), .S(n10047), .Z(n8916) );
  NAND2_X1 U10343 ( .A1(n8914), .A2(n8943), .ZN(n8915) );
  OAI211_X1 U10344 ( .C1(n8917), .C2(n8947), .A(n8916), .B(n8915), .ZN(
        P2_U3449) );
  INV_X1 U10345 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8919) );
  MUX2_X1 U10346 ( .A(n8919), .B(n8918), .S(n10047), .Z(n8920) );
  OAI21_X1 U10347 ( .B1(n8921), .B2(n8952), .A(n8920), .ZN(P2_U3448) );
  INV_X1 U10348 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8923) );
  MUX2_X1 U10349 ( .A(n8923), .B(n8922), .S(n10047), .Z(n8924) );
  OAI21_X1 U10350 ( .B1(n8925), .B2(n8952), .A(n8924), .ZN(P2_U3447) );
  MUX2_X1 U10351 ( .A(n8926), .B(P2_REG0_REG_19__SCAN_IN), .S(n10049), .Z(
        n8930) );
  OAI22_X1 U10352 ( .A1(n8928), .A2(n8947), .B1(n8927), .B2(n8952), .ZN(n8929)
         );
  INV_X1 U10353 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8932) );
  MUX2_X1 U10354 ( .A(n8932), .B(n8931), .S(n10047), .Z(n8933) );
  OAI21_X1 U10355 ( .B1(n8934), .B2(n8947), .A(n8933), .ZN(P2_U3444) );
  INV_X1 U10356 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8935) );
  MUX2_X1 U10357 ( .A(n8936), .B(n8935), .S(n10049), .Z(n8939) );
  NAND2_X1 U10358 ( .A1(n8937), .A2(n8943), .ZN(n8938) );
  OAI211_X1 U10359 ( .C1(n8940), .C2(n8947), .A(n8939), .B(n8938), .ZN(
        P2_U3441) );
  INV_X1 U10360 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8942) );
  MUX2_X1 U10361 ( .A(n8942), .B(n8941), .S(n10047), .Z(n8946) );
  NAND2_X1 U10362 ( .A1(n8944), .A2(n8943), .ZN(n8945) );
  OAI211_X1 U10363 ( .C1(n8948), .C2(n8947), .A(n8946), .B(n8945), .ZN(
        P2_U3438) );
  INV_X1 U10364 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8950) );
  MUX2_X1 U10365 ( .A(n8950), .B(n8949), .S(n10047), .Z(n8951) );
  OAI21_X1 U10366 ( .B1(n8953), .B2(n8952), .A(n8951), .ZN(P2_U3435) );
  INV_X1 U10367 ( .A(n9626), .ZN(n8958) );
  NOR4_X1 U10368 ( .A1(n8954), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n8955), .ZN(n8956) );
  AOI21_X1 U10369 ( .B1(n8963), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8956), .ZN(
        n8957) );
  OAI21_X1 U10370 ( .B1(n8958), .B2(n8965), .A(n8957), .ZN(P2_U3264) );
  AOI21_X1 U10371 ( .B1(n8963), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8959), .ZN(
        n8960) );
  OAI21_X1 U10372 ( .B1(n8961), .B2(n8965), .A(n8960), .ZN(P2_U3267) );
  AOI21_X1 U10373 ( .B1(n8963), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8962), .ZN(
        n8964) );
  OAI21_X1 U10374 ( .B1(n8966), .B2(n8965), .A(n8964), .ZN(P2_U3268) );
  MUX2_X1 U10375 ( .A(n8967), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10376 ( .A(n8968), .ZN(n8969) );
  NAND2_X1 U10377 ( .A1(n8970), .A2(n8969), .ZN(n8982) );
  NAND2_X1 U10378 ( .A1(n9543), .A2(n8971), .ZN(n8973) );
  NAND2_X1 U10379 ( .A1(n9174), .A2(n6152), .ZN(n8972) );
  NAND2_X1 U10380 ( .A1(n8973), .A2(n8972), .ZN(n8974) );
  XNOR2_X1 U10381 ( .A(n8974), .B(n5963), .ZN(n8978) );
  INV_X1 U10382 ( .A(n8978), .ZN(n8980) );
  AND2_X1 U10383 ( .A1(n9174), .A2(n8975), .ZN(n8976) );
  AOI21_X1 U10384 ( .B1(n9543), .B2(n6152), .A(n8976), .ZN(n8977) );
  INV_X1 U10385 ( .A(n8977), .ZN(n8979) );
  AOI21_X1 U10386 ( .B1(n8980), .B2(n8979), .A(n9030), .ZN(n8981) );
  AOI21_X1 U10387 ( .B1(n8986), .B2(n8982), .A(n8981), .ZN(n8987) );
  INV_X1 U10388 ( .A(n8981), .ZN(n8984) );
  INV_X1 U10389 ( .A(n8982), .ZN(n8983) );
  NOR2_X1 U10390 ( .A1(n8984), .A2(n8983), .ZN(n8985) );
  AND2_X2 U10391 ( .A1(n8986), .A2(n8985), .ZN(n9026) );
  AND2_X1 U10392 ( .A1(n9175), .A2(n9131), .ZN(n8988) );
  AOI21_X1 U10393 ( .B1(n9173), .B2(n4509), .A(n8988), .ZN(n9377) );
  INV_X1 U10394 ( .A(n9708), .ZN(n9156) );
  AOI22_X1 U10395 ( .A1(n9381), .A2(n9156), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n8989) );
  OAI21_X1 U10396 ( .B1(n9377), .B2(n9153), .A(n8989), .ZN(n8990) );
  AOI21_X1 U10397 ( .B1(n9543), .B2(n9167), .A(n8990), .ZN(n8991) );
  NAND2_X1 U10398 ( .A1(n8992), .A2(n8991), .ZN(P1_U3214) );
  XNOR2_X1 U10399 ( .A(n8994), .B(n8993), .ZN(n8995) );
  XNOR2_X1 U10400 ( .A(n8996), .B(n8995), .ZN(n9002) );
  NAND2_X1 U10401 ( .A1(n9188), .A2(n9131), .ZN(n8998) );
  NAND2_X1 U10402 ( .A1(n9186), .A2(n4509), .ZN(n8997) );
  NAND2_X1 U10403 ( .A1(n8998), .A2(n8997), .ZN(n9599) );
  AOI22_X1 U10404 ( .A1(n9702), .A2(n9599), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n8999) );
  OAI21_X1 U10405 ( .B1(n9733), .B2(n9708), .A(n8999), .ZN(n9000) );
  AOI21_X1 U10406 ( .B1(n9735), .B2(n9167), .A(n9000), .ZN(n9001) );
  OAI21_X1 U10407 ( .B1(n9002), .B2(n9693), .A(n9001), .ZN(P1_U3215) );
  OAI21_X1 U10408 ( .B1(n9005), .B2(n9003), .A(n9004), .ZN(n9006) );
  NAND2_X1 U10409 ( .A1(n9006), .A2(n9096), .ZN(n9012) );
  INV_X1 U10410 ( .A(n9007), .ZN(n9421) );
  AND2_X1 U10411 ( .A1(n9179), .A2(n9131), .ZN(n9008) );
  AOI21_X1 U10412 ( .B1(n9177), .B2(n4509), .A(n9008), .ZN(n9418) );
  OAI22_X1 U10413 ( .A1(n9418), .A2(n9153), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9009), .ZN(n9010) );
  AOI21_X1 U10414 ( .B1(n9421), .B2(n9156), .A(n9010), .ZN(n9011) );
  OAI211_X1 U10415 ( .C1(n9424), .C2(n9704), .A(n9012), .B(n9011), .ZN(
        P1_U3216) );
  XOR2_X1 U10416 ( .A(n9014), .B(n9013), .Z(n9020) );
  NAND2_X1 U10417 ( .A1(n9181), .A2(n4509), .ZN(n9016) );
  NAND2_X1 U10418 ( .A1(n9183), .A2(n9131), .ZN(n9015) );
  NAND2_X1 U10419 ( .A1(n9016), .A2(n9015), .ZN(n9481) );
  AOI22_X1 U10420 ( .A1(n9702), .A2(n9481), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n9017) );
  OAI21_X1 U10421 ( .B1(n9475), .B2(n9708), .A(n9017), .ZN(n9018) );
  AOI21_X1 U10422 ( .B1(n9582), .B2(n9167), .A(n9018), .ZN(n9019) );
  OAI21_X1 U10423 ( .B1(n9020), .B2(n9693), .A(n9019), .ZN(P1_U3219) );
  NAND2_X1 U10424 ( .A1(n9538), .A2(n6152), .ZN(n9022) );
  NAND2_X1 U10425 ( .A1(n9173), .A2(n8975), .ZN(n9021) );
  NAND2_X1 U10426 ( .A1(n9022), .A2(n9021), .ZN(n9023) );
  XNOR2_X1 U10427 ( .A(n9023), .B(n5983), .ZN(n9025) );
  AOI22_X1 U10428 ( .A1(n9538), .A2(n8971), .B1(n6152), .B2(n9173), .ZN(n9024)
         );
  XNOR2_X1 U10429 ( .A(n9025), .B(n9024), .ZN(n9031) );
  OR4_X2 U10430 ( .A1(n9026), .A2(n9030), .A3(n9031), .A4(n9693), .ZN(n9035)
         );
  NAND3_X1 U10431 ( .A1(n9026), .A2(n9096), .A3(n9031), .ZN(n9034) );
  AOI22_X1 U10432 ( .A1(n9172), .A2(n4509), .B1(n9174), .B2(n9131), .ZN(n9362)
         );
  NOR2_X1 U10433 ( .A1(n9362), .A2(n9153), .ZN(n9029) );
  OAI22_X1 U10434 ( .A1(n9367), .A2(n9708), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9027), .ZN(n9028) );
  AOI211_X1 U10435 ( .C1(n9538), .C2(n6200), .A(n9029), .B(n9028), .ZN(n9033)
         );
  NAND3_X1 U10436 ( .A1(n9031), .A2(n9096), .A3(n9030), .ZN(n9032) );
  NAND4_X1 U10437 ( .A1(n9035), .A2(n9034), .A3(n9033), .A4(n9032), .ZN(
        P1_U3220) );
  XNOR2_X1 U10438 ( .A(n9036), .B(n9037), .ZN(n9043) );
  NAND2_X1 U10439 ( .A1(n9179), .A2(n4509), .ZN(n9039) );
  NAND2_X1 U10440 ( .A1(n9181), .A2(n9131), .ZN(n9038) );
  NAND2_X1 U10441 ( .A1(n9039), .A2(n9038), .ZN(n9451) );
  AOI22_X1 U10442 ( .A1(n9451), .A2(n9702), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9040) );
  OAI21_X1 U10443 ( .B1(n9445), .B2(n9708), .A(n9040), .ZN(n9041) );
  AOI21_X1 U10444 ( .B1(n9572), .B2(n6200), .A(n9041), .ZN(n9042) );
  OAI21_X1 U10445 ( .B1(n9043), .B2(n9693), .A(n9042), .ZN(P1_U3223) );
  XOR2_X1 U10446 ( .A(n9045), .B(n9044), .Z(n9053) );
  NAND2_X1 U10447 ( .A1(n9702), .A2(n9046), .ZN(n9048) );
  OAI211_X1 U10448 ( .C1(n9708), .C2(n9049), .A(n9048), .B(n9047), .ZN(n9050)
         );
  AOI21_X1 U10449 ( .B1(n9051), .B2(n6200), .A(n9050), .ZN(n9052) );
  OAI21_X1 U10450 ( .B1(n9053), .B2(n9693), .A(n9052), .ZN(P1_U3224) );
  OAI21_X1 U10451 ( .B1(n9055), .B2(n9054), .A(n6182), .ZN(n9056) );
  NAND2_X1 U10452 ( .A1(n9056), .A2(n9096), .ZN(n9061) );
  NAND2_X1 U10453 ( .A1(n9175), .A2(n4509), .ZN(n9058) );
  NAND2_X1 U10454 ( .A1(n9177), .A2(n9131), .ZN(n9057) );
  NAND2_X1 U10455 ( .A1(n9058), .A2(n9057), .ZN(n9396) );
  OAI22_X1 U10456 ( .A1(n9389), .A2(n9708), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10359), .ZN(n9059) );
  AOI21_X1 U10457 ( .B1(n9396), .B2(n9702), .A(n9059), .ZN(n9060) );
  OAI211_X1 U10458 ( .C1(n4754), .C2(n9704), .A(n9061), .B(n9060), .ZN(
        P1_U3225) );
  XOR2_X1 U10459 ( .A(n9064), .B(n9063), .Z(n9070) );
  NAND2_X1 U10460 ( .A1(n9184), .A2(n4509), .ZN(n9066) );
  NAND2_X1 U10461 ( .A1(n9186), .A2(n9131), .ZN(n9065) );
  NAND2_X1 U10462 ( .A1(n9066), .A2(n9065), .ZN(n9650) );
  NAND2_X1 U10463 ( .A1(n9702), .A2(n9650), .ZN(n9067) );
  NAND2_X1 U10464 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9281) );
  OAI211_X1 U10465 ( .C1(n9708), .C2(n9652), .A(n9067), .B(n9281), .ZN(n9068)
         );
  AOI21_X1 U10466 ( .B1(n9654), .B2(n9167), .A(n9068), .ZN(n9069) );
  OAI21_X1 U10467 ( .B1(n9070), .B2(n9693), .A(n9069), .ZN(P1_U3226) );
  XOR2_X1 U10468 ( .A(n9071), .B(n9072), .Z(n9078) );
  NAND2_X1 U10469 ( .A1(n9183), .A2(n4509), .ZN(n9074) );
  NAND2_X1 U10470 ( .A1(n9185), .A2(n9131), .ZN(n9073) );
  NAND2_X1 U10471 ( .A1(n9074), .A2(n9073), .ZN(n9509) );
  NAND2_X1 U10472 ( .A1(n9702), .A2(n9509), .ZN(n9075) );
  NAND2_X1 U10473 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9309) );
  OAI211_X1 U10474 ( .C1(n9708), .C2(n9514), .A(n9075), .B(n9309), .ZN(n9076)
         );
  AOI21_X1 U10475 ( .B1(n9521), .B2(n6200), .A(n9076), .ZN(n9077) );
  OAI21_X1 U10476 ( .B1(n9078), .B2(n9693), .A(n9077), .ZN(P1_U3228) );
  INV_X1 U10477 ( .A(n9004), .ZN(n9081) );
  NOR3_X1 U10478 ( .A1(n9081), .A2(n9080), .A3(n9079), .ZN(n9084) );
  INV_X1 U10479 ( .A(n9082), .ZN(n9083) );
  OAI21_X1 U10480 ( .B1(n9084), .B2(n9083), .A(n9096), .ZN(n9091) );
  NAND2_X1 U10481 ( .A1(n9176), .A2(n4509), .ZN(n9086) );
  NAND2_X1 U10482 ( .A1(n9178), .A2(n9131), .ZN(n9085) );
  NAND2_X1 U10483 ( .A1(n9086), .A2(n9085), .ZN(n9410) );
  INV_X1 U10484 ( .A(n9404), .ZN(n9088) );
  OAI22_X1 U10485 ( .A1(n9088), .A2(n9708), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9087), .ZN(n9089) );
  AOI21_X1 U10486 ( .B1(n9410), .B2(n9702), .A(n9089), .ZN(n9090) );
  OAI211_X1 U10487 ( .C1(n9406), .C2(n9704), .A(n9091), .B(n9090), .ZN(
        P1_U3229) );
  AOI21_X1 U10488 ( .B1(n9094), .B2(n9093), .A(n9092), .ZN(n9098) );
  OAI211_X1 U10489 ( .C1(n9098), .C2(n9097), .A(n9096), .B(n9095), .ZN(n9108)
         );
  NAND2_X1 U10490 ( .A1(n9100), .A2(n9099), .ZN(n9102) );
  INV_X1 U10491 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9101) );
  NOR2_X1 U10492 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9101), .ZN(n9264) );
  AOI21_X1 U10493 ( .B1(n9702), .B2(n9102), .A(n9264), .ZN(n9107) );
  NAND2_X1 U10494 ( .A1(n9167), .A2(n9883), .ZN(n9106) );
  INV_X1 U10495 ( .A(n9103), .ZN(n9104) );
  NAND2_X1 U10496 ( .A1(n9156), .A2(n9104), .ZN(n9105) );
  NAND4_X1 U10497 ( .A1(n9108), .A2(n9107), .A3(n9106), .A4(n9105), .ZN(
        P1_U3231) );
  XOR2_X1 U10498 ( .A(n9111), .B(n9110), .Z(n9112) );
  XNOR2_X1 U10499 ( .A(n9109), .B(n9112), .ZN(n9118) );
  NOR2_X1 U10500 ( .A1(n9708), .A2(n9466), .ZN(n9116) );
  AND2_X1 U10501 ( .A1(n9182), .A2(n9131), .ZN(n9113) );
  AOI21_X1 U10502 ( .B1(n9180), .B2(n4509), .A(n9113), .ZN(n9461) );
  OAI22_X1 U10503 ( .A1(n9461), .A2(n9153), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9114), .ZN(n9115) );
  AOI211_X1 U10504 ( .C1(n9578), .C2(n6200), .A(n9116), .B(n9115), .ZN(n9117)
         );
  OAI21_X1 U10505 ( .B1(n9118), .B2(n9693), .A(n9117), .ZN(P1_U3233) );
  XOR2_X1 U10506 ( .A(n9119), .B(n9120), .Z(n9127) );
  AOI22_X1 U10507 ( .A1(n9702), .A2(n9121), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n9122) );
  OAI21_X1 U10508 ( .B1(n9123), .B2(n9708), .A(n9122), .ZN(n9124) );
  AOI21_X1 U10509 ( .B1(n9125), .B2(n6200), .A(n9124), .ZN(n9126) );
  OAI21_X1 U10510 ( .B1(n9127), .B2(n9693), .A(n9126), .ZN(P1_U3234) );
  XNOR2_X1 U10511 ( .A(n4596), .B(n9128), .ZN(n9129) );
  XNOR2_X1 U10512 ( .A(n9130), .B(n9129), .ZN(n9137) );
  NAND2_X1 U10513 ( .A1(n9178), .A2(n4509), .ZN(n9133) );
  NAND2_X1 U10514 ( .A1(n9180), .A2(n9131), .ZN(n9132) );
  NAND2_X1 U10515 ( .A1(n9133), .A2(n9132), .ZN(n9438) );
  AOI22_X1 U10516 ( .A1(n9438), .A2(n9702), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9134) );
  OAI21_X1 U10517 ( .B1(n9432), .B2(n9708), .A(n9134), .ZN(n9135) );
  AOI21_X1 U10518 ( .B1(n9567), .B2(n9167), .A(n9135), .ZN(n9136) );
  OAI21_X1 U10519 ( .B1(n9137), .B2(n9693), .A(n9136), .ZN(P1_U3235) );
  INV_X1 U10520 ( .A(n9139), .ZN(n9142) );
  OR2_X1 U10521 ( .A1(n9140), .A2(n9139), .ZN(n9141) );
  AOI22_X1 U10522 ( .A1(n9138), .A2(n9142), .B1(n4607), .B2(n9141), .ZN(n9148)
         );
  AOI22_X1 U10523 ( .A1(n9702), .A2(n9143), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n9144) );
  OAI21_X1 U10524 ( .B1(n9145), .B2(n9708), .A(n9144), .ZN(n9146) );
  AOI21_X1 U10525 ( .B1(n9897), .B2(n6200), .A(n9146), .ZN(n9147) );
  OAI21_X1 U10526 ( .B1(n9148), .B2(n9693), .A(n9147), .ZN(P1_U3236) );
  XNOR2_X1 U10527 ( .A(n4826), .B(n9149), .ZN(n9150) );
  XNOR2_X1 U10528 ( .A(n9151), .B(n9150), .ZN(n9158) );
  AOI22_X1 U10529 ( .A1(n9182), .A2(n4509), .B1(n9131), .B2(n9184), .ZN(n9492)
         );
  OAI22_X1 U10530 ( .A1(n9153), .A2(n9492), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9152), .ZN(n9155) );
  NOR2_X1 U10531 ( .A1(n9501), .A2(n9704), .ZN(n9154) );
  AOI211_X1 U10532 ( .C1(n9156), .C2(n9497), .A(n9155), .B(n9154), .ZN(n9157)
         );
  OAI21_X1 U10533 ( .B1(n9158), .B2(n9693), .A(n9157), .ZN(P1_U3238) );
  XNOR2_X1 U10534 ( .A(n9161), .B(n9160), .ZN(n9162) );
  XNOR2_X1 U10535 ( .A(n9159), .B(n9162), .ZN(n9170) );
  AOI22_X1 U10536 ( .A1(n9702), .A2(n9163), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n9164) );
  OAI21_X1 U10537 ( .B1(n9165), .B2(n9708), .A(n9164), .ZN(n9166) );
  AOI21_X1 U10538 ( .B1(n9168), .B2(n9167), .A(n9166), .ZN(n9169) );
  OAI21_X1 U10539 ( .B1(n9170), .B2(n9693), .A(n9169), .ZN(P1_U3241) );
  MUX2_X1 U10540 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9171), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10541 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n5878), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10542 ( .A(n9172), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9198), .Z(
        P1_U3583) );
  MUX2_X1 U10543 ( .A(n9173), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9198), .Z(
        P1_U3582) );
  MUX2_X1 U10544 ( .A(n9174), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9198), .Z(
        P1_U3581) );
  MUX2_X1 U10545 ( .A(n9175), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9198), .Z(
        P1_U3580) );
  MUX2_X1 U10546 ( .A(n9176), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9198), .Z(
        P1_U3579) );
  MUX2_X1 U10547 ( .A(n9177), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9198), .Z(
        P1_U3578) );
  MUX2_X1 U10548 ( .A(n9178), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9198), .Z(
        P1_U3577) );
  MUX2_X1 U10549 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9179), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10550 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9180), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10551 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9181), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10552 ( .A(n9182), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9198), .Z(
        P1_U3573) );
  MUX2_X1 U10553 ( .A(n9183), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9198), .Z(
        P1_U3572) );
  MUX2_X1 U10554 ( .A(n9184), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9198), .Z(
        P1_U3571) );
  MUX2_X1 U10555 ( .A(n9185), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9198), .Z(
        P1_U3570) );
  MUX2_X1 U10556 ( .A(n9186), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9198), .Z(
        P1_U3569) );
  MUX2_X1 U10557 ( .A(n9187), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9198), .Z(
        P1_U3568) );
  MUX2_X1 U10558 ( .A(n9188), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9198), .Z(
        P1_U3567) );
  MUX2_X1 U10559 ( .A(n9189), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9198), .Z(
        P1_U3566) );
  MUX2_X1 U10560 ( .A(n9190), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9198), .Z(
        P1_U3565) );
  MUX2_X1 U10561 ( .A(n9191), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9198), .Z(
        P1_U3564) );
  MUX2_X1 U10562 ( .A(n9192), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9198), .Z(
        P1_U3563) );
  MUX2_X1 U10563 ( .A(n9193), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9198), .Z(
        P1_U3562) );
  MUX2_X1 U10564 ( .A(n9697), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9198), .Z(
        P1_U3561) );
  MUX2_X1 U10565 ( .A(n9194), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9198), .Z(
        P1_U3560) );
  MUX2_X1 U10566 ( .A(n9695), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9198), .Z(
        P1_U3559) );
  MUX2_X1 U10567 ( .A(n9195), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9198), .Z(
        P1_U3558) );
  MUX2_X1 U10568 ( .A(n9196), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9198), .Z(
        P1_U3557) );
  MUX2_X1 U10569 ( .A(n9197), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9198), .Z(
        P1_U3556) );
  MUX2_X1 U10570 ( .A(n5979), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9198), .Z(
        P1_U3555) );
  INV_X1 U10571 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9200) );
  OAI22_X1 U10572 ( .A1(n9344), .A2(n9200), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9199), .ZN(n9201) );
  AOI21_X1 U10573 ( .B1(n9202), .B2(n9724), .A(n9201), .ZN(n9210) );
  OAI211_X1 U10574 ( .C1(n9205), .C2(n9204), .A(n9338), .B(n9203), .ZN(n9209)
         );
  OAI211_X1 U10575 ( .C1(n9207), .C2(n9228), .A(n9720), .B(n9206), .ZN(n9208)
         );
  NAND3_X1 U10576 ( .A1(n9210), .A2(n9209), .A3(n9208), .ZN(P1_U3244) );
  OAI211_X1 U10577 ( .C1(n9213), .C2(n9212), .A(n9338), .B(n9211), .ZN(n9224)
         );
  INV_X1 U10578 ( .A(n9214), .ZN(n9218) );
  INV_X1 U10579 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9216) );
  NAND2_X1 U10580 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9215) );
  OAI21_X1 U10581 ( .B1(n9344), .B2(n9216), .A(n9215), .ZN(n9217) );
  AOI21_X1 U10582 ( .B1(n9724), .B2(n9218), .A(n9217), .ZN(n9223) );
  OAI211_X1 U10583 ( .C1(n9221), .C2(n9220), .A(n9720), .B(n9219), .ZN(n9222)
         );
  NAND3_X1 U10584 ( .A1(n9224), .A2(n9223), .A3(n9222), .ZN(P1_U3246) );
  NAND3_X1 U10585 ( .A1(n9225), .A2(n4511), .A3(n9226), .ZN(n9232) );
  OAI21_X1 U10586 ( .B1(n4511), .B2(P1_REG2_REG_0__SCAN_IN), .A(n9226), .ZN(
        n9709) );
  INV_X1 U10587 ( .A(n9227), .ZN(n9229) );
  AOI22_X1 U10588 ( .A1(n9230), .A2(n9709), .B1(n9229), .B2(n9228), .ZN(n9231)
         );
  NAND3_X1 U10589 ( .A1(n9232), .A2(P1_U3973), .A3(n9231), .ZN(n9730) );
  INV_X1 U10590 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9234) );
  OAI22_X1 U10591 ( .A1(n9344), .A2(n9234), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9233), .ZN(n9235) );
  AOI21_X1 U10592 ( .B1(n9724), .B2(n9236), .A(n9235), .ZN(n9245) );
  OAI211_X1 U10593 ( .C1(n9239), .C2(n9238), .A(n9338), .B(n9237), .ZN(n9244)
         );
  OAI211_X1 U10594 ( .C1(n9242), .C2(n9241), .A(n9720), .B(n9240), .ZN(n9243)
         );
  NAND4_X1 U10595 ( .A1(n9730), .A2(n9245), .A3(n9244), .A4(n9243), .ZN(
        P1_U3247) );
  OAI211_X1 U10596 ( .C1(n9248), .C2(n9247), .A(n9338), .B(n9246), .ZN(n9259)
         );
  INV_X1 U10597 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9250) );
  OAI21_X1 U10598 ( .B1(n9344), .B2(n9250), .A(n9249), .ZN(n9251) );
  AOI21_X1 U10599 ( .B1(n9724), .B2(n9252), .A(n9251), .ZN(n9258) );
  INV_X1 U10600 ( .A(n9253), .ZN(n9254) );
  OAI211_X1 U10601 ( .C1(n9256), .C2(n9255), .A(n9720), .B(n9254), .ZN(n9257)
         );
  NAND3_X1 U10602 ( .A1(n9259), .A2(n9258), .A3(n9257), .ZN(P1_U3248) );
  OAI21_X1 U10603 ( .B1(n9262), .B2(n9261), .A(n9260), .ZN(n9263) );
  NAND2_X1 U10604 ( .A1(n9263), .A2(n9720), .ZN(n9273) );
  AOI21_X1 U10605 ( .B1(n9715), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9264), .ZN(
        n9272) );
  OAI21_X1 U10606 ( .B1(n9267), .B2(n9266), .A(n9265), .ZN(n9268) );
  NAND2_X1 U10607 ( .A1(n9268), .A2(n9338), .ZN(n9271) );
  NAND2_X1 U10608 ( .A1(n9724), .A2(n9269), .ZN(n9270) );
  NAND4_X1 U10609 ( .A1(n9273), .A2(n9272), .A3(n9271), .A4(n9270), .ZN(
        P1_U3252) );
  NOR2_X1 U10610 ( .A1(n9274), .A2(n9283), .ZN(n9276) );
  NOR2_X1 U10611 ( .A1(n9276), .A2(n9275), .ZN(n9279) );
  MUX2_X1 U10612 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9277), .S(n9305), .Z(n9278) );
  NAND2_X1 U10613 ( .A1(n9279), .A2(n9278), .ZN(n9304) );
  OAI21_X1 U10614 ( .B1(n9279), .B2(n9278), .A(n9304), .ZN(n9294) );
  NAND2_X1 U10615 ( .A1(n9715), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9280) );
  OAI211_X1 U10616 ( .C1(n9311), .C2(n9282), .A(n9281), .B(n9280), .ZN(n9293)
         );
  NOR2_X1 U10617 ( .A1(n9284), .A2(n9283), .ZN(n9286) );
  MUX2_X1 U10618 ( .A(n9287), .B(P1_REG2_REG_16__SCAN_IN), .S(n9305), .Z(n9290) );
  OR2_X1 U10619 ( .A1(n9291), .A2(n9290), .ZN(n9298) );
  INV_X1 U10620 ( .A(n9298), .ZN(n9288) );
  AOI211_X1 U10621 ( .C1(n9291), .C2(n9290), .A(n9289), .B(n9288), .ZN(n9292)
         );
  AOI211_X1 U10622 ( .C1(n9338), .C2(n9294), .A(n9293), .B(n9292), .ZN(n9295)
         );
  INV_X1 U10623 ( .A(n9295), .ZN(P1_U3259) );
  OR2_X1 U10624 ( .A1(n9318), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9323) );
  NAND2_X1 U10625 ( .A1(n9318), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9296) );
  AND2_X1 U10626 ( .A1(n9323), .A2(n9296), .ZN(n9300) );
  NAND2_X1 U10627 ( .A1(n9305), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9297) );
  NAND2_X1 U10628 ( .A1(n9299), .A2(n9300), .ZN(n9324) );
  OAI21_X1 U10629 ( .B1(n9300), .B2(n9299), .A(n9324), .ZN(n9301) );
  NAND2_X1 U10630 ( .A1(n9301), .A2(n9720), .ZN(n9315) );
  NOR2_X1 U10631 ( .A1(n9310), .A2(n9302), .ZN(n9303) );
  AOI21_X1 U10632 ( .B1(n9302), .B2(n9310), .A(n9303), .ZN(n9307) );
  OAI21_X1 U10633 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n9305), .A(n9304), .ZN(
        n9306) );
  NAND2_X1 U10634 ( .A1(n9306), .A2(n9307), .ZN(n9317) );
  OAI21_X1 U10635 ( .B1(n9307), .B2(n9306), .A(n9317), .ZN(n9313) );
  NAND2_X1 U10636 ( .A1(n9715), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9308) );
  OAI211_X1 U10637 ( .C1(n9311), .C2(n9310), .A(n9309), .B(n9308), .ZN(n9312)
         );
  AOI21_X1 U10638 ( .B1(n9313), .B2(n9338), .A(n9312), .ZN(n9314) );
  NAND2_X1 U10639 ( .A1(n9315), .A2(n9314), .ZN(P1_U3260) );
  NAND2_X1 U10640 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9316) );
  OAI21_X1 U10641 ( .B1(n9344), .B2(n10067), .A(n9316), .ZN(n9322) );
  OAI21_X1 U10642 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9318), .A(n9317), .ZN(
        n9320) );
  NAND2_X1 U10643 ( .A1(n9325), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9334) );
  OAI21_X1 U10644 ( .B1(n9325), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9334), .ZN(
        n9319) );
  NOR2_X1 U10645 ( .A1(n9320), .A2(n9319), .ZN(n9336) );
  AOI211_X1 U10646 ( .C1(n9320), .C2(n9319), .A(n9727), .B(n9336), .ZN(n9321)
         );
  AOI211_X1 U10647 ( .C1(n9724), .C2(n9325), .A(n9322), .B(n9321), .ZN(n9330)
         );
  AND2_X1 U10648 ( .A1(n9324), .A2(n9323), .ZN(n9328) );
  NAND2_X1 U10649 ( .A1(n9325), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9331) );
  OR2_X1 U10650 ( .A1(n9325), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9326) );
  AND2_X1 U10651 ( .A1(n9331), .A2(n9326), .ZN(n9327) );
  NAND2_X1 U10652 ( .A1(n9328), .A2(n9327), .ZN(n9332) );
  OAI211_X1 U10653 ( .C1(n9328), .C2(n9327), .A(n9332), .B(n9720), .ZN(n9329)
         );
  NAND2_X1 U10654 ( .A1(n9330), .A2(n9329), .ZN(P1_U3261) );
  NAND2_X1 U10655 ( .A1(n9332), .A2(n9331), .ZN(n9333) );
  XNOR2_X1 U10656 ( .A(n9333), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9341) );
  INV_X1 U10657 ( .A(n9341), .ZN(n9339) );
  INV_X1 U10658 ( .A(n9334), .ZN(n9335) );
  NOR2_X1 U10659 ( .A1(n9336), .A2(n9335), .ZN(n9337) );
  XNOR2_X1 U10660 ( .A(n9337), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9340) );
  AOI22_X1 U10661 ( .A1(n9339), .A2(n9720), .B1(n9338), .B2(n9340), .ZN(n9342)
         );
  NAND2_X1 U10662 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9343) );
  NAND2_X1 U10663 ( .A1(n4656), .A2(n9353), .ZN(n9352) );
  XNOR2_X1 U10664 ( .A(n9524), .B(n9352), .ZN(n9526) );
  INV_X1 U10665 ( .A(n9345), .ZN(n9351) );
  NOR2_X1 U10666 ( .A1(n9347), .A2(n9346), .ZN(n9528) );
  NAND2_X1 U10667 ( .A1(n9516), .A2(n9528), .ZN(n9354) );
  OAI21_X1 U10668 ( .B1(n9516), .B2(n9348), .A(n9354), .ZN(n9349) );
  AOI21_X1 U10669 ( .B1(n9524), .B2(n9788), .A(n9349), .ZN(n9350) );
  OAI21_X1 U10670 ( .B1(n9526), .B2(n9351), .A(n9350), .ZN(P1_U3263) );
  OAI211_X1 U10671 ( .C1(n4656), .C2(n9353), .A(n9793), .B(n9352), .ZN(n9530)
         );
  OAI21_X1 U10672 ( .B1(n9516), .B2(n9355), .A(n9354), .ZN(n9356) );
  AOI21_X1 U10673 ( .B1(n9357), .B2(n9788), .A(n9356), .ZN(n9358) );
  OAI21_X1 U10674 ( .B1(n9530), .B2(n9661), .A(n9358), .ZN(P1_U3264) );
  XNOR2_X1 U10675 ( .A(n9359), .B(n9361), .ZN(n9540) );
  XOR2_X1 U10676 ( .A(n9361), .B(n9360), .Z(n9363) );
  OAI21_X1 U10677 ( .B1(n9363), .B2(n9765), .A(n9362), .ZN(n9536) );
  INV_X1 U10678 ( .A(n9379), .ZN(n9366) );
  INV_X1 U10679 ( .A(n9364), .ZN(n9365) );
  AOI211_X1 U10680 ( .C1(n9538), .C2(n9366), .A(n9600), .B(n9365), .ZN(n9537)
         );
  NAND2_X1 U10681 ( .A1(n9537), .A2(n9757), .ZN(n9370) );
  INV_X1 U10682 ( .A(n9367), .ZN(n9368) );
  AOI22_X1 U10683 ( .A1(n9368), .A2(n9786), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9785), .ZN(n9369) );
  OAI211_X1 U10684 ( .C1(n9371), .C2(n9500), .A(n9370), .B(n9369), .ZN(n9372)
         );
  AOI21_X1 U10685 ( .B1(n9536), .B2(n9516), .A(n9372), .ZN(n9373) );
  OAI21_X1 U10686 ( .B1(n9540), .B2(n9662), .A(n9373), .ZN(P1_U3265) );
  XNOR2_X1 U10687 ( .A(n9376), .B(n9375), .ZN(n9378) );
  OAI21_X1 U10688 ( .B1(n9378), .B2(n9765), .A(n9377), .ZN(n9541) );
  INV_X1 U10689 ( .A(n9543), .ZN(n9384) );
  AOI211_X1 U10690 ( .C1(n9543), .C2(n9380), .A(n9600), .B(n9379), .ZN(n9542)
         );
  NAND2_X1 U10691 ( .A1(n9542), .A2(n9757), .ZN(n9383) );
  AOI22_X1 U10692 ( .A1(n9381), .A2(n9786), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9785), .ZN(n9382) );
  OAI211_X1 U10693 ( .C1(n9384), .C2(n9500), .A(n9383), .B(n9382), .ZN(n9385)
         );
  AOI21_X1 U10694 ( .B1(n9541), .B2(n9516), .A(n9385), .ZN(n9386) );
  OAI21_X1 U10695 ( .B1(n9545), .B2(n9662), .A(n9386), .ZN(P1_U3266) );
  XNOR2_X1 U10696 ( .A(n9387), .B(n9394), .ZN(n9555) );
  AOI211_X1 U10697 ( .C1(n9552), .C2(n9402), .A(n9600), .B(n9388), .ZN(n9551)
         );
  INV_X1 U10698 ( .A(n9389), .ZN(n9390) );
  AOI22_X1 U10699 ( .A1(n9390), .A2(n9786), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9785), .ZN(n9391) );
  OAI21_X1 U10700 ( .B1(n4754), .B2(n9500), .A(n9391), .ZN(n9399) );
  INV_X1 U10701 ( .A(n9392), .ZN(n9393) );
  NOR2_X1 U10702 ( .A1(n9407), .A2(n9393), .ZN(n9395) );
  XNOR2_X1 U10703 ( .A(n9395), .B(n9394), .ZN(n9397) );
  AOI21_X1 U10704 ( .B1(n9397), .B2(n9782), .A(n9396), .ZN(n9554) );
  NOR2_X1 U10705 ( .A1(n9554), .A2(n9785), .ZN(n9398) );
  AOI211_X1 U10706 ( .C1(n9551), .C2(n9757), .A(n9399), .B(n9398), .ZN(n9400)
         );
  OAI21_X1 U10707 ( .B1(n9555), .B2(n9662), .A(n9400), .ZN(P1_U3268) );
  XNOR2_X1 U10708 ( .A(n9401), .B(n9408), .ZN(n9560) );
  INV_X1 U10709 ( .A(n9402), .ZN(n9403) );
  AOI211_X1 U10710 ( .C1(n9557), .C2(n4758), .A(n9600), .B(n9403), .ZN(n9556)
         );
  AOI22_X1 U10711 ( .A1(n9404), .A2(n9786), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9785), .ZN(n9405) );
  OAI21_X1 U10712 ( .B1(n9406), .B2(n9500), .A(n9405), .ZN(n9414) );
  NOR2_X1 U10713 ( .A1(n9407), .A2(n9765), .ZN(n9412) );
  OAI21_X1 U10714 ( .B1(n4555), .B2(n9409), .A(n9408), .ZN(n9411) );
  AOI21_X1 U10715 ( .B1(n9412), .B2(n9411), .A(n9410), .ZN(n9559) );
  NOR2_X1 U10716 ( .A1(n9559), .A2(n9785), .ZN(n9413) );
  AOI211_X1 U10717 ( .C1(n9556), .C2(n9757), .A(n9414), .B(n9413), .ZN(n9415)
         );
  OAI21_X1 U10718 ( .B1(n9560), .B2(n9662), .A(n9415), .ZN(P1_U3269) );
  XNOR2_X1 U10719 ( .A(n4586), .B(n9416), .ZN(n9565) );
  AOI21_X1 U10720 ( .B1(n9417), .B2(n9416), .A(n4555), .ZN(n9419) );
  OAI21_X1 U10721 ( .B1(n9419), .B2(n9765), .A(n9418), .ZN(n9561) );
  AOI211_X1 U10722 ( .C1(n9563), .C2(n9429), .A(n9600), .B(n9420), .ZN(n9562)
         );
  NAND2_X1 U10723 ( .A1(n9562), .A2(n9757), .ZN(n9423) );
  AOI22_X1 U10724 ( .A1(n9421), .A2(n9786), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9785), .ZN(n9422) );
  OAI211_X1 U10725 ( .C1(n9424), .C2(n9500), .A(n9423), .B(n9422), .ZN(n9425)
         );
  AOI21_X1 U10726 ( .B1(n9561), .B2(n9516), .A(n9425), .ZN(n9426) );
  OAI21_X1 U10727 ( .B1(n9565), .B2(n9662), .A(n9426), .ZN(P1_U3270) );
  XNOR2_X1 U10728 ( .A(n9428), .B(n9427), .ZN(n9570) );
  INV_X1 U10729 ( .A(n9444), .ZN(n9431) );
  INV_X1 U10730 ( .A(n9429), .ZN(n9430) );
  AOI211_X1 U10731 ( .C1(n9567), .C2(n9431), .A(n9600), .B(n9430), .ZN(n9566)
         );
  INV_X1 U10732 ( .A(n9432), .ZN(n9433) );
  AOI22_X1 U10733 ( .A1(n9433), .A2(n9786), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9785), .ZN(n9434) );
  OAI21_X1 U10734 ( .B1(n9435), .B2(n9500), .A(n9434), .ZN(n9441) );
  XNOR2_X1 U10735 ( .A(n9437), .B(n9436), .ZN(n9439) );
  AOI21_X1 U10736 ( .B1(n9439), .B2(n9782), .A(n9438), .ZN(n9569) );
  NOR2_X1 U10737 ( .A1(n9569), .A2(n9785), .ZN(n9440) );
  AOI211_X1 U10738 ( .C1(n9566), .C2(n9757), .A(n9441), .B(n9440), .ZN(n9442)
         );
  OAI21_X1 U10739 ( .B1(n9570), .B2(n9662), .A(n9442), .ZN(P1_U3271) );
  XNOR2_X1 U10740 ( .A(n9443), .B(n9449), .ZN(n9575) );
  AOI211_X1 U10741 ( .C1(n9572), .C2(n9463), .A(n9600), .B(n9444), .ZN(n9571)
         );
  INV_X1 U10742 ( .A(n9445), .ZN(n9446) );
  AOI22_X1 U10743 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(n9785), .B1(n9446), .B2(
        n9786), .ZN(n9447) );
  OAI21_X1 U10744 ( .B1(n9448), .B2(n9500), .A(n9447), .ZN(n9454) );
  XNOR2_X1 U10745 ( .A(n9450), .B(n9449), .ZN(n9452) );
  AOI21_X1 U10746 ( .B1(n9452), .B2(n9782), .A(n9451), .ZN(n9574) );
  NOR2_X1 U10747 ( .A1(n9574), .A2(n9785), .ZN(n9453) );
  AOI211_X1 U10748 ( .C1(n9571), .C2(n9757), .A(n9454), .B(n9453), .ZN(n9455)
         );
  OAI21_X1 U10749 ( .B1(n9575), .B2(n9662), .A(n9455), .ZN(P1_U3272) );
  XNOR2_X1 U10750 ( .A(n9457), .B(n9456), .ZN(n9580) );
  OAI211_X1 U10751 ( .C1(n9460), .C2(n9459), .A(n9458), .B(n9782), .ZN(n9462)
         );
  NAND2_X1 U10752 ( .A1(n9462), .A2(n9461), .ZN(n9577) );
  INV_X1 U10753 ( .A(n9474), .ZN(n9465) );
  INV_X1 U10754 ( .A(n9463), .ZN(n9464) );
  AOI211_X1 U10755 ( .C1(n9578), .C2(n9465), .A(n9600), .B(n9464), .ZN(n9576)
         );
  NAND2_X1 U10756 ( .A1(n9576), .A2(n9757), .ZN(n9469) );
  INV_X1 U10757 ( .A(n9466), .ZN(n9467) );
  AOI22_X1 U10758 ( .A1(n9785), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9467), .B2(
        n9786), .ZN(n9468) );
  OAI211_X1 U10759 ( .C1(n9470), .C2(n9500), .A(n9469), .B(n9468), .ZN(n9471)
         );
  AOI21_X1 U10760 ( .B1(n9516), .B2(n9577), .A(n9471), .ZN(n9472) );
  OAI21_X1 U10761 ( .B1(n9580), .B2(n9662), .A(n9472), .ZN(P1_U3273) );
  XOR2_X1 U10762 ( .A(n9479), .B(n9473), .Z(n9585) );
  AOI211_X1 U10763 ( .C1(n9582), .C2(n9495), .A(n9600), .B(n9474), .ZN(n9581)
         );
  INV_X1 U10764 ( .A(n9475), .ZN(n9476) );
  AOI22_X1 U10765 ( .A1(n9785), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9476), .B2(
        n9786), .ZN(n9477) );
  OAI21_X1 U10766 ( .B1(n9478), .B2(n9500), .A(n9477), .ZN(n9484) );
  XNOR2_X1 U10767 ( .A(n9480), .B(n9479), .ZN(n9482) );
  AOI21_X1 U10768 ( .B1(n9482), .B2(n9782), .A(n9481), .ZN(n9584) );
  NOR2_X1 U10769 ( .A1(n9584), .A2(n9785), .ZN(n9483) );
  AOI211_X1 U10770 ( .C1(n9581), .C2(n9757), .A(n9484), .B(n9483), .ZN(n9485)
         );
  OAI21_X1 U10771 ( .B1(n9585), .B2(n9662), .A(n9485), .ZN(P1_U3274) );
  XOR2_X1 U10772 ( .A(n9486), .B(n9488), .Z(n9590) );
  INV_X1 U10773 ( .A(n9487), .ZN(n9491) );
  AOI21_X1 U10774 ( .B1(n9504), .B2(n9489), .A(n9488), .ZN(n9490) );
  OAI21_X1 U10775 ( .B1(n9491), .B2(n9490), .A(n9782), .ZN(n9493) );
  NAND2_X1 U10776 ( .A1(n9493), .A2(n9492), .ZN(n9587) );
  INV_X1 U10777 ( .A(n9494), .ZN(n9517) );
  INV_X1 U10778 ( .A(n9495), .ZN(n9496) );
  AOI211_X1 U10779 ( .C1(n9588), .C2(n9517), .A(n9600), .B(n9496), .ZN(n9586)
         );
  NAND2_X1 U10780 ( .A1(n9586), .A2(n9757), .ZN(n9499) );
  AOI22_X1 U10781 ( .A1(n9785), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9497), .B2(
        n9786), .ZN(n9498) );
  OAI211_X1 U10782 ( .C1(n9501), .C2(n9500), .A(n9499), .B(n9498), .ZN(n9502)
         );
  AOI21_X1 U10783 ( .B1(n9516), .B2(n9587), .A(n9502), .ZN(n9503) );
  OAI21_X1 U10784 ( .B1(n9590), .B2(n9662), .A(n9503), .ZN(P1_U3275) );
  INV_X1 U10785 ( .A(n9504), .ZN(n9508) );
  AOI21_X1 U10786 ( .B1(n9647), .B2(n9506), .A(n9505), .ZN(n9507) );
  NOR3_X1 U10787 ( .A1(n9508), .A2(n9507), .A3(n9765), .ZN(n9510) );
  NOR2_X1 U10788 ( .A1(n9510), .A2(n9509), .ZN(n9667) );
  XNOR2_X1 U10789 ( .A(n9512), .B(n9511), .ZN(n9670) );
  NAND2_X1 U10790 ( .A1(n9670), .A2(n9797), .ZN(n9523) );
  OAI22_X1 U10791 ( .A1(n9516), .A2(n9515), .B1(n9514), .B2(n9513), .ZN(n9520)
         );
  INV_X1 U10792 ( .A(n9521), .ZN(n9668) );
  INV_X1 U10793 ( .A(n9659), .ZN(n9518) );
  OAI211_X1 U10794 ( .C1(n9668), .C2(n9518), .A(n9517), .B(n9793), .ZN(n9666)
         );
  NOR2_X1 U10795 ( .A1(n9666), .A2(n9661), .ZN(n9519) );
  AOI211_X1 U10796 ( .C1(n9788), .C2(n9521), .A(n9520), .B(n9519), .ZN(n9522)
         );
  OAI211_X1 U10797 ( .C1(n9785), .C2(n9667), .A(n9523), .B(n9522), .ZN(
        P1_U3276) );
  AOI21_X1 U10798 ( .B1(n9524), .B2(n9898), .A(n9528), .ZN(n9525) );
  OAI21_X1 U10799 ( .B1(n9526), .B2(n9600), .A(n9525), .ZN(n9605) );
  MUX2_X1 U10800 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9605), .S(n9936), .Z(
        P1_U3553) );
  INV_X1 U10801 ( .A(n9528), .ZN(n9529) );
  OAI211_X1 U10802 ( .C1(n4656), .C2(n9913), .A(n9530), .B(n9529), .ZN(n9606)
         );
  MUX2_X1 U10803 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9606), .S(n9936), .Z(
        P1_U3552) );
  NAND2_X1 U10804 ( .A1(n9531), .A2(n9916), .ZN(n9535) );
  MUX2_X1 U10805 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9607), .S(n9936), .Z(
        P1_U3551) );
  AOI211_X1 U10806 ( .C1(n9898), .C2(n9538), .A(n9537), .B(n9536), .ZN(n9539)
         );
  OAI21_X1 U10807 ( .B1(n9540), .B2(n9862), .A(n9539), .ZN(n9608) );
  MUX2_X1 U10808 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9608), .S(n9936), .Z(
        P1_U3550) );
  AOI211_X1 U10809 ( .C1(n9898), .C2(n9543), .A(n9542), .B(n9541), .ZN(n9544)
         );
  OAI21_X1 U10810 ( .B1(n9545), .B2(n9862), .A(n9544), .ZN(n9609) );
  MUX2_X1 U10811 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9609), .S(n9936), .Z(
        P1_U3549) );
  AOI22_X1 U10812 ( .A1(n9547), .A2(n9793), .B1(n9898), .B2(n9546), .ZN(n9548)
         );
  OAI211_X1 U10813 ( .C1(n9550), .C2(n9862), .A(n9549), .B(n9548), .ZN(n9610)
         );
  MUX2_X1 U10814 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9610), .S(n9936), .Z(
        P1_U3548) );
  AOI21_X1 U10815 ( .B1(n9898), .B2(n9552), .A(n9551), .ZN(n9553) );
  OAI211_X1 U10816 ( .C1(n9555), .C2(n9862), .A(n9554), .B(n9553), .ZN(n9611)
         );
  MUX2_X1 U10817 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9611), .S(n9936), .Z(
        P1_U3547) );
  AOI21_X1 U10818 ( .B1(n9898), .B2(n9557), .A(n9556), .ZN(n9558) );
  OAI211_X1 U10819 ( .C1(n9560), .C2(n9862), .A(n9559), .B(n9558), .ZN(n9612)
         );
  MUX2_X1 U10820 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9612), .S(n9936), .Z(
        P1_U3546) );
  AOI211_X1 U10821 ( .C1(n9898), .C2(n9563), .A(n9562), .B(n9561), .ZN(n9564)
         );
  OAI21_X1 U10822 ( .B1(n9565), .B2(n9862), .A(n9564), .ZN(n9613) );
  MUX2_X1 U10823 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9613), .S(n9936), .Z(
        P1_U3545) );
  AOI21_X1 U10824 ( .B1(n9898), .B2(n9567), .A(n9566), .ZN(n9568) );
  OAI211_X1 U10825 ( .C1(n9570), .C2(n9862), .A(n9569), .B(n9568), .ZN(n9614)
         );
  MUX2_X1 U10826 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9614), .S(n9936), .Z(
        P1_U3544) );
  AOI21_X1 U10827 ( .B1(n9898), .B2(n9572), .A(n9571), .ZN(n9573) );
  OAI211_X1 U10828 ( .C1(n9575), .C2(n9862), .A(n9574), .B(n9573), .ZN(n9615)
         );
  MUX2_X1 U10829 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9615), .S(n9936), .Z(
        P1_U3543) );
  AOI211_X1 U10830 ( .C1(n9898), .C2(n9578), .A(n9577), .B(n9576), .ZN(n9579)
         );
  OAI21_X1 U10831 ( .B1(n9580), .B2(n9862), .A(n9579), .ZN(n9616) );
  MUX2_X1 U10832 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9616), .S(n9936), .Z(
        P1_U3542) );
  AOI21_X1 U10833 ( .B1(n9898), .B2(n9582), .A(n9581), .ZN(n9583) );
  OAI211_X1 U10834 ( .C1(n9585), .C2(n9862), .A(n9584), .B(n9583), .ZN(n9617)
         );
  MUX2_X1 U10835 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9617), .S(n9936), .Z(
        P1_U3541) );
  AOI211_X1 U10836 ( .C1(n9898), .C2(n9588), .A(n9587), .B(n9586), .ZN(n9589)
         );
  OAI21_X1 U10837 ( .B1(n9590), .B2(n9862), .A(n9589), .ZN(n9618) );
  MUX2_X1 U10838 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9618), .S(n9936), .Z(
        P1_U3540) );
  AND2_X1 U10839 ( .A1(n9592), .A2(n9591), .ZN(n9594) );
  OAI21_X1 U10840 ( .B1(n9594), .B2(n9597), .A(n9593), .ZN(n9739) );
  INV_X1 U10841 ( .A(n9739), .ZN(n9603) );
  INV_X1 U10842 ( .A(n9595), .ZN(n9596) );
  AOI211_X1 U10843 ( .C1(n9597), .C2(n4603), .A(n9765), .B(n9596), .ZN(n9598)
         );
  AOI211_X1 U10844 ( .C1(n9739), .C2(n9905), .A(n9599), .B(n9598), .ZN(n9742)
         );
  AOI211_X1 U10845 ( .C1(n9735), .C2(n9601), .A(n9600), .B(n4595), .ZN(n9737)
         );
  AOI21_X1 U10846 ( .B1(n9898), .B2(n9735), .A(n9737), .ZN(n9602) );
  OAI211_X1 U10847 ( .C1(n9603), .C2(n9901), .A(n9742), .B(n9602), .ZN(n9619)
         );
  MUX2_X1 U10848 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9619), .S(n9936), .Z(
        P1_U3536) );
  MUX2_X1 U10849 ( .A(n9604), .B(P1_REG1_REG_0__SCAN_IN), .S(n9934), .Z(
        P1_U3522) );
  MUX2_X1 U10850 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9605), .S(n9919), .Z(
        P1_U3521) );
  MUX2_X1 U10851 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9606), .S(n9919), .Z(
        P1_U3520) );
  MUX2_X1 U10852 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9608), .S(n9919), .Z(
        P1_U3518) );
  MUX2_X1 U10853 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9609), .S(n9919), .Z(
        P1_U3517) );
  MUX2_X1 U10854 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9610), .S(n9919), .Z(
        P1_U3516) );
  MUX2_X1 U10855 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9611), .S(n9919), .Z(
        P1_U3515) );
  MUX2_X1 U10856 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9612), .S(n9919), .Z(
        P1_U3514) );
  MUX2_X1 U10857 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9613), .S(n9919), .Z(
        P1_U3513) );
  MUX2_X1 U10858 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9614), .S(n9919), .Z(
        P1_U3512) );
  MUX2_X1 U10859 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9615), .S(n9919), .Z(
        P1_U3511) );
  MUX2_X1 U10860 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9616), .S(n9919), .Z(
        P1_U3510) );
  MUX2_X1 U10861 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9617), .S(n9919), .Z(
        P1_U3509) );
  MUX2_X1 U10862 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9618), .S(n9919), .Z(
        P1_U3507) );
  MUX2_X1 U10863 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9619), .S(n9919), .Z(
        P1_U3495) );
  MUX2_X1 U10864 ( .A(n9620), .B(P1_D_REG_0__SCAN_IN), .S(n9833), .Z(P1_U3439)
         );
  NAND3_X1 U10865 ( .A1(n9622), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n9623) );
  OAI22_X1 U10866 ( .A1(n9621), .A2(n9623), .B1(n10265), .B2(n9633), .ZN(n9624) );
  AOI21_X1 U10867 ( .B1(n9626), .B2(n9625), .A(n9624), .ZN(n9627) );
  INV_X1 U10868 ( .A(n9627), .ZN(P1_U3324) );
  OAI222_X1 U10869 ( .A1(n9633), .A2(n9630), .B1(n9629), .B2(n9628), .C1(n5292), .C2(P1_U3086), .ZN(P1_U3325) );
  OAI222_X1 U10870 ( .A1(n9633), .A2(n9632), .B1(P1_U3086), .B2(n5294), .C1(
        n9629), .C2(n9631), .ZN(P1_U3326) );
  MUX2_X1 U10871 ( .A(n9634), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI21_X1 U10872 ( .B1(n9637), .B2(n9636), .A(n9635), .ZN(n9643) );
  INV_X1 U10873 ( .A(n9638), .ZN(n9640) );
  NOR2_X1 U10874 ( .A1(n9892), .A2(n9704), .ZN(n9639) );
  AOI211_X1 U10875 ( .C1(n9702), .C2(n9641), .A(n9640), .B(n9639), .ZN(n9642)
         );
  OAI21_X1 U10876 ( .B1(n9643), .B2(n9693), .A(n9642), .ZN(n9644) );
  INV_X1 U10877 ( .A(n9644), .ZN(n9645) );
  OAI21_X1 U10878 ( .B1(n9646), .B2(n9708), .A(n9645), .ZN(P1_U3217) );
  OAI21_X1 U10879 ( .B1(n9649), .B2(n9648), .A(n9647), .ZN(n9651) );
  AOI21_X1 U10880 ( .B1(n9651), .B2(n9782), .A(n9650), .ZN(n9672) );
  INV_X1 U10881 ( .A(n9652), .ZN(n9653) );
  AOI222_X1 U10882 ( .A1(n9654), .A2(n9788), .B1(n9653), .B2(n9786), .C1(
        P1_REG2_REG_16__SCAN_IN), .C2(n9785), .ZN(n9665) );
  NOR2_X1 U10883 ( .A1(n9656), .A2(n9655), .ZN(n9657) );
  OR2_X1 U10884 ( .A1(n9658), .A2(n9657), .ZN(n9671) );
  OAI211_X1 U10885 ( .C1(n9660), .C2(n9674), .A(n9793), .B(n9659), .ZN(n9673)
         );
  OAI22_X1 U10886 ( .A1(n9671), .A2(n9662), .B1(n9673), .B2(n9661), .ZN(n9663)
         );
  INV_X1 U10887 ( .A(n9663), .ZN(n9664) );
  OAI211_X1 U10888 ( .C1(n9785), .C2(n9672), .A(n9665), .B(n9664), .ZN(
        P1_U3277) );
  OAI211_X1 U10889 ( .C1(n9668), .C2(n9913), .A(n9667), .B(n9666), .ZN(n9669)
         );
  AOI21_X1 U10890 ( .B1(n9670), .B2(n9916), .A(n9669), .ZN(n9685) );
  AOI22_X1 U10891 ( .A1(n9936), .A2(n9685), .B1(n9302), .B2(n9934), .ZN(
        P1_U3539) );
  INV_X1 U10892 ( .A(n9671), .ZN(n9677) );
  INV_X1 U10893 ( .A(n9672), .ZN(n9676) );
  OAI21_X1 U10894 ( .B1(n9674), .B2(n9913), .A(n9673), .ZN(n9675) );
  AOI211_X1 U10895 ( .C1(n9677), .C2(n9916), .A(n9676), .B(n9675), .ZN(n9687)
         );
  AOI22_X1 U10896 ( .A1(n9936), .A2(n9687), .B1(n9277), .B2(n9934), .ZN(
        P1_U3538) );
  OAI211_X1 U10897 ( .C1(n9680), .C2(n9913), .A(n9679), .B(n9678), .ZN(n9681)
         );
  AOI21_X1 U10898 ( .B1(n9682), .B2(n9916), .A(n9681), .ZN(n9688) );
  AOI22_X1 U10899 ( .A1(n9936), .A2(n9688), .B1(n9683), .B2(n9934), .ZN(
        P1_U3537) );
  INV_X1 U10900 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9684) );
  AOI22_X1 U10901 ( .A1(n9919), .A2(n9685), .B1(n9684), .B2(n9918), .ZN(
        P1_U3504) );
  INV_X1 U10902 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9686) );
  AOI22_X1 U10903 ( .A1(n9919), .A2(n9687), .B1(n9686), .B2(n9918), .ZN(
        P1_U3501) );
  AOI22_X1 U10904 ( .A1(n9919), .A2(n9688), .B1(n5500), .B2(n9918), .ZN(
        P1_U3498) );
  XNOR2_X1 U10905 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10906 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10907 ( .A(n9690), .ZN(n9691) );
  NAND3_X1 U10908 ( .A1(n7512), .A2(n9692), .A3(n9691), .ZN(n9694) );
  AOI21_X1 U10909 ( .B1(n9689), .B2(n9694), .A(n9693), .ZN(n9706) );
  NAND2_X1 U10910 ( .A1(n9695), .A2(n9131), .ZN(n9699) );
  NAND2_X1 U10911 ( .A1(n9697), .A2(n4509), .ZN(n9698) );
  NAND2_X1 U10912 ( .A1(n9699), .A2(n9698), .ZN(n9767) );
  INV_X1 U10913 ( .A(n9700), .ZN(n9701) );
  AOI21_X1 U10914 ( .B1(n9702), .B2(n9767), .A(n9701), .ZN(n9703) );
  OAI21_X1 U10915 ( .B1(n9867), .B2(n9704), .A(n9703), .ZN(n9705) );
  NOR2_X1 U10916 ( .A1(n9706), .A2(n9705), .ZN(n9707) );
  OAI21_X1 U10917 ( .B1(n9769), .B2(n9708), .A(n9707), .ZN(P1_U3239) );
  AOI21_X1 U10918 ( .B1(n4511), .B2(n9710), .A(n9709), .ZN(n9711) );
  XNOR2_X1 U10919 ( .A(n9711), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9714) );
  AOI22_X1 U10920 ( .A1(n9715), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9712) );
  OAI21_X1 U10921 ( .B1(n9714), .B2(n9713), .A(n9712), .ZN(P1_U3243) );
  AOI22_X1 U10922 ( .A1(n9715), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n9732) );
  OAI21_X1 U10923 ( .B1(n9718), .B2(n9717), .A(n9716), .ZN(n9728) );
  OAI211_X1 U10924 ( .C1(n9722), .C2(n9721), .A(n9720), .B(n9719), .ZN(n9726)
         );
  NAND2_X1 U10925 ( .A1(n9724), .A2(n9723), .ZN(n9725) );
  OAI211_X1 U10926 ( .C1(n9728), .C2(n9727), .A(n9726), .B(n9725), .ZN(n9729)
         );
  INV_X1 U10927 ( .A(n9729), .ZN(n9731) );
  NAND3_X1 U10928 ( .A1(n9732), .A2(n9731), .A3(n9730), .ZN(P1_U3245) );
  INV_X1 U10929 ( .A(n9733), .ZN(n9734) );
  AOI222_X1 U10930 ( .A1(n9735), .A2(n9788), .B1(P1_REG2_REG_14__SCAN_IN), 
        .B2(n9785), .C1(n9786), .C2(n9734), .ZN(n9741) );
  INV_X1 U10931 ( .A(n9736), .ZN(n9738) );
  AOI22_X1 U10932 ( .A1(n9739), .A2(n9738), .B1(n9757), .B2(n9737), .ZN(n9740)
         );
  OAI211_X1 U10933 ( .C1(n9785), .C2(n9742), .A(n9741), .B(n9740), .ZN(
        P1_U3279) );
  INV_X1 U10934 ( .A(n9743), .ZN(n9748) );
  AOI21_X1 U10935 ( .B1(n9746), .B2(n9745), .A(n9744), .ZN(n9747) );
  NOR3_X1 U10936 ( .A1(n9748), .A2(n9747), .A3(n9765), .ZN(n9750) );
  NOR2_X1 U10937 ( .A1(n9750), .A2(n9749), .ZN(n9880) );
  INV_X1 U10938 ( .A(n9751), .ZN(n9752) );
  AOI222_X1 U10939 ( .A1(n9755), .A2(n9788), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n9785), .C1(n9786), .C2(n9752), .ZN(n9760) );
  XNOR2_X1 U10940 ( .A(n9753), .B(n9754), .ZN(n9882) );
  OAI211_X1 U10941 ( .C1(n4760), .C2(n4759), .A(n9793), .B(n9756), .ZN(n9879)
         );
  INV_X1 U10942 ( .A(n9879), .ZN(n9758) );
  AOI22_X1 U10943 ( .A1(n9882), .A2(n9797), .B1(n9758), .B2(n9757), .ZN(n9759)
         );
  OAI211_X1 U10944 ( .C1(n9785), .C2(n9880), .A(n9760), .B(n9759), .ZN(
        P1_U3285) );
  INV_X1 U10945 ( .A(n9761), .ZN(n9762) );
  NOR2_X1 U10946 ( .A1(n9763), .A2(n9762), .ZN(n9764) );
  AOI211_X1 U10947 ( .C1(n9772), .C2(n9766), .A(n9765), .B(n9764), .ZN(n9768)
         );
  NOR2_X1 U10948 ( .A1(n9768), .A2(n9767), .ZN(n9866) );
  INV_X1 U10949 ( .A(n9769), .ZN(n9770) );
  AOI222_X1 U10950 ( .A1(n9771), .A2(n9788), .B1(P1_REG2_REG_6__SCAN_IN), .B2(
        n9785), .C1(n9786), .C2(n9770), .ZN(n9778) );
  XNOR2_X1 U10951 ( .A(n9773), .B(n9772), .ZN(n9869) );
  OAI211_X1 U10952 ( .C1(n9775), .C2(n9867), .A(n9793), .B(n9774), .ZN(n9865)
         );
  INV_X1 U10953 ( .A(n9865), .ZN(n9776) );
  AOI22_X1 U10954 ( .A1(n9869), .A2(n9797), .B1(n9776), .B2(n9757), .ZN(n9777)
         );
  OAI211_X1 U10955 ( .C1(n9785), .C2(n9866), .A(n9778), .B(n9777), .ZN(
        P1_U3287) );
  XNOR2_X1 U10956 ( .A(n9779), .B(n9791), .ZN(n9783) );
  INV_X1 U10957 ( .A(n9780), .ZN(n9781) );
  AOI21_X1 U10958 ( .B1(n9783), .B2(n9782), .A(n9781), .ZN(n9853) );
  INV_X1 U10959 ( .A(n9784), .ZN(n9787) );
  XNOR2_X1 U10960 ( .A(n9790), .B(n9791), .ZN(n9856) );
  INV_X1 U10961 ( .A(n9792), .ZN(n9795) );
  OAI211_X1 U10962 ( .C1(n4839), .C2(n9795), .A(n9794), .B(n9793), .ZN(n9852)
         );
  INV_X1 U10963 ( .A(n9852), .ZN(n9796) );
  AOI22_X1 U10964 ( .A1(n9856), .A2(n9797), .B1(n9796), .B2(n9757), .ZN(n9798)
         );
  OAI211_X1 U10965 ( .C1(n9785), .C2(n9853), .A(n9799), .B(n9798), .ZN(
        P1_U3289) );
  INV_X1 U10966 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10120) );
  NOR2_X1 U10967 ( .A1(n9822), .A2(n10120), .ZN(P1_U3294) );
  INV_X1 U10968 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n9801) );
  NOR2_X1 U10969 ( .A1(n9822), .A2(n9801), .ZN(P1_U3295) );
  INV_X1 U10970 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n9802) );
  NOR2_X1 U10971 ( .A1(n9822), .A2(n9802), .ZN(P1_U3296) );
  INV_X1 U10972 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9803) );
  NOR2_X1 U10973 ( .A1(n9822), .A2(n9803), .ZN(P1_U3297) );
  INV_X1 U10974 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9804) );
  NOR2_X1 U10975 ( .A1(n9822), .A2(n9804), .ZN(P1_U3298) );
  INV_X1 U10976 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9805) );
  NOR2_X1 U10977 ( .A1(n9822), .A2(n9805), .ZN(P1_U3299) );
  INV_X1 U10978 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n9806) );
  NOR2_X1 U10979 ( .A1(n9830), .A2(n9806), .ZN(P1_U3300) );
  INV_X1 U10980 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9807) );
  NOR2_X1 U10981 ( .A1(n9830), .A2(n9807), .ZN(P1_U3301) );
  INV_X1 U10982 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9808) );
  NOR2_X1 U10983 ( .A1(n9822), .A2(n9808), .ZN(P1_U3302) );
  INV_X1 U10984 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9809) );
  NOR2_X1 U10985 ( .A1(n9822), .A2(n9809), .ZN(P1_U3303) );
  INV_X1 U10986 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9810) );
  NOR2_X1 U10987 ( .A1(n9822), .A2(n9810), .ZN(P1_U3304) );
  INV_X1 U10988 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9811) );
  NOR2_X1 U10989 ( .A1(n9822), .A2(n9811), .ZN(P1_U3305) );
  INV_X1 U10990 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9812) );
  NOR2_X1 U10991 ( .A1(n9822), .A2(n9812), .ZN(P1_U3306) );
  INV_X1 U10992 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n9813) );
  NOR2_X1 U10993 ( .A1(n9822), .A2(n9813), .ZN(P1_U3307) );
  INV_X1 U10994 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9814) );
  NOR2_X1 U10995 ( .A1(n9822), .A2(n9814), .ZN(P1_U3308) );
  INV_X1 U10996 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10283) );
  NOR2_X1 U10997 ( .A1(n9822), .A2(n10283), .ZN(P1_U3309) );
  INV_X1 U10998 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n9815) );
  NOR2_X1 U10999 ( .A1(n9822), .A2(n9815), .ZN(P1_U3310) );
  INV_X1 U11000 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9816) );
  NOR2_X1 U11001 ( .A1(n9822), .A2(n9816), .ZN(P1_U3311) );
  INV_X1 U11002 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9817) );
  NOR2_X1 U11003 ( .A1(n9822), .A2(n9817), .ZN(P1_U3312) );
  INV_X1 U11004 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9818) );
  NOR2_X1 U11005 ( .A1(n9822), .A2(n9818), .ZN(P1_U3313) );
  INV_X1 U11006 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9819) );
  NOR2_X1 U11007 ( .A1(n9830), .A2(n9819), .ZN(P1_U3314) );
  INV_X1 U11008 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n9820) );
  NOR2_X1 U11009 ( .A1(n9830), .A2(n9820), .ZN(P1_U3315) );
  INV_X1 U11010 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9821) );
  NOR2_X1 U11011 ( .A1(n9822), .A2(n9821), .ZN(P1_U3316) );
  INV_X1 U11012 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9823) );
  NOR2_X1 U11013 ( .A1(n9830), .A2(n9823), .ZN(P1_U3317) );
  INV_X1 U11014 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n9824) );
  NOR2_X1 U11015 ( .A1(n9830), .A2(n9824), .ZN(P1_U3318) );
  INV_X1 U11016 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9825) );
  NOR2_X1 U11017 ( .A1(n9830), .A2(n9825), .ZN(P1_U3319) );
  INV_X1 U11018 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9826) );
  NOR2_X1 U11019 ( .A1(n9830), .A2(n9826), .ZN(P1_U3320) );
  INV_X1 U11020 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9827) );
  NOR2_X1 U11021 ( .A1(n9830), .A2(n9827), .ZN(P1_U3321) );
  INV_X1 U11022 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9828) );
  NOR2_X1 U11023 ( .A1(n9830), .A2(n9828), .ZN(P1_U3322) );
  INV_X1 U11024 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n9829) );
  NOR2_X1 U11025 ( .A1(n9830), .A2(n9829), .ZN(P1_U3323) );
  AOI21_X1 U11026 ( .B1(n9833), .B2(n9832), .A(n9831), .ZN(P1_U3440) );
  AOI21_X1 U11027 ( .B1(n9898), .B2(n9835), .A(n9834), .ZN(n9839) );
  INV_X1 U11028 ( .A(n9901), .ZN(n9837) );
  OAI21_X1 U11029 ( .B1(n9837), .B2(n9905), .A(n9836), .ZN(n9838) );
  AND3_X1 U11030 ( .A1(n9840), .A2(n9839), .A3(n9838), .ZN(n9921) );
  INV_X1 U11031 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9841) );
  AOI22_X1 U11032 ( .A1(n9919), .A2(n9921), .B1(n9841), .B2(n9918), .ZN(
        P1_U3456) );
  OAI211_X1 U11033 ( .C1(n9844), .C2(n9913), .A(n9843), .B(n9842), .ZN(n9845)
         );
  AOI21_X1 U11034 ( .B1(n9846), .B2(n9916), .A(n9845), .ZN(n9922) );
  AOI22_X1 U11035 ( .A1(n9919), .A2(n9922), .B1(n5616), .B2(n9918), .ZN(
        P1_U3459) );
  OAI21_X1 U11036 ( .B1(n5754), .B2(n9913), .A(n9847), .ZN(n9849) );
  AOI211_X1 U11037 ( .C1(n9850), .C2(n9916), .A(n9849), .B(n9848), .ZN(n9923)
         );
  INV_X1 U11038 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9851) );
  AOI22_X1 U11039 ( .A1(n9919), .A2(n9923), .B1(n9851), .B2(n9918), .ZN(
        P1_U3462) );
  OAI21_X1 U11040 ( .B1(n4839), .B2(n9913), .A(n9852), .ZN(n9855) );
  INV_X1 U11041 ( .A(n9853), .ZN(n9854) );
  AOI211_X1 U11042 ( .C1(n9916), .C2(n9856), .A(n9855), .B(n9854), .ZN(n9924)
         );
  INV_X1 U11043 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9857) );
  AOI22_X1 U11044 ( .A1(n9919), .A2(n9924), .B1(n9857), .B2(n9918), .ZN(
        P1_U3465) );
  AOI21_X1 U11045 ( .B1(n9898), .B2(n9859), .A(n9858), .ZN(n9860) );
  OAI211_X1 U11046 ( .C1(n9863), .C2(n9862), .A(n9861), .B(n9860), .ZN(n9864)
         );
  INV_X1 U11047 ( .A(n9864), .ZN(n9926) );
  AOI22_X1 U11048 ( .A1(n9919), .A2(n9926), .B1(n5652), .B2(n9918), .ZN(
        P1_U3468) );
  OAI211_X1 U11049 ( .C1(n9867), .C2(n9913), .A(n9866), .B(n9865), .ZN(n9868)
         );
  AOI21_X1 U11050 ( .B1(n9916), .B2(n9869), .A(n9868), .ZN(n9927) );
  INV_X1 U11051 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9870) );
  AOI22_X1 U11052 ( .A1(n9919), .A2(n9927), .B1(n9870), .B2(n9918), .ZN(
        P1_U3471) );
  AOI21_X1 U11053 ( .B1(n9901), .B2(n9872), .A(n9871), .ZN(n9876) );
  NOR2_X1 U11054 ( .A1(n9873), .A2(n9913), .ZN(n9874) );
  NOR4_X1 U11055 ( .A1(n9877), .A2(n9876), .A3(n9875), .A4(n9874), .ZN(n9928)
         );
  INV_X1 U11056 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9878) );
  AOI22_X1 U11057 ( .A1(n9919), .A2(n9928), .B1(n9878), .B2(n9918), .ZN(
        P1_U3474) );
  OAI211_X1 U11058 ( .C1(n4759), .C2(n9913), .A(n9880), .B(n9879), .ZN(n9881)
         );
  AOI21_X1 U11059 ( .B1(n9916), .B2(n9882), .A(n9881), .ZN(n9929) );
  AOI22_X1 U11060 ( .A1(n9919), .A2(n9929), .B1(n5674), .B2(n9918), .ZN(
        P1_U3477) );
  INV_X1 U11061 ( .A(n9883), .ZN(n9885) );
  OAI21_X1 U11062 ( .B1(n9885), .B2(n9913), .A(n9884), .ZN(n9887) );
  AOI211_X1 U11063 ( .C1(n9916), .C2(n9888), .A(n9887), .B(n9886), .ZN(n9930)
         );
  INV_X1 U11064 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9889) );
  AOI22_X1 U11065 ( .A1(n9919), .A2(n9930), .B1(n9889), .B2(n9918), .ZN(
        P1_U3480) );
  OAI211_X1 U11066 ( .C1(n9892), .C2(n9913), .A(n9891), .B(n9890), .ZN(n9893)
         );
  AOI21_X1 U11067 ( .B1(n9894), .B2(n9916), .A(n9893), .ZN(n9931) );
  INV_X1 U11068 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9895) );
  AOI22_X1 U11069 ( .A1(n9919), .A2(n9931), .B1(n9895), .B2(n9918), .ZN(
        P1_U3483) );
  AOI21_X1 U11070 ( .B1(n9898), .B2(n9897), .A(n9896), .ZN(n9899) );
  OAI211_X1 U11071 ( .C1(n9902), .C2(n9901), .A(n9900), .B(n9899), .ZN(n9903)
         );
  AOI21_X1 U11072 ( .B1(n9905), .B2(n9904), .A(n9903), .ZN(n9932) );
  INV_X1 U11073 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10325) );
  AOI22_X1 U11074 ( .A1(n9919), .A2(n9932), .B1(n10325), .B2(n9918), .ZN(
        P1_U3486) );
  OAI211_X1 U11075 ( .C1(n5062), .C2(n9913), .A(n9907), .B(n9906), .ZN(n9908)
         );
  AOI21_X1 U11076 ( .B1(n9909), .B2(n9916), .A(n9908), .ZN(n9933) );
  INV_X1 U11077 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9910) );
  AOI22_X1 U11078 ( .A1(n9919), .A2(n9933), .B1(n9910), .B2(n9918), .ZN(
        P1_U3489) );
  OAI211_X1 U11079 ( .C1(n9914), .C2(n9913), .A(n9912), .B(n9911), .ZN(n9915)
         );
  AOI21_X1 U11080 ( .B1(n9917), .B2(n9916), .A(n9915), .ZN(n9935) );
  AOI22_X1 U11081 ( .A1(n9919), .A2(n9935), .B1(n5517), .B2(n9918), .ZN(
        P1_U3492) );
  AOI22_X1 U11082 ( .A1(n9936), .A2(n9921), .B1(n9920), .B2(n9934), .ZN(
        P1_U3523) );
  AOI22_X1 U11083 ( .A1(n9936), .A2(n9922), .B1(n6886), .B2(n9934), .ZN(
        P1_U3524) );
  AOI22_X1 U11084 ( .A1(n9936), .A2(n9923), .B1(n6887), .B2(n9934), .ZN(
        P1_U3525) );
  AOI22_X1 U11085 ( .A1(n9936), .A2(n9924), .B1(n6888), .B2(n9934), .ZN(
        P1_U3526) );
  AOI22_X1 U11086 ( .A1(n9936), .A2(n9926), .B1(n9925), .B2(n9934), .ZN(
        P1_U3527) );
  AOI22_X1 U11087 ( .A1(n9936), .A2(n9927), .B1(n6890), .B2(n9934), .ZN(
        P1_U3528) );
  AOI22_X1 U11088 ( .A1(n9936), .A2(n9928), .B1(n6891), .B2(n9934), .ZN(
        P1_U3529) );
  AOI22_X1 U11089 ( .A1(n9936), .A2(n9929), .B1(n6892), .B2(n9934), .ZN(
        P1_U3530) );
  AOI22_X1 U11090 ( .A1(n9936), .A2(n9930), .B1(n5666), .B2(n9934), .ZN(
        P1_U3531) );
  AOI22_X1 U11091 ( .A1(n9936), .A2(n9931), .B1(n6965), .B2(n9934), .ZN(
        P1_U3532) );
  AOI22_X1 U11092 ( .A1(n9936), .A2(n9932), .B1(n7135), .B2(n9934), .ZN(
        P1_U3533) );
  AOI22_X1 U11093 ( .A1(n9936), .A2(n9933), .B1(n5534), .B2(n9934), .ZN(
        P1_U3534) );
  AOI22_X1 U11094 ( .A1(n9936), .A2(n9935), .B1(n7421), .B2(n9934), .ZN(
        P1_U3535) );
  AOI22_X1 U11095 ( .A1(n9938), .A2(n9937), .B1(n9973), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n9953) );
  OAI21_X1 U11096 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n9940), .A(n9939), .ZN(
        n9951) );
  INV_X1 U11097 ( .A(n9941), .ZN(n9942) );
  NAND3_X1 U11098 ( .A1(n9944), .A2(n9943), .A3(n9942), .ZN(n9945) );
  AOI21_X1 U11099 ( .B1(n9960), .B2(n9945), .A(n9981), .ZN(n9950) );
  AOI21_X1 U11100 ( .B1(n10217), .B2(n9947), .A(n9946), .ZN(n9948) );
  NOR2_X1 U11101 ( .A1(n9948), .A2(n9986), .ZN(n9949) );
  AOI211_X1 U11102 ( .C1(n9991), .C2(n9951), .A(n9950), .B(n9949), .ZN(n9952)
         );
  OAI211_X1 U11103 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6406), .A(n9953), .B(
        n9952), .ZN(P2_U3195) );
  AOI22_X1 U11104 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n9973), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3151), .ZN(n9970) );
  OAI21_X1 U11105 ( .B1(n9956), .B2(n9955), .A(n9954), .ZN(n9968) );
  INV_X1 U11106 ( .A(n9957), .ZN(n9958) );
  NAND3_X1 U11107 ( .A1(n9960), .A2(n9959), .A3(n9958), .ZN(n9961) );
  AOI21_X1 U11108 ( .B1(n9962), .B2(n9961), .A(n9981), .ZN(n9967) );
  AOI21_X1 U11109 ( .B1(n4559), .B2(n9964), .A(n9963), .ZN(n9965) );
  NOR2_X1 U11110 ( .A1(n9965), .A2(n9986), .ZN(n9966) );
  AOI211_X1 U11111 ( .C1(n9991), .C2(n9968), .A(n9967), .B(n9966), .ZN(n9969)
         );
  OAI211_X1 U11112 ( .C1(n9995), .C2(n9971), .A(n9970), .B(n9969), .ZN(
        P2_U3196) );
  AOI22_X1 U11113 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n9973), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(P2_U3151), .ZN(n9993) );
  OAI21_X1 U11114 ( .B1(n9976), .B2(n9975), .A(n9974), .ZN(n9990) );
  INV_X1 U11115 ( .A(n9977), .ZN(n9978) );
  NAND3_X1 U11116 ( .A1(n9980), .A2(n9979), .A3(n9978), .ZN(n9982) );
  AOI21_X1 U11117 ( .B1(n9983), .B2(n9982), .A(n9981), .ZN(n9989) );
  AOI21_X1 U11118 ( .B1(n4560), .B2(n9985), .A(n9984), .ZN(n9987) );
  NOR2_X1 U11119 ( .A1(n9987), .A2(n9986), .ZN(n9988) );
  AOI211_X1 U11120 ( .C1(n9991), .C2(n9990), .A(n9989), .B(n9988), .ZN(n9992)
         );
  OAI211_X1 U11121 ( .C1(n9995), .C2(n9994), .A(n9993), .B(n9992), .ZN(
        P2_U3198) );
  INV_X1 U11122 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10001) );
  AOI22_X1 U11123 ( .A1(n9998), .A2(n9997), .B1(n10046), .B2(n9996), .ZN(n9999) );
  AND2_X1 U11124 ( .A1(n10000), .A2(n9999), .ZN(n10050) );
  AOI22_X1 U11125 ( .A1(n10049), .A2(n10001), .B1(n10050), .B2(n10047), .ZN(
        P2_U3396) );
  INV_X1 U11126 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10006) );
  OAI21_X1 U11127 ( .B1(n10003), .B2(n10029), .A(n10002), .ZN(n10004) );
  AOI21_X1 U11128 ( .B1(n10005), .B2(n10021), .A(n10004), .ZN(n10052) );
  AOI22_X1 U11129 ( .A1(n10049), .A2(n10006), .B1(n10052), .B2(n10047), .ZN(
        P2_U3399) );
  INV_X1 U11130 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10011) );
  OAI21_X1 U11131 ( .B1(n10008), .B2(n10029), .A(n10007), .ZN(n10009) );
  AOI21_X1 U11132 ( .B1(n10010), .B2(n10021), .A(n10009), .ZN(n10465) );
  AOI22_X1 U11133 ( .A1(n10049), .A2(n10011), .B1(n10465), .B2(n10047), .ZN(
        P2_U3402) );
  INV_X1 U11134 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10016) );
  NOR2_X1 U11135 ( .A1(n10029), .A2(n10012), .ZN(n10014) );
  AOI211_X1 U11136 ( .C1(n10021), .C2(n10015), .A(n10014), .B(n10013), .ZN(
        n10054) );
  AOI22_X1 U11137 ( .A1(n10049), .A2(n10016), .B1(n10054), .B2(n10047), .ZN(
        P2_U3405) );
  INV_X1 U11138 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10023) );
  INV_X1 U11139 ( .A(n10017), .ZN(n10022) );
  OAI21_X1 U11140 ( .B1(n10019), .B2(n10029), .A(n10018), .ZN(n10020) );
  AOI21_X1 U11141 ( .B1(n10022), .B2(n10021), .A(n10020), .ZN(n10056) );
  AOI22_X1 U11142 ( .A1(n10049), .A2(n10023), .B1(n10056), .B2(n10047), .ZN(
        P2_U3408) );
  INV_X1 U11143 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10028) );
  OAI22_X1 U11144 ( .A1(n10025), .A2(n10041), .B1(n10024), .B2(n10029), .ZN(
        n10026) );
  NOR2_X1 U11145 ( .A1(n10027), .A2(n10026), .ZN(n10057) );
  AOI22_X1 U11146 ( .A1(n10049), .A2(n10028), .B1(n10057), .B2(n10047), .ZN(
        P2_U3411) );
  INV_X1 U11147 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10035) );
  OAI22_X1 U11148 ( .A1(n10032), .A2(n10031), .B1(n10030), .B2(n10029), .ZN(
        n10033) );
  NOR2_X1 U11149 ( .A1(n10034), .A2(n10033), .ZN(n10058) );
  AOI22_X1 U11150 ( .A1(n10049), .A2(n10035), .B1(n10058), .B2(n10047), .ZN(
        P2_U3414) );
  INV_X1 U11151 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10040) );
  NOR2_X1 U11152 ( .A1(n10036), .A2(n10041), .ZN(n10038) );
  AOI211_X1 U11153 ( .C1(n10046), .C2(n10039), .A(n10038), .B(n10037), .ZN(
        n10059) );
  AOI22_X1 U11154 ( .A1(n10049), .A2(n10040), .B1(n10059), .B2(n10047), .ZN(
        P2_U3417) );
  INV_X1 U11155 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10048) );
  NOR2_X1 U11156 ( .A1(n10042), .A2(n10041), .ZN(n10044) );
  AOI211_X1 U11157 ( .C1(n10046), .C2(n10045), .A(n10044), .B(n10043), .ZN(
        n10060) );
  AOI22_X1 U11158 ( .A1(n10049), .A2(n10048), .B1(n10060), .B2(n10047), .ZN(
        P2_U3420) );
  AOI22_X1 U11159 ( .A1(n10466), .A2(n10050), .B1(n7013), .B2(n10463), .ZN(
        P2_U3461) );
  INV_X1 U11160 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10051) );
  AOI22_X1 U11161 ( .A1(n10466), .A2(n10052), .B1(n10051), .B2(n10463), .ZN(
        P2_U3462) );
  INV_X1 U11162 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10053) );
  AOI22_X1 U11163 ( .A1(n10466), .A2(n10054), .B1(n10053), .B2(n10463), .ZN(
        P2_U3464) );
  AOI22_X1 U11164 ( .A1(n10466), .A2(n10056), .B1(n10055), .B2(n10463), .ZN(
        P2_U3465) );
  AOI22_X1 U11165 ( .A1(n10466), .A2(n10057), .B1(n7064), .B2(n10463), .ZN(
        P2_U3466) );
  AOI22_X1 U11166 ( .A1(n10466), .A2(n10058), .B1(n7205), .B2(n10463), .ZN(
        P2_U3467) );
  AOI22_X1 U11167 ( .A1(n10466), .A2(n10059), .B1(n7225), .B2(n10463), .ZN(
        P2_U3468) );
  AOI22_X1 U11168 ( .A1(n10466), .A2(n10060), .B1(n7336), .B2(n10463), .ZN(
        P2_U3469) );
  OAI222_X1 U11169 ( .A1(n10065), .A2(n10064), .B1(n10065), .B2(n10063), .C1(
        n10062), .C2(n10061), .ZN(ADD_1068_U5) );
  XOR2_X1 U11170 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11171 ( .B1(n10068), .B2(n10067), .A(n10066), .ZN(n10069) );
  INV_X1 U11172 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10340) );
  XNOR2_X1 U11173 ( .A(n10069), .B(n10340), .ZN(ADD_1068_U55) );
  OAI21_X1 U11174 ( .B1(n10072), .B2(n10071), .A(n10070), .ZN(ADD_1068_U56) );
  OAI21_X1 U11175 ( .B1(n10075), .B2(n10074), .A(n10073), .ZN(ADD_1068_U57) );
  OAI21_X1 U11176 ( .B1(n10078), .B2(n10077), .A(n10076), .ZN(ADD_1068_U58) );
  OAI21_X1 U11177 ( .B1(n10081), .B2(n10080), .A(n10079), .ZN(ADD_1068_U59) );
  OAI21_X1 U11178 ( .B1(n10084), .B2(n10083), .A(n10082), .ZN(ADD_1068_U60) );
  OAI21_X1 U11179 ( .B1(n10087), .B2(n10086), .A(n10085), .ZN(ADD_1068_U61) );
  OAI21_X1 U11180 ( .B1(n10090), .B2(n10089), .A(n10088), .ZN(ADD_1068_U62) );
  OAI21_X1 U11181 ( .B1(n10093), .B2(n10092), .A(n10091), .ZN(ADD_1068_U63) );
  AOI22_X1 U11182 ( .A1(n7637), .A2(keyinput210), .B1(keyinput217), .B2(n5592), 
        .ZN(n10094) );
  OAI221_X1 U11183 ( .B1(n7637), .B2(keyinput210), .C1(n5592), .C2(keyinput217), .A(n10094), .ZN(n10104) );
  AOI22_X1 U11184 ( .A1(n10268), .A2(keyinput196), .B1(keyinput188), .B2(
        n10340), .ZN(n10095) );
  OAI221_X1 U11185 ( .B1(n10268), .B2(keyinput196), .C1(n10340), .C2(
        keyinput188), .A(n10095), .ZN(n10103) );
  AOI22_X1 U11186 ( .A1(n10098), .A2(keyinput216), .B1(keyinput147), .B2(
        n10097), .ZN(n10096) );
  OAI221_X1 U11187 ( .B1(n10098), .B2(keyinput216), .C1(n10097), .C2(
        keyinput147), .A(n10096), .ZN(n10102) );
  AOI22_X1 U11188 ( .A1(n10293), .A2(keyinput234), .B1(keyinput243), .B2(
        n10100), .ZN(n10099) );
  OAI221_X1 U11189 ( .B1(n10293), .B2(keyinput234), .C1(n10100), .C2(
        keyinput243), .A(n10099), .ZN(n10101) );
  NOR4_X1 U11190 ( .A1(n10104), .A2(n10103), .A3(n10102), .A4(n10101), .ZN(
        n10139) );
  AOI22_X1 U11191 ( .A1(n10328), .A2(keyinput149), .B1(keyinput246), .B2(
        n10283), .ZN(n10105) );
  OAI221_X1 U11192 ( .B1(n10328), .B2(keyinput149), .C1(n10283), .C2(
        keyinput246), .A(n10105), .ZN(n10115) );
  AOI22_X1 U11193 ( .A1(n10356), .A2(keyinput223), .B1(n10107), .B2(
        keyinput170), .ZN(n10106) );
  OAI221_X1 U11194 ( .B1(n10356), .B2(keyinput223), .C1(n10107), .C2(
        keyinput170), .A(n10106), .ZN(n10114) );
  AOI22_X1 U11195 ( .A1(n10358), .A2(keyinput220), .B1(keyinput237), .B2(
        n10109), .ZN(n10108) );
  OAI221_X1 U11196 ( .B1(n10358), .B2(keyinput220), .C1(n10109), .C2(
        keyinput237), .A(n10108), .ZN(n10113) );
  XNOR2_X1 U11197 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(keyinput222), .ZN(n10111)
         );
  XNOR2_X1 U11198 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput235), .ZN(n10110)
         );
  NAND2_X1 U11199 ( .A1(n10111), .A2(n10110), .ZN(n10112) );
  NOR4_X1 U11200 ( .A1(n10115), .A2(n10114), .A3(n10113), .A4(n10112), .ZN(
        n10138) );
  AOI22_X1 U11201 ( .A1(n8143), .A2(keyinput181), .B1(keyinput194), .B2(n5605), 
        .ZN(n10116) );
  OAI221_X1 U11202 ( .B1(n8143), .B2(keyinput181), .C1(n5605), .C2(keyinput194), .A(n10116), .ZN(n10126) );
  INV_X1 U11203 ( .A(SI_30_), .ZN(n10118) );
  AOI22_X1 U11204 ( .A1(n10118), .A2(keyinput205), .B1(n7619), .B2(keyinput169), .ZN(n10117) );
  OAI221_X1 U11205 ( .B1(n10118), .B2(keyinput205), .C1(n7619), .C2(
        keyinput169), .A(n10117), .ZN(n10125) );
  AOI22_X1 U11206 ( .A1(n10120), .A2(keyinput157), .B1(keyinput182), .B2(
        n10312), .ZN(n10119) );
  OAI221_X1 U11207 ( .B1(n10120), .B2(keyinput157), .C1(n10312), .C2(
        keyinput182), .A(n10119), .ZN(n10124) );
  AOI22_X1 U11208 ( .A1(n10122), .A2(keyinput195), .B1(keyinput155), .B2(n5616), .ZN(n10121) );
  OAI221_X1 U11209 ( .B1(n10122), .B2(keyinput195), .C1(n5616), .C2(
        keyinput155), .A(n10121), .ZN(n10123) );
  NOR4_X1 U11210 ( .A1(n10126), .A2(n10125), .A3(n10124), .A4(n10123), .ZN(
        n10137) );
  AOI22_X1 U11211 ( .A1(n10349), .A2(keyinput138), .B1(n10306), .B2(
        keyinput166), .ZN(n10127) );
  OAI221_X1 U11212 ( .B1(n10349), .B2(keyinput138), .C1(n10306), .C2(
        keyinput166), .A(n10127), .ZN(n10135) );
  AOI22_X1 U11213 ( .A1(n10311), .A2(keyinput135), .B1(keyinput219), .B2(n5565), .ZN(n10128) );
  OAI221_X1 U11214 ( .B1(n10311), .B2(keyinput135), .C1(n5565), .C2(
        keyinput219), .A(n10128), .ZN(n10134) );
  INV_X1 U11215 ( .A(SI_31_), .ZN(n10370) );
  AOI22_X1 U11216 ( .A1(n10308), .A2(keyinput143), .B1(keyinput227), .B2(
        n10370), .ZN(n10129) );
  OAI221_X1 U11217 ( .B1(n10308), .B2(keyinput143), .C1(n10370), .C2(
        keyinput227), .A(n10129), .ZN(n10133) );
  INV_X1 U11218 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10131) );
  AOI22_X1 U11219 ( .A1(n5254), .A2(keyinput183), .B1(keyinput207), .B2(n10131), .ZN(n10130) );
  OAI221_X1 U11220 ( .B1(n5254), .B2(keyinput183), .C1(n10131), .C2(
        keyinput207), .A(n10130), .ZN(n10132) );
  NOR4_X1 U11221 ( .A1(n10135), .A2(n10134), .A3(n10133), .A4(n10132), .ZN(
        n10136) );
  NAND4_X1 U11222 ( .A1(n10139), .A2(n10138), .A3(n10137), .A4(n10136), .ZN(
        n10462) );
  OAI22_X1 U11223 ( .A1(P1_D_REG_20__SCAN_IN), .A2(keyinput185), .B1(
        P1_REG3_REG_27__SCAN_IN), .B2(keyinput226), .ZN(n10140) );
  AOI221_X1 U11224 ( .B1(P1_D_REG_20__SCAN_IN), .B2(keyinput185), .C1(
        keyinput226), .C2(P1_REG3_REG_27__SCAN_IN), .A(n10140), .ZN(n10147) );
  OAI22_X1 U11225 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput228), .B1(
        P2_REG3_REG_7__SCAN_IN), .B2(keyinput152), .ZN(n10141) );
  AOI221_X1 U11226 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput228), .C1(
        keyinput152), .C2(P2_REG3_REG_7__SCAN_IN), .A(n10141), .ZN(n10146) );
  OAI22_X1 U11227 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput129), .B1(
        P1_IR_REG_3__SCAN_IN), .B2(keyinput224), .ZN(n10142) );
  AOI221_X1 U11228 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput129), .C1(
        keyinput224), .C2(P1_IR_REG_3__SCAN_IN), .A(n10142), .ZN(n10145) );
  OAI22_X1 U11229 ( .A1(SI_24_), .A2(keyinput203), .B1(P2_REG1_REG_10__SCAN_IN), .B2(keyinput168), .ZN(n10143) );
  AOI221_X1 U11230 ( .B1(SI_24_), .B2(keyinput203), .C1(keyinput168), .C2(
        P2_REG1_REG_10__SCAN_IN), .A(n10143), .ZN(n10144) );
  NAND4_X1 U11231 ( .A1(n10147), .A2(n10146), .A3(n10145), .A4(n10144), .ZN(
        n10175) );
  OAI22_X1 U11232 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(keyinput174), .B1(
        keyinput225), .B2(P1_REG3_REG_3__SCAN_IN), .ZN(n10148) );
  AOI221_X1 U11233 ( .B1(P2_IR_REG_8__SCAN_IN), .B2(keyinput174), .C1(
        P1_REG3_REG_3__SCAN_IN), .C2(keyinput225), .A(n10148), .ZN(n10155) );
  OAI22_X1 U11234 ( .A1(P2_REG0_REG_25__SCAN_IN), .A2(keyinput144), .B1(
        P1_REG2_REG_3__SCAN_IN), .B2(keyinput175), .ZN(n10149) );
  AOI221_X1 U11235 ( .B1(P2_REG0_REG_25__SCAN_IN), .B2(keyinput144), .C1(
        keyinput175), .C2(P1_REG2_REG_3__SCAN_IN), .A(n10149), .ZN(n10154) );
  OAI22_X1 U11236 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(keyinput130), .B1(
        P1_REG3_REG_14__SCAN_IN), .B2(keyinput201), .ZN(n10150) );
  AOI221_X1 U11237 ( .B1(P2_DATAO_REG_14__SCAN_IN), .B2(keyinput130), .C1(
        keyinput201), .C2(P1_REG3_REG_14__SCAN_IN), .A(n10150), .ZN(n10153) );
  OAI22_X1 U11238 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(keyinput197), .B1(
        keyinput137), .B2(P1_REG3_REG_5__SCAN_IN), .ZN(n10151) );
  AOI221_X1 U11239 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(keyinput197), .C1(
        P1_REG3_REG_5__SCAN_IN), .C2(keyinput137), .A(n10151), .ZN(n10152) );
  NAND4_X1 U11240 ( .A1(n10155), .A2(n10154), .A3(n10153), .A4(n10152), .ZN(
        n10174) );
  OAI22_X1 U11241 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(keyinput167), .B1(
        P1_REG0_REG_11__SCAN_IN), .B2(keyinput218), .ZN(n10156) );
  AOI221_X1 U11242 ( .B1(P2_IR_REG_5__SCAN_IN), .B2(keyinput167), .C1(
        keyinput218), .C2(P1_REG0_REG_11__SCAN_IN), .A(n10156), .ZN(n10163) );
  OAI22_X1 U11243 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(keyinput186), .B1(
        keyinput128), .B2(P1_REG2_REG_5__SCAN_IN), .ZN(n10157) );
  AOI221_X1 U11244 ( .B1(P2_IR_REG_2__SCAN_IN), .B2(keyinput186), .C1(
        P1_REG2_REG_5__SCAN_IN), .C2(keyinput128), .A(n10157), .ZN(n10162) );
  OAI22_X1 U11245 ( .A1(P1_REG0_REG_13__SCAN_IN), .A2(keyinput244), .B1(
        keyinput209), .B2(P2_DATAO_REG_31__SCAN_IN), .ZN(n10158) );
  AOI221_X1 U11246 ( .B1(P1_REG0_REG_13__SCAN_IN), .B2(keyinput244), .C1(
        P2_DATAO_REG_31__SCAN_IN), .C2(keyinput209), .A(n10158), .ZN(n10161)
         );
  OAI22_X1 U11247 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(keyinput229), .B1(
        P1_REG2_REG_19__SCAN_IN), .B2(keyinput142), .ZN(n10159) );
  AOI221_X1 U11248 ( .B1(P1_REG3_REG_28__SCAN_IN), .B2(keyinput229), .C1(
        keyinput142), .C2(P1_REG2_REG_19__SCAN_IN), .A(n10159), .ZN(n10160) );
  NAND4_X1 U11249 ( .A1(n10163), .A2(n10162), .A3(n10161), .A4(n10160), .ZN(
        n10173) );
  OAI22_X1 U11250 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput151), .B1(
        P2_REG1_REG_13__SCAN_IN), .B2(keyinput255), .ZN(n10164) );
  AOI221_X1 U11251 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput151), .C1(
        keyinput255), .C2(P2_REG1_REG_13__SCAN_IN), .A(n10164), .ZN(n10171) );
  OAI22_X1 U11252 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(keyinput198), .B1(
        keyinput238), .B2(P1_REG0_REG_5__SCAN_IN), .ZN(n10165) );
  AOI221_X1 U11253 ( .B1(P2_IR_REG_14__SCAN_IN), .B2(keyinput198), .C1(
        P1_REG0_REG_5__SCAN_IN), .C2(keyinput238), .A(n10165), .ZN(n10170) );
  OAI22_X1 U11254 ( .A1(P1_RD_REG_SCAN_IN), .A2(keyinput213), .B1(
        P1_D_REG_3__SCAN_IN), .B2(keyinput231), .ZN(n10166) );
  AOI221_X1 U11255 ( .B1(P1_RD_REG_SCAN_IN), .B2(keyinput213), .C1(keyinput231), .C2(P1_D_REG_3__SCAN_IN), .A(n10166), .ZN(n10169) );
  OAI22_X1 U11256 ( .A1(P1_D_REG_18__SCAN_IN), .A2(keyinput178), .B1(
        keyinput247), .B2(P1_ADDR_REG_11__SCAN_IN), .ZN(n10167) );
  AOI221_X1 U11257 ( .B1(P1_D_REG_18__SCAN_IN), .B2(keyinput178), .C1(
        P1_ADDR_REG_11__SCAN_IN), .C2(keyinput247), .A(n10167), .ZN(n10168) );
  NAND4_X1 U11258 ( .A1(n10171), .A2(n10170), .A3(n10169), .A4(n10168), .ZN(
        n10172) );
  NOR4_X1 U11259 ( .A1(n10175), .A2(n10174), .A3(n10173), .A4(n10172), .ZN(
        n10262) );
  OAI22_X1 U11260 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(keyinput211), .B1(
        keyinput199), .B2(P2_WR_REG_SCAN_IN), .ZN(n10176) );
  AOI221_X1 U11261 ( .B1(P2_REG2_REG_28__SCAN_IN), .B2(keyinput211), .C1(
        P2_WR_REG_SCAN_IN), .C2(keyinput199), .A(n10176), .ZN(n10183) );
  OAI22_X1 U11262 ( .A1(P2_REG0_REG_29__SCAN_IN), .A2(keyinput190), .B1(
        keyinput252), .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n10177) );
  AOI221_X1 U11263 ( .B1(P2_REG0_REG_29__SCAN_IN), .B2(keyinput190), .C1(
        P1_DATAO_REG_17__SCAN_IN), .C2(keyinput252), .A(n10177), .ZN(n10182)
         );
  OAI22_X1 U11264 ( .A1(P1_REG1_REG_23__SCAN_IN), .A2(keyinput251), .B1(
        P1_ADDR_REG_7__SCAN_IN), .B2(keyinput236), .ZN(n10178) );
  AOI221_X1 U11265 ( .B1(P1_REG1_REG_23__SCAN_IN), .B2(keyinput251), .C1(
        keyinput236), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n10178), .ZN(n10181) );
  OAI22_X1 U11266 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput187), .B1(
        P1_REG0_REG_15__SCAN_IN), .B2(keyinput240), .ZN(n10179) );
  AOI221_X1 U11267 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput187), .C1(
        keyinput240), .C2(P1_REG0_REG_15__SCAN_IN), .A(n10179), .ZN(n10180) );
  NAND4_X1 U11268 ( .A1(n10183), .A2(n10182), .A3(n10181), .A4(n10180), .ZN(
        n10211) );
  OAI22_X1 U11269 ( .A1(SI_20_), .A2(keyinput162), .B1(keyinput159), .B2(
        P1_REG0_REG_28__SCAN_IN), .ZN(n10184) );
  AOI221_X1 U11270 ( .B1(SI_20_), .B2(keyinput162), .C1(
        P1_REG0_REG_28__SCAN_IN), .C2(keyinput159), .A(n10184), .ZN(n10191) );
  OAI22_X1 U11271 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput184), .B1(
        keyinput141), .B2(P2_REG0_REG_0__SCAN_IN), .ZN(n10185) );
  AOI221_X1 U11272 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput184), .C1(
        P2_REG0_REG_0__SCAN_IN), .C2(keyinput141), .A(n10185), .ZN(n10190) );
  OAI22_X1 U11273 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(keyinput249), .B1(
        keyinput208), .B2(P1_REG0_REG_27__SCAN_IN), .ZN(n10186) );
  AOI221_X1 U11274 ( .B1(P2_DATAO_REG_15__SCAN_IN), .B2(keyinput249), .C1(
        P1_REG0_REG_27__SCAN_IN), .C2(keyinput208), .A(n10186), .ZN(n10189) );
  OAI22_X1 U11275 ( .A1(P2_D_REG_5__SCAN_IN), .A2(keyinput233), .B1(
        P2_REG1_REG_20__SCAN_IN), .B2(keyinput179), .ZN(n10187) );
  AOI221_X1 U11276 ( .B1(P2_D_REG_5__SCAN_IN), .B2(keyinput233), .C1(
        keyinput179), .C2(P2_REG1_REG_20__SCAN_IN), .A(n10187), .ZN(n10188) );
  NAND4_X1 U11277 ( .A1(n10191), .A2(n10190), .A3(n10189), .A4(n10188), .ZN(
        n10210) );
  OAI22_X1 U11278 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(keyinput136), .B1(
        keyinput215), .B2(P2_REG1_REG_17__SCAN_IN), .ZN(n10192) );
  AOI221_X1 U11279 ( .B1(P1_DATAO_REG_5__SCAN_IN), .B2(keyinput136), .C1(
        P2_REG1_REG_17__SCAN_IN), .C2(keyinput215), .A(n10192), .ZN(n10199) );
  OAI22_X1 U11280 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(keyinput165), .B1(
        P1_REG2_REG_14__SCAN_IN), .B2(keyinput202), .ZN(n10193) );
  AOI221_X1 U11281 ( .B1(P1_IR_REG_15__SCAN_IN), .B2(keyinput165), .C1(
        keyinput202), .C2(P1_REG2_REG_14__SCAN_IN), .A(n10193), .ZN(n10198) );
  OAI22_X1 U11282 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(keyinput254), .B1(
        keyinput230), .B2(P1_IR_REG_29__SCAN_IN), .ZN(n10194) );
  AOI221_X1 U11283 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(keyinput254), .C1(
        P1_IR_REG_29__SCAN_IN), .C2(keyinput230), .A(n10194), .ZN(n10197) );
  OAI22_X1 U11284 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput156), .B1(
        P2_REG0_REG_14__SCAN_IN), .B2(keyinput139), .ZN(n10195) );
  AOI221_X1 U11285 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput156), .C1(
        keyinput139), .C2(P2_REG0_REG_14__SCAN_IN), .A(n10195), .ZN(n10196) );
  NAND4_X1 U11286 ( .A1(n10199), .A2(n10198), .A3(n10197), .A4(n10196), .ZN(
        n10209) );
  OAI22_X1 U11287 ( .A1(SI_14_), .A2(keyinput172), .B1(keyinput145), .B2(
        P2_REG2_REG_12__SCAN_IN), .ZN(n10200) );
  AOI221_X1 U11288 ( .B1(SI_14_), .B2(keyinput172), .C1(
        P2_REG2_REG_12__SCAN_IN), .C2(keyinput145), .A(n10200), .ZN(n10207) );
  OAI22_X1 U11289 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(keyinput242), .B1(
        P2_ADDR_REG_2__SCAN_IN), .B2(keyinput193), .ZN(n10201) );
  AOI221_X1 U11290 ( .B1(P2_DATAO_REG_2__SCAN_IN), .B2(keyinput242), .C1(
        keyinput193), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n10201), .ZN(n10206) );
  OAI22_X1 U11291 ( .A1(P2_REG0_REG_24__SCAN_IN), .A2(keyinput250), .B1(
        P1_ADDR_REG_3__SCAN_IN), .B2(keyinput245), .ZN(n10202) );
  AOI221_X1 U11292 ( .B1(P2_REG0_REG_24__SCAN_IN), .B2(keyinput250), .C1(
        keyinput245), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n10202), .ZN(n10205) );
  OAI22_X1 U11293 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(keyinput212), .B1(
        P2_ADDR_REG_17__SCAN_IN), .B2(keyinput150), .ZN(n10203) );
  AOI221_X1 U11294 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(keyinput212), .C1(
        keyinput150), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n10203), .ZN(n10204) );
  NAND4_X1 U11295 ( .A1(n10207), .A2(n10206), .A3(n10205), .A4(n10204), .ZN(
        n10208) );
  NOR4_X1 U11296 ( .A1(n10211), .A2(n10210), .A3(n10209), .A4(n10208), .ZN(
        n10261) );
  AOI22_X1 U11297 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(keyinput146), .B1(n5930), 
        .B2(keyinput221), .ZN(n10212) );
  OAI221_X1 U11298 ( .B1(P2_IR_REG_1__SCAN_IN), .B2(keyinput146), .C1(n5930), 
        .C2(keyinput221), .A(n10212), .ZN(n10223) );
  AOI22_X1 U11299 ( .A1(n10281), .A2(keyinput161), .B1(keyinput189), .B2(
        n10214), .ZN(n10213) );
  OAI221_X1 U11300 ( .B1(n10281), .B2(keyinput161), .C1(n10214), .C2(
        keyinput189), .A(n10213), .ZN(n10222) );
  INV_X1 U11301 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n10216) );
  AOI22_X1 U11302 ( .A1(n10217), .A2(keyinput163), .B1(keyinput248), .B2(
        n10216), .ZN(n10215) );
  OAI221_X1 U11303 ( .B1(n10217), .B2(keyinput163), .C1(n10216), .C2(
        keyinput248), .A(n10215), .ZN(n10221) );
  AOI22_X1 U11304 ( .A1(n10219), .A2(keyinput180), .B1(keyinput239), .B2(
        n10267), .ZN(n10218) );
  OAI221_X1 U11305 ( .B1(n10219), .B2(keyinput180), .C1(n10267), .C2(
        keyinput239), .A(n10218), .ZN(n10220) );
  NOR4_X1 U11306 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        n10260) );
  OAI22_X1 U11307 ( .A1(n10339), .A2(keyinput192), .B1(n10291), .B2(
        keyinput132), .ZN(n10224) );
  AOI221_X1 U11308 ( .B1(n10339), .B2(keyinput192), .C1(keyinput132), .C2(
        n10291), .A(n10224), .ZN(n10228) );
  OAI22_X1 U11309 ( .A1(n10226), .A2(keyinput253), .B1(n5558), .B2(keyinput134), .ZN(n10225) );
  AOI221_X1 U11310 ( .B1(n10226), .B2(keyinput253), .C1(keyinput134), .C2(
        n5558), .A(n10225), .ZN(n10227) );
  AND2_X1 U11311 ( .A1(n10228), .A2(n10227), .ZN(n10258) );
  OAI22_X1 U11312 ( .A1(n8029), .A2(keyinput214), .B1(n5534), .B2(keyinput148), 
        .ZN(n10229) );
  AOI221_X1 U11313 ( .B1(n8029), .B2(keyinput214), .C1(keyinput148), .C2(n5534), .A(n10229), .ZN(n10257) );
  INV_X1 U11314 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10231) );
  OAI22_X1 U11315 ( .A1(n6891), .A2(keyinput133), .B1(n10231), .B2(keyinput200), .ZN(n10230) );
  AOI221_X1 U11316 ( .B1(n6891), .B2(keyinput133), .C1(keyinput200), .C2(
        n10231), .A(n10230), .ZN(n10256) );
  OAI22_X1 U11317 ( .A1(n10294), .A2(keyinput158), .B1(n10233), .B2(
        keyinput140), .ZN(n10232) );
  AOI221_X1 U11318 ( .B1(n10294), .B2(keyinput158), .C1(keyinput140), .C2(
        n10233), .A(n10232), .ZN(n10243) );
  OAI22_X1 U11319 ( .A1(n6238), .A2(keyinput171), .B1(n10235), .B2(keyinput160), .ZN(n10234) );
  AOI221_X1 U11320 ( .B1(n6238), .B2(keyinput171), .C1(keyinput160), .C2(
        n10235), .A(n10234), .ZN(n10242) );
  OAI22_X1 U11321 ( .A1(n10238), .A2(keyinput206), .B1(n10237), .B2(
        keyinput177), .ZN(n10236) );
  AOI221_X1 U11322 ( .B1(n10238), .B2(keyinput206), .C1(keyinput177), .C2(
        n10237), .A(n10236), .ZN(n10241) );
  OAI22_X1 U11323 ( .A1(n10364), .A2(keyinput131), .B1(n10361), .B2(
        keyinput204), .ZN(n10239) );
  AOI221_X1 U11324 ( .B1(n10364), .B2(keyinput131), .C1(keyinput204), .C2(
        n10361), .A(n10239), .ZN(n10240) );
  NAND4_X1 U11325 ( .A1(n10243), .A2(n10242), .A3(n10241), .A4(n10240), .ZN(
        n10254) );
  XNOR2_X1 U11326 ( .A(P2_IR_REG_23__SCAN_IN), .B(keyinput153), .ZN(n10247) );
  XNOR2_X1 U11327 ( .A(SI_0_), .B(keyinput176), .ZN(n10246) );
  XNOR2_X1 U11328 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput173), .ZN(n10245) );
  XNOR2_X1 U11329 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput232), .ZN(n10244) );
  NAND4_X1 U11330 ( .A1(n10247), .A2(n10246), .A3(n10245), .A4(n10244), .ZN(
        n10253) );
  XNOR2_X1 U11331 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput154), .ZN(n10251)
         );
  XNOR2_X1 U11332 ( .A(P1_REG3_REG_13__SCAN_IN), .B(keyinput164), .ZN(n10250)
         );
  XNOR2_X1 U11333 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput241), .ZN(n10249) );
  XNOR2_X1 U11334 ( .A(keyinput191), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n10248)
         );
  NAND4_X1 U11335 ( .A1(n10251), .A2(n10250), .A3(n10249), .A4(n10248), .ZN(
        n10252) );
  NOR3_X1 U11336 ( .A1(n10254), .A2(n10253), .A3(n10252), .ZN(n10255) );
  AND4_X1 U11337 ( .A1(n10258), .A2(n10257), .A3(n10256), .A4(n10255), .ZN(
        n10259) );
  NAND4_X1 U11338 ( .A1(n10262), .A2(n10261), .A3(n10260), .A4(n10259), .ZN(
        n10461) );
  AOI22_X1 U11339 ( .A1(P1_REG0_REG_13__SCAN_IN), .A2(keyinput116), .B1(
        P1_RD_REG_SCAN_IN), .B2(keyinput85), .ZN(n10263) );
  OAI221_X1 U11340 ( .B1(P1_REG0_REG_13__SCAN_IN), .B2(keyinput116), .C1(
        P1_RD_REG_SCAN_IN), .C2(keyinput85), .A(n10263), .ZN(n10275) );
  AOI22_X1 U11341 ( .A1(P1_REG0_REG_15__SCAN_IN), .A2(keyinput112), .B1(n10265), .B2(keyinput81), .ZN(n10264) );
  OAI221_X1 U11342 ( .B1(P1_REG0_REG_15__SCAN_IN), .B2(keyinput112), .C1(
        n10265), .C2(keyinput81), .A(n10264), .ZN(n10274) );
  AOI22_X1 U11343 ( .A1(n10268), .A2(keyinput68), .B1(keyinput111), .B2(n10267), .ZN(n10266) );
  OAI221_X1 U11344 ( .B1(n10268), .B2(keyinput68), .C1(n10267), .C2(
        keyinput111), .A(n10266), .ZN(n10273) );
  AOI22_X1 U11345 ( .A1(n10271), .A2(keyinput62), .B1(keyinput34), .B2(n10270), 
        .ZN(n10269) );
  OAI221_X1 U11346 ( .B1(n10271), .B2(keyinput62), .C1(n10270), .C2(keyinput34), .A(n10269), .ZN(n10272) );
  NOR4_X1 U11347 ( .A1(n10275), .A2(n10274), .A3(n10273), .A4(n10272), .ZN(
        n10323) );
  AOI22_X1 U11348 ( .A1(n10278), .A2(keyinput123), .B1(keyinput22), .B2(n10277), .ZN(n10276) );
  OAI221_X1 U11349 ( .B1(n10278), .B2(keyinput123), .C1(n10277), .C2(
        keyinput22), .A(n10276), .ZN(n10289) );
  AOI22_X1 U11350 ( .A1(n10281), .A2(keyinput33), .B1(keyinput11), .B2(n10280), 
        .ZN(n10279) );
  OAI221_X1 U11351 ( .B1(n10281), .B2(keyinput33), .C1(n10280), .C2(keyinput11), .A(n10279), .ZN(n10288) );
  AOI22_X1 U11352 ( .A1(n10284), .A2(keyinput124), .B1(keyinput118), .B2(
        n10283), .ZN(n10282) );
  OAI221_X1 U11353 ( .B1(n10284), .B2(keyinput124), .C1(n10283), .C2(
        keyinput118), .A(n10282), .ZN(n10287) );
  AOI22_X1 U11354 ( .A1(n8143), .A2(keyinput53), .B1(keyinput82), .B2(n7637), 
        .ZN(n10285) );
  OAI221_X1 U11355 ( .B1(n8143), .B2(keyinput53), .C1(n7637), .C2(keyinput82), 
        .A(n10285), .ZN(n10286) );
  NOR4_X1 U11356 ( .A1(n10289), .A2(n10288), .A3(n10287), .A4(n10286), .ZN(
        n10322) );
  AOI22_X1 U11357 ( .A1(n10291), .A2(keyinput4), .B1(n5254), .B2(keyinput55), 
        .ZN(n10290) );
  OAI221_X1 U11358 ( .B1(n10291), .B2(keyinput4), .C1(n5254), .C2(keyinput55), 
        .A(n10290), .ZN(n10303) );
  AOI22_X1 U11359 ( .A1(n10294), .A2(keyinput30), .B1(keyinput106), .B2(n10293), .ZN(n10292) );
  OAI221_X1 U11360 ( .B1(n10294), .B2(keyinput30), .C1(n10293), .C2(
        keyinput106), .A(n10292), .ZN(n10302) );
  AOI22_X1 U11361 ( .A1(n10297), .A2(keyinput87), .B1(n10296), .B2(keyinput59), 
        .ZN(n10295) );
  OAI221_X1 U11362 ( .B1(n10297), .B2(keyinput87), .C1(n10296), .C2(keyinput59), .A(n10295), .ZN(n10301) );
  XNOR2_X1 U11363 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput107), .ZN(n10299)
         );
  XNOR2_X1 U11364 ( .A(SI_0_), .B(keyinput48), .ZN(n10298) );
  NAND2_X1 U11365 ( .A1(n10299), .A2(n10298), .ZN(n10300) );
  NOR4_X1 U11366 ( .A1(n10303), .A2(n10302), .A3(n10301), .A4(n10300), .ZN(
        n10321) );
  AOI22_X1 U11367 ( .A1(n10306), .A2(keyinput38), .B1(keyinput108), .B2(n10305), .ZN(n10304) );
  OAI221_X1 U11368 ( .B1(n10306), .B2(keyinput38), .C1(n10305), .C2(
        keyinput108), .A(n10304), .ZN(n10319) );
  AOI22_X1 U11369 ( .A1(n10309), .A2(keyinput127), .B1(n10308), .B2(keyinput15), .ZN(n10307) );
  OAI221_X1 U11370 ( .B1(n10309), .B2(keyinput127), .C1(n10308), .C2(
        keyinput15), .A(n10307), .ZN(n10318) );
  AOI22_X1 U11371 ( .A1(n10312), .A2(keyinput54), .B1(n10311), .B2(keyinput7), 
        .ZN(n10310) );
  OAI221_X1 U11372 ( .B1(n10312), .B2(keyinput54), .C1(n10311), .C2(keyinput7), 
        .A(n10310), .ZN(n10317) );
  INV_X1 U11373 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10315) );
  AOI22_X1 U11374 ( .A1(n10315), .A2(keyinput74), .B1(keyinput65), .B2(n10314), 
        .ZN(n10313) );
  OAI221_X1 U11375 ( .B1(n10315), .B2(keyinput74), .C1(n10314), .C2(keyinput65), .A(n10313), .ZN(n10316) );
  NOR4_X1 U11376 ( .A1(n10319), .A2(n10318), .A3(n10317), .A4(n10316), .ZN(
        n10320) );
  NAND4_X1 U11377 ( .A1(n10323), .A2(n10322), .A3(n10321), .A4(n10320), .ZN(
        n10459) );
  AOI22_X1 U11378 ( .A1(n10326), .A2(keyinput121), .B1(keyinput90), .B2(n10325), .ZN(n10324) );
  OAI221_X1 U11379 ( .B1(n10326), .B2(keyinput121), .C1(n10325), .C2(
        keyinput90), .A(n10324), .ZN(n10337) );
  INV_X1 U11380 ( .A(SI_14_), .ZN(n10329) );
  AOI22_X1 U11381 ( .A1(n10329), .A2(keyinput44), .B1(n10328), .B2(keyinput21), 
        .ZN(n10327) );
  OAI221_X1 U11382 ( .B1(n10329), .B2(keyinput44), .C1(n10328), .C2(keyinput21), .A(n10327), .ZN(n10336) );
  AOI22_X1 U11383 ( .A1(n10331), .A2(keyinput1), .B1(keyinput14), .B2(n5431), 
        .ZN(n10330) );
  OAI221_X1 U11384 ( .B1(n10331), .B2(keyinput1), .C1(n5431), .C2(keyinput14), 
        .A(n10330), .ZN(n10335) );
  XNOR2_X1 U11385 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput102), .ZN(n10333) );
  XNOR2_X1 U11386 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput104), .ZN(n10332) );
  NAND2_X1 U11387 ( .A1(n10333), .A2(n10332), .ZN(n10334) );
  NOR4_X1 U11388 ( .A1(n10337), .A2(n10336), .A3(n10335), .A4(n10334), .ZN(
        n10383) );
  AOI22_X1 U11389 ( .A1(n10340), .A2(keyinput60), .B1(n10339), .B2(keyinput64), 
        .ZN(n10338) );
  OAI221_X1 U11390 ( .B1(n10340), .B2(keyinput60), .C1(n10339), .C2(keyinput64), .A(n10338), .ZN(n10354) );
  AOI22_X1 U11391 ( .A1(n10343), .A2(keyinput94), .B1(n10342), .B2(keyinput126), .ZN(n10341) );
  OAI221_X1 U11392 ( .B1(n10343), .B2(keyinput94), .C1(n10342), .C2(
        keyinput126), .A(n10341), .ZN(n10344) );
  INV_X1 U11393 ( .A(n10344), .ZN(n10346) );
  XNOR2_X1 U11394 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput18), .ZN(n10345) );
  NAND2_X1 U11395 ( .A1(n10346), .A2(n10345), .ZN(n10353) );
  AOI22_X1 U11396 ( .A1(n10349), .A2(keyinput10), .B1(keyinput56), .B2(n10348), 
        .ZN(n10347) );
  OAI221_X1 U11397 ( .B1(n10349), .B2(keyinput10), .C1(n10348), .C2(keyinput56), .A(n10347), .ZN(n10352) );
  XNOR2_X1 U11398 ( .A(n10350), .B(keyinput119), .ZN(n10351) );
  NOR4_X1 U11399 ( .A1(n10354), .A2(n10353), .A3(n10352), .A4(n10351), .ZN(
        n10382) );
  AOI22_X1 U11400 ( .A1(n5629), .A2(keyinput96), .B1(keyinput95), .B2(n10356), 
        .ZN(n10355) );
  OAI221_X1 U11401 ( .B1(n5629), .B2(keyinput96), .C1(n10356), .C2(keyinput95), 
        .A(n10355), .ZN(n10368) );
  AOI22_X1 U11402 ( .A1(n10359), .A2(keyinput69), .B1(n10358), .B2(keyinput92), 
        .ZN(n10357) );
  OAI221_X1 U11403 ( .B1(n10359), .B2(keyinput69), .C1(n10358), .C2(keyinput92), .A(n10357), .ZN(n10367) );
  AOI22_X1 U11404 ( .A1(n5534), .A2(keyinput20), .B1(n10361), .B2(keyinput76), 
        .ZN(n10360) );
  OAI221_X1 U11405 ( .B1(n5534), .B2(keyinput20), .C1(n10361), .C2(keyinput76), 
        .A(n10360), .ZN(n10366) );
  AOI22_X1 U11406 ( .A1(n10364), .A2(keyinput3), .B1(keyinput36), .B2(n10363), 
        .ZN(n10362) );
  OAI221_X1 U11407 ( .B1(n10364), .B2(keyinput3), .C1(n10363), .C2(keyinput36), 
        .A(n10362), .ZN(n10365) );
  NOR4_X1 U11408 ( .A1(n10368), .A2(n10367), .A3(n10366), .A4(n10365), .ZN(
        n10381) );
  AOI22_X1 U11409 ( .A1(n10371), .A2(keyinput2), .B1(keyinput99), .B2(n10370), 
        .ZN(n10369) );
  OAI221_X1 U11410 ( .B1(n10371), .B2(keyinput2), .C1(n10370), .C2(keyinput99), 
        .A(n10369), .ZN(n10379) );
  AOI22_X1 U11411 ( .A1(n5592), .A2(keyinput89), .B1(n8029), .B2(keyinput86), 
        .ZN(n10372) );
  OAI221_X1 U11412 ( .B1(n5592), .B2(keyinput89), .C1(n8029), .C2(keyinput86), 
        .A(n10372), .ZN(n10378) );
  AOI22_X1 U11413 ( .A1(n5484), .A2(keyinput73), .B1(n6238), .B2(keyinput43), 
        .ZN(n10373) );
  OAI221_X1 U11414 ( .B1(n5484), .B2(keyinput73), .C1(n6238), .C2(keyinput43), 
        .A(n10373), .ZN(n10377) );
  XOR2_X1 U11415 ( .A(n5565), .B(keyinput91), .Z(n10375) );
  XNOR2_X1 U11416 ( .A(P2_IR_REG_23__SCAN_IN), .B(keyinput25), .ZN(n10374) );
  NAND2_X1 U11417 ( .A1(n10375), .A2(n10374), .ZN(n10376) );
  NOR4_X1 U11418 ( .A1(n10379), .A2(n10378), .A3(n10377), .A4(n10376), .ZN(
        n10380) );
  NAND4_X1 U11419 ( .A1(n10383), .A2(n10382), .A3(n10381), .A4(n10380), .ZN(
        n10458) );
  AOI22_X1 U11420 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(keyinput9), .B1(
        P1_D_REG_31__SCAN_IN), .B2(keyinput29), .ZN(n10384) );
  OAI221_X1 U11421 ( .B1(P1_REG3_REG_5__SCAN_IN), .B2(keyinput9), .C1(
        P1_D_REG_31__SCAN_IN), .C2(keyinput29), .A(n10384), .ZN(n10391) );
  AOI22_X1 U11422 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(keyinput101), .B1(
        P2_REG0_REG_25__SCAN_IN), .B2(keyinput16), .ZN(n10385) );
  OAI221_X1 U11423 ( .B1(P1_REG3_REG_28__SCAN_IN), .B2(keyinput101), .C1(
        P2_REG0_REG_25__SCAN_IN), .C2(keyinput16), .A(n10385), .ZN(n10390) );
  AOI22_X1 U11424 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(keyinput114), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(keyinput26), .ZN(n10386) );
  OAI221_X1 U11425 ( .B1(P2_DATAO_REG_2__SCAN_IN), .B2(keyinput114), .C1(
        P2_DATAO_REG_6__SCAN_IN), .C2(keyinput26), .A(n10386), .ZN(n10389) );
  AOI22_X1 U11426 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(keyinput115), .B1(
        P1_D_REG_18__SCAN_IN), .B2(keyinput50), .ZN(n10387) );
  OAI221_X1 U11427 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(keyinput115), .C1(
        P1_D_REG_18__SCAN_IN), .C2(keyinput50), .A(n10387), .ZN(n10388) );
  NOR4_X1 U11428 ( .A1(n10391), .A2(n10390), .A3(n10389), .A4(n10388), .ZN(
        n10419) );
  AOI22_X1 U11429 ( .A1(P2_REG1_REG_20__SCAN_IN), .A2(keyinput51), .B1(
        P2_REG0_REG_24__SCAN_IN), .B2(keyinput122), .ZN(n10392) );
  OAI221_X1 U11430 ( .B1(P2_REG1_REG_20__SCAN_IN), .B2(keyinput51), .C1(
        P2_REG0_REG_24__SCAN_IN), .C2(keyinput122), .A(n10392), .ZN(n10399) );
  AOI22_X1 U11431 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(keyinput40), .B1(
        P2_REG3_REG_4__SCAN_IN), .B2(keyinput32), .ZN(n10393) );
  OAI221_X1 U11432 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(keyinput40), .C1(
        P2_REG3_REG_4__SCAN_IN), .C2(keyinput32), .A(n10393), .ZN(n10398) );
  AOI22_X1 U11433 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(keyinput125), .B1(SI_23_), .B2(keyinput52), .ZN(n10394) );
  OAI221_X1 U11434 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(keyinput125), .C1(
        SI_23_), .C2(keyinput52), .A(n10394), .ZN(n10397) );
  AOI22_X1 U11435 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput93), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(keyinput23), .ZN(n10395) );
  OAI221_X1 U11436 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput93), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput23), .A(n10395), .ZN(n10396) );
  NOR4_X1 U11437 ( .A1(n10399), .A2(n10398), .A3(n10397), .A4(n10396), .ZN(
        n10418) );
  AOI22_X1 U11438 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(keyinput39), .B1(
        P2_IR_REG_7__SCAN_IN), .B2(keyinput113), .ZN(n10400) );
  OAI221_X1 U11439 ( .B1(P2_IR_REG_5__SCAN_IN), .B2(keyinput39), .C1(
        P2_IR_REG_7__SCAN_IN), .C2(keyinput113), .A(n10400), .ZN(n10407) );
  AOI22_X1 U11440 ( .A1(P1_REG0_REG_28__SCAN_IN), .A2(keyinput31), .B1(SI_10_), 
        .B2(keyinput19), .ZN(n10401) );
  OAI221_X1 U11441 ( .B1(P1_REG0_REG_28__SCAN_IN), .B2(keyinput31), .C1(SI_10_), .C2(keyinput19), .A(n10401), .ZN(n10406) );
  AOI22_X1 U11442 ( .A1(SI_30_), .A2(keyinput77), .B1(P1_REG3_REG_10__SCAN_IN), 
        .B2(keyinput6), .ZN(n10402) );
  OAI221_X1 U11443 ( .B1(SI_30_), .B2(keyinput77), .C1(P1_REG3_REG_10__SCAN_IN), .C2(keyinput6), .A(n10402), .ZN(n10405) );
  AOI22_X1 U11444 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(keyinput12), .B1(
        P2_D_REG_5__SCAN_IN), .B2(keyinput105), .ZN(n10403) );
  OAI221_X1 U11445 ( .B1(P1_DATAO_REG_18__SCAN_IN), .B2(keyinput12), .C1(
        P2_D_REG_5__SCAN_IN), .C2(keyinput105), .A(n10403), .ZN(n10404) );
  NOR4_X1 U11446 ( .A1(n10407), .A2(n10406), .A3(n10405), .A4(n10404), .ZN(
        n10417) );
  AOI22_X1 U11447 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(keyinput5), .B1(
        P2_IR_REG_14__SCAN_IN), .B2(keyinput70), .ZN(n10408) );
  OAI221_X1 U11448 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(keyinput5), .C1(
        P2_IR_REG_14__SCAN_IN), .C2(keyinput70), .A(n10408), .ZN(n10415) );
  AOI22_X1 U11449 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(keyinput45), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(keyinput8), .ZN(n10409) );
  OAI221_X1 U11450 ( .B1(P1_IR_REG_24__SCAN_IN), .B2(keyinput45), .C1(
        P1_DATAO_REG_5__SCAN_IN), .C2(keyinput8), .A(n10409), .ZN(n10414) );
  AOI22_X1 U11451 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput28), .B1(
        P2_D_REG_2__SCAN_IN), .B2(keyinput88), .ZN(n10410) );
  OAI221_X1 U11452 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput28), .C1(
        P2_D_REG_2__SCAN_IN), .C2(keyinput88), .A(n10410), .ZN(n10413) );
  AOI22_X1 U11453 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput71), .B1(
        P2_ADDR_REG_16__SCAN_IN), .B2(keyinput79), .ZN(n10411) );
  OAI221_X1 U11454 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput71), .C1(
        P2_ADDR_REG_16__SCAN_IN), .C2(keyinput79), .A(n10411), .ZN(n10412) );
  NOR4_X1 U11455 ( .A1(n10415), .A2(n10414), .A3(n10413), .A4(n10412), .ZN(
        n10416) );
  NAND4_X1 U11456 ( .A1(n10419), .A2(n10418), .A3(n10417), .A4(n10416), .ZN(
        n10457) );
  AOI22_X1 U11457 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput103), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(keyinput61), .ZN(n10420) );
  OAI221_X1 U11458 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput103), .C1(
        P1_DATAO_REG_23__SCAN_IN), .C2(keyinput61), .A(n10420), .ZN(n10427) );
  AOI22_X1 U11459 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(keyinput47), .B1(
        P2_REG2_REG_10__SCAN_IN), .B2(keyinput84), .ZN(n10421) );
  OAI221_X1 U11460 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(keyinput47), .C1(
        P2_REG2_REG_10__SCAN_IN), .C2(keyinput84), .A(n10421), .ZN(n10426) );
  AOI22_X1 U11461 ( .A1(P1_REG1_REG_28__SCAN_IN), .A2(keyinput49), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(keyinput97), .ZN(n10422) );
  OAI221_X1 U11462 ( .B1(P1_REG1_REG_28__SCAN_IN), .B2(keyinput49), .C1(
        P1_REG3_REG_3__SCAN_IN), .C2(keyinput97), .A(n10422), .ZN(n10425) );
  AOI22_X1 U11463 ( .A1(P1_REG0_REG_30__SCAN_IN), .A2(keyinput72), .B1(
        P2_REG3_REG_23__SCAN_IN), .B2(keyinput100), .ZN(n10423) );
  OAI221_X1 U11464 ( .B1(P1_REG0_REG_30__SCAN_IN), .B2(keyinput72), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput100), .A(n10423), .ZN(n10424) );
  NOR4_X1 U11465 ( .A1(n10427), .A2(n10426), .A3(n10425), .A4(n10424), .ZN(
        n10455) );
  AOI22_X1 U11466 ( .A1(P1_REG2_REG_1__SCAN_IN), .A2(keyinput66), .B1(
        P2_REG2_REG_12__SCAN_IN), .B2(keyinput17), .ZN(n10428) );
  OAI221_X1 U11467 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(keyinput66), .C1(
        P2_REG2_REG_12__SCAN_IN), .C2(keyinput17), .A(n10428), .ZN(n10435) );
  AOI22_X1 U11468 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(keyinput117), .B1(
        P1_REG0_REG_27__SCAN_IN), .B2(keyinput80), .ZN(n10429) );
  OAI221_X1 U11469 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(keyinput117), .C1(
        P1_REG0_REG_27__SCAN_IN), .C2(keyinput80), .A(n10429), .ZN(n10434) );
  AOI22_X1 U11470 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(keyinput67), .B1(SI_24_), 
        .B2(keyinput75), .ZN(n10430) );
  OAI221_X1 U11471 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(keyinput67), .C1(SI_24_), .C2(keyinput75), .A(n10430), .ZN(n10433) );
  AOI22_X1 U11472 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(keyinput35), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(keyinput78), .ZN(n10431) );
  OAI221_X1 U11473 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(keyinput35), .C1(
        P1_DATAO_REG_29__SCAN_IN), .C2(keyinput78), .A(n10431), .ZN(n10432) );
  NOR4_X1 U11474 ( .A1(n10435), .A2(n10434), .A3(n10433), .A4(n10432), .ZN(
        n10454) );
  AOI22_X1 U11475 ( .A1(P2_REG1_REG_31__SCAN_IN), .A2(keyinput120), .B1(
        P1_REG0_REG_5__SCAN_IN), .B2(keyinput110), .ZN(n10436) );
  OAI221_X1 U11476 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(keyinput120), .C1(
        P1_REG0_REG_5__SCAN_IN), .C2(keyinput110), .A(n10436), .ZN(n10443) );
  AOI22_X1 U11477 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(keyinput63), .B1(
        P2_IR_REG_2__SCAN_IN), .B2(keyinput58), .ZN(n10437) );
  OAI221_X1 U11478 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(keyinput63), .C1(
        P2_IR_REG_2__SCAN_IN), .C2(keyinput58), .A(n10437), .ZN(n10442) );
  AOI22_X1 U11479 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(keyinput0), .B1(
        P2_REG3_REG_7__SCAN_IN), .B2(keyinput24), .ZN(n10438) );
  OAI221_X1 U11480 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(keyinput0), .C1(
        P2_REG3_REG_7__SCAN_IN), .C2(keyinput24), .A(n10438), .ZN(n10441) );
  AOI22_X1 U11481 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(keyinput98), .B1(
        P2_REG0_REG_0__SCAN_IN), .B2(keyinput13), .ZN(n10439) );
  OAI221_X1 U11482 ( .B1(P1_REG3_REG_27__SCAN_IN), .B2(keyinput98), .C1(
        P2_REG0_REG_0__SCAN_IN), .C2(keyinput13), .A(n10439), .ZN(n10440) );
  NOR4_X1 U11483 ( .A1(n10443), .A2(n10442), .A3(n10441), .A4(n10440), .ZN(
        n10453) );
  AOI22_X1 U11484 ( .A1(P1_REG0_REG_2__SCAN_IN), .A2(keyinput27), .B1(
        P1_IR_REG_15__SCAN_IN), .B2(keyinput37), .ZN(n10444) );
  OAI221_X1 U11485 ( .B1(P1_REG0_REG_2__SCAN_IN), .B2(keyinput27), .C1(
        P1_IR_REG_15__SCAN_IN), .C2(keyinput37), .A(n10444), .ZN(n10451) );
  AOI22_X1 U11486 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(keyinput83), .B1(
        P2_IR_REG_8__SCAN_IN), .B2(keyinput46), .ZN(n10445) );
  OAI221_X1 U11487 ( .B1(P2_REG2_REG_28__SCAN_IN), .B2(keyinput83), .C1(
        P2_IR_REG_8__SCAN_IN), .C2(keyinput46), .A(n10445), .ZN(n10450) );
  AOI22_X1 U11488 ( .A1(P1_REG1_REG_14__SCAN_IN), .A2(keyinput41), .B1(
        P1_REG1_REG_18__SCAN_IN), .B2(keyinput109), .ZN(n10446) );
  OAI221_X1 U11489 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(keyinput41), .C1(
        P1_REG1_REG_18__SCAN_IN), .C2(keyinput109), .A(n10446), .ZN(n10449) );
  AOI22_X1 U11490 ( .A1(P1_REG1_REG_27__SCAN_IN), .A2(keyinput42), .B1(
        P1_D_REG_20__SCAN_IN), .B2(keyinput57), .ZN(n10447) );
  OAI221_X1 U11491 ( .B1(P1_REG1_REG_27__SCAN_IN), .B2(keyinput42), .C1(
        P1_D_REG_20__SCAN_IN), .C2(keyinput57), .A(n10447), .ZN(n10448) );
  NOR4_X1 U11492 ( .A1(n10451), .A2(n10450), .A3(n10449), .A4(n10448), .ZN(
        n10452) );
  NAND4_X1 U11493 ( .A1(n10455), .A2(n10454), .A3(n10453), .A4(n10452), .ZN(
        n10456) );
  NOR4_X1 U11494 ( .A1(n10459), .A2(n10458), .A3(n10457), .A4(n10456), .ZN(
        n10460) );
  OAI21_X1 U11495 ( .B1(n10462), .B2(n10461), .A(n10460), .ZN(n10468) );
  AOI22_X1 U11496 ( .A1(n10466), .A2(n10465), .B1(n10464), .B2(n10463), .ZN(
        n10467) );
  XNOR2_X1 U11497 ( .A(n10468), .B(n10467), .ZN(P2_U3463) );
  OAI21_X1 U11498 ( .B1(n10471), .B2(n10470), .A(n10469), .ZN(ADD_1068_U50) );
  OAI21_X1 U11499 ( .B1(n10474), .B2(n10473), .A(n10472), .ZN(ADD_1068_U51) );
  OAI21_X1 U11500 ( .B1(n10477), .B2(n10476), .A(n10475), .ZN(ADD_1068_U47) );
  OAI21_X1 U11501 ( .B1(n10480), .B2(n10479), .A(n10478), .ZN(ADD_1068_U49) );
  OAI21_X1 U11502 ( .B1(n10483), .B2(n10482), .A(n10481), .ZN(ADD_1068_U48) );
  AOI21_X1 U11503 ( .B1(n10486), .B2(n10485), .A(n10484), .ZN(ADD_1068_U54) );
  AOI21_X1 U11504 ( .B1(n10489), .B2(n10488), .A(n10487), .ZN(ADD_1068_U53) );
  OAI21_X1 U11505 ( .B1(n10492), .B2(n10491), .A(n10490), .ZN(ADD_1068_U52) );
  CLKBUF_X3 U5752 ( .A(n5985), .Z(n8975) );
  CLKBUF_X1 U7457 ( .A(n5740), .Z(n5695) );
endmodule

