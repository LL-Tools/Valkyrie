

module b21_C_AntiSAT_k_128_2 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072;

  AND4_X1 U4809 ( .A1(n4349), .A2(n4409), .A3(n4492), .A4(n4408), .ZN(n8031)
         );
  NAND2_X1 U4810 ( .A1(n5747), .A2(n5746), .ZN(n5791) );
  OR2_X1 U4811 ( .A1(n7434), .A2(n4861), .ZN(n8105) );
  INV_X1 U4812 ( .A(n9913), .ZN(n7444) );
  CLKBUF_X1 U4813 ( .A(n4937), .Z(n5460) );
  INV_X2 U4814 ( .A(n8043), .ZN(n5783) );
  NAND2_X2 U4815 ( .A1(n5509), .A2(n9136), .ZN(n6572) );
  INV_X1 U4816 ( .A(n5550), .ZN(n6571) );
  AOI21_X1 U4817 ( .B1(n4784), .B2(n8353), .A(n4782), .ZN(n4781) );
  OR2_X1 U4818 ( .A1(n8027), .A2(n7848), .ZN(n7975) );
  BUF_X1 U4819 ( .A(n5560), .Z(n4311) );
  AND2_X1 U4820 ( .A1(n9293), .A2(n9061), .ZN(n7775) );
  NOR2_X1 U4821 ( .A1(n8342), .A2(n4785), .ZN(n4784) );
  NAND2_X1 U4822 ( .A1(n7957), .A2(n7958), .ZN(n8342) );
  INV_X1 U4823 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5919) );
  INV_X1 U4824 ( .A(n8964), .ZN(n4931) );
  AND4_X1 U4825 ( .A1(n4965), .A2(n4964), .A3(n4963), .A4(n4962), .ZN(n9748)
         );
  AND2_X1 U4827 ( .A1(n6571), .A2(n5841), .ZN(n5625) );
  NAND2_X2 U4828 ( .A1(n4882), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4877) );
  OAI21_X2 U4829 ( .B1(n5118), .B2(n4341), .A(n4742), .ZN(n5172) );
  OAI21_X2 U4830 ( .B1(n8434), .B2(n8433), .A(n7940), .ZN(n8424) );
  OAI21_X2 U4831 ( .B1(n8454), .B2(n7821), .A(n7986), .ZN(n8434) );
  MUX2_X2 U4832 ( .A(n7623), .B(n7622), .S(n7704), .Z(n7645) );
  MUX2_X2 U4833 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4899), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n4902) );
  BUF_X4 U4834 ( .A(n7825), .Z(n4304) );
  NAND2_X1 U4835 ( .A1(n6501), .A2(n6103), .ZN(n7825) );
  XNOR2_X1 U4837 ( .A(n7434), .B(n4861), .ZN(n8107) );
  INV_X1 U4838 ( .A(n7182), .ZN(n7180) );
  OAI21_X1 U4839 ( .B1(n4444), .B2(n4443), .A(n4442), .ZN(n4441) );
  INV_X2 U4840 ( .A(n5625), .ZN(n5739) );
  NAND2_X1 U4841 ( .A1(n4932), .A2(n4931), .ZN(n7528) );
  AND4_X2 U4842 ( .A1(n4943), .A2(n4942), .A3(n4941), .A4(n4940), .ZN(n4956)
         );
  INV_X2 U4843 ( .A(n6476), .ZN(n9950) );
  NAND2_X2 U4844 ( .A1(n7864), .A2(n7863), .ZN(n6396) );
  INV_X1 U4845 ( .A(n6616), .ZN(n9942) );
  AND3_X1 U4846 ( .A1(n6136), .A2(n6137), .A3(n4345), .ZN(n9936) );
  NAND2_X1 U4847 ( .A1(n7331), .A2(n9385), .ZN(n5006) );
  NAND2_X1 U4848 ( .A1(n6501), .A2(n7501), .ZN(n6790) );
  NAND2_X2 U4849 ( .A1(n6264), .A2(n6052), .ZN(n6501) );
  CLKBUF_X2 U4850 ( .A(n4895), .Z(n7501) );
  AOI21_X1 U4851 ( .B1(n9303), .B2(n9720), .A(n4568), .ZN(n4567) );
  OR3_X1 U4852 ( .A1(n8024), .A2(n8023), .A3(n8022), .ZN(n4349) );
  AOI211_X1 U4853 ( .C1(n9489), .C2(n9122), .A(n9094), .B(n9093), .ZN(n9310)
         );
  NOR2_X1 U4854 ( .A1(n8535), .A2(n4368), .ZN(n4459) );
  NAND2_X1 U4855 ( .A1(n8906), .A2(n5683), .ZN(n8870) );
  INV_X1 U4856 ( .A(n7460), .ZN(n8084) );
  NAND2_X1 U4857 ( .A1(n9148), .A2(n4404), .ZN(n9152) );
  OAI211_X1 U4858 ( .C1(n8107), .C2(n7447), .A(n4343), .B(n4440), .ZN(n7460)
         );
  NAND2_X1 U4859 ( .A1(n8362), .A2(n8363), .ZN(n8361) );
  AND2_X1 U4860 ( .A1(n7506), .A2(n7505), .ZN(n9293) );
  NAND2_X1 U4861 ( .A1(n8328), .A2(n7961), .ZN(n8303) );
  NAND2_X1 U4862 ( .A1(n9165), .A2(n9166), .ZN(n9148) );
  NAND2_X1 U4863 ( .A1(n8123), .A2(n7429), .ZN(n7434) );
  NAND2_X1 U4864 ( .A1(n8125), .A2(n8124), .ZN(n8123) );
  OR2_X1 U4865 ( .A1(n8336), .A2(n8537), .ZN(n8318) );
  AND2_X1 U4866 ( .A1(n5748), .A2(n5749), .ZN(n5746) );
  NAND2_X1 U4867 ( .A1(n4430), .A2(n4652), .ZN(n8076) );
  NAND2_X1 U4868 ( .A1(n7797), .A2(n7796), .ZN(n8537) );
  NAND2_X1 U4869 ( .A1(n7770), .A2(n7554), .ZN(n9092) );
  NOR2_X1 U4870 ( .A1(n8239), .A2(n8238), .ZN(n8255) );
  XNOR2_X1 U4871 ( .A(n4754), .B(n8247), .ZN(n8239) );
  XNOR2_X1 U4872 ( .A(n5434), .B(n5433), .ZN(n8831) );
  NAND2_X1 U4873 ( .A1(n5422), .A2(n5421), .ZN(n5434) );
  NAND2_X1 U4874 ( .A1(n7449), .A2(n7448), .ZN(n8554) );
  INV_X1 U4875 ( .A(n9713), .ZN(n4612) );
  AOI21_X1 U4876 ( .B1(n9499), .B2(n5151), .A(n4327), .ZN(n4614) );
  AND2_X1 U4877 ( .A1(n4529), .A2(n4527), .ZN(n6757) );
  NAND2_X1 U4878 ( .A1(n7587), .A2(n5515), .ZN(n9769) );
  NAND2_X1 U4879 ( .A1(n5233), .A2(n5232), .ZN(n5256) );
  NAND2_X1 U4880 ( .A1(n4600), .A2(n6705), .ZN(n6758) );
  NAND2_X1 U4881 ( .A1(n5768), .A2(n5986), .ZN(n8997) );
  AND2_X1 U4882 ( .A1(n7729), .A2(n7757), .ZN(n7595) );
  AND2_X1 U4883 ( .A1(n7588), .A2(n7590), .ZN(n9747) );
  XNOR2_X1 U4884 ( .A(n4566), .B(n5060), .ZN(n6594) );
  INV_X2 U4885 ( .A(n9441), .ZN(n4305) );
  AND2_X1 U4886 ( .A1(n6514), .A2(n7868), .ZN(n4316) );
  NAND2_X1 U4887 ( .A1(n4741), .A2(n5054), .ZN(n4566) );
  NAND2_X1 U4888 ( .A1(n6576), .A2(n5511), .ZN(n7530) );
  NAND2_X1 U4889 ( .A1(n5531), .A2(n7786), .ZN(n9770) );
  NAND2_X1 U4890 ( .A1(n5052), .A2(n5051), .ZN(n4741) );
  INV_X1 U4891 ( .A(n5509), .ZN(n7788) );
  NOR2_X1 U4892 ( .A1(n5553), .A2(n6582), .ZN(n6577) );
  AND4_X1 U4893 ( .A1(n4985), .A2(n4984), .A3(n4983), .A4(n4982), .ZN(n9773)
         );
  CLKBUF_X1 U4894 ( .A(n5510), .Z(n7752) );
  NAND2_X1 U4895 ( .A1(n5016), .A2(n5015), .ZN(n5033) );
  NAND2_X1 U4896 ( .A1(n4884), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n4890) );
  AND2_X1 U4897 ( .A1(n5471), .A2(n5470), .ZN(n5510) );
  NAND2_X1 U4898 ( .A1(n4417), .A2(n4990), .ZN(n5012) );
  AND4_X1 U4899 ( .A1(n6056), .A2(n6055), .A3(n6054), .A4(n6053), .ZN(n6402)
         );
  INV_X2 U4900 ( .A(n7390), .ZN(n7798) );
  AND4_X1 U4901 ( .A1(n6120), .A2(n6119), .A3(n6118), .A4(n6117), .ZN(n6550)
         );
  CLKBUF_X3 U4902 ( .A(n5844), .Z(n4307) );
  AND4_X1 U4903 ( .A1(n6133), .A2(n6132), .A3(n6131), .A4(n6130), .ZN(n6611)
         );
  NAND2_X1 U4904 ( .A1(n4883), .A2(n4882), .ZN(n9385) );
  NAND2_X1 U4906 ( .A1(n5505), .A2(n5504), .ZN(n5841) );
  INV_X2 U4907 ( .A(n6790), .ZN(n7839) );
  NAND2_X1 U4908 ( .A1(n4418), .A2(n4970), .ZN(n4987) );
  XNOR2_X1 U4909 ( .A(n5475), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5504) );
  AND2_X2 U4910 ( .A1(n8824), .A2(n5978), .ZN(n7832) );
  XNOR2_X1 U4912 ( .A(n5483), .B(n5482), .ZN(n7126) );
  OR2_X1 U4913 ( .A1(n5089), .A2(n5088), .ZN(n5108) );
  OR2_X1 U4914 ( .A1(n5935), .A2(n5919), .ZN(n5937) );
  XNOR2_X1 U4915 ( .A(n4547), .B(n5938), .ZN(n6052) );
  OAI21_X1 U4916 ( .B1(n4922), .B2(n4801), .A(n4924), .ZN(n4945) );
  NOR2_X1 U4917 ( .A1(n5831), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n5935) );
  OAI21_X1 U4918 ( .B1(n5831), .B2(n4788), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n4547) );
  XNOR2_X1 U4919 ( .A(n4923), .B(SI_1_), .ZN(n4922) );
  NAND2_X1 U4920 ( .A1(n4906), .A2(n6061), .ZN(n4923) );
  CLKBUF_X1 U4921 ( .A(n5081), .Z(n5082) );
  NAND2_X2 U4922 ( .A1(n6103), .A2(P1_U3084), .ZN(n9397) );
  NOR2_X1 U4923 ( .A1(n4643), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4642) );
  OR2_X1 U4924 ( .A1(n4994), .A2(n4878), .ZN(n4951) );
  CLKBUF_X1 U4925 ( .A(n4920), .Z(n4994) );
  NOR2_X1 U4926 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4833) );
  INV_X1 U4927 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5468) );
  INV_X1 U4928 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6189) );
  INV_X1 U4929 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n8726) );
  INV_X1 U4930 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4876) );
  NOR2_X2 U4931 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4972) );
  INV_X1 U4932 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4891) );
  INV_X1 U4933 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5945) );
  NOR2_X1 U4934 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4778) );
  INV_X1 U4935 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5803) );
  INV_X1 U4936 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5944) );
  INV_X4 U4937 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NAND2_X1 U4938 ( .A1(n9179), .A2(n7673), .ZN(n9165) );
  NAND2_X1 U4939 ( .A1(n5553), .A2(n6565), .ZN(n6569) );
  AND2_X1 U4940 ( .A1(n5791), .A2(n4306), .ZN(n8060) );
  NOR2_X1 U4941 ( .A1(n5793), .A2(n5792), .ZN(n4306) );
  NOR2_X2 U4942 ( .A1(n5824), .A2(n5823), .ZN(n5828) );
  NAND2_X1 U4943 ( .A1(n5552), .A2(n5551), .ZN(n5988) );
  NAND2_X1 U4944 ( .A1(n5471), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5467) );
  AND2_X1 U4945 ( .A1(n4821), .A2(n4824), .ZN(n8916) );
  OAI22_X2 U4946 ( .A1(n7204), .A2(n5186), .B1(n9275), .B2(n8848), .ZN(n9271)
         );
  BUF_X4 U4947 ( .A(n5560), .Z(n4310) );
  OAI21_X2 U4948 ( .B1(n7180), .B2(n4342), .A(n4665), .ZN(n8095) );
  NOR4_X2 U4949 ( .A1(n7775), .A2(n7751), .A3(n7750), .A4(n7749), .ZN(n7754)
         );
  AND2_X2 U4950 ( .A1(n5841), .A2(n5550), .ZN(n5560) );
  AND2_X1 U4951 ( .A1(n4868), .A2(n4867), .ZN(n4845) );
  NAND2_X2 U4952 ( .A1(n8870), .A2(n5695), .ZN(n5709) );
  NOR2_X2 U4953 ( .A1(n5279), .A2(n4860), .ZN(n5283) );
  BUF_X1 U4954 ( .A(n5560), .Z(n4309) );
  INV_X1 U4955 ( .A(n4313), .ZN(n4312) );
  AND2_X1 U4956 ( .A1(n6571), .A2(n5841), .ZN(n4313) );
  NAND2_X1 U4957 ( .A1(n7934), .A2(n7989), .ZN(n4464) );
  OR2_X1 U4958 ( .A1(n8588), .A2(n8287), .ZN(n7989) );
  NAND2_X1 U4959 ( .A1(n5209), .A2(n5208), .ZN(n4608) );
  INV_X1 U4960 ( .A(n4626), .ZN(n4623) );
  AND2_X1 U4961 ( .A1(n8024), .A2(n6109), .ZN(n4495) );
  XNOR2_X1 U4962 ( .A(n5918), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U4963 ( .A1(n5922), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5918) );
  NAND2_X1 U4964 ( .A1(n7936), .A2(n4391), .ZN(n4483) );
  NOR2_X1 U4965 ( .A1(n7821), .A2(n7975), .ZN(n4484) );
  AND2_X1 U4966 ( .A1(n7937), .A2(n4482), .ZN(n4481) );
  AND2_X1 U4967 ( .A1(n7986), .A2(n7975), .ZN(n4482) );
  AOI21_X1 U4968 ( .B1(n4808), .B2(n4806), .A(n4805), .ZN(n4804) );
  INV_X1 U4969 ( .A(n7947), .ZN(n4805) );
  INV_X1 U4970 ( .A(n7943), .ZN(n4806) );
  AOI21_X1 U4971 ( .B1(n8371), .B2(n4491), .A(n7978), .ZN(n4490) );
  INV_X1 U4972 ( .A(n8985), .ZN(n4830) );
  INV_X1 U4973 ( .A(n4339), .ZN(n4836) );
  OR2_X1 U4974 ( .A1(n9302), .A2(n9090), .ZN(n7705) );
  INV_X1 U4975 ( .A(n5296), .ZN(n4718) );
  INV_X1 U4976 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5236) );
  INV_X1 U4977 ( .A(n8116), .ZN(n4653) );
  INV_X1 U4978 ( .A(n4403), .ZN(n7970) );
  INV_X1 U4979 ( .A(n8829), .ZN(n5978) );
  OR2_X1 U4980 ( .A1(n5913), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5947) );
  NAND2_X1 U4981 ( .A1(n8422), .A2(n8293), .ZN(n4456) );
  AOI21_X1 U4982 ( .B1(n4453), .B2(n4451), .A(n4450), .ZN(n4449) );
  INV_X1 U4983 ( .A(n4454), .ZN(n4451) );
  NAND2_X1 U4984 ( .A1(n9950), .A2(n8188), .ZN(n7868) );
  AND2_X1 U4985 ( .A1(n7921), .A2(n7239), .ZN(n4585) );
  INV_X1 U4986 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5950) );
  INV_X1 U4987 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5804) );
  INV_X1 U4988 ( .A(n9385), .ZN(n4886) );
  NAND2_X1 U4989 ( .A1(n7650), .A2(n7651), .ZN(n4564) );
  NAND2_X1 U4990 ( .A1(n4416), .A2(n4415), .ZN(n7092) );
  INV_X1 U4991 ( .A(n4340), .ZN(n4622) );
  AND2_X1 U4992 ( .A1(n6726), .A2(n9136), .ZN(n5751) );
  NAND2_X1 U4993 ( .A1(n5436), .A2(n5435), .ZN(n5451) );
  NAND2_X1 U4994 ( .A1(n5434), .A2(n5433), .ZN(n5436) );
  OAI21_X1 U4995 ( .B1(n5402), .B2(n5401), .A(n5400), .ZN(n5420) );
  INV_X1 U4996 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n4869) );
  AOI21_X1 U4997 ( .B1(n4729), .B2(n4337), .A(n4728), .ZN(n4727) );
  NOR2_X1 U4998 ( .A1(n5191), .A2(n4734), .ZN(n4733) );
  INV_X1 U4999 ( .A(n5173), .ZN(n4734) );
  INV_X1 U5000 ( .A(n4743), .ZN(n4742) );
  OAI21_X1 U5001 ( .B1(n4746), .B2(n4341), .A(n5152), .ZN(n4743) );
  INV_X1 U5002 ( .A(n7359), .ZN(n4436) );
  NAND2_X1 U5003 ( .A1(n8023), .A2(n8020), .ZN(n7845) );
  OR2_X1 U5004 ( .A1(n8567), .A2(n8293), .ZN(n8409) );
  OR2_X1 U5005 ( .A1(n8453), .A2(n8289), .ZN(n4856) );
  AOI21_X1 U5006 ( .B1(n4685), .B2(n4683), .A(n4371), .ZN(n4682) );
  INV_X1 U5007 ( .A(n8489), .ZN(n4683) );
  INV_X1 U5008 ( .A(n4685), .ZN(n4684) );
  AOI21_X1 U5009 ( .B1(n4712), .B2(n8001), .A(n4370), .ZN(n4457) );
  INV_X1 U5010 ( .A(n6501), .ZN(n7369) );
  INV_X1 U5011 ( .A(n4304), .ZN(n7370) );
  NAND2_X1 U5012 ( .A1(n7841), .A2(n7840), .ZN(n8522) );
  NOR2_X1 U5013 ( .A1(n4788), .A2(n4787), .ZN(n4786) );
  NAND2_X1 U5014 ( .A1(n5827), .A2(n5938), .ZN(n4787) );
  NAND2_X1 U5015 ( .A1(n5813), .A2(n4676), .ZN(n4674) );
  OR2_X1 U5016 ( .A1(n8917), .A2(n5731), .ZN(n4823) );
  CLKBUF_X3 U5017 ( .A(n4939), .Z(n7507) );
  AND2_X1 U5018 ( .A1(n4886), .A2(n7331), .ZN(n4939) );
  XNOR2_X1 U5019 ( .A(n9033), .B(n9045), .ZN(n9656) );
  NOR2_X1 U5020 ( .A1(n4510), .A2(n9307), .ZN(n4507) );
  NOR2_X1 U5021 ( .A1(n9512), .A2(n4509), .ZN(n4508) );
  OR2_X1 U5022 ( .A1(n4510), .A2(n9307), .ZN(n4509) );
  AND2_X1 U5023 ( .A1(n4631), .A2(n5418), .ZN(n4626) );
  NAND2_X1 U5024 ( .A1(n9313), .A2(n9122), .ZN(n4629) );
  AOI21_X1 U5025 ( .B1(n4323), .B2(n4606), .A(n4365), .ZN(n4602) );
  NAND2_X1 U5026 ( .A1(n5200), .A2(n5199), .ZN(n9286) );
  BUF_X1 U5027 ( .A(n5278), .Z(n7512) );
  AOI21_X1 U5028 ( .B1(n4612), .B2(n4329), .A(n4609), .ZN(n7078) );
  NAND2_X1 U5029 ( .A1(n4376), .A2(n4610), .ZN(n4609) );
  INV_X1 U5030 ( .A(n5278), .ZN(n5104) );
  INV_X1 U5031 ( .A(n4919), .ZN(n5844) );
  AND2_X1 U5032 ( .A1(n4919), .A2(n6103), .ZN(n5278) );
  NAND2_X1 U5033 ( .A1(n7726), .A2(n6577), .ZN(n6576) );
  NAND2_X2 U5034 ( .A1(n5532), .A2(n7492), .ZN(n4919) );
  INV_X1 U5035 ( .A(n9104), .ZN(n9313) );
  NAND2_X1 U5036 ( .A1(n4493), .A2(n4355), .ZN(n4492) );
  INV_X1 U5037 ( .A(n4495), .ZN(n4493) );
  AOI211_X1 U5038 ( .C1(n8264), .C2(n9892), .A(n9895), .B(n8481), .ZN(n4769)
         );
  NOR2_X1 U5039 ( .A1(n4318), .A2(n7990), .ZN(n4473) );
  NAND2_X1 U5040 ( .A1(n5518), .A2(n7595), .ZN(n7601) );
  NOR2_X1 U5041 ( .A1(n4477), .A2(n7888), .ZN(n4476) );
  INV_X1 U5042 ( .A(n7886), .ZN(n4477) );
  AND2_X1 U5043 ( .A1(n7989), .A2(n7929), .ZN(n4799) );
  NAND2_X1 U5044 ( .A1(n4479), .A2(n4328), .ZN(n4803) );
  AOI21_X1 U5045 ( .B1(n4804), .B2(n4807), .A(n4348), .ZN(n4802) );
  INV_X1 U5046 ( .A(n4808), .ZN(n4807) );
  NAND2_X1 U5047 ( .A1(n4490), .A2(n7950), .ZN(n4489) );
  AND2_X1 U5048 ( .A1(n8014), .A2(n7956), .ZN(n4814) );
  OR2_X1 U5049 ( .A1(n4379), .A2(n4816), .ZN(n4488) );
  INV_X1 U5050 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4714) );
  AND2_X1 U5051 ( .A1(n8109), .A2(n7433), .ZN(n4664) );
  NAND2_X1 U5052 ( .A1(n4546), .A2(n4545), .ZN(n4544) );
  INV_X1 U5053 ( .A(n4593), .ZN(n4591) );
  INV_X1 U5054 ( .A(n4781), .ZN(n4587) );
  INV_X1 U5055 ( .A(n4594), .ZN(n4588) );
  NAND2_X1 U5056 ( .A1(n8371), .A2(n7951), .ZN(n4593) );
  AND2_X1 U5057 ( .A1(n7951), .A2(n7947), .ZN(n4594) );
  NAND2_X1 U5058 ( .A1(n4449), .A2(n4452), .ZN(n4446) );
  OR2_X1 U5059 ( .A1(n8558), .A2(n8061), .ZN(n7947) );
  NOR2_X1 U5060 ( .A1(n8296), .A2(n4697), .ZN(n4693) );
  OR2_X1 U5061 ( .A1(n8554), .A2(n8173), .ZN(n7951) );
  OR2_X1 U5062 ( .A1(n7421), .A2(n8128), .ZN(n7435) );
  NOR2_X1 U5063 ( .A1(n8567), .A2(n8573), .ZN(n4539) );
  OR2_X1 U5064 ( .A1(n8578), .A2(n8289), .ZN(n7986) );
  OR2_X1 U5065 ( .A1(n8584), .A2(n8456), .ZN(n7988) );
  OR2_X1 U5066 ( .A1(n8594), .A2(n8098), .ZN(n7929) );
  NAND2_X1 U5067 ( .A1(n9458), .A2(n4535), .ZN(n4534) );
  NOR2_X1 U5068 ( .A1(n4531), .A2(n4528), .ZN(n4527) );
  NAND2_X1 U5069 ( .A1(n9966), .A2(n9956), .ZN(n4528) );
  OR2_X1 U5070 ( .A1(n8280), .A2(n8606), .ZN(n8281) );
  NAND2_X1 U5071 ( .A1(n4710), .A2(n8281), .ZN(n4709) );
  OR2_X1 U5072 ( .A1(n4531), .A2(n6477), .ZN(n4530) );
  NAND2_X1 U5073 ( .A1(n6033), .A2(n6032), .ZN(n8526) );
  NAND2_X1 U5074 ( .A1(n6382), .A2(n6381), .ZN(n8527) );
  NOR2_X1 U5075 ( .A1(n4827), .A2(n4830), .ZN(n4826) );
  INV_X1 U5076 ( .A(n5662), .ZN(n4827) );
  OR2_X1 U5077 ( .A1(n5657), .A2(n4830), .ZN(n4829) );
  INV_X1 U5078 ( .A(n4835), .ZN(n4834) );
  OAI21_X1 U5079 ( .B1(n4319), .B2(n4836), .A(n4372), .ZN(n4835) );
  XNOR2_X1 U5080 ( .A(n5568), .B(n5783), .ZN(n5569) );
  INV_X1 U5081 ( .A(n5660), .ZN(n4831) );
  NAND2_X1 U5082 ( .A1(n7778), .A2(n7581), .ZN(n7584) );
  AND2_X1 U5083 ( .A1(n7580), .A2(n7704), .ZN(n7581) );
  NOR2_X1 U5084 ( .A1(n4628), .A2(n4617), .ZN(n4616) );
  INV_X1 U5085 ( .A(n9121), .ZN(n4617) );
  NAND2_X1 U5086 ( .A1(n9071), .A2(n4622), .ZN(n4621) );
  INV_X1 U5087 ( .A(n7770), .ZN(n4554) );
  INV_X1 U5088 ( .A(n4557), .ZN(n4555) );
  OAI21_X1 U5089 ( .B1(n7566), .B2(n7694), .A(n7699), .ZN(n4559) );
  NOR2_X1 U5090 ( .A1(n9327), .A2(n9323), .ZN(n4503) );
  INV_X1 U5091 ( .A(n9173), .ZN(n5325) );
  NAND2_X1 U5092 ( .A1(n9520), .A2(n9532), .ZN(n4498) );
  NAND2_X1 U5093 ( .A1(n7788), .A2(n9745), .ZN(n7704) );
  OAI21_X1 U5094 ( .B1(n5383), .B2(n5382), .A(n5386), .ZN(n5402) );
  NAND2_X1 U5095 ( .A1(n5370), .A2(n5369), .ZN(n5383) );
  OAI21_X1 U5096 ( .B1(n5327), .B2(n4748), .A(n5331), .ZN(n5348) );
  INV_X1 U5097 ( .A(n5328), .ZN(n4748) );
  OR2_X1 U5098 ( .A1(n5469), .A2(n5468), .ZN(n5470) );
  NAND2_X1 U5099 ( .A1(n4715), .A2(n4716), .ZN(n5313) );
  AOI21_X1 U5100 ( .B1(n4317), .B2(n4724), .A(n4717), .ZN(n4716) );
  INV_X1 U5101 ( .A(n5295), .ZN(n4717) );
  AND2_X1 U5102 ( .A1(n5314), .A2(n5301), .ZN(n5312) );
  INV_X1 U5103 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5218) );
  INV_X1 U5104 ( .A(n5190), .ZN(n4731) );
  INV_X1 U5105 ( .A(n4730), .ZN(n4729) );
  OAI21_X1 U5106 ( .B1(n4733), .B2(n4337), .A(n5210), .ZN(n4730) );
  NOR2_X1 U5107 ( .A1(n5136), .A2(n4747), .ZN(n4746) );
  INV_X1 U5108 ( .A(n5117), .ZN(n4747) );
  NAND2_X1 U5109 ( .A1(n5116), .A2(n5115), .ZN(n5118) );
  NOR2_X1 U5110 ( .A1(n5073), .A2(n4740), .ZN(n4739) );
  INV_X1 U5111 ( .A(n5054), .ZN(n4740) );
  AND2_X1 U5112 ( .A1(n4994), .A2(n4865), .ZN(n4866) );
  OR2_X1 U5113 ( .A1(n8152), .A2(n7475), .ZN(n4427) );
  OR2_X1 U5114 ( .A1(n7153), .A2(n7152), .ZN(n7242) );
  INV_X1 U5115 ( .A(n6702), .ZN(n4444) );
  NOR2_X1 U5116 ( .A1(n7056), .A2(n4660), .ZN(n4442) );
  INV_X1 U5117 ( .A(n4662), .ZN(n4443) );
  XNOR2_X1 U5118 ( .A(n6973), .B(n7798), .ZN(n7003) );
  AND2_X1 U5119 ( .A1(n6423), .A2(n6422), .ZN(n4670) );
  OR2_X1 U5120 ( .A1(n7143), .A2(n5835), .ZN(n6259) );
  AND4_X1 U5121 ( .A1(n7248), .A2(n7247), .A3(n7246), .A4(n7245), .ZN(n8177)
         );
  OR2_X1 U5122 ( .A1(n6266), .A2(n6265), .ZN(n4752) );
  NOR2_X1 U5123 ( .A1(n5947), .A2(n5946), .ZN(n5951) );
  OR2_X1 U5124 ( .A1(n6732), .A2(n6731), .ZN(n4765) );
  INV_X1 U5125 ( .A(n4544), .ZN(n4543) );
  NAND2_X1 U5126 ( .A1(n7831), .A2(n7830), .ZN(n8276) );
  AND2_X1 U5127 ( .A1(n7342), .A2(n7341), .ZN(n8325) );
  OR2_X1 U5128 ( .A1(n7477), .A2(n7453), .ZN(n7342) );
  INV_X1 U5129 ( .A(n7955), .ZN(n4785) );
  NAND2_X1 U5130 ( .A1(n8361), .A2(n7955), .ZN(n8343) );
  OR2_X1 U5131 ( .A1(n8548), .A2(n8297), .ZN(n8298) );
  NAND2_X1 U5132 ( .A1(n4592), .A2(n4593), .ZN(n8362) );
  NAND2_X1 U5133 ( .A1(n8397), .A2(n4594), .ZN(n4592) );
  NAND2_X1 U5134 ( .A1(n8397), .A2(n7947), .ZN(n8376) );
  NAND2_X1 U5135 ( .A1(n8402), .A2(n4693), .ZN(n4689) );
  NAND2_X1 U5136 ( .A1(n4695), .A2(n8061), .ZN(n4694) );
  INV_X1 U5137 ( .A(n4691), .ZN(n4690) );
  OAI21_X1 U5138 ( .B1(n4693), .B2(n4692), .A(n8371), .ZN(n4691) );
  INV_X1 U5139 ( .A(n4694), .ZN(n4692) );
  NAND2_X1 U5140 ( .A1(n8439), .A2(n4330), .ZN(n8389) );
  AND2_X1 U5141 ( .A1(n4456), .A2(n8292), .ZN(n4454) );
  NAND2_X1 U5142 ( .A1(n4378), .A2(n4456), .ZN(n4453) );
  NAND2_X1 U5143 ( .A1(n4445), .A2(n4449), .ZN(n8402) );
  OR2_X1 U5144 ( .A1(n8432), .A2(n4452), .ZN(n4445) );
  AND3_X1 U5145 ( .A1(n7411), .A2(n7410), .A3(n7409), .ZN(n8458) );
  NAND2_X1 U5146 ( .A1(n4681), .A2(n4679), .ZN(n8447) );
  AOI21_X1 U5147 ( .B1(n4682), .B2(n4684), .A(n4680), .ZN(n4679) );
  AND2_X1 U5148 ( .A1(n4351), .A2(n8466), .ZN(n4685) );
  NAND2_X1 U5149 ( .A1(n8502), .A2(n8286), .ZN(n8488) );
  NAND2_X1 U5150 ( .A1(n8285), .A2(n8098), .ZN(n8286) );
  INV_X1 U5151 ( .A(n4585), .ZN(n4584) );
  AOI21_X1 U5152 ( .B1(n4585), .B2(n4583), .A(n4582), .ZN(n4581) );
  NAND2_X1 U5153 ( .A1(n4704), .A2(n4702), .ZN(n8502) );
  NOR2_X1 U5154 ( .A1(n4705), .A2(n4703), .ZN(n4702) );
  INV_X1 U5155 ( .A(n8514), .ZN(n4703) );
  NOR2_X1 U5156 ( .A1(n7235), .A2(n7234), .ZN(n8283) );
  AND2_X1 U5157 ( .A1(n7921), .A2(n8600), .ZN(n8282) );
  NAND2_X1 U5158 ( .A1(n7151), .A2(n8008), .ZN(n7240) );
  NAND2_X1 U5159 ( .A1(n4700), .A2(n4698), .ZN(n6946) );
  AND2_X1 U5160 ( .A1(n4699), .A2(n8004), .ZN(n4698) );
  NAND2_X1 U5161 ( .A1(n8000), .A2(n6843), .ZN(n4699) );
  OAI21_X1 U5162 ( .B1(n6859), .B2(n6860), .A(n4595), .ZN(n6956) );
  INV_X1 U5163 ( .A(n4596), .ZN(n4595) );
  OR2_X1 U5164 ( .A1(n6795), .A2(n8000), .ZN(n6844) );
  NOR2_X1 U5165 ( .A1(n7999), .A2(n4713), .ZN(n4712) );
  INV_X1 U5166 ( .A(n6748), .ZN(n4713) );
  AND2_X1 U5167 ( .A1(n6157), .A2(n6052), .ZN(n8603) );
  NAND2_X1 U5168 ( .A1(n6654), .A2(n7997), .ZN(n6636) );
  OR2_X1 U5169 ( .A1(n6638), .A2(n8001), .ZN(n6749) );
  NOR2_X1 U5170 ( .A1(n7996), .A2(n4773), .ZN(n4772) );
  NOR2_X1 U5171 ( .A1(n4316), .A2(n4776), .ZN(n4773) );
  NAND2_X1 U5172 ( .A1(n6545), .A2(n7857), .ZN(n6515) );
  AND4_X1 U5173 ( .A1(n6170), .A2(n6169), .A3(n6168), .A4(n6167), .ZN(n6467)
         );
  NAND2_X1 U5174 ( .A1(n7850), .A2(n7860), .ZN(n6400) );
  INV_X1 U5175 ( .A(n6109), .ZN(n8023) );
  INV_X1 U5176 ( .A(n8603), .ZN(n8457) );
  NOR2_X1 U5177 ( .A1(n4580), .A2(n9996), .ZN(n4460) );
  INV_X1 U5178 ( .A(n8536), .ZN(n4580) );
  NAND2_X1 U5179 ( .A1(n7274), .A2(n7273), .ZN(n8610) );
  INV_X1 U5180 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5936) );
  XNOR2_X1 U5181 ( .A(n5934), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8020) );
  NAND2_X1 U5182 ( .A1(n4649), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n4648) );
  NAND2_X1 U5183 ( .A1(n6047), .A2(n5919), .ZN(n4647) );
  NOR2_X1 U5184 ( .A1(n6047), .A2(n5919), .ZN(n4649) );
  AND2_X1 U5185 ( .A1(n5812), .A2(n4780), .ZN(n4779) );
  AND2_X1 U5186 ( .A1(n5911), .A2(n5928), .ZN(n6792) );
  NAND2_X1 U5187 ( .A1(n5709), .A2(n4319), .ZN(n4838) );
  NAND2_X1 U5188 ( .A1(n4842), .A2(n4840), .ZN(n7037) );
  NOR2_X1 U5189 ( .A1(n7039), .A2(n4841), .ZN(n4840) );
  INV_X1 U5190 ( .A(n4843), .ZN(n4841) );
  AND2_X1 U5191 ( .A1(n5642), .A2(n5641), .ZN(n8935) );
  OR2_X1 U5192 ( .A1(n7756), .A2(n5751), .ZN(n6088) );
  NAND2_X1 U5193 ( .A1(n5480), .A2(n4846), .ZN(n4901) );
  AND2_X1 U5194 ( .A1(n4848), .A2(n4847), .ZN(n4846) );
  INV_X1 U5195 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4847) );
  AND3_X1 U5196 ( .A1(n5399), .A2(n5398), .A3(n5397), .ZN(n5733) );
  NOR2_X1 U5197 ( .A1(n9642), .A2(n9032), .ZN(n9033) );
  OR2_X1 U5198 ( .A1(n9656), .A2(n9655), .ZN(n4518) );
  AND2_X1 U5199 ( .A1(n5442), .A2(n5459), .ZN(n9075) );
  OR2_X1 U5200 ( .A1(n9317), .A2(n5733), .ZN(n9105) );
  NAND2_X1 U5201 ( .A1(n9119), .A2(n5733), .ZN(n4631) );
  AND2_X1 U5202 ( .A1(n9161), .A2(n4501), .ZN(n9116) );
  NOR2_X1 U5203 ( .A1(n4502), .A2(n9317), .ZN(n4501) );
  INV_X1 U5204 ( .A(n4503), .ZN(n4502) );
  AND2_X1 U5205 ( .A1(n7746), .A2(n7675), .ZN(n4404) );
  OR2_X1 U5206 ( .A1(n9332), .A2(n9182), .ZN(n5344) );
  NOR2_X1 U5207 ( .A1(n9186), .A2(n9332), .ZN(n9161) );
  AND2_X1 U5208 ( .A1(n7672), .A2(n7673), .ZN(n9173) );
  AOI21_X1 U5209 ( .B1(n5294), .B2(n4637), .A(n4359), .ZN(n4636) );
  INV_X1 U5210 ( .A(n5269), .ZN(n4637) );
  OR2_X1 U5211 ( .A1(n7722), .A2(n7721), .ZN(n9199) );
  NAND2_X1 U5212 ( .A1(n4563), .A2(n4561), .ZN(n9214) );
  AOI21_X1 U5213 ( .B1(n7657), .B2(n4564), .A(n4562), .ZN(n4561) );
  INV_X1 U5214 ( .A(n7665), .ZN(n4562) );
  NOR2_X1 U5215 ( .A1(n4315), .A2(n9359), .ZN(n9243) );
  AND2_X1 U5216 ( .A1(n9225), .A2(n7650), .ZN(n9247) );
  AOI21_X1 U5217 ( .B1(n4320), .B2(n4605), .A(n4362), .ZN(n4604) );
  INV_X1 U5218 ( .A(n5208), .ZN(n4605) );
  INV_X1 U5219 ( .A(n4320), .ZN(n4606) );
  NAND2_X1 U5220 ( .A1(n5178), .A2(n5177), .ZN(n8848) );
  NAND2_X1 U5221 ( .A1(n5522), .A2(n4332), .ZN(n7207) );
  AND2_X1 U5222 ( .A1(n7609), .A2(n7626), .ZN(n7733) );
  AND2_X1 U5223 ( .A1(n9714), .A2(n7602), .ZN(n4548) );
  OR2_X1 U5224 ( .A1(n9759), .A2(n9758), .ZN(n9761) );
  NOR2_X1 U5225 ( .A1(n7524), .A2(n6565), .ZN(n6671) );
  NAND2_X1 U5226 ( .A1(n7514), .A2(n7513), .ZN(n9512) );
  INV_X1 U5227 ( .A(n4618), .ZN(n9072) );
  AOI22_X1 U5228 ( .A1(n4632), .A2(n4619), .B1(n4628), .B2(n4622), .ZN(n4618)
         );
  NOR2_X1 U5229 ( .A1(n4340), .A2(n4623), .ZN(n4619) );
  AND3_X1 U5230 ( .A1(n5086), .A2(n5085), .A3(n5084), .ZN(n9850) );
  AND2_X1 U5231 ( .A1(n6093), .A2(n5752), .ZN(n9827) );
  OR2_X1 U5232 ( .A1(n7704), .A2(n7783), .ZN(n9832) );
  INV_X1 U5233 ( .A(n9828), .ZN(n9851) );
  INV_X1 U5234 ( .A(n7524), .ZN(n9795) );
  XNOR2_X1 U5235 ( .A(n7504), .B(n7503), .ZN(n8818) );
  NAND2_X1 U5236 ( .A1(n5479), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5475) );
  XNOR2_X1 U5237 ( .A(n5507), .B(n5506), .ZN(n6985) );
  OR2_X1 U5238 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n4860) );
  NAND2_X1 U5239 ( .A1(n4719), .A2(n4721), .ZN(n5297) );
  NAND2_X1 U5240 ( .A1(n4720), .A2(n4723), .ZN(n4719) );
  INV_X1 U5241 ( .A(n5256), .ZN(n4720) );
  NAND2_X1 U5242 ( .A1(n4732), .A2(n5190), .ZN(n5212) );
  NAND2_X1 U5243 ( .A1(n5174), .A2(n4733), .ZN(n4732) );
  OAI21_X2 U5244 ( .B1(n5052), .B2(n4738), .A(n4735), .ZN(n5116) );
  NAND2_X1 U5245 ( .A1(n4858), .A2(n4739), .ZN(n4738) );
  INV_X1 U5246 ( .A(n4736), .ZN(n4735) );
  OAI21_X1 U5247 ( .B1(n4737), .B2(n4813), .A(n4810), .ZN(n4736) );
  INV_X1 U5248 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4864) );
  INV_X1 U5249 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4865) );
  INV_X1 U5250 ( .A(n4921), .ZN(n4801) );
  AOI21_X1 U5251 ( .B1(n4425), .B2(n7475), .A(n4422), .ZN(n4421) );
  OAI21_X1 U5252 ( .B1(n7476), .B2(n4423), .A(n8150), .ZN(n4422) );
  OR2_X1 U5253 ( .A1(n8152), .A2(n7475), .ZN(n4423) );
  OR2_X1 U5254 ( .A1(n7476), .A2(n7475), .ZN(n4424) );
  NAND2_X1 U5255 ( .A1(n8542), .A2(n9886), .ZN(n4429) );
  NAND2_X1 U5256 ( .A1(n7173), .A2(n7172), .ZN(n7178) );
  INV_X1 U5257 ( .A(n8584), .ZN(n8288) );
  AND4_X1 U5258 ( .A1(n7298), .A2(n7297), .A3(n7296), .A4(n7295), .ZN(n8287)
         );
  OR2_X1 U5259 ( .A1(n6790), .A2(n6105), .ZN(n6106) );
  AOI21_X1 U5260 ( .B1(n4375), .B2(n4654), .A(n4331), .ZN(n4652) );
  AND2_X1 U5261 ( .A1(n7469), .A2(n7468), .ZN(n8358) );
  NAND2_X1 U5262 ( .A1(n8084), .A2(n7461), .ZN(n4650) );
  NAND2_X1 U5263 ( .A1(n7463), .A2(n7462), .ZN(n4651) );
  NAND2_X1 U5264 ( .A1(n4495), .A2(n4494), .ZN(n4408) );
  NOR2_X1 U5265 ( .A1(n7982), .A2(n9913), .ZN(n4494) );
  OR2_X1 U5266 ( .A1(n6385), .A2(n6052), .ZN(n8455) );
  INV_X1 U5267 ( .A(n8458), .ZN(n8291) );
  AND2_X1 U5268 ( .A1(n4765), .A2(n4764), .ZN(n7019) );
  NAND2_X1 U5269 ( .A1(n6941), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4764) );
  INV_X1 U5270 ( .A(n4754), .ZN(n8253) );
  NAND2_X1 U5271 ( .A1(n4579), .A2(n4577), .ZN(n8535) );
  INV_X1 U5272 ( .A(n4578), .ZN(n4577) );
  NAND2_X1 U5273 ( .A1(n4321), .A2(n8608), .ZN(n4579) );
  OAI22_X1 U5274 ( .A1(n8345), .A2(n8455), .B1(n8306), .B2(n8305), .ZN(n4578)
         );
  OR2_X1 U5275 ( .A1(n9904), .A2(n8525), .ZN(n8437) );
  AND2_X1 U5276 ( .A1(n7143), .A2(n8836), .ZN(n9908) );
  INV_X1 U5277 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U5278 ( .A1(n6048), .A2(n6046), .ZN(n6050) );
  OAI21_X1 U5279 ( .B1(n6594), .B2(n5104), .A(n4565), .ZN(n6826) );
  NOR2_X1 U5280 ( .A1(n4353), .A2(n4325), .ZN(n4565) );
  NOR2_X1 U5281 ( .A1(n6726), .A2(n4414), .ZN(n4413) );
  INV_X1 U5282 ( .A(n7784), .ZN(n4414) );
  OR2_X1 U5283 ( .A1(n7792), .A2(n4412), .ZN(n4411) );
  AND2_X1 U5284 ( .A1(n7785), .A2(n6726), .ZN(n4412) );
  MUX2_X1 U5285 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4903), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n4904) );
  INV_X1 U5286 ( .A(n5635), .ZN(n9004) );
  NAND2_X1 U5287 ( .A1(n4937), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4888) );
  AOI21_X1 U5288 ( .B1(n5541), .B2(n9770), .A(n5540), .ZN(n9300) );
  INV_X1 U5289 ( .A(n5539), .ZN(n5540) );
  XNOR2_X1 U5290 ( .A(n5530), .B(n5529), .ZN(n5541) );
  AOI22_X1 U5291 ( .A1(n9002), .A2(n9489), .B1(n9060), .B2(n9001), .ZN(n5539)
         );
  AOI21_X1 U5292 ( .B1(n9298), .B2(n9720), .A(n5545), .ZN(n5546) );
  XNOR2_X1 U5293 ( .A(n5464), .B(n7750), .ZN(n9301) );
  OR2_X1 U5294 ( .A1(n9306), .A2(n9290), .ZN(n4570) );
  AOI21_X1 U5295 ( .B1(n9081), .B2(n9770), .A(n4571), .ZN(n9305) );
  NAND2_X1 U5296 ( .A1(n4573), .A2(n4572), .ZN(n4571) );
  NAND2_X1 U5297 ( .A1(n9080), .A2(n9742), .ZN(n4573) );
  AND2_X1 U5298 ( .A1(n5409), .A2(n5408), .ZN(n9104) );
  NAND2_X1 U5299 ( .A1(n9779), .A2(n9740), .ZN(n9765) );
  OR3_X1 U5300 ( .A1(n9832), .A2(n7752), .A3(n9791), .ZN(n9283) );
  AND2_X1 U5301 ( .A1(n9235), .A2(n9828), .ZN(n9720) );
  INV_X1 U5302 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4878) );
  AOI21_X1 U5303 ( .B1(n4469), .B2(n4467), .A(n7867), .ZN(n7879) );
  NAND2_X1 U5304 ( .A1(n4818), .A2(n4361), .ZN(n4474) );
  NAND2_X1 U5305 ( .A1(n4478), .A2(n4476), .ZN(n4475) );
  MUX2_X1 U5306 ( .A(n7608), .B(n7607), .S(n7704), .Z(n7628) );
  NAND2_X1 U5307 ( .A1(n4800), .A2(n7978), .ZN(n4465) );
  NAND2_X1 U5308 ( .A1(n7930), .A2(n4799), .ZN(n4798) );
  MUX2_X1 U5309 ( .A(n7671), .B(n7670), .S(n7704), .Z(n7680) );
  AOI21_X1 U5310 ( .B1(n7943), .B2(n7944), .A(n4809), .ZN(n4808) );
  OR2_X1 U5311 ( .A1(n7951), .A2(n7975), .ZN(n4817) );
  AOI21_X1 U5312 ( .B1(n4487), .B2(n7966), .A(n4335), .ZN(n4485) );
  NAND2_X1 U5313 ( .A1(n4377), .A2(n7966), .ZN(n4486) );
  NAND2_X1 U5314 ( .A1(n4803), .A2(n4802), .ZN(n7953) );
  AND2_X1 U5315 ( .A1(n6528), .A2(n6473), .ZN(n6470) );
  NAND2_X1 U5316 ( .A1(n9960), .A2(n9950), .ZN(n4531) );
  AOI21_X1 U5317 ( .B1(n7701), .B2(n7700), .A(n9092), .ZN(n7709) );
  OAI21_X1 U5318 ( .B1(n7327), .B2(n7326), .A(n7330), .ZN(n7498) );
  INV_X1 U5319 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5235) );
  INV_X1 U5320 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5234) );
  INV_X1 U5321 ( .A(n5230), .ZN(n4728) );
  INV_X1 U5322 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5213) );
  INV_X1 U5323 ( .A(SI_15_), .ZN(n5193) );
  INV_X1 U5324 ( .A(n5140), .ZN(n4744) );
  NAND2_X1 U5325 ( .A1(n6977), .A2(n4439), .ZN(n7050) );
  INV_X1 U5326 ( .A(n6990), .ZN(n4439) );
  NAND2_X1 U5327 ( .A1(n4793), .A2(n7837), .ZN(n4792) );
  INV_X1 U5328 ( .A(n7973), .ZN(n4793) );
  NAND2_X1 U5329 ( .A1(n4792), .A2(n4794), .ZN(n4791) );
  AND2_X1 U5330 ( .A1(n8276), .A2(n4795), .ZN(n4794) );
  INV_X1 U5331 ( .A(n7837), .ZN(n4795) );
  INV_X1 U5332 ( .A(n8017), .ZN(n7984) );
  OAI21_X1 U5333 ( .B1(n8522), .B2(n8272), .A(n7971), .ZN(n8017) );
  OR2_X1 U5334 ( .A1(n7479), .A2(n7478), .ZN(n7481) );
  OR2_X1 U5335 ( .A1(n8537), .A2(n8345), .ZN(n7961) );
  NOR2_X1 U5336 ( .A1(n8562), .A2(n4538), .ZN(n4537) );
  INV_X1 U5337 ( .A(n4539), .ZN(n4538) );
  INV_X1 U5338 ( .A(n4453), .ZN(n4452) );
  INV_X1 U5339 ( .A(n8008), .ZN(n4583) );
  INV_X1 U5340 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7152) );
  INV_X1 U5341 ( .A(n7858), .ZN(n4776) );
  AOI21_X1 U5342 ( .B1(n4316), .B2(n4777), .A(n4776), .ZN(n4775) );
  AND2_X1 U5343 ( .A1(n6524), .A2(n6468), .ZN(n6469) );
  AND2_X1 U5344 ( .A1(n6526), .A2(n6470), .ZN(n6468) );
  NOR2_X1 U5345 ( .A1(n9929), .A2(n9920), .ZN(n4536) );
  INV_X1 U5346 ( .A(SI_25_), .ZN(n8779) );
  NOR2_X1 U5347 ( .A1(n8283), .A2(n8282), .ZN(n4711) );
  NAND2_X1 U5348 ( .A1(n6534), .A2(n6446), .ZN(n6444) );
  NAND2_X1 U5349 ( .A1(n5816), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U5350 ( .A1(n5933), .A2(n5815), .ZN(n5816) );
  INV_X1 U5351 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U5352 ( .A1(n4673), .A2(n5814), .ZN(n4672) );
  NOR2_X1 U5353 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5814) );
  INV_X1 U5354 ( .A(n4675), .ZN(n4673) );
  INV_X1 U5355 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4676) );
  INV_X1 U5356 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5813) );
  INV_X1 U5357 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5805) );
  INV_X1 U5358 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5806) );
  INV_X1 U5359 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5807) );
  NOR2_X1 U5360 ( .A1(n4849), .A2(n4326), .ZN(n4848) );
  NAND2_X1 U5361 ( .A1(n4850), .A2(n5482), .ZN(n4849) );
  INV_X1 U5362 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4850) );
  NAND2_X1 U5363 ( .A1(n5466), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5469) );
  NOR2_X1 U5364 ( .A1(n9629), .A2(n4522), .ZN(n9031) );
  AND2_X1 U5365 ( .A1(n9634), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4522) );
  NAND2_X1 U5366 ( .A1(n4512), .A2(n4511), .ZN(n4510) );
  AND2_X1 U5367 ( .A1(n7686), .A2(n7545), .ZN(n7746) );
  NOR2_X1 U5368 ( .A1(n9350), .A2(n9356), .ZN(n4514) );
  INV_X1 U5369 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5088) );
  NAND2_X1 U5370 ( .A1(n4611), .A2(n5087), .ZN(n4610) );
  INV_X1 U5371 ( .A(n5065), .ZN(n4611) );
  INV_X1 U5372 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U5373 ( .A1(n5519), .A2(n5518), .ZN(n6916) );
  NAND2_X1 U5374 ( .A1(n5509), .A2(n7752), .ZN(n7756) );
  NAND2_X1 U5375 ( .A1(n6909), .A2(n9821), .ZN(n4506) );
  XNOR2_X1 U5376 ( .A(n7498), .B(n7497), .ZN(n7495) );
  AND2_X1 U5377 ( .A1(n5435), .A2(n5427), .ZN(n5433) );
  AND2_X1 U5378 ( .A1(n5421), .A2(n5406), .ZN(n5419) );
  INV_X1 U5379 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4644) );
  NAND2_X1 U5380 ( .A1(n5315), .A2(n5314), .ZN(n5327) );
  AOI21_X1 U5381 ( .B1(n4723), .B2(n4722), .A(n4394), .ZN(n4721) );
  INV_X1 U5382 ( .A(n5254), .ZN(n4722) );
  INV_X1 U5383 ( .A(SI_13_), .ZN(n5156) );
  NAND2_X1 U5384 ( .A1(n4739), .A2(n5050), .ZN(n4737) );
  AOI21_X1 U5385 ( .B1(n4858), .B2(n4812), .A(n4811), .ZN(n4810) );
  INV_X1 U5386 ( .A(n5096), .ZN(n4811) );
  INV_X1 U5387 ( .A(n5074), .ZN(n4812) );
  OAI21_X1 U5388 ( .B1(n6103), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n4926), .ZN(
        n4946) );
  NAND2_X1 U5389 ( .A1(n6103), .A2(n4925), .ZN(n4926) );
  INV_X1 U5390 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4892) );
  NAND2_X1 U5391 ( .A1(n7180), .A2(n7179), .ZN(n7270) );
  AND2_X1 U5392 ( .A1(n4380), .A2(n4434), .ZN(n4433) );
  NAND2_X1 U5393 ( .A1(n4435), .A2(n7359), .ZN(n4434) );
  INV_X1 U5394 ( .A(n4437), .ZN(n4435) );
  OR2_X1 U5395 ( .A1(n8109), .A2(n7433), .ZN(n4440) );
  AOI21_X1 U5396 ( .B1(n4657), .B2(n4656), .A(n4655), .ZN(n4654) );
  INV_X1 U5397 ( .A(n7385), .ZN(n4655) );
  INV_X1 U5398 ( .A(n8141), .ZN(n4656) );
  INV_X1 U5399 ( .A(n6977), .ZN(n6975) );
  NOR2_X1 U5400 ( .A1(n7360), .A2(n4438), .ZN(n4437) );
  INV_X1 U5401 ( .A(n7282), .ZN(n4438) );
  INV_X1 U5402 ( .A(n4666), .ZN(n4665) );
  OAI21_X1 U5403 ( .B1(n7179), .B2(n4342), .A(n7278), .ZN(n4666) );
  INV_X1 U5404 ( .A(n7293), .ZN(n5971) );
  OR2_X1 U5405 ( .A1(n6417), .A2(n6416), .ZN(n4671) );
  OR2_X1 U5406 ( .A1(n7467), .A2(n7466), .ZN(n7469) );
  OR2_X1 U5407 ( .A1(n9904), .A2(n6157), .ZN(n6262) );
  OAI21_X1 U5408 ( .B1(n4338), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5933) );
  AND3_X1 U5409 ( .A1(n7425), .A2(n7424), .A3(n7423), .ZN(n8293) );
  AND4_X1 U5410 ( .A1(n7397), .A2(n7396), .A3(n7395), .A4(n7394), .ZN(n8289)
         );
  AND4_X1 U5411 ( .A1(n6148), .A2(n6147), .A3(n6146), .A4(n6145), .ZN(n6548)
         );
  NOR3_X1 U5412 ( .A1(n9901), .A2(n9896), .A3(n9404), .ZN(n9403) );
  NOR2_X1 U5413 ( .A1(n9417), .A2(n9416), .ZN(n9415) );
  NAND2_X1 U5414 ( .A1(n4752), .A2(n4751), .ZN(n4750) );
  NAND2_X1 U5415 ( .A1(n6283), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4751) );
  NAND2_X1 U5416 ( .A1(n4407), .A2(n4406), .ZN(n4760) );
  INV_X1 U5417 ( .A(n6300), .ZN(n4406) );
  INV_X1 U5418 ( .A(n6301), .ZN(n4407) );
  OR2_X1 U5419 ( .A1(n6317), .A2(n6316), .ZN(n4758) );
  NOR2_X1 U5420 ( .A1(n6729), .A2(n4766), .ZN(n8194) );
  AND2_X1 U5421 ( .A1(n6792), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4766) );
  NAND2_X1 U5422 ( .A1(n8194), .A2(n8195), .ZN(n8193) );
  OR2_X1 U5423 ( .A1(n5959), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n5960) );
  OR2_X1 U5424 ( .A1(n8223), .A2(n8222), .ZN(n4756) );
  NAND2_X1 U5425 ( .A1(n4756), .A2(n4755), .ZN(n4754) );
  NAND2_X1 U5426 ( .A1(n8240), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4755) );
  INV_X1 U5427 ( .A(n4590), .ZN(n4589) );
  AOI21_X1 U5428 ( .B1(n4590), .B2(n4588), .A(n4587), .ZN(n4586) );
  NOR2_X1 U5429 ( .A1(n4591), .A2(n4783), .ZN(n4590) );
  NAND2_X1 U5430 ( .A1(n7961), .A2(n7959), .ZN(n8323) );
  OR2_X1 U5431 ( .A1(n8542), .A2(n8364), .ZN(n8299) );
  NAND2_X1 U5432 ( .A1(n4688), .A2(n4687), .ZN(n8354) );
  AOI21_X1 U5433 ( .B1(n4690), .B2(n4692), .A(n4367), .ZN(n4687) );
  NAND2_X1 U5434 ( .A1(n4447), .A2(n4360), .ZN(n4688) );
  NAND2_X1 U5435 ( .A1(n4597), .A2(n4598), .ZN(n8395) );
  AOI21_X1 U5436 ( .B1(n7823), .B2(n8423), .A(n4599), .ZN(n4598) );
  INV_X1 U5437 ( .A(n7945), .ZN(n4599) );
  NAND2_X1 U5438 ( .A1(n8439), .A2(n4537), .ZN(n8404) );
  OR2_X1 U5439 ( .A1(n8424), .A2(n8423), .ZN(n8427) );
  NAND2_X1 U5440 ( .A1(n8439), .A2(n8290), .ZN(n8441) );
  NAND2_X1 U5441 ( .A1(n8508), .A2(n7816), .ZN(n8510) );
  NAND2_X1 U5442 ( .A1(n8283), .A2(n4707), .ZN(n4704) );
  INV_X1 U5443 ( .A(n4709), .ZN(n4707) );
  OAI21_X1 U5444 ( .B1(n4709), .B2(n4706), .A(n4393), .ZN(n4705) );
  INV_X1 U5445 ( .A(n8282), .ZN(n4706) );
  OR2_X1 U5446 ( .A1(n4534), .A2(n8610), .ZN(n4533) );
  OR2_X1 U5447 ( .A1(n4535), .A2(n8179), .ZN(n4863) );
  NOR2_X1 U5448 ( .A1(n7148), .A2(n8008), .ZN(n7235) );
  NOR3_X1 U5449 ( .A1(n7117), .A2(n7913), .A3(n7116), .ZN(n7252) );
  NOR2_X1 U5450 ( .A1(n7117), .A2(n7116), .ZN(n7162) );
  AND4_X1 U5451 ( .A1(n6855), .A2(n6854), .A3(n6853), .A4(n6852), .ZN(n7112)
         );
  CLKBUF_X1 U5452 ( .A(n6860), .Z(n6752) );
  OR2_X1 U5453 ( .A1(n6474), .A2(n7995), .ZN(n6631) );
  NOR2_X1 U5454 ( .A1(n6613), .A2(n6476), .ZN(n6646) );
  AND2_X1 U5455 ( .A1(n4536), .A2(n6534), .ZN(n6554) );
  INV_X1 U5456 ( .A(n6396), .ZN(n6397) );
  NAND2_X1 U5457 ( .A1(n6535), .A2(n7862), .ZN(n7850) );
  NAND2_X1 U5458 ( .A1(n8038), .A2(n9914), .ZN(n6535) );
  NAND2_X1 U5459 ( .A1(n7465), .A2(n7464), .ZN(n8548) );
  NAND2_X1 U5460 ( .A1(n7420), .A2(n7419), .ZN(n8567) );
  NAND2_X1 U5461 ( .A1(n7364), .A2(n7363), .ZN(n8588) );
  NOR2_X1 U5462 ( .A1(n4711), .A2(n4709), .ZN(n9446) );
  NAND2_X1 U5463 ( .A1(n7240), .A2(n4585), .ZN(n8601) );
  NOR3_X1 U5464 ( .A1(n6477), .A2(n6613), .A3(n6476), .ZN(n6660) );
  OR2_X1 U5465 ( .A1(n7444), .A2(n6159), .ZN(n9994) );
  INV_X1 U5466 ( .A(n9994), .ZN(n9930) );
  INV_X1 U5467 ( .A(n8529), .ZN(n8613) );
  NOR2_X1 U5468 ( .A1(n8528), .A2(n8527), .ZN(n8614) );
  AND2_X1 U5469 ( .A1(n6031), .A2(n6030), .ZN(n9903) );
  NAND2_X1 U5470 ( .A1(n6259), .A2(n9912), .ZN(n9904) );
  NAND2_X1 U5471 ( .A1(n4789), .A2(n5936), .ZN(n4788) );
  INV_X1 U5472 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4789) );
  NAND2_X1 U5473 ( .A1(n5837), .A2(n5836), .ZN(n5839) );
  NOR2_X1 U5474 ( .A1(n5824), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n6200) );
  AND2_X1 U5475 ( .A1(n5893), .A2(n5804), .ZN(n5900) );
  AND2_X1 U5476 ( .A1(n5895), .A2(n5894), .ZN(n6304) );
  INV_X2 U5477 ( .A(n8045), .ZN(n5785) );
  INV_X1 U5478 ( .A(n8878), .ZN(n4837) );
  NAND2_X1 U5479 ( .A1(n5710), .A2(n8923), .ZN(n4839) );
  NAND2_X1 U5480 ( .A1(n4825), .A2(n4352), .ZN(n8895) );
  NAND2_X1 U5481 ( .A1(n5664), .A2(n4831), .ZN(n4828) );
  OR2_X1 U5482 ( .A1(n5446), .A2(n4961), .ZN(n4963) );
  NAND2_X1 U5483 ( .A1(n6821), .A2(n6822), .ZN(n4843) );
  OR2_X1 U5484 ( .A1(n6821), .A2(n6822), .ZN(n4844) );
  NAND2_X1 U5485 ( .A1(n5553), .A2(n4313), .ZN(n5556) );
  AND2_X1 U5486 ( .A1(n5700), .A2(n5699), .ZN(n8925) );
  NOR2_X1 U5487 ( .A1(n5694), .A2(n5693), .ZN(n5695) );
  OR2_X1 U5488 ( .A1(n5319), .A2(n5318), .ZN(n5338) );
  OR2_X1 U5489 ( .A1(n5338), .A2(n8954), .ZN(n5361) );
  NAND2_X1 U5490 ( .A1(n5628), .A2(n5627), .ZN(n7220) );
  NAND2_X1 U5491 ( .A1(n4832), .A2(n5657), .ZN(n8986) );
  NAND2_X1 U5492 ( .A1(n8843), .A2(n5662), .ZN(n4832) );
  OAI21_X1 U5493 ( .B1(n8843), .B2(n4831), .A(n5664), .ZN(n8987) );
  OR2_X1 U5494 ( .A1(n5202), .A2(n5201), .ZN(n5224) );
  NAND2_X1 U5495 ( .A1(n4410), .A2(n7717), .ZN(n7790) );
  NAND2_X1 U5496 ( .A1(n5469), .A2(n5468), .ZN(n5471) );
  AOI21_X1 U5497 ( .B1(n9087), .B2(n5460), .A(n5432), .ZN(n9003) );
  AND3_X1 U5498 ( .A1(n5417), .A2(n5416), .A3(n5415), .ZN(n5796) );
  AND4_X1 U5499 ( .A1(n5134), .A2(n5133), .A3(n5132), .A4(n5131), .ZN(n5635)
         );
  NOR2_X1 U5500 ( .A1(n6237), .A2(n6238), .ZN(n6236) );
  OR2_X1 U5501 ( .A1(n6236), .A2(n4517), .ZN(n9596) );
  NOR2_X1 U5502 ( .A1(n6242), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4517) );
  NAND2_X1 U5503 ( .A1(n9596), .A2(n9597), .ZN(n9595) );
  NAND2_X1 U5504 ( .A1(n6008), .A2(n4519), .ZN(n9616) );
  NAND2_X1 U5505 ( .A1(n4521), .A2(n4520), .ZN(n4519) );
  INV_X1 U5506 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n4520) );
  NAND2_X1 U5507 ( .A1(n9616), .A2(n9617), .ZN(n9615) );
  OR2_X1 U5508 ( .A1(n5841), .A2(n5842), .ZN(n5872) );
  NOR2_X1 U5509 ( .A1(n9029), .A2(n4523), .ZN(n9631) );
  AND2_X1 U5510 ( .A1(n9030), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4523) );
  NOR2_X1 U5511 ( .A1(n9631), .A2(n9630), .ZN(n9629) );
  XNOR2_X1 U5512 ( .A(n9031), .B(n9043), .ZN(n9643) );
  NOR2_X1 U5513 ( .A1(n9679), .A2(n4526), .ZN(n9695) );
  AND2_X1 U5514 ( .A1(n9039), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4526) );
  NOR2_X1 U5515 ( .A1(n9695), .A2(n9696), .ZN(n9694) );
  NAND2_X1 U5516 ( .A1(n4615), .A2(n4620), .ZN(n9070) );
  AOI21_X1 U5517 ( .B1(n4627), .B2(n4623), .A(n4621), .ZN(n4620) );
  OR2_X1 U5518 ( .A1(n9084), .A2(n9302), .ZN(n9073) );
  INV_X1 U5519 ( .A(n4553), .ZN(n4551) );
  NOR2_X1 U5520 ( .A1(n9120), .A2(n4555), .ZN(n4552) );
  AOI21_X1 U5521 ( .B1(n4557), .B2(n7566), .A(n4554), .ZN(n4553) );
  NAND2_X1 U5522 ( .A1(n9110), .A2(n9489), .ZN(n4572) );
  NOR2_X1 U5523 ( .A1(n4559), .A2(n9092), .ZN(n4557) );
  NAND2_X1 U5524 ( .A1(n4558), .A2(n4556), .ZN(n9091) );
  INV_X1 U5525 ( .A(n4559), .ZN(n4556) );
  AND2_X1 U5526 ( .A1(n5449), .A2(n5448), .ZN(n9090) );
  AND2_X1 U5527 ( .A1(n9116), .A2(n9104), .ZN(n9100) );
  NAND2_X1 U5528 ( .A1(n9161), .A2(n4503), .ZN(n9133) );
  NAND2_X1 U5529 ( .A1(n9161), .A2(n9147), .ZN(n9142) );
  INV_X1 U5530 ( .A(n7746), .ZN(n9149) );
  AND2_X1 U5531 ( .A1(n7676), .A2(n7675), .ZN(n9166) );
  NAND2_X1 U5532 ( .A1(n9243), .A2(n4513), .ZN(n9186) );
  AND2_X1 U5533 ( .A1(n4322), .A2(n9339), .ZN(n4513) );
  AOI21_X1 U5534 ( .B1(n4324), .B2(n4638), .A(n4369), .ZN(n4634) );
  NAND2_X1 U5535 ( .A1(n9177), .A2(n5527), .ZN(n9179) );
  NAND2_X1 U5536 ( .A1(n9213), .A2(n7664), .ZN(n9200) );
  NAND2_X1 U5537 ( .A1(n9243), .A2(n4322), .ZN(n9194) );
  AND2_X1 U5538 ( .A1(n9243), .A2(n9239), .ZN(n9233) );
  NAND2_X1 U5539 ( .A1(n9243), .A2(n4514), .ZN(n9207) );
  AND2_X1 U5540 ( .A1(n7660), .A2(n7664), .ZN(n9215) );
  INV_X1 U5541 ( .A(n5263), .ZN(n5261) );
  OR2_X1 U5542 ( .A1(n9255), .A2(n4564), .ZN(n9226) );
  INV_X1 U5543 ( .A(n4498), .ZN(n4497) );
  NOR3_X1 U5544 ( .A1(n9502), .A2(n8848), .A3(n8938), .ZN(n9279) );
  INV_X1 U5545 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5163) );
  NOR2_X1 U5546 ( .A1(n9502), .A2(n8938), .ZN(n7211) );
  NAND2_X1 U5547 ( .A1(n5522), .A2(n7616), .ZN(n7193) );
  OR2_X1 U5548 ( .A1(n9501), .A2(n9495), .ZN(n9502) );
  OAI211_X1 U5549 ( .C1(n5061), .C2(n5931), .A(n5123), .B(n5122), .ZN(n7226)
         );
  NOR2_X1 U5550 ( .A1(n7082), .A2(n7133), .ZN(n7098) );
  OR2_X1 U5551 ( .A1(n9717), .A2(n7046), .ZN(n7082) );
  AND4_X1 U5552 ( .A1(n5094), .A2(n5093), .A3(n5092), .A4(n5091), .ZN(n6932)
         );
  NAND4_X1 U5553 ( .A1(n4505), .A2(n9837), .A3(n9842), .A4(n4504), .ZN(n9717)
         );
  INV_X1 U5554 ( .A(n9761), .ZN(n4504) );
  INV_X1 U5555 ( .A(n4506), .ZN(n4505) );
  AND4_X1 U5556 ( .A1(n5072), .A2(n5071), .A3(n5070), .A4(n5069), .ZN(n9721)
         );
  NAND2_X1 U5557 ( .A1(n6920), .A2(n9837), .ZN(n9716) );
  INV_X1 U5558 ( .A(n5518), .ZN(n7594) );
  OAI21_X1 U5559 ( .B1(n9737), .B2(n9747), .A(n5002), .ZN(n6832) );
  NOR2_X1 U5560 ( .A1(n4506), .A2(n9761), .ZN(n6920) );
  AND2_X1 U5561 ( .A1(n6671), .A2(n4931), .ZN(n6688) );
  INV_X1 U5562 ( .A(n9772), .ZN(n9742) );
  NAND2_X1 U5563 ( .A1(n5391), .A2(n5390), .ZN(n9317) );
  NAND2_X1 U5564 ( .A1(n5372), .A2(n5371), .ZN(n9323) );
  NAND2_X1 U5565 ( .A1(n5337), .A2(n5336), .ZN(n9332) );
  NAND2_X1 U5566 ( .A1(n5242), .A2(n5241), .ZN(n9359) );
  AND2_X1 U5567 ( .A1(n9730), .A2(n9832), .ZN(n9514) );
  INV_X1 U5568 ( .A(n9495), .ZN(n9541) );
  INV_X1 U5569 ( .A(n7226), .ZN(n9545) );
  INV_X1 U5570 ( .A(n9827), .ZN(n9849) );
  AND2_X1 U5571 ( .A1(n6090), .A2(n6089), .ZN(n6100) );
  AND2_X1 U5572 ( .A1(n7788), .A2(n7776), .ZN(n6093) );
  NAND2_X1 U5573 ( .A1(n5504), .A2(n5487), .ZN(n9378) );
  XNOR2_X1 U5574 ( .A(n7327), .B(n5456), .ZN(n8828) );
  XNOR2_X1 U5575 ( .A(n5451), .B(n5450), .ZN(n8039) );
  INV_X1 U5576 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5476) );
  XNOR2_X1 U5577 ( .A(n5383), .B(n5381), .ZN(n7353) );
  OAI21_X1 U5578 ( .B1(n5348), .B2(n5347), .A(n5346), .ZN(n5355) );
  AND2_X1 U5579 ( .A1(n5369), .A2(n5353), .ZN(n5354) );
  INV_X1 U5580 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5473) );
  INV_X1 U5581 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5217) );
  OAI21_X1 U5582 ( .B1(n5174), .B2(n4337), .A(n4729), .ZN(n5231) );
  NAND2_X1 U5583 ( .A1(n4745), .A2(n5140), .ZN(n5154) );
  NAND2_X1 U5584 ( .A1(n5118), .A2(n4746), .ZN(n4745) );
  XNOR2_X1 U5585 ( .A(n5095), .B(n4858), .ZN(n6703) );
  NAND2_X1 U5586 ( .A1(n4741), .A2(n4739), .ZN(n5075) );
  INV_X1 U5587 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4868) );
  AND3_X1 U5588 ( .A1(n4866), .A2(n4993), .A3(n4867), .ZN(n5037) );
  XNOR2_X1 U5589 ( .A(n5052), .B(n5050), .ZN(n6496) );
  NAND2_X1 U5590 ( .A1(n6103), .A2(n4896), .ZN(n4906) );
  AND4_X1 U5591 ( .A1(n6220), .A2(n6219), .A3(n6218), .A4(n6217), .ZN(n6657)
         );
  NAND2_X1 U5592 ( .A1(n4669), .A2(n4667), .ZN(n6593) );
  AOI21_X1 U5593 ( .B1(n4670), .B2(n6416), .A(n4668), .ZN(n4667) );
  INV_X1 U5594 ( .A(n6494), .ZN(n4668) );
  NAND2_X1 U5595 ( .A1(n4661), .A2(n6967), .ZN(n7057) );
  NAND2_X1 U5596 ( .A1(n6702), .A2(n4662), .ZN(n4661) );
  AND4_X1 U5597 ( .A1(n6806), .A2(n6805), .A3(n6804), .A4(n6803), .ZN(n6993)
         );
  INV_X1 U5598 ( .A(n8129), .ZN(n9881) );
  NAND2_X1 U5599 ( .A1(n4659), .A2(n4657), .ZN(n8067) );
  AND2_X1 U5600 ( .A1(n4659), .A2(n4347), .ZN(n8069) );
  NAND2_X1 U5601 ( .A1(n8142), .A2(n8141), .ZN(n4659) );
  AND4_X1 U5602 ( .A1(n6429), .A2(n6428), .A3(n6427), .A4(n6426), .ZN(n6634)
         );
  OAI22_X1 U5603 ( .A1(n6593), .A2(n6592), .B1(n6591), .B2(n6590), .ZN(n6697)
         );
  INV_X1 U5604 ( .A(n8192), .ZN(n8038) );
  NAND2_X1 U5605 ( .A1(n8034), .A2(n8033), .ZN(n8032) );
  AND4_X1 U5606 ( .A1(n7158), .A2(n7157), .A3(n7156), .A4(n7155), .ZN(n8101)
         );
  NAND2_X1 U5607 ( .A1(n8095), .A2(n7282), .ZN(n7361) );
  NAND2_X1 U5608 ( .A1(n7285), .A2(n7284), .ZN(n8594) );
  AND4_X1 U5609 ( .A1(n6508), .A2(n6507), .A3(n6506), .A4(n6505), .ZN(n6719)
         );
  OAI21_X1 U5610 ( .B1(n8142), .B2(n4658), .A(n4654), .ZN(n8117) );
  NAND2_X1 U5611 ( .A1(n7389), .A2(n7388), .ZN(n8578) );
  NAND2_X1 U5612 ( .A1(n7055), .A2(n4441), .ZN(n7173) );
  AND4_X1 U5613 ( .A1(n6718), .A2(n6717), .A3(n6716), .A4(n6715), .ZN(n6979)
         );
  XNOR2_X1 U5614 ( .A(n7003), .B(n7004), .ZN(n6977) );
  AND4_X1 U5615 ( .A1(n7379), .A2(n7378), .A3(n7377), .A4(n7376), .ZN(n8456)
         );
  OR2_X1 U5616 ( .A1(n8129), .A2(n8457), .ZN(n8145) );
  NAND2_X1 U5617 ( .A1(n4432), .A2(n7359), .ZN(n8142) );
  NAND2_X1 U5618 ( .A1(n8095), .A2(n4437), .ZN(n4432) );
  NAND2_X1 U5619 ( .A1(n4671), .A2(n4670), .ZN(n6495) );
  OR2_X1 U5620 ( .A1(n8129), .A2(n8455), .ZN(n8156) );
  INV_X1 U5621 ( .A(n9882), .ZN(n8150) );
  INV_X1 U5622 ( .A(n9891), .ZN(n8158) );
  OR3_X1 U5623 ( .A1(n6063), .A2(n9930), .A3(n6262), .ZN(n9882) );
  NAND2_X1 U5624 ( .A1(n7238), .A2(n7237), .ZN(n8280) );
  INV_X1 U5625 ( .A(n8025), .ZN(n4409) );
  OR2_X1 U5626 ( .A1(n9904), .A2(n6057), .ZN(n8026) );
  XNOR2_X1 U5627 ( .A(n5933), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8027) );
  AND3_X1 U5628 ( .A1(n5926), .A2(n5925), .A3(n5924), .ZN(n8305) );
  INV_X1 U5629 ( .A(n8325), .ZN(n8364) );
  OR2_X1 U5630 ( .A1(n6259), .A2(n5840), .ZN(n8175) );
  INV_X1 U5631 ( .A(n8101), .ZN(n8606) );
  NOR2_X1 U5632 ( .A1(n6336), .A2(n6257), .ZN(n4753) );
  INV_X1 U5633 ( .A(n4752), .ZN(n6282) );
  AND2_X1 U5634 ( .A1(n4750), .A2(n4749), .ZN(n6298) );
  INV_X1 U5635 ( .A(n6285), .ZN(n4749) );
  INV_X1 U5636 ( .A(n4750), .ZN(n6286) );
  INV_X1 U5637 ( .A(n4760), .ZN(n6314) );
  AND2_X1 U5638 ( .A1(n4760), .A2(n4759), .ZN(n6317) );
  NAND2_X1 U5639 ( .A1(n6315), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4759) );
  INV_X1 U5640 ( .A(n4758), .ZN(n6339) );
  NOR2_X1 U5641 ( .A1(n6371), .A2(n6370), .ZN(n6369) );
  AND2_X1 U5642 ( .A1(n4758), .A2(n4757), .ZN(n6371) );
  NAND2_X1 U5643 ( .A1(n6345), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4757) );
  AND2_X1 U5644 ( .A1(n6704), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4767) );
  NOR2_X1 U5645 ( .A1(n6358), .A2(n6357), .ZN(n6729) );
  AND2_X1 U5646 ( .A1(n5952), .A2(n5959), .ZN(n6941) );
  NAND2_X1 U5647 ( .A1(n8193), .A2(n4405), .ZN(n6732) );
  OR2_X1 U5648 ( .A1(n8199), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4405) );
  INV_X1 U5649 ( .A(n4765), .ZN(n6777) );
  OR2_X1 U5650 ( .A1(n7059), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4761) );
  NAND2_X1 U5651 ( .A1(n7019), .A2(n4763), .ZN(n4762) );
  INV_X1 U5652 ( .A(n7020), .ZN(n4763) );
  NOR2_X1 U5653 ( .A1(n8262), .A2(n6052), .ZN(n9897) );
  AND2_X1 U5654 ( .A1(n6275), .A2(n6264), .ZN(n9892) );
  INV_X1 U5655 ( .A(n8228), .ZN(n8220) );
  INV_X1 U5656 ( .A(n4756), .ZN(n8237) );
  NOR2_X1 U5657 ( .A1(n8276), .A2(n4542), .ZN(n4541) );
  NAND2_X1 U5658 ( .A1(n4543), .A2(n8341), .ZN(n4542) );
  NAND2_X1 U5659 ( .A1(n8361), .A2(n4784), .ZN(n8347) );
  NAND2_X1 U5660 ( .A1(n8376), .A2(n8375), .ZN(n8374) );
  OAI21_X1 U5661 ( .B1(n8402), .B2(n4692), .A(n4690), .ZN(n8370) );
  NAND2_X1 U5662 ( .A1(n4689), .A2(n4694), .ZN(n8372) );
  NAND2_X1 U5663 ( .A1(n8402), .A2(n4696), .ZN(n8388) );
  NAND2_X1 U5664 ( .A1(n4448), .A2(n4453), .ZN(n8403) );
  NAND2_X1 U5665 ( .A1(n8432), .A2(n4454), .ZN(n4448) );
  AND2_X1 U5666 ( .A1(n4455), .A2(n4346), .ZN(n8418) );
  NAND2_X1 U5667 ( .A1(n8432), .A2(n8292), .ZN(n4455) );
  NAND2_X1 U5668 ( .A1(n4678), .A2(n4682), .ZN(n8449) );
  OR2_X1 U5669 ( .A1(n8488), .A2(n4684), .ZN(n4678) );
  NAND2_X1 U5670 ( .A1(n7372), .A2(n7371), .ZN(n8584) );
  NAND2_X1 U5671 ( .A1(n4686), .A2(n4685), .ZN(n8464) );
  AND2_X1 U5672 ( .A1(n4686), .A2(n4351), .ZN(n8465) );
  NAND2_X1 U5673 ( .A1(n8488), .A2(n8489), .ZN(n4686) );
  INV_X1 U5674 ( .A(n8588), .ZN(n8498) );
  NAND2_X1 U5675 ( .A1(n7240), .A2(n7239), .ZN(n7813) );
  INV_X1 U5676 ( .A(n8437), .ZN(n9435) );
  NAND2_X1 U5677 ( .A1(n6844), .A2(n6843), .ZN(n6848) );
  NAND2_X1 U5678 ( .A1(n6794), .A2(n6793), .ZN(n6994) );
  OR2_X1 U5679 ( .A1(n6791), .A2(n6790), .ZN(n6794) );
  NAND2_X1 U5680 ( .A1(n6749), .A2(n6748), .ZN(n6750) );
  OR2_X1 U5681 ( .A1(n6594), .A2(n6790), .ZN(n6597) );
  NAND2_X1 U5682 ( .A1(n6515), .A2(n4316), .ZN(n6463) );
  INV_X1 U5683 ( .A(n9936), .ZN(n9885) );
  NAND2_X1 U5684 ( .A1(n9441), .A2(n6389), .ZN(n9438) );
  INV_X1 U5685 ( .A(n9438), .ZN(n8484) );
  AND2_X1 U5686 ( .A1(n9448), .A2(n9456), .ZN(n8494) );
  AND2_X2 U5687 ( .A1(n8614), .A2(n8529), .ZN(n10023) );
  NAND2_X1 U5688 ( .A1(n4461), .A2(n4459), .ZN(n8616) );
  NAND2_X1 U5689 ( .A1(n8534), .A2(n10001), .ZN(n4461) );
  AND2_X1 U5690 ( .A1(n6158), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9912) );
  NAND2_X1 U5691 ( .A1(n5923), .A2(n5922), .ZN(n8829) );
  OR2_X1 U5692 ( .A1(n5920), .A2(n5919), .ZN(n5921) );
  NAND2_X1 U5693 ( .A1(n5833), .A2(n5832), .ZN(n8836) );
  XNOR2_X1 U5694 ( .A(n5818), .B(n5817), .ZN(n7143) );
  INV_X1 U5695 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5817) );
  NAND2_X1 U5696 ( .A1(n5839), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5818) );
  INV_X1 U5697 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8702) );
  INV_X1 U5698 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7418) );
  INV_X1 U5699 ( .A(n8027), .ZN(n8531) );
  INV_X1 U5700 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7401) );
  INV_X1 U5701 ( .A(n8020), .ZN(n7836) );
  INV_X1 U5702 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7387) );
  AOI21_X1 U5703 ( .B1(n4314), .B2(n4649), .A(n4646), .ZN(n4645) );
  NAND2_X1 U5704 ( .A1(n4648), .A2(n4647), .ZN(n4646) );
  INV_X1 U5705 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6587) );
  INV_X1 U5706 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6198) );
  INV_X1 U5707 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6194) );
  INV_X1 U5708 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n5962) );
  INV_X1 U5709 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5912) );
  INV_X1 U5710 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5916) );
  INV_X1 U5711 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6407) );
  INV_X1 U5712 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6209) );
  INV_X1 U5713 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6150) );
  INV_X1 U5714 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U5715 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4771) );
  AND2_X1 U5716 ( .A1(n8048), .A2(n8977), .ZN(n8049) );
  NAND2_X1 U5717 ( .A1(n4838), .A2(n4839), .ZN(n8879) );
  AND4_X1 U5718 ( .A1(n5169), .A2(n5168), .A3(n5167), .A4(n5166), .ZN(n7264)
         );
  NAND2_X1 U5719 ( .A1(n7220), .A2(n5633), .ZN(n7260) );
  NAND2_X1 U5720 ( .A1(n8915), .A2(n5732), .ZN(n8886) );
  AND4_X1 U5721 ( .A1(n5010), .A2(n5009), .A3(n5008), .A4(n5007), .ZN(n6919)
         );
  AND4_X1 U5722 ( .A1(n5268), .A2(n5267), .A3(n5266), .A4(n5265), .ZN(n8911)
         );
  OAI211_X1 U5723 ( .C1(n5104), .C2(n6149), .A(n4976), .B(n4975), .ZN(n9758)
         );
  AND4_X1 U5724 ( .A1(n5049), .A2(n5048), .A3(n5047), .A4(n5046), .ZN(n7044)
         );
  INV_X1 U5725 ( .A(n9850), .ZN(n7046) );
  AOI21_X1 U5726 ( .B1(n5709), .B2(n5708), .A(n8923), .ZN(n8927) );
  NAND3_X1 U5727 ( .A1(n4930), .A2(n4929), .A3(n4928), .ZN(n8964) );
  NAND2_X1 U5728 ( .A1(n5278), .A2(n4927), .ZN(n4928) );
  INV_X1 U5729 ( .A(n9000), .ZN(n8965) );
  INV_X1 U5730 ( .A(n8994), .ZN(n8966) );
  AND4_X1 U5731 ( .A1(n5031), .A2(n5030), .A3(n5029), .A4(n5028), .ZN(n9722)
         );
  INV_X1 U5732 ( .A(n9286), .ZN(n9520) );
  INV_X1 U5733 ( .A(n9090), .ZN(n9002) );
  INV_X1 U5734 ( .A(n5733), .ZN(n9131) );
  INV_X1 U5735 ( .A(n5668), .ZN(n9276) );
  INV_X1 U5736 ( .A(n7264), .ZN(n9491) );
  INV_X1 U5737 ( .A(n6932), .ZN(n9005) );
  INV_X1 U5738 ( .A(n9721), .ZN(n9006) );
  INV_X1 U5739 ( .A(n9773), .ZN(n9009) );
  NAND2_X1 U5740 ( .A1(n9020), .A2(n9019), .ZN(n9024) );
  NOR2_X1 U5741 ( .A1(n9607), .A2(n4344), .ZN(n6009) );
  NAND2_X1 U5742 ( .A1(n6009), .A2(n6010), .ZN(n6008) );
  INV_X1 U5743 ( .A(n4518), .ZN(n9654) );
  AND2_X1 U5744 ( .A1(n4518), .A2(n4381), .ZN(n9668) );
  XNOR2_X1 U5745 ( .A(n4524), .B(n9037), .ZN(n9055) );
  OR2_X1 U5746 ( .A1(n9694), .A2(n4525), .ZN(n4524) );
  AND2_X1 U5747 ( .A1(n9038), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4525) );
  INV_X1 U5748 ( .A(n9708), .ZN(n9688) );
  NAND2_X1 U5749 ( .A1(n4632), .A2(n4626), .ZN(n4630) );
  NOR2_X1 U5750 ( .A1(n4625), .A2(n4624), .ZN(n9099) );
  INV_X1 U5751 ( .A(n4631), .ZN(n4624) );
  INV_X1 U5752 ( .A(n4632), .ZN(n4625) );
  INV_X1 U5753 ( .A(n9323), .ZN(n9128) );
  NAND2_X1 U5754 ( .A1(n4635), .A2(n4636), .ZN(n9193) );
  OR2_X1 U5755 ( .A1(n9223), .A2(n4638), .ZN(n4635) );
  NAND2_X1 U5756 ( .A1(n4603), .A2(n4604), .ZN(n9242) );
  OR2_X1 U5757 ( .A1(n9271), .A2(n4606), .ZN(n4603) );
  NAND2_X1 U5758 ( .A1(n4607), .A2(n5208), .ZN(n9254) );
  OR2_X1 U5759 ( .A1(n9271), .A2(n5209), .ZN(n4607) );
  NAND2_X1 U5760 ( .A1(n9497), .A2(n5151), .ZN(n7191) );
  NAND2_X1 U5761 ( .A1(n9712), .A2(n5065), .ZN(n6933) );
  OAI211_X1 U5762 ( .C1(n5104), .C2(n6134), .A(n4955), .B(n4954), .ZN(n6692)
         );
  NAND2_X1 U5763 ( .A1(n4992), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4516) );
  NAND2_X1 U5764 ( .A1(n5278), .A2(n5882), .ZN(n4515) );
  INV_X2 U5765 ( .A(n9779), .ZN(n9755) );
  INV_X1 U5766 ( .A(n9765), .ZN(n9494) );
  AND2_X2 U5767 ( .A1(n6100), .A2(n6099), .ZN(n9879) );
  AOI211_X1 U5768 ( .C1(n9827), .C2(n9512), .A(n9511), .B(n9510), .ZN(n9552)
         );
  NAND2_X1 U5769 ( .A1(n5841), .A2(n5508), .ZN(n9791) );
  NAND2_X1 U5770 ( .A1(n4875), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4880) );
  INV_X1 U5771 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n6929) );
  INV_X1 U5772 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6789) );
  INV_X1 U5773 ( .A(n7752), .ZN(n7776) );
  INV_X1 U5774 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6725) );
  INV_X1 U5775 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6589) );
  NAND2_X1 U5776 ( .A1(n5465), .A2(n5284), .ZN(n9136) );
  INV_X1 U5777 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6188) );
  INV_X1 U5778 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5958) );
  INV_X1 U5779 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8710) );
  INV_X1 U5780 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5931) );
  INV_X1 U5781 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5908) );
  XNOR2_X1 U5782 ( .A(n5116), .B(n5114), .ZN(n6791) );
  INV_X1 U5783 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5907) );
  NOR2_X1 U5784 ( .A1(n6893), .A2(n10057), .ZN(n10052) );
  AOI21_X1 U5785 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10050), .ZN(n10049) );
  NOR2_X1 U5786 ( .A1(n10049), .A2(n10048), .ZN(n10047) );
  AOI21_X1 U5787 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10047), .ZN(n10046) );
  AND2_X1 U5788 ( .A1(n7491), .A2(n4429), .ZN(n4428) );
  NAND2_X1 U5789 ( .A1(n4421), .A2(n4424), .ZN(n4420) );
  NAND2_X1 U5790 ( .A1(n4770), .A2(n4768), .ZN(n8267) );
  OAI21_X1 U5791 ( .B1(n8263), .B2(n8262), .A(n4769), .ZN(n4768) );
  NAND2_X1 U5792 ( .A1(n4576), .A2(n4575), .ZN(P2_U3549) );
  OR2_X1 U5793 ( .A1(n10023), .A2(n5981), .ZN(n4575) );
  NAND2_X1 U5794 ( .A1(n8616), .A2(n10023), .ZN(n4576) );
  OAI21_X1 U5795 ( .B1(n9089), .B2(n9000), .A(n5799), .ZN(n5800) );
  OAI21_X1 U5796 ( .B1(n9104), .B2(n9000), .A(n5774), .ZN(n5775) );
  OAI21_X1 U5797 ( .B1(n4413), .B2(n4411), .A(n7791), .ZN(n7793) );
  NOR2_X1 U5798 ( .A1(n5548), .A2(n5547), .ZN(n5549) );
  INV_X1 U5799 ( .A(n5546), .ZN(n5547) );
  OAI21_X1 U5800 ( .B1(n9305), .B2(n9755), .A(n4567), .ZN(P1_U3263) );
  NAND2_X1 U5801 ( .A1(n4570), .A2(n4569), .ZN(n4568) );
  INV_X1 U5802 ( .A(n9082), .ZN(n4569) );
  OR2_X1 U5803 ( .A1(n5824), .A2(n4675), .ZN(n4314) );
  NAND2_X1 U5804 ( .A1(n4725), .A2(n5271), .ZN(n4724) );
  OR2_X1 U5805 ( .A1(n9502), .A2(n4496), .ZN(n4315) );
  AND2_X1 U5806 ( .A1(n4721), .A2(n4718), .ZN(n4317) );
  XNOR2_X1 U5807 ( .A(n4771), .B(n5896), .ZN(n6271) );
  AND2_X1 U5808 ( .A1(n7853), .A2(n7975), .ZN(n4318) );
  AND2_X1 U5809 ( .A1(n5708), .A2(n5710), .ZN(n4319) );
  INV_X1 U5810 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6046) );
  INV_X2 U5811 ( .A(n5006), .ZN(n5246) );
  AND2_X1 U5812 ( .A1(n4608), .A2(n9256), .ZN(n4320) );
  XNOR2_X1 U5813 ( .A(n8304), .B(n8303), .ZN(n4321) );
  NAND2_X1 U5814 ( .A1(n7885), .A2(n7884), .ZN(n6637) );
  INV_X1 U5815 ( .A(n6637), .ZN(n8001) );
  AND2_X1 U5816 ( .A1(n4514), .A2(n9198), .ZN(n4322) );
  AND2_X1 U5817 ( .A1(n4604), .A2(n4358), .ZN(n4323) );
  AND2_X1 U5818 ( .A1(n4636), .A2(n4356), .ZN(n4324) );
  AND2_X1 U5819 ( .A1(n4307), .A2(n9624), .ZN(n4325) );
  OR2_X1 U5820 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4326) );
  NAND2_X1 U5821 ( .A1(n5438), .A2(n5437), .ZN(n9302) );
  INV_X1 U5822 ( .A(n9302), .ZN(n4511) );
  INV_X1 U5823 ( .A(n7611), .ZN(n4415) );
  AND2_X1 U5824 ( .A1(n9532), .A2(n7264), .ZN(n4327) );
  AND2_X1 U5825 ( .A1(n4804), .A2(n7941), .ZN(n4328) );
  INV_X1 U5826 ( .A(n7566), .ZN(n4560) );
  AND2_X1 U5827 ( .A1(n5064), .A2(n5087), .ZN(n4329) );
  AND2_X1 U5828 ( .A1(n4537), .A2(n4695), .ZN(n4330) );
  AND2_X1 U5829 ( .A1(n7399), .A2(n7398), .ZN(n4331) );
  NAND2_X1 U5830 ( .A1(n5286), .A2(n5285), .ZN(n9350) );
  AND2_X1 U5831 ( .A1(n7432), .A2(n7431), .ZN(n8408) );
  INV_X1 U5832 ( .A(n8408), .ZN(n8562) );
  AND2_X1 U5833 ( .A1(n4550), .A2(n7616), .ZN(n4332) );
  NAND2_X1 U5834 ( .A1(n7954), .A2(n4817), .ZN(n4816) );
  OR3_X1 U5835 ( .A1(n4314), .A2(P2_IR_REG_19__SCAN_IN), .A3(
        P2_IR_REG_20__SCAN_IN), .ZN(n4333) );
  NAND2_X1 U5836 ( .A1(n7827), .A2(n7826), .ZN(n8308) );
  INV_X1 U5837 ( .A(n8308), .ZN(n4546) );
  AND4_X1 U5838 ( .A1(n5238), .A2(n5218), .A3(n5236), .A4(n5468), .ZN(n4334)
         );
  AND2_X1 U5839 ( .A1(n7964), .A2(n7965), .ZN(n4335) );
  INV_X1 U5840 ( .A(n9167), .ZN(n8952) );
  INV_X1 U5841 ( .A(n4724), .ZN(n4723) );
  OR3_X1 U5842 ( .A1(n7117), .A2(n7913), .A3(n4534), .ZN(n4336) );
  OR2_X1 U5843 ( .A1(n9496), .A2(n9499), .ZN(n9497) );
  NAND2_X1 U5844 ( .A1(n5222), .A2(n5221), .ZN(n8894) );
  INV_X1 U5845 ( .A(n8894), .ZN(n4499) );
  INV_X1 U5846 ( .A(n4937), .ZN(n5414) );
  INV_X1 U5847 ( .A(n6758), .ZN(n9973) );
  INV_X1 U5848 ( .A(n7913), .ZN(n9465) );
  NAND2_X1 U5849 ( .A1(n7146), .A2(n7145), .ZN(n7913) );
  OR2_X1 U5850 ( .A1(n5211), .A2(n4731), .ZN(n4337) );
  OR2_X1 U5851 ( .A1(n5824), .A2(n4672), .ZN(n4338) );
  INV_X1 U5852 ( .A(n6402), .ZN(n6387) );
  NAND2_X1 U5853 ( .A1(n5455), .A2(n5454), .ZN(n7327) );
  NAND2_X1 U5854 ( .A1(n8986), .A2(n8985), .ZN(n8896) );
  INV_X1 U5855 ( .A(n7116), .ZN(n4535) );
  INV_X2 U5856 ( .A(n5061), .ZN(n5407) );
  AND2_X1 U5857 ( .A1(n4837), .A2(n4839), .ZN(n4339) );
  AND2_X1 U5858 ( .A1(n9089), .A2(n9003), .ZN(n4340) );
  INV_X1 U5859 ( .A(n6826), .ZN(n9842) );
  OR2_X1 U5860 ( .A1(n5153), .A2(n4744), .ZN(n4341) );
  NAND2_X1 U5861 ( .A1(n7269), .A2(n7271), .ZN(n4342) );
  OR2_X1 U5862 ( .A1(n8105), .A2(n4664), .ZN(n4343) );
  INV_X1 U5863 ( .A(n4628), .ZN(n4627) );
  NAND2_X1 U5864 ( .A1(n9092), .A2(n4629), .ZN(n4628) );
  AND2_X1 U5865 ( .A1(n4866), .A2(n4993), .ZN(n4997) );
  INV_X1 U5866 ( .A(n4658), .ZN(n4657) );
  NAND2_X1 U5867 ( .A1(n4347), .A2(n8068), .ZN(n4658) );
  NAND2_X1 U5868 ( .A1(n5893), .A2(n4780), .ZN(n5904) );
  INV_X1 U5869 ( .A(n8296), .ZN(n8394) );
  AND2_X1 U5870 ( .A1(n7947), .A2(n7952), .ZN(n8296) );
  AND2_X1 U5871 ( .A1(n9602), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4344) );
  AND2_X1 U5872 ( .A1(n4630), .A2(n4629), .ZN(n9083) );
  OR2_X1 U5873 ( .A1(n6501), .A2(n6336), .ZN(n4345) );
  NAND2_X1 U5874 ( .A1(n8573), .A2(n8291), .ZN(n4346) );
  NAND2_X1 U5875 ( .A1(n5174), .A2(n5173), .ZN(n5192) );
  INV_X1 U5876 ( .A(n8410), .ZN(n4450) );
  NAND2_X1 U5877 ( .A1(n7367), .A2(n7366), .ZN(n4347) );
  AND2_X1 U5878 ( .A1(n7948), .A2(n7978), .ZN(n4348) );
  INV_X1 U5879 ( .A(n8600), .ZN(n4582) );
  NAND2_X1 U5880 ( .A1(n6211), .A2(n4462), .ZN(n6476) );
  NAND2_X1 U5881 ( .A1(n8510), .A2(n7929), .ZN(n8467) );
  OR3_X1 U5882 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4350) );
  NAND2_X1 U5883 ( .A1(n8916), .A2(n8917), .ZN(n8915) );
  AND2_X1 U5884 ( .A1(n4972), .A2(n4864), .ZN(n4993) );
  NAND2_X1 U5885 ( .A1(n8498), .A2(n8287), .ZN(n4351) );
  INV_X1 U5886 ( .A(n7857), .ZN(n4777) );
  AND3_X1 U5887 ( .A1(n4829), .A2(n8897), .A3(n4828), .ZN(n4352) );
  INV_X1 U5888 ( .A(n8448), .ZN(n4680) );
  AND2_X1 U5889 ( .A1(n5407), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n4353) );
  NAND2_X1 U5890 ( .A1(n5877), .A2(n4778), .ZN(n5886) );
  AND2_X1 U5891 ( .A1(n4558), .A2(n4557), .ZN(n4354) );
  NAND2_X1 U5892 ( .A1(n6597), .A2(n6596), .ZN(n6747) );
  NOR2_X1 U5893 ( .A1(n8021), .A2(n8020), .ZN(n4355) );
  NAND2_X1 U5894 ( .A1(n5260), .A2(n5259), .ZN(n9356) );
  NAND2_X1 U5895 ( .A1(n9344), .A2(n9216), .ZN(n4356) );
  OR2_X1 U5896 ( .A1(n4511), .A2(n9090), .ZN(n4357) );
  NAND2_X1 U5897 ( .A1(n9359), .A2(n9261), .ZN(n4358) );
  NAND2_X1 U5898 ( .A1(n8439), .A2(n4539), .ZN(n4540) );
  AND2_X1 U5899 ( .A1(n9350), .A2(n9230), .ZN(n4359) );
  AND2_X1 U5900 ( .A1(n7403), .A2(n7402), .ZN(n8290) );
  INV_X1 U5901 ( .A(n8290), .ZN(n8573) );
  XNOR2_X1 U5902 ( .A(n8302), .B(n8304), .ZN(n8534) );
  INV_X1 U5903 ( .A(n8061), .ZN(n8295) );
  AND2_X1 U5904 ( .A1(n7352), .A2(n7351), .ZN(n8061) );
  AND2_X1 U5905 ( .A1(n4690), .A2(n4446), .ZN(n4360) );
  INV_X1 U5906 ( .A(n4992), .ZN(n5061) );
  INV_X1 U5907 ( .A(n7192), .ZN(n4550) );
  NAND2_X1 U5908 ( .A1(n7896), .A2(n7978), .ZN(n4361) );
  INV_X1 U5909 ( .A(n8276), .ZN(n9453) );
  INV_X1 U5910 ( .A(n4697), .ZN(n4696) );
  AND2_X1 U5911 ( .A1(n8894), .A2(n9276), .ZN(n4362) );
  AND2_X1 U5912 ( .A1(n4823), .A2(n8887), .ZN(n4363) );
  NAND2_X1 U5913 ( .A1(n6608), .A2(n7869), .ZN(n7990) );
  INV_X1 U5914 ( .A(n7950), .ZN(n4491) );
  INV_X1 U5915 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5938) );
  NOR2_X1 U5916 ( .A1(n4546), .A2(n9994), .ZN(n4364) );
  INV_X1 U5917 ( .A(n4426), .ZN(n4425) );
  NAND2_X1 U5918 ( .A1(n7476), .A2(n4427), .ZN(n4426) );
  NOR2_X1 U5919 ( .A1(n9359), .A2(n9261), .ZN(n4365) );
  AND2_X1 U5920 ( .A1(n4838), .A2(n4339), .ZN(n4366) );
  NOR2_X1 U5921 ( .A1(n8554), .A2(n8365), .ZN(n4367) );
  INV_X1 U5922 ( .A(n4816), .ZN(n4815) );
  OR2_X1 U5923 ( .A1(n4460), .A2(n4364), .ZN(n4368) );
  NOR2_X1 U5924 ( .A1(n9344), .A2(n9216), .ZN(n4369) );
  INV_X1 U5925 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5482) );
  AND2_X1 U5926 ( .A1(n9973), .A2(n6807), .ZN(n4370) );
  NOR2_X1 U5927 ( .A1(n8288), .A2(n8456), .ZN(n4371) );
  NAND2_X1 U5928 ( .A1(n5717), .A2(n5716), .ZN(n4372) );
  AND2_X1 U5929 ( .A1(n4642), .A2(n4640), .ZN(n5480) );
  INV_X1 U5930 ( .A(n4858), .ZN(n4813) );
  NAND2_X1 U5931 ( .A1(n4642), .A2(n4641), .ZN(n4373) );
  AND4_X1 U5932 ( .A1(n4873), .A2(n4872), .A3(n4874), .A4(n4644), .ZN(n4374)
         );
  INV_X1 U5933 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5506) );
  OAI21_X1 U5934 ( .B1(n4490), .B2(n4488), .A(n4814), .ZN(n4487) );
  AND2_X1 U5935 ( .A1(n4658), .A2(n4653), .ZN(n4375) );
  NOR2_X1 U5936 ( .A1(n6965), .A2(n4663), .ZN(n4662) );
  NAND2_X1 U5937 ( .A1(n9006), .A2(n7046), .ZN(n4376) );
  OR2_X1 U5938 ( .A1(n9307), .A2(n9003), .ZN(n7770) );
  AND2_X1 U5939 ( .A1(n4489), .A2(n4815), .ZN(n4377) );
  AND2_X1 U5940 ( .A1(n7908), .A2(n7907), .ZN(n8003) );
  NAND2_X1 U5941 ( .A1(n8423), .A2(n4346), .ZN(n4378) );
  AND2_X1 U5942 ( .A1(n8375), .A2(n7952), .ZN(n4379) );
  NAND2_X1 U5943 ( .A1(n6807), .A2(n6758), .ZN(n7887) );
  AND2_X1 U5944 ( .A1(n4654), .A2(n4653), .ZN(n4380) );
  OR2_X1 U5945 ( .A1(n8542), .A2(n8325), .ZN(n7957) );
  INV_X1 U5946 ( .A(n7957), .ZN(n4782) );
  AND2_X1 U5947 ( .A1(n7614), .A2(n7635), .ZN(n9499) );
  OR2_X1 U5948 ( .A1(n9033), .A2(n9045), .ZN(n4381) );
  AND2_X1 U5949 ( .A1(n7892), .A2(n7895), .ZN(n8000) );
  AND2_X1 U5950 ( .A1(n4421), .A2(n4426), .ZN(n4382) );
  INV_X1 U5951 ( .A(n9307), .ZN(n9089) );
  OR2_X1 U5952 ( .A1(n5664), .A2(n4826), .ZN(n4383) );
  AND2_X1 U5953 ( .A1(n5636), .A2(n5633), .ZN(n4384) );
  AND2_X1 U5954 ( .A1(n8006), .A2(n7106), .ZN(n4385) );
  AND2_X1 U5955 ( .A1(n7984), .A2(n4791), .ZN(n4386) );
  NAND2_X1 U5956 ( .A1(n6468), .A2(n7856), .ZN(n4387) );
  AND2_X1 U5957 ( .A1(n5804), .A2(n5805), .ZN(n4780) );
  OR2_X1 U5958 ( .A1(n4326), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4388) );
  INV_X1 U5959 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6541) );
  NAND2_X1 U5960 ( .A1(n4333), .A2(n4645), .ZN(n6109) );
  OAI211_X1 U5961 ( .C1(n5104), .C2(n6208), .A(n5001), .B(n5000), .ZN(n9739)
         );
  INV_X1 U5962 ( .A(n8537), .ZN(n4545) );
  NOR2_X1 U5963 ( .A1(n6752), .A2(n6637), .ZN(n4389) );
  NAND2_X1 U5964 ( .A1(n7270), .A2(n7269), .ZN(n4390) );
  NAND2_X1 U5965 ( .A1(n7356), .A2(n7355), .ZN(n8558) );
  INV_X1 U5966 ( .A(n8558), .ZN(n4695) );
  NAND2_X1 U5967 ( .A1(n5303), .A2(n5302), .ZN(n9344) );
  NOR2_X1 U5968 ( .A1(n8477), .A2(n8578), .ZN(n8439) );
  NAND2_X1 U5969 ( .A1(n5458), .A2(n5457), .ZN(n9297) );
  INV_X1 U5970 ( .A(n9297), .ZN(n4512) );
  NOR3_X1 U5971 ( .A1(n7117), .A2(n4533), .A3(n7913), .ZN(n4532) );
  NAND2_X1 U5972 ( .A1(n4708), .A2(n8281), .ZN(n8598) );
  NAND2_X1 U5973 ( .A1(n5120), .A2(n4871), .ZN(n5145) );
  NAND2_X1 U5974 ( .A1(n5358), .A2(n5357), .ZN(n9327) );
  INV_X1 U5975 ( .A(n9327), .ZN(n9147) );
  INV_X1 U5976 ( .A(n9532), .ZN(n8938) );
  AND2_X1 U5977 ( .A1(n5162), .A2(n5161), .ZN(n9532) );
  AND2_X1 U5978 ( .A1(n7940), .A2(n4484), .ZN(n4391) );
  AND2_X1 U5979 ( .A1(n7925), .A2(n8509), .ZN(n8599) );
  AND2_X1 U5980 ( .A1(n6749), .A2(n4712), .ZN(n4392) );
  INV_X1 U5981 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6047) );
  NAND2_X1 U5982 ( .A1(n8610), .A2(n8284), .ZN(n4393) );
  AND2_X1 U5983 ( .A1(n5273), .A2(SI_18_), .ZN(n4394) );
  NAND2_X1 U5984 ( .A1(n6798), .A2(n6797), .ZN(n4395) );
  OR2_X1 U5985 ( .A1(n5824), .A2(n4674), .ZN(n4396) );
  NOR2_X1 U5986 ( .A1(n9255), .A2(n5525), .ZN(n4397) );
  NAND2_X1 U5987 ( .A1(n5317), .A2(n5316), .ZN(n9185) );
  INV_X1 U5988 ( .A(n9185), .ZN(n9339) );
  AND2_X1 U5989 ( .A1(n4865), .A2(n4864), .ZN(n4398) );
  AND2_X1 U5990 ( .A1(n6162), .A2(n6058), .ZN(n9886) );
  NAND2_X1 U5991 ( .A1(n5828), .A2(n5827), .ZN(n5831) );
  OR2_X1 U5992 ( .A1(n4530), .A2(n6613), .ZN(n4399) );
  NAND2_X1 U5993 ( .A1(n4463), .A2(n6633), .ZN(n6654) );
  INV_X1 U5994 ( .A(n6967), .ZN(n4660) );
  NAND2_X1 U5995 ( .A1(n4842), .A2(n4843), .ZN(n7036) );
  OR2_X1 U5996 ( .A1(n9761), .A2(n9739), .ZN(n4400) );
  OR2_X1 U5997 ( .A1(n5082), .A2(n4643), .ZN(n4401) );
  NAND2_X1 U5998 ( .A1(n4612), .A2(n5064), .ZN(n9712) );
  AND2_X1 U5999 ( .A1(n7624), .A2(n7625), .ZN(n9714) );
  INV_X1 U6001 ( .A(n4960), .ZN(n5446) );
  INV_X1 U6002 ( .A(n4500), .ZN(n9281) );
  NOR3_X1 U6003 ( .A1(n9502), .A2(n8848), .A3(n4498), .ZN(n4500) );
  AND2_X1 U6004 ( .A1(n4671), .A2(n6422), .ZN(n4402) );
  INV_X1 U6005 ( .A(n9920), .ZN(n6446) );
  AND2_X1 U6006 ( .A1(n8022), .A2(n7845), .ZN(n8512) );
  INV_X1 U6007 ( .A(n8512), .ZN(n8608) );
  INV_X1 U6008 ( .A(n8481), .ZN(n8530) );
  NAND2_X1 U6009 ( .A1(n6051), .A2(n6050), .ZN(n8481) );
  AND2_X1 U6010 ( .A1(n9913), .A2(n6109), .ZN(n9456) );
  INV_X1 U6011 ( .A(n9456), .ZN(n9996) );
  INV_X1 U6012 ( .A(n5902), .ZN(n4521) );
  INV_X1 U6013 ( .A(n6726), .ZN(n7783) );
  NAND2_X1 U6014 ( .A1(n4798), .A2(n7975), .ZN(n4466) );
  NAND2_X1 U6015 ( .A1(n6703), .A2(n7839), .ZN(n4600) );
  NAND2_X1 U6016 ( .A1(n7933), .A2(n4481), .ZN(n4480) );
  OR2_X1 U6017 ( .A1(n7918), .A2(n7917), .ZN(n7914) );
  NAND2_X1 U6018 ( .A1(n7891), .A2(n7895), .ZN(n7894) );
  AOI21_X1 U6019 ( .B1(n7897), .B2(n4475), .A(n4474), .ZN(n7906) );
  OAI21_X1 U6020 ( .B1(n7953), .B2(n4486), .A(n4485), .ZN(n4403) );
  NAND2_X1 U6021 ( .A1(n4819), .A2(n7975), .ZN(n4818) );
  NOR3_X2 U6022 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .A3(
        P1_IR_REG_8__SCAN_IN), .ZN(n4639) );
  INV_X1 U6023 ( .A(n4901), .ZN(n4900) );
  NAND2_X1 U6024 ( .A1(n4549), .A2(n7662), .ZN(n9177) );
  INV_X1 U6025 ( .A(n6930), .ZN(n4416) );
  NAND2_X1 U6026 ( .A1(n4881), .A2(n4880), .ZN(n4883) );
  INV_X1 U6027 ( .A(n5562), .ZN(n7525) );
  NAND4_X2 U6028 ( .A1(n4910), .A2(n4909), .A3(n4911), .A4(n4912), .ZN(n5562)
         );
  NOR2_X2 U6029 ( .A1(n9257), .A2(n9256), .ZN(n9255) );
  AOI21_X2 U6030 ( .B1(n9130), .B2(n7683), .A(n7684), .ZN(n9120) );
  NAND2_X1 U6031 ( .A1(n4762), .A2(n4761), .ZN(n7021) );
  NAND2_X1 U6032 ( .A1(n8265), .A2(n8481), .ZN(n4770) );
  NAND2_X1 U6033 ( .A1(n5355), .A2(n5354), .ZN(n5370) );
  INV_X1 U6034 ( .A(n4784), .ZN(n4783) );
  NOR2_X1 U6035 ( .A1(n6355), .A2(n4767), .ZN(n6358) );
  NOR2_X1 U6036 ( .A1(n6327), .A2(n4753), .ZN(n6266) );
  XNOR2_X1 U6037 ( .A(n8256), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8263) );
  OAI21_X2 U6038 ( .B1(n5709), .B2(n4836), .A(n4834), .ZN(n5724) );
  INV_X1 U6039 ( .A(n8395), .ZN(n7824) );
  NAND3_X1 U6040 ( .A1(n7711), .A2(n7712), .A3(n7772), .ZN(n4410) );
  INV_X2 U6041 ( .A(n6922), .ZN(n9837) );
  AND2_X2 U6042 ( .A1(n7764), .A2(n7602), .ZN(n5518) );
  AOI21_X2 U6043 ( .B1(n5727), .B2(n8948), .A(n5726), .ZN(n8858) );
  NAND2_X2 U6044 ( .A1(n5510), .A2(n6726), .ZN(n5550) );
  NAND2_X1 U6045 ( .A1(n5033), .A2(n5032), .ZN(n4574) );
  NAND2_X2 U6046 ( .A1(n9008), .A2(n9837), .ZN(n7764) );
  INV_X1 U6047 ( .A(n9200), .ZN(n4549) );
  NAND2_X1 U6048 ( .A1(n7205), .A2(n7620), .ZN(n9273) );
  NAND2_X1 U6049 ( .A1(n4945), .A2(n4944), .ZN(n4949) );
  NAND2_X1 U6050 ( .A1(n4987), .A2(n4986), .ZN(n4417) );
  NAND2_X1 U6051 ( .A1(n4967), .A2(n4966), .ZN(n4418) );
  NAND2_X1 U6052 ( .A1(n8153), .A2(n4382), .ZN(n4419) );
  OAI211_X1 U6053 ( .C1(n8153), .C2(n4420), .A(n4419), .B(n4428), .ZN(P2_U3216) );
  NAND2_X1 U6054 ( .A1(n8153), .A2(n8152), .ZN(n8151) );
  OAI21_X1 U6055 ( .B1(n8153), .B2(n7475), .A(n4425), .ZN(n7811) );
  OR2_X1 U6056 ( .A1(n8095), .A2(n4436), .ZN(n4431) );
  NAND2_X1 U6057 ( .A1(n4433), .A2(n4431), .ZN(n4430) );
  NAND2_X2 U6058 ( .A1(n4574), .A2(n5036), .ZN(n5052) );
  NAND2_X1 U6059 ( .A1(n8432), .A2(n4449), .ZN(n4447) );
  NAND2_X1 U6060 ( .A1(n4458), .A2(n4457), .ZN(n6795) );
  NAND2_X1 U6061 ( .A1(n6638), .A2(n4712), .ZN(n4458) );
  OR2_X1 U6062 ( .A1(n6208), .A2(n6790), .ZN(n4462) );
  XNOR2_X1 U6063 ( .A(n5012), .B(n5011), .ZN(n6208) );
  NAND3_X1 U6064 ( .A1(n6632), .A2(n6631), .A3(n7996), .ZN(n4463) );
  NAND2_X1 U6065 ( .A1(n4464), .A2(n7987), .ZN(n7935) );
  NAND2_X1 U6066 ( .A1(n4466), .A2(n4465), .ZN(n7934) );
  NAND2_X1 U6067 ( .A1(n4468), .A2(n7866), .ZN(n4467) );
  INV_X1 U6068 ( .A(n4472), .ZN(n4468) );
  NAND2_X1 U6069 ( .A1(n4470), .A2(n7975), .ZN(n4469) );
  NAND4_X1 U6070 ( .A1(n4472), .A2(n7875), .A3(n4471), .A4(n7858), .ZN(n4470)
         );
  NAND2_X1 U6071 ( .A1(n7872), .A2(n4777), .ZN(n4471) );
  NAND2_X1 U6072 ( .A1(n7872), .A2(n4473), .ZN(n4472) );
  NAND3_X1 U6073 ( .A1(n7883), .A2(n7882), .A3(n8001), .ZN(n4478) );
  NAND3_X1 U6074 ( .A1(n4483), .A2(n4480), .A3(n7939), .ZN(n4479) );
  NAND3_X1 U6075 ( .A1(n9527), .A2(n4499), .A3(n4497), .ZN(n4496) );
  NAND2_X1 U6076 ( .A1(n9100), .A2(n9089), .ZN(n9084) );
  AND2_X1 U6077 ( .A1(n9100), .A2(n4507), .ZN(n9065) );
  NAND2_X1 U6078 ( .A1(n9100), .A2(n4508), .ZN(n9064) );
  OAI211_X2 U6079 ( .C1(n4919), .C2(n4908), .A(n4516), .B(n4515), .ZN(n7524)
         );
  AND2_X2 U6080 ( .A1(n4919), .A2(n7501), .ZN(n4992) );
  NAND3_X1 U6081 ( .A1(n4374), .A2(n4833), .A3(n4334), .ZN(n4643) );
  MUX2_X1 U6082 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n5847), .S(n9018), .Z(n9019)
         );
  XNOR2_X2 U6083 ( .A(n4951), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9018) );
  INV_X1 U6084 ( .A(n6613), .ZN(n4529) );
  INV_X1 U6085 ( .A(n4532), .ZN(n8609) );
  NAND3_X1 U6086 ( .A1(n4536), .A2(n6534), .A3(n9936), .ZN(n6612) );
  NAND3_X2 U6087 ( .A1(n6107), .A2(n6106), .A3(n4852), .ZN(n9920) );
  INV_X1 U6088 ( .A(n4540), .ZN(n8419) );
  NAND2_X1 U6089 ( .A1(n8356), .A2(n4541), .ZN(n8269) );
  NAND2_X1 U6090 ( .A1(n8356), .A2(n8341), .ZN(n8336) );
  NOR2_X2 U6091 ( .A1(n8336), .A2(n4544), .ZN(n8307) );
  NAND2_X1 U6092 ( .A1(n6916), .A2(n4548), .ZN(n9726) );
  NAND2_X1 U6093 ( .A1(n9726), .A2(n7625), .ZN(n6930) );
  NAND2_X1 U6094 ( .A1(n7207), .A2(n5523), .ZN(n7205) );
  NAND2_X1 U6095 ( .A1(n9120), .A2(n4560), .ZN(n4558) );
  NOR2_X1 U6096 ( .A1(n4552), .A2(n4551), .ZN(n9078) );
  NOR2_X1 U6097 ( .A1(n9120), .A2(n5528), .ZN(n9107) );
  NAND2_X1 U6098 ( .A1(n9255), .A2(n7657), .ZN(n4563) );
  OAI21_X1 U6099 ( .B1(n7151), .B2(n4584), .A(n4581), .ZN(n7814) );
  OAI21_X2 U6100 ( .B1(n4589), .B2(n8397), .A(n4586), .ZN(n8322) );
  OAI21_X1 U6101 ( .B1(n6856), .B2(n6857), .A(n7895), .ZN(n4596) );
  AND2_X1 U6102 ( .A1(n6797), .A2(n7887), .ZN(n6856) );
  NAND2_X1 U6103 ( .A1(n8424), .A2(n7823), .ZN(n4597) );
  NAND2_X1 U6104 ( .A1(n4601), .A2(n4602), .ZN(n9221) );
  NAND2_X1 U6105 ( .A1(n9271), .A2(n4323), .ZN(n4601) );
  NAND2_X1 U6106 ( .A1(n4613), .A2(n4614), .ZN(n5171) );
  NAND2_X1 U6107 ( .A1(n9496), .A2(n5151), .ZN(n4613) );
  NAND2_X1 U6108 ( .A1(n9115), .A2(n9121), .ZN(n4632) );
  NAND2_X1 U6109 ( .A1(n9115), .A2(n4616), .ZN(n4615) );
  NAND2_X1 U6110 ( .A1(n9223), .A2(n4324), .ZN(n4633) );
  NAND2_X1 U6111 ( .A1(n4633), .A2(n4634), .ZN(n9174) );
  NAND2_X1 U6112 ( .A1(n9223), .A2(n5269), .ZN(n9206) );
  INV_X1 U6113 ( .A(n5294), .ZN(n4638) );
  NAND4_X1 U6114 ( .A1(n4639), .A2(n4845), .A3(n4972), .A4(n4920), .ZN(n5079)
         );
  NAND4_X1 U6115 ( .A1(n4845), .A2(n4398), .A3(n4972), .A4(n4920), .ZN(n5062)
         );
  INV_X1 U6116 ( .A(n5081), .ZN(n4640) );
  NOR2_X1 U6117 ( .A1(n5082), .A2(n4388), .ZN(n4641) );
  NOR2_X2 U6118 ( .A1(n5081), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5120) );
  NAND2_X1 U6119 ( .A1(n4314), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6048) );
  AND2_X2 U6120 ( .A1(n4651), .A2(n4650), .ZN(n8153) );
  NAND2_X1 U6121 ( .A1(n6702), .A2(n6701), .ZN(n6966) );
  INV_X1 U6122 ( .A(n6701), .ZN(n4663) );
  NAND2_X1 U6123 ( .A1(n6417), .A2(n4670), .ZN(n4669) );
  NAND3_X1 U6124 ( .A1(n5813), .A2(n4676), .A3(n6541), .ZN(n4675) );
  AND3_X1 U6125 ( .A1(n4677), .A2(n4387), .A3(n6472), .ZN(n6632) );
  NAND2_X1 U6126 ( .A1(n6469), .A2(n6525), .ZN(n4677) );
  NAND2_X1 U6127 ( .A1(n8488), .A2(n4682), .ZN(n4681) );
  NOR2_X1 U6128 ( .A1(n8408), .A2(n8294), .ZN(n4697) );
  NAND2_X1 U6129 ( .A1(n6795), .A2(n6843), .ZN(n4700) );
  NOR2_X1 U6130 ( .A1(n4701), .A2(n4705), .ZN(n8503) );
  INV_X1 U6131 ( .A(n4704), .ZN(n4701) );
  INV_X1 U6132 ( .A(n4711), .ZN(n4708) );
  INV_X1 U6133 ( .A(n8599), .ZN(n4710) );
  NAND2_X1 U6134 ( .A1(n7107), .A2(n4385), .ZN(n7147) );
  NAND2_X1 U6135 ( .A1(n7147), .A2(n4863), .ZN(n7148) );
  NAND2_X1 U6136 ( .A1(n7107), .A2(n7106), .ZN(n7108) );
  NAND2_X1 U6137 ( .A1(n9936), .A2(n8190), .ZN(n7869) );
  NAND3_X1 U6138 ( .A1(n4891), .A2(n6898), .A3(n4714), .ZN(n4797) );
  INV_X2 U6139 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6898) );
  NAND2_X1 U6140 ( .A1(n5256), .A2(n4317), .ZN(n4715) );
  OAI21_X1 U6141 ( .B1(n5256), .B2(n5255), .A(n5254), .ZN(n5272) );
  NAND2_X1 U6142 ( .A1(n5255), .A2(n5254), .ZN(n4725) );
  NAND2_X1 U6143 ( .A1(n5174), .A2(n4729), .ZN(n4726) );
  NAND2_X1 U6144 ( .A1(n4726), .A2(n4727), .ZN(n5233) );
  NAND2_X1 U6145 ( .A1(n5118), .A2(n5117), .ZN(n5137) );
  MUX2_X1 U6146 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6254), .S(n6271), .Z(n9404)
         );
  NAND2_X1 U6147 ( .A1(n6545), .A2(n4775), .ZN(n4774) );
  NAND2_X1 U6148 ( .A1(n4774), .A2(n4772), .ZN(n6640) );
  NAND3_X1 U6149 ( .A1(n5877), .A2(n4778), .A3(n5803), .ZN(n5891) );
  NOR2_X2 U6150 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5877) );
  NAND2_X1 U6151 ( .A1(n5893), .A2(n4779), .ZN(n5824) );
  AND2_X1 U6152 ( .A1(n5828), .A2(n4786), .ZN(n5920) );
  NAND2_X1 U6153 ( .A1(n4790), .A2(n4386), .ZN(n7842) );
  NAND2_X1 U6154 ( .A1(n7838), .A2(n4792), .ZN(n4790) );
  OAI21_X2 U6155 ( .B1(n8467), .B2(n7817), .A(n7820), .ZN(n8454) );
  OAI21_X2 U6156 ( .B1(n7111), .B2(n7110), .A(n7903), .ZN(n7150) );
  OAI21_X2 U6157 ( .B1(n6956), .B2(n6955), .A(n7899), .ZN(n7111) );
  AND2_X2 U6158 ( .A1(n4797), .A2(n4796), .ZN(n4895) );
  NAND3_X1 U6159 ( .A1(n4892), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4796) );
  INV_X8 U6160 ( .A(n4895), .ZN(n6103) );
  NAND3_X1 U6161 ( .A1(n7926), .A2(n7927), .A3(n8469), .ZN(n4800) );
  OAI21_X1 U6162 ( .B1(n7978), .B2(n7945), .A(n7952), .ZN(n4809) );
  NAND2_X1 U6163 ( .A1(n5075), .A2(n5074), .ZN(n5095) );
  OAI21_X1 U6164 ( .B1(n7894), .B2(n7893), .A(n4820), .ZN(n4819) );
  AND2_X1 U6165 ( .A1(n7899), .A2(n7892), .ZN(n4820) );
  INV_X1 U6166 ( .A(n8858), .ZN(n4821) );
  OAI211_X2 U6167 ( .C1(n4824), .C2(n5731), .A(n4822), .B(n4363), .ZN(n5747)
         );
  NAND2_X1 U6168 ( .A1(n8858), .A2(n5732), .ZN(n4822) );
  NAND2_X1 U6169 ( .A1(n8857), .A2(n8860), .ZN(n4824) );
  NAND2_X1 U6170 ( .A1(n8843), .A2(n4383), .ZN(n4825) );
  NAND2_X1 U6171 ( .A1(n5120), .A2(n4833), .ZN(n5147) );
  NAND2_X1 U6172 ( .A1(n7220), .A2(n4384), .ZN(n7258) );
  NAND2_X1 U6173 ( .A1(n6820), .A2(n4844), .ZN(n4842) );
  NAND2_X1 U6174 ( .A1(n5480), .A2(n4848), .ZN(n4898) );
  NAND2_X1 U6175 ( .A1(n5480), .A2(n5482), .ZN(n5474) );
  INV_X1 U6176 ( .A(n5750), .ZN(n5760) );
  NAND2_X1 U6177 ( .A1(n9296), .A2(n9295), .ZN(n9364) );
  NAND2_X1 U6178 ( .A1(n9292), .A2(n9828), .ZN(n9296) );
  INV_X1 U6179 ( .A(n5977), .ZN(n8824) );
  NAND2_X1 U6180 ( .A1(n8967), .A2(n9805), .ZN(n7532) );
  INV_X1 U6181 ( .A(n6400), .ZN(n6398) );
  OAI211_X2 U6182 ( .C1(n6501), .C2(n6272), .A(n6124), .B(n6123), .ZN(n9929)
         );
  NAND2_X1 U6183 ( .A1(n9077), .A2(n7706), .ZN(n5530) );
  NAND2_X1 U6184 ( .A1(n4960), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4889) );
  INV_X1 U6185 ( .A(n9255), .ZN(n9259) );
  OAI21_X1 U6186 ( .B1(n9293), .B2(n9849), .A(n9508), .ZN(n9294) );
  NAND2_X1 U6187 ( .A1(n5515), .A2(n9766), .ZN(n9756) );
  NOR2_X2 U6188 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4920) );
  NAND2_X1 U6189 ( .A1(n5451), .A2(n5450), .ZN(n5455) );
  NAND4_X1 U6190 ( .A1(n6067), .A2(n6066), .A3(n6065), .A4(n6064), .ZN(n8192)
         );
  OAI21_X1 U6191 ( .B1(n6569), .B2(n9795), .A(n7525), .ZN(n4914) );
  NAND2_X1 U6192 ( .A1(n7887), .A2(n7893), .ZN(n6753) );
  NAND2_X2 U6193 ( .A1(n5647), .A2(n5646), .ZN(n8843) );
  NAND2_X1 U6194 ( .A1(n5724), .A2(n5723), .ZN(n8947) );
  INV_X1 U6195 ( .A(n5724), .ZN(n5718) );
  OAI222_X1 U6196 ( .A1(P2_U3152), .A2(n6736), .B1(n8835), .B2(n6791), .C1(
        n5912), .C2(n8827), .ZN(P2_U3348) );
  OAI222_X1 U6197 ( .A1(n9397), .A2(n6791), .B1(n6184), .B2(P1_U3084), .C1(
        n5908), .C2(n9401), .ZN(P1_U3343) );
  NAND2_X1 U6198 ( .A1(n4934), .A2(n8964), .ZN(n7526) );
  INV_X1 U6199 ( .A(n4934), .ZN(n4932) );
  XNOR2_X1 U6200 ( .A(n7495), .B(SI_30_), .ZN(n7829) );
  AND2_X1 U6201 ( .A1(n6092), .A2(n8043), .ZN(n9752) );
  NAND2_X2 U6202 ( .A1(n6383), .A2(n8437), .ZN(n9441) );
  OR2_X1 U6203 ( .A1(n6501), .A2(n6295), .ZN(n4851) );
  OR2_X1 U6204 ( .A1(n6501), .A2(n6271), .ZN(n4852) );
  INV_X1 U6205 ( .A(n7704), .ZN(n7582) );
  OR2_X1 U6206 ( .A1(n8952), .A2(n9147), .ZN(n4853) );
  OR2_X1 U6207 ( .A1(n9339), .A2(n8955), .ZN(n4854) );
  NOR2_X1 U6208 ( .A1(n7052), .A2(n7051), .ZN(n4855) );
  OR2_X1 U6209 ( .A1(n9164), .A2(n8882), .ZN(n4857) );
  AND4_X1 U6210 ( .A1(n7291), .A2(n7290), .A3(n7289), .A4(n7288), .ZN(n8098)
         );
  AND2_X1 U6211 ( .A1(n5096), .A2(n5078), .ZN(n4858) );
  AND2_X1 U6212 ( .A1(n5173), .A2(n5159), .ZN(n4859) );
  INV_X1 U6213 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4875) );
  NAND2_X1 U6214 ( .A1(n9010), .A2(n9813), .ZN(n5515) );
  INV_X1 U6215 ( .A(n8977), .ZN(n8988) );
  INV_X1 U6216 ( .A(n7651), .ZN(n5525) );
  INV_X1 U6217 ( .A(n8594), .ZN(n8285) );
  XOR2_X1 U6218 ( .A(n8408), .B(n7798), .Z(n4861) );
  INV_X1 U6219 ( .A(n8345), .ZN(n8300) );
  AND2_X1 U6220 ( .A1(n7488), .A2(n7487), .ZN(n8345) );
  AND2_X1 U6221 ( .A1(n6436), .A2(n6388), .ZN(n4862) );
  INV_X1 U6222 ( .A(n8871), .ZN(n5694) );
  OR2_X2 U6223 ( .A1(n5872), .A2(P1_U3084), .ZN(n9011) );
  INV_X1 U6224 ( .A(n5841), .ZN(n5554) );
  INV_X1 U6225 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5809) );
  INV_X1 U6226 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5808) );
  OR2_X1 U6227 ( .A1(n8172), .A2(n7836), .ZN(n7837) );
  INV_X1 U6228 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n4871) );
  INV_X1 U6229 ( .A(n8106), .ZN(n7445) );
  NOR2_X1 U6230 ( .A1(n5811), .A2(n5810), .ZN(n5812) );
  NAND2_X1 U6231 ( .A1(n9490), .A2(n7226), .ZN(n5124) );
  NAND2_X1 U6232 ( .A1(n7446), .A2(n7445), .ZN(n7447) );
  INV_X1 U6233 ( .A(n7392), .ZN(n5972) );
  AOI22_X1 U6234 ( .A1(n6565), .A2(n4311), .B1(n5554), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U6235 ( .A1(n7771), .A2(n7582), .ZN(n7583) );
  AND2_X1 U6236 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5966) );
  NAND2_X1 U6237 ( .A1(n5972), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7405) );
  NAND2_X1 U6238 ( .A1(n4545), .A2(n8345), .ZN(n8301) );
  INV_X1 U6239 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8712) );
  INV_X1 U6240 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5827) );
  NAND2_X1 U6241 ( .A1(n5556), .A2(n5555), .ZN(n5987) );
  NAND2_X1 U6242 ( .A1(n7584), .A2(n7583), .ZN(n7712) );
  OR2_X1 U6243 ( .A1(n5164), .A2(n5163), .ZN(n5180) );
  OR2_X1 U6244 ( .A1(n5067), .A2(n5066), .ZN(n5089) );
  INV_X1 U6245 ( .A(n9714), .ZN(n5064) );
  INV_X1 U6246 ( .A(SI_20_), .ZN(n5298) );
  INV_X1 U6247 ( .A(SI_16_), .ZN(n8628) );
  INV_X1 U6248 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4867) );
  INV_X1 U6249 ( .A(n7183), .ZN(n7179) );
  INV_X1 U6250 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6849) );
  INV_X1 U6251 ( .A(n7242), .ZN(n5970) );
  INV_X1 U6252 ( .A(n7053), .ZN(n7054) );
  OR2_X1 U6253 ( .A1(n7286), .A2(n8224), .ZN(n7293) );
  OR2_X1 U6254 ( .A1(n7435), .A2(n8712), .ZN(n7437) );
  INV_X1 U6255 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8224) );
  AND2_X1 U6256 ( .A1(n7481), .A2(n7480), .ZN(n8320) );
  INV_X1 U6257 ( .A(n8439), .ZN(n8450) );
  INV_X1 U6258 ( .A(n8172), .ZN(n8272) );
  INV_X1 U6259 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8698) );
  NOR2_X1 U6260 ( .A1(n7913), .A2(n8178), .ZN(n7234) );
  NAND2_X1 U6261 ( .A1(n6757), .A2(n9973), .ZN(n6813) );
  NAND2_X1 U6262 ( .A1(n9456), .A2(n8530), .ZN(n8525) );
  INV_X1 U6263 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5836) );
  INV_X1 U6264 ( .A(n7261), .ZN(n5636) );
  INV_X1 U6265 ( .A(n5224), .ZN(n5223) );
  INV_X1 U6266 ( .A(n5306), .ZN(n5304) );
  INV_X1 U6267 ( .A(n6122), .ZN(n4927) );
  AND2_X1 U6268 ( .A1(n5758), .A2(n6099), .ZN(n5769) );
  INV_X1 U6269 ( .A(n7595), .ZN(n5021) );
  INV_X1 U6270 ( .A(n7750), .ZN(n5529) );
  AND2_X1 U6271 ( .A1(n7526), .A2(n7528), .ZN(n7723) );
  AND2_X1 U6272 ( .A1(n5486), .A2(n5485), .ZN(n5487) );
  INV_X1 U6273 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5238) );
  INV_X1 U6274 ( .A(SI_9_), .ZN(n8624) );
  OR2_X1 U6275 ( .A1(n4304), .A2(n8832), .ZN(n7333) );
  OR2_X1 U6276 ( .A1(n7374), .A2(n7373), .ZN(n7392) );
  OR2_X1 U6277 ( .A1(n6850), .A2(n6849), .ZN(n6949) );
  NOR2_X1 U6278 ( .A1(n4855), .A2(n7054), .ZN(n7055) );
  OR2_X1 U6279 ( .A1(n6800), .A2(n8197), .ZN(n6850) );
  NAND2_X1 U6280 ( .A1(n5971), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7374) );
  AND2_X1 U6281 ( .A1(n8027), .A2(n8020), .ZN(n6157) );
  INV_X1 U6282 ( .A(n6157), .ZN(n6385) );
  INV_X1 U6283 ( .A(n7832), .ZN(n7485) );
  INV_X1 U6284 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8197) );
  INV_X1 U6285 ( .A(n8455), .ZN(n8605) );
  NAND2_X1 U6286 ( .A1(n4862), .A2(n6396), .ZN(n6525) );
  INV_X1 U6287 ( .A(n8836), .ZN(n6030) );
  OR2_X1 U6288 ( .A1(n5288), .A2(n5287), .ZN(n5306) );
  AND2_X1 U6289 ( .A1(n5780), .A2(n5779), .ZN(n5792) );
  INV_X1 U6290 ( .A(n9182), .ZN(n8882) );
  OR2_X1 U6291 ( .A1(n5393), .A2(n5392), .ZN(n5412) );
  OR2_X1 U6292 ( .A1(n5244), .A2(n5243), .ZN(n5263) );
  OR2_X1 U6293 ( .A1(n5771), .A2(n6229), .ZN(n8953) );
  OR2_X1 U6294 ( .A1(n5771), .A2(n5532), .ZN(n8994) );
  NOR2_X1 U6295 ( .A1(n5859), .A2(n9392), .ZN(n9052) );
  AND2_X1 U6296 ( .A1(n7661), .A2(n7665), .ZN(n9222) );
  INV_X1 U6297 ( .A(n9136), .ZN(n9745) );
  AND2_X1 U6298 ( .A1(n6093), .A2(n6726), .ZN(n9828) );
  OR2_X1 U6299 ( .A1(n7756), .A2(n6229), .ZN(n9772) );
  AND2_X1 U6300 ( .A1(n6088), .A2(n6087), .ZN(n6090) );
  INV_X1 U6301 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5282) );
  AND2_X1 U6302 ( .A1(n5232), .A2(n5216), .ZN(n5230) );
  INV_X1 U6303 ( .A(n8145), .ZN(n8154) );
  AND2_X1 U6304 ( .A1(n7459), .A2(n7458), .ZN(n8173) );
  AND4_X1 U6305 ( .A1(n6954), .A2(n6953), .A3(n6952), .A4(n6951), .ZN(n8179)
         );
  AND2_X1 U6306 ( .A1(n6267), .A2(n6052), .ZN(n9895) );
  INV_X1 U6307 ( .A(n9895), .ZN(n8234) );
  INV_X1 U6308 ( .A(n6753), .ZN(n7999) );
  AND2_X1 U6309 ( .A1(n8192), .A2(n9914), .ZN(n6437) );
  AOI21_X1 U6310 ( .B1(n9903), .B2(n9907), .A(n9908), .ZN(n8529) );
  INV_X1 U6311 ( .A(n10001), .ZN(n9924) );
  AND2_X1 U6312 ( .A1(n6749), .A2(n6639), .ZN(n9970) );
  NAND2_X1 U6313 ( .A1(n8533), .A2(n9471), .ZN(n10001) );
  INV_X1 U6314 ( .A(n8953), .ZN(n8992) );
  NOR2_X2 U6315 ( .A1(n5764), .A2(n5759), .ZN(n8977) );
  OR2_X1 U6316 ( .A1(n5766), .A2(n5984), .ZN(n5761) );
  AND3_X1 U6317 ( .A1(n5463), .A2(n5462), .A3(n5461), .ZN(n8050) );
  AND4_X1 U6318 ( .A1(n5324), .A2(n5323), .A3(n5322), .A4(n5321), .ZN(n8955)
         );
  AND4_X1 U6319 ( .A1(n5229), .A2(n5228), .A3(n5227), .A4(n5226), .ZN(n5668)
         );
  INV_X1 U6320 ( .A(n9698), .ZN(n9665) );
  NOR2_X1 U6321 ( .A1(n5855), .A2(n5532), .ZN(n9698) );
  INV_X1 U6322 ( .A(n9702), .ZN(n9671) );
  NOR2_X1 U6323 ( .A1(P1_U3083), .A2(n5873), .ZN(n9603) );
  INV_X1 U6324 ( .A(n9512), .ZN(n9066) );
  AND2_X1 U6325 ( .A1(n7720), .A2(n7719), .ZN(n9129) );
  AND2_X1 U6326 ( .A1(n5753), .A2(n6229), .ZN(n9489) );
  INV_X1 U6327 ( .A(n9283), .ZN(n9783) );
  AND2_X1 U6328 ( .A1(n9779), .A2(n6570), .ZN(n9764) );
  AND2_X1 U6329 ( .A1(n5757), .A2(n9380), .ZN(n6099) );
  INV_X1 U6330 ( .A(n9294), .ZN(n9295) );
  INV_X1 U6331 ( .A(n9514), .ZN(n9855) );
  AND2_X1 U6332 ( .A1(n5500), .A2(n5499), .ZN(n6091) );
  AND2_X1 U6333 ( .A1(n5257), .A2(n5240), .ZN(n9039) );
  AND2_X1 U6334 ( .A1(n4999), .A2(n4998), .ZN(n9599) );
  INV_X1 U6335 ( .A(n9401), .ZN(n9390) );
  NAND2_X1 U6336 ( .A1(n5942), .A2(n5941), .ZN(n9898) );
  NAND2_X1 U6337 ( .A1(n6163), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9891) );
  INV_X1 U6338 ( .A(n9886), .ZN(n8161) );
  INV_X1 U6339 ( .A(n8173), .ZN(n8365) );
  INV_X1 U6340 ( .A(n8098), .ZN(n8604) );
  INV_X1 U6341 ( .A(n6719), .ZN(n8185) );
  INV_X1 U6342 ( .A(n9897), .ZN(n9414) );
  INV_X1 U6343 ( .A(n8494), .ZN(n8443) );
  OR2_X1 U6344 ( .A1(n4305), .A2(n6558), .ZN(n8487) );
  NAND2_X1 U6345 ( .A1(n9441), .A2(n6386), .ZN(n9444) );
  INV_X1 U6346 ( .A(n10023), .ZN(n10021) );
  INV_X1 U6347 ( .A(n10004), .ZN(n10002) );
  AND2_X2 U6348 ( .A1(n8614), .A2(n8613), .ZN(n10004) );
  NOR2_X1 U6349 ( .A1(n9904), .A2(n9903), .ZN(n9906) );
  INV_X1 U6350 ( .A(n9906), .ZN(n9909) );
  INV_X1 U6351 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n5954) );
  OR2_X1 U6352 ( .A1(n5859), .A2(n4307), .ZN(n9569) );
  INV_X1 U6353 ( .A(n9317), .ZN(n9119) );
  INV_X1 U6354 ( .A(n9332), .ZN(n9164) );
  AND2_X1 U6355 ( .A1(n5761), .A2(n9283), .ZN(n9000) );
  INV_X1 U6356 ( .A(n5796), .ZN(n9122) );
  INV_X1 U6357 ( .A(n8911), .ZN(n9248) );
  INV_X1 U6358 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n8626) );
  OR2_X1 U6359 ( .A1(n5859), .A2(n5858), .ZN(n9708) );
  INV_X1 U6360 ( .A(n9603), .ZN(n9711) );
  NAND2_X1 U6361 ( .A1(n9779), .A2(n9752), .ZN(n9290) );
  NAND2_X1 U6362 ( .A1(n5542), .A2(n9283), .ZN(n9779) );
  INV_X1 U6363 ( .A(n9879), .ZN(n9876) );
  INV_X1 U6364 ( .A(n9859), .ZN(n9857) );
  AND2_X2 U6365 ( .A1(n6100), .A2(n6091), .ZN(n9859) );
  OR2_X1 U6366 ( .A1(n9791), .A2(n9379), .ZN(n9789) );
  INV_X1 U6367 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9394) );
  INV_X1 U6368 ( .A(n9659), .ZN(n9045) );
  INV_X1 U6369 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5943) );
  NOR2_X1 U6370 ( .A1(n10052), .A2(n10051), .ZN(n10050) );
  INV_X2 U6371 ( .A(n8175), .ZN(P2_U3966) );
  INV_X1 U6372 ( .A(n9011), .ZN(P1_U4006) );
  INV_X1 U6373 ( .A(n5079), .ZN(n4870) );
  NAND2_X1 U6374 ( .A1(n4870), .A2(n4869), .ZN(n5081) );
  NOR2_X1 U6375 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n4874) );
  NOR2_X1 U6376 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4873) );
  NOR2_X1 U6377 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4872) );
  NAND2_X1 U6378 ( .A1(n4900), .A2(n4875), .ZN(n4882) );
  XNOR2_X2 U6379 ( .A(n4877), .B(n4876), .ZN(n7331) );
  OR2_X1 U6380 ( .A1(n4900), .A2(n4878), .ZN(n4879) );
  NAND2_X1 U6381 ( .A1(n4879), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n4881) );
  INV_X1 U6382 ( .A(n5006), .ZN(n4884) );
  INV_X1 U6383 ( .A(n7331), .ZN(n4885) );
  AND2_X2 U6384 ( .A1(n4885), .A2(n9385), .ZN(n4960) );
  AND2_X2 U6385 ( .A1(n4886), .A2(n4885), .ZN(n4937) );
  NAND2_X1 U6386 ( .A1(n4939), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4887) );
  NAND4_X2 U6387 ( .A1(n4890), .A2(n4889), .A3(n4888), .A4(n4887), .ZN(n5553)
         );
  INV_X1 U6388 ( .A(SI_0_), .ZN(n4894) );
  INV_X1 U6389 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n4893) );
  OAI21_X1 U6390 ( .B1(n7501), .B2(n4894), .A(n4893), .ZN(n4897) );
  AND2_X1 U6391 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4896) );
  AND2_X1 U6392 ( .A1(n4906), .A2(n4897), .ZN(n9402) );
  NAND2_X1 U6393 ( .A1(n4898), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4899) );
  NAND2_X2 U6394 ( .A1(n4902), .A2(n4901), .ZN(n5532) );
  NAND2_X1 U6395 ( .A1(n4373), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4903) );
  NAND2_X2 U6396 ( .A1(n4898), .A2(n4904), .ZN(n7492) );
  MUX2_X1 U6397 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9402), .S(n4919), .Z(n6565) );
  AND2_X1 U6398 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4905) );
  NAND2_X1 U6399 ( .A1(n7501), .A2(n4905), .ZN(n6061) );
  MUX2_X1 U6400 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n6103), .Z(n4921) );
  XNOR2_X1 U6401 ( .A(n4922), .B(n4921), .ZN(n5882) );
  NAND2_X1 U6402 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4907) );
  XNOR2_X1 U6403 ( .A(n4907), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9577) );
  INV_X1 U6404 ( .A(n9577), .ZN(n4908) );
  NAND2_X1 U6405 ( .A1(n4937), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4912) );
  NAND2_X1 U6406 ( .A1(n4960), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4911) );
  NAND2_X1 U6407 ( .A1(n5246), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4910) );
  NAND2_X1 U6408 ( .A1(n4939), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4909) );
  NAND2_X1 U6409 ( .A1(n6569), .A2(n9795), .ZN(n4913) );
  NAND2_X1 U6410 ( .A1(n4914), .A2(n4913), .ZN(n6669) );
  NAND2_X1 U6411 ( .A1(n4937), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n4918) );
  NAND2_X1 U6412 ( .A1(n4960), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4917) );
  NAND2_X1 U6413 ( .A1(n4939), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4916) );
  NAND2_X1 U6414 ( .A1(n5246), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n4915) );
  AND4_X2 U6415 ( .A1(n4918), .A2(n4917), .A3(n4916), .A4(n4915), .ZN(n4934)
         );
  INV_X1 U6416 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4950) );
  NAND2_X1 U6417 ( .A1(n4307), .A2(n9018), .ZN(n4930) );
  NAND2_X1 U6418 ( .A1(n4992), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4929) );
  NAND2_X1 U6419 ( .A1(n4923), .A2(SI_1_), .ZN(n4924) );
  INV_X1 U6420 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6121) );
  INV_X1 U6421 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4925) );
  XNOR2_X1 U6422 ( .A(n4946), .B(SI_2_), .ZN(n4944) );
  XNOR2_X1 U6423 ( .A(n4945), .B(n4944), .ZN(n6122) );
  NAND2_X1 U6424 ( .A1(n7528), .A2(n7526), .ZN(n4933) );
  NAND2_X1 U6425 ( .A1(n6669), .A2(n4933), .ZN(n4936) );
  NAND2_X1 U6426 ( .A1(n4934), .A2(n4931), .ZN(n4935) );
  NAND2_X1 U6427 ( .A1(n4936), .A2(n4935), .ZN(n6681) );
  INV_X1 U6428 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n4938) );
  NAND2_X1 U6429 ( .A1(n4937), .A2(n4938), .ZN(n4943) );
  NAND2_X1 U6430 ( .A1(n7507), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4942) );
  NAND2_X1 U6431 ( .A1(n4960), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4941) );
  NAND2_X1 U6432 ( .A1(n5246), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n4940) );
  INV_X1 U6433 ( .A(n4956), .ZN(n8967) );
  INV_X1 U6434 ( .A(n4946), .ZN(n4947) );
  NAND2_X1 U6435 ( .A1(n4947), .A2(SI_2_), .ZN(n4948) );
  NAND2_X1 U6436 ( .A1(n4949), .A2(n4948), .ZN(n4967) );
  INV_X1 U6437 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5889) );
  MUX2_X1 U6438 ( .A(n6135), .B(n5889), .S(n6103), .Z(n4968) );
  XNOR2_X1 U6439 ( .A(n4968), .B(SI_3_), .ZN(n4966) );
  XNOR2_X1 U6440 ( .A(n4967), .B(n4966), .ZN(n6134) );
  NAND2_X1 U6441 ( .A1(n4992), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4955) );
  NAND2_X1 U6442 ( .A1(n4951), .A2(n4950), .ZN(n4952) );
  NAND2_X1 U6443 ( .A1(n4952), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4953) );
  XNOR2_X1 U6444 ( .A(n4953), .B(P1_IR_REG_3__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U6445 ( .A1(n4307), .A2(n5888), .ZN(n4954) );
  INV_X1 U6446 ( .A(n6692), .ZN(n9805) );
  NAND2_X1 U6447 ( .A1(n4956), .A2(n6692), .ZN(n7727) );
  NAND2_X1 U6448 ( .A1(n7532), .A2(n7727), .ZN(n5513) );
  NAND2_X1 U6449 ( .A1(n6681), .A2(n5513), .ZN(n4958) );
  NAND2_X1 U6450 ( .A1(n4956), .A2(n9805), .ZN(n4957) );
  NAND2_X1 U6451 ( .A1(n4958), .A2(n4957), .ZN(n9757) );
  INV_X1 U6452 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n4959) );
  XNOR2_X1 U6453 ( .A(n4959), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n9782) );
  NAND2_X1 U6454 ( .A1(n4937), .A2(n9782), .ZN(n4965) );
  NAND2_X1 U6455 ( .A1(n7507), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n4964) );
  INV_X1 U6456 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n4961) );
  NAND2_X1 U6457 ( .A1(n5246), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n4962) );
  INV_X1 U6458 ( .A(n9748), .ZN(n9010) );
  INV_X1 U6459 ( .A(n4968), .ZN(n4969) );
  NAND2_X1 U6460 ( .A1(n4969), .A2(SI_3_), .ZN(n4970) );
  INV_X1 U6461 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n4971) );
  MUX2_X1 U6462 ( .A(n6150), .B(n4971), .S(n6103), .Z(n4988) );
  XNOR2_X1 U6463 ( .A(n4988), .B(SI_4_), .ZN(n4986) );
  XNOR2_X1 U6464 ( .A(n4987), .B(n4986), .ZN(n6149) );
  NAND2_X1 U6465 ( .A1(n4992), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U6466 ( .A1(n4994), .A2(n4972), .ZN(n4973) );
  NAND2_X1 U6467 ( .A1(n4973), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4974) );
  XNOR2_X1 U6468 ( .A(n4974), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U6469 ( .A1(n4307), .A2(n6242), .ZN(n4975) );
  INV_X1 U6470 ( .A(n9758), .ZN(n9813) );
  NAND2_X1 U6471 ( .A1(n9748), .A2(n9758), .ZN(n9766) );
  NAND2_X1 U6472 ( .A1(n9757), .A2(n9756), .ZN(n4978) );
  NAND2_X1 U6473 ( .A1(n9748), .A2(n9813), .ZN(n4977) );
  NAND2_X1 U6474 ( .A1(n4978), .A2(n4977), .ZN(n9737) );
  NAND2_X1 U6475 ( .A1(n7507), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4985) );
  NAND3_X1 U6476 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5004) );
  INV_X1 U6477 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n4980) );
  NAND2_X1 U6478 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n4979) );
  NAND2_X1 U6479 ( .A1(n4980), .A2(n4979), .ZN(n4981) );
  AND2_X1 U6480 ( .A1(n5004), .A2(n4981), .ZN(n9741) );
  NAND2_X1 U6481 ( .A1(n4937), .A2(n9741), .ZN(n4984) );
  NAND2_X1 U6482 ( .A1(n4960), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4983) );
  NAND2_X1 U6483 ( .A1(n4884), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n4982) );
  INV_X1 U6484 ( .A(n4988), .ZN(n4989) );
  NAND2_X1 U6485 ( .A1(n4989), .A2(SI_4_), .ZN(n4990) );
  INV_X1 U6486 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n4991) );
  MUX2_X1 U6487 ( .A(n6209), .B(n4991), .S(n6103), .Z(n5013) );
  XNOR2_X1 U6488 ( .A(n5013), .B(SI_5_), .ZN(n5011) );
  NAND2_X1 U6489 ( .A1(n5407), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5001) );
  NAND2_X1 U6490 ( .A1(n4994), .A2(n4993), .ZN(n4995) );
  NAND2_X1 U6491 ( .A1(n4995), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4996) );
  MUX2_X1 U6492 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4996), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n4999) );
  INV_X1 U6493 ( .A(n4997), .ZN(n4998) );
  NAND2_X1 U6494 ( .A1(n4307), .A2(n9599), .ZN(n5000) );
  NAND2_X1 U6495 ( .A1(n9773), .A2(n9739), .ZN(n7588) );
  INV_X1 U6496 ( .A(n9739), .ZN(n9821) );
  NAND2_X1 U6497 ( .A1(n9009), .A2(n9821), .ZN(n7590) );
  NAND2_X1 U6498 ( .A1(n9009), .A2(n9739), .ZN(n5002) );
  INV_X1 U6499 ( .A(n6832), .ZN(n5022) );
  INV_X1 U6500 ( .A(n5004), .ZN(n5003) );
  NAND2_X1 U6501 ( .A1(n5003), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5026) );
  INV_X1 U6502 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6907) );
  NAND2_X1 U6503 ( .A1(n5004), .A2(n6907), .ZN(n5005) );
  AND2_X1 U6504 ( .A1(n5026), .A2(n5005), .ZN(n6912) );
  NAND2_X1 U6505 ( .A1(n4937), .A2(n6912), .ZN(n5010) );
  NAND2_X1 U6506 ( .A1(n7507), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5009) );
  NAND2_X1 U6507 ( .A1(n4960), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5008) );
  NAND2_X1 U6508 ( .A1(n4884), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5007) );
  NAND2_X1 U6509 ( .A1(n5012), .A2(n5011), .ZN(n5016) );
  INV_X1 U6510 ( .A(n5013), .ZN(n5014) );
  NAND2_X1 U6511 ( .A1(n5014), .A2(SI_5_), .ZN(n5015) );
  INV_X1 U6512 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5017) );
  MUX2_X1 U6513 ( .A(n6407), .B(n5017), .S(n6103), .Z(n5034) );
  XNOR2_X1 U6514 ( .A(n5034), .B(SI_6_), .ZN(n5032) );
  XNOR2_X1 U6515 ( .A(n5033), .B(n5032), .ZN(n6406) );
  NAND2_X1 U6516 ( .A1(n5407), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5020) );
  OR2_X1 U6517 ( .A1(n4997), .A2(n4878), .ZN(n5018) );
  XNOR2_X1 U6518 ( .A(n5018), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9602) );
  NAND2_X1 U6519 ( .A1(n4307), .A2(n9602), .ZN(n5019) );
  OAI211_X1 U6520 ( .C1(n5104), .C2(n6406), .A(n5020), .B(n5019), .ZN(n9826)
         );
  NAND2_X1 U6521 ( .A1(n6919), .A2(n9826), .ZN(n7729) );
  INV_X1 U6522 ( .A(n6919), .ZN(n9743) );
  INV_X1 U6523 ( .A(n9826), .ZN(n6909) );
  NAND2_X1 U6524 ( .A1(n9743), .A2(n6909), .ZN(n7757) );
  NAND2_X1 U6525 ( .A1(n5022), .A2(n5021), .ZN(n6830) );
  NAND2_X1 U6526 ( .A1(n6919), .A2(n6909), .ZN(n5023) );
  NAND2_X1 U6527 ( .A1(n6830), .A2(n5023), .ZN(n6915) );
  NAND2_X1 U6528 ( .A1(n7507), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5031) );
  INV_X1 U6529 ( .A(n5026), .ZN(n5024) );
  NAND2_X1 U6530 ( .A1(n5024), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5044) );
  INV_X1 U6531 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5025) );
  NAND2_X1 U6532 ( .A1(n5026), .A2(n5025), .ZN(n5027) );
  AND2_X1 U6533 ( .A1(n5044), .A2(n5027), .ZN(n6921) );
  NAND2_X1 U6534 ( .A1(n4937), .A2(n6921), .ZN(n5030) );
  NAND2_X1 U6535 ( .A1(n5535), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5029) );
  NAND2_X1 U6536 ( .A1(n4884), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5028) );
  INV_X1 U6537 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n8784) );
  INV_X1 U6538 ( .A(n5034), .ZN(n5035) );
  NAND2_X1 U6539 ( .A1(n5035), .A2(SI_6_), .ZN(n5036) );
  MUX2_X1 U6540 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6103), .Z(n5053) );
  XNOR2_X1 U6541 ( .A(n5053), .B(SI_7_), .ZN(n5050) );
  NAND2_X1 U6542 ( .A1(n7512), .A2(n6496), .ZN(n5040) );
  OR2_X1 U6543 ( .A1(n5037), .A2(n4878), .ZN(n5038) );
  XNOR2_X1 U6544 ( .A(n5038), .B(P1_IR_REG_7__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U6545 ( .A1(n4307), .A2(n5902), .ZN(n5039) );
  OAI211_X1 U6546 ( .C1(n5061), .C2(n8784), .A(n5040), .B(n5039), .ZN(n6922)
         );
  NAND2_X1 U6547 ( .A1(n9722), .A2(n6922), .ZN(n7602) );
  INV_X1 U6548 ( .A(n9722), .ZN(n9008) );
  NAND2_X1 U6549 ( .A1(n6915), .A2(n7594), .ZN(n5042) );
  NAND2_X1 U6550 ( .A1(n9722), .A2(n9837), .ZN(n5041) );
  NAND2_X1 U6551 ( .A1(n5042), .A2(n5041), .ZN(n9713) );
  NAND2_X1 U6552 ( .A1(n7507), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5049) );
  INV_X1 U6553 ( .A(n5044), .ZN(n5043) );
  NAND2_X1 U6554 ( .A1(n5043), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5067) );
  INV_X1 U6555 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6824) );
  NAND2_X1 U6556 ( .A1(n5044), .A2(n6824), .ZN(n5045) );
  AND2_X1 U6557 ( .A1(n5067), .A2(n5045), .ZN(n9732) );
  NAND2_X1 U6558 ( .A1(n5460), .A2(n9732), .ZN(n5048) );
  NAND2_X1 U6559 ( .A1(n5535), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5047) );
  NAND2_X1 U6560 ( .A1(n5246), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5046) );
  INV_X1 U6561 ( .A(n5050), .ZN(n5051) );
  NAND2_X1 U6562 ( .A1(n5053), .A2(SI_7_), .ZN(n5054) );
  INV_X1 U6563 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5906) );
  INV_X1 U6564 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5055) );
  MUX2_X1 U6565 ( .A(n5906), .B(n5055), .S(n6103), .Z(n5057) );
  INV_X1 U6566 ( .A(SI_8_), .ZN(n5056) );
  NAND2_X1 U6567 ( .A1(n5057), .A2(n5056), .ZN(n5074) );
  INV_X1 U6568 ( .A(n5057), .ZN(n5058) );
  NAND2_X1 U6569 ( .A1(n5058), .A2(SI_8_), .ZN(n5059) );
  NAND2_X1 U6570 ( .A1(n5074), .A2(n5059), .ZN(n5073) );
  INV_X1 U6571 ( .A(n5073), .ZN(n5060) );
  NAND2_X1 U6572 ( .A1(n5062), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5063) );
  XNOR2_X1 U6573 ( .A(n5063), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9624) );
  NAND2_X1 U6574 ( .A1(n7044), .A2(n6826), .ZN(n7624) );
  INV_X1 U6575 ( .A(n7044), .ZN(n9007) );
  NAND2_X1 U6576 ( .A1(n9007), .A2(n9842), .ZN(n7625) );
  NAND2_X1 U6577 ( .A1(n9007), .A2(n6826), .ZN(n5065) );
  NAND2_X1 U6578 ( .A1(n5067), .A2(n5066), .ZN(n5068) );
  AND2_X1 U6579 ( .A1(n5089), .A2(n5068), .ZN(n7041) );
  NAND2_X1 U6580 ( .A1(n5460), .A2(n7041), .ZN(n5072) );
  NAND2_X1 U6581 ( .A1(n7507), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5071) );
  NAND2_X1 U6582 ( .A1(n5535), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5070) );
  NAND2_X1 U6583 ( .A1(n5246), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5069) );
  MUX2_X1 U6584 ( .A(n5916), .B(n5907), .S(n6103), .Z(n5076) );
  NAND2_X1 U6585 ( .A1(n5076), .A2(n8624), .ZN(n5096) );
  INV_X1 U6586 ( .A(n5076), .ZN(n5077) );
  NAND2_X1 U6587 ( .A1(n5077), .A2(SI_9_), .ZN(n5078) );
  NAND2_X1 U6588 ( .A1(n7512), .A2(n6703), .ZN(n5086) );
  NAND2_X1 U6589 ( .A1(n5407), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n5085) );
  NAND2_X1 U6590 ( .A1(n5079), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5080) );
  MUX2_X1 U6591 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5080), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n5083) );
  AND2_X1 U6592 ( .A1(n5083), .A2(n5082), .ZN(n5998) );
  NAND2_X1 U6593 ( .A1(n4307), .A2(n5998), .ZN(n5084) );
  NAND2_X1 U6594 ( .A1(n9721), .A2(n9850), .ZN(n5087) );
  NAND2_X1 U6595 ( .A1(n5089), .A2(n5088), .ZN(n5090) );
  AND2_X1 U6596 ( .A1(n5108), .A2(n5090), .ZN(n7134) );
  NAND2_X1 U6597 ( .A1(n5460), .A2(n7134), .ZN(n5094) );
  NAND2_X1 U6598 ( .A1(n7507), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5093) );
  NAND2_X1 U6599 ( .A1(n5535), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5092) );
  NAND2_X1 U6600 ( .A1(n5246), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5091) );
  MUX2_X1 U6601 ( .A(n5912), .B(n5908), .S(n6103), .Z(n5098) );
  INV_X1 U6602 ( .A(SI_10_), .ZN(n5097) );
  NAND2_X1 U6603 ( .A1(n5098), .A2(n5097), .ZN(n5117) );
  INV_X1 U6604 ( .A(n5098), .ZN(n5099) );
  NAND2_X1 U6605 ( .A1(n5099), .A2(SI_10_), .ZN(n5100) );
  NAND2_X1 U6606 ( .A1(n5117), .A2(n5100), .ZN(n5114) );
  NAND2_X1 U6607 ( .A1(n5407), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U6608 ( .A1(n5082), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5101) );
  XNOR2_X1 U6609 ( .A(n5101), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U6610 ( .A1(n4307), .A2(n6000), .ZN(n5102) );
  OAI211_X1 U6611 ( .C1(n5104), .C2(n6791), .A(n5103), .B(n5102), .ZN(n7133)
         );
  NAND2_X1 U6612 ( .A1(n6932), .A2(n7133), .ZN(n7613) );
  INV_X1 U6613 ( .A(n7133), .ZN(n9427) );
  NAND2_X1 U6614 ( .A1(n9005), .A2(n9427), .ZN(n7630) );
  NAND2_X1 U6615 ( .A1(n7613), .A2(n7630), .ZN(n7736) );
  NAND2_X1 U6616 ( .A1(n7078), .A2(n7736), .ZN(n7077) );
  NAND2_X1 U6617 ( .A1(n6932), .A2(n9427), .ZN(n5105) );
  NAND2_X1 U6618 ( .A1(n7077), .A2(n5105), .ZN(n7090) );
  NAND2_X1 U6619 ( .A1(n7507), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5113) );
  INV_X1 U6620 ( .A(n5108), .ZN(n5106) );
  NAND2_X1 U6621 ( .A1(n5106), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5129) );
  INV_X1 U6622 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5107) );
  NAND2_X1 U6623 ( .A1(n5108), .A2(n5107), .ZN(n5109) );
  AND2_X1 U6624 ( .A1(n5129), .A2(n5109), .ZN(n7227) );
  NAND2_X1 U6625 ( .A1(n5460), .A2(n7227), .ZN(n5112) );
  NAND2_X1 U6626 ( .A1(n5535), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5111) );
  NAND2_X1 U6627 ( .A1(n5246), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5110) );
  NAND4_X1 U6628 ( .A1(n5113), .A2(n5112), .A3(n5111), .A4(n5110), .ZN(n9490)
         );
  INV_X1 U6629 ( .A(n5114), .ZN(n5115) );
  INV_X1 U6630 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5119) );
  MUX2_X1 U6631 ( .A(n5119), .B(n5931), .S(n6103), .Z(n5138) );
  XNOR2_X1 U6632 ( .A(n5138), .B(SI_11_), .ZN(n5135) );
  XNOR2_X1 U6633 ( .A(n5137), .B(n5135), .ZN(n6845) );
  NAND2_X1 U6634 ( .A1(n5278), .A2(n6845), .ZN(n5123) );
  OR2_X1 U6635 ( .A1(n5120), .A2(n4878), .ZN(n5121) );
  XNOR2_X1 U6636 ( .A(n5121), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6455) );
  NAND2_X1 U6637 ( .A1(n4307), .A2(n6455), .ZN(n5122) );
  NAND2_X1 U6638 ( .A1(n7090), .A2(n5124), .ZN(n5126) );
  INV_X1 U6639 ( .A(n9490), .ZN(n5520) );
  NAND2_X1 U6640 ( .A1(n5520), .A2(n9545), .ZN(n5125) );
  NAND2_X1 U6641 ( .A1(n5126), .A2(n5125), .ZN(n9496) );
  INV_X1 U6642 ( .A(n5129), .ZN(n5127) );
  NAND2_X1 U6643 ( .A1(n5127), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5164) );
  INV_X1 U6644 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5128) );
  NAND2_X1 U6645 ( .A1(n5129), .A2(n5128), .ZN(n5130) );
  AND2_X1 U6646 ( .A1(n5164), .A2(n5130), .ZN(n9493) );
  NAND2_X1 U6647 ( .A1(n5460), .A2(n9493), .ZN(n5134) );
  NAND2_X1 U6648 ( .A1(n7507), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5133) );
  NAND2_X1 U6649 ( .A1(n5535), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5132) );
  NAND2_X1 U6650 ( .A1(n5246), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5131) );
  INV_X1 U6651 ( .A(n5135), .ZN(n5136) );
  INV_X1 U6652 ( .A(n5138), .ZN(n5139) );
  NAND2_X1 U6653 ( .A1(n5139), .A2(SI_11_), .ZN(n5140) );
  MUX2_X1 U6654 ( .A(n5954), .B(n5943), .S(n6103), .Z(n5142) );
  INV_X1 U6655 ( .A(SI_12_), .ZN(n5141) );
  NAND2_X1 U6656 ( .A1(n5142), .A2(n5141), .ZN(n5152) );
  INV_X1 U6657 ( .A(n5142), .ZN(n5143) );
  NAND2_X1 U6658 ( .A1(n5143), .A2(SI_12_), .ZN(n5144) );
  NAND2_X1 U6659 ( .A1(n5152), .A2(n5144), .ZN(n5153) );
  XNOR2_X1 U6660 ( .A(n5154), .B(n5153), .ZN(n6940) );
  NAND2_X1 U6661 ( .A1(n6940), .A2(n7512), .ZN(n5150) );
  NAND2_X1 U6662 ( .A1(n5145), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5146) );
  MUX2_X1 U6663 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5146), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5148) );
  AND2_X1 U6664 ( .A1(n5148), .A2(n5147), .ZN(n9030) );
  AOI22_X1 U6665 ( .A1(n5407), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n4307), .B2(
        n9030), .ZN(n5149) );
  NAND2_X1 U6666 ( .A1(n5150), .A2(n5149), .ZN(n9495) );
  NAND2_X1 U6667 ( .A1(n5635), .A2(n9495), .ZN(n7614) );
  NAND2_X1 U6668 ( .A1(n9004), .A2(n9541), .ZN(n7635) );
  NAND2_X1 U6669 ( .A1(n9004), .A2(n9495), .ZN(n5151) );
  INV_X1 U6670 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n5155) );
  MUX2_X1 U6671 ( .A(n5155), .B(n8710), .S(n6103), .Z(n5157) );
  NAND2_X1 U6672 ( .A1(n5157), .A2(n5156), .ZN(n5173) );
  INV_X1 U6673 ( .A(n5157), .ZN(n5158) );
  NAND2_X1 U6674 ( .A1(n5158), .A2(SI_13_), .ZN(n5159) );
  XNOR2_X1 U6675 ( .A(n5172), .B(n4859), .ZN(n7058) );
  NAND2_X1 U6676 ( .A1(n7058), .A2(n7512), .ZN(n5162) );
  NAND2_X1 U6677 ( .A1(n5147), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5160) );
  XNOR2_X1 U6678 ( .A(n5160), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9634) );
  AOI22_X1 U6679 ( .A1(n5407), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n4307), .B2(
        n9634), .ZN(n5161) );
  NAND2_X1 U6680 ( .A1(n5164), .A2(n5163), .ZN(n5165) );
  AND2_X1 U6681 ( .A1(n5180), .A2(n5165), .ZN(n8939) );
  NAND2_X1 U6682 ( .A1(n5460), .A2(n8939), .ZN(n5169) );
  NAND2_X1 U6683 ( .A1(n7507), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U6684 ( .A1(n5535), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6685 ( .A1(n5246), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6686 ( .A1(n8938), .A2(n9491), .ZN(n5170) );
  NAND2_X1 U6687 ( .A1(n5171), .A2(n5170), .ZN(n7204) );
  NAND2_X1 U6688 ( .A1(n5172), .A2(n4859), .ZN(n5174) );
  MUX2_X1 U6689 ( .A(n5962), .B(n5958), .S(n6103), .Z(n5188) );
  XNOR2_X1 U6690 ( .A(n5188), .B(SI_14_), .ZN(n5187) );
  XNOR2_X1 U6691 ( .A(n5192), .B(n5187), .ZN(n7144) );
  NAND2_X1 U6692 ( .A1(n7144), .A2(n7512), .ZN(n5178) );
  OAI21_X1 U6693 ( .B1(n5147), .B2(P1_IR_REG_13__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5175) );
  NAND2_X1 U6694 ( .A1(n5175), .A2(n8726), .ZN(n5197) );
  OR2_X1 U6695 ( .A1(n5175), .A2(n8726), .ZN(n5176) );
  NAND2_X1 U6696 ( .A1(n5197), .A2(n5176), .ZN(n9043) );
  INV_X1 U6697 ( .A(n9043), .ZN(n9646) );
  AOI22_X1 U6698 ( .A1(n5407), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n4307), .B2(
        n9646), .ZN(n5177) );
  NAND2_X1 U6699 ( .A1(n7507), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5185) );
  INV_X1 U6700 ( .A(n5180), .ZN(n5179) );
  NAND2_X1 U6701 ( .A1(n5179), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5202) );
  INV_X1 U6702 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8847) );
  NAND2_X1 U6703 ( .A1(n5180), .A2(n8847), .ZN(n5181) );
  AND2_X1 U6704 ( .A1(n5202), .A2(n5181), .ZN(n8849) );
  NAND2_X1 U6705 ( .A1(n5460), .A2(n8849), .ZN(n5184) );
  NAND2_X1 U6706 ( .A1(n5535), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6707 ( .A1(n5246), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5182) );
  NAND4_X1 U6708 ( .A1(n5185), .A2(n5184), .A3(n5183), .A4(n5182), .ZN(n9275)
         );
  AND2_X1 U6709 ( .A1(n8848), .A2(n9275), .ZN(n5186) );
  INV_X1 U6710 ( .A(n5187), .ZN(n5191) );
  INV_X1 U6711 ( .A(n5188), .ZN(n5189) );
  NAND2_X1 U6712 ( .A1(n5189), .A2(SI_14_), .ZN(n5190) );
  MUX2_X1 U6713 ( .A(n6194), .B(n6188), .S(n6103), .Z(n5194) );
  NAND2_X1 U6714 ( .A1(n5194), .A2(n5193), .ZN(n5210) );
  INV_X1 U6715 ( .A(n5194), .ZN(n5195) );
  NAND2_X1 U6716 ( .A1(n5195), .A2(SI_15_), .ZN(n5196) );
  NAND2_X1 U6717 ( .A1(n5210), .A2(n5196), .ZN(n5211) );
  XNOR2_X1 U6718 ( .A(n5212), .B(n5211), .ZN(n7236) );
  NAND2_X1 U6719 ( .A1(n7236), .A2(n7512), .ZN(n5200) );
  NAND2_X1 U6720 ( .A1(n5197), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5198) );
  XNOR2_X1 U6721 ( .A(n5198), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9659) );
  AOI22_X1 U6722 ( .A1(n5407), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n4307), .B2(
        n9659), .ZN(n5199) );
  NAND2_X1 U6723 ( .A1(n7507), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5207) );
  INV_X1 U6724 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U6725 ( .A1(n5202), .A2(n5201), .ZN(n5203) );
  AND2_X1 U6726 ( .A1(n5224), .A2(n5203), .ZN(n9282) );
  NAND2_X1 U6727 ( .A1(n5460), .A2(n9282), .ZN(n5206) );
  NAND2_X1 U6728 ( .A1(n5535), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5205) );
  NAND2_X1 U6729 ( .A1(n5246), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5204) );
  NAND4_X1 U6730 ( .A1(n5207), .A2(n5206), .A3(n5205), .A4(n5204), .ZN(n9262)
         );
  NOR2_X1 U6731 ( .A1(n9286), .A2(n9262), .ZN(n5209) );
  NAND2_X1 U6732 ( .A1(n9286), .A2(n9262), .ZN(n5208) );
  MUX2_X1 U6733 ( .A(n6198), .B(n5213), .S(n6103), .Z(n5214) );
  NAND2_X1 U6734 ( .A1(n5214), .A2(n8628), .ZN(n5232) );
  INV_X1 U6735 ( .A(n5214), .ZN(n5215) );
  NAND2_X1 U6736 ( .A1(n5215), .A2(SI_16_), .ZN(n5216) );
  XNOR2_X1 U6737 ( .A(n5231), .B(n5230), .ZN(n7272) );
  NAND2_X1 U6738 ( .A1(n7272), .A2(n5278), .ZN(n5222) );
  NAND3_X1 U6739 ( .A1(n8726), .A2(n5218), .A3(n5217), .ZN(n5219) );
  NOR2_X2 U6740 ( .A1(n5147), .A2(n5219), .ZN(n5237) );
  OR2_X1 U6741 ( .A1(n5237), .A2(n4878), .ZN(n5220) );
  XNOR2_X1 U6742 ( .A(n5220), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9672) );
  AOI22_X1 U6743 ( .A1(n5407), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n4307), .B2(
        n9672), .ZN(n5221) );
  NAND2_X1 U6744 ( .A1(n7507), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5229) );
  NAND2_X1 U6745 ( .A1(n5223), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5244) );
  INV_X1 U6746 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8900) );
  NAND2_X1 U6747 ( .A1(n5224), .A2(n8900), .ZN(n5225) );
  AND2_X1 U6748 ( .A1(n5244), .A2(n5225), .ZN(n9265) );
  NAND2_X1 U6749 ( .A1(n5460), .A2(n9265), .ZN(n5228) );
  NAND2_X1 U6750 ( .A1(n5535), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6751 ( .A1(n5246), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5226) );
  OR2_X1 U6752 ( .A1(n8894), .A2(n5668), .ZN(n7652) );
  NAND2_X1 U6753 ( .A1(n8894), .A2(n5668), .ZN(n7651) );
  NAND2_X1 U6754 ( .A1(n7652), .A2(n7651), .ZN(n9256) );
  MUX2_X1 U6755 ( .A(n5235), .B(n5234), .S(n6103), .Z(n5252) );
  XNOR2_X1 U6756 ( .A(n5252), .B(SI_17_), .ZN(n5251) );
  XNOR2_X1 U6757 ( .A(n5256), .B(n5251), .ZN(n7283) );
  NAND2_X1 U6758 ( .A1(n7283), .A2(n7512), .ZN(n5242) );
  NAND2_X1 U6759 ( .A1(n5237), .A2(n5236), .ZN(n5279) );
  NAND2_X1 U6760 ( .A1(n5279), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6761 ( .A1(n5239), .A2(n5238), .ZN(n5257) );
  OR2_X1 U6762 ( .A1(n5239), .A2(n5238), .ZN(n5240) );
  AOI22_X1 U6763 ( .A1(n5407), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n4307), .B2(
        n9039), .ZN(n5241) );
  NAND2_X1 U6764 ( .A1(n7507), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5250) );
  INV_X1 U6765 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U6766 ( .A1(n5244), .A2(n5243), .ZN(n5245) );
  AND2_X1 U6767 ( .A1(n5263), .A2(n5245), .ZN(n9244) );
  NAND2_X1 U6768 ( .A1(n5460), .A2(n9244), .ZN(n5249) );
  NAND2_X1 U6769 ( .A1(n4960), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U6770 ( .A1(n5246), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5247) );
  NAND4_X1 U6771 ( .A1(n5250), .A2(n5249), .A3(n5248), .A4(n5247), .ZN(n9261)
         );
  INV_X1 U6772 ( .A(n5251), .ZN(n5255) );
  INV_X1 U6773 ( .A(n5252), .ZN(n5253) );
  NAND2_X1 U6774 ( .A1(n5253), .A2(SI_17_), .ZN(n5254) );
  MUX2_X1 U6775 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6103), .Z(n5273) );
  XNOR2_X1 U6776 ( .A(n5273), .B(SI_18_), .ZN(n5270) );
  XNOR2_X1 U6777 ( .A(n5272), .B(n5270), .ZN(n7362) );
  NAND2_X1 U6778 ( .A1(n7362), .A2(n7512), .ZN(n5260) );
  NAND2_X1 U6779 ( .A1(n5257), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5258) );
  XNOR2_X1 U6780 ( .A(n5258), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9038) );
  AOI22_X1 U6781 ( .A1(n5407), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n4307), .B2(
        n9038), .ZN(n5259) );
  NAND2_X1 U6782 ( .A1(n7507), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6783 ( .A1(n5261), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5288) );
  INV_X1 U6784 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U6785 ( .A1(n5263), .A2(n5262), .ZN(n5264) );
  AND2_X1 U6786 ( .A1(n5288), .A2(n5264), .ZN(n9236) );
  NAND2_X1 U6787 ( .A1(n5460), .A2(n9236), .ZN(n5267) );
  NAND2_X1 U6788 ( .A1(n5535), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5266) );
  NAND2_X1 U6789 ( .A1(n4884), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5265) );
  OR2_X1 U6790 ( .A1(n9356), .A2(n8911), .ZN(n7661) );
  NAND2_X1 U6791 ( .A1(n9356), .A2(n8911), .ZN(n7665) );
  OR2_X2 U6792 ( .A1(n9221), .A2(n9222), .ZN(n9223) );
  NAND2_X1 U6793 ( .A1(n9356), .A2(n9248), .ZN(n5269) );
  INV_X1 U6794 ( .A(n5270), .ZN(n5271) );
  MUX2_X1 U6795 ( .A(n6587), .B(n6589), .S(n6103), .Z(n5275) );
  INV_X1 U6796 ( .A(SI_19_), .ZN(n5274) );
  NAND2_X1 U6797 ( .A1(n5275), .A2(n5274), .ZN(n5295) );
  INV_X1 U6798 ( .A(n5275), .ZN(n5276) );
  NAND2_X1 U6799 ( .A1(n5276), .A2(SI_19_), .ZN(n5277) );
  NAND2_X1 U6800 ( .A1(n5295), .A2(n5277), .ZN(n5296) );
  XNOR2_X1 U6801 ( .A(n5297), .B(n5296), .ZN(n7368) );
  NAND2_X1 U6802 ( .A1(n7368), .A2(n5278), .ZN(n5286) );
  INV_X1 U6803 ( .A(n5283), .ZN(n5280) );
  NAND2_X1 U6804 ( .A1(n5280), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5281) );
  MUX2_X1 U6805 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5281), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n5284) );
  NAND2_X1 U6806 ( .A1(n5283), .A2(n5282), .ZN(n5465) );
  AOI22_X1 U6807 ( .A1(n5407), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9745), .B2(
        n4307), .ZN(n5285) );
  NAND2_X1 U6808 ( .A1(n7507), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5293) );
  INV_X1 U6809 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5287) );
  NAND2_X1 U6810 ( .A1(n5288), .A2(n5287), .ZN(n5289) );
  AND2_X1 U6811 ( .A1(n5306), .A2(n5289), .ZN(n9210) );
  NAND2_X1 U6812 ( .A1(n5460), .A2(n9210), .ZN(n5292) );
  NAND2_X1 U6813 ( .A1(n4960), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6814 ( .A1(n4884), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5290) );
  NAND4_X1 U6815 ( .A1(n5293), .A2(n5292), .A3(n5291), .A4(n5290), .ZN(n9230)
         );
  OR2_X1 U6816 ( .A1(n9350), .A2(n9230), .ZN(n5294) );
  MUX2_X1 U6817 ( .A(n7387), .B(n6725), .S(n6103), .Z(n5299) );
  NAND2_X1 U6818 ( .A1(n5299), .A2(n5298), .ZN(n5314) );
  INV_X1 U6819 ( .A(n5299), .ZN(n5300) );
  NAND2_X1 U6820 ( .A1(n5300), .A2(SI_20_), .ZN(n5301) );
  XNOR2_X1 U6821 ( .A(n5313), .B(n5312), .ZN(n7386) );
  NAND2_X1 U6822 ( .A1(n7386), .A2(n7512), .ZN(n5303) );
  NAND2_X1 U6823 ( .A1(n5407), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5302) );
  NAND2_X1 U6824 ( .A1(n7507), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U6825 ( .A1(n5304), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5319) );
  INV_X1 U6826 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U6827 ( .A1(n5306), .A2(n5305), .ZN(n5307) );
  AND2_X1 U6828 ( .A1(n5319), .A2(n5307), .ZN(n9196) );
  NAND2_X1 U6829 ( .A1(n5460), .A2(n9196), .ZN(n5310) );
  NAND2_X1 U6830 ( .A1(n4960), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U6831 ( .A1(n4884), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5308) );
  NAND4_X1 U6832 ( .A1(n5311), .A2(n5310), .A3(n5309), .A4(n5308), .ZN(n9216)
         );
  INV_X1 U6833 ( .A(n9174), .ZN(n5326) );
  NAND2_X1 U6834 ( .A1(n5313), .A2(n5312), .ZN(n5315) );
  MUX2_X1 U6835 ( .A(n7401), .B(n6789), .S(n6103), .Z(n5329) );
  XNOR2_X1 U6836 ( .A(n5329), .B(SI_21_), .ZN(n5328) );
  XNOR2_X1 U6837 ( .A(n5327), .B(n5328), .ZN(n7400) );
  NAND2_X1 U6838 ( .A1(n7400), .A2(n7512), .ZN(n5317) );
  NAND2_X1 U6839 ( .A1(n5407), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6840 ( .A1(n7507), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5324) );
  INV_X1 U6841 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5318) );
  NAND2_X1 U6842 ( .A1(n5319), .A2(n5318), .ZN(n5320) );
  AND2_X1 U6843 ( .A1(n5338), .A2(n5320), .ZN(n9188) );
  NAND2_X1 U6844 ( .A1(n5460), .A2(n9188), .ZN(n5323) );
  NAND2_X1 U6845 ( .A1(n5535), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6846 ( .A1(n4884), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5321) );
  OR2_X1 U6847 ( .A1(n9185), .A2(n8955), .ZN(n7672) );
  NAND2_X1 U6848 ( .A1(n9185), .A2(n8955), .ZN(n7673) );
  NAND2_X1 U6849 ( .A1(n5326), .A2(n5325), .ZN(n9172) );
  NAND2_X1 U6850 ( .A1(n9172), .A2(n4854), .ZN(n9160) );
  INV_X1 U6851 ( .A(n5329), .ZN(n5330) );
  NAND2_X1 U6852 ( .A1(n5330), .A2(SI_21_), .ZN(n5331) );
  MUX2_X1 U6853 ( .A(n7418), .B(n6929), .S(n6103), .Z(n5333) );
  INV_X1 U6854 ( .A(SI_22_), .ZN(n5332) );
  NAND2_X1 U6855 ( .A1(n5333), .A2(n5332), .ZN(n5346) );
  INV_X1 U6856 ( .A(n5333), .ZN(n5334) );
  NAND2_X1 U6857 ( .A1(n5334), .A2(SI_22_), .ZN(n5335) );
  NAND2_X1 U6858 ( .A1(n5346), .A2(n5335), .ZN(n5347) );
  XNOR2_X1 U6859 ( .A(n5348), .B(n5347), .ZN(n7417) );
  NAND2_X1 U6860 ( .A1(n7417), .A2(n7512), .ZN(n5337) );
  NAND2_X1 U6861 ( .A1(n5407), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U6862 ( .A1(n7507), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5343) );
  INV_X1 U6863 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8954) );
  NAND2_X1 U6864 ( .A1(n5338), .A2(n8954), .ZN(n5339) );
  AND2_X1 U6865 ( .A1(n5361), .A2(n5339), .ZN(n9162) );
  NAND2_X1 U6866 ( .A1(n5460), .A2(n9162), .ZN(n5342) );
  NAND2_X1 U6867 ( .A1(n5535), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U6868 ( .A1(n4884), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5340) );
  NAND4_X1 U6869 ( .A1(n5343), .A2(n5342), .A3(n5341), .A4(n5340), .ZN(n9182)
         );
  NAND2_X1 U6870 ( .A1(n9160), .A2(n5344), .ZN(n5345) );
  NAND2_X1 U6871 ( .A1(n5345), .A2(n4857), .ZN(n9141) );
  INV_X1 U6872 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5349) );
  MUX2_X1 U6873 ( .A(n8702), .B(n5349), .S(n6103), .Z(n5351) );
  INV_X1 U6874 ( .A(SI_23_), .ZN(n5350) );
  NAND2_X1 U6875 ( .A1(n5351), .A2(n5350), .ZN(n5369) );
  INV_X1 U6876 ( .A(n5351), .ZN(n5352) );
  NAND2_X1 U6877 ( .A1(n5352), .A2(SI_23_), .ZN(n5353) );
  OR2_X1 U6878 ( .A1(n5355), .A2(n5354), .ZN(n5356) );
  NAND2_X1 U6879 ( .A1(n5370), .A2(n5356), .ZN(n7430) );
  NAND2_X1 U6880 ( .A1(n7430), .A2(n7512), .ZN(n5358) );
  NAND2_X1 U6881 ( .A1(n5407), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5357) );
  NAND2_X1 U6882 ( .A1(n7507), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5366) );
  INV_X1 U6883 ( .A(n5361), .ZN(n5359) );
  NAND2_X1 U6884 ( .A1(n5359), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5375) );
  INV_X1 U6885 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U6886 ( .A1(n5361), .A2(n5360), .ZN(n5362) );
  AND2_X1 U6887 ( .A1(n5375), .A2(n5362), .ZN(n9145) );
  NAND2_X1 U6888 ( .A1(n5460), .A2(n9145), .ZN(n5365) );
  NAND2_X1 U6889 ( .A1(n5535), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U6890 ( .A1(n4884), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5363) );
  NAND4_X1 U6891 ( .A1(n5366), .A2(n5365), .A3(n5364), .A4(n5363), .ZN(n9167)
         );
  NAND2_X1 U6892 ( .A1(n9147), .A2(n8952), .ZN(n5367) );
  NAND2_X1 U6893 ( .A1(n9141), .A2(n5367), .ZN(n5368) );
  NAND2_X1 U6894 ( .A1(n5368), .A2(n4853), .ZN(n9127) );
  INV_X1 U6895 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7354) );
  INV_X1 U6896 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7125) );
  MUX2_X1 U6897 ( .A(n7354), .B(n7125), .S(n6103), .Z(n5384) );
  XNOR2_X1 U6898 ( .A(n5384), .B(SI_24_), .ZN(n5381) );
  NAND2_X1 U6899 ( .A1(n7353), .A2(n7512), .ZN(n5372) );
  NAND2_X1 U6900 ( .A1(n5407), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5371) );
  INV_X1 U6901 ( .A(n5375), .ZN(n5373) );
  NAND2_X1 U6902 ( .A1(n5373), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5393) );
  INV_X1 U6903 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6904 ( .A1(n5375), .A2(n5374), .ZN(n5376) );
  AND2_X1 U6905 ( .A1(n5393), .A2(n5376), .ZN(n9135) );
  NAND2_X1 U6906 ( .A1(n9135), .A2(n5460), .ZN(n5380) );
  NAND2_X1 U6907 ( .A1(n7507), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6908 ( .A1(n4960), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U6909 ( .A1(n4884), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5377) );
  NAND4_X1 U6910 ( .A1(n5380), .A2(n5379), .A3(n5378), .A4(n5377), .ZN(n9154)
         );
  AND2_X1 U6911 ( .A1(n9323), .A2(n9154), .ZN(n7718) );
  OR2_X1 U6912 ( .A1(n9323), .A2(n9154), .ZN(n7719) );
  OAI21_X2 U6913 ( .B1(n9127), .B2(n7718), .A(n7719), .ZN(n9115) );
  INV_X1 U6914 ( .A(n5381), .ZN(n5382) );
  INV_X1 U6915 ( .A(n5384), .ZN(n5385) );
  NAND2_X1 U6916 ( .A1(n5385), .A2(SI_24_), .ZN(n5386) );
  INV_X1 U6917 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8841) );
  INV_X1 U6918 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n9400) );
  MUX2_X1 U6919 ( .A(n8841), .B(n9400), .S(n6103), .Z(n5387) );
  NAND2_X1 U6920 ( .A1(n5387), .A2(n8779), .ZN(n5400) );
  INV_X1 U6921 ( .A(n5387), .ZN(n5388) );
  NAND2_X1 U6922 ( .A1(n5388), .A2(SI_25_), .ZN(n5389) );
  NAND2_X1 U6923 ( .A1(n5400), .A2(n5389), .ZN(n5401) );
  XNOR2_X1 U6924 ( .A(n5402), .B(n5401), .ZN(n8837) );
  NAND2_X1 U6925 ( .A1(n8837), .A2(n7512), .ZN(n5391) );
  NAND2_X1 U6926 ( .A1(n4992), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5390) );
  INV_X1 U6927 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U6928 ( .A1(n5393), .A2(n5392), .ZN(n5394) );
  AND2_X1 U6929 ( .A1(n5412), .A2(n5394), .ZN(n9117) );
  NAND2_X1 U6930 ( .A1(n9117), .A2(n5460), .ZN(n5399) );
  NAND2_X1 U6931 ( .A1(n7507), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5396) );
  NAND2_X1 U6932 ( .A1(n4960), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5395) );
  AND2_X1 U6933 ( .A1(n5396), .A2(n5395), .ZN(n5398) );
  NAND2_X1 U6934 ( .A1(n4884), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6935 ( .A1(n9317), .A2(n5733), .ZN(n7694) );
  NAND2_X1 U6936 ( .A1(n9105), .A2(n7694), .ZN(n9121) );
  INV_X1 U6937 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8834) );
  MUX2_X1 U6938 ( .A(n8834), .B(n9394), .S(n6103), .Z(n5404) );
  INV_X1 U6939 ( .A(SI_26_), .ZN(n5403) );
  NAND2_X1 U6940 ( .A1(n5404), .A2(n5403), .ZN(n5421) );
  INV_X1 U6941 ( .A(n5404), .ZN(n5405) );
  NAND2_X1 U6942 ( .A1(n5405), .A2(SI_26_), .ZN(n5406) );
  XNOR2_X1 U6943 ( .A(n5420), .B(n5419), .ZN(n8833) );
  NAND2_X1 U6944 ( .A1(n8833), .A2(n7512), .ZN(n5409) );
  NAND2_X1 U6945 ( .A1(n5407), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5408) );
  INV_X1 U6946 ( .A(n5412), .ZN(n5410) );
  NAND2_X1 U6947 ( .A1(n5410), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5441) );
  INV_X1 U6948 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U6949 ( .A1(n5412), .A2(n5411), .ZN(n5413) );
  NAND2_X1 U6950 ( .A1(n5441), .A2(n5413), .ZN(n5762) );
  OR2_X1 U6951 ( .A1(n5762), .A2(n5414), .ZN(n5417) );
  AOI22_X1 U6952 ( .A1(n4960), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n4884), .B2(
        P1_REG0_REG_26__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U6953 ( .A1(n7507), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U6954 ( .A1(n9104), .A2(n5796), .ZN(n5418) );
  NAND2_X1 U6955 ( .A1(n5420), .A2(n5419), .ZN(n5422) );
  INV_X1 U6956 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8832) );
  INV_X1 U6957 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5423) );
  MUX2_X1 U6958 ( .A(n8832), .B(n5423), .S(n6103), .Z(n5425) );
  INV_X1 U6959 ( .A(SI_27_), .ZN(n5424) );
  NAND2_X1 U6960 ( .A1(n5425), .A2(n5424), .ZN(n5435) );
  INV_X1 U6961 ( .A(n5425), .ZN(n5426) );
  NAND2_X1 U6962 ( .A1(n5426), .A2(SI_27_), .ZN(n5427) );
  NAND2_X1 U6963 ( .A1(n8831), .A2(n7512), .ZN(n5429) );
  NAND2_X1 U6964 ( .A1(n5407), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5428) );
  NAND2_X2 U6965 ( .A1(n5429), .A2(n5428), .ZN(n9307) );
  XNOR2_X1 U6966 ( .A(n5441), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9087) );
  INV_X1 U6967 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U6968 ( .A1(n7507), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6969 ( .A1(n4960), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5430) );
  OAI211_X1 U6970 ( .C1(n5006), .C2(n8723), .A(n5431), .B(n5430), .ZN(n5432)
         );
  NAND2_X1 U6971 ( .A1(n9307), .A2(n9003), .ZN(n7554) );
  INV_X1 U6972 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8040) );
  MUX2_X1 U6973 ( .A(n8040), .B(n8698), .S(n6103), .Z(n5453) );
  XNOR2_X1 U6974 ( .A(n5453), .B(SI_28_), .ZN(n5450) );
  NAND2_X1 U6975 ( .A1(n8039), .A2(n7512), .ZN(n5438) );
  NAND2_X1 U6976 ( .A1(n5407), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5437) );
  INV_X1 U6977 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5795) );
  INV_X1 U6978 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5439) );
  OAI21_X1 U6979 ( .B1(n5441), .B2(n5795), .A(n5439), .ZN(n5442) );
  NAND2_X1 U6980 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5440) );
  OR2_X1 U6981 ( .A1(n5441), .A2(n5440), .ZN(n5459) );
  NAND2_X1 U6982 ( .A1(n9075), .A2(n5460), .ZN(n5449) );
  INV_X1 U6983 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U6984 ( .A1(n7507), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U6985 ( .A1(n4884), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5443) );
  OAI211_X1 U6986 ( .C1(n5446), .C2(n5445), .A(n5444), .B(n5443), .ZN(n5447)
         );
  INV_X1 U6987 ( .A(n5447), .ZN(n5448) );
  NAND2_X1 U6988 ( .A1(n9302), .A2(n9090), .ZN(n7706) );
  NAND2_X1 U6989 ( .A1(n7705), .A2(n7706), .ZN(n9071) );
  NAND2_X1 U6990 ( .A1(n9070), .A2(n4357), .ZN(n5464) );
  INV_X1 U6991 ( .A(SI_28_), .ZN(n5452) );
  NAND2_X1 U6992 ( .A1(n5453), .A2(n5452), .ZN(n5454) );
  INV_X1 U6993 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8830) );
  INV_X1 U6994 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9384) );
  MUX2_X1 U6995 ( .A(n8830), .B(n9384), .S(n6103), .Z(n7328) );
  XNOR2_X1 U6996 ( .A(n7328), .B(SI_29_), .ZN(n5456) );
  NAND2_X1 U6997 ( .A1(n8828), .A2(n7512), .ZN(n5458) );
  NAND2_X1 U6998 ( .A1(n4992), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5457) );
  INV_X1 U6999 ( .A(n5459), .ZN(n5543) );
  NAND2_X1 U7000 ( .A1(n5543), .A2(n5460), .ZN(n5463) );
  AOI22_X1 U7001 ( .A1(n4960), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n4884), .B2(
        P1_REG0_REG_29__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U7002 ( .A1(n7507), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5461) );
  OR2_X1 U7003 ( .A1(n9297), .A2(n8050), .ZN(n7580) );
  NAND2_X1 U7004 ( .A1(n9297), .A2(n8050), .ZN(n7771) );
  NAND2_X1 U7005 ( .A1(n7580), .A2(n7771), .ZN(n7750) );
  NAND2_X2 U7006 ( .A1(n5465), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U7007 ( .A1(n5472), .A2(n5473), .ZN(n5466) );
  XNOR2_X2 U7008 ( .A(n5467), .B(P1_IR_REG_22__SCAN_IN), .ZN(n5509) );
  XNOR2_X2 U7009 ( .A(n5472), .B(n5473), .ZN(n6726) );
  NAND2_X1 U7010 ( .A1(n5474), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U7011 ( .A1(n5477), .A2(n5476), .ZN(n5479) );
  OR2_X1 U7012 ( .A1(n5477), .A2(n5476), .ZN(n5478) );
  NAND2_X1 U7013 ( .A1(n5479), .A2(n5478), .ZN(n9398) );
  INV_X1 U7014 ( .A(n5480), .ZN(n5481) );
  NAND2_X1 U7015 ( .A1(n5481), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5483) );
  NAND3_X1 U7016 ( .A1(n9398), .A2(P1_B_REG_SCAN_IN), .A3(n7126), .ZN(n5486)
         );
  INV_X1 U7017 ( .A(n7126), .ZN(n5484) );
  INV_X1 U7018 ( .A(P1_B_REG_SCAN_IN), .ZN(n5533) );
  NAND2_X1 U7019 ( .A1(n5484), .A2(n5533), .ZN(n5485) );
  INV_X1 U7020 ( .A(n5504), .ZN(n9395) );
  NAND2_X1 U7021 ( .A1(n9395), .A2(n7126), .ZN(n9380) );
  OAI21_X1 U7022 ( .B1(n9378), .B2(P1_D_REG_0__SCAN_IN), .A(n9380), .ZN(n5500)
         );
  NOR4_X1 U7023 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5491) );
  NOR4_X1 U7024 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5490) );
  NOR4_X1 U7025 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5489) );
  NOR4_X1 U7026 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5488) );
  AND4_X1 U7027 ( .A1(n5491), .A2(n5490), .A3(n5489), .A4(n5488), .ZN(n5497)
         );
  NOR2_X1 U7028 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .ZN(
        n5495) );
  NOR4_X1 U7029 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5494) );
  NOR4_X1 U7030 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5493) );
  NOR4_X1 U7031 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5492) );
  AND4_X1 U7032 ( .A1(n5495), .A2(n5494), .A3(n5493), .A4(n5492), .ZN(n5496)
         );
  NAND2_X1 U7033 ( .A1(n5497), .A2(n5496), .ZN(n5755) );
  INV_X1 U7034 ( .A(n5755), .ZN(n5498) );
  OR2_X1 U7035 ( .A1(n9378), .A2(n5498), .ZN(n5499) );
  OR2_X1 U7036 ( .A1(n9378), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5503) );
  INV_X1 U7037 ( .A(n9398), .ZN(n5501) );
  OR2_X1 U7038 ( .A1(n5504), .A2(n5501), .ZN(n5502) );
  NAND2_X1 U7039 ( .A1(n5503), .A2(n5502), .ZN(n6085) );
  NOR2_X1 U7040 ( .A1(n9398), .A2(n7126), .ZN(n5505) );
  NAND2_X1 U7041 ( .A1(n4401), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5507) );
  AND2_X1 U7042 ( .A1(n6985), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5508) );
  NOR2_X1 U7043 ( .A1(n6085), .A2(n9791), .ZN(n9790) );
  NAND3_X1 U7044 ( .A1(n6088), .A2(n6091), .A3(n9790), .ZN(n5542) );
  OR2_X1 U7045 ( .A1(n6572), .A2(n5550), .ZN(n6092) );
  NAND2_X4 U7046 ( .A1(n6572), .A2(n5550), .ZN(n8043) );
  XNOR2_X2 U7047 ( .A(n5562), .B(n7524), .ZN(n7726) );
  INV_X1 U7048 ( .A(n6565), .ZN(n6582) );
  NAND2_X1 U7049 ( .A1(n7525), .A2(n7524), .ZN(n5511) );
  NAND2_X1 U7050 ( .A1(n7530), .A2(n7723), .ZN(n5512) );
  NAND2_X1 U7051 ( .A1(n5512), .A2(n7526), .ZN(n6683) );
  INV_X1 U7052 ( .A(n5513), .ZN(n6684) );
  NAND2_X1 U7053 ( .A1(n6683), .A2(n6684), .ZN(n5514) );
  NAND2_X1 U7054 ( .A1(n5514), .A2(n7727), .ZN(n7587) );
  AND3_X1 U7055 ( .A1(n7588), .A2(n9766), .A3(n7729), .ZN(n7728) );
  NAND2_X1 U7056 ( .A1(n9769), .A2(n7728), .ZN(n5517) );
  INV_X1 U7057 ( .A(n7590), .ZN(n7600) );
  NAND2_X1 U7058 ( .A1(n7729), .A2(n7600), .ZN(n5516) );
  AND2_X1 U7059 ( .A1(n5516), .A2(n7757), .ZN(n7535) );
  NAND2_X1 U7060 ( .A1(n5517), .A2(n7535), .ZN(n6917) );
  INV_X1 U7061 ( .A(n6917), .ZN(n5519) );
  INV_X1 U7062 ( .A(n7602), .ZN(n9724) );
  NAND2_X1 U7063 ( .A1(n9006), .A2(n9850), .ZN(n7626) );
  NAND2_X1 U7064 ( .A1(n7630), .A2(n7626), .ZN(n7611) );
  NAND2_X1 U7065 ( .A1(n9721), .A2(n7046), .ZN(n7609) );
  NAND2_X1 U7066 ( .A1(n7609), .A2(n7613), .ZN(n7629) );
  NAND2_X1 U7067 ( .A1(n7629), .A2(n7630), .ZN(n7091) );
  NAND2_X1 U7068 ( .A1(n5520), .A2(n7226), .ZN(n9486) );
  AND2_X1 U7069 ( .A1(n7614), .A2(n9486), .ZN(n7637) );
  AND2_X1 U7070 ( .A1(n7091), .A2(n7637), .ZN(n7540) );
  NAND2_X1 U7071 ( .A1(n7092), .A2(n7540), .ZN(n5522) );
  NAND3_X1 U7072 ( .A1(n7614), .A2(n9545), .A3(n9490), .ZN(n5521) );
  AND2_X1 U7073 ( .A1(n5521), .A2(n7635), .ZN(n7616) );
  NAND2_X1 U7074 ( .A1(n9532), .A2(n9491), .ZN(n7518) );
  NAND2_X1 U7075 ( .A1(n7264), .A2(n8938), .ZN(n7538) );
  NAND2_X1 U7076 ( .A1(n7518), .A2(n7538), .ZN(n7192) );
  INV_X1 U7077 ( .A(n9275), .ZN(n8995) );
  OR2_X1 U7078 ( .A1(n8848), .A2(n8995), .ZN(n7620) );
  NAND2_X1 U7079 ( .A1(n8848), .A2(n8995), .ZN(n7586) );
  NAND2_X1 U7080 ( .A1(n7620), .A2(n7586), .ZN(n7740) );
  INV_X1 U7081 ( .A(n7538), .ZN(n7516) );
  NOR2_X1 U7082 ( .A1(n7740), .A2(n7516), .ZN(n5523) );
  INV_X1 U7083 ( .A(n9262), .ZN(n8902) );
  NAND2_X1 U7084 ( .A1(n9286), .A2(n8902), .ZN(n7647) );
  NAND2_X1 U7085 ( .A1(n9273), .A2(n7647), .ZN(n5524) );
  OR2_X1 U7086 ( .A1(n9286), .A2(n8902), .ZN(n7646) );
  NAND2_X1 U7087 ( .A1(n5524), .A2(n7646), .ZN(n9257) );
  INV_X1 U7088 ( .A(n9261), .ZN(n8981) );
  NAND2_X1 U7089 ( .A1(n9359), .A2(n8981), .ZN(n7650) );
  OR2_X1 U7090 ( .A1(n9359), .A2(n8981), .ZN(n9225) );
  AND2_X1 U7091 ( .A1(n7661), .A2(n9225), .ZN(n7657) );
  INV_X1 U7092 ( .A(n9230), .ZN(n8930) );
  OR2_X1 U7093 ( .A1(n9350), .A2(n8930), .ZN(n7660) );
  NAND2_X1 U7094 ( .A1(n9350), .A2(n8930), .ZN(n7664) );
  NAND2_X1 U7095 ( .A1(n9214), .A2(n9215), .ZN(n9213) );
  INV_X1 U7096 ( .A(n9216), .ZN(n5526) );
  AND2_X1 U7097 ( .A1(n9344), .A2(n5526), .ZN(n7721) );
  INV_X1 U7098 ( .A(n9344), .ZN(n9198) );
  AND2_X1 U7099 ( .A1(n9198), .A2(n9216), .ZN(n7722) );
  NOR2_X1 U7100 ( .A1(n5325), .A2(n7722), .ZN(n5527) );
  OR2_X1 U7101 ( .A1(n9332), .A2(n8882), .ZN(n7676) );
  NAND2_X1 U7102 ( .A1(n9332), .A2(n8882), .ZN(n7675) );
  NAND2_X1 U7103 ( .A1(n9147), .A2(n9167), .ZN(n7686) );
  NAND2_X1 U7104 ( .A1(n9327), .A2(n8952), .ZN(n7545) );
  NAND2_X1 U7105 ( .A1(n9152), .A2(n7686), .ZN(n9130) );
  INV_X1 U7106 ( .A(n9154), .ZN(n8890) );
  NAND2_X1 U7107 ( .A1(n9323), .A2(n8890), .ZN(n7683) );
  AND2_X1 U7108 ( .A1(n9128), .A2(n9154), .ZN(n7684) );
  INV_X1 U7109 ( .A(n7694), .ZN(n5528) );
  OR2_X1 U7110 ( .A1(n9313), .A2(n5796), .ZN(n7698) );
  NAND2_X1 U7111 ( .A1(n7698), .A2(n9105), .ZN(n7566) );
  NAND2_X1 U7112 ( .A1(n9313), .A2(n5796), .ZN(n7699) );
  INV_X1 U7113 ( .A(n9071), .ZN(n9079) );
  NAND2_X1 U7114 ( .A1(n9078), .A2(n9079), .ZN(n9077) );
  NAND2_X1 U7115 ( .A1(n5509), .A2(n9745), .ZN(n5531) );
  OR2_X1 U7116 ( .A1(n7776), .A2(n6726), .ZN(n7786) );
  INV_X1 U7117 ( .A(n7756), .ZN(n5753) );
  INV_X1 U7118 ( .A(n5532), .ZN(n6229) );
  NOR2_X1 U7119 ( .A1(n7492), .A2(n5533), .ZN(n5534) );
  NOR2_X1 U7120 ( .A1(n9772), .A2(n5534), .ZN(n9060) );
  INV_X1 U7121 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U7122 ( .A1(n7507), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U7123 ( .A1(n4884), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5536) );
  OAI211_X1 U7124 ( .C1(n5446), .C2(n5538), .A(n5537), .B(n5536), .ZN(n9001)
         );
  NOR2_X1 U7125 ( .A1(n9300), .A2(n9755), .ZN(n5548) );
  NAND2_X1 U7126 ( .A1(n6688), .A2(n9805), .ZN(n9759) );
  NAND2_X1 U7127 ( .A1(n7098), .A2(n9545), .ZN(n9501) );
  INV_X1 U7128 ( .A(n8848), .ZN(n9527) );
  INV_X1 U7129 ( .A(n9356), .ZN(n9239) );
  INV_X1 U7130 ( .A(n9350), .ZN(n9212) );
  AOI21_X1 U7131 ( .B1(n9297), .B2(n9073), .A(n9065), .ZN(n9298) );
  OR2_X1 U7132 ( .A1(n5542), .A2(n9745), .ZN(n9500) );
  INV_X1 U7133 ( .A(n9500), .ZN(n9235) );
  AND2_X1 U7134 ( .A1(n6093), .A2(n7783), .ZN(n9740) );
  AOI22_X1 U7135 ( .A1(P1_REG2_REG_29__SCAN_IN), .A2(n9755), .B1(n5543), .B2(
        n9783), .ZN(n5544) );
  OAI21_X1 U7136 ( .B1(n4512), .B2(n9765), .A(n5544), .ZN(n5545) );
  OAI21_X1 U7137 ( .B1(n9301), .B2(n9290), .A(n5549), .ZN(P1_U3355) );
  INV_X2 U7138 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NAND2_X1 U7139 ( .A1(n7788), .A2(n5751), .ZN(n6573) );
  AND2_X4 U7140 ( .A1(n6573), .A2(n4310), .ZN(n8045) );
  OAI22_X1 U7141 ( .A1(n9147), .A2(n5739), .B1(n8952), .B2(n5785), .ZN(n8860)
         );
  NAND2_X1 U7142 ( .A1(n5553), .A2(n8045), .ZN(n5552) );
  AOI22_X1 U7143 ( .A1(n6565), .A2(n4313), .B1(n5554), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U7144 ( .A1(n5988), .A2(n5987), .ZN(n5559) );
  INV_X1 U7145 ( .A(n5987), .ZN(n5557) );
  NAND2_X1 U7146 ( .A1(n5557), .A2(n5783), .ZN(n5558) );
  NAND2_X1 U7147 ( .A1(n5559), .A2(n5558), .ZN(n5564) );
  INV_X2 U7148 ( .A(n4309), .ZN(n5737) );
  OAI22_X1 U7149 ( .A1(n7525), .A2(n4312), .B1(n9795), .B2(n5737), .ZN(n5561)
         );
  XNOR2_X1 U7150 ( .A(n5561), .B(n8043), .ZN(n5565) );
  NAND2_X1 U7151 ( .A1(n5564), .A2(n5565), .ZN(n6021) );
  NOR2_X1 U7152 ( .A1(n9795), .A2(n4312), .ZN(n5563) );
  AOI21_X1 U7153 ( .B1(n5562), .B2(n8045), .A(n5563), .ZN(n6022) );
  NAND2_X1 U7154 ( .A1(n6021), .A2(n6022), .ZN(n6020) );
  INV_X1 U7155 ( .A(n5564), .ZN(n5567) );
  INV_X1 U7156 ( .A(n5565), .ZN(n5566) );
  NAND2_X1 U7157 ( .A1(n5567), .A2(n5566), .ZN(n6024) );
  NAND2_X1 U7158 ( .A1(n6020), .A2(n6024), .ZN(n8960) );
  OAI22_X1 U7159 ( .A1(n4934), .A2(n4312), .B1(n4931), .B2(n5737), .ZN(n5568)
         );
  OAI22_X1 U7160 ( .A1(n4934), .A2(n5785), .B1(n4931), .B2(n4312), .ZN(n5570)
         );
  XNOR2_X1 U7161 ( .A(n5569), .B(n5570), .ZN(n8962) );
  NAND2_X1 U7162 ( .A1(n8960), .A2(n8962), .ZN(n8961) );
  INV_X1 U7163 ( .A(n5569), .ZN(n5571) );
  OR2_X1 U7164 ( .A1(n5571), .A2(n5570), .ZN(n5572) );
  NAND2_X1 U7165 ( .A1(n8961), .A2(n5572), .ZN(n6248) );
  OAI22_X1 U7166 ( .A1(n4956), .A2(n5739), .B1(n9805), .B2(n5737), .ZN(n5573)
         );
  XNOR2_X1 U7167 ( .A(n5573), .B(n5783), .ZN(n5577) );
  OR2_X1 U7168 ( .A1(n4956), .A2(n5785), .ZN(n5575) );
  NAND2_X1 U7169 ( .A1(n6692), .A2(n5625), .ZN(n5574) );
  NAND2_X1 U7170 ( .A1(n5575), .A2(n5574), .ZN(n5578) );
  INV_X1 U7171 ( .A(n5578), .ZN(n5576) );
  AND2_X1 U7172 ( .A1(n5577), .A2(n5576), .ZN(n6245) );
  INV_X1 U7173 ( .A(n5577), .ZN(n5579) );
  NAND2_X1 U7174 ( .A1(n5579), .A2(n5578), .ZN(n6244) );
  OAI21_X1 U7175 ( .B1(n6248), .B2(n6245), .A(n6244), .ZN(n6487) );
  OAI22_X1 U7176 ( .A1(n9748), .A2(n5739), .B1(n9813), .B2(n5737), .ZN(n5580)
         );
  XNOR2_X1 U7177 ( .A(n5580), .B(n5783), .ZN(n5581) );
  OAI22_X1 U7178 ( .A1(n9748), .A2(n5785), .B1(n9813), .B2(n5739), .ZN(n5582)
         );
  XNOR2_X1 U7179 ( .A(n5581), .B(n5582), .ZN(n6486) );
  NAND2_X1 U7180 ( .A1(n6487), .A2(n6486), .ZN(n6485) );
  INV_X1 U7181 ( .A(n5581), .ZN(n5583) );
  NAND2_X1 U7182 ( .A1(n5583), .A2(n5582), .ZN(n5584) );
  NAND2_X1 U7183 ( .A1(n6485), .A2(n5584), .ZN(n6767) );
  OAI22_X1 U7184 ( .A1(n6919), .A2(n5739), .B1(n6909), .B2(n5737), .ZN(n5585)
         );
  XNOR2_X1 U7185 ( .A(n5585), .B(n8043), .ZN(n6904) );
  OR2_X1 U7186 ( .A1(n6919), .A2(n5785), .ZN(n5587) );
  NAND2_X1 U7187 ( .A1(n9826), .A2(n4308), .ZN(n5586) );
  NAND2_X1 U7188 ( .A1(n5587), .A2(n5586), .ZN(n6903) );
  NAND2_X1 U7189 ( .A1(n6904), .A2(n6903), .ZN(n5595) );
  OAI22_X1 U7190 ( .A1(n9773), .A2(n5739), .B1(n9821), .B2(n5737), .ZN(n5588)
         );
  XNOR2_X1 U7191 ( .A(n5588), .B(n5783), .ZN(n6768) );
  INV_X1 U7192 ( .A(n6768), .ZN(n6902) );
  OR2_X1 U7193 ( .A1(n9773), .A2(n5785), .ZN(n5590) );
  NAND2_X1 U7194 ( .A1(n9739), .A2(n4308), .ZN(n5589) );
  NAND2_X1 U7195 ( .A1(n5590), .A2(n5589), .ZN(n5592) );
  NAND2_X1 U7196 ( .A1(n6902), .A2(n5592), .ZN(n5591) );
  NAND2_X1 U7197 ( .A1(n5595), .A2(n5591), .ZN(n5598) );
  INV_X1 U7198 ( .A(n5592), .ZN(n6770) );
  AND2_X1 U7199 ( .A1(n6768), .A2(n6770), .ZN(n5596) );
  INV_X1 U7200 ( .A(n6903), .ZN(n5594) );
  INV_X1 U7201 ( .A(n6904), .ZN(n5593) );
  AOI22_X1 U7202 ( .A1(n5596), .A2(n5595), .B1(n5594), .B2(n5593), .ZN(n5597)
         );
  OAI21_X2 U7203 ( .B1(n6767), .B2(n5598), .A(n5597), .ZN(n6625) );
  OR2_X1 U7204 ( .A1(n9722), .A2(n5785), .ZN(n5600) );
  NAND2_X1 U7205 ( .A1(n6922), .A2(n4308), .ZN(n5599) );
  NAND2_X1 U7206 ( .A1(n5600), .A2(n5599), .ZN(n6622) );
  INV_X1 U7207 ( .A(n6622), .ZN(n5601) );
  NAND2_X1 U7208 ( .A1(n6625), .A2(n5601), .ZN(n5603) );
  OAI22_X1 U7209 ( .A1(n9722), .A2(n5739), .B1(n9837), .B2(n5737), .ZN(n5602)
         );
  XNOR2_X1 U7210 ( .A(n5602), .B(n8043), .ZN(n6623) );
  NAND2_X1 U7211 ( .A1(n5603), .A2(n6623), .ZN(n5606) );
  INV_X1 U7212 ( .A(n6625), .ZN(n5604) );
  NAND2_X1 U7213 ( .A1(n5604), .A2(n6622), .ZN(n5605) );
  NAND2_X1 U7214 ( .A1(n5606), .A2(n5605), .ZN(n6820) );
  OR2_X1 U7215 ( .A1(n7044), .A2(n5785), .ZN(n5608) );
  NAND2_X1 U7216 ( .A1(n6826), .A2(n4308), .ZN(n5607) );
  NAND2_X1 U7217 ( .A1(n5608), .A2(n5607), .ZN(n6822) );
  OAI22_X1 U7218 ( .A1(n7044), .A2(n5739), .B1(n9842), .B2(n5737), .ZN(n5609)
         );
  XNOR2_X1 U7219 ( .A(n5609), .B(n8043), .ZN(n6821) );
  OAI22_X1 U7220 ( .A1(n9721), .A2(n5739), .B1(n9850), .B2(n5737), .ZN(n5610)
         );
  XNOR2_X1 U7221 ( .A(n5610), .B(n5783), .ZN(n5612) );
  NOR2_X1 U7222 ( .A1(n9850), .A2(n5739), .ZN(n5611) );
  AOI21_X1 U7223 ( .B1(n9006), .B2(n8045), .A(n5611), .ZN(n5613) );
  NAND2_X1 U7224 ( .A1(n5612), .A2(n5613), .ZN(n5617) );
  INV_X1 U7225 ( .A(n5612), .ZN(n5615) );
  INV_X1 U7226 ( .A(n5613), .ZN(n5614) );
  NAND2_X1 U7227 ( .A1(n5615), .A2(n5614), .ZN(n5616) );
  NAND2_X1 U7228 ( .A1(n5617), .A2(n5616), .ZN(n7039) );
  NAND2_X1 U7229 ( .A1(n7037), .A2(n5617), .ZN(n7129) );
  OAI22_X1 U7230 ( .A1(n6932), .A2(n5739), .B1(n9427), .B2(n5737), .ZN(n5618)
         );
  XNOR2_X1 U7231 ( .A(n5618), .B(n8043), .ZN(n5620) );
  OAI22_X1 U7232 ( .A1(n6932), .A2(n5785), .B1(n9427), .B2(n5739), .ZN(n5619)
         );
  NAND2_X1 U7233 ( .A1(n5620), .A2(n5619), .ZN(n7127) );
  NAND2_X1 U7234 ( .A1(n7129), .A2(n7127), .ZN(n5621) );
  OR2_X1 U7235 ( .A1(n5620), .A2(n5619), .ZN(n7128) );
  NAND2_X1 U7236 ( .A1(n5621), .A2(n7128), .ZN(n7222) );
  INV_X1 U7237 ( .A(n7222), .ZN(n5628) );
  NAND2_X1 U7238 ( .A1(n9490), .A2(n4308), .ZN(n5623) );
  NAND2_X1 U7239 ( .A1(n7226), .A2(n4310), .ZN(n5622) );
  NAND2_X1 U7240 ( .A1(n5623), .A2(n5622), .ZN(n5624) );
  XNOR2_X1 U7241 ( .A(n5624), .B(n5783), .ZN(n5629) );
  AND2_X1 U7242 ( .A1(n7226), .A2(n4308), .ZN(n5626) );
  AOI21_X1 U7243 ( .B1(n9490), .B2(n8045), .A(n5626), .ZN(n5630) );
  XNOR2_X1 U7244 ( .A(n5629), .B(n5630), .ZN(n7223) );
  INV_X1 U7245 ( .A(n7223), .ZN(n5627) );
  INV_X1 U7246 ( .A(n5629), .ZN(n5632) );
  INV_X1 U7247 ( .A(n5630), .ZN(n5631) );
  NAND2_X1 U7248 ( .A1(n5632), .A2(n5631), .ZN(n5633) );
  OAI22_X1 U7249 ( .A1(n5635), .A2(n5739), .B1(n9541), .B2(n5737), .ZN(n5634)
         );
  XNOR2_X1 U7250 ( .A(n5634), .B(n8043), .ZN(n5638) );
  OAI22_X1 U7251 ( .A1(n5635), .A2(n5785), .B1(n9541), .B2(n5739), .ZN(n5637)
         );
  XNOR2_X1 U7252 ( .A(n5638), .B(n5637), .ZN(n7261) );
  OR2_X1 U7253 ( .A1(n5638), .A2(n5637), .ZN(n5639) );
  AND2_X2 U7254 ( .A1(n7258), .A2(n5639), .ZN(n8934) );
  OAI22_X1 U7255 ( .A1(n9532), .A2(n5737), .B1(n7264), .B2(n5739), .ZN(n5640)
         );
  XNOR2_X1 U7256 ( .A(n5640), .B(n5783), .ZN(n8936) );
  OR2_X1 U7257 ( .A1(n7264), .A2(n5785), .ZN(n5642) );
  OR2_X1 U7258 ( .A1(n9532), .A2(n5739), .ZN(n5641) );
  NAND2_X1 U7259 ( .A1(n8936), .A2(n8935), .ZN(n5643) );
  NAND2_X1 U7260 ( .A1(n8934), .A2(n5643), .ZN(n5647) );
  INV_X1 U7261 ( .A(n8936), .ZN(n5645) );
  INV_X1 U7262 ( .A(n8935), .ZN(n5644) );
  NAND2_X1 U7263 ( .A1(n5645), .A2(n5644), .ZN(n5646) );
  NAND2_X1 U7264 ( .A1(n8848), .A2(n4311), .ZN(n5649) );
  NAND2_X1 U7265 ( .A1(n9275), .A2(n4308), .ZN(n5648) );
  NAND2_X1 U7266 ( .A1(n5649), .A2(n5648), .ZN(n5650) );
  XNOR2_X1 U7267 ( .A(n5650), .B(n5783), .ZN(n8845) );
  AND2_X1 U7268 ( .A1(n9275), .A2(n8045), .ZN(n5651) );
  AOI21_X1 U7269 ( .B1(n8848), .B2(n4308), .A(n5651), .ZN(n8844) );
  NAND2_X1 U7270 ( .A1(n8845), .A2(n8844), .ZN(n5662) );
  NAND2_X1 U7271 ( .A1(n9286), .A2(n4310), .ZN(n5653) );
  NAND2_X1 U7272 ( .A1(n9262), .A2(n4308), .ZN(n5652) );
  NAND2_X1 U7273 ( .A1(n5653), .A2(n5652), .ZN(n5654) );
  XNOR2_X1 U7274 ( .A(n5654), .B(n5783), .ZN(n5661) );
  INV_X1 U7275 ( .A(n8845), .ZN(n5656) );
  INV_X1 U7276 ( .A(n8844), .ZN(n5655) );
  NAND2_X1 U7277 ( .A1(n5656), .A2(n5655), .ZN(n5660) );
  AND2_X1 U7278 ( .A1(n5661), .A2(n5660), .ZN(n5657) );
  NAND2_X1 U7279 ( .A1(n9286), .A2(n4308), .ZN(n5659) );
  NAND2_X1 U7280 ( .A1(n9262), .A2(n8045), .ZN(n5658) );
  NAND2_X1 U7281 ( .A1(n5659), .A2(n5658), .ZN(n8985) );
  INV_X1 U7282 ( .A(n5661), .ZN(n5663) );
  AND2_X1 U7283 ( .A1(n5663), .A2(n5662), .ZN(n5664) );
  NAND2_X1 U7284 ( .A1(n8894), .A2(n4311), .ZN(n5666) );
  NAND2_X1 U7285 ( .A1(n9276), .A2(n4308), .ZN(n5665) );
  NAND2_X1 U7286 ( .A1(n5666), .A2(n5665), .ZN(n5667) );
  XNOR2_X1 U7287 ( .A(n5667), .B(n5783), .ZN(n5670) );
  NOR2_X1 U7288 ( .A1(n5668), .A2(n5785), .ZN(n5669) );
  AOI21_X1 U7289 ( .B1(n8894), .B2(n4308), .A(n5669), .ZN(n5671) );
  NAND2_X1 U7290 ( .A1(n5670), .A2(n5671), .ZN(n5675) );
  INV_X1 U7291 ( .A(n5670), .ZN(n5673) );
  INV_X1 U7292 ( .A(n5671), .ZN(n5672) );
  NAND2_X1 U7293 ( .A1(n5673), .A2(n5672), .ZN(n5674) );
  AND2_X1 U7294 ( .A1(n5675), .A2(n5674), .ZN(n8897) );
  NAND2_X1 U7295 ( .A1(n8895), .A2(n5675), .ZN(n8907) );
  NAND2_X1 U7296 ( .A1(n9359), .A2(n4310), .ZN(n5677) );
  NAND2_X1 U7297 ( .A1(n9261), .A2(n4308), .ZN(n5676) );
  NAND2_X1 U7298 ( .A1(n5677), .A2(n5676), .ZN(n5678) );
  XNOR2_X1 U7299 ( .A(n5678), .B(n8043), .ZN(n5680) );
  AND2_X1 U7300 ( .A1(n9261), .A2(n8045), .ZN(n5679) );
  AOI21_X1 U7301 ( .B1(n9359), .B2(n4308), .A(n5679), .ZN(n5681) );
  XNOR2_X1 U7302 ( .A(n5680), .B(n5681), .ZN(n8908) );
  NAND2_X1 U7303 ( .A1(n8907), .A2(n8908), .ZN(n8906) );
  INV_X1 U7304 ( .A(n5680), .ZN(n5682) );
  NAND2_X1 U7305 ( .A1(n5682), .A2(n5681), .ZN(n5683) );
  NAND2_X1 U7306 ( .A1(n9350), .A2(n4311), .ZN(n5685) );
  NAND2_X1 U7307 ( .A1(n9230), .A2(n4308), .ZN(n5684) );
  NAND2_X1 U7308 ( .A1(n5685), .A2(n5684), .ZN(n5686) );
  XNOR2_X1 U7309 ( .A(n5686), .B(n8043), .ZN(n5697) );
  NAND2_X1 U7310 ( .A1(n9350), .A2(n4308), .ZN(n5688) );
  NAND2_X1 U7311 ( .A1(n9230), .A2(n8045), .ZN(n5687) );
  NAND2_X1 U7312 ( .A1(n5688), .A2(n5687), .ZN(n5698) );
  NAND2_X1 U7313 ( .A1(n5697), .A2(n5698), .ZN(n8871) );
  NAND2_X1 U7314 ( .A1(n9356), .A2(n4310), .ZN(n5690) );
  NAND2_X1 U7315 ( .A1(n9248), .A2(n4308), .ZN(n5689) );
  NAND2_X1 U7316 ( .A1(n5690), .A2(n5689), .ZN(n5691) );
  XNOR2_X1 U7317 ( .A(n5691), .B(n5783), .ZN(n8869) );
  NOR2_X1 U7318 ( .A1(n8911), .A2(n5785), .ZN(n5692) );
  AOI21_X1 U7319 ( .B1(n9356), .B2(n4308), .A(n5692), .ZN(n8974) );
  NOR2_X1 U7320 ( .A1(n8869), .A2(n8974), .ZN(n5693) );
  INV_X1 U7321 ( .A(n8869), .ZN(n8867) );
  INV_X1 U7322 ( .A(n8974), .ZN(n5696) );
  NOR2_X1 U7323 ( .A1(n8867), .A2(n5696), .ZN(n5701) );
  INV_X1 U7324 ( .A(n5697), .ZN(n5700) );
  INV_X1 U7325 ( .A(n5698), .ZN(n5699) );
  AOI21_X1 U7326 ( .B1(n5701), .B2(n8871), .A(n8925), .ZN(n5708) );
  NAND2_X1 U7327 ( .A1(n9344), .A2(n4310), .ZN(n5703) );
  NAND2_X1 U7328 ( .A1(n9216), .A2(n4308), .ZN(n5702) );
  NAND2_X1 U7329 ( .A1(n5703), .A2(n5702), .ZN(n5704) );
  XNOR2_X1 U7330 ( .A(n5704), .B(n5783), .ZN(n5707) );
  AND2_X1 U7331 ( .A1(n9216), .A2(n8045), .ZN(n5705) );
  AOI21_X1 U7332 ( .B1(n9344), .B2(n4308), .A(n5705), .ZN(n5706) );
  NAND2_X1 U7333 ( .A1(n5707), .A2(n5706), .ZN(n5710) );
  OAI21_X1 U7334 ( .B1(n5707), .B2(n5706), .A(n5710), .ZN(n8923) );
  NAND2_X1 U7335 ( .A1(n9185), .A2(n4311), .ZN(n5712) );
  OR2_X1 U7336 ( .A1(n8955), .A2(n5739), .ZN(n5711) );
  NAND2_X1 U7337 ( .A1(n5712), .A2(n5711), .ZN(n5713) );
  XNOR2_X1 U7338 ( .A(n5713), .B(n8043), .ZN(n5714) );
  OAI22_X1 U7339 ( .A1(n9339), .A2(n5739), .B1(n8955), .B2(n5785), .ZN(n5715)
         );
  XNOR2_X1 U7340 ( .A(n5714), .B(n5715), .ZN(n8878) );
  INV_X1 U7341 ( .A(n5714), .ZN(n5717) );
  INV_X1 U7342 ( .A(n5715), .ZN(n5716) );
  OAI22_X1 U7343 ( .A1(n9164), .A2(n5739), .B1(n8882), .B2(n5785), .ZN(n5722)
         );
  NAND2_X1 U7344 ( .A1(n5718), .A2(n5722), .ZN(n8948) );
  NAND2_X1 U7345 ( .A1(n9327), .A2(n4310), .ZN(n5720) );
  NAND2_X1 U7346 ( .A1(n9167), .A2(n4308), .ZN(n5719) );
  NAND2_X1 U7347 ( .A1(n5720), .A2(n5719), .ZN(n5721) );
  XNOR2_X1 U7348 ( .A(n5721), .B(n5783), .ZN(n5726) );
  INV_X1 U7349 ( .A(n5722), .ZN(n5723) );
  OAI22_X1 U7350 ( .A1(n9164), .A2(n5737), .B1(n8882), .B2(n5739), .ZN(n5725)
         );
  XNOR2_X1 U7351 ( .A(n5725), .B(n8043), .ZN(n8949) );
  NAND2_X1 U7352 ( .A1(n8947), .A2(n8949), .ZN(n5727) );
  NAND3_X1 U7353 ( .A1(n8948), .A2(n5726), .A3(n5727), .ZN(n8857) );
  OAI22_X1 U7354 ( .A1(n9128), .A2(n5737), .B1(n8890), .B2(n5739), .ZN(n5728)
         );
  XNOR2_X1 U7355 ( .A(n5728), .B(n8043), .ZN(n5730) );
  OAI22_X1 U7356 ( .A1(n9128), .A2(n5739), .B1(n8890), .B2(n5785), .ZN(n5729)
         );
  NOR2_X1 U7357 ( .A1(n5730), .A2(n5729), .ZN(n5731) );
  AOI21_X1 U7358 ( .B1(n5730), .B2(n5729), .A(n5731), .ZN(n8917) );
  INV_X1 U7359 ( .A(n5731), .ZN(n5732) );
  OAI22_X1 U7360 ( .A1(n9119), .A2(n5739), .B1(n5733), .B2(n5785), .ZN(n5743)
         );
  NAND2_X1 U7361 ( .A1(n9317), .A2(n4311), .ZN(n5735) );
  NAND2_X1 U7362 ( .A1(n9131), .A2(n4308), .ZN(n5734) );
  NAND2_X1 U7363 ( .A1(n5735), .A2(n5734), .ZN(n5736) );
  XNOR2_X1 U7364 ( .A(n5736), .B(n8043), .ZN(n5742) );
  XOR2_X1 U7365 ( .A(n5743), .B(n5742), .Z(n8887) );
  OAI22_X1 U7366 ( .A1(n9104), .A2(n5737), .B1(n5796), .B2(n5739), .ZN(n5738)
         );
  XNOR2_X1 U7367 ( .A(n5738), .B(n5783), .ZN(n5778) );
  OR2_X1 U7368 ( .A1(n9104), .A2(n5739), .ZN(n5741) );
  NAND2_X1 U7369 ( .A1(n9122), .A2(n8045), .ZN(n5740) );
  NAND2_X1 U7370 ( .A1(n5741), .A2(n5740), .ZN(n5779) );
  XNOR2_X1 U7371 ( .A(n5778), .B(n5779), .ZN(n5748) );
  INV_X1 U7372 ( .A(n5742), .ZN(n5745) );
  INV_X1 U7373 ( .A(n5743), .ZN(n5744) );
  NAND2_X1 U7374 ( .A1(n5745), .A2(n5744), .ZN(n5749) );
  AOI21_X1 U7375 ( .B1(n5747), .B2(n5749), .A(n5748), .ZN(n5750) );
  INV_X1 U7376 ( .A(n5751), .ZN(n5752) );
  OR2_X1 U7377 ( .A1(n9827), .A2(n5753), .ZN(n5764) );
  INV_X1 U7378 ( .A(n6085), .ZN(n5758) );
  INV_X1 U7379 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5754) );
  NOR2_X1 U7380 ( .A1(n5755), .A2(n5754), .ZN(n5756) );
  OR2_X1 U7381 ( .A1(n9378), .A2(n5756), .ZN(n5757) );
  INV_X1 U7382 ( .A(n9791), .ZN(n6086) );
  NAND2_X1 U7383 ( .A1(n5769), .A2(n6086), .ZN(n5759) );
  NAND3_X1 U7384 ( .A1(n5791), .A2(n5760), .A3(n8977), .ZN(n5777) );
  NAND2_X1 U7385 ( .A1(n9740), .A2(n6086), .ZN(n5766) );
  INV_X1 U7386 ( .A(n5769), .ZN(n5984) );
  INV_X1 U7387 ( .A(n5762), .ZN(n9102) );
  AND3_X1 U7388 ( .A1(n6088), .A2(n5841), .A3(n6985), .ZN(n5763) );
  OAI21_X1 U7389 ( .B1(n5764), .B2(n5769), .A(n5763), .ZN(n5765) );
  NAND2_X1 U7390 ( .A1(n5765), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5768) );
  NOR2_X1 U7391 ( .A1(n6092), .A2(n9791), .ZN(n5770) );
  INV_X1 U7392 ( .A(n5770), .ZN(n7493) );
  NAND2_X1 U7393 ( .A1(n7493), .A2(n5766), .ZN(n5767) );
  NAND2_X1 U7394 ( .A1(n5767), .A2(n5984), .ZN(n5986) );
  NAND2_X1 U7395 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  AOI22_X1 U7396 ( .A1(n8966), .A2(n9131), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n5772) );
  OAI21_X1 U7397 ( .B1(n9003), .B2(n8953), .A(n5772), .ZN(n5773) );
  AOI21_X1 U7398 ( .B1(n9102), .B2(n8997), .A(n5773), .ZN(n5774) );
  INV_X1 U7399 ( .A(n5775), .ZN(n5776) );
  NAND2_X1 U7400 ( .A1(n5777), .A2(n5776), .ZN(P1_U3238) );
  INV_X1 U7401 ( .A(n5778), .ZN(n5780) );
  INV_X1 U7402 ( .A(n5792), .ZN(n5790) );
  NAND2_X1 U7403 ( .A1(n9307), .A2(n4311), .ZN(n5782) );
  OR2_X1 U7404 ( .A1(n9003), .A2(n5739), .ZN(n5781) );
  NAND2_X1 U7405 ( .A1(n5782), .A2(n5781), .ZN(n5784) );
  XNOR2_X1 U7406 ( .A(n5784), .B(n5783), .ZN(n5788) );
  NOR2_X1 U7407 ( .A1(n9003), .A2(n5785), .ZN(n5786) );
  AOI21_X1 U7408 ( .B1(n9307), .B2(n5625), .A(n5786), .ZN(n5787) );
  NAND2_X1 U7409 ( .A1(n5788), .A2(n5787), .ZN(n8053) );
  OAI21_X1 U7410 ( .B1(n5788), .B2(n5787), .A(n8053), .ZN(n5793) );
  INV_X1 U7411 ( .A(n5793), .ZN(n5789) );
  AOI21_X1 U7412 ( .B1(n5791), .B2(n5790), .A(n5789), .ZN(n5794) );
  OAI21_X1 U7413 ( .B1(n5794), .B2(n8060), .A(n8977), .ZN(n5802) );
  OAI22_X1 U7414 ( .A1(n5796), .A2(n8994), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5795), .ZN(n5798) );
  NOR2_X1 U7415 ( .A1(n9090), .A2(n8953), .ZN(n5797) );
  AOI211_X1 U7416 ( .C1(n9087), .C2(n8997), .A(n5798), .B(n5797), .ZN(n5799)
         );
  INV_X1 U7417 ( .A(n5800), .ZN(n5801) );
  NAND2_X1 U7418 ( .A1(n5802), .A2(n5801), .ZN(P1_U3212) );
  NOR2_X2 U7419 ( .A1(n5891), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5893) );
  NAND4_X1 U7420 ( .A1(n5808), .A2(n5807), .A3(n5945), .A4(n5806), .ZN(n5811)
         );
  NAND4_X1 U7421 ( .A1(n6189), .A2(n5944), .A3(n5950), .A4(n5809), .ZN(n5810)
         );
  NOR3_X1 U7422 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .A3(
        P2_IR_REG_21__SCAN_IN), .ZN(n5822) );
  NOR2_X1 U7423 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5821) );
  NOR2_X1 U7424 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5820) );
  NOR2_X1 U7425 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5819) );
  NAND4_X1 U7426 ( .A1(n5822), .A2(n5821), .A3(n5820), .A4(n5819), .ZN(n5823)
         );
  NOR2_X1 U7427 ( .A1(n5828), .A2(n5919), .ZN(n5825) );
  MUX2_X1 U7428 ( .A(n5919), .B(n5825), .S(P2_IR_REG_25__SCAN_IN), .Z(n5826)
         );
  INV_X1 U7429 ( .A(n5826), .ZN(n5829) );
  NAND2_X1 U7430 ( .A1(n5829), .A2(n5831), .ZN(n8839) );
  INV_X1 U7431 ( .A(n8839), .ZN(n5834) );
  NAND2_X1 U7432 ( .A1(n5831), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5830) );
  MUX2_X1 U7433 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5830), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5833) );
  INV_X1 U7434 ( .A(n5935), .ZN(n5832) );
  NAND2_X1 U7435 ( .A1(n5834), .A2(n6030), .ZN(n5835) );
  OR2_X1 U7436 ( .A1(n5837), .A2(n5836), .ZN(n5838) );
  NAND2_X1 U7437 ( .A1(n5839), .A2(n5838), .ZN(n6158) );
  INV_X1 U7438 ( .A(n9912), .ZN(n5840) );
  INV_X1 U7439 ( .A(n6985), .ZN(n5842) );
  OR2_X1 U7440 ( .A1(n7756), .A2(n5842), .ZN(n5843) );
  NAND2_X1 U7441 ( .A1(n5843), .A2(n5872), .ZN(n5859) );
  NAND2_X1 U7442 ( .A1(n9569), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AND2_X1 U7443 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7040) );
  NOR2_X1 U7444 ( .A1(n9624), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5845) );
  AOI21_X1 U7445 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9624), .A(n5845), .ZN(
        n9617) );
  NOR2_X1 U7446 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n5902), .ZN(n5846) );
  AOI21_X1 U7447 ( .B1(n5902), .B2(P1_REG2_REG_7__SCAN_IN), .A(n5846), .ZN(
        n6010) );
  INV_X1 U7448 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U7449 ( .A1(n9577), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U7450 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9585) );
  INV_X1 U7451 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5848) );
  MUX2_X1 U7452 ( .A(n5848), .B(P1_REG2_REG_1__SCAN_IN), .S(n9577), .Z(n9584)
         );
  NOR2_X1 U7453 ( .A1(n9585), .A2(n9584), .ZN(n9583) );
  INV_X1 U7454 ( .A(n9583), .ZN(n5849) );
  NAND2_X1 U7455 ( .A1(n5850), .A2(n5849), .ZN(n9020) );
  NAND2_X1 U7456 ( .A1(n9018), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U7457 ( .A1(n9024), .A2(n5851), .ZN(n6081) );
  INV_X1 U7458 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6690) );
  MUX2_X1 U7459 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6690), .S(n5888), .Z(n6082)
         );
  NAND2_X1 U7460 ( .A1(n6081), .A2(n6082), .ZN(n6080) );
  NAND2_X1 U7461 ( .A1(n5888), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U7462 ( .A1(n6080), .A2(n5852), .ZN(n6237) );
  MUX2_X1 U7463 ( .A(n4961), .B(P1_REG2_REG_4__SCAN_IN), .S(n6242), .Z(n6238)
         );
  NOR2_X1 U7464 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9599), .ZN(n5853) );
  AOI21_X1 U7465 ( .B1(n9599), .B2(P1_REG2_REG_5__SCAN_IN), .A(n5853), .ZN(
        n9597) );
  OAI21_X1 U7466 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n9599), .A(n9595), .ZN(
        n9609) );
  INV_X1 U7467 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6837) );
  MUX2_X1 U7468 ( .A(n6837), .B(P1_REG2_REG_6__SCAN_IN), .S(n9602), .Z(n9608)
         );
  NOR2_X1 U7469 ( .A1(n9609), .A2(n9608), .ZN(n9607) );
  OAI21_X1 U7470 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9624), .A(n9615), .ZN(
        n5857) );
  NAND2_X1 U7471 ( .A1(n5998), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5854) );
  OAI21_X1 U7472 ( .B1(n5998), .B2(P1_REG2_REG_9__SCAN_IN), .A(n5854), .ZN(
        n5856) );
  NOR2_X1 U7473 ( .A1(n5856), .A2(n5857), .ZN(n5997) );
  INV_X1 U7474 ( .A(n7492), .ZN(n9567) );
  NAND2_X1 U7475 ( .A1(n9567), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9392) );
  INV_X1 U7476 ( .A(n9052), .ZN(n5855) );
  AOI211_X1 U7477 ( .C1(n5857), .C2(n5856), .A(n5997), .B(n9665), .ZN(n5876)
         );
  NOR2_X1 U7478 ( .A1(n5532), .A2(P1_U3084), .ZN(n9387) );
  NAND2_X1 U7479 ( .A1(n9387), .A2(n7492), .ZN(n5858) );
  NOR2_X1 U7480 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n5902), .ZN(n5860) );
  AOI21_X1 U7481 ( .B1(n5902), .B2(P1_REG1_REG_7__SCAN_IN), .A(n5860), .ZN(
        n6013) );
  INV_X1 U7482 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9862) );
  MUX2_X1 U7483 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9862), .S(n9018), .Z(n9014)
         );
  INV_X1 U7484 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9860) );
  MUX2_X1 U7485 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9860), .S(n9577), .Z(n9578)
         );
  NAND2_X1 U7486 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9582) );
  INV_X1 U7487 ( .A(n9582), .ZN(n5861) );
  NAND2_X1 U7488 ( .A1(n9578), .A2(n5861), .ZN(n9579) );
  NAND2_X1 U7489 ( .A1(n9577), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U7490 ( .A1(n9579), .A2(n5862), .ZN(n9013) );
  NAND2_X1 U7491 ( .A1(n9014), .A2(n9013), .ZN(n9012) );
  NAND2_X1 U7492 ( .A1(n9018), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U7493 ( .A1(n9012), .A2(n5863), .ZN(n6074) );
  INV_X1 U7494 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9864) );
  MUX2_X1 U7495 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9864), .S(n5888), .Z(n6075)
         );
  NAND2_X1 U7496 ( .A1(n6074), .A2(n6075), .ZN(n6073) );
  NAND2_X1 U7497 ( .A1(n5888), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U7498 ( .A1(n6073), .A2(n5864), .ZN(n6232) );
  INV_X1 U7499 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9866) );
  MUX2_X1 U7500 ( .A(n9866), .B(P1_REG1_REG_4__SCAN_IN), .S(n6242), .Z(n6233)
         );
  NOR2_X1 U7501 ( .A1(n6232), .A2(n6233), .ZN(n6231) );
  INV_X1 U7502 ( .A(n6231), .ZN(n5865) );
  OAI21_X1 U7503 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n6242), .A(n5865), .ZN(
        n9592) );
  NAND2_X1 U7504 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9599), .ZN(n5866) );
  OAI21_X1 U7505 ( .B1(n9599), .B2(P1_REG1_REG_5__SCAN_IN), .A(n5866), .ZN(
        n9591) );
  NOR2_X1 U7506 ( .A1(n9592), .A2(n9591), .ZN(n9590) );
  AOI21_X1 U7507 ( .B1(n9599), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9590), .ZN(
        n9606) );
  NOR2_X1 U7508 ( .A1(n9602), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5867) );
  AOI21_X1 U7509 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n9602), .A(n5867), .ZN(
        n9605) );
  NAND2_X1 U7510 ( .A1(n9606), .A2(n9605), .ZN(n9604) );
  OAI21_X1 U7511 ( .B1(n9602), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9604), .ZN(
        n6012) );
  NAND2_X1 U7512 ( .A1(n6013), .A2(n6012), .ZN(n6011) );
  OR2_X1 U7513 ( .A1(n5902), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7514 ( .A1(n6011), .A2(n5868), .ZN(n9623) );
  NAND2_X1 U7515 ( .A1(n9624), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5869) );
  NOR2_X1 U7516 ( .A1(n9624), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9619) );
  AOI21_X1 U7517 ( .B1(n9623), .B2(n5869), .A(n9619), .ZN(n9618) );
  INV_X1 U7518 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9877) );
  INV_X1 U7519 ( .A(n5998), .ZN(n5993) );
  AOI22_X1 U7520 ( .A1(n5998), .A2(n9877), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n5993), .ZN(n5870) );
  NOR2_X1 U7521 ( .A1(n9618), .A2(n5870), .ZN(n5992) );
  AOI21_X1 U7522 ( .B1(n9618), .B2(n5870), .A(n5992), .ZN(n5871) );
  NOR2_X1 U7523 ( .A1(n9708), .A2(n5871), .ZN(n5875) );
  INV_X1 U7524 ( .A(n5872), .ZN(n5873) );
  INV_X1 U7525 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10058) );
  NAND2_X1 U7526 ( .A1(n9052), .A2(n5532), .ZN(n9702) );
  OAI22_X1 U7527 ( .A1(n9711), .A2(n10058), .B1(n5993), .B2(n9702), .ZN(n5874)
         );
  OR4_X1 U7528 ( .A1(n7040), .A2(n5876), .A3(n5875), .A4(n5874), .ZN(P1_U3250)
         );
  AND2_X1 U7529 ( .A1(n6103), .A2(P2_U3152), .ZN(n6204) );
  INV_X2 U7530 ( .A(n6204), .ZN(n8827) );
  NAND2_X1 U7531 ( .A1(n7501), .A2(P2_U3152), .ZN(n8840) );
  OR2_X1 U7532 ( .A1(n5877), .A2(n5919), .ZN(n5879) );
  INV_X1 U7533 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5878) );
  XNOR2_X1 U7534 ( .A(n5879), .B(n5878), .ZN(n6272) );
  OAI222_X1 U7535 ( .A1(n8827), .A2(n6121), .B1(n8840), .B2(n6122), .C1(
        P2_U3152), .C2(n6272), .ZN(P2_U3356) );
  INV_X1 U7536 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U7537 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4350), .ZN(n5880) );
  XNOR2_X1 U7538 ( .A(n5881), .B(n5880), .ZN(n6336) );
  OAI222_X1 U7539 ( .A1(n8827), .A2(n6135), .B1(n8840), .B2(n6134), .C1(
        P2_U3152), .C2(n6336), .ZN(P2_U3355) );
  INV_X1 U7540 ( .A(n5882), .ZN(n6105) );
  NAND2_X1 U7541 ( .A1(n7501), .A2(P1_U3084), .ZN(n9401) );
  AOI22_X1 U7542 ( .A1(n9390), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n9577), .ZN(n5883) );
  OAI21_X1 U7543 ( .B1(n6105), .B2(n9397), .A(n5883), .ZN(P1_U3352) );
  AOI22_X1 U7544 ( .A1(n9390), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n9018), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n5884) );
  OAI21_X1 U7545 ( .B1(n6122), .B2(n9397), .A(n5884), .ZN(P1_U3351) );
  AOI22_X1 U7546 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6242), .B1(n9390), .B2(
        P2_DATAO_REG_4__SCAN_IN), .ZN(n5885) );
  OAI21_X1 U7547 ( .B1(n6149), .B2(n9397), .A(n5885), .ZN(P1_U3349) );
  NAND2_X1 U7548 ( .A1(n5886), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5887) );
  XNOR2_X1 U7549 ( .A(n5887), .B(n5803), .ZN(n6290) );
  OAI222_X1 U7550 ( .A1(n8827), .A2(n6150), .B1(n8840), .B2(n6149), .C1(
        P2_U3152), .C2(n6290), .ZN(P2_U3354) );
  INV_X1 U7551 ( .A(n5888), .ZN(n6078) );
  OAI222_X1 U7552 ( .A1(n9401), .A2(n5889), .B1(n9397), .B2(n6134), .C1(
        P1_U3084), .C2(n6078), .ZN(P1_U3350) );
  AOI22_X1 U7553 ( .A1(n9599), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9390), .ZN(n5890) );
  OAI21_X1 U7554 ( .B1(n6208), .B2(n9397), .A(n5890), .ZN(P1_U3348) );
  NAND2_X1 U7555 ( .A1(n5891), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5892) );
  MUX2_X1 U7556 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5892), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5895) );
  INV_X1 U7557 ( .A(n5893), .ZN(n5894) );
  INV_X1 U7558 ( .A(n6304), .ZN(n6295) );
  OAI222_X1 U7559 ( .A1(n8827), .A2(n6209), .B1(n8840), .B2(n6208), .C1(
        P2_U3152), .C2(n6295), .ZN(P2_U3353) );
  INV_X1 U7560 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6104) );
  INV_X1 U7561 ( .A(n8840), .ZN(n7034) );
  INV_X1 U7562 ( .A(n7034), .ZN(n8835) );
  INV_X1 U7563 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5896) );
  OAI222_X1 U7564 ( .A1(n8827), .A2(n6104), .B1(n8835), .B2(n6105), .C1(
        P2_U3152), .C2(n6271), .ZN(P2_U3357) );
  AOI22_X1 U7565 ( .A1(n9602), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9390), .ZN(n5897) );
  OAI21_X1 U7566 ( .B1(n6406), .B2(n9397), .A(n5897), .ZN(P1_U3347) );
  OR2_X1 U7567 ( .A1(n5893), .A2(n5919), .ZN(n5898) );
  XNOR2_X1 U7568 ( .A(n5898), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6315) );
  INV_X1 U7569 ( .A(n6315), .ZN(n6410) );
  OAI222_X1 U7570 ( .A1(n8827), .A2(n6407), .B1(n8840), .B2(n6406), .C1(
        P2_U3152), .C2(n6410), .ZN(P2_U3352) );
  AOI22_X1 U7571 ( .A1(n9624), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9390), .ZN(n5899) );
  OAI21_X1 U7572 ( .B1(n6594), .B2(n9397), .A(n5899), .ZN(P1_U3345) );
  INV_X1 U7573 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6497) );
  INV_X1 U7574 ( .A(n6496), .ZN(n5903) );
  OR2_X1 U7575 ( .A1(n5900), .A2(n5919), .ZN(n5901) );
  XNOR2_X1 U7576 ( .A(n5901), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6345) );
  INV_X1 U7577 ( .A(n6345), .ZN(n6500) );
  OAI222_X1 U7578 ( .A1(n8827), .A2(n6497), .B1(n8835), .B2(n5903), .C1(
        P2_U3152), .C2(n6500), .ZN(P2_U3351) );
  OAI222_X1 U7579 ( .A1(n9401), .A2(n8784), .B1(n9397), .B2(n5903), .C1(
        P1_U3084), .C2(n4521), .ZN(P1_U3346) );
  NAND2_X1 U7580 ( .A1(n5904), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5905) );
  XNOR2_X1 U7581 ( .A(n5905), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6595) );
  INV_X1 U7582 ( .A(n6595), .ZN(n6378) );
  OAI222_X1 U7583 ( .A1(n8827), .A2(n5906), .B1(n8840), .B2(n6594), .C1(
        P2_U3152), .C2(n6378), .ZN(P2_U3350) );
  INV_X1 U7584 ( .A(n6703), .ZN(n5915) );
  OAI222_X1 U7585 ( .A1(n9397), .A2(n5915), .B1(n5993), .B2(P1_U3084), .C1(
        n5907), .C2(n9401), .ZN(P1_U3344) );
  INV_X1 U7586 ( .A(n6000), .ZN(n6184) );
  OR2_X1 U7587 ( .A1(n5904), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U7588 ( .A1(n5947), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5910) );
  INV_X1 U7589 ( .A(n5910), .ZN(n5909) );
  NAND2_X1 U7590 ( .A1(n5909), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5911) );
  NAND2_X1 U7591 ( .A1(n5910), .A2(n5945), .ZN(n5928) );
  INV_X1 U7592 ( .A(n6792), .ZN(n6736) );
  NAND2_X1 U7593 ( .A1(n5913), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5914) );
  XNOR2_X1 U7594 ( .A(n5914), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6704) );
  INV_X1 U7595 ( .A(n6704), .ZN(n6361) );
  OAI222_X1 U7596 ( .A1(n8827), .A2(n5916), .B1(n8835), .B2(n5915), .C1(n6361), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  NAND2_X1 U7597 ( .A1(n5920), .A2(n5917), .ZN(n5922) );
  MUX2_X1 U7598 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5921), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5923) );
  NAND2_X1 U7599 ( .A1(n7832), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5926) );
  AND2_X2 U7600 ( .A1(n5977), .A2(n8829), .ZN(n6802) );
  NAND2_X1 U7601 ( .A1(n6802), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5925) );
  AND2_X2 U7602 ( .A1(n8824), .A2(n8829), .ZN(n7244) );
  NAND2_X1 U7603 ( .A1(n7244), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7604 ( .A1(n8175), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5927) );
  OAI21_X1 U7605 ( .B1(n8175), .B2(n8305), .A(n5927), .ZN(P2_U3582) );
  INV_X1 U7606 ( .A(n6845), .ZN(n5932) );
  NAND2_X1 U7607 ( .A1(n5928), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5929) );
  XNOR2_X1 U7608 ( .A(n5929), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8199) );
  AOI22_X1 U7609 ( .A1(n8199), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n6204), .ZN(n5930) );
  OAI21_X1 U7610 ( .B1(n5932), .B2(n8840), .A(n5930), .ZN(P2_U3347) );
  INV_X1 U7611 ( .A(n6455), .ZN(n6451) );
  OAI222_X1 U7612 ( .A1(n9397), .A2(n5932), .B1(n6451), .B2(P1_U3084), .C1(
        n5931), .C2(n9401), .ZN(P1_U3342) );
  NAND2_X1 U7613 ( .A1(n4338), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5934) );
  XNOR2_X2 U7614 ( .A(n5937), .B(n5936), .ZN(n6264) );
  NOR2_X1 U7615 ( .A1(n6157), .A2(n7369), .ZN(n5939) );
  OR2_X1 U7616 ( .A1(n9904), .A2(n5939), .ZN(n5942) );
  INV_X1 U7617 ( .A(n6158), .ZN(n5940) );
  NAND2_X1 U7618 ( .A1(n5940), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8030) );
  OR2_X1 U7619 ( .A1(n8030), .A2(n6501), .ZN(n5941) );
  NOR2_X1 U7620 ( .A1(n9898), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7621 ( .A(n6940), .ZN(n5953) );
  INV_X1 U7622 ( .A(n9030), .ZN(n9041) );
  OAI222_X1 U7623 ( .A1(n9401), .A2(n5943), .B1(n9397), .B2(n5953), .C1(
        P1_U3084), .C2(n9041), .ZN(P1_U3341) );
  NAND2_X1 U7624 ( .A1(n5945), .A2(n5944), .ZN(n5946) );
  NOR2_X1 U7625 ( .A1(n5951), .A2(n5919), .ZN(n5948) );
  MUX2_X1 U7626 ( .A(n5919), .B(n5948), .S(P2_IR_REG_12__SCAN_IN), .Z(n5949)
         );
  INV_X1 U7627 ( .A(n5949), .ZN(n5952) );
  NAND2_X1 U7628 ( .A1(n5951), .A2(n5950), .ZN(n5959) );
  INV_X1 U7629 ( .A(n6941), .ZN(n6779) );
  OAI222_X1 U7630 ( .A1(n8827), .A2(n5954), .B1(n8835), .B2(n5953), .C1(
        P2_U3152), .C2(n6779), .ZN(P2_U3346) );
  INV_X1 U7631 ( .A(n7058), .ZN(n5957) );
  NAND2_X1 U7632 ( .A1(n5959), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5955) );
  XNOR2_X1 U7633 ( .A(n5955), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7059) );
  AOI22_X1 U7634 ( .A1(n7059), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n6204), .ZN(n5956) );
  OAI21_X1 U7635 ( .B1(n5957), .B2(n8840), .A(n5956), .ZN(P2_U3345) );
  INV_X1 U7636 ( .A(n9634), .ZN(n9042) );
  OAI222_X1 U7637 ( .A1(n9401), .A2(n8710), .B1(n9042), .B2(P1_U3084), .C1(
        n9397), .C2(n5957), .ZN(P1_U3340) );
  INV_X1 U7638 ( .A(n7144), .ZN(n5961) );
  OAI222_X1 U7639 ( .A1(n9397), .A2(n5961), .B1(n9043), .B2(P1_U3084), .C1(
        n5958), .C2(n9401), .ZN(P1_U3339) );
  NAND2_X1 U7640 ( .A1(n5960), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6190) );
  XNOR2_X1 U7641 ( .A(n6190), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7306) );
  INV_X1 U7642 ( .A(n7306), .ZN(n7313) );
  OAI222_X1 U7643 ( .A1(n8827), .A2(n5962), .B1(n8835), .B2(n5961), .C1(n7313), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  NAND3_X1 U7644 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n6215) );
  INV_X1 U7645 ( .A(n6215), .ZN(n5963) );
  NAND2_X1 U7646 ( .A1(n5963), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6424) );
  INV_X1 U7647 ( .A(n6424), .ZN(n5964) );
  NAND2_X1 U7648 ( .A1(n5964), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6503) );
  INV_X1 U7649 ( .A(n6503), .ZN(n5965) );
  NAND2_X1 U7650 ( .A1(n5965), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6713) );
  INV_X1 U7651 ( .A(n6713), .ZN(n5967) );
  NAND2_X1 U7652 ( .A1(n5967), .A2(n5966), .ZN(n6800) );
  INV_X1 U7653 ( .A(n6949), .ZN(n5968) );
  NAND2_X1 U7654 ( .A1(n5968), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7063) );
  INV_X1 U7655 ( .A(n7063), .ZN(n5969) );
  NAND2_X1 U7656 ( .A1(n5969), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7153) );
  NAND2_X1 U7657 ( .A1(n5970), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7286) );
  INV_X1 U7658 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7373) );
  INV_X1 U7659 ( .A(n7405), .ZN(n5973) );
  NAND2_X1 U7660 ( .A1(n5973), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n7421) );
  INV_X1 U7661 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8128) );
  INV_X1 U7662 ( .A(n7437), .ZN(n5974) );
  NAND2_X1 U7663 ( .A1(n5974), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n7451) );
  INV_X1 U7664 ( .A(n7451), .ZN(n5975) );
  NAND2_X1 U7665 ( .A1(n5975), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n7467) );
  INV_X1 U7666 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7466) );
  INV_X1 U7667 ( .A(n7469), .ZN(n5976) );
  NAND2_X1 U7668 ( .A1(n5976), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n7479) );
  INV_X1 U7669 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7478) );
  INV_X1 U7670 ( .A(n7481), .ZN(n8309) );
  AND2_X2 U7671 ( .A1(n5978), .A2(n5977), .ZN(n6143) );
  INV_X1 U7672 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7673 ( .A1(n7244), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U7674 ( .A1(n6802), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5979) );
  OAI211_X1 U7675 ( .C1(n5981), .C2(n7485), .A(n5980), .B(n5979), .ZN(n5982)
         );
  AOI21_X1 U7676 ( .B1(n8309), .B2(n6143), .A(n5982), .ZN(n8326) );
  NAND2_X1 U7677 ( .A1(n8175), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5983) );
  OAI21_X1 U7678 ( .B1(n8326), .B2(n8175), .A(n5983), .ZN(P2_U3581) );
  NAND2_X1 U7679 ( .A1(n9849), .A2(n5984), .ZN(n5985) );
  NAND4_X1 U7680 ( .A1(n5986), .A2(n6086), .A3(n6088), .A4(n5985), .ZN(n8968)
         );
  INV_X1 U7681 ( .A(n8968), .ZN(n5991) );
  INV_X1 U7682 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6563) );
  XOR2_X1 U7683 ( .A(n5988), .B(n5987), .Z(n6228) );
  NAND2_X1 U7684 ( .A1(n6228), .A2(n8977), .ZN(n5990) );
  AOI22_X1 U7685 ( .A1(n8992), .A2(n5562), .B1(n8965), .B2(n6565), .ZN(n5989)
         );
  OAI211_X1 U7686 ( .C1(n5991), .C2(n6563), .A(n5990), .B(n5989), .ZN(P1_U3230) );
  INV_X1 U7687 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9432) );
  AOI21_X1 U7688 ( .B1(n5993), .B2(n9877), .A(n5992), .ZN(n6178) );
  AOI22_X1 U7689 ( .A1(n6000), .A2(n9432), .B1(P1_REG1_REG_10__SCAN_IN), .B2(
        n6184), .ZN(n6177) );
  NOR2_X1 U7690 ( .A1(n6178), .A2(n6177), .ZN(n6176) );
  AOI21_X1 U7691 ( .B1(n6184), .B2(n9432), .A(n6176), .ZN(n5995) );
  INV_X1 U7692 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9550) );
  AOI22_X1 U7693 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n6451), .B1(n6455), .B2(
        n9550), .ZN(n5994) );
  NOR2_X1 U7694 ( .A1(n5995), .A2(n5994), .ZN(n6450) );
  AOI21_X1 U7695 ( .B1(n5995), .B2(n5994), .A(n6450), .ZN(n6007) );
  INV_X1 U7696 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5996) );
  AOI22_X1 U7697 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6455), .B1(n6451), .B2(
        n5996), .ZN(n6002) );
  AOI21_X1 U7698 ( .B1(n5998), .B2(P1_REG2_REG_9__SCAN_IN), .A(n5997), .ZN(
        n6180) );
  NAND2_X1 U7699 ( .A1(n6000), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5999) );
  OAI21_X1 U7700 ( .B1(n6000), .B2(P1_REG2_REG_10__SCAN_IN), .A(n5999), .ZN(
        n6181) );
  NOR2_X1 U7701 ( .A1(n6180), .A2(n6181), .ZN(n6179) );
  AOI21_X1 U7702 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n6000), .A(n6179), .ZN(
        n6001) );
  NAND2_X1 U7703 ( .A1(n6002), .A2(n6001), .ZN(n6454) );
  OAI21_X1 U7704 ( .B1(n6002), .B2(n6001), .A(n6454), .ZN(n6005) );
  NAND2_X1 U7705 ( .A1(n9603), .A2(P1_ADDR_REG_11__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7706 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7224) );
  OAI211_X1 U7707 ( .C1(n9702), .C2(n6451), .A(n6003), .B(n7224), .ZN(n6004)
         );
  AOI21_X1 U7708 ( .B1(n9698), .B2(n6005), .A(n6004), .ZN(n6006) );
  OAI21_X1 U7709 ( .B1(n6007), .B2(n9708), .A(n6006), .ZN(P1_U3252) );
  INV_X1 U7710 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6019) );
  OAI21_X1 U7711 ( .B1(n6010), .B2(n6009), .A(n6008), .ZN(n6017) );
  OAI21_X1 U7712 ( .B1(n6013), .B2(n6012), .A(n6011), .ZN(n6014) );
  NOR2_X1 U7713 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5025), .ZN(n6627) );
  AOI21_X1 U7714 ( .B1(n9688), .B2(n6014), .A(n6627), .ZN(n6015) );
  OAI21_X1 U7715 ( .B1(n9702), .B2(n4521), .A(n6015), .ZN(n6016) );
  AOI21_X1 U7716 ( .B1(n9698), .B2(n6017), .A(n6016), .ZN(n6018) );
  OAI21_X1 U7717 ( .B1(n9711), .B2(n6019), .A(n6018), .ZN(P1_U3248) );
  INV_X1 U7718 ( .A(n6020), .ZN(n6025) );
  AOI21_X1 U7719 ( .B1(n6024), .B2(n6021), .A(n6022), .ZN(n6023) );
  AOI21_X1 U7720 ( .B1(n6025), .B2(n6024), .A(n6023), .ZN(n6028) );
  AOI22_X1 U7721 ( .A1(n8966), .A2(n5553), .B1(n8965), .B2(n7524), .ZN(n6027)
         );
  AOI22_X1 U7722 ( .A1(n8992), .A2(n4932), .B1(n8968), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6026) );
  OAI211_X1 U7723 ( .C1(n6028), .C2(n8988), .A(n6027), .B(n6026), .ZN(P1_U3220) );
  XNOR2_X1 U7724 ( .A(n7143), .B(P2_B_REG_SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7725 ( .A1(n6029), .A2(n8839), .ZN(n6031) );
  INV_X1 U7726 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9910) );
  NAND2_X1 U7727 ( .A1(n9903), .A2(n9910), .ZN(n6033) );
  AND2_X1 U7728 ( .A1(n8839), .A2(n8836), .ZN(n9911) );
  INV_X1 U7729 ( .A(n9911), .ZN(n6032) );
  INV_X1 U7730 ( .A(n8526), .ZN(n6045) );
  INV_X1 U7731 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9907) );
  NOR2_X1 U7732 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .ZN(
        n6037) );
  NOR4_X1 U7733 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n6036) );
  NOR4_X1 U7734 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n6035) );
  NOR4_X1 U7735 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n6034) );
  AND4_X1 U7736 ( .A1(n6037), .A2(n6036), .A3(n6035), .A4(n6034), .ZN(n6043)
         );
  NOR4_X1 U7737 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6041) );
  NOR4_X1 U7738 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6040) );
  NOR4_X1 U7739 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6039) );
  NOR4_X1 U7740 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6038) );
  AND4_X1 U7741 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), .ZN(n6042)
         );
  NAND2_X1 U7742 ( .A1(n6043), .A2(n6042), .ZN(n6044) );
  NAND2_X1 U7743 ( .A1(n9903), .A2(n6044), .ZN(n6382) );
  NAND3_X1 U7744 ( .A1(n6045), .A2(n8529), .A3(n6382), .ZN(n6063) );
  INV_X1 U7745 ( .A(n6048), .ZN(n6049) );
  NAND2_X1 U7746 ( .A1(n6049), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7747 ( .A1(n6063), .A2(n8525), .ZN(n6162) );
  NAND2_X1 U7748 ( .A1(n6109), .A2(n8481), .ZN(n6057) );
  NAND2_X1 U7749 ( .A1(n8026), .A2(n6262), .ZN(n6381) );
  NAND2_X1 U7750 ( .A1(n6162), .A2(n6381), .ZN(n8133) );
  INV_X1 U7751 ( .A(n8133), .ZN(n6072) );
  INV_X1 U7752 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6071) );
  OR2_X1 U7753 ( .A1(n6063), .A2(n8026), .ZN(n8129) );
  NAND2_X1 U7754 ( .A1(n7832), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U7755 ( .A1(n6143), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7756 ( .A1(n7244), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U7757 ( .A1(n6802), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6053) );
  INV_X1 U7758 ( .A(n6057), .ZN(n6159) );
  NOR2_X1 U7759 ( .A1(n9904), .A2(n9994), .ZN(n6058) );
  NAND2_X1 U7760 ( .A1(n7501), .A2(SI_0_), .ZN(n6060) );
  INV_X1 U7761 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7762 ( .A1(n6060), .A2(n6059), .ZN(n6062) );
  AND2_X1 U7763 ( .A1(n6062), .A2(n6061), .ZN(n8842) );
  MUX2_X1 U7764 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8842), .S(n6501), .Z(n9914) );
  AOI22_X1 U7765 ( .A1(n8154), .A2(n6387), .B1(n9886), .B2(n9914), .ZN(n6070)
         );
  NAND2_X1 U7766 ( .A1(n6143), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7767 ( .A1(n7832), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U7768 ( .A1(n7244), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7769 ( .A1(n6802), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7770 ( .A1(n6437), .A2(n7444), .ZN(n6112) );
  INV_X1 U7771 ( .A(n9914), .ZN(n6534) );
  OAI21_X1 U7772 ( .B1(n8038), .B2(n9913), .A(n6534), .ZN(n6068) );
  NAND3_X1 U7773 ( .A1(n8150), .A2(n6112), .A3(n6068), .ZN(n6069) );
  OAI211_X1 U7774 ( .C1(n6072), .C2(n6071), .A(n6070), .B(n6069), .ZN(P2_U3234) );
  AND2_X1 U7775 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6251) );
  INV_X1 U7776 ( .A(n6251), .ZN(n6077) );
  OAI211_X1 U7777 ( .C1(n6075), .C2(n6074), .A(n9688), .B(n6073), .ZN(n6076)
         );
  OAI211_X1 U7778 ( .C1(n9702), .C2(n6078), .A(n6077), .B(n6076), .ZN(n6079)
         );
  INV_X1 U7779 ( .A(n6079), .ZN(n6084) );
  OAI211_X1 U7780 ( .C1(n6082), .C2(n6081), .A(n9698), .B(n6080), .ZN(n6083)
         );
  OAI211_X1 U7781 ( .C1(n9711), .C2(n8626), .A(n6084), .B(n6083), .ZN(P1_U3244) );
  AND2_X1 U7782 ( .A1(n6086), .A2(n6085), .ZN(n6087) );
  OR2_X1 U7783 ( .A1(n9832), .A2(n7752), .ZN(n6089) );
  INV_X1 U7784 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6098) );
  INV_X1 U7785 ( .A(n6093), .ZN(n6096) );
  AND2_X1 U7786 ( .A1(n5553), .A2(n6582), .ZN(n7522) );
  NOR2_X1 U7787 ( .A1(n6577), .A2(n7522), .ZN(n7724) );
  INV_X1 U7788 ( .A(n6092), .ZN(n6094) );
  NOR3_X1 U7789 ( .A1(n7724), .A2(n6094), .A3(n6093), .ZN(n6095) );
  AOI21_X1 U7790 ( .B1(n9742), .B2(n5562), .A(n6095), .ZN(n6562) );
  OAI21_X1 U7791 ( .B1(n6582), .B2(n6096), .A(n6562), .ZN(n6101) );
  NAND2_X1 U7792 ( .A1(n6101), .A2(n9859), .ZN(n6097) );
  OAI21_X1 U7793 ( .B1(n9859), .B2(n6098), .A(n6097), .ZN(P1_U3454) );
  INV_X1 U7794 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9574) );
  NAND2_X1 U7795 ( .A1(n6101), .A2(n9879), .ZN(n6102) );
  OAI21_X1 U7796 ( .B1(n9879), .B2(n9574), .A(n6102), .ZN(P1_U3523) );
  OR2_X1 U7797 ( .A1(n6402), .A2(n9913), .ZN(n6115) );
  OR2_X1 U7798 ( .A1(n7825), .A2(n6104), .ZN(n6107) );
  NAND2_X1 U7799 ( .A1(n8027), .A2(n8481), .ZN(n6108) );
  NAND2_X1 U7800 ( .A1(n6108), .A2(n7836), .ZN(n6110) );
  XNOR2_X1 U7801 ( .A(n9920), .B(n7390), .ZN(n6113) );
  XNOR2_X1 U7802 ( .A(n6115), .B(n6113), .ZN(n8034) );
  OR2_X1 U7803 ( .A1(n7390), .A2(n9914), .ZN(n6111) );
  AND2_X1 U7804 ( .A1(n6112), .A2(n6111), .ZN(n8033) );
  INV_X1 U7805 ( .A(n6113), .ZN(n6114) );
  NAND2_X1 U7806 ( .A1(n6115), .A2(n6114), .ZN(n6116) );
  NAND2_X1 U7807 ( .A1(n8032), .A2(n6116), .ZN(n8135) );
  NAND2_X1 U7808 ( .A1(n6143), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7809 ( .A1(n7832), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7810 ( .A1(n7244), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U7811 ( .A1(n6802), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6117) );
  OR2_X1 U7812 ( .A1(n6550), .A2(n9913), .ZN(n6127) );
  OR2_X1 U7813 ( .A1(n4304), .A2(n6121), .ZN(n6124) );
  OR2_X1 U7814 ( .A1(n6790), .A2(n6122), .ZN(n6123) );
  XNOR2_X1 U7815 ( .A(n9929), .B(n7390), .ZN(n6125) );
  XNOR2_X1 U7816 ( .A(n6127), .B(n6125), .ZN(n8136) );
  NAND2_X1 U7817 ( .A1(n8135), .A2(n8136), .ZN(n8134) );
  INV_X1 U7818 ( .A(n6125), .ZN(n6126) );
  NAND2_X1 U7819 ( .A1(n6127), .A2(n6126), .ZN(n6128) );
  NAND2_X1 U7820 ( .A1(n8134), .A2(n6128), .ZN(n9884) );
  INV_X1 U7821 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7822 ( .A1(n6143), .A2(n6129), .ZN(n6133) );
  NAND2_X1 U7823 ( .A1(n7832), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7824 ( .A1(n7244), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7825 ( .A1(n6802), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6130) );
  OR2_X1 U7826 ( .A1(n6611), .A2(n9913), .ZN(n6138) );
  OR2_X1 U7827 ( .A1(n6790), .A2(n6134), .ZN(n6137) );
  OR2_X1 U7828 ( .A1(n4304), .A2(n6135), .ZN(n6136) );
  XNOR2_X1 U7829 ( .A(n9885), .B(n7798), .ZN(n6139) );
  XNOR2_X1 U7830 ( .A(n6138), .B(n6139), .ZN(n9883) );
  OR2_X1 U7831 ( .A1(n9884), .A2(n9883), .ZN(n9887) );
  INV_X1 U7832 ( .A(n6138), .ZN(n6141) );
  INV_X1 U7833 ( .A(n6139), .ZN(n6140) );
  NAND2_X1 U7834 ( .A1(n6141), .A2(n6140), .ZN(n6142) );
  NAND2_X1 U7835 ( .A1(n9887), .A2(n6142), .ZN(n6214) );
  NAND2_X1 U7836 ( .A1(n7832), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6148) );
  INV_X1 U7837 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6144) );
  XNOR2_X1 U7838 ( .A(n6144), .B(P2_REG3_REG_3__SCAN_IN), .ZN(n6615) );
  NAND2_X1 U7839 ( .A1(n6143), .A2(n6615), .ZN(n6147) );
  NAND2_X1 U7840 ( .A1(n7244), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7841 ( .A1(n6802), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6145) );
  OR2_X1 U7842 ( .A1(n6548), .A2(n9913), .ZN(n6154) );
  OR2_X1 U7843 ( .A1(n6790), .A2(n6149), .ZN(n6152) );
  OR2_X1 U7844 ( .A1(n4304), .A2(n6150), .ZN(n6151) );
  OAI211_X1 U7845 ( .C1(n6501), .C2(n6290), .A(n6152), .B(n6151), .ZN(n6616)
         );
  XNOR2_X1 U7846 ( .A(n6616), .B(n7798), .ZN(n6153) );
  NOR2_X1 U7847 ( .A1(n6154), .A2(n6153), .ZN(n6213) );
  NAND2_X1 U7848 ( .A1(n6154), .A2(n6153), .ZN(n6212) );
  INV_X1 U7849 ( .A(n6212), .ZN(n6155) );
  NOR2_X1 U7850 ( .A1(n6213), .A2(n6155), .ZN(n6156) );
  XNOR2_X1 U7851 ( .A(n6214), .B(n6156), .ZN(n6174) );
  OAI211_X1 U7852 ( .C1(n6159), .C2(n6385), .A(n6259), .B(n6158), .ZN(n6160)
         );
  INV_X1 U7853 ( .A(n6160), .ZN(n6161) );
  NAND2_X1 U7854 ( .A1(n6162), .A2(n6161), .ZN(n6163) );
  NAND2_X1 U7855 ( .A1(n7832), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6170) );
  INV_X1 U7856 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7857 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6164) );
  NAND2_X1 U7858 ( .A1(n6165), .A2(n6164), .ZN(n6166) );
  AND2_X1 U7859 ( .A1(n6215), .A2(n6166), .ZN(n6520) );
  NAND2_X1 U7860 ( .A1(n6143), .A2(n6520), .ZN(n6169) );
  NAND2_X1 U7861 ( .A1(n7244), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7862 ( .A1(n6802), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6167) );
  OAI22_X1 U7863 ( .A1(n6611), .A2(n8156), .B1(n8145), .B2(n6467), .ZN(n6172)
         );
  NAND2_X1 U7864 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n6268) );
  OAI21_X1 U7865 ( .B1(n8161), .B2(n9942), .A(n6268), .ZN(n6171) );
  AOI211_X1 U7866 ( .C1(n6615), .C2(n8158), .A(n6172), .B(n6171), .ZN(n6173)
         );
  OAI21_X1 U7867 ( .B1(n6174), .B2(n9882), .A(n6173), .ZN(P2_U3232) );
  INV_X1 U7868 ( .A(n7272), .ZN(n6199) );
  AOI22_X1 U7869 ( .A1(n9672), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9390), .ZN(n6175) );
  OAI21_X1 U7870 ( .B1(n6199), .B2(n9397), .A(n6175), .ZN(P1_U3337) );
  AOI21_X1 U7871 ( .B1(n6178), .B2(n6177), .A(n6176), .ZN(n6187) );
  AOI21_X1 U7872 ( .B1(n6181), .B2(n6180), .A(n6179), .ZN(n6182) );
  NAND2_X1 U7873 ( .A1(n9698), .A2(n6182), .ZN(n6183) );
  NAND2_X1 U7874 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7131) );
  OAI211_X1 U7875 ( .C1(n9702), .C2(n6184), .A(n6183), .B(n7131), .ZN(n6185)
         );
  AOI21_X1 U7876 ( .B1(n9603), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n6185), .ZN(
        n6186) );
  OAI21_X1 U7877 ( .B1(n6187), .B2(n9708), .A(n6186), .ZN(P1_U3251) );
  INV_X1 U7878 ( .A(n7236), .ZN(n6193) );
  OAI222_X1 U7879 ( .A1(n9401), .A2(n6188), .B1(n9397), .B2(n6193), .C1(
        P1_U3084), .C2(n9045), .ZN(P1_U3338) );
  NAND2_X1 U7880 ( .A1(n6190), .A2(n6189), .ZN(n6191) );
  NAND2_X1 U7881 ( .A1(n6191), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6192) );
  XNOR2_X1 U7882 ( .A(n6192), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8214) );
  INV_X1 U7883 ( .A(n8214), .ZN(n7314) );
  OAI222_X1 U7884 ( .A1(n8827), .A2(n6194), .B1(n8835), .B2(n6193), .C1(
        P2_U3152), .C2(n7314), .ZN(P2_U3343) );
  NAND2_X1 U7885 ( .A1(n5824), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6195) );
  MUX2_X1 U7886 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6195), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6197) );
  INV_X1 U7887 ( .A(n6200), .ZN(n6196) );
  NAND2_X1 U7888 ( .A1(n6197), .A2(n6196), .ZN(n8228) );
  OAI222_X1 U7889 ( .A1(P2_U3152), .A2(n8228), .B1(n8835), .B2(n6199), .C1(
        n6198), .C2(n8827), .ZN(P2_U3342) );
  INV_X1 U7890 ( .A(n7283), .ZN(n6207) );
  NOR2_X1 U7891 ( .A1(n6200), .A2(n5919), .ZN(n6201) );
  MUX2_X1 U7892 ( .A(n5919), .B(n6201), .S(P2_IR_REG_17__SCAN_IN), .Z(n6202)
         );
  INV_X1 U7893 ( .A(n6202), .ZN(n6203) );
  AND2_X1 U7894 ( .A1(n6203), .A2(n4396), .ZN(n8240) );
  AOI22_X1 U7895 ( .A1(n8240), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n6204), .ZN(n6205) );
  OAI21_X1 U7896 ( .B1(n6207), .B2(n8840), .A(n6205), .ZN(P2_U3341) );
  AOI22_X1 U7897 ( .A1(n9039), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9390), .ZN(n6206) );
  OAI21_X1 U7898 ( .B1(n6207), .B2(n9397), .A(n6206), .ZN(P1_U3336) );
  OR2_X1 U7899 ( .A1(n6467), .A2(n9913), .ZN(n6418) );
  OR2_X1 U7900 ( .A1(n4304), .A2(n6209), .ZN(n6210) );
  AND2_X1 U7901 ( .A1(n6210), .A2(n4851), .ZN(n6211) );
  XNOR2_X1 U7902 ( .A(n6476), .B(n7798), .ZN(n6419) );
  XNOR2_X1 U7903 ( .A(n6418), .B(n6419), .ZN(n6416) );
  OAI21_X1 U7904 ( .B1(n6214), .B2(n6213), .A(n6212), .ZN(n6417) );
  XOR2_X1 U7905 ( .A(n6416), .B(n6417), .Z(n6226) );
  INV_X1 U7906 ( .A(n6520), .ZN(n6224) );
  INV_X1 U7907 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U7908 ( .A1(n6215), .A2(n6302), .ZN(n6216) );
  AND2_X1 U7909 ( .A1(n6424), .A2(n6216), .ZN(n6479) );
  NAND2_X1 U7910 ( .A1(n6143), .A2(n6479), .ZN(n6220) );
  NAND2_X1 U7911 ( .A1(n7832), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7912 ( .A1(n7244), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U7913 ( .A1(n6802), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6217) );
  OR2_X1 U7914 ( .A1(n6548), .A2(n8455), .ZN(n6221) );
  OAI21_X1 U7915 ( .B1(n6657), .B2(n8457), .A(n6221), .ZN(n6517) );
  AND2_X1 U7916 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6287) );
  AOI21_X1 U7917 ( .B1(n9881), .B2(n6517), .A(n6287), .ZN(n6223) );
  NAND2_X1 U7918 ( .A1(n9886), .A2(n6476), .ZN(n6222) );
  OAI211_X1 U7919 ( .C1(n9891), .C2(n6224), .A(n6223), .B(n6222), .ZN(n6225)
         );
  AOI21_X1 U7920 ( .B1(n6226), .B2(n8150), .A(n6225), .ZN(n6227) );
  INV_X1 U7921 ( .A(n6227), .ZN(P2_U3229) );
  INV_X1 U7922 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6872) );
  MUX2_X1 U7923 ( .A(n6228), .B(n9585), .S(n9567), .Z(n6230) );
  OAI21_X1 U7924 ( .B1(n7492), .B2(P1_REG2_REG_0__SCAN_IN), .A(n6229), .ZN(
        n9565) );
  INV_X1 U7925 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9566) );
  NAND2_X1 U7926 ( .A1(n9565), .A2(n9566), .ZN(n9568) );
  OAI211_X1 U7927 ( .C1(n6230), .C2(n5532), .A(P1_U4006), .B(n9568), .ZN(n9028) );
  AOI21_X1 U7928 ( .B1(n6233), .B2(n6232), .A(n6231), .ZN(n6235) );
  AND2_X1 U7929 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n6489) );
  INV_X1 U7930 ( .A(n6489), .ZN(n6234) );
  OAI21_X1 U7931 ( .B1(n9708), .B2(n6235), .A(n6234), .ZN(n6241) );
  AOI21_X1 U7932 ( .B1(n6238), .B2(n6237), .A(n6236), .ZN(n6239) );
  NOR2_X1 U7933 ( .A1(n9665), .A2(n6239), .ZN(n6240) );
  AOI211_X1 U7934 ( .C1(n9671), .C2(n6242), .A(n6241), .B(n6240), .ZN(n6243)
         );
  OAI211_X1 U7935 ( .C1(n6872), .C2(n9711), .A(n9028), .B(n6243), .ZN(P1_U3245) );
  INV_X1 U7936 ( .A(n8997), .ZN(n6493) );
  INV_X1 U7937 ( .A(n6244), .ZN(n6246) );
  NOR2_X1 U7938 ( .A1(n6246), .A2(n6245), .ZN(n6247) );
  XNOR2_X1 U7939 ( .A(n6248), .B(n6247), .ZN(n6249) );
  NAND2_X1 U7940 ( .A1(n6249), .A2(n8977), .ZN(n6253) );
  OAI22_X1 U7941 ( .A1(n4934), .A2(n8994), .B1(n8953), .B2(n9748), .ZN(n6250)
         );
  AOI211_X1 U7942 ( .C1(n6692), .C2(n8965), .A(n6251), .B(n6250), .ZN(n6252)
         );
  OAI211_X1 U7943 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n6493), .A(n6253), .B(
        n6252), .ZN(P1_U3216) );
  INV_X1 U7944 ( .A(n6272), .ZN(n9419) );
  INV_X1 U7945 ( .A(n6271), .ZN(n9407) );
  INV_X1 U7946 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9901) );
  INV_X1 U7947 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9896) );
  INV_X1 U7948 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6254) );
  AOI21_X1 U7949 ( .B1(n9407), .B2(P2_REG2_REG_1__SCAN_IN), .A(n9403), .ZN(
        n9417) );
  INV_X1 U7950 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6255) );
  MUX2_X1 U7951 ( .A(n6255), .B(P2_REG2_REG_2__SCAN_IN), .S(n6272), .Z(n6256)
         );
  INV_X1 U7952 ( .A(n6256), .ZN(n9416) );
  AOI21_X1 U7953 ( .B1(n9419), .B2(P2_REG2_REG_2__SCAN_IN), .A(n9415), .ZN(
        n6329) );
  INV_X1 U7954 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6257) );
  MUX2_X1 U7955 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6257), .S(n6336), .Z(n6328)
         );
  NOR2_X1 U7956 ( .A1(n6329), .A2(n6328), .ZN(n6327) );
  INV_X1 U7957 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6258) );
  MUX2_X1 U7958 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6258), .S(n6290), .Z(n6265)
         );
  OAI21_X1 U7959 ( .B1(n6259), .B2(P2_U3152), .A(n8030), .ZN(n6260) );
  INV_X1 U7960 ( .A(n6260), .ZN(n6261) );
  NAND2_X1 U7961 ( .A1(n6262), .A2(n6261), .ZN(n6263) );
  NAND2_X1 U7962 ( .A1(n6263), .A2(n6501), .ZN(n6274) );
  NAND2_X1 U7963 ( .A1(n6274), .A2(n8175), .ZN(n6267) );
  INV_X1 U7964 ( .A(n6264), .ZN(n8270) );
  NAND2_X1 U7965 ( .A1(n6267), .A2(n8270), .ZN(n8262) );
  AOI211_X1 U7966 ( .C1(n6266), .C2(n6265), .A(n6282), .B(n9414), .ZN(n6281)
         );
  INV_X1 U7967 ( .A(n6268), .ZN(n6269) );
  AOI21_X1 U7968 ( .B1(n9898), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6269), .ZN(
        n6279) );
  INV_X1 U7969 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10010) );
  MUX2_X1 U7970 ( .A(n10010), .B(P2_REG1_REG_3__SCAN_IN), .S(n6336), .Z(n6332)
         );
  INV_X1 U7971 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6270) );
  MUX2_X1 U7972 ( .A(n6270), .B(P2_REG1_REG_2__SCAN_IN), .S(n6272), .Z(n9421)
         );
  INV_X1 U7973 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10007) );
  MUX2_X1 U7974 ( .A(n10007), .B(P2_REG1_REG_1__SCAN_IN), .S(n6271), .Z(n9409)
         );
  NAND3_X1 U7975 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n9409), .ZN(n9408) );
  OAI21_X1 U7976 ( .B1(n6271), .B2(n10007), .A(n9408), .ZN(n9422) );
  NAND2_X1 U7977 ( .A1(n9421), .A2(n9422), .ZN(n9420) );
  OAI21_X1 U7978 ( .B1(n6272), .B2(n6270), .A(n9420), .ZN(n6333) );
  NAND2_X1 U7979 ( .A1(n6332), .A2(n6333), .ZN(n6331) );
  OAI21_X1 U7980 ( .B1(n6336), .B2(n10010), .A(n6331), .ZN(n6277) );
  INV_X1 U7981 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6273) );
  MUX2_X1 U7982 ( .A(n6273), .B(P2_REG1_REG_4__SCAN_IN), .S(n6290), .Z(n6276)
         );
  INV_X1 U7983 ( .A(n6274), .ZN(n6275) );
  NAND2_X1 U7984 ( .A1(n6276), .A2(n6277), .ZN(n6289) );
  OAI211_X1 U7985 ( .C1(n6277), .C2(n6276), .A(n9892), .B(n6289), .ZN(n6278)
         );
  OAI211_X1 U7986 ( .C1(n8234), .C2(n6290), .A(n6279), .B(n6278), .ZN(n6280)
         );
  OR2_X1 U7987 ( .A1(n6281), .A2(n6280), .ZN(P2_U3249) );
  INV_X1 U7988 ( .A(n6290), .ZN(n6283) );
  NAND2_X1 U7989 ( .A1(n6304), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6284) );
  OAI21_X1 U7990 ( .B1(n6304), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6284), .ZN(
        n6285) );
  AOI211_X1 U7991 ( .C1(n6286), .C2(n6285), .A(n6298), .B(n9414), .ZN(n6297)
         );
  AOI21_X1 U7992 ( .B1(n9898), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6287), .ZN(
        n6294) );
  INV_X1 U7993 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6288) );
  MUX2_X1 U7994 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6288), .S(n6304), .Z(n6292)
         );
  OAI21_X1 U7995 ( .B1(n6290), .B2(n6273), .A(n6289), .ZN(n6291) );
  NAND2_X1 U7996 ( .A1(n6292), .A2(n6291), .ZN(n6305) );
  OAI211_X1 U7997 ( .C1(n6292), .C2(n6291), .A(n9892), .B(n6305), .ZN(n6293)
         );
  OAI211_X1 U7998 ( .C1(n8234), .C2(n6295), .A(n6294), .B(n6293), .ZN(n6296)
         );
  OR2_X1 U7999 ( .A1(n6297), .A2(n6296), .ZN(P2_U3250) );
  AOI21_X1 U8000 ( .B1(n6304), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6298), .ZN(
        n6301) );
  NAND2_X1 U8001 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(n6315), .ZN(n6299) );
  OAI21_X1 U8002 ( .B1(n6315), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6299), .ZN(
        n6300) );
  AOI211_X1 U8003 ( .C1(n6301), .C2(n6300), .A(n6314), .B(n9414), .ZN(n6313)
         );
  NOR2_X1 U8004 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6302), .ZN(n6303) );
  AOI21_X1 U8005 ( .B1(n9898), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6303), .ZN(
        n6311) );
  NAND2_X1 U8006 ( .A1(n6304), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U8007 ( .A1(n6306), .A2(n6305), .ZN(n6309) );
  INV_X1 U8008 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6307) );
  MUX2_X1 U8009 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6307), .S(n6315), .Z(n6308)
         );
  NAND2_X1 U8010 ( .A1(n6308), .A2(n6309), .ZN(n6320) );
  OAI211_X1 U8011 ( .C1(n6309), .C2(n6308), .A(n9892), .B(n6320), .ZN(n6310)
         );
  OAI211_X1 U8012 ( .C1(n8234), .C2(n6410), .A(n6311), .B(n6310), .ZN(n6312)
         );
  OR2_X1 U8013 ( .A1(n6313), .A2(n6312), .ZN(P2_U3251) );
  INV_X1 U8014 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6659) );
  MUX2_X1 U8015 ( .A(n6659), .B(P2_REG2_REG_7__SCAN_IN), .S(n6345), .Z(n6316)
         );
  AOI211_X1 U8016 ( .C1(n6317), .C2(n6316), .A(n6339), .B(n9414), .ZN(n6326)
         );
  INV_X1 U8017 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6509) );
  NOR2_X1 U8018 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6509), .ZN(n6318) );
  AOI21_X1 U8019 ( .B1(n9898), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6318), .ZN(
        n6324) );
  INV_X1 U8020 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6319) );
  MUX2_X1 U8021 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6319), .S(n6345), .Z(n6322)
         );
  OAI21_X1 U8022 ( .B1(n6410), .B2(n6307), .A(n6320), .ZN(n6321) );
  NAND2_X1 U8023 ( .A1(n6322), .A2(n6321), .ZN(n6346) );
  OAI211_X1 U8024 ( .C1(n6322), .C2(n6321), .A(n9892), .B(n6346), .ZN(n6323)
         );
  OAI211_X1 U8025 ( .C1(n8234), .C2(n6500), .A(n6324), .B(n6323), .ZN(n6325)
         );
  OR2_X1 U8026 ( .A1(n6326), .A2(n6325), .ZN(P2_U3252) );
  AOI211_X1 U8027 ( .C1(n6329), .C2(n6328), .A(n6327), .B(n9414), .ZN(n6338)
         );
  AND2_X1 U8028 ( .A1(P2_U3152), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6330) );
  AOI21_X1 U8029 ( .B1(n9898), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6330), .ZN(
        n6335) );
  OAI211_X1 U8030 ( .C1(n6333), .C2(n6332), .A(n9892), .B(n6331), .ZN(n6334)
         );
  OAI211_X1 U8031 ( .C1(n8234), .C2(n6336), .A(n6335), .B(n6334), .ZN(n6337)
         );
  OR2_X1 U8032 ( .A1(n6338), .A2(n6337), .ZN(P2_U3248) );
  NAND2_X1 U8033 ( .A1(n6595), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6340) );
  OAI21_X1 U8034 ( .B1(n6595), .B2(P2_REG2_REG_8__SCAN_IN), .A(n6340), .ZN(
        n6370) );
  AOI21_X1 U8035 ( .B1(n6595), .B2(P2_REG2_REG_8__SCAN_IN), .A(n6369), .ZN(
        n6343) );
  NAND2_X1 U8036 ( .A1(P2_REG2_REG_9__SCAN_IN), .A2(n6704), .ZN(n6341) );
  OAI21_X1 U8037 ( .B1(n6704), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6341), .ZN(
        n6342) );
  NOR2_X1 U8038 ( .A1(n6343), .A2(n6342), .ZN(n6355) );
  AOI211_X1 U8039 ( .C1(n6343), .C2(n6342), .A(n6355), .B(n9414), .ZN(n6354)
         );
  NAND2_X1 U8040 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n6720) );
  INV_X1 U8041 ( .A(n6720), .ZN(n6344) );
  AOI21_X1 U8042 ( .B1(n9898), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n6344), .ZN(
        n6352) );
  INV_X1 U8043 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10016) );
  MUX2_X1 U8044 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10016), .S(n6595), .Z(n6374)
         );
  NAND2_X1 U8045 ( .A1(n6345), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6347) );
  NAND2_X1 U8046 ( .A1(n6347), .A2(n6346), .ZN(n6375) );
  NAND2_X1 U8047 ( .A1(n6374), .A2(n6375), .ZN(n6373) );
  OAI21_X1 U8048 ( .B1(n6378), .B2(n10016), .A(n6373), .ZN(n6350) );
  INV_X1 U8049 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6348) );
  MUX2_X1 U8050 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6348), .S(n6704), .Z(n6349)
         );
  NAND2_X1 U8051 ( .A1(n6349), .A2(n6350), .ZN(n6360) );
  OAI211_X1 U8052 ( .C1(n6350), .C2(n6349), .A(n9892), .B(n6360), .ZN(n6351)
         );
  OAI211_X1 U8053 ( .C1(n8234), .C2(n6361), .A(n6352), .B(n6351), .ZN(n6353)
         );
  OR2_X1 U8054 ( .A1(n6354), .A2(n6353), .ZN(P2_U3254) );
  NAND2_X1 U8055 ( .A1(n6792), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6356) );
  OAI21_X1 U8056 ( .B1(n6792), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6356), .ZN(
        n6357) );
  AOI211_X1 U8057 ( .C1(n6358), .C2(n6357), .A(n6729), .B(n9414), .ZN(n6368)
         );
  NAND2_X1 U8058 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n6991) );
  INV_X1 U8059 ( .A(n6991), .ZN(n6359) );
  AOI21_X1 U8060 ( .B1(n9898), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n6359), .ZN(
        n6366) );
  OAI21_X1 U8061 ( .B1(n6361), .B2(n6348), .A(n6360), .ZN(n6364) );
  INV_X1 U8062 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6362) );
  MUX2_X1 U8063 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6362), .S(n6792), .Z(n6363)
         );
  NAND2_X1 U8064 ( .A1(n6363), .A2(n6364), .ZN(n6735) );
  OAI211_X1 U8065 ( .C1(n6364), .C2(n6363), .A(n9892), .B(n6735), .ZN(n6365)
         );
  OAI211_X1 U8066 ( .C1(n8234), .C2(n6736), .A(n6366), .B(n6365), .ZN(n6367)
         );
  OR2_X1 U8067 ( .A1(n6368), .A2(n6367), .ZN(P2_U3255) );
  AOI211_X1 U8068 ( .C1(n6371), .C2(n6370), .A(n6369), .B(n9414), .ZN(n6380)
         );
  NAND2_X1 U8069 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n6602) );
  INV_X1 U8070 ( .A(n6602), .ZN(n6372) );
  AOI21_X1 U8071 ( .B1(n9898), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6372), .ZN(
        n6377) );
  OAI211_X1 U8072 ( .C1(n6375), .C2(n6374), .A(n9892), .B(n6373), .ZN(n6376)
         );
  OAI211_X1 U8073 ( .C1(n8234), .C2(n6378), .A(n6377), .B(n6376), .ZN(n6379)
         );
  OR2_X1 U8074 ( .A1(n6380), .A2(n6379), .ZN(P2_U3253) );
  NOR2_X1 U8075 ( .A1(n8527), .A2(n8526), .ZN(n6392) );
  NAND2_X1 U8076 ( .A1(n6392), .A2(n8613), .ZN(n6383) );
  NAND2_X1 U8077 ( .A1(n8531), .A2(n8023), .ZN(n6384) );
  NAND4_X1 U8078 ( .A1(n7444), .A2(n6385), .A3(n8481), .A4(n6384), .ZN(n8533)
         );
  NAND2_X1 U8079 ( .A1(n8020), .A2(n8530), .ZN(n7848) );
  OR2_X1 U8080 ( .A1(n8023), .A2(n7848), .ZN(n6558) );
  NAND2_X1 U8081 ( .A1(n8533), .A2(n6558), .ZN(n6386) );
  INV_X1 U8082 ( .A(n9444), .ZN(n6531) );
  NAND2_X1 U8083 ( .A1(n6387), .A2(n6446), .ZN(n7860) );
  NAND2_X1 U8084 ( .A1(n6402), .A2(n9920), .ZN(n7862) );
  NAND2_X1 U8085 ( .A1(n7860), .A2(n7862), .ZN(n6438) );
  NAND2_X1 U8086 ( .A1(n6438), .A2(n6437), .ZN(n6436) );
  NAND2_X1 U8087 ( .A1(n6387), .A2(n9920), .ZN(n6388) );
  INV_X1 U8088 ( .A(n6550), .ZN(n8191) );
  INV_X1 U8089 ( .A(n9929), .ZN(n6390) );
  NAND2_X1 U8090 ( .A1(n8191), .A2(n6390), .ZN(n7864) );
  NAND2_X1 U8091 ( .A1(n6550), .A2(n9929), .ZN(n7863) );
  OAI21_X1 U8092 ( .B1(n4862), .B2(n6396), .A(n6525), .ZN(n9933) );
  AND2_X1 U8093 ( .A1(n9913), .A2(n8023), .ZN(n6389) );
  NOR2_X1 U8094 ( .A1(n8529), .A2(n8530), .ZN(n6391) );
  AND2_X1 U8095 ( .A1(n6392), .A2(n6391), .ZN(n9448) );
  NAND2_X1 U8096 ( .A1(n6444), .A2(n9929), .ZN(n6393) );
  NAND2_X1 U8097 ( .A1(n6393), .A2(n9456), .ZN(n6394) );
  NOR2_X1 U8098 ( .A1(n6554), .A2(n6394), .ZN(n9928) );
  AOI22_X1 U8099 ( .A1(n9448), .A2(n9928), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n9435), .ZN(n6395) );
  OAI21_X1 U8100 ( .B1(n9438), .B2(n6390), .A(n6395), .ZN(n6404) );
  NAND2_X1 U8101 ( .A1(n8027), .A2(n8530), .ZN(n8022) );
  NAND2_X1 U8102 ( .A1(n6398), .A2(n6397), .ZN(n6546) );
  INV_X1 U8103 ( .A(n6546), .ZN(n6399) );
  AOI21_X1 U8104 ( .B1(n6396), .B2(n6400), .A(n6399), .ZN(n6401) );
  OAI222_X1 U8105 ( .A1(n8455), .A2(n6402), .B1(n8457), .B2(n6611), .C1(n8512), 
        .C2(n6401), .ZN(n9927) );
  MUX2_X1 U8106 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9927), .S(n9441), .Z(n6403)
         );
  AOI211_X1 U8107 ( .C1(n6531), .C2(n9933), .A(n6404), .B(n6403), .ZN(n6405)
         );
  INV_X1 U8108 ( .A(n6405), .ZN(P2_U3294) );
  NOR2_X1 U8109 ( .A1(n6657), .A2(n9913), .ZN(n6411) );
  OR2_X1 U8110 ( .A1(n6790), .A2(n6406), .ZN(n6409) );
  OR2_X1 U8111 ( .A1(n4304), .A2(n6407), .ZN(n6408) );
  OAI211_X1 U8112 ( .C1(n6501), .C2(n6410), .A(n6409), .B(n6408), .ZN(n6477)
         );
  XNOR2_X1 U8113 ( .A(n6477), .B(n7390), .ZN(n6412) );
  NAND2_X1 U8114 ( .A1(n6411), .A2(n6412), .ZN(n6415) );
  INV_X1 U8115 ( .A(n6411), .ZN(n6414) );
  INV_X1 U8116 ( .A(n6412), .ZN(n6413) );
  NAND2_X1 U8117 ( .A1(n6414), .A2(n6413), .ZN(n6494) );
  AND2_X1 U8118 ( .A1(n6415), .A2(n6494), .ZN(n6423) );
  INV_X1 U8119 ( .A(n6418), .ZN(n6421) );
  INV_X1 U8120 ( .A(n6419), .ZN(n6420) );
  NAND2_X1 U8121 ( .A1(n6421), .A2(n6420), .ZN(n6422) );
  OAI21_X1 U8122 ( .B1(n6423), .B2(n4402), .A(n6495), .ZN(n6434) );
  INV_X1 U8123 ( .A(n6477), .ZN(n9956) );
  NAND2_X1 U8124 ( .A1(n8158), .A2(n6479), .ZN(n6432) );
  NAND2_X1 U8125 ( .A1(n7832), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6429) );
  NAND2_X1 U8126 ( .A1(n6424), .A2(n6509), .ZN(n6425) );
  AND2_X1 U8127 ( .A1(n6503), .A2(n6425), .ZN(n6662) );
  NAND2_X1 U8128 ( .A1(n6143), .A2(n6662), .ZN(n6428) );
  NAND2_X1 U8129 ( .A1(n7244), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6427) );
  NAND2_X1 U8130 ( .A1(n6802), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6426) );
  OR2_X1 U8131 ( .A1(n6634), .A2(n8457), .ZN(n6430) );
  OAI21_X1 U8132 ( .B1(n6467), .B2(n8455), .A(n6430), .ZN(n6465) );
  AOI22_X1 U8133 ( .A1(n9881), .A2(n6465), .B1(P2_REG3_REG_6__SCAN_IN), .B2(
        P2_U3152), .ZN(n6431) );
  OAI211_X1 U8134 ( .C1(n9956), .C2(n8161), .A(n6432), .B(n6431), .ZN(n6433)
         );
  AOI21_X1 U8135 ( .B1(n6434), .B2(n8150), .A(n6433), .ZN(n6435) );
  INV_X1 U8136 ( .A(n6435), .ZN(P2_U3241) );
  OAI21_X1 U8137 ( .B1(n6438), .B2(n6437), .A(n6436), .ZN(n9923) );
  NOR2_X1 U8138 ( .A1(n6550), .A2(n8457), .ZN(n6442) );
  INV_X1 U8139 ( .A(n7850), .ZN(n6440) );
  INV_X1 U8140 ( .A(n6438), .ZN(n7992) );
  NOR2_X1 U8141 ( .A1(n7992), .A2(n6535), .ZN(n6439) );
  AOI211_X1 U8142 ( .C1(n6440), .C2(n7860), .A(n8512), .B(n6439), .ZN(n6441)
         );
  AOI211_X1 U8143 ( .C1(n8605), .C2(n8192), .A(n6442), .B(n6441), .ZN(n9922)
         );
  MUX2_X1 U8144 ( .A(n6254), .B(n9922), .S(n9441), .Z(n6449) );
  NAND2_X1 U8145 ( .A1(n9920), .A2(n9914), .ZN(n6443) );
  AND3_X1 U8146 ( .A1(n6444), .A2(n9456), .A3(n6443), .ZN(n9919) );
  AOI22_X1 U8147 ( .A1(n9448), .A2(n9919), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9435), .ZN(n6445) );
  OAI21_X1 U8148 ( .B1(n9438), .B2(n6446), .A(n6445), .ZN(n6447) );
  INV_X1 U8149 ( .A(n6447), .ZN(n6448) );
  OAI211_X1 U8150 ( .C1(n9444), .C2(n9923), .A(n6449), .B(n6448), .ZN(P2_U3295) );
  AOI21_X1 U8151 ( .B1(n9550), .B2(n6451), .A(n6450), .ZN(n6453) );
  MUX2_X1 U8152 ( .A(n9544), .B(P1_REG1_REG_12__SCAN_IN), .S(n9030), .Z(n6452)
         );
  NOR2_X1 U8153 ( .A1(n6453), .A2(n6452), .ZN(n9040) );
  AOI21_X1 U8154 ( .B1(n6453), .B2(n6452), .A(n9040), .ZN(n6461) );
  NAND2_X1 U8155 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7262) );
  OAI21_X1 U8156 ( .B1(n9702), .B2(n9041), .A(n7262), .ZN(n6459) );
  OAI21_X1 U8157 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6455), .A(n6454), .ZN(
        n6457) );
  XNOR2_X1 U8158 ( .A(n9030), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n6456) );
  NOR2_X1 U8159 ( .A1(n6457), .A2(n6456), .ZN(n9029) );
  AOI211_X1 U8160 ( .C1(n6457), .C2(n6456), .A(n9665), .B(n9029), .ZN(n6458)
         );
  AOI211_X1 U8161 ( .C1(n9603), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n6459), .B(
        n6458), .ZN(n6460) );
  OAI21_X1 U8162 ( .B1(n6461), .B2(n9708), .A(n6460), .ZN(P1_U3253) );
  NAND2_X1 U8163 ( .A1(n6546), .A2(n7863), .ZN(n6462) );
  NAND2_X1 U8164 ( .A1(n6611), .A2(n9885), .ZN(n6608) );
  INV_X1 U8165 ( .A(n6611), .ZN(n8190) );
  INV_X1 U8166 ( .A(n7990), .ZN(n7856) );
  NAND2_X1 U8167 ( .A1(n6462), .A2(n7856), .ZN(n6545) );
  NAND2_X1 U8168 ( .A1(n6548), .A2(n6616), .ZN(n7854) );
  AND2_X1 U8169 ( .A1(n7854), .A2(n6608), .ZN(n7857) );
  INV_X1 U8170 ( .A(n6467), .ZN(n8188) );
  INV_X1 U8171 ( .A(n6548), .ZN(n8189) );
  NAND2_X1 U8172 ( .A1(n8189), .A2(n9942), .ZN(n6514) );
  NAND2_X1 U8173 ( .A1(n6467), .A2(n6476), .ZN(n7858) );
  NAND2_X1 U8174 ( .A1(n6657), .A2(n6477), .ZN(n7875) );
  INV_X1 U8175 ( .A(n6657), .ZN(n8187) );
  NAND2_X1 U8176 ( .A1(n8187), .A2(n9956), .ZN(n7873) );
  NAND2_X1 U8177 ( .A1(n7875), .A2(n7873), .ZN(n7996) );
  NAND3_X1 U8178 ( .A1(n6463), .A2(n7858), .A3(n7996), .ZN(n6464) );
  AOI21_X1 U8179 ( .B1(n6640), .B2(n6464), .A(n8512), .ZN(n6466) );
  NOR2_X1 U8180 ( .A1(n6466), .A2(n6465), .ZN(n9955) );
  NAND2_X1 U8181 ( .A1(n6550), .A2(n6390), .ZN(n6524) );
  NAND2_X1 U8182 ( .A1(n6611), .A2(n9936), .ZN(n6526) );
  NAND2_X1 U8183 ( .A1(n6548), .A2(n9942), .ZN(n6528) );
  NAND2_X1 U8184 ( .A1(n6467), .A2(n9950), .ZN(n6473) );
  INV_X1 U8185 ( .A(n6470), .ZN(n6471) );
  NAND2_X1 U8186 ( .A1(n7854), .A2(n6514), .ZN(n7991) );
  OR2_X1 U8187 ( .A1(n6471), .A2(n7991), .ZN(n6472) );
  INV_X1 U8188 ( .A(n6473), .ZN(n6474) );
  NAND2_X1 U8189 ( .A1(n7858), .A2(n7868), .ZN(n7995) );
  AND2_X1 U8190 ( .A1(n6632), .A2(n6631), .ZN(n6475) );
  XNOR2_X1 U8191 ( .A(n6475), .B(n7996), .ZN(n9958) );
  NAND2_X1 U8192 ( .A1(n9958), .A2(n6531), .ZN(n6484) );
  NOR2_X1 U8193 ( .A1(n9438), .A2(n9956), .ZN(n6482) );
  INV_X1 U8194 ( .A(n9448), .ZN(n6555) );
  OR2_X1 U8195 ( .A1(n6612), .A2(n6616), .ZN(n6613) );
  XNOR2_X1 U8196 ( .A(n6646), .B(n6477), .ZN(n6478) );
  NAND2_X1 U8197 ( .A1(n6478), .A2(n9456), .ZN(n9954) );
  INV_X1 U8198 ( .A(n6479), .ZN(n6480) );
  OAI22_X1 U8199 ( .A1(n6555), .A2(n9954), .B1(n6480), .B2(n8437), .ZN(n6481)
         );
  AOI211_X1 U8200 ( .C1(n4305), .C2(P2_REG2_REG_6__SCAN_IN), .A(n6482), .B(
        n6481), .ZN(n6483) );
  OAI211_X1 U8201 ( .C1(n9955), .C2(n4305), .A(n6484), .B(n6483), .ZN(P2_U3290) );
  INV_X1 U8202 ( .A(n9782), .ZN(n6492) );
  OAI211_X1 U8203 ( .C1(n6487), .C2(n6486), .A(n6485), .B(n8977), .ZN(n6491)
         );
  OAI22_X1 U8204 ( .A1(n4956), .A2(n8994), .B1(n8953), .B2(n9773), .ZN(n6488)
         );
  AOI211_X1 U8205 ( .C1(n9758), .C2(n8965), .A(n6489), .B(n6488), .ZN(n6490)
         );
  OAI211_X1 U8206 ( .C1(n6493), .C2(n6492), .A(n6491), .B(n6490), .ZN(P1_U3228) );
  OR2_X1 U8207 ( .A1(n6634), .A2(n9913), .ZN(n6590) );
  NAND2_X1 U8208 ( .A1(n7839), .A2(n6496), .ZN(n6499) );
  OR2_X1 U8209 ( .A1(n4304), .A2(n6497), .ZN(n6498) );
  OAI211_X1 U8210 ( .C1(n6501), .C2(n6500), .A(n6499), .B(n6498), .ZN(n6665)
         );
  XNOR2_X1 U8211 ( .A(n6665), .B(n7798), .ZN(n6591) );
  XNOR2_X1 U8212 ( .A(n6590), .B(n6591), .ZN(n6592) );
  XNOR2_X1 U8213 ( .A(n6593), .B(n6592), .ZN(n6513) );
  NAND2_X1 U8214 ( .A1(n7832), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6508) );
  INV_X1 U8215 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6502) );
  NAND2_X1 U8216 ( .A1(n6503), .A2(n6502), .ZN(n6504) );
  AND2_X1 U8217 ( .A1(n6713), .A2(n6504), .ZN(n6648) );
  NAND2_X1 U8218 ( .A1(n6143), .A2(n6648), .ZN(n6507) );
  NAND2_X1 U8219 ( .A1(n7244), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U8220 ( .A1(n6802), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6505) );
  OAI22_X1 U8221 ( .A1(n6719), .A2(n8145), .B1(n8156), .B2(n6657), .ZN(n6511)
         );
  INV_X1 U8222 ( .A(n6665), .ZN(n9960) );
  OAI22_X1 U8223 ( .A1(n8161), .A2(n9960), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6509), .ZN(n6510) );
  AOI211_X1 U8224 ( .C1(n6662), .C2(n8158), .A(n6511), .B(n6510), .ZN(n6512)
         );
  OAI21_X1 U8225 ( .B1(n6513), .B2(n9882), .A(n6512), .ZN(P2_U3215) );
  NAND2_X1 U8226 ( .A1(n6515), .A2(n6514), .ZN(n6516) );
  XNOR2_X1 U8227 ( .A(n6516), .B(n7995), .ZN(n6518) );
  AOI21_X1 U8228 ( .B1(n6518), .B2(n8608), .A(n6517), .ZN(n9949) );
  NOR2_X1 U8229 ( .A1(n4305), .A2(n8530), .ZN(n8519) );
  INV_X1 U8230 ( .A(n6646), .ZN(n6519) );
  OAI211_X1 U8231 ( .C1(n9950), .C2(n4529), .A(n6519), .B(n9456), .ZN(n9948)
         );
  INV_X1 U8232 ( .A(n9948), .ZN(n6523) );
  AOI22_X1 U8233 ( .A1(n4305), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n6520), .B2(
        n9435), .ZN(n6521) );
  OAI21_X1 U8234 ( .B1(n9950), .B2(n9438), .A(n6521), .ZN(n6522) );
  AOI21_X1 U8235 ( .B1(n8519), .B2(n6523), .A(n6522), .ZN(n6533) );
  NAND2_X1 U8236 ( .A1(n6525), .A2(n6524), .ZN(n6544) );
  NAND2_X1 U8237 ( .A1(n6544), .A2(n7990), .ZN(n6527) );
  NAND2_X1 U8238 ( .A1(n6527), .A2(n6526), .ZN(n6607) );
  NAND2_X1 U8239 ( .A1(n6607), .A2(n7991), .ZN(n6529) );
  NAND2_X1 U8240 ( .A1(n6529), .A2(n6528), .ZN(n6530) );
  XNOR2_X1 U8241 ( .A(n7995), .B(n6530), .ZN(n9952) );
  NAND2_X1 U8242 ( .A1(n9952), .A2(n6531), .ZN(n6532) );
  OAI211_X1 U8243 ( .C1(n9949), .C2(n4305), .A(n6533), .B(n6532), .ZN(P2_U3291) );
  NAND2_X1 U8244 ( .A1(n8192), .A2(n6534), .ZN(n7859) );
  NAND2_X1 U8245 ( .A1(n6535), .A2(n7859), .ZN(n9915) );
  INV_X1 U8246 ( .A(n9915), .ZN(n6540) );
  AOI22_X1 U8247 ( .A1(n9915), .A2(n8608), .B1(n8603), .B2(n6387), .ZN(n9917)
         );
  OAI21_X1 U8248 ( .B1(n6071), .B2(n8437), .A(n9917), .ZN(n6537) );
  NOR2_X1 U8249 ( .A1(n9441), .A2(n9896), .ZN(n6536) );
  AOI21_X1 U8250 ( .B1(n9441), .B2(n6537), .A(n6536), .ZN(n6539) );
  OAI21_X1 U8251 ( .B1(n8484), .B2(n8494), .A(n9914), .ZN(n6538) );
  OAI211_X1 U8252 ( .C1(n6540), .C2(n9444), .A(n6539), .B(n6538), .ZN(P2_U3296) );
  INV_X1 U8253 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n8700) );
  INV_X1 U8254 ( .A(n7362), .ZN(n6543) );
  INV_X1 U8255 ( .A(n9038), .ZN(n9701) );
  OAI222_X1 U8256 ( .A1(n9401), .A2(n8700), .B1(n9397), .B2(n6543), .C1(
        P1_U3084), .C2(n9701), .ZN(P1_U3335) );
  INV_X1 U8257 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U8258 ( .A1(n4396), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6542) );
  XNOR2_X1 U8259 ( .A(n6542), .B(n6541), .ZN(n8258) );
  OAI222_X1 U8260 ( .A1(n8827), .A2(n8704), .B1(n8835), .B2(n6543), .C1(
        P2_U3152), .C2(n8258), .ZN(P2_U3340) );
  XNOR2_X1 U8261 ( .A(n6544), .B(n7990), .ZN(n9938) );
  INV_X1 U8262 ( .A(n8533), .ZN(n6642) );
  NAND2_X1 U8263 ( .A1(n9938), .A2(n6642), .ZN(n6553) );
  NAND3_X1 U8264 ( .A1(n6546), .A2(n7863), .A3(n7990), .ZN(n6547) );
  NAND2_X1 U8265 ( .A1(n6545), .A2(n6547), .ZN(n6551) );
  OR2_X1 U8266 ( .A1(n6548), .A2(n8457), .ZN(n6549) );
  OAI21_X1 U8267 ( .B1(n6550), .B2(n8455), .A(n6549), .ZN(n9880) );
  AOI21_X1 U8268 ( .B1(n6551), .B2(n8608), .A(n9880), .ZN(n6552) );
  AND2_X1 U8269 ( .A1(n6553), .A2(n6552), .ZN(n9940) );
  OAI211_X1 U8270 ( .C1(n6554), .C2(n9936), .A(n9456), .B(n6612), .ZN(n9935)
         );
  OAI22_X1 U8271 ( .A1(n6555), .A2(n9935), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8437), .ZN(n6557) );
  NOR2_X1 U8272 ( .A1(n9441), .A2(n6257), .ZN(n6556) );
  AOI211_X1 U8273 ( .C1(n8484), .C2(n9885), .A(n6557), .B(n6556), .ZN(n6561)
         );
  INV_X1 U8274 ( .A(n8487), .ZN(n6559) );
  NAND2_X1 U8275 ( .A1(n6559), .A2(n9938), .ZN(n6560) );
  OAI211_X1 U8276 ( .C1(n4305), .C2(n9940), .A(n6561), .B(n6560), .ZN(P2_U3293) );
  INV_X1 U8277 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6568) );
  OAI21_X1 U8278 ( .B1(n6563), .B2(n9283), .A(n6562), .ZN(n6564) );
  NAND2_X1 U8279 ( .A1(n6564), .A2(n9779), .ZN(n6567) );
  OAI21_X1 U8280 ( .B1(n9720), .B2(n9494), .A(n6565), .ZN(n6566) );
  OAI211_X1 U8281 ( .C1(n6568), .C2(n9779), .A(n6567), .B(n6566), .ZN(P1_U3291) );
  XNOR2_X1 U8282 ( .A(n6569), .B(n7726), .ZN(n9793) );
  AND2_X1 U8283 ( .A1(n6571), .A2(n9745), .ZN(n6570) );
  INV_X1 U8284 ( .A(n9764), .ZN(n6842) );
  OR2_X1 U8285 ( .A1(n6572), .A2(n6571), .ZN(n6575) );
  OR2_X1 U8286 ( .A1(n6573), .A2(n7776), .ZN(n6574) );
  AND2_X1 U8287 ( .A1(n6575), .A2(n6574), .ZN(n9730) );
  AOI22_X1 U8288 ( .A1(n4932), .A2(n9742), .B1(n9489), .B2(n5553), .ZN(n6580)
         );
  OAI21_X1 U8289 ( .B1(n6577), .B2(n7726), .A(n6576), .ZN(n6578) );
  NAND2_X1 U8290 ( .A1(n6578), .A2(n9770), .ZN(n6579) );
  OAI211_X1 U8291 ( .C1(n9793), .C2(n9730), .A(n6580), .B(n6579), .ZN(n9796)
         );
  INV_X1 U8292 ( .A(n6671), .ZN(n6581) );
  OAI211_X1 U8293 ( .C1(n9795), .C2(n6582), .A(n6581), .B(n9828), .ZN(n9794)
         );
  INV_X1 U8294 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6583) );
  OAI22_X1 U8295 ( .A1(n9794), .A2(n9745), .B1(n9283), .B2(n6583), .ZN(n6584)
         );
  OAI21_X1 U8296 ( .B1(n9796), .B2(n6584), .A(n9779), .ZN(n6586) );
  AOI22_X1 U8297 ( .A1(n9494), .A2(n7524), .B1(n9755), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6585) );
  OAI211_X1 U8298 ( .C1(n9793), .C2(n6842), .A(n6586), .B(n6585), .ZN(P1_U3290) );
  INV_X1 U8299 ( .A(n7368), .ZN(n6588) );
  OAI222_X1 U8300 ( .A1(n8827), .A2(n6587), .B1(n8835), .B2(n6588), .C1(
        P2_U3152), .C2(n8481), .ZN(P2_U3339) );
  OAI222_X1 U8301 ( .A1(n9401), .A2(n6589), .B1(n9397), .B2(n6588), .C1(
        P1_U3084), .C2(n9136), .ZN(P1_U3334) );
  OR2_X1 U8302 ( .A1(n6719), .A2(n9913), .ZN(n6698) );
  AOI22_X1 U8303 ( .A1(n7370), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7369), .B2(
        n6595), .ZN(n6596) );
  XNOR2_X1 U8304 ( .A(n6747), .B(n7390), .ZN(n6699) );
  XNOR2_X1 U8305 ( .A(n6698), .B(n6699), .ZN(n6696) );
  XNOR2_X1 U8306 ( .A(n6697), .B(n6696), .ZN(n6606) );
  NAND2_X1 U8307 ( .A1(n7832), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6601) );
  XNOR2_X1 U8308 ( .A(n6713), .B(P2_REG3_REG_9__SCAN_IN), .ZN(n6761) );
  NAND2_X1 U8309 ( .A1(n6143), .A2(n6761), .ZN(n6600) );
  NAND2_X1 U8310 ( .A1(n7244), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U8311 ( .A1(n6802), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6598) );
  NAND4_X1 U8312 ( .A1(n6601), .A2(n6600), .A3(n6599), .A4(n6598), .ZN(n8184)
         );
  INV_X1 U8313 ( .A(n8184), .ZN(n6807) );
  OAI22_X1 U8314 ( .A1(n6634), .A2(n8156), .B1(n8145), .B2(n6807), .ZN(n6604)
         );
  INV_X1 U8315 ( .A(n6747), .ZN(n9966) );
  OAI21_X1 U8316 ( .B1(n8161), .B2(n9966), .A(n6602), .ZN(n6603) );
  AOI211_X1 U8317 ( .C1(n6648), .C2(n8158), .A(n6604), .B(n6603), .ZN(n6605)
         );
  OAI21_X1 U8318 ( .B1(n6606), .B2(n9882), .A(n6605), .ZN(P2_U3223) );
  XNOR2_X1 U8319 ( .A(n6607), .B(n7991), .ZN(n9946) );
  INV_X1 U8320 ( .A(n9946), .ZN(n6621) );
  NAND2_X1 U8321 ( .A1(n6545), .A2(n6608), .ZN(n6609) );
  XNOR2_X1 U8322 ( .A(n6609), .B(n7991), .ZN(n6610) );
  OAI222_X1 U8323 ( .A1(n8457), .A2(n6467), .B1(n8455), .B2(n6611), .C1(n6610), 
        .C2(n8512), .ZN(n9944) );
  INV_X1 U8324 ( .A(n6612), .ZN(n6614) );
  OAI21_X1 U8325 ( .B1(n6614), .B2(n9942), .A(n6613), .ZN(n9943) );
  AOI22_X1 U8326 ( .A1(n4305), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n6615), .B2(
        n9435), .ZN(n6618) );
  NAND2_X1 U8327 ( .A1(n8484), .A2(n6616), .ZN(n6617) );
  OAI211_X1 U8328 ( .C1(n8443), .C2(n9943), .A(n6618), .B(n6617), .ZN(n6619)
         );
  AOI21_X1 U8329 ( .B1(n9944), .B2(n9441), .A(n6619), .ZN(n6620) );
  OAI21_X1 U8330 ( .B1(n6621), .B2(n9444), .A(n6620), .ZN(P2_U3292) );
  XNOR2_X1 U8331 ( .A(n6623), .B(n6622), .ZN(n6624) );
  XNOR2_X1 U8332 ( .A(n6625), .B(n6624), .ZN(n6630) );
  OAI22_X1 U8333 ( .A1(n6919), .A2(n8994), .B1(n8953), .B2(n7044), .ZN(n6626)
         );
  AOI211_X1 U8334 ( .C1(n6922), .C2(n8965), .A(n6627), .B(n6626), .ZN(n6629)
         );
  NAND2_X1 U8335 ( .A1(n8997), .A2(n6921), .ZN(n6628) );
  OAI211_X1 U8336 ( .C1(n6630), .C2(n8988), .A(n6629), .B(n6628), .ZN(P1_U3211) );
  NAND2_X1 U8337 ( .A1(n6657), .A2(n9956), .ZN(n6633) );
  NAND2_X1 U8338 ( .A1(n6634), .A2(n6665), .ZN(n7880) );
  INV_X1 U8339 ( .A(n6634), .ZN(n8186) );
  NAND2_X1 U8340 ( .A1(n8186), .A2(n9960), .ZN(n7881) );
  NAND2_X1 U8341 ( .A1(n7880), .A2(n7881), .ZN(n7997) );
  NAND2_X1 U8342 ( .A1(n6634), .A2(n9960), .ZN(n6635) );
  NAND2_X1 U8343 ( .A1(n6636), .A2(n6635), .ZN(n6638) );
  NAND2_X1 U8344 ( .A1(n6719), .A2(n6747), .ZN(n7884) );
  NAND2_X1 U8345 ( .A1(n8185), .A2(n9966), .ZN(n7885) );
  NAND2_X1 U8346 ( .A1(n6638), .A2(n8001), .ZN(n6639) );
  INV_X1 U8347 ( .A(n9970), .ZN(n6653) );
  NAND3_X1 U8348 ( .A1(n6640), .A2(n7875), .A3(n7880), .ZN(n6641) );
  NAND2_X1 U8349 ( .A1(n6641), .A2(n7881), .ZN(n6860) );
  AOI21_X1 U8350 ( .B1(n6637), .B2(n6752), .A(n4389), .ZN(n6645) );
  NAND2_X1 U8351 ( .A1(n9970), .A2(n6642), .ZN(n6644) );
  AOI22_X1 U8352 ( .A1(n8186), .A2(n8605), .B1(n8603), .B2(n8184), .ZN(n6643)
         );
  OAI211_X1 U8353 ( .C1(n8512), .C2(n6645), .A(n6644), .B(n6643), .ZN(n9968)
         );
  NAND2_X1 U8354 ( .A1(n9968), .A2(n9441), .ZN(n6652) );
  INV_X1 U8355 ( .A(n6757), .ZN(n6759) );
  NAND2_X1 U8356 ( .A1(n4399), .A2(n6747), .ZN(n6647) );
  NAND2_X1 U8357 ( .A1(n6759), .A2(n6647), .ZN(n9967) );
  AOI22_X1 U8358 ( .A1(n4305), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n6648), .B2(
        n9435), .ZN(n6649) );
  OAI21_X1 U8359 ( .B1(n8443), .B2(n9967), .A(n6649), .ZN(n6650) );
  AOI21_X1 U8360 ( .B1(n8484), .B2(n6747), .A(n6650), .ZN(n6651) );
  OAI211_X1 U8361 ( .C1(n6653), .C2(n8487), .A(n6652), .B(n6651), .ZN(P2_U3288) );
  XNOR2_X1 U8362 ( .A(n6654), .B(n7997), .ZN(n9964) );
  INV_X1 U8363 ( .A(n9964), .ZN(n6668) );
  NAND2_X1 U8364 ( .A1(n6640), .A2(n7875), .ZN(n6655) );
  XNOR2_X1 U8365 ( .A(n6655), .B(n7997), .ZN(n6656) );
  OAI222_X1 U8366 ( .A1(n8455), .A2(n6657), .B1(n8457), .B2(n6719), .C1(n6656), 
        .C2(n8512), .ZN(n9962) );
  INV_X1 U8367 ( .A(n9962), .ZN(n6658) );
  MUX2_X1 U8368 ( .A(n6659), .B(n6658), .S(n9441), .Z(n6667) );
  OR2_X1 U8369 ( .A1(n6660), .A2(n9960), .ZN(n6661) );
  NAND2_X1 U8370 ( .A1(n4399), .A2(n6661), .ZN(n9961) );
  INV_X1 U8371 ( .A(n6662), .ZN(n6663) );
  OAI22_X1 U8372 ( .A1(n8443), .A2(n9961), .B1(n6663), .B2(n8437), .ZN(n6664)
         );
  AOI21_X1 U8373 ( .B1(n8484), .B2(n6665), .A(n6664), .ZN(n6666) );
  OAI211_X1 U8374 ( .C1(n6668), .C2(n9444), .A(n6667), .B(n6666), .ZN(P2_U3289) );
  INV_X1 U8375 ( .A(n7723), .ZN(n6670) );
  XNOR2_X1 U8376 ( .A(n6669), .B(n6670), .ZN(n9803) );
  INV_X1 U8377 ( .A(n9720), .ZN(n9762) );
  NOR2_X1 U8378 ( .A1(n6671), .A2(n4931), .ZN(n6672) );
  OR2_X1 U8379 ( .A1(n6688), .A2(n6672), .ZN(n9800) );
  AOI22_X1 U8380 ( .A1(n9494), .A2(n8964), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9783), .ZN(n6673) );
  OAI21_X1 U8381 ( .B1(n9762), .B2(n9800), .A(n6673), .ZN(n6679) );
  INV_X1 U8382 ( .A(n9730), .ZN(n9776) );
  INV_X1 U8383 ( .A(n9489), .ZN(n9774) );
  OAI22_X1 U8384 ( .A1(n7525), .A2(n9774), .B1(n4956), .B2(n9772), .ZN(n6674)
         );
  AOI21_X1 U8385 ( .B1(n9803), .B2(n9776), .A(n6674), .ZN(n6677) );
  XNOR2_X1 U8386 ( .A(n7530), .B(n7723), .ZN(n6675) );
  NAND2_X1 U8387 ( .A1(n6675), .A2(n9770), .ZN(n6676) );
  NAND2_X1 U8388 ( .A1(n6677), .A2(n6676), .ZN(n9801) );
  MUX2_X1 U8389 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9801), .S(n9779), .Z(n6678)
         );
  AOI211_X1 U8390 ( .C1(n9764), .C2(n9803), .A(n6679), .B(n6678), .ZN(n6680)
         );
  INV_X1 U8391 ( .A(n6680), .ZN(P1_U3289) );
  XNOR2_X1 U8392 ( .A(n5513), .B(n6681), .ZN(n9808) );
  OAI22_X1 U8393 ( .A1(n4934), .A2(n9774), .B1(n9748), .B2(n9772), .ZN(n6682)
         );
  AOI21_X1 U8394 ( .B1(n9808), .B2(n9776), .A(n6682), .ZN(n6687) );
  XNOR2_X1 U8395 ( .A(n6683), .B(n6684), .ZN(n6685) );
  NAND2_X1 U8396 ( .A1(n6685), .A2(n9770), .ZN(n6686) );
  AND2_X1 U8397 ( .A1(n6687), .A2(n6686), .ZN(n9810) );
  OR2_X1 U8398 ( .A1(n6688), .A2(n9805), .ZN(n6689) );
  NAND2_X1 U8399 ( .A1(n9759), .A2(n6689), .ZN(n9806) );
  OAI22_X1 U8400 ( .A1(n9779), .A2(n6690), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9283), .ZN(n6691) );
  AOI21_X1 U8401 ( .B1(n9494), .B2(n6692), .A(n6691), .ZN(n6693) );
  OAI21_X1 U8402 ( .B1(n9762), .B2(n9806), .A(n6693), .ZN(n6694) );
  AOI21_X1 U8403 ( .B1(n9808), .B2(n9764), .A(n6694), .ZN(n6695) );
  OAI21_X1 U8404 ( .B1(n9810), .B2(n9755), .A(n6695), .ZN(P1_U3288) );
  INV_X1 U8405 ( .A(n6698), .ZN(n6700) );
  NAND2_X1 U8406 ( .A1(n6700), .A2(n6699), .ZN(n6701) );
  AOI22_X1 U8407 ( .A1(n7370), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7369), .B2(
        n6704), .ZN(n6705) );
  XNOR2_X1 U8408 ( .A(n9973), .B(n7798), .ZN(n6709) );
  INV_X1 U8409 ( .A(n6709), .ZN(n6707) );
  AND2_X1 U8410 ( .A1(n8184), .A2(n7444), .ZN(n6708) );
  INV_X1 U8411 ( .A(n6708), .ZN(n6706) );
  NAND2_X1 U8412 ( .A1(n6707), .A2(n6706), .ZN(n6967) );
  AND2_X1 U8413 ( .A1(n6709), .A2(n6708), .ZN(n6965) );
  NOR2_X1 U8414 ( .A1(n4660), .A2(n6965), .ZN(n6710) );
  XNOR2_X1 U8415 ( .A(n6966), .B(n6710), .ZN(n6724) );
  NAND2_X1 U8416 ( .A1(n7832), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6718) );
  INV_X1 U8417 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6712) );
  INV_X1 U8418 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6711) );
  OAI21_X1 U8419 ( .B1(n6713), .B2(n6712), .A(n6711), .ZN(n6714) );
  AND2_X1 U8420 ( .A1(n6714), .A2(n6800), .ZN(n6811) );
  NAND2_X1 U8421 ( .A1(n6143), .A2(n6811), .ZN(n6717) );
  NAND2_X1 U8422 ( .A1(n7244), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6716) );
  NAND2_X1 U8423 ( .A1(n6802), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6715) );
  OAI22_X1 U8424 ( .A1(n6719), .A2(n8156), .B1(n8145), .B2(n6979), .ZN(n6722)
         );
  OAI21_X1 U8425 ( .B1(n8161), .B2(n9973), .A(n6720), .ZN(n6721) );
  AOI211_X1 U8426 ( .C1(n6761), .C2(n8158), .A(n6722), .B(n6721), .ZN(n6723)
         );
  OAI21_X1 U8427 ( .B1(n6724), .B2(n9882), .A(n6723), .ZN(P2_U3233) );
  INV_X1 U8428 ( .A(n7386), .ZN(n6746) );
  OAI222_X1 U8429 ( .A1(n9397), .A2(n6746), .B1(n6726), .B2(P1_U3084), .C1(
        n6725), .C2(n9401), .ZN(P1_U3333) );
  INV_X1 U8430 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6727) );
  MUX2_X1 U8431 ( .A(n6727), .B(P2_REG2_REG_11__SCAN_IN), .S(n8199), .Z(n6728)
         );
  INV_X1 U8432 ( .A(n6728), .ZN(n8195) );
  NAND2_X1 U8433 ( .A1(n6941), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6730) );
  OAI21_X1 U8434 ( .B1(n6941), .B2(P2_REG2_REG_12__SCAN_IN), .A(n6730), .ZN(
        n6731) );
  AOI211_X1 U8435 ( .C1(n6732), .C2(n6731), .A(n6777), .B(n9414), .ZN(n6745)
         );
  INV_X1 U8436 ( .A(n9892), .ZN(n9893) );
  INV_X1 U8437 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6733) );
  MUX2_X1 U8438 ( .A(n6733), .B(P2_REG1_REG_12__SCAN_IN), .S(n6941), .Z(n6739)
         );
  NAND2_X1 U8439 ( .A1(n8199), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6737) );
  INV_X1 U8440 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6734) );
  MUX2_X1 U8441 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n6734), .S(n8199), .Z(n8201)
         );
  OAI21_X1 U8442 ( .B1(n6736), .B2(n6362), .A(n6735), .ZN(n8202) );
  NAND2_X1 U8443 ( .A1(n8201), .A2(n8202), .ZN(n8200) );
  NAND2_X1 U8444 ( .A1(n6737), .A2(n8200), .ZN(n6738) );
  NOR2_X1 U8445 ( .A1(n6738), .A2(n6739), .ZN(n6778) );
  AOI21_X1 U8446 ( .B1(n6739), .B2(n6738), .A(n6778), .ZN(n6743) );
  NAND2_X1 U8447 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7011) );
  INV_X1 U8448 ( .A(n7011), .ZN(n6740) );
  AOI21_X1 U8449 ( .B1(n9898), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n6740), .ZN(
        n6742) );
  NAND2_X1 U8450 ( .A1(n9895), .A2(n6941), .ZN(n6741) );
  OAI211_X1 U8451 ( .C1(n9893), .C2(n6743), .A(n6742), .B(n6741), .ZN(n6744)
         );
  OR2_X1 U8452 ( .A1(n6745), .A2(n6744), .ZN(P2_U3257) );
  OAI222_X1 U8453 ( .A1(n8827), .A2(n7387), .B1(n8835), .B2(n6746), .C1(n6109), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  NAND2_X1 U8454 ( .A1(n9973), .A2(n8184), .ZN(n7893) );
  NAND2_X1 U8455 ( .A1(n8185), .A2(n6747), .ZN(n6748) );
  AOI21_X1 U8456 ( .B1(n7999), .B2(n6750), .A(n4392), .ZN(n9972) );
  INV_X1 U8457 ( .A(n6979), .ZN(n8183) );
  AOI22_X1 U8458 ( .A1(n8605), .A2(n8185), .B1(n8183), .B2(n8603), .ZN(n6756)
         );
  INV_X1 U8459 ( .A(n7884), .ZN(n6751) );
  NOR3_X1 U8460 ( .A1(n4389), .A2(n6751), .A3(n7999), .ZN(n6754) );
  OR2_X1 U8461 ( .A1(n6637), .A2(n6753), .ZN(n6858) );
  OR2_X1 U8462 ( .A1(n6752), .A2(n6858), .ZN(n6798) );
  OR2_X1 U8463 ( .A1(n6753), .A2(n7884), .ZN(n6797) );
  OAI21_X1 U8464 ( .B1(n6754), .B2(n4395), .A(n8608), .ZN(n6755) );
  OAI211_X1 U8465 ( .C1(n9972), .C2(n8533), .A(n6756), .B(n6755), .ZN(n9975)
         );
  NAND2_X1 U8466 ( .A1(n9975), .A2(n9441), .ZN(n6766) );
  NAND2_X1 U8467 ( .A1(n6759), .A2(n6758), .ZN(n6760) );
  NAND2_X1 U8468 ( .A1(n6813), .A2(n6760), .ZN(n9974) );
  INV_X1 U8469 ( .A(n9974), .ZN(n6764) );
  AOI22_X1 U8470 ( .A1(n4305), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n6761), .B2(
        n9435), .ZN(n6762) );
  OAI21_X1 U8471 ( .B1(n9973), .B2(n9438), .A(n6762), .ZN(n6763) );
  AOI21_X1 U8472 ( .B1(n6764), .B2(n8494), .A(n6763), .ZN(n6765) );
  OAI211_X1 U8473 ( .C1(n9972), .C2(n8487), .A(n6766), .B(n6765), .ZN(P2_U3287) );
  XNOR2_X1 U8474 ( .A(n6767), .B(n6768), .ZN(n6769) );
  NAND2_X1 U8475 ( .A1(n6769), .A2(n6770), .ZN(n6901) );
  OAI21_X1 U8476 ( .B1(n6770), .B2(n6769), .A(n6901), .ZN(n6771) );
  NAND2_X1 U8477 ( .A1(n6771), .A2(n8977), .ZN(n6776) );
  AND2_X1 U8478 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9594) );
  INV_X1 U8479 ( .A(n9594), .ZN(n6772) );
  OAI21_X1 U8480 ( .B1(n9000), .B2(n9821), .A(n6772), .ZN(n6774) );
  OAI22_X1 U8481 ( .A1(n6919), .A2(n8953), .B1(n8994), .B2(n9748), .ZN(n6773)
         );
  AOI211_X1 U8482 ( .C1(n9741), .C2(n8997), .A(n6774), .B(n6773), .ZN(n6775)
         );
  NAND2_X1 U8483 ( .A1(n6776), .A2(n6775), .ZN(P1_U3225) );
  XNOR2_X1 U8484 ( .A(n7059), .B(P2_REG2_REG_13__SCAN_IN), .ZN(n7020) );
  XNOR2_X1 U8485 ( .A(n7020), .B(n7019), .ZN(n6788) );
  AOI21_X1 U8486 ( .B1(n6779), .B2(n6733), .A(n6778), .ZN(n6783) );
  INV_X1 U8487 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9477) );
  MUX2_X1 U8488 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9477), .S(n7059), .Z(n6781)
         );
  INV_X1 U8489 ( .A(n6781), .ZN(n6782) );
  INV_X1 U8490 ( .A(n6783), .ZN(n6780) );
  AND2_X1 U8491 ( .A1(n6781), .A2(n6780), .ZN(n7024) );
  AOI21_X1 U8492 ( .B1(n6783), .B2(n6782), .A(n7024), .ZN(n6785) );
  NAND2_X1 U8493 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7069) );
  NAND2_X1 U8494 ( .A1(n9898), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6784) );
  OAI211_X1 U8495 ( .C1(n9893), .C2(n6785), .A(n7069), .B(n6784), .ZN(n6786)
         );
  AOI21_X1 U8496 ( .B1(n7059), .B2(n9895), .A(n6786), .ZN(n6787) );
  OAI21_X1 U8497 ( .B1(n6788), .B2(n9414), .A(n6787), .ZN(P2_U3258) );
  INV_X1 U8498 ( .A(n7400), .ZN(n6819) );
  OAI222_X1 U8499 ( .A1(n9397), .A2(n6819), .B1(n7776), .B2(P1_U3084), .C1(
        n6789), .C2(n9401), .ZN(P1_U3332) );
  AOI22_X1 U8500 ( .A1(n7370), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7369), .B2(
        n6792), .ZN(n6793) );
  OR2_X1 U8501 ( .A1(n6994), .A2(n6979), .ZN(n7892) );
  NAND2_X1 U8502 ( .A1(n6994), .A2(n6979), .ZN(n7895) );
  NAND2_X1 U8503 ( .A1(n6795), .A2(n8000), .ZN(n6796) );
  NAND2_X1 U8504 ( .A1(n6844), .A2(n6796), .ZN(n9979) );
  NAND2_X1 U8505 ( .A1(n6798), .A2(n6856), .ZN(n6799) );
  XNOR2_X1 U8506 ( .A(n6799), .B(n8000), .ZN(n6809) );
  NAND2_X1 U8507 ( .A1(n7832), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6806) );
  NAND2_X1 U8508 ( .A1(n6800), .A2(n8197), .ZN(n6801) );
  AND2_X1 U8509 ( .A1(n6850), .A2(n6801), .ZN(n6982) );
  NAND2_X1 U8510 ( .A1(n6143), .A2(n6982), .ZN(n6805) );
  NAND2_X1 U8511 ( .A1(n7244), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U8512 ( .A1(n6802), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6803) );
  OAI22_X1 U8513 ( .A1(n6807), .A2(n8455), .B1(n6993), .B2(n8457), .ZN(n6808)
         );
  AOI21_X1 U8514 ( .B1(n6809), .B2(n8608), .A(n6808), .ZN(n6810) );
  OAI21_X1 U8515 ( .B1(n9979), .B2(n8533), .A(n6810), .ZN(n9982) );
  NAND2_X1 U8516 ( .A1(n9982), .A2(n9441), .ZN(n6818) );
  INV_X1 U8517 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6812) );
  INV_X1 U8518 ( .A(n6811), .ZN(n6995) );
  OAI22_X1 U8519 ( .A1(n9441), .A2(n6812), .B1(n6995), .B2(n8437), .ZN(n6816)
         );
  AND2_X1 U8520 ( .A1(n6813), .A2(n6994), .ZN(n6814) );
  NOR2_X1 U8521 ( .A1(n6813), .A2(n6994), .ZN(n6862) );
  OR2_X1 U8522 ( .A1(n6814), .A2(n6862), .ZN(n9981) );
  NOR2_X1 U8523 ( .A1(n9981), .A2(n8443), .ZN(n6815) );
  AOI211_X1 U8524 ( .C1(n8484), .C2(n6994), .A(n6816), .B(n6815), .ZN(n6817)
         );
  OAI211_X1 U8525 ( .C1(n9979), .C2(n8487), .A(n6818), .B(n6817), .ZN(P2_U3286) );
  OAI222_X1 U8526 ( .A1(n8827), .A2(n7401), .B1(n8835), .B2(n6819), .C1(n7836), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  XOR2_X1 U8527 ( .A(n6822), .B(n6821), .Z(n6823) );
  XNOR2_X1 U8528 ( .A(n6820), .B(n6823), .ZN(n6829) );
  NOR2_X1 U8529 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6824), .ZN(n9621) );
  OAI22_X1 U8530 ( .A1(n9722), .A2(n8994), .B1(n8953), .B2(n9721), .ZN(n6825)
         );
  AOI211_X1 U8531 ( .C1(n6826), .C2(n8965), .A(n9621), .B(n6825), .ZN(n6828)
         );
  NAND2_X1 U8532 ( .A1(n8997), .A2(n9732), .ZN(n6827) );
  OAI211_X1 U8533 ( .C1(n6829), .C2(n8988), .A(n6828), .B(n6827), .ZN(P1_U3219) );
  INV_X1 U8534 ( .A(n6830), .ZN(n6831) );
  AOI21_X1 U8535 ( .B1(n7595), .B2(n6832), .A(n6831), .ZN(n9833) );
  NAND2_X1 U8536 ( .A1(n9769), .A2(n9766), .ZN(n9746) );
  INV_X1 U8537 ( .A(n7588), .ZN(n7599) );
  AOI21_X1 U8538 ( .B1(n9746), .B2(n9747), .A(n7599), .ZN(n6833) );
  XOR2_X1 U8539 ( .A(n7595), .B(n6833), .Z(n6836) );
  AOI22_X1 U8540 ( .A1(n9742), .A2(n9008), .B1(n9009), .B2(n9489), .ZN(n6834)
         );
  OAI21_X1 U8541 ( .B1(n9833), .B2(n9730), .A(n6834), .ZN(n6835) );
  AOI21_X1 U8542 ( .B1(n6836), .B2(n9770), .A(n6835), .ZN(n9831) );
  MUX2_X1 U8543 ( .A(n6837), .B(n9831), .S(n9779), .Z(n6841) );
  AOI21_X1 U8544 ( .B1(n9826), .B2(n4400), .A(n6920), .ZN(n9829) );
  INV_X1 U8545 ( .A(n6912), .ZN(n6838) );
  OAI22_X1 U8546 ( .A1(n9765), .A2(n6909), .B1(n6838), .B2(n9283), .ZN(n6839)
         );
  AOI21_X1 U8547 ( .B1(n9829), .B2(n9720), .A(n6839), .ZN(n6840) );
  OAI211_X1 U8548 ( .C1(n9833), .C2(n6842), .A(n6841), .B(n6840), .ZN(P1_U3285) );
  NAND2_X1 U8549 ( .A1(n6994), .A2(n8183), .ZN(n6843) );
  NAND2_X1 U8550 ( .A1(n6845), .A2(n7839), .ZN(n6847) );
  AOI22_X1 U8551 ( .A1(n7370), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7369), .B2(
        n8199), .ZN(n6846) );
  NAND2_X1 U8552 ( .A1(n6847), .A2(n6846), .ZN(n6973) );
  OR2_X1 U8553 ( .A1(n6973), .A2(n6993), .ZN(n7899) );
  NAND2_X1 U8554 ( .A1(n6973), .A2(n6993), .ZN(n7898) );
  NAND2_X1 U8555 ( .A1(n7899), .A2(n7898), .ZN(n8004) );
  OAI21_X1 U8556 ( .B1(n6848), .B2(n8004), .A(n6946), .ZN(n9987) );
  NAND2_X1 U8557 ( .A1(n6850), .A2(n6849), .ZN(n6851) );
  AND2_X1 U8558 ( .A1(n6949), .A2(n6851), .ZN(n7014) );
  NAND2_X1 U8559 ( .A1(n6143), .A2(n7014), .ZN(n6855) );
  NAND2_X1 U8560 ( .A1(n7832), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6854) );
  NAND2_X1 U8561 ( .A1(n7244), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6853) );
  NAND2_X1 U8562 ( .A1(n6802), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6852) );
  INV_X1 U8563 ( .A(n7892), .ZN(n6857) );
  OR2_X1 U8564 ( .A1(n6858), .A2(n6857), .ZN(n6859) );
  XNOR2_X1 U8565 ( .A(n6956), .B(n8004), .ZN(n6861) );
  OAI222_X1 U8566 ( .A1(n8457), .A2(n7112), .B1(n8455), .B2(n6979), .C1(n6861), 
        .C2(n8512), .ZN(n9990) );
  INV_X1 U8567 ( .A(n6973), .ZN(n9988) );
  NAND2_X1 U8568 ( .A1(n6862), .A2(n9988), .ZN(n6958) );
  OAI21_X1 U8569 ( .B1(n6862), .B2(n9988), .A(n6958), .ZN(n9989) );
  AOI22_X1 U8570 ( .A1(n4305), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n6982), .B2(
        n9435), .ZN(n6864) );
  NAND2_X1 U8571 ( .A1(n8484), .A2(n6973), .ZN(n6863) );
  OAI211_X1 U8572 ( .C1(n9989), .C2(n8443), .A(n6864), .B(n6863), .ZN(n6865)
         );
  AOI21_X1 U8573 ( .B1(n9990), .B2(n9441), .A(n6865), .ZN(n6866) );
  OAI21_X1 U8574 ( .B1(n9444), .B2(n9987), .A(n6866), .ZN(P2_U3285) );
  INV_X1 U8575 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10062) );
  NOR2_X1 U8576 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(P2_ADDR_REG_17__SCAN_IN), 
        .ZN(n6867) );
  AOI21_X1 U8577 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n6867), .ZN(n10031) );
  NOR2_X1 U8578 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .ZN(n6868) );
  AOI21_X1 U8579 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n6868), .ZN(n10034) );
  NOR2_X1 U8580 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n6869) );
  AOI21_X1 U8581 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n6869), .ZN(n10037) );
  NOR2_X1 U8582 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n6870) );
  AOI21_X1 U8583 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n6870), .ZN(n10040) );
  NOR2_X1 U8584 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .ZN(n6871) );
  AOI21_X1 U8585 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n6871), .ZN(n10043) );
  NOR2_X1 U8586 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n6880) );
  XOR2_X1 U8587 ( .A(n6872), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10072) );
  NAND2_X1 U8588 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n6878) );
  INV_X1 U8589 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6873) );
  AOI22_X1 U8590 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .B1(n6873), .B2(n8626), .ZN(n10070) );
  NAND2_X1 U8591 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n6876) );
  INV_X1 U8592 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6874) );
  XNOR2_X1 U8593 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n6874), .ZN(n10066) );
  AOI21_X1 U8594 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10024) );
  INV_X1 U8595 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10028) );
  NAND3_X1 U8596 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10026) );
  OAI21_X1 U8597 ( .B1(n10024), .B2(n10028), .A(n10026), .ZN(n10065) );
  NAND2_X1 U8598 ( .A1(n10066), .A2(n10065), .ZN(n6875) );
  NAND2_X1 U8599 ( .A1(n6876), .A2(n6875), .ZN(n10069) );
  NAND2_X1 U8600 ( .A1(n10070), .A2(n10069), .ZN(n6877) );
  NAND2_X1 U8601 ( .A1(n6878), .A2(n6877), .ZN(n10071) );
  NOR2_X1 U8602 ( .A1(n10072), .A2(n10071), .ZN(n6879) );
  NOR2_X1 U8603 ( .A1(n6880), .A2(n6879), .ZN(n6881) );
  NOR2_X1 U8604 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n6881), .ZN(n10055) );
  AND2_X1 U8605 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n6881), .ZN(n10054) );
  NOR2_X1 U8606 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10054), .ZN(n6882) );
  NOR2_X1 U8607 ( .A1(n10055), .A2(n6882), .ZN(n6883) );
  NAND2_X1 U8608 ( .A1(n6883), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n6885) );
  XOR2_X1 U8609 ( .A(n6883), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10053) );
  NAND2_X1 U8610 ( .A1(n10053), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n6884) );
  NAND2_X1 U8611 ( .A1(n6885), .A2(n6884), .ZN(n6886) );
  NAND2_X1 U8612 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n6886), .ZN(n6888) );
  XOR2_X1 U8613 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n6886), .Z(n10067) );
  NAND2_X1 U8614 ( .A1(n10067), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n6887) );
  NAND2_X1 U8615 ( .A1(n6888), .A2(n6887), .ZN(n6889) );
  NAND2_X1 U8616 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n6889), .ZN(n6891) );
  INV_X1 U8617 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9628) );
  XNOR2_X1 U8618 ( .A(n9628), .B(n6889), .ZN(n10068) );
  NAND2_X1 U8619 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10068), .ZN(n6890) );
  NAND2_X1 U8620 ( .A1(n6891), .A2(n6890), .ZN(n6892) );
  AND2_X1 U8621 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n6892), .ZN(n6893) );
  XNOR2_X1 U8622 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n6892), .ZN(n10059) );
  NOR2_X1 U8623 ( .A1(n10059), .A2(n10058), .ZN(n10057) );
  NAND2_X1 U8624 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n6894) );
  OAI21_X1 U8625 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n6894), .ZN(n10051) );
  NAND2_X1 U8626 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n6895) );
  OAI21_X1 U8627 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n6895), .ZN(n10048) );
  NOR2_X1 U8628 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n6896) );
  AOI21_X1 U8629 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n6896), .ZN(n10045) );
  NAND2_X1 U8630 ( .A1(n10046), .A2(n10045), .ZN(n10044) );
  OAI21_X1 U8631 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10044), .ZN(n10042) );
  NAND2_X1 U8632 ( .A1(n10043), .A2(n10042), .ZN(n10041) );
  OAI21_X1 U8633 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10041), .ZN(n10039) );
  NAND2_X1 U8634 ( .A1(n10040), .A2(n10039), .ZN(n10038) );
  OAI21_X1 U8635 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10038), .ZN(n10036) );
  NAND2_X1 U8636 ( .A1(n10037), .A2(n10036), .ZN(n10035) );
  OAI21_X1 U8637 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10035), .ZN(n10033) );
  NAND2_X1 U8638 ( .A1(n10034), .A2(n10033), .ZN(n10032) );
  OAI21_X1 U8639 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n10032), .ZN(n10030) );
  NAND2_X1 U8640 ( .A1(n10031), .A2(n10030), .ZN(n10029) );
  OAI21_X1 U8641 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10029), .ZN(n10061) );
  NOR2_X1 U8642 ( .A1(n10062), .A2(n10061), .ZN(n6897) );
  NAND2_X1 U8643 ( .A1(n10062), .A2(n10061), .ZN(n10060) );
  OAI21_X1 U8644 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n6897), .A(n10060), .ZN(
        n6900) );
  XNOR2_X1 U8645 ( .A(n6898), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n6899) );
  XNOR2_X1 U8646 ( .A(n6900), .B(n6899), .ZN(ADD_1071_U4) );
  OAI21_X1 U8647 ( .B1(n6902), .B2(n6767), .A(n6901), .ZN(n6906) );
  XNOR2_X1 U8648 ( .A(n6904), .B(n6903), .ZN(n6905) );
  XNOR2_X1 U8649 ( .A(n6906), .B(n6905), .ZN(n6914) );
  NOR2_X1 U8650 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6907), .ZN(n9611) );
  INV_X1 U8651 ( .A(n9611), .ZN(n6908) );
  OAI21_X1 U8652 ( .B1(n9000), .B2(n6909), .A(n6908), .ZN(n6911) );
  OAI22_X1 U8653 ( .A1(n9722), .A2(n8953), .B1(n8994), .B2(n9773), .ZN(n6910)
         );
  AOI211_X1 U8654 ( .C1(n6912), .C2(n8997), .A(n6911), .B(n6910), .ZN(n6913)
         );
  OAI21_X1 U8655 ( .B1(n6914), .B2(n8988), .A(n6913), .ZN(P1_U3237) );
  XNOR2_X1 U8656 ( .A(n6915), .B(n7594), .ZN(n9840) );
  INV_X1 U8657 ( .A(n9840), .ZN(n6927) );
  INV_X1 U8658 ( .A(n9770), .ZN(n9749) );
  INV_X1 U8659 ( .A(n6916), .ZN(n9725) );
  AOI21_X1 U8660 ( .B1(n7594), .B2(n6917), .A(n9725), .ZN(n6918) );
  OAI222_X1 U8661 ( .A1(n9772), .A2(n7044), .B1(n9774), .B2(n6919), .C1(n9749), 
        .C2(n6918), .ZN(n9838) );
  OAI211_X1 U8662 ( .C1(n6920), .C2(n9837), .A(n9828), .B(n9716), .ZN(n9836)
         );
  AOI22_X1 U8663 ( .A1(n9755), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n6921), .B2(
        n9783), .ZN(n6924) );
  NAND2_X1 U8664 ( .A1(n9494), .A2(n6922), .ZN(n6923) );
  OAI211_X1 U8665 ( .C1(n9836), .C2(n9500), .A(n6924), .B(n6923), .ZN(n6925)
         );
  AOI21_X1 U8666 ( .B1(n9838), .B2(n9779), .A(n6925), .ZN(n6926) );
  OAI21_X1 U8667 ( .B1(n6927), .B2(n9290), .A(n6926), .ZN(P1_U3284) );
  INV_X1 U8668 ( .A(n7417), .ZN(n6928) );
  OAI222_X1 U8669 ( .A1(n8827), .A2(n7418), .B1(n8835), .B2(n6928), .C1(
        P2_U3152), .C2(n8531), .ZN(P2_U3336) );
  OAI222_X1 U8670 ( .A1(n9401), .A2(n6929), .B1(n9397), .B2(n6928), .C1(
        P1_U3084), .C2(n7788), .ZN(P1_U3331) );
  XNOR2_X1 U8671 ( .A(n6930), .B(n7733), .ZN(n6931) );
  OAI222_X1 U8672 ( .A1(n9772), .A2(n6932), .B1(n9774), .B2(n7044), .C1(n9749), 
        .C2(n6931), .ZN(n9853) );
  INV_X1 U8673 ( .A(n9853), .ZN(n6939) );
  XNOR2_X1 U8674 ( .A(n6933), .B(n7733), .ZN(n9856) );
  INV_X1 U8675 ( .A(n9290), .ZN(n9505) );
  INV_X1 U8676 ( .A(n9717), .ZN(n6934) );
  OAI21_X1 U8677 ( .B1(n6934), .B2(n9850), .A(n7082), .ZN(n9852) );
  AOI22_X1 U8678 ( .A1(n9755), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7041), .B2(
        n9783), .ZN(n6936) );
  NAND2_X1 U8679 ( .A1(n9494), .A2(n7046), .ZN(n6935) );
  OAI211_X1 U8680 ( .C1(n9852), .C2(n9762), .A(n6936), .B(n6935), .ZN(n6937)
         );
  AOI21_X1 U8681 ( .B1(n9856), .B2(n9505), .A(n6937), .ZN(n6938) );
  OAI21_X1 U8682 ( .B1(n6939), .B2(n9755), .A(n6938), .ZN(P1_U3282) );
  INV_X1 U8683 ( .A(n6993), .ZN(n8182) );
  NAND2_X1 U8684 ( .A1(n6973), .A2(n8182), .ZN(n6944) );
  AND2_X1 U8685 ( .A1(n6946), .A2(n6944), .ZN(n6947) );
  NAND2_X1 U8686 ( .A1(n6940), .A2(n7839), .ZN(n6943) );
  AOI22_X1 U8687 ( .A1(n7370), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7369), .B2(
        n6941), .ZN(n6942) );
  NAND2_X1 U8688 ( .A1(n6943), .A2(n6942), .ZN(n7105) );
  OR2_X1 U8689 ( .A1(n7105), .A2(n7112), .ZN(n7902) );
  NAND2_X1 U8690 ( .A1(n7105), .A2(n7112), .ZN(n7903) );
  NAND2_X1 U8691 ( .A1(n7902), .A2(n7903), .ZN(n8005) );
  AND2_X1 U8692 ( .A1(n8005), .A2(n6944), .ZN(n6945) );
  NAND2_X1 U8693 ( .A1(n6946), .A2(n6945), .ZN(n7107) );
  OAI21_X1 U8694 ( .B1(n6947), .B2(n8005), .A(n7107), .ZN(n10000) );
  INV_X1 U8695 ( .A(n10000), .ZN(n6964) );
  NAND2_X1 U8696 ( .A1(n7832), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6954) );
  INV_X1 U8697 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6948) );
  NAND2_X1 U8698 ( .A1(n6949), .A2(n6948), .ZN(n6950) );
  AND2_X1 U8699 ( .A1(n7063), .A2(n6950), .ZN(n7119) );
  NAND2_X1 U8700 ( .A1(n6143), .A2(n7119), .ZN(n6953) );
  NAND2_X1 U8701 ( .A1(n7244), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6952) );
  NAND2_X1 U8702 ( .A1(n6802), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6951) );
  INV_X1 U8703 ( .A(n7898), .ZN(n6955) );
  XOR2_X1 U8704 ( .A(n8005), .B(n7111), .Z(n6957) );
  OAI222_X1 U8705 ( .A1(n8455), .A2(n6993), .B1(n8457), .B2(n8179), .C1(n8512), 
        .C2(n6957), .ZN(n9998) );
  INV_X1 U8706 ( .A(n6958), .ZN(n6959) );
  INV_X1 U8707 ( .A(n7105), .ZN(n9995) );
  OR2_X2 U8708 ( .A1(n6958), .A2(n7105), .ZN(n7117) );
  OAI21_X1 U8709 ( .B1(n6959), .B2(n9995), .A(n7117), .ZN(n9997) );
  AOI22_X1 U8710 ( .A1(n4305), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7014), .B2(
        n9435), .ZN(n6961) );
  NAND2_X1 U8711 ( .A1(n8484), .A2(n7105), .ZN(n6960) );
  OAI211_X1 U8712 ( .C1(n9997), .C2(n8443), .A(n6961), .B(n6960), .ZN(n6962)
         );
  AOI21_X1 U8713 ( .B1(n9998), .B2(n9441), .A(n6962), .ZN(n6963) );
  OAI21_X1 U8714 ( .B1(n6964), .B2(n9444), .A(n6963), .ZN(P2_U3284) );
  XNOR2_X1 U8715 ( .A(n6994), .B(n7390), .ZN(n6968) );
  NOR2_X1 U8716 ( .A1(n6979), .A2(n9913), .ZN(n6969) );
  NAND2_X1 U8717 ( .A1(n6968), .A2(n6969), .ZN(n6974) );
  INV_X1 U8718 ( .A(n6968), .ZN(n6971) );
  INV_X1 U8719 ( .A(n6969), .ZN(n6970) );
  NAND2_X1 U8720 ( .A1(n6971), .A2(n6970), .ZN(n6972) );
  NAND2_X1 U8721 ( .A1(n6974), .A2(n6972), .ZN(n6990) );
  OR2_X1 U8722 ( .A1(n7057), .A2(n6990), .ZN(n6988) );
  NAND2_X1 U8723 ( .A1(n6988), .A2(n6974), .ZN(n6978) );
  NOR2_X1 U8724 ( .A1(n6993), .A2(n9913), .ZN(n7004) );
  OR2_X1 U8725 ( .A1(n7057), .A2(n7050), .ZN(n7008) );
  OR2_X1 U8726 ( .A1(n6975), .A2(n6974), .ZN(n7006) );
  AND2_X1 U8727 ( .A1(n7008), .A2(n7006), .ZN(n6976) );
  OAI211_X1 U8728 ( .C1(n6978), .C2(n6977), .A(n6976), .B(n8150), .ZN(n6984)
         );
  NOR2_X1 U8729 ( .A1(n8156), .A2(n6979), .ZN(n6981) );
  OAI22_X1 U8730 ( .A1(n8145), .A2(n7112), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8197), .ZN(n6980) );
  AOI211_X1 U8731 ( .C1(n8158), .C2(n6982), .A(n6981), .B(n6980), .ZN(n6983)
         );
  OAI211_X1 U8732 ( .C1(n9988), .C2(n8161), .A(n6984), .B(n6983), .ZN(P2_U3238) );
  INV_X1 U8733 ( .A(n7430), .ZN(n6987) );
  NOR2_X1 U8734 ( .A1(n6985), .A2(P1_U3084), .ZN(n7791) );
  AOI21_X1 U8735 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9390), .A(n7791), .ZN(
        n6986) );
  OAI21_X1 U8736 ( .B1(n6987), .B2(n9397), .A(n6986), .ZN(P1_U3330) );
  INV_X1 U8737 ( .A(n6988), .ZN(n6989) );
  AOI211_X1 U8738 ( .C1(n6990), .C2(n7057), .A(n9882), .B(n6989), .ZN(n6998)
         );
  INV_X1 U8739 ( .A(n8156), .ZN(n8143) );
  NAND2_X1 U8740 ( .A1(n8143), .A2(n8184), .ZN(n6992) );
  OAI211_X1 U8741 ( .C1(n6993), .C2(n8145), .A(n6992), .B(n6991), .ZN(n6997)
         );
  INV_X1 U8742 ( .A(n6994), .ZN(n9980) );
  OAI22_X1 U8743 ( .A1(n8161), .A2(n9980), .B1(n9891), .B2(n6995), .ZN(n6996)
         );
  OR3_X1 U8744 ( .A1(n6998), .A2(n6997), .A3(n6996), .ZN(P2_U3219) );
  XNOR2_X1 U8745 ( .A(n7105), .B(n7798), .ZN(n6999) );
  OR2_X1 U8746 ( .A1(n7112), .A2(n9913), .ZN(n7000) );
  NAND2_X1 U8747 ( .A1(n6999), .A2(n7000), .ZN(n7049) );
  INV_X1 U8748 ( .A(n6999), .ZN(n7002) );
  INV_X1 U8749 ( .A(n7000), .ZN(n7001) );
  NAND2_X1 U8750 ( .A1(n7002), .A2(n7001), .ZN(n7053) );
  NAND2_X1 U8751 ( .A1(n7049), .A2(n7053), .ZN(n7010) );
  INV_X1 U8752 ( .A(n7003), .ZN(n7005) );
  NAND2_X1 U8753 ( .A1(n7005), .A2(n7004), .ZN(n7007) );
  AND2_X1 U8754 ( .A1(n7007), .A2(n7006), .ZN(n7051) );
  NAND2_X1 U8755 ( .A1(n7008), .A2(n7051), .ZN(n7009) );
  XOR2_X1 U8756 ( .A(n7010), .B(n7009), .Z(n7017) );
  NAND2_X1 U8757 ( .A1(n8143), .A2(n8182), .ZN(n7012) );
  OAI211_X1 U8758 ( .C1(n8179), .C2(n8145), .A(n7012), .B(n7011), .ZN(n7013)
         );
  AOI21_X1 U8759 ( .B1(n7014), .B2(n8158), .A(n7013), .ZN(n7016) );
  NAND2_X1 U8760 ( .A1(n9886), .A2(n7105), .ZN(n7015) );
  OAI211_X1 U8761 ( .C1(n7017), .C2(n9882), .A(n7016), .B(n7015), .ZN(P2_U3226) );
  INV_X1 U8762 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7018) );
  AOI22_X1 U8763 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7306), .B1(n7313), .B2(
        n7018), .ZN(n7022) );
  NAND2_X1 U8764 ( .A1(n7022), .A2(n7021), .ZN(n7305) );
  OAI21_X1 U8765 ( .B1(n7022), .B2(n7021), .A(n7305), .ZN(n7032) );
  NOR2_X1 U8766 ( .A1(n7059), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7023) );
  NOR2_X1 U8767 ( .A1(n7024), .A2(n7023), .ZN(n7026) );
  INV_X1 U8768 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9470) );
  AOI22_X1 U8769 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n7313), .B1(n7306), .B2(
        n9470), .ZN(n7025) );
  NOR2_X1 U8770 ( .A1(n7026), .A2(n7025), .ZN(n7312) );
  AOI21_X1 U8771 ( .B1(n7026), .B2(n7025), .A(n7312), .ZN(n7030) );
  NAND2_X1 U8772 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7184) );
  INV_X1 U8773 ( .A(n7184), .ZN(n7027) );
  AOI21_X1 U8774 ( .B1(n9898), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n7027), .ZN(
        n7029) );
  NAND2_X1 U8775 ( .A1(n9895), .A2(n7306), .ZN(n7028) );
  OAI211_X1 U8776 ( .C1(n9893), .C2(n7030), .A(n7029), .B(n7028), .ZN(n7031)
         );
  AOI21_X1 U8777 ( .B1(n9897), .B2(n7032), .A(n7031), .ZN(n7033) );
  INV_X1 U8778 ( .A(n7033), .ZN(P2_U3259) );
  NAND2_X1 U8779 ( .A1(n7430), .A2(n7034), .ZN(n7035) );
  OAI211_X1 U8780 ( .C1(n8702), .C2(n8827), .A(n7035), .B(n8030), .ZN(P2_U3335) );
  INV_X1 U8781 ( .A(n7037), .ZN(n7038) );
  AOI21_X1 U8782 ( .B1(n7039), .B2(n7036), .A(n7038), .ZN(n7048) );
  AOI21_X1 U8783 ( .B1(n8992), .B2(n9005), .A(n7040), .ZN(n7043) );
  NAND2_X1 U8784 ( .A1(n8997), .A2(n7041), .ZN(n7042) );
  OAI211_X1 U8785 ( .C1(n7044), .C2(n8994), .A(n7043), .B(n7042), .ZN(n7045)
         );
  AOI21_X1 U8786 ( .B1(n7046), .B2(n8965), .A(n7045), .ZN(n7047) );
  OAI21_X1 U8787 ( .B1(n7048), .B2(n8988), .A(n7047), .ZN(P1_U3229) );
  INV_X1 U8788 ( .A(n7049), .ZN(n7052) );
  OR2_X1 U8789 ( .A1(n7050), .A2(n7052), .ZN(n7056) );
  NAND2_X1 U8790 ( .A1(n7058), .A2(n7839), .ZN(n7061) );
  AOI22_X1 U8791 ( .A1(n7370), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7369), .B2(
        n7059), .ZN(n7060) );
  NAND2_X1 U8792 ( .A1(n7061), .A2(n7060), .ZN(n7116) );
  XNOR2_X1 U8793 ( .A(n7116), .B(n7798), .ZN(n7174) );
  NOR2_X1 U8794 ( .A1(n8179), .A2(n9913), .ZN(n7175) );
  XNOR2_X1 U8795 ( .A(n7174), .B(n7175), .ZN(n7172) );
  XNOR2_X1 U8796 ( .A(n7173), .B(n7172), .ZN(n7074) );
  NOR2_X1 U8797 ( .A1(n8161), .A2(n4535), .ZN(n7072) );
  INV_X1 U8798 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7062) );
  NAND2_X1 U8799 ( .A1(n7063), .A2(n7062), .ZN(n7064) );
  AND2_X1 U8800 ( .A1(n7153), .A2(n7064), .ZN(n7188) );
  NAND2_X1 U8801 ( .A1(n6143), .A2(n7188), .ZN(n7068) );
  NAND2_X1 U8802 ( .A1(n7832), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7067) );
  NAND2_X1 U8803 ( .A1(n7244), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7066) );
  NAND2_X1 U8804 ( .A1(n6802), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7065) );
  NAND4_X1 U8805 ( .A1(n7068), .A2(n7067), .A3(n7066), .A4(n7065), .ZN(n8178)
         );
  INV_X1 U8806 ( .A(n8178), .ZN(n7911) );
  INV_X1 U8807 ( .A(n7112), .ZN(n8181) );
  NAND2_X1 U8808 ( .A1(n8143), .A2(n8181), .ZN(n7070) );
  OAI211_X1 U8809 ( .C1(n7911), .C2(n8145), .A(n7070), .B(n7069), .ZN(n7071)
         );
  AOI211_X1 U8810 ( .C1(n8158), .C2(n7119), .A(n7072), .B(n7071), .ZN(n7073)
         );
  OAI21_X1 U8811 ( .B1(n7074), .B2(n9882), .A(n7073), .ZN(P2_U3236) );
  INV_X1 U8812 ( .A(n7626), .ZN(n7075) );
  AOI21_X1 U8813 ( .B1(n6930), .B2(n7609), .A(n7075), .ZN(n7076) );
  XNOR2_X1 U8814 ( .A(n7076), .B(n7736), .ZN(n7081) );
  OAI21_X1 U8815 ( .B1(n7078), .B2(n7736), .A(n7077), .ZN(n9430) );
  NAND2_X1 U8816 ( .A1(n9430), .A2(n9776), .ZN(n7080) );
  AOI22_X1 U8817 ( .A1(n9006), .A2(n9489), .B1(n9742), .B2(n9490), .ZN(n7079)
         );
  OAI211_X1 U8818 ( .C1(n9749), .C2(n7081), .A(n7080), .B(n7079), .ZN(n9428)
         );
  INV_X1 U8819 ( .A(n9428), .ZN(n7089) );
  INV_X1 U8820 ( .A(n7082), .ZN(n7084) );
  INV_X1 U8821 ( .A(n7098), .ZN(n7083) );
  OAI211_X1 U8822 ( .C1(n9427), .C2(n7084), .A(n7083), .B(n9828), .ZN(n9426)
         );
  AOI22_X1 U8823 ( .A1(n9755), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7134), .B2(
        n9783), .ZN(n7086) );
  NAND2_X1 U8824 ( .A1(n9494), .A2(n7133), .ZN(n7085) );
  OAI211_X1 U8825 ( .C1(n9426), .C2(n9500), .A(n7086), .B(n7085), .ZN(n7087)
         );
  AOI21_X1 U8826 ( .B1(n9430), .B2(n9764), .A(n7087), .ZN(n7088) );
  OAI21_X1 U8827 ( .B1(n7089), .B2(n9755), .A(n7088), .ZN(P1_U3281) );
  XNOR2_X1 U8828 ( .A(n9490), .B(n7226), .ZN(n7738) );
  XNOR2_X1 U8829 ( .A(n7090), .B(n7738), .ZN(n7097) );
  AOI22_X1 U8830 ( .A1(n9742), .A2(n9004), .B1(n9005), .B2(n9489), .ZN(n7096)
         );
  NAND2_X1 U8831 ( .A1(n7092), .A2(n7091), .ZN(n7093) );
  NAND2_X1 U8832 ( .A1(n7093), .A2(n7738), .ZN(n9487) );
  OAI21_X1 U8833 ( .B1(n7093), .B2(n7738), .A(n9487), .ZN(n7094) );
  NAND2_X1 U8834 ( .A1(n7094), .A2(n9770), .ZN(n7095) );
  OAI211_X1 U8835 ( .C1(n7097), .C2(n9730), .A(n7096), .B(n7095), .ZN(n9547)
         );
  INV_X1 U8836 ( .A(n9547), .ZN(n7104) );
  INV_X1 U8837 ( .A(n7097), .ZN(n9549) );
  OR2_X1 U8838 ( .A1(n7098), .A2(n9545), .ZN(n7099) );
  NAND2_X1 U8839 ( .A1(n9501), .A2(n7099), .ZN(n9546) );
  AOI22_X1 U8840 ( .A1(n9755), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7227), .B2(
        n9783), .ZN(n7101) );
  NAND2_X1 U8841 ( .A1(n9494), .A2(n7226), .ZN(n7100) );
  OAI211_X1 U8842 ( .C1(n9546), .C2(n9762), .A(n7101), .B(n7100), .ZN(n7102)
         );
  AOI21_X1 U8843 ( .B1(n9549), .B2(n9764), .A(n7102), .ZN(n7103) );
  OAI21_X1 U8844 ( .B1(n7104), .B2(n9755), .A(n7103), .ZN(P1_U3280) );
  OR2_X1 U8845 ( .A1(n7105), .A2(n8181), .ZN(n7106) );
  OR2_X1 U8846 ( .A1(n7116), .A2(n8179), .ZN(n7908) );
  NAND2_X1 U8847 ( .A1(n7116), .A2(n8179), .ZN(n7907) );
  NAND2_X1 U8848 ( .A1(n7108), .A2(n8003), .ZN(n7109) );
  NAND2_X1 U8849 ( .A1(n7147), .A2(n7109), .ZN(n9472) );
  INV_X1 U8850 ( .A(n7902), .ZN(n7110) );
  XNOR2_X1 U8851 ( .A(n7150), .B(n8003), .ZN(n7114) );
  OAI22_X1 U8852 ( .A1(n7911), .A2(n8457), .B1(n7112), .B2(n8455), .ZN(n7113)
         );
  AOI21_X1 U8853 ( .B1(n7114), .B2(n8608), .A(n7113), .ZN(n7115) );
  OAI21_X1 U8854 ( .B1(n9472), .B2(n8533), .A(n7115), .ZN(n9474) );
  NAND2_X1 U8855 ( .A1(n9474), .A2(n9441), .ZN(n7124) );
  AND2_X1 U8856 ( .A1(n7117), .A2(n7116), .ZN(n7118) );
  OR2_X1 U8857 ( .A1(n7118), .A2(n7162), .ZN(n9473) );
  INV_X1 U8858 ( .A(n9473), .ZN(n7122) );
  AOI22_X1 U8859 ( .A1(n4305), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7119), .B2(
        n9435), .ZN(n7120) );
  OAI21_X1 U8860 ( .B1(n4535), .B2(n9438), .A(n7120), .ZN(n7121) );
  AOI21_X1 U8861 ( .B1(n7122), .B2(n8494), .A(n7121), .ZN(n7123) );
  OAI211_X1 U8862 ( .C1(n9472), .C2(n8487), .A(n7124), .B(n7123), .ZN(P2_U3283) );
  INV_X1 U8863 ( .A(n7353), .ZN(n7142) );
  OAI222_X1 U8864 ( .A1(n9397), .A2(n7142), .B1(P1_U3084), .B2(n7126), .C1(
        n7125), .C2(n9401), .ZN(P1_U3329) );
  NAND2_X1 U8865 ( .A1(n7128), .A2(n7127), .ZN(n7130) );
  XOR2_X1 U8866 ( .A(n7130), .B(n7129), .Z(n7140) );
  INV_X1 U8867 ( .A(n7131), .ZN(n7132) );
  AOI21_X1 U8868 ( .B1(n8992), .B2(n9490), .A(n7132), .ZN(n7138) );
  NAND2_X1 U8869 ( .A1(n8965), .A2(n7133), .ZN(n7137) );
  NAND2_X1 U8870 ( .A1(n8997), .A2(n7134), .ZN(n7136) );
  NAND2_X1 U8871 ( .A1(n8966), .A2(n9006), .ZN(n7135) );
  NAND4_X1 U8872 ( .A1(n7138), .A2(n7137), .A3(n7136), .A4(n7135), .ZN(n7139)
         );
  AOI21_X1 U8873 ( .B1(n7140), .B2(n8977), .A(n7139), .ZN(n7141) );
  INV_X1 U8874 ( .A(n7141), .ZN(P1_U3215) );
  OAI222_X1 U8875 ( .A1(n7143), .A2(P2_U3152), .B1(n8835), .B2(n7142), .C1(
        n7354), .C2(n8827), .ZN(P2_U3334) );
  NAND2_X1 U8876 ( .A1(n7144), .A2(n7839), .ZN(n7146) );
  AOI22_X1 U8877 ( .A1(n7370), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7369), .B2(
        n7306), .ZN(n7145) );
  XNOR2_X1 U8878 ( .A(n7913), .B(n8178), .ZN(n8008) );
  AOI21_X1 U8879 ( .B1(n8008), .B2(n7148), .A(n7235), .ZN(n9464) );
  INV_X1 U8880 ( .A(n7907), .ZN(n7149) );
  AOI21_X1 U8881 ( .B1(n7150), .B2(n8003), .A(n7149), .ZN(n7151) );
  OAI211_X1 U8882 ( .C1(n7151), .C2(n8008), .A(n7240), .B(n8608), .ZN(n7160)
         );
  NAND2_X1 U8883 ( .A1(n7832), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7158) );
  NAND2_X1 U8884 ( .A1(n7153), .A2(n7152), .ZN(n7154) );
  AND2_X1 U8885 ( .A1(n7242), .A2(n7154), .ZN(n8165) );
  NAND2_X1 U8886 ( .A1(n6143), .A2(n8165), .ZN(n7157) );
  NAND2_X1 U8887 ( .A1(n7244), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7156) );
  NAND2_X1 U8888 ( .A1(n6802), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7155) );
  NAND2_X1 U8889 ( .A1(n8606), .A2(n8603), .ZN(n7159) );
  OAI211_X1 U8890 ( .C1(n8179), .C2(n8455), .A(n7160), .B(n7159), .ZN(n9468)
         );
  INV_X1 U8891 ( .A(n7252), .ZN(n7161) );
  OAI21_X1 U8892 ( .B1(n9465), .B2(n7162), .A(n7161), .ZN(n9466) );
  AOI22_X1 U8893 ( .A1(n4305), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7188), .B2(
        n9435), .ZN(n7164) );
  NAND2_X1 U8894 ( .A1(n8484), .A2(n7913), .ZN(n7163) );
  OAI211_X1 U8895 ( .C1(n9466), .C2(n8443), .A(n7164), .B(n7163), .ZN(n7165)
         );
  AOI21_X1 U8896 ( .B1(n9468), .B2(n9441), .A(n7165), .ZN(n7166) );
  OAI21_X1 U8897 ( .B1(n9464), .B2(n9444), .A(n7166), .ZN(P2_U3282) );
  XNOR2_X1 U8898 ( .A(n7913), .B(n7798), .ZN(n7167) );
  NAND2_X1 U8899 ( .A1(n8178), .A2(n7444), .ZN(n7168) );
  NAND2_X1 U8900 ( .A1(n7167), .A2(n7168), .ZN(n7269) );
  INV_X1 U8901 ( .A(n7167), .ZN(n7170) );
  INV_X1 U8902 ( .A(n7168), .ZN(n7169) );
  NAND2_X1 U8903 ( .A1(n7170), .A2(n7169), .ZN(n7171) );
  NAND2_X1 U8904 ( .A1(n7269), .A2(n7171), .ZN(n7183) );
  INV_X1 U8905 ( .A(n7174), .ZN(n7176) );
  NAND2_X1 U8906 ( .A1(n7176), .A2(n7175), .ZN(n7177) );
  NAND2_X1 U8907 ( .A1(n7178), .A2(n7177), .ZN(n7182) );
  INV_X1 U8908 ( .A(n7270), .ZN(n7181) );
  AOI21_X1 U8909 ( .B1(n7183), .B2(n7182), .A(n7181), .ZN(n7190) );
  NAND2_X1 U8910 ( .A1(n8154), .A2(n8606), .ZN(n7185) );
  OAI211_X1 U8911 ( .C1(n8179), .C2(n8156), .A(n7185), .B(n7184), .ZN(n7187)
         );
  NOR2_X1 U8912 ( .A1(n9465), .A2(n8161), .ZN(n7186) );
  AOI211_X1 U8913 ( .C1(n8158), .C2(n7188), .A(n7187), .B(n7186), .ZN(n7189)
         );
  OAI21_X1 U8914 ( .B1(n7190), .B2(n9882), .A(n7189), .ZN(P2_U3217) );
  XNOR2_X1 U8915 ( .A(n7191), .B(n4550), .ZN(n9535) );
  NAND2_X1 U8916 ( .A1(n7193), .A2(n7192), .ZN(n7194) );
  NAND2_X1 U8917 ( .A1(n7207), .A2(n7194), .ZN(n7195) );
  NAND2_X1 U8918 ( .A1(n7195), .A2(n9770), .ZN(n7197) );
  AOI22_X1 U8919 ( .A1(n9004), .A2(n9489), .B1(n9742), .B2(n9275), .ZN(n7196)
         );
  NAND2_X1 U8920 ( .A1(n7197), .A2(n7196), .ZN(n7198) );
  AOI21_X1 U8921 ( .B1(n9535), .B2(n9776), .A(n7198), .ZN(n9537) );
  AND2_X1 U8922 ( .A1(n9502), .A2(n8938), .ZN(n7199) );
  OR2_X1 U8923 ( .A1(n7199), .A2(n7211), .ZN(n9533) );
  AOI22_X1 U8924 ( .A1(n9755), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8939), .B2(
        n9783), .ZN(n7201) );
  NAND2_X1 U8925 ( .A1(n8938), .A2(n9494), .ZN(n7200) );
  OAI211_X1 U8926 ( .C1(n9533), .C2(n9762), .A(n7201), .B(n7200), .ZN(n7202)
         );
  AOI21_X1 U8927 ( .B1(n9535), .B2(n9764), .A(n7202), .ZN(n7203) );
  OAI21_X1 U8928 ( .B1(n9537), .B2(n9755), .A(n7203), .ZN(P1_U3278) );
  XOR2_X1 U8929 ( .A(n7204), .B(n7740), .Z(n9530) );
  INV_X1 U8930 ( .A(n9530), .ZN(n7219) );
  NAND2_X1 U8931 ( .A1(n7205), .A2(n9770), .ZN(n7210) );
  INV_X1 U8932 ( .A(n7740), .ZN(n7206) );
  AOI21_X1 U8933 ( .B1(n7207), .B2(n7538), .A(n7206), .ZN(n7209) );
  AOI22_X1 U8934 ( .A1(n9491), .A2(n9489), .B1(n9742), .B2(n9262), .ZN(n7208)
         );
  OAI21_X1 U8935 ( .B1(n7210), .B2(n7209), .A(n7208), .ZN(n9529) );
  OAI21_X1 U8936 ( .B1(n7211), .B2(n9527), .A(n9828), .ZN(n7212) );
  OR2_X1 U8937 ( .A1(n7212), .A2(n9279), .ZN(n9526) );
  INV_X1 U8938 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7214) );
  INV_X1 U8939 ( .A(n8849), .ZN(n7213) );
  OAI22_X1 U8940 ( .A1(n9779), .A2(n7214), .B1(n7213), .B2(n9283), .ZN(n7215)
         );
  AOI21_X1 U8941 ( .B1(n8848), .B2(n9494), .A(n7215), .ZN(n7216) );
  OAI21_X1 U8942 ( .B1(n9526), .B2(n9500), .A(n7216), .ZN(n7217) );
  AOI21_X1 U8943 ( .B1(n9529), .B2(n9779), .A(n7217), .ZN(n7218) );
  OAI21_X1 U8944 ( .B1(n7219), .B2(n9290), .A(n7218), .ZN(P1_U3277) );
  INV_X1 U8945 ( .A(n7220), .ZN(n7221) );
  AOI211_X1 U8946 ( .C1(n7223), .C2(n7222), .A(n8988), .B(n7221), .ZN(n7233)
         );
  INV_X1 U8947 ( .A(n7224), .ZN(n7225) );
  AOI21_X1 U8948 ( .B1(n8992), .B2(n9004), .A(n7225), .ZN(n7231) );
  NAND2_X1 U8949 ( .A1(n8965), .A2(n7226), .ZN(n7230) );
  NAND2_X1 U8950 ( .A1(n8997), .A2(n7227), .ZN(n7229) );
  NAND2_X1 U8951 ( .A1(n8966), .A2(n9005), .ZN(n7228) );
  NAND4_X1 U8952 ( .A1(n7231), .A2(n7230), .A3(n7229), .A4(n7228), .ZN(n7232)
         );
  OR2_X1 U8953 ( .A1(n7233), .A2(n7232), .ZN(P1_U3234) );
  NAND2_X1 U8954 ( .A1(n7236), .A2(n7839), .ZN(n7238) );
  AOI22_X1 U8955 ( .A1(n7370), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7369), .B2(
        n8214), .ZN(n7237) );
  OR2_X1 U8956 ( .A1(n8280), .A2(n8101), .ZN(n7921) );
  NAND2_X1 U8957 ( .A1(n8280), .A2(n8101), .ZN(n8600) );
  XNOR2_X1 U8958 ( .A(n8283), .B(n8282), .ZN(n9462) );
  INV_X1 U8959 ( .A(n9462), .ZN(n7257) );
  OR2_X1 U8960 ( .A1(n7913), .A2(n7911), .ZN(n7239) );
  XNOR2_X1 U8961 ( .A(n7813), .B(n8282), .ZN(n7251) );
  NAND2_X1 U8962 ( .A1(n7832), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7248) );
  INV_X1 U8963 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7241) );
  NAND2_X1 U8964 ( .A1(n7242), .A2(n7241), .ZN(n7243) );
  AND2_X1 U8965 ( .A1(n7286), .A2(n7243), .ZN(n9436) );
  NAND2_X1 U8966 ( .A1(n6143), .A2(n9436), .ZN(n7247) );
  NAND2_X1 U8967 ( .A1(n7244), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7246) );
  NAND2_X1 U8968 ( .A1(n6802), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7245) );
  NAND2_X1 U8969 ( .A1(n8178), .A2(n8605), .ZN(n7249) );
  OAI21_X1 U8970 ( .B1(n8177), .B2(n8457), .A(n7249), .ZN(n8166) );
  INV_X1 U8971 ( .A(n8166), .ZN(n7250) );
  OAI21_X1 U8972 ( .B1(n7251), .B2(n8512), .A(n7250), .ZN(n9461) );
  INV_X1 U8973 ( .A(n8280), .ZN(n9458) );
  OAI21_X1 U8974 ( .B1(n7252), .B2(n9458), .A(n4336), .ZN(n9459) );
  AOI22_X1 U8975 ( .A1(n4305), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8165), .B2(
        n9435), .ZN(n7254) );
  NAND2_X1 U8976 ( .A1(n8280), .A2(n8484), .ZN(n7253) );
  OAI211_X1 U8977 ( .C1(n9459), .C2(n8443), .A(n7254), .B(n7253), .ZN(n7255)
         );
  AOI21_X1 U8978 ( .B1(n9461), .B2(n9441), .A(n7255), .ZN(n7256) );
  OAI21_X1 U8979 ( .B1(n7257), .B2(n9444), .A(n7256), .ZN(P2_U3281) );
  INV_X1 U8980 ( .A(n7258), .ZN(n7259) );
  AOI21_X1 U8981 ( .B1(n7261), .B2(n7260), .A(n7259), .ZN(n7268) );
  NOR2_X1 U8982 ( .A1(n9000), .A2(n9541), .ZN(n7266) );
  NAND2_X1 U8983 ( .A1(n8966), .A2(n9490), .ZN(n7263) );
  OAI211_X1 U8984 ( .C1(n7264), .C2(n8953), .A(n7263), .B(n7262), .ZN(n7265)
         );
  AOI211_X1 U8985 ( .C1(n9493), .C2(n8997), .A(n7266), .B(n7265), .ZN(n7267)
         );
  OAI21_X1 U8986 ( .B1(n7268), .B2(n8988), .A(n7267), .ZN(P1_U3222) );
  XNOR2_X1 U8987 ( .A(n8280), .B(n7798), .ZN(n8091) );
  OR2_X1 U8988 ( .A1(n8101), .A2(n9913), .ZN(n7275) );
  NAND2_X1 U8989 ( .A1(n8091), .A2(n7275), .ZN(n7271) );
  NAND2_X1 U8990 ( .A1(n7272), .A2(n7839), .ZN(n7274) );
  AOI22_X1 U8991 ( .A1(n7370), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7369), .B2(
        n8220), .ZN(n7273) );
  XNOR2_X1 U8992 ( .A(n8610), .B(n7798), .ZN(n7281) );
  NOR2_X1 U8993 ( .A1(n8177), .A2(n9913), .ZN(n7279) );
  XNOR2_X1 U8994 ( .A(n7281), .B(n7279), .ZN(n8094) );
  INV_X1 U8995 ( .A(n8091), .ZN(n7276) );
  INV_X1 U8996 ( .A(n7275), .ZN(n8164) );
  NAND2_X1 U8997 ( .A1(n7276), .A2(n8164), .ZN(n7277) );
  AND2_X1 U8998 ( .A1(n8094), .A2(n7277), .ZN(n7278) );
  INV_X1 U8999 ( .A(n7279), .ZN(n7280) );
  NAND2_X1 U9000 ( .A1(n7281), .A2(n7280), .ZN(n7282) );
  NAND2_X1 U9001 ( .A1(n7283), .A2(n7839), .ZN(n7285) );
  AOI22_X1 U9002 ( .A1(n7370), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7369), .B2(
        n8240), .ZN(n7284) );
  XNOR2_X1 U9003 ( .A(n8594), .B(n7390), .ZN(n7358) );
  NAND2_X1 U9004 ( .A1(n7286), .A2(n8224), .ZN(n7287) );
  AND2_X1 U9005 ( .A1(n7293), .A2(n7287), .ZN(n8506) );
  NAND2_X1 U9006 ( .A1(n6143), .A2(n8506), .ZN(n7291) );
  NAND2_X1 U9007 ( .A1(n7832), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7290) );
  NAND2_X1 U9008 ( .A1(n7244), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7289) );
  NAND2_X1 U9009 ( .A1(n6802), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n7288) );
  NOR2_X1 U9010 ( .A1(n8098), .A2(n9913), .ZN(n7357) );
  XNOR2_X1 U9011 ( .A(n7358), .B(n7357), .ZN(n7360) );
  XNOR2_X1 U9012 ( .A(n7361), .B(n7360), .ZN(n7304) );
  INV_X1 U9013 ( .A(n8506), .ZN(n7301) );
  NAND2_X1 U9014 ( .A1(n7832), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7298) );
  INV_X1 U9015 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7292) );
  NAND2_X1 U9016 ( .A1(n7293), .A2(n7292), .ZN(n7294) );
  AND2_X1 U9017 ( .A1(n7374), .A2(n7294), .ZN(n8495) );
  NAND2_X1 U9018 ( .A1(n6143), .A2(n8495), .ZN(n7297) );
  NAND2_X1 U9019 ( .A1(n7244), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7296) );
  NAND2_X1 U9020 ( .A1(n6802), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7295) );
  OR2_X1 U9021 ( .A1(n8177), .A2(n8455), .ZN(n7299) );
  OAI21_X1 U9022 ( .B1(n8287), .B2(n8457), .A(n7299), .ZN(n8515) );
  AOI22_X1 U9023 ( .A1(n9881), .A2(n8515), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n7300) );
  OAI21_X1 U9024 ( .B1(n7301), .B2(n9891), .A(n7300), .ZN(n7302) );
  AOI21_X1 U9025 ( .B1(n8594), .B2(n9886), .A(n7302), .ZN(n7303) );
  OAI21_X1 U9026 ( .B1(n7304), .B2(n9882), .A(n7303), .ZN(P2_U3230) );
  OAI21_X1 U9027 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7306), .A(n7305), .ZN(
        n7307) );
  NAND2_X1 U9028 ( .A1(n7314), .A2(n7307), .ZN(n7308) );
  XNOR2_X1 U9029 ( .A(n8214), .B(n7307), .ZN(n8212) );
  INV_X1 U9030 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8211) );
  NAND2_X1 U9031 ( .A1(n8212), .A2(n8211), .ZN(n8210) );
  NAND2_X1 U9032 ( .A1(n7308), .A2(n8210), .ZN(n7311) );
  NAND2_X1 U9033 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8220), .ZN(n7309) );
  OAI21_X1 U9034 ( .B1(n8220), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7309), .ZN(
        n7310) );
  NOR2_X1 U9035 ( .A1(n7310), .A2(n7311), .ZN(n8219) );
  AOI211_X1 U9036 ( .C1(n7311), .C2(n7310), .A(n8219), .B(n9414), .ZN(n7324)
         );
  AOI21_X1 U9037 ( .B1(n9470), .B2(n7313), .A(n7312), .ZN(n7315) );
  NAND2_X1 U9038 ( .A1(n8214), .A2(n7315), .ZN(n7316) );
  XNOR2_X1 U9039 ( .A(n7315), .B(n7314), .ZN(n8208) );
  NAND2_X1 U9040 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8208), .ZN(n8207) );
  NAND2_X1 U9041 ( .A1(n7316), .A2(n8207), .ZN(n7318) );
  XNOR2_X1 U9042 ( .A(n8220), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n7317) );
  NOR2_X1 U9043 ( .A1(n7317), .A2(n7318), .ZN(n8226) );
  AOI21_X1 U9044 ( .B1(n7318), .B2(n7317), .A(n8226), .ZN(n7322) );
  NAND2_X1 U9045 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8099) );
  INV_X1 U9046 ( .A(n8099), .ZN(n7319) );
  AOI21_X1 U9047 ( .B1(n9898), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7319), .ZN(
        n7321) );
  NAND2_X1 U9048 ( .A1(n9895), .A2(n8220), .ZN(n7320) );
  OAI211_X1 U9049 ( .C1(n7322), .C2(n9893), .A(n7321), .B(n7320), .ZN(n7323)
         );
  OR2_X1 U9050 ( .A1(n7324), .A2(n7323), .ZN(P2_U3261) );
  INV_X1 U9051 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7332) );
  INV_X1 U9052 ( .A(SI_29_), .ZN(n7325) );
  AND2_X1 U9053 ( .A1(n7328), .A2(n7325), .ZN(n7326) );
  INV_X1 U9054 ( .A(n7328), .ZN(n7329) );
  NAND2_X1 U9055 ( .A1(n7329), .A2(SI_29_), .ZN(n7330) );
  MUX2_X1 U9056 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7501), .Z(n7497) );
  INV_X1 U9057 ( .A(n7829), .ZN(n8825) );
  OAI222_X1 U9058 ( .A1(n9401), .A2(n7332), .B1(n9397), .B2(n8825), .C1(
        P1_U3084), .C2(n7331), .ZN(P1_U3323) );
  NAND2_X1 U9059 ( .A1(n8831), .A2(n7839), .ZN(n7334) );
  NAND2_X2 U9060 ( .A1(n7334), .A2(n7333), .ZN(n8542) );
  INV_X1 U9061 ( .A(n8542), .ZN(n8341) );
  XNOR2_X1 U9062 ( .A(n8542), .B(n7798), .ZN(n7344) );
  INV_X1 U9063 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7335) );
  NAND2_X1 U9064 ( .A1(n7469), .A2(n7335), .ZN(n7336) );
  NAND2_X1 U9065 ( .A1(n7479), .A2(n7336), .ZN(n7477) );
  INV_X1 U9066 ( .A(n6143), .ZN(n7453) );
  INV_X1 U9067 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n7339) );
  NAND2_X1 U9068 ( .A1(n6802), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n7338) );
  NAND2_X1 U9069 ( .A1(n7244), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7337) );
  OAI211_X1 U9070 ( .C1(n7485), .C2(n7339), .A(n7338), .B(n7337), .ZN(n7340)
         );
  INV_X1 U9071 ( .A(n7340), .ZN(n7341) );
  NAND2_X1 U9072 ( .A1(n8364), .A2(n7444), .ZN(n7343) );
  NOR2_X1 U9073 ( .A1(n7344), .A2(n7343), .ZN(n7802) );
  AOI21_X1 U9074 ( .B1(n7344), .B2(n7343), .A(n7802), .ZN(n7476) );
  INV_X1 U9075 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n7345) );
  NAND2_X1 U9076 ( .A1(n7437), .A2(n7345), .ZN(n7346) );
  NAND2_X1 U9077 ( .A1(n7451), .A2(n7346), .ZN(n8391) );
  OR2_X1 U9078 ( .A1(n8391), .A2(n7453), .ZN(n7352) );
  INV_X1 U9079 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n7349) );
  NAND2_X1 U9080 ( .A1(n7244), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n7348) );
  NAND2_X1 U9081 ( .A1(n6802), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n7347) );
  OAI211_X1 U9082 ( .C1(n7349), .C2(n7485), .A(n7348), .B(n7347), .ZN(n7350)
         );
  INV_X1 U9083 ( .A(n7350), .ZN(n7351) );
  NAND2_X1 U9084 ( .A1(n8295), .A2(n7444), .ZN(n7433) );
  INV_X1 U9085 ( .A(n7433), .ZN(n8108) );
  NAND2_X1 U9086 ( .A1(n7353), .A2(n7839), .ZN(n7356) );
  OR2_X1 U9087 ( .A1(n4304), .A2(n7354), .ZN(n7355) );
  XNOR2_X1 U9088 ( .A(n8558), .B(n7798), .ZN(n8109) );
  NAND2_X1 U9089 ( .A1(n7358), .A2(n7357), .ZN(n7359) );
  NAND2_X1 U9090 ( .A1(n7362), .A2(n7839), .ZN(n7364) );
  INV_X1 U9091 ( .A(n8258), .ZN(n8247) );
  AOI22_X1 U9092 ( .A1(n7370), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7369), .B2(
        n8247), .ZN(n7363) );
  XNOR2_X1 U9093 ( .A(n8588), .B(n7798), .ZN(n7365) );
  NOR2_X1 U9094 ( .A1(n8287), .A2(n9913), .ZN(n7366) );
  XNOR2_X1 U9095 ( .A(n7365), .B(n7366), .ZN(n8141) );
  INV_X1 U9096 ( .A(n7365), .ZN(n7367) );
  NAND2_X1 U9097 ( .A1(n7368), .A2(n7839), .ZN(n7372) );
  AOI22_X1 U9098 ( .A1(n7370), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7369), .B2(
        n8530), .ZN(n7371) );
  XNOR2_X1 U9099 ( .A(n8584), .B(n7798), .ZN(n7380) );
  NAND2_X1 U9100 ( .A1(n7832), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n7379) );
  NAND2_X1 U9101 ( .A1(n7374), .A2(n7373), .ZN(n7375) );
  AND2_X1 U9102 ( .A1(n7392), .A2(n7375), .ZN(n8480) );
  NAND2_X1 U9103 ( .A1(n6143), .A2(n8480), .ZN(n7378) );
  NAND2_X1 U9104 ( .A1(n7244), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n7377) );
  NAND2_X1 U9105 ( .A1(n6802), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n7376) );
  OR2_X1 U9106 ( .A1(n8456), .A2(n9913), .ZN(n7381) );
  NAND2_X1 U9107 ( .A1(n7380), .A2(n7381), .ZN(n7385) );
  INV_X1 U9108 ( .A(n7380), .ZN(n7383) );
  INV_X1 U9109 ( .A(n7381), .ZN(n7382) );
  NAND2_X1 U9110 ( .A1(n7383), .A2(n7382), .ZN(n7384) );
  AND2_X1 U9111 ( .A1(n7385), .A2(n7384), .ZN(n8068) );
  NAND2_X1 U9112 ( .A1(n7386), .A2(n7839), .ZN(n7389) );
  OR2_X1 U9113 ( .A1(n4304), .A2(n7387), .ZN(n7388) );
  XNOR2_X1 U9114 ( .A(n8578), .B(n7390), .ZN(n7399) );
  INV_X1 U9115 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7391) );
  NAND2_X1 U9116 ( .A1(n7392), .A2(n7391), .ZN(n7393) );
  AND2_X1 U9117 ( .A1(n7405), .A2(n7393), .ZN(n8451) );
  NAND2_X1 U9118 ( .A1(n8451), .A2(n6143), .ZN(n7397) );
  NAND2_X1 U9119 ( .A1(n7244), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n7396) );
  NAND2_X1 U9120 ( .A1(n6802), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n7395) );
  NAND2_X1 U9121 ( .A1(n7832), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n7394) );
  NOR2_X1 U9122 ( .A1(n8289), .A2(n9913), .ZN(n7398) );
  XNOR2_X1 U9123 ( .A(n7399), .B(n7398), .ZN(n8116) );
  NAND2_X1 U9124 ( .A1(n7400), .A2(n7839), .ZN(n7403) );
  OR2_X1 U9125 ( .A1(n4304), .A2(n7401), .ZN(n7402) );
  XNOR2_X1 U9126 ( .A(n8290), .B(n7798), .ZN(n7414) );
  INV_X1 U9127 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7404) );
  NAND2_X1 U9128 ( .A1(n7405), .A2(n7404), .ZN(n7406) );
  NAND2_X1 U9129 ( .A1(n7421), .A2(n7406), .ZN(n8438) );
  OR2_X1 U9130 ( .A1(n7453), .A2(n8438), .ZN(n7411) );
  NAND2_X1 U9131 ( .A1(n7832), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n7408) );
  NAND2_X1 U9132 ( .A1(n7244), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7407) );
  AND2_X1 U9133 ( .A1(n7408), .A2(n7407), .ZN(n7410) );
  NAND2_X1 U9134 ( .A1(n6802), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7409) );
  NAND2_X1 U9135 ( .A1(n8291), .A2(n7444), .ZN(n7412) );
  XNOR2_X1 U9136 ( .A(n7414), .B(n7412), .ZN(n8075) );
  NAND2_X1 U9137 ( .A1(n8076), .A2(n8075), .ZN(n7416) );
  INV_X1 U9138 ( .A(n7412), .ZN(n7413) );
  NAND2_X1 U9139 ( .A1(n7414), .A2(n7413), .ZN(n7415) );
  NAND2_X1 U9140 ( .A1(n7416), .A2(n7415), .ZN(n7428) );
  NAND2_X1 U9141 ( .A1(n7417), .A2(n7839), .ZN(n7420) );
  OR2_X1 U9142 ( .A1(n4304), .A2(n7418), .ZN(n7419) );
  XNOR2_X1 U9143 ( .A(n8567), .B(n7798), .ZN(n7426) );
  XNOR2_X1 U9144 ( .A(n7428), .B(n7426), .ZN(n8125) );
  NAND2_X1 U9145 ( .A1(n7421), .A2(n8128), .ZN(n7422) );
  NAND2_X1 U9146 ( .A1(n7435), .A2(n7422), .ZN(n8127) );
  OR2_X1 U9147 ( .A1(n8127), .A2(n7453), .ZN(n7425) );
  AOI22_X1 U9148 ( .A1(n7832), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n7244), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n7424) );
  NAND2_X1 U9149 ( .A1(n6802), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n7423) );
  INV_X1 U9150 ( .A(n8293), .ZN(n8176) );
  NAND2_X1 U9151 ( .A1(n8176), .A2(n7444), .ZN(n8124) );
  INV_X1 U9152 ( .A(n7426), .ZN(n7427) );
  OR2_X1 U9153 ( .A1(n7428), .A2(n7427), .ZN(n7429) );
  NAND2_X1 U9154 ( .A1(n7430), .A2(n7839), .ZN(n7432) );
  OR2_X1 U9155 ( .A1(n4304), .A2(n8702), .ZN(n7431) );
  NAND2_X1 U9156 ( .A1(n8109), .A2(n8061), .ZN(n7446) );
  NAND2_X1 U9157 ( .A1(n7435), .A2(n8712), .ZN(n7436) );
  AND2_X1 U9158 ( .A1(n7437), .A2(n7436), .ZN(n8406) );
  NAND2_X1 U9159 ( .A1(n8406), .A2(n6143), .ZN(n7443) );
  INV_X1 U9160 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n7440) );
  NAND2_X1 U9161 ( .A1(n7244), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n7439) );
  NAND2_X1 U9162 ( .A1(n6802), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n7438) );
  OAI211_X1 U9163 ( .C1(n7485), .C2(n7440), .A(n7439), .B(n7438), .ZN(n7441)
         );
  INV_X1 U9164 ( .A(n7441), .ZN(n7442) );
  NAND2_X1 U9165 ( .A1(n7443), .A2(n7442), .ZN(n8174) );
  NAND2_X1 U9166 ( .A1(n8174), .A2(n7444), .ZN(n8106) );
  NAND2_X1 U9167 ( .A1(n8837), .A2(n7839), .ZN(n7449) );
  OR2_X1 U9168 ( .A1(n4304), .A2(n8841), .ZN(n7448) );
  XOR2_X1 U9169 ( .A(n7798), .B(n8554), .Z(n8082) );
  NAND2_X1 U9170 ( .A1(n7460), .A2(n8082), .ZN(n7463) );
  INV_X1 U9171 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n7450) );
  NAND2_X1 U9172 ( .A1(n7451), .A2(n7450), .ZN(n7452) );
  NAND2_X1 U9173 ( .A1(n7467), .A2(n7452), .ZN(n8381) );
  OR2_X1 U9174 ( .A1(n8381), .A2(n7453), .ZN(n7459) );
  INV_X1 U9175 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n7456) );
  NAND2_X1 U9176 ( .A1(n6802), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n7455) );
  NAND2_X1 U9177 ( .A1(n7244), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n7454) );
  OAI211_X1 U9178 ( .C1(n7485), .C2(n7456), .A(n7455), .B(n7454), .ZN(n7457)
         );
  INV_X1 U9179 ( .A(n7457), .ZN(n7458) );
  NOR2_X1 U9180 ( .A1(n8173), .A2(n9913), .ZN(n8081) );
  INV_X1 U9181 ( .A(n8081), .ZN(n7462) );
  INV_X1 U9182 ( .A(n8082), .ZN(n7461) );
  NAND2_X1 U9183 ( .A1(n8833), .A2(n7839), .ZN(n7465) );
  OR2_X1 U9184 ( .A1(n4304), .A2(n8834), .ZN(n7464) );
  XNOR2_X1 U9185 ( .A(n8548), .B(n7798), .ZN(n7474) );
  NAND2_X1 U9186 ( .A1(n7467), .A2(n7466), .ZN(n7468) );
  INV_X1 U9187 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8713) );
  NAND2_X1 U9188 ( .A1(n6802), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n7471) );
  NAND2_X1 U9189 ( .A1(n7244), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7470) );
  OAI211_X1 U9190 ( .C1(n7485), .C2(n8713), .A(n7471), .B(n7470), .ZN(n7472)
         );
  AOI21_X1 U9191 ( .B1(n8358), .B2(n6143), .A(n7472), .ZN(n8344) );
  OR2_X1 U9192 ( .A1(n8344), .A2(n9913), .ZN(n7473) );
  NOR2_X1 U9193 ( .A1(n7474), .A2(n7473), .ZN(n7475) );
  AOI21_X1 U9194 ( .B1(n7474), .B2(n7473), .A(n7475), .ZN(n8152) );
  INV_X1 U9195 ( .A(n7477), .ZN(n8339) );
  NAND2_X1 U9196 ( .A1(n7479), .A2(n7478), .ZN(n7480) );
  NAND2_X1 U9197 ( .A1(n8320), .A2(n6143), .ZN(n7488) );
  INV_X1 U9198 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n7484) );
  NAND2_X1 U9199 ( .A1(n7244), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7483) );
  NAND2_X1 U9200 ( .A1(n6802), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n7482) );
  OAI211_X1 U9201 ( .C1(n7485), .C2(n7484), .A(n7483), .B(n7482), .ZN(n7486)
         );
  INV_X1 U9202 ( .A(n7486), .ZN(n7487) );
  AOI22_X1 U9203 ( .A1(n8300), .A2(n8154), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n7489) );
  OAI21_X1 U9204 ( .B1(n8344), .B2(n8156), .A(n7489), .ZN(n7490) );
  AOI21_X1 U9205 ( .B1(n8339), .B2(n8158), .A(n7490), .ZN(n7491) );
  NOR3_X1 U9206 ( .A1(n7493), .A2(n5532), .A3(n7492), .ZN(n7795) );
  INV_X1 U9207 ( .A(n7791), .ZN(n7494) );
  OAI21_X1 U9208 ( .B1(n5509), .B2(n7494), .A(P1_B_REG_SCAN_IN), .ZN(n7794) );
  INV_X1 U9209 ( .A(n7495), .ZN(n7496) );
  NAND2_X1 U9210 ( .A1(n7496), .A2(SI_30_), .ZN(n7500) );
  NAND2_X1 U9211 ( .A1(n7498), .A2(n7497), .ZN(n7499) );
  NAND2_X1 U9212 ( .A1(n7500), .A2(n7499), .ZN(n7504) );
  MUX2_X1 U9213 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7501), .Z(n7502) );
  XNOR2_X1 U9214 ( .A(n7502), .B(SI_31_), .ZN(n7503) );
  NAND2_X1 U9215 ( .A1(n8818), .A2(n7512), .ZN(n7506) );
  NAND2_X1 U9216 ( .A1(n5407), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7505) );
  INV_X1 U9217 ( .A(n9293), .ZN(n7578) );
  NAND2_X1 U9218 ( .A1(n7507), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n7510) );
  NAND2_X1 U9219 ( .A1(n4960), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n7509) );
  NAND2_X1 U9220 ( .A1(n4884), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n7508) );
  NAND3_X1 U9221 ( .A1(n7510), .A2(n7509), .A3(n7508), .ZN(n9061) );
  INV_X1 U9222 ( .A(n9061), .ZN(n7511) );
  AND2_X1 U9223 ( .A1(n7578), .A2(n7511), .ZN(n7713) );
  NAND2_X1 U9224 ( .A1(n7829), .A2(n7512), .ZN(n7514) );
  NAND2_X1 U9225 ( .A1(n5407), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7513) );
  INV_X1 U9226 ( .A(n9001), .ZN(n7515) );
  NOR2_X1 U9227 ( .A1(n9512), .A2(n7515), .ZN(n7576) );
  NOR2_X1 U9228 ( .A1(n7713), .A2(n7576), .ZN(n7753) );
  AND2_X1 U9229 ( .A1(n9512), .A2(n7515), .ZN(n7751) );
  INV_X1 U9230 ( .A(n7751), .ZN(n7573) );
  NAND2_X1 U9231 ( .A1(n7665), .A2(n7650), .ZN(n7655) );
  OR2_X1 U9232 ( .A1(n7655), .A2(n5525), .ZN(n7542) );
  INV_X1 U9233 ( .A(n7625), .ZN(n7610) );
  OAI21_X1 U9234 ( .B1(n7610), .B2(n7611), .A(n7540), .ZN(n7517) );
  AOI21_X1 U9235 ( .B1(n7517), .B2(n7616), .A(n7516), .ZN(n7519) );
  NAND2_X1 U9236 ( .A1(n7620), .A2(n7518), .ZN(n7617) );
  OAI211_X1 U9237 ( .C1(n7519), .C2(n7617), .A(n7647), .B(n7586), .ZN(n7520)
         );
  AND3_X1 U9238 ( .A1(n7520), .A2(n7646), .A3(n7652), .ZN(n7521) );
  NOR2_X1 U9239 ( .A1(n7542), .A2(n7521), .ZN(n7767) );
  INV_X1 U9240 ( .A(n7767), .ZN(n7552) );
  INV_X1 U9241 ( .A(n7764), .ZN(n7603) );
  INV_X1 U9242 ( .A(n7522), .ZN(n7523) );
  OAI211_X1 U9243 ( .C1(n7525), .C2(n7524), .A(n7752), .B(n7523), .ZN(n7527)
         );
  NAND2_X1 U9244 ( .A1(n7527), .A2(n7526), .ZN(n7529) );
  OAI21_X1 U9245 ( .B1(n7530), .B2(n7529), .A(n7528), .ZN(n7531) );
  NAND2_X1 U9246 ( .A1(n7531), .A2(n7727), .ZN(n7537) );
  AND2_X1 U9247 ( .A1(n5515), .A2(n7532), .ZN(n7533) );
  NAND2_X1 U9248 ( .A1(n7535), .A2(n7533), .ZN(n7760) );
  INV_X1 U9249 ( .A(n7760), .ZN(n7536) );
  INV_X1 U9250 ( .A(n7728), .ZN(n7534) );
  AOI22_X1 U9251 ( .A1(n7537), .A2(n7536), .B1(n7535), .B2(n7534), .ZN(n7544)
         );
  AND2_X1 U9252 ( .A1(n7586), .A2(n7538), .ZN(n7636) );
  AND2_X1 U9253 ( .A1(n7602), .A2(n7624), .ZN(n7539) );
  NAND4_X1 U9254 ( .A1(n7540), .A2(n7647), .A3(n7636), .A4(n7539), .ZN(n7541)
         );
  OR2_X1 U9255 ( .A1(n7542), .A2(n7541), .ZN(n7762) );
  INV_X1 U9256 ( .A(n7762), .ZN(n7543) );
  OAI21_X1 U9257 ( .B1(n7603), .B2(n7544), .A(n7543), .ZN(n7551) );
  OR2_X1 U9258 ( .A1(n7684), .A2(n7545), .ZN(n7546) );
  NAND3_X1 U9259 ( .A1(n7546), .A2(n7694), .A3(n7683), .ZN(n7688) );
  NAND2_X1 U9260 ( .A1(n7672), .A2(n7721), .ZN(n7547) );
  AND2_X1 U9261 ( .A1(n7547), .A2(n7673), .ZN(n7548) );
  AND2_X1 U9262 ( .A1(n7675), .A2(n7548), .ZN(n7679) );
  NAND2_X1 U9263 ( .A1(n7679), .A2(n7664), .ZN(n7549) );
  NOR2_X1 U9264 ( .A1(n7688), .A2(n7549), .ZN(n7765) );
  INV_X1 U9265 ( .A(n7765), .ZN(n7550) );
  AOI21_X1 U9266 ( .B1(n7552), .B2(n7551), .A(n7550), .ZN(n7553) );
  NOR2_X1 U9267 ( .A1(n9092), .A2(n7553), .ZN(n7571) );
  NAND2_X1 U9268 ( .A1(n7706), .A2(n7554), .ZN(n7702) );
  INV_X1 U9269 ( .A(n7699), .ZN(n7555) );
  AND2_X1 U9270 ( .A1(n7770), .A2(n7555), .ZN(n7556) );
  OR2_X1 U9271 ( .A1(n7702), .A2(n7556), .ZN(n7768) );
  AND2_X1 U9272 ( .A1(n7580), .A2(n7705), .ZN(n7569) );
  INV_X1 U9273 ( .A(n7679), .ZN(n7561) );
  INV_X1 U9274 ( .A(n7660), .ZN(n7557) );
  OR2_X1 U9275 ( .A1(n7722), .A2(n7557), .ZN(n7667) );
  INV_X1 U9276 ( .A(n7657), .ZN(n7558) );
  AND3_X1 U9277 ( .A1(n7558), .A2(n7665), .A3(n7664), .ZN(n7559) );
  NOR2_X1 U9278 ( .A1(n7667), .A2(n7559), .ZN(n7560) );
  OAI21_X1 U9279 ( .B1(n7561), .B2(n7560), .A(n7686), .ZN(n7562) );
  OAI21_X1 U9280 ( .B1(n7561), .B2(n7672), .A(n7676), .ZN(n7678) );
  OR2_X1 U9281 ( .A1(n7562), .A2(n7678), .ZN(n7563) );
  NOR2_X1 U9282 ( .A1(n7684), .A2(n7563), .ZN(n7564) );
  NOR2_X1 U9283 ( .A1(n7688), .A2(n7564), .ZN(n7565) );
  NOR2_X1 U9284 ( .A1(n7566), .A2(n7565), .ZN(n7567) );
  OR2_X1 U9285 ( .A1(n7768), .A2(n7567), .ZN(n7568) );
  NAND2_X1 U9286 ( .A1(n7569), .A2(n7568), .ZN(n7773) );
  INV_X1 U9287 ( .A(n7773), .ZN(n7570) );
  OAI21_X1 U9288 ( .B1(n7571), .B2(n7768), .A(n7570), .ZN(n7572) );
  NAND3_X1 U9289 ( .A1(n7573), .A2(n7771), .A3(n7572), .ZN(n7574) );
  AOI21_X1 U9290 ( .B1(n7753), .B2(n7574), .A(n7775), .ZN(n7575) );
  XNOR2_X1 U9291 ( .A(n7575), .B(n9745), .ZN(n7785) );
  INV_X1 U9292 ( .A(n7576), .ZN(n7577) );
  NAND2_X1 U9293 ( .A1(n7577), .A2(n9061), .ZN(n7579) );
  NAND2_X1 U9294 ( .A1(n7579), .A2(n7578), .ZN(n7778) );
  NAND2_X1 U9295 ( .A1(n9061), .A2(n9001), .ZN(n7585) );
  NAND2_X1 U9296 ( .A1(n9512), .A2(n7585), .ZN(n7772) );
  NAND2_X1 U9297 ( .A1(n7617), .A2(n7586), .ZN(n7623) );
  NAND2_X1 U9298 ( .A1(n7588), .A2(n9766), .ZN(n7593) );
  INV_X1 U9299 ( .A(n5515), .ZN(n7589) );
  NAND2_X1 U9300 ( .A1(n7589), .A2(n7588), .ZN(n7591) );
  NAND2_X1 U9301 ( .A1(n7591), .A2(n7590), .ZN(n7730) );
  INV_X1 U9302 ( .A(n7730), .ZN(n7592) );
  OAI21_X1 U9303 ( .B1(n7587), .B2(n7593), .A(n7592), .ZN(n7598) );
  INV_X1 U9304 ( .A(n7601), .ZN(n7597) );
  NAND2_X1 U9305 ( .A1(n7764), .A2(n7757), .ZN(n7596) );
  AOI22_X1 U9306 ( .A1(n7598), .A2(n7597), .B1(n7602), .B2(n7596), .ZN(n7608)
         );
  OR2_X1 U9307 ( .A1(n9746), .A2(n7599), .ZN(n7606) );
  NOR2_X1 U9308 ( .A1(n7601), .A2(n7600), .ZN(n7605) );
  OAI21_X1 U9309 ( .B1(n7603), .B2(n7729), .A(n7602), .ZN(n7604) );
  AOI21_X1 U9310 ( .B1(n7606), .B2(n7605), .A(n7604), .ZN(n7607) );
  OAI211_X1 U9311 ( .C1(n7628), .C2(n7610), .A(n7609), .B(n7624), .ZN(n7612)
         );
  NAND2_X1 U9312 ( .A1(n7612), .A2(n4415), .ZN(n7615) );
  NAND3_X1 U9313 ( .A1(n7615), .A2(n7614), .A3(n7613), .ZN(n7621) );
  NAND2_X1 U9314 ( .A1(n7616), .A2(n7704), .ZN(n7618) );
  NOR2_X1 U9315 ( .A1(n7618), .A2(n7617), .ZN(n7639) );
  INV_X1 U9316 ( .A(n7636), .ZN(n7619) );
  AOI22_X1 U9317 ( .A1(n7621), .A2(n7639), .B1(n7620), .B2(n7619), .ZN(n7622)
         );
  INV_X1 U9318 ( .A(n7624), .ZN(n7627) );
  OAI211_X1 U9319 ( .C1(n7628), .C2(n7627), .A(n7626), .B(n7625), .ZN(n7633)
         );
  INV_X1 U9320 ( .A(n7629), .ZN(n7632) );
  NAND2_X1 U9321 ( .A1(n7630), .A2(n7635), .ZN(n7631) );
  AOI21_X1 U9322 ( .B1(n7633), .B2(n7632), .A(n7631), .ZN(n7634) );
  OAI21_X1 U9323 ( .B1(n7634), .B2(n7704), .A(n7738), .ZN(n7643) );
  INV_X1 U9324 ( .A(n7635), .ZN(n7638) );
  OAI211_X1 U9325 ( .C1(n7638), .C2(n7637), .A(n7636), .B(n7582), .ZN(n7641)
         );
  INV_X1 U9326 ( .A(n7639), .ZN(n7640) );
  NAND2_X1 U9327 ( .A1(n7641), .A2(n7640), .ZN(n7642) );
  NAND2_X1 U9328 ( .A1(n7646), .A2(n7647), .ZN(n9272) );
  AOI21_X1 U9329 ( .B1(n7643), .B2(n7642), .A(n9272), .ZN(n7644) );
  NAND2_X1 U9330 ( .A1(n7645), .A2(n7644), .ZN(n7649) );
  INV_X1 U9331 ( .A(n9256), .ZN(n9253) );
  MUX2_X1 U9332 ( .A(n7647), .B(n7646), .S(n7704), .Z(n7648) );
  NAND3_X1 U9333 ( .A1(n7649), .A2(n9253), .A3(n7648), .ZN(n7654) );
  MUX2_X1 U9334 ( .A(n7652), .B(n7651), .S(n7704), .Z(n7653) );
  NAND3_X1 U9335 ( .A1(n7654), .A2(n9247), .A3(n7653), .ZN(n7659) );
  INV_X1 U9336 ( .A(n7655), .ZN(n7656) );
  MUX2_X1 U9337 ( .A(n7657), .B(n7656), .S(n7582), .Z(n7658) );
  NAND2_X1 U9338 ( .A1(n7659), .A2(n7658), .ZN(n7666) );
  NAND3_X1 U9339 ( .A1(n7666), .A2(n7661), .A3(n7660), .ZN(n7663) );
  INV_X1 U9340 ( .A(n7721), .ZN(n7662) );
  NAND3_X1 U9341 ( .A1(n7663), .A2(n7664), .A3(n7662), .ZN(n7671) );
  NAND3_X1 U9342 ( .A1(n7666), .A2(n7665), .A3(n7664), .ZN(n7669) );
  INV_X1 U9343 ( .A(n7667), .ZN(n7668) );
  NAND2_X1 U9344 ( .A1(n7669), .A2(n7668), .ZN(n7670) );
  INV_X1 U9345 ( .A(n7722), .ZN(n9176) );
  NAND3_X1 U9346 ( .A1(n7680), .A2(n9176), .A3(n7672), .ZN(n7674) );
  NAND2_X1 U9347 ( .A1(n7674), .A2(n7673), .ZN(n7677) );
  INV_X1 U9348 ( .A(n7675), .ZN(n9150) );
  AOI21_X1 U9349 ( .B1(n7677), .B2(n7676), .A(n9150), .ZN(n7682) );
  AOI21_X1 U9350 ( .B1(n7680), .B2(n7679), .A(n7678), .ZN(n7681) );
  MUX2_X1 U9351 ( .A(n7682), .B(n7681), .S(n7704), .Z(n7693) );
  INV_X1 U9352 ( .A(n7683), .ZN(n7687) );
  OR3_X1 U9353 ( .A1(n9149), .A2(n7684), .A3(n7687), .ZN(n7692) );
  INV_X1 U9354 ( .A(n7684), .ZN(n7685) );
  OAI211_X1 U9355 ( .C1(n7687), .C2(n7686), .A(n7685), .B(n9105), .ZN(n7689)
         );
  MUX2_X1 U9356 ( .A(n7689), .B(n7688), .S(n7582), .Z(n7690) );
  INV_X1 U9357 ( .A(n7690), .ZN(n7691) );
  OAI21_X1 U9358 ( .B1(n7693), .B2(n7692), .A(n7691), .ZN(n7696) );
  MUX2_X1 U9359 ( .A(n9105), .B(n7694), .S(n7704), .Z(n7695) );
  NAND2_X1 U9360 ( .A1(n7696), .A2(n7695), .ZN(n7697) );
  XNOR2_X1 U9361 ( .A(n9104), .B(n9122), .ZN(n9098) );
  INV_X1 U9362 ( .A(n9098), .ZN(n9108) );
  NAND2_X1 U9363 ( .A1(n7697), .A2(n9108), .ZN(n7701) );
  MUX2_X1 U9364 ( .A(n7699), .B(n7698), .S(n7582), .Z(n7700) );
  NAND2_X1 U9365 ( .A1(n7705), .A2(n7770), .ZN(n7703) );
  MUX2_X1 U9366 ( .A(n7703), .B(n7702), .S(n7704), .Z(n7708) );
  MUX2_X1 U9367 ( .A(n7706), .B(n7705), .S(n7704), .Z(n7707) );
  OAI21_X1 U9368 ( .B1(n7709), .B2(n7708), .A(n7707), .ZN(n7710) );
  NAND2_X1 U9369 ( .A1(n7710), .A2(n5529), .ZN(n7711) );
  INV_X1 U9370 ( .A(n7775), .ZN(n7787) );
  OAI21_X1 U9371 ( .B1(n7582), .B2(n7772), .A(n7787), .ZN(n7716) );
  INV_X1 U9372 ( .A(n7713), .ZN(n7715) );
  INV_X1 U9373 ( .A(n7778), .ZN(n7714) );
  AOI22_X1 U9374 ( .A1(n7716), .A2(n7715), .B1(n7714), .B2(n7582), .ZN(n7717)
         );
  INV_X1 U9375 ( .A(n7718), .ZN(n7720) );
  NAND3_X1 U9376 ( .A1(n5518), .A2(n7724), .A3(n7723), .ZN(n7725) );
  NOR2_X1 U9377 ( .A1(n7760), .A2(n7725), .ZN(n7735) );
  AND2_X1 U9378 ( .A1(n9714), .A2(n7726), .ZN(n7734) );
  NAND2_X1 U9379 ( .A1(n7728), .A2(n7727), .ZN(n7732) );
  NAND2_X1 U9380 ( .A1(n7730), .A2(n7729), .ZN(n7731) );
  NAND2_X1 U9381 ( .A1(n7732), .A2(n7731), .ZN(n7758) );
  NAND4_X1 U9382 ( .A1(n7735), .A2(n7734), .A3(n7733), .A4(n7758), .ZN(n7737)
         );
  NOR2_X1 U9383 ( .A1(n7737), .A2(n7736), .ZN(n7739) );
  NAND4_X1 U9384 ( .A1(n7739), .A2(n4550), .A3(n9499), .A4(n7738), .ZN(n7741)
         );
  OR3_X1 U9385 ( .A1(n7741), .A2(n9272), .A3(n7740), .ZN(n7742) );
  NOR2_X1 U9386 ( .A1(n7742), .A2(n9256), .ZN(n7743) );
  NAND4_X1 U9387 ( .A1(n9215), .A2(n9247), .A3(n9222), .A4(n7743), .ZN(n7744)
         );
  NOR2_X1 U9388 ( .A1(n9199), .A2(n7744), .ZN(n7745) );
  NAND4_X1 U9389 ( .A1(n7746), .A2(n9166), .A3(n9173), .A4(n7745), .ZN(n7747)
         );
  NOR4_X1 U9390 ( .A1(n9092), .A2(n9129), .A3(n9121), .A4(n7747), .ZN(n7748)
         );
  NAND3_X1 U9391 ( .A1(n9079), .A2(n7748), .A3(n9108), .ZN(n7749) );
  AOI21_X1 U9392 ( .B1(n7754), .B2(n7753), .A(n7752), .ZN(n7780) );
  INV_X1 U9393 ( .A(n7780), .ZN(n7755) );
  OAI21_X1 U9394 ( .B1(n7790), .B2(n7756), .A(n7755), .ZN(n7782) );
  INV_X1 U9395 ( .A(n6683), .ZN(n7761) );
  INV_X1 U9396 ( .A(n7757), .ZN(n7759) );
  OAI22_X1 U9397 ( .A1(n7761), .A2(n7760), .B1(n7759), .B2(n7758), .ZN(n7763)
         );
  AOI21_X1 U9398 ( .B1(n7764), .B2(n7763), .A(n7762), .ZN(n7766) );
  OAI21_X1 U9399 ( .B1(n7767), .B2(n7766), .A(n7765), .ZN(n7769) );
  AOI21_X1 U9400 ( .B1(n7770), .B2(n7769), .A(n7768), .ZN(n7774) );
  OAI211_X1 U9401 ( .C1(n7774), .C2(n7773), .A(n7772), .B(n7771), .ZN(n7777)
         );
  AOI211_X1 U9402 ( .C1(n7778), .C2(n7777), .A(n7776), .B(n7775), .ZN(n7779)
         );
  NOR2_X1 U9403 ( .A1(n7780), .A2(n7779), .ZN(n7781) );
  MUX2_X1 U9404 ( .A(n7782), .B(n7781), .S(n9136), .Z(n7784) );
  INV_X1 U9405 ( .A(n7786), .ZN(n7789) );
  AND4_X1 U9406 ( .A1(n7790), .A2(n7789), .A3(n7788), .A4(n7787), .ZN(n7792)
         );
  OAI21_X1 U9407 ( .B1(n7795), .B2(n7794), .A(n7793), .ZN(P1_U3240) );
  NAND2_X1 U9408 ( .A1(n8039), .A2(n7839), .ZN(n7797) );
  OR2_X1 U9409 ( .A1(n4304), .A2(n8040), .ZN(n7796) );
  NOR2_X1 U9410 ( .A1(n8345), .A2(n9913), .ZN(n7799) );
  XNOR2_X1 U9411 ( .A(n7799), .B(n7798), .ZN(n7800) );
  XNOR2_X1 U9412 ( .A(n8537), .B(n7800), .ZN(n7806) );
  INV_X1 U9413 ( .A(n7806), .ZN(n7801) );
  NAND2_X1 U9414 ( .A1(n7801), .A2(n8150), .ZN(n7812) );
  INV_X1 U9415 ( .A(n7802), .ZN(n7805) );
  NAND4_X1 U9416 ( .A1(n7811), .A2(n8150), .A3(n7806), .A4(n7805), .ZN(n7810)
         );
  AOI22_X1 U9417 ( .A1(n8364), .A2(n8143), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n7804) );
  NAND2_X1 U9418 ( .A1(n8158), .A2(n8320), .ZN(n7803) );
  OAI211_X1 U9419 ( .C1(n8326), .C2(n8145), .A(n7804), .B(n7803), .ZN(n7808)
         );
  NOR3_X1 U9420 ( .A1(n7806), .A2(n7805), .A3(n9882), .ZN(n7807) );
  AOI211_X1 U9421 ( .C1(n9886), .C2(n8537), .A(n7808), .B(n7807), .ZN(n7809)
         );
  OAI211_X1 U9422 ( .C1(n7812), .C2(n7811), .A(n7810), .B(n7809), .ZN(P2_U3222) );
  NAND2_X1 U9423 ( .A1(n8558), .A2(n8061), .ZN(n7952) );
  INV_X1 U9424 ( .A(n7921), .ZN(n7912) );
  OR2_X1 U9425 ( .A1(n8610), .A2(n8177), .ZN(n7925) );
  NAND2_X1 U9426 ( .A1(n8610), .A2(n8177), .ZN(n8509) );
  NAND2_X1 U9427 ( .A1(n7814), .A2(n8599), .ZN(n8508) );
  NAND2_X1 U9428 ( .A1(n8594), .A2(n8098), .ZN(n7927) );
  NAND2_X1 U9429 ( .A1(n7929), .A2(n7927), .ZN(n8514) );
  INV_X1 U9430 ( .A(n8509), .ZN(n7815) );
  NOR2_X1 U9431 ( .A1(n8514), .A2(n7815), .ZN(n7816) );
  INV_X1 U9432 ( .A(n7989), .ZN(n8468) );
  INV_X1 U9433 ( .A(n7988), .ZN(n7819) );
  OR2_X1 U9434 ( .A1(n8468), .A2(n7819), .ZN(n7817) );
  NAND2_X1 U9435 ( .A1(n8588), .A2(n8287), .ZN(n8469) );
  NAND2_X1 U9436 ( .A1(n8584), .A2(n8456), .ZN(n7987) );
  AND2_X1 U9437 ( .A1(n8469), .A2(n7987), .ZN(n7818) );
  OR2_X1 U9438 ( .A1(n7819), .A2(n7818), .ZN(n7820) );
  NAND2_X1 U9439 ( .A1(n8578), .A2(n8289), .ZN(n7985) );
  INV_X1 U9440 ( .A(n7985), .ZN(n7821) );
  XNOR2_X1 U9441 ( .A(n8573), .B(n8458), .ZN(n8433) );
  NAND2_X1 U9442 ( .A1(n8573), .A2(n8458), .ZN(n7940) );
  NAND2_X1 U9443 ( .A1(n8567), .A2(n8293), .ZN(n7941) );
  NAND2_X1 U9444 ( .A1(n8409), .A2(n7941), .ZN(n8423) );
  NAND2_X1 U9445 ( .A1(n8408), .A2(n8174), .ZN(n7946) );
  INV_X1 U9446 ( .A(n8174), .ZN(n8294) );
  NAND2_X1 U9447 ( .A1(n8562), .A2(n8294), .ZN(n7945) );
  NAND2_X1 U9448 ( .A1(n7946), .A2(n7945), .ZN(n8410) );
  INV_X1 U9449 ( .A(n8409), .ZN(n7822) );
  NOR2_X1 U9450 ( .A1(n8410), .A2(n7822), .ZN(n7823) );
  NAND2_X2 U9451 ( .A1(n8296), .A2(n7824), .ZN(n8397) );
  NAND2_X1 U9452 ( .A1(n8554), .A2(n8173), .ZN(n7949) );
  NAND2_X1 U9453 ( .A1(n7951), .A2(n7949), .ZN(n8371) );
  INV_X1 U9454 ( .A(n8371), .ZN(n8375) );
  OR2_X1 U9455 ( .A1(n8548), .A2(n8344), .ZN(n7954) );
  NAND2_X1 U9456 ( .A1(n8548), .A2(n8344), .ZN(n7955) );
  NAND2_X1 U9457 ( .A1(n7954), .A2(n7955), .ZN(n8353) );
  INV_X1 U9458 ( .A(n8353), .ZN(n8363) );
  NAND2_X1 U9459 ( .A1(n8542), .A2(n8325), .ZN(n7958) );
  NAND2_X1 U9460 ( .A1(n8537), .A2(n8345), .ZN(n7959) );
  INV_X1 U9461 ( .A(n8323), .ZN(n8015) );
  NAND2_X1 U9462 ( .A1(n8322), .A2(n8015), .ZN(n8328) );
  NAND2_X1 U9463 ( .A1(n8828), .A2(n7839), .ZN(n7827) );
  OR2_X1 U9464 ( .A1(n4304), .A2(n8830), .ZN(n7826) );
  OR2_X1 U9465 ( .A1(n8308), .A2(n8326), .ZN(n7967) );
  INV_X1 U9466 ( .A(n7967), .ZN(n7828) );
  NAND2_X1 U9467 ( .A1(n8308), .A2(n8326), .ZN(n7968) );
  OAI21_X1 U9468 ( .B1(n8303), .B2(n7828), .A(n7968), .ZN(n7838) );
  NAND2_X1 U9469 ( .A1(n7829), .A2(n7839), .ZN(n7831) );
  INV_X1 U9470 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8826) );
  OR2_X1 U9471 ( .A1(n4304), .A2(n8826), .ZN(n7830) );
  OR2_X1 U9472 ( .A1(n8276), .A2(n8305), .ZN(n7973) );
  NAND2_X1 U9473 ( .A1(n7832), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7835) );
  NAND2_X1 U9474 ( .A1(n6802), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7834) );
  NAND2_X1 U9475 ( .A1(n7244), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7833) );
  NAND3_X1 U9476 ( .A1(n7835), .A2(n7834), .A3(n7833), .ZN(n8172) );
  NAND2_X1 U9477 ( .A1(n8818), .A2(n7839), .ZN(n7841) );
  INV_X1 U9478 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8820) );
  OR2_X1 U9479 ( .A1(n4304), .A2(n8820), .ZN(n7840) );
  NAND2_X1 U9480 ( .A1(n8276), .A2(n8305), .ZN(n7971) );
  NAND2_X1 U9481 ( .A1(n8522), .A2(n8272), .ZN(n7974) );
  NAND2_X1 U9482 ( .A1(n7842), .A2(n7974), .ZN(n7844) );
  INV_X1 U9483 ( .A(n7845), .ZN(n7843) );
  AND2_X1 U9484 ( .A1(n7844), .A2(n7843), .ZN(n7847) );
  AOI21_X1 U9485 ( .B1(n7845), .B2(n9996), .A(n7844), .ZN(n7846) );
  MUX2_X2 U9486 ( .A(n7847), .B(n7846), .S(n8481), .Z(n8025) );
  INV_X1 U9487 ( .A(n7975), .ZN(n7978) );
  AND2_X1 U9488 ( .A1(n7859), .A2(n8020), .ZN(n7849) );
  OAI21_X1 U9489 ( .B1(n7850), .B2(n7849), .A(n7860), .ZN(n7851) );
  NAND2_X1 U9490 ( .A1(n7851), .A2(n7863), .ZN(n7852) );
  NAND2_X1 U9491 ( .A1(n7852), .A2(n7864), .ZN(n7853) );
  AND2_X1 U9492 ( .A1(n7858), .A2(n7854), .ZN(n7855) );
  MUX2_X1 U9493 ( .A(n7855), .B(n4316), .S(n7975), .Z(n7872) );
  NAND2_X1 U9494 ( .A1(n7860), .A2(n7859), .ZN(n7861) );
  NAND3_X1 U9495 ( .A1(n7863), .A2(n7862), .A3(n7861), .ZN(n7865) );
  NAND2_X1 U9496 ( .A1(n7865), .A2(n7864), .ZN(n7866) );
  INV_X1 U9497 ( .A(n7873), .ZN(n7867) );
  INV_X1 U9498 ( .A(n7868), .ZN(n7871) );
  NAND2_X1 U9499 ( .A1(n4316), .A2(n7869), .ZN(n7870) );
  OAI21_X1 U9500 ( .B1(n7872), .B2(n7871), .A(n7870), .ZN(n7874) );
  AOI21_X1 U9501 ( .B1(n7874), .B2(n7873), .A(n7975), .ZN(n7878) );
  NOR2_X1 U9502 ( .A1(n7875), .A2(n7975), .ZN(n7876) );
  NOR2_X1 U9503 ( .A1(n7876), .A2(n7997), .ZN(n7877) );
  OAI21_X1 U9504 ( .B1(n7879), .B2(n7878), .A(n7877), .ZN(n7883) );
  MUX2_X1 U9505 ( .A(n7881), .B(n7880), .S(n7975), .Z(n7882) );
  MUX2_X1 U9506 ( .A(n7885), .B(n7884), .S(n7978), .Z(n7886) );
  NAND2_X1 U9507 ( .A1(n7892), .A2(n7893), .ZN(n7889) );
  INV_X1 U9508 ( .A(n7887), .ZN(n7888) );
  MUX2_X1 U9509 ( .A(n7889), .B(n7888), .S(n7975), .Z(n7890) );
  INV_X1 U9510 ( .A(n7890), .ZN(n7891) );
  INV_X1 U9511 ( .A(n7894), .ZN(n7897) );
  NAND2_X1 U9512 ( .A1(n7898), .A2(n7895), .ZN(n7896) );
  NAND2_X1 U9513 ( .A1(n7903), .A2(n7898), .ZN(n7901) );
  NAND2_X1 U9514 ( .A1(n7902), .A2(n7899), .ZN(n7900) );
  MUX2_X1 U9515 ( .A(n7901), .B(n7900), .S(n7978), .Z(n7905) );
  MUX2_X1 U9516 ( .A(n7903), .B(n7902), .S(n7975), .Z(n7904) );
  OAI211_X1 U9517 ( .C1(n7906), .C2(n7905), .A(n8003), .B(n7904), .ZN(n7910)
         );
  MUX2_X1 U9518 ( .A(n7908), .B(n7907), .S(n7975), .Z(n7909) );
  NAND2_X1 U9519 ( .A1(n7910), .A2(n7909), .ZN(n7918) );
  MUX2_X1 U9520 ( .A(n7911), .B(n9465), .S(n7978), .Z(n7917) );
  AOI21_X1 U9521 ( .B1(n7914), .B2(n8178), .A(n7912), .ZN(n7916) );
  AOI21_X1 U9522 ( .B1(n7914), .B2(n7913), .A(n4582), .ZN(n7915) );
  MUX2_X1 U9523 ( .A(n7916), .B(n7915), .S(n7975), .Z(n7920) );
  NAND2_X1 U9524 ( .A1(n7918), .A2(n7917), .ZN(n7919) );
  NAND2_X1 U9525 ( .A1(n7920), .A2(n7919), .ZN(n7924) );
  MUX2_X1 U9526 ( .A(n7921), .B(n8600), .S(n7978), .Z(n7922) );
  AND2_X1 U9527 ( .A1(n7922), .A2(n8599), .ZN(n7923) );
  NAND2_X1 U9528 ( .A1(n7924), .A2(n7923), .ZN(n7928) );
  NAND3_X1 U9529 ( .A1(n7928), .A2(n7925), .A3(n7929), .ZN(n7926) );
  NAND3_X1 U9530 ( .A1(n7928), .A2(n8509), .A3(n7927), .ZN(n7930) );
  NAND2_X1 U9531 ( .A1(n7934), .A2(n8469), .ZN(n7931) );
  NAND2_X1 U9532 ( .A1(n7931), .A2(n7988), .ZN(n7932) );
  NAND3_X1 U9533 ( .A1(n7932), .A2(n7987), .A3(n7985), .ZN(n7933) );
  NAND2_X1 U9534 ( .A1(n8290), .A2(n8291), .ZN(n7937) );
  NAND3_X1 U9535 ( .A1(n7935), .A2(n7988), .A3(n7986), .ZN(n7936) );
  NAND2_X1 U9536 ( .A1(n8409), .A2(n7937), .ZN(n7938) );
  NAND2_X1 U9537 ( .A1(n7938), .A2(n7978), .ZN(n7939) );
  AOI21_X1 U9538 ( .B1(n7941), .B2(n7940), .A(n7978), .ZN(n7944) );
  NOR2_X1 U9539 ( .A1(n8409), .A2(n7978), .ZN(n7942) );
  NOR2_X1 U9540 ( .A1(n8410), .A2(n7942), .ZN(n7943) );
  NAND2_X1 U9541 ( .A1(n7947), .A2(n7946), .ZN(n7948) );
  NAND2_X1 U9542 ( .A1(n7955), .A2(n7949), .ZN(n7950) );
  INV_X1 U9543 ( .A(n8342), .ZN(n8014) );
  MUX2_X1 U9544 ( .A(n7955), .B(n7954), .S(n7975), .Z(n7956) );
  NAND2_X1 U9545 ( .A1(n7959), .A2(n7958), .ZN(n7960) );
  MUX2_X1 U9546 ( .A(n4782), .B(n7960), .S(n7975), .Z(n7963) );
  INV_X1 U9547 ( .A(n7961), .ZN(n7962) );
  NOR2_X1 U9548 ( .A1(n7963), .A2(n7962), .ZN(n7966) );
  NAND2_X1 U9549 ( .A1(n8537), .A2(n8300), .ZN(n7965) );
  MUX2_X1 U9550 ( .A(n8300), .B(n8537), .S(n7978), .Z(n7964) );
  NAND2_X1 U9551 ( .A1(n7967), .A2(n7968), .ZN(n8304) );
  MUX2_X1 U9552 ( .A(n7968), .B(n7967), .S(n7975), .Z(n7969) );
  OAI21_X1 U9553 ( .B1(n7970), .B2(n8304), .A(n7969), .ZN(n7972) );
  NAND3_X1 U9554 ( .A1(n7972), .A2(n7973), .A3(n7971), .ZN(n7977) );
  AND2_X1 U9555 ( .A1(n7974), .A2(n7973), .ZN(n7983) );
  MUX2_X1 U9556 ( .A(n7984), .B(n7983), .S(n7975), .Z(n7976) );
  NAND2_X1 U9557 ( .A1(n7977), .A2(n7976), .ZN(n7981) );
  INV_X1 U9558 ( .A(n8522), .ZN(n8273) );
  MUX2_X1 U9559 ( .A(n8172), .B(n8522), .S(n7978), .Z(n7979) );
  OAI21_X1 U9560 ( .B1(n8273), .B2(n8272), .A(n7979), .ZN(n7980) );
  NAND2_X1 U9561 ( .A1(n7981), .A2(n7980), .ZN(n8024) );
  INV_X1 U9562 ( .A(n8022), .ZN(n7982) );
  INV_X1 U9563 ( .A(n7983), .ZN(n8018) );
  INV_X1 U9564 ( .A(n8423), .ZN(n8417) );
  NAND2_X1 U9565 ( .A1(n7986), .A2(n7985), .ZN(n8448) );
  NAND2_X1 U9566 ( .A1(n7988), .A2(n7987), .ZN(n8466) );
  NAND2_X1 U9567 ( .A1(n7989), .A2(n8469), .ZN(n8489) );
  NOR4_X1 U9568 ( .A1(n6396), .A2(n7990), .A3(n9915), .A4(n6109), .ZN(n7994)
         );
  INV_X1 U9569 ( .A(n7991), .ZN(n7993) );
  NAND3_X1 U9570 ( .A1(n7994), .A2(n7993), .A3(n7992), .ZN(n7998) );
  NOR4_X1 U9571 ( .A1(n7998), .A2(n7997), .A3(n7996), .A4(n7995), .ZN(n8002)
         );
  NAND4_X1 U9572 ( .A1(n8002), .A2(n8001), .A3(n8000), .A4(n7999), .ZN(n8007)
         );
  INV_X1 U9573 ( .A(n8003), .ZN(n8006) );
  NOR4_X1 U9574 ( .A1(n8007), .A2(n8006), .A3(n8005), .A4(n8004), .ZN(n8009)
         );
  NAND4_X1 U9575 ( .A1(n8599), .A2(n8282), .A3(n8009), .A4(n8008), .ZN(n8010)
         );
  NOR4_X1 U9576 ( .A1(n8466), .A2(n8489), .A3(n8514), .A4(n8010), .ZN(n8011)
         );
  NAND4_X1 U9577 ( .A1(n4450), .A2(n8417), .A3(n4680), .A4(n8011), .ZN(n8012)
         );
  NOR4_X1 U9578 ( .A1(n8371), .A2(n8394), .A3(n8433), .A4(n8012), .ZN(n8013)
         );
  NAND4_X1 U9579 ( .A1(n8015), .A2(n8014), .A3(n8363), .A4(n8013), .ZN(n8016)
         );
  NOR4_X1 U9580 ( .A1(n8018), .A2(n8017), .A3(n8304), .A4(n8016), .ZN(n8019)
         );
  XNOR2_X1 U9581 ( .A(n8019), .B(n8530), .ZN(n8021) );
  NOR3_X1 U9582 ( .A1(n8026), .A2(n6264), .A3(n8455), .ZN(n8029) );
  OAI21_X1 U9583 ( .B1(n8030), .B2(n8027), .A(P2_B_REG_SCAN_IN), .ZN(n8028) );
  OAI22_X1 U9584 ( .A1(n8031), .A2(n8030), .B1(n8029), .B2(n8028), .ZN(
        P2_U3244) );
  AOI22_X1 U9585 ( .A1(n8154), .A2(n8191), .B1(n9886), .B2(n9920), .ZN(n8037)
         );
  OAI21_X1 U9586 ( .B1(n8034), .B2(n8033), .A(n8032), .ZN(n8035) );
  AOI22_X1 U9587 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(n8133), .B1(n8150), .B2(
        n8035), .ZN(n8036) );
  OAI211_X1 U9588 ( .C1(n8038), .C2(n8156), .A(n8037), .B(n8036), .ZN(P2_U3224) );
  INV_X1 U9589 ( .A(n8039), .ZN(n9389) );
  OAI222_X1 U9590 ( .A1(n8827), .A2(n8040), .B1(n8840), .B2(n9389), .C1(n6052), 
        .C2(P2_U3152), .ZN(P2_U3330) );
  NAND2_X1 U9591 ( .A1(n9302), .A2(n4310), .ZN(n8042) );
  NAND2_X1 U9592 ( .A1(n9002), .A2(n4308), .ZN(n8041) );
  NAND2_X1 U9593 ( .A1(n8042), .A2(n8041), .ZN(n8044) );
  XNOR2_X1 U9594 ( .A(n8044), .B(n8043), .ZN(n8047) );
  AOI22_X1 U9595 ( .A1(n9302), .A2(n5625), .B1(n8045), .B2(n9002), .ZN(n8046)
         );
  XNOR2_X1 U9596 ( .A(n8047), .B(n8046), .ZN(n8048) );
  INV_X1 U9597 ( .A(n8048), .ZN(n8054) );
  NAND3_X1 U9598 ( .A1(n8054), .A2(n8977), .A3(n8053), .ZN(n8059) );
  NAND2_X1 U9599 ( .A1(n8060), .A2(n8049), .ZN(n8058) );
  INV_X1 U9600 ( .A(n8050), .ZN(n9080) );
  AOI22_X1 U9601 ( .A1(n9080), .A2(n8992), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8052) );
  NAND2_X1 U9602 ( .A1(n8997), .A2(n9075), .ZN(n8051) );
  OAI211_X1 U9603 ( .C1(n9003), .C2(n8994), .A(n8052), .B(n8051), .ZN(n8056)
         );
  NOR3_X1 U9604 ( .A1(n8054), .A2(n8988), .A3(n8053), .ZN(n8055) );
  AOI211_X1 U9605 ( .C1(n9302), .C2(n8965), .A(n8056), .B(n8055), .ZN(n8057)
         );
  OAI211_X1 U9606 ( .C1(n8060), .C2(n8059), .A(n8058), .B(n8057), .ZN(P1_U3218) );
  XNOR2_X1 U9607 ( .A(n8107), .B(n8106), .ZN(n8066) );
  INV_X1 U9608 ( .A(n8406), .ZN(n8063) );
  OAI22_X1 U9609 ( .A1(n8061), .A2(n8457), .B1(n8293), .B2(n8455), .ZN(n8412)
         );
  AOI22_X1 U9610 ( .A1(n9881), .A2(n8412), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8062) );
  OAI21_X1 U9611 ( .B1(n8063), .B2(n9891), .A(n8062), .ZN(n8064) );
  AOI21_X1 U9612 ( .B1(n8562), .B2(n9886), .A(n8064), .ZN(n8065) );
  OAI21_X1 U9613 ( .B1(n8066), .B2(n9882), .A(n8065), .ZN(P2_U3218) );
  OAI21_X1 U9614 ( .B1(n8069), .B2(n8068), .A(n8067), .ZN(n8070) );
  NAND2_X1 U9615 ( .A1(n8070), .A2(n8150), .ZN(n8074) );
  INV_X1 U9616 ( .A(n8289), .ZN(n8474) );
  NAND2_X1 U9617 ( .A1(n8154), .A2(n8474), .ZN(n8071) );
  NAND2_X1 U9618 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8266) );
  OAI211_X1 U9619 ( .C1(n8287), .C2(n8156), .A(n8071), .B(n8266), .ZN(n8072)
         );
  AOI21_X1 U9620 ( .B1(n8480), .B2(n8158), .A(n8072), .ZN(n8073) );
  OAI211_X1 U9621 ( .C1(n8288), .C2(n8161), .A(n8074), .B(n8073), .ZN(P2_U3221) );
  XNOR2_X1 U9622 ( .A(n8076), .B(n8075), .ZN(n8080) );
  OAI22_X1 U9623 ( .A1(n8293), .A2(n8457), .B1(n8289), .B2(n8455), .ZN(n8435)
         );
  AOI22_X1 U9624 ( .A1(n9881), .A2(n8435), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8077) );
  OAI21_X1 U9625 ( .B1(n8438), .B2(n9891), .A(n8077), .ZN(n8078) );
  AOI21_X1 U9626 ( .B1(n8573), .B2(n9886), .A(n8078), .ZN(n8079) );
  OAI21_X1 U9627 ( .B1(n8080), .B2(n9882), .A(n8079), .ZN(P2_U3225) );
  XNOR2_X1 U9628 ( .A(n8082), .B(n8081), .ZN(n8083) );
  XNOR2_X1 U9629 ( .A(n8084), .B(n8083), .ZN(n8090) );
  OR2_X1 U9630 ( .A1(n8344), .A2(n8457), .ZN(n8086) );
  NAND2_X1 U9631 ( .A1(n8295), .A2(n8605), .ZN(n8085) );
  NAND2_X1 U9632 ( .A1(n8086), .A2(n8085), .ZN(n8377) );
  AOI22_X1 U9633 ( .A1(n8377), .A2(n9881), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8087) );
  OAI21_X1 U9634 ( .B1(n8381), .B2(n9891), .A(n8087), .ZN(n8088) );
  AOI21_X1 U9635 ( .B1(n8554), .B2(n9886), .A(n8088), .ZN(n8089) );
  OAI21_X1 U9636 ( .B1(n8090), .B2(n9882), .A(n8089), .ZN(P2_U3227) );
  INV_X1 U9637 ( .A(n8610), .ZN(n9439) );
  NAND2_X1 U9638 ( .A1(n4390), .A2(n8091), .ZN(n8092) );
  OAI21_X1 U9639 ( .B1(n4390), .B2(n8091), .A(n8092), .ZN(n8163) );
  NOR2_X1 U9640 ( .A1(n8163), .A2(n8164), .ZN(n8162) );
  INV_X1 U9641 ( .A(n8092), .ZN(n8093) );
  NOR3_X1 U9642 ( .A1(n8162), .A2(n8094), .A3(n8093), .ZN(n8097) );
  INV_X1 U9643 ( .A(n8095), .ZN(n8096) );
  OAI21_X1 U9644 ( .B1(n8097), .B2(n8096), .A(n8150), .ZN(n8104) );
  NAND2_X1 U9645 ( .A1(n8154), .A2(n8604), .ZN(n8100) );
  OAI211_X1 U9646 ( .C1(n8101), .C2(n8156), .A(n8100), .B(n8099), .ZN(n8102)
         );
  AOI21_X1 U9647 ( .B1(n9436), .B2(n8158), .A(n8102), .ZN(n8103) );
  OAI211_X1 U9648 ( .C1(n9439), .C2(n8161), .A(n8104), .B(n8103), .ZN(P2_U3228) );
  OAI21_X1 U9649 ( .B1(n8107), .B2(n8106), .A(n8105), .ZN(n8111) );
  XNOR2_X1 U9650 ( .A(n8109), .B(n8108), .ZN(n8110) );
  XNOR2_X1 U9651 ( .A(n8111), .B(n8110), .ZN(n8115) );
  OAI22_X1 U9652 ( .A1(n8173), .A2(n8457), .B1(n8294), .B2(n8455), .ZN(n8396)
         );
  AOI22_X1 U9653 ( .A1(n8396), .A2(n9881), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n8112) );
  OAI21_X1 U9654 ( .B1(n8391), .B2(n9891), .A(n8112), .ZN(n8113) );
  AOI21_X1 U9655 ( .B1(n8558), .B2(n9886), .A(n8113), .ZN(n8114) );
  OAI21_X1 U9656 ( .B1(n8115), .B2(n9882), .A(n8114), .ZN(P2_U3231) );
  XNOR2_X1 U9657 ( .A(n8117), .B(n8116), .ZN(n8122) );
  AOI22_X1 U9658 ( .A1(n8154), .A2(n8291), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8119) );
  NAND2_X1 U9659 ( .A1(n8158), .A2(n8451), .ZN(n8118) );
  OAI211_X1 U9660 ( .C1(n8456), .C2(n8156), .A(n8119), .B(n8118), .ZN(n8120)
         );
  AOI21_X1 U9661 ( .B1(n8578), .B2(n9886), .A(n8120), .ZN(n8121) );
  OAI21_X1 U9662 ( .B1(n8122), .B2(n9882), .A(n8121), .ZN(P2_U3235) );
  INV_X1 U9663 ( .A(n8567), .ZN(n8422) );
  OAI21_X1 U9664 ( .B1(n8125), .B2(n8124), .A(n8123), .ZN(n8126) );
  NAND2_X1 U9665 ( .A1(n8126), .A2(n8150), .ZN(n8132) );
  INV_X1 U9666 ( .A(n8127), .ZN(n8420) );
  AOI22_X1 U9667 ( .A1(n8174), .A2(n8603), .B1(n8291), .B2(n8605), .ZN(n8425)
         );
  OAI22_X1 U9668 ( .A1(n8129), .A2(n8425), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8128), .ZN(n8130) );
  AOI21_X1 U9669 ( .B1(n8158), .B2(n8420), .A(n8130), .ZN(n8131) );
  OAI211_X1 U9670 ( .C1(n8422), .C2(n8161), .A(n8132), .B(n8131), .ZN(P2_U3237) );
  AOI22_X1 U9671 ( .A1(n8154), .A2(n8190), .B1(n8143), .B2(n6387), .ZN(n8140)
         );
  AOI22_X1 U9672 ( .A1(n9886), .A2(n9929), .B1(n8133), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n8139) );
  OAI21_X1 U9673 ( .B1(n8136), .B2(n8135), .A(n8134), .ZN(n8137) );
  NAND2_X1 U9674 ( .A1(n8137), .A2(n8150), .ZN(n8138) );
  NAND3_X1 U9675 ( .A1(n8140), .A2(n8139), .A3(n8138), .ZN(P2_U3239) );
  XNOR2_X1 U9676 ( .A(n8142), .B(n8141), .ZN(n8149) );
  NAND2_X1 U9677 ( .A1(n8143), .A2(n8604), .ZN(n8144) );
  NAND2_X1 U9678 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8245) );
  OAI211_X1 U9679 ( .C1(n8456), .C2(n8145), .A(n8144), .B(n8245), .ZN(n8147)
         );
  NOR2_X1 U9680 ( .A1(n8498), .A2(n8161), .ZN(n8146) );
  AOI211_X1 U9681 ( .C1(n8158), .C2(n8495), .A(n8147), .B(n8146), .ZN(n8148)
         );
  OAI21_X1 U9682 ( .B1(n8149), .B2(n9882), .A(n8148), .ZN(P2_U3240) );
  INV_X1 U9683 ( .A(n8548), .ZN(n8360) );
  OAI211_X1 U9684 ( .C1(n8153), .C2(n8152), .A(n8151), .B(n8150), .ZN(n8160)
         );
  AOI22_X1 U9685 ( .A1(n8364), .A2(n8154), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8155) );
  OAI21_X1 U9686 ( .B1(n8173), .B2(n8156), .A(n8155), .ZN(n8157) );
  AOI21_X1 U9687 ( .B1(n8358), .B2(n8158), .A(n8157), .ZN(n8159) );
  OAI211_X1 U9688 ( .C1(n8360), .C2(n8161), .A(n8160), .B(n8159), .ZN(P2_U3242) );
  AOI21_X1 U9689 ( .B1(n8164), .B2(n8163), .A(n8162), .ZN(n8171) );
  INV_X1 U9690 ( .A(n8165), .ZN(n8168) );
  AND2_X1 U9691 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8209) );
  AOI21_X1 U9692 ( .B1(n9881), .B2(n8166), .A(n8209), .ZN(n8167) );
  OAI21_X1 U9693 ( .B1(n9891), .B2(n8168), .A(n8167), .ZN(n8169) );
  AOI21_X1 U9694 ( .B1(n8280), .B2(n9886), .A(n8169), .ZN(n8170) );
  OAI21_X1 U9695 ( .B1(n8171), .B2(n9882), .A(n8170), .ZN(P2_U3243) );
  MUX2_X1 U9696 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8172), .S(P2_U3966), .Z(
        P2_U3583) );
  MUX2_X1 U9697 ( .A(n8300), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8175), .Z(
        P2_U3580) );
  MUX2_X1 U9698 ( .A(n8364), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8175), .Z(
        P2_U3579) );
  INV_X1 U9699 ( .A(n8344), .ZN(n8297) );
  MUX2_X1 U9700 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8297), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U9701 ( .A(n8365), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8175), .Z(
        P2_U3577) );
  MUX2_X1 U9702 ( .A(n8295), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8175), .Z(
        P2_U3576) );
  MUX2_X1 U9703 ( .A(n8174), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8175), .Z(
        P2_U3575) );
  MUX2_X1 U9704 ( .A(n8176), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8175), .Z(
        P2_U3574) );
  MUX2_X1 U9705 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8291), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9706 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8474), .S(P2_U3966), .Z(
        P2_U3572) );
  INV_X1 U9707 ( .A(n8456), .ZN(n8490) );
  MUX2_X1 U9708 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8490), .S(P2_U3966), .Z(
        P2_U3571) );
  INV_X1 U9709 ( .A(n8287), .ZN(n8475) );
  MUX2_X1 U9710 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8475), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9711 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8604), .S(P2_U3966), .Z(
        P2_U3569) );
  INV_X1 U9712 ( .A(n8177), .ZN(n8284) );
  MUX2_X1 U9713 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8284), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9714 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8606), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9715 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8178), .S(P2_U3966), .Z(
        P2_U3566) );
  INV_X1 U9716 ( .A(n8179), .ZN(n8180) );
  MUX2_X1 U9717 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8180), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9718 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8181), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9719 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8182), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9720 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8183), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9721 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8184), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9722 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8185), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9723 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8186), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9724 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8187), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9725 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8188), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9726 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8189), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9727 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8190), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U9728 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8191), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U9729 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6387), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U9730 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8192), .S(P2_U3966), .Z(
        P2_U3552) );
  OAI21_X1 U9731 ( .B1(n8195), .B2(n8194), .A(n8193), .ZN(n8196) );
  NAND2_X1 U9732 ( .A1(n9897), .A2(n8196), .ZN(n8206) );
  NOR2_X1 U9733 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8197), .ZN(n8198) );
  AOI21_X1 U9734 ( .B1(n9898), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8198), .ZN(
        n8205) );
  NAND2_X1 U9735 ( .A1(n9895), .A2(n8199), .ZN(n8204) );
  OAI211_X1 U9736 ( .C1(n8202), .C2(n8201), .A(n9892), .B(n8200), .ZN(n8203)
         );
  NAND4_X1 U9737 ( .A1(n8206), .A2(n8205), .A3(n8204), .A4(n8203), .ZN(
        P2_U3256) );
  OAI211_X1 U9738 ( .C1(n8208), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9892), .B(
        n8207), .ZN(n8218) );
  AOI21_X1 U9739 ( .B1(n9898), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8209), .ZN(
        n8217) );
  OAI21_X1 U9740 ( .B1(n8212), .B2(n8211), .A(n8210), .ZN(n8213) );
  NAND2_X1 U9741 ( .A1(n9897), .A2(n8213), .ZN(n8216) );
  NAND2_X1 U9742 ( .A1(n9895), .A2(n8214), .ZN(n8215) );
  NAND4_X1 U9743 ( .A1(n8218), .A2(n8217), .A3(n8216), .A4(n8215), .ZN(
        P2_U3260) );
  AOI21_X1 U9744 ( .B1(n8220), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8219), .ZN(
        n8223) );
  NAND2_X1 U9745 ( .A1(n8240), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8221) );
  OAI21_X1 U9746 ( .B1(n8240), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8221), .ZN(
        n8222) );
  AOI211_X1 U9747 ( .C1(n8223), .C2(n8222), .A(n8237), .B(n9414), .ZN(n8236)
         );
  INV_X1 U9748 ( .A(n8240), .ZN(n8233) );
  NOR2_X1 U9749 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8224), .ZN(n8225) );
  AOI21_X1 U9750 ( .B1(n9898), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8225), .ZN(
        n8232) );
  XOR2_X1 U9751 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8240), .Z(n8230) );
  INV_X1 U9752 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8227) );
  AOI21_X1 U9753 ( .B1(n8228), .B2(n8227), .A(n8226), .ZN(n8229) );
  NAND2_X1 U9754 ( .A1(n8230), .A2(n8229), .ZN(n8241) );
  OAI211_X1 U9755 ( .C1(n8230), .C2(n8229), .A(n9892), .B(n8241), .ZN(n8231)
         );
  OAI211_X1 U9756 ( .C1(n8234), .C2(n8233), .A(n8232), .B(n8231), .ZN(n8235)
         );
  OR2_X1 U9757 ( .A1(n8236), .A2(n8235), .ZN(P2_U3262) );
  INV_X1 U9758 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8238) );
  AOI211_X1 U9759 ( .C1(n8239), .C2(n8238), .A(n8255), .B(n9414), .ZN(n8252)
         );
  INV_X1 U9760 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8259) );
  XNOR2_X1 U9761 ( .A(n8258), .B(n8259), .ZN(n8244) );
  NAND2_X1 U9762 ( .A1(n8240), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8242) );
  NAND2_X1 U9763 ( .A1(n8242), .A2(n8241), .ZN(n8243) );
  NOR2_X1 U9764 ( .A1(n8243), .A2(n8244), .ZN(n8257) );
  AOI21_X1 U9765 ( .B1(n8244), .B2(n8243), .A(n8257), .ZN(n8250) );
  INV_X1 U9766 ( .A(n8245), .ZN(n8246) );
  AOI21_X1 U9767 ( .B1(n9898), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8246), .ZN(
        n8249) );
  NAND2_X1 U9768 ( .A1(n9895), .A2(n8247), .ZN(n8248) );
  OAI211_X1 U9769 ( .C1(n9893), .C2(n8250), .A(n8249), .B(n8248), .ZN(n8251)
         );
  OR2_X1 U9770 ( .A1(n8252), .A2(n8251), .ZN(P2_U3263) );
  INV_X1 U9771 ( .A(n9898), .ZN(n8268) );
  NOR2_X1 U9772 ( .A1(n8253), .A2(n8258), .ZN(n8254) );
  NOR2_X1 U9773 ( .A1(n8255), .A2(n8254), .ZN(n8256) );
  INV_X1 U9774 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8722) );
  AOI21_X1 U9775 ( .B1(n8259), .B2(n8258), .A(n8257), .ZN(n8260) );
  XOR2_X1 U9776 ( .A(n8260), .B(P2_REG1_REG_19__SCAN_IN), .Z(n8261) );
  AOI22_X1 U9777 ( .A1(n8263), .A2(n9897), .B1(n9892), .B2(n8261), .ZN(n8265)
         );
  INV_X1 U9778 ( .A(n8261), .ZN(n8264) );
  OAI211_X1 U9779 ( .C1(n8268), .C2(n6898), .A(n8267), .B(n8266), .ZN(P2_U3264) );
  NOR2_X2 U9780 ( .A1(n8609), .A2(n8594), .ZN(n8505) );
  AND2_X2 U9781 ( .A1(n8505), .A2(n8498), .ZN(n8492) );
  NAND2_X1 U9782 ( .A1(n8492), .A2(n8288), .ZN(n8477) );
  NOR2_X2 U9783 ( .A1(n8389), .A2(n8554), .ZN(n8380) );
  AND2_X2 U9784 ( .A1(n8380), .A2(n8360), .ZN(n8356) );
  XNOR2_X1 U9785 ( .A(n8269), .B(n8522), .ZN(n8524) );
  NAND2_X1 U9786 ( .A1(n8270), .A2(P2_B_REG_SCAN_IN), .ZN(n8271) );
  NAND2_X1 U9787 ( .A1(n8603), .A2(n8271), .ZN(n8306) );
  NOR2_X1 U9788 ( .A1(n8272), .A2(n8306), .ZN(n8521) );
  INV_X1 U9789 ( .A(n8521), .ZN(n9452) );
  NOR2_X1 U9790 ( .A1(n4305), .A2(n9452), .ZN(n8277) );
  NOR2_X1 U9791 ( .A1(n8273), .A2(n9438), .ZN(n8274) );
  AOI211_X1 U9792 ( .C1(n4305), .C2(P2_REG2_REG_31__SCAN_IN), .A(n8277), .B(
        n8274), .ZN(n8275) );
  OAI21_X1 U9793 ( .B1(n8443), .B2(n8524), .A(n8275), .ZN(P2_U3265) );
  XNOR2_X1 U9794 ( .A(n8276), .B(n8307), .ZN(n9455) );
  NAND2_X1 U9795 ( .A1(n9455), .A2(n8494), .ZN(n8279) );
  AOI21_X1 U9796 ( .B1(n4305), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8277), .ZN(
        n8278) );
  OAI211_X1 U9797 ( .C1(n9453), .C2(n9438), .A(n8279), .B(n8278), .ZN(P2_U3266) );
  INV_X1 U9798 ( .A(n8578), .ZN(n8453) );
  NAND2_X1 U9799 ( .A1(n8447), .A2(n4856), .ZN(n8432) );
  NAND2_X1 U9800 ( .A1(n8290), .A2(n8458), .ZN(n8292) );
  NAND2_X1 U9801 ( .A1(n8354), .A2(n8353), .ZN(n8352) );
  NAND2_X1 U9802 ( .A1(n8352), .A2(n8298), .ZN(n8334) );
  NAND2_X1 U9803 ( .A1(n8334), .A2(n8342), .ZN(n8333) );
  NAND2_X1 U9804 ( .A1(n8333), .A2(n8299), .ZN(n8316) );
  NAND2_X1 U9805 ( .A1(n8316), .A2(n8323), .ZN(n8315) );
  NAND2_X1 U9806 ( .A1(n8315), .A2(n8301), .ZN(n8302) );
  INV_X1 U9807 ( .A(n8534), .ZN(n8314) );
  AOI21_X1 U9808 ( .B1(n8308), .B2(n8318), .A(n8307), .ZN(n8536) );
  NAND2_X1 U9809 ( .A1(n8536), .A2(n8494), .ZN(n8311) );
  AOI22_X1 U9810 ( .A1(n4305), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8309), .B2(
        n9435), .ZN(n8310) );
  OAI211_X1 U9811 ( .C1(n4546), .C2(n9438), .A(n8311), .B(n8310), .ZN(n8312)
         );
  AOI21_X1 U9812 ( .B1(n8535), .B2(n9441), .A(n8312), .ZN(n8313) );
  OAI21_X1 U9813 ( .B1(n8314), .B2(n9444), .A(n8313), .ZN(P2_U3267) );
  OAI21_X1 U9814 ( .B1(n8316), .B2(n8323), .A(n8315), .ZN(n8317) );
  INV_X1 U9815 ( .A(n8317), .ZN(n8541) );
  INV_X1 U9816 ( .A(n8318), .ZN(n8319) );
  AOI21_X1 U9817 ( .B1(n8537), .B2(n8336), .A(n8319), .ZN(n8538) );
  AOI22_X1 U9818 ( .A1(n8320), .A2(n9435), .B1(n4305), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8321) );
  OAI21_X1 U9819 ( .B1(n4545), .B2(n9438), .A(n8321), .ZN(n8331) );
  INV_X1 U9820 ( .A(n8322), .ZN(n8324) );
  AOI21_X1 U9821 ( .B1(n8324), .B2(n8323), .A(n8512), .ZN(n8329) );
  OAI22_X1 U9822 ( .A1(n8326), .A2(n8457), .B1(n8325), .B2(n8455), .ZN(n8327)
         );
  AOI21_X1 U9823 ( .B1(n8329), .B2(n8328), .A(n8327), .ZN(n8540) );
  NOR2_X1 U9824 ( .A1(n8540), .A2(n4305), .ZN(n8330) );
  AOI211_X1 U9825 ( .C1(n8538), .C2(n8494), .A(n8331), .B(n8330), .ZN(n8332)
         );
  OAI21_X1 U9826 ( .B1(n8541), .B2(n9444), .A(n8332), .ZN(P2_U3268) );
  OAI21_X1 U9827 ( .B1(n8334), .B2(n8342), .A(n8333), .ZN(n8335) );
  INV_X1 U9828 ( .A(n8335), .ZN(n8546) );
  INV_X1 U9829 ( .A(n8356), .ZN(n8338) );
  INV_X1 U9830 ( .A(n8336), .ZN(n8337) );
  AOI21_X1 U9831 ( .B1(n8542), .B2(n8338), .A(n8337), .ZN(n8543) );
  AOI22_X1 U9832 ( .A1(n4305), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8339), .B2(
        n9435), .ZN(n8340) );
  OAI21_X1 U9833 ( .B1(n8341), .B2(n9438), .A(n8340), .ZN(n8350) );
  AOI21_X1 U9834 ( .B1(n8343), .B2(n8342), .A(n8512), .ZN(n8348) );
  OAI22_X1 U9835 ( .A1(n8345), .A2(n8457), .B1(n8344), .B2(n8455), .ZN(n8346)
         );
  AOI21_X1 U9836 ( .B1(n8348), .B2(n8347), .A(n8346), .ZN(n8545) );
  NOR2_X1 U9837 ( .A1(n8545), .A2(n4305), .ZN(n8349) );
  AOI211_X1 U9838 ( .C1(n8543), .C2(n8494), .A(n8350), .B(n8349), .ZN(n8351)
         );
  OAI21_X1 U9839 ( .B1(n8546), .B2(n9444), .A(n8351), .ZN(P2_U3269) );
  OAI21_X1 U9840 ( .B1(n8354), .B2(n8353), .A(n8352), .ZN(n8355) );
  INV_X1 U9841 ( .A(n8355), .ZN(n8551) );
  INV_X1 U9842 ( .A(n8380), .ZN(n8357) );
  AOI211_X1 U9843 ( .C1(n8548), .C2(n8357), .A(n9996), .B(n8356), .ZN(n8547)
         );
  AOI22_X1 U9844 ( .A1(n4305), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8358), .B2(
        n9435), .ZN(n8359) );
  OAI21_X1 U9845 ( .B1(n8360), .B2(n9438), .A(n8359), .ZN(n8368) );
  OAI21_X1 U9846 ( .B1(n8363), .B2(n8362), .A(n8361), .ZN(n8366) );
  AOI222_X1 U9847 ( .A1(n8608), .A2(n8366), .B1(n8365), .B2(n8605), .C1(n8364), 
        .C2(n8603), .ZN(n8550) );
  NOR2_X1 U9848 ( .A1(n8550), .A2(n4305), .ZN(n8367) );
  AOI211_X1 U9849 ( .C1(n8547), .C2(n8519), .A(n8368), .B(n8367), .ZN(n8369)
         );
  OAI21_X1 U9850 ( .B1(n8551), .B2(n9444), .A(n8369), .ZN(P2_U3270) );
  OAI21_X1 U9851 ( .B1(n8372), .B2(n8371), .A(n8370), .ZN(n8373) );
  INV_X1 U9852 ( .A(n8373), .ZN(n8556) );
  OAI211_X1 U9853 ( .C1(n8376), .C2(n8375), .A(n8374), .B(n8608), .ZN(n8379)
         );
  INV_X1 U9854 ( .A(n8377), .ZN(n8378) );
  NAND2_X1 U9855 ( .A1(n8379), .A2(n8378), .ZN(n8552) );
  INV_X1 U9856 ( .A(n8554), .ZN(n8385) );
  AOI211_X1 U9857 ( .C1(n8554), .C2(n8389), .A(n9996), .B(n8380), .ZN(n8553)
         );
  NAND2_X1 U9858 ( .A1(n8553), .A2(n8519), .ZN(n8384) );
  INV_X1 U9859 ( .A(n8381), .ZN(n8382) );
  AOI22_X1 U9860 ( .A1(n4305), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8382), .B2(
        n9435), .ZN(n8383) );
  OAI211_X1 U9861 ( .C1(n8385), .C2(n9438), .A(n8384), .B(n8383), .ZN(n8386)
         );
  AOI21_X1 U9862 ( .B1(n8552), .B2(n9441), .A(n8386), .ZN(n8387) );
  OAI21_X1 U9863 ( .B1(n8556), .B2(n9444), .A(n8387), .ZN(P2_U3271) );
  XNOR2_X1 U9864 ( .A(n8388), .B(n8394), .ZN(n8561) );
  INV_X1 U9865 ( .A(n8389), .ZN(n8390) );
  AOI211_X1 U9866 ( .C1(n8558), .C2(n8404), .A(n9996), .B(n8390), .ZN(n8557)
         );
  INV_X1 U9867 ( .A(n8391), .ZN(n8392) );
  AOI22_X1 U9868 ( .A1(n4305), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8392), .B2(
        n9435), .ZN(n8393) );
  OAI21_X1 U9869 ( .B1(n4695), .B2(n9438), .A(n8393), .ZN(n8400) );
  AOI21_X1 U9870 ( .B1(n8395), .B2(n8394), .A(n8512), .ZN(n8398) );
  AOI21_X1 U9871 ( .B1(n8398), .B2(n8397), .A(n8396), .ZN(n8560) );
  NOR2_X1 U9872 ( .A1(n8560), .A2(n4305), .ZN(n8399) );
  AOI211_X1 U9873 ( .C1(n8557), .C2(n9448), .A(n8400), .B(n8399), .ZN(n8401)
         );
  OAI21_X1 U9874 ( .B1(n8561), .B2(n9444), .A(n8401), .ZN(P2_U3272) );
  OAI21_X1 U9875 ( .B1(n8403), .B2(n8410), .A(n8402), .ZN(n8566) );
  INV_X1 U9876 ( .A(n8404), .ZN(n8405) );
  AOI21_X1 U9877 ( .B1(n8562), .B2(n4540), .A(n8405), .ZN(n8563) );
  AOI22_X1 U9878 ( .A1(n4305), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8406), .B2(
        n9435), .ZN(n8407) );
  OAI21_X1 U9879 ( .B1(n8408), .B2(n9438), .A(n8407), .ZN(n8415) );
  NAND2_X1 U9880 ( .A1(n8427), .A2(n8409), .ZN(n8411) );
  XNOR2_X1 U9881 ( .A(n8411), .B(n8410), .ZN(n8413) );
  AOI21_X1 U9882 ( .B1(n8413), .B2(n8608), .A(n8412), .ZN(n8565) );
  NOR2_X1 U9883 ( .A1(n8565), .A2(n4305), .ZN(n8414) );
  AOI211_X1 U9884 ( .C1(n8563), .C2(n8494), .A(n8415), .B(n8414), .ZN(n8416)
         );
  OAI21_X1 U9885 ( .B1(n8566), .B2(n9444), .A(n8416), .ZN(P2_U3273) );
  XNOR2_X1 U9886 ( .A(n8418), .B(n8417), .ZN(n8571) );
  AOI21_X1 U9887 ( .B1(n8567), .B2(n8441), .A(n8419), .ZN(n8568) );
  AOI22_X1 U9888 ( .A1(n4305), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8420), .B2(
        n9435), .ZN(n8421) );
  OAI21_X1 U9889 ( .B1(n8422), .B2(n9438), .A(n8421), .ZN(n8430) );
  AOI21_X1 U9890 ( .B1(n8424), .B2(n8423), .A(n8512), .ZN(n8428) );
  INV_X1 U9891 ( .A(n8425), .ZN(n8426) );
  AOI21_X1 U9892 ( .B1(n8428), .B2(n8427), .A(n8426), .ZN(n8570) );
  NOR2_X1 U9893 ( .A1(n8570), .A2(n4305), .ZN(n8429) );
  AOI211_X1 U9894 ( .C1(n8568), .C2(n8494), .A(n8430), .B(n8429), .ZN(n8431)
         );
  OAI21_X1 U9895 ( .B1(n8571), .B2(n9444), .A(n8431), .ZN(P2_U3274) );
  XNOR2_X1 U9896 ( .A(n8432), .B(n8433), .ZN(n8577) );
  XNOR2_X1 U9897 ( .A(n8434), .B(n8433), .ZN(n8436) );
  AOI21_X1 U9898 ( .B1(n8436), .B2(n8608), .A(n8435), .ZN(n8576) );
  OAI21_X1 U9899 ( .B1(n8438), .B2(n8437), .A(n8576), .ZN(n8445) );
  NAND2_X1 U9900 ( .A1(n8450), .A2(n8573), .ZN(n8440) );
  NAND2_X1 U9901 ( .A1(n8441), .A2(n8440), .ZN(n8572) );
  AOI22_X1 U9902 ( .A1(n8573), .A2(n8484), .B1(P2_REG2_REG_21__SCAN_IN), .B2(
        n4305), .ZN(n8442) );
  OAI21_X1 U9903 ( .B1(n8572), .B2(n8443), .A(n8442), .ZN(n8444) );
  AOI21_X1 U9904 ( .B1(n8445), .B2(n9441), .A(n8444), .ZN(n8446) );
  OAI21_X1 U9905 ( .B1(n8577), .B2(n9444), .A(n8446), .ZN(P2_U3275) );
  OAI21_X1 U9906 ( .B1(n8449), .B2(n8448), .A(n8447), .ZN(n8582) );
  AOI21_X1 U9907 ( .B1(n8578), .B2(n8477), .A(n8439), .ZN(n8579) );
  AOI22_X1 U9908 ( .A1(n4305), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8451), .B2(
        n9435), .ZN(n8452) );
  OAI21_X1 U9909 ( .B1(n8453), .B2(n9438), .A(n8452), .ZN(n8462) );
  XNOR2_X1 U9910 ( .A(n8454), .B(n4680), .ZN(n8460) );
  OAI22_X1 U9911 ( .A1(n8458), .A2(n8457), .B1(n8456), .B2(n8455), .ZN(n8459)
         );
  AOI21_X1 U9912 ( .B1(n8460), .B2(n8608), .A(n8459), .ZN(n8581) );
  NOR2_X1 U9913 ( .A1(n8581), .A2(n4305), .ZN(n8461) );
  AOI211_X1 U9914 ( .C1(n8579), .C2(n8494), .A(n8462), .B(n8461), .ZN(n8463)
         );
  OAI21_X1 U9915 ( .B1(n8582), .B2(n9444), .A(n8463), .ZN(P2_U3276) );
  OAI21_X1 U9916 ( .B1(n8465), .B2(n8466), .A(n8464), .ZN(n8587) );
  INV_X1 U9917 ( .A(n8466), .ZN(n8473) );
  OR2_X1 U9918 ( .A1(n8467), .A2(n8468), .ZN(n8470) );
  NAND2_X1 U9919 ( .A1(n8470), .A2(n8469), .ZN(n8472) );
  NAND2_X1 U9920 ( .A1(n8472), .A2(n8473), .ZN(n8471) );
  OAI21_X1 U9921 ( .B1(n8473), .B2(n8472), .A(n8471), .ZN(n8476) );
  AOI222_X1 U9922 ( .A1(n8608), .A2(n8476), .B1(n8475), .B2(n8605), .C1(n8474), 
        .C2(n8603), .ZN(n8586) );
  INV_X1 U9923 ( .A(n8492), .ZN(n8479) );
  INV_X1 U9924 ( .A(n8477), .ZN(n8478) );
  AOI211_X1 U9925 ( .C1(n8584), .C2(n8479), .A(n9996), .B(n8478), .ZN(n8583)
         );
  AOI22_X1 U9926 ( .A1(n8583), .A2(n8481), .B1(n9435), .B2(n8480), .ZN(n8482)
         );
  OAI211_X1 U9927 ( .C1(n8587), .C2(n8533), .A(n8586), .B(n8482), .ZN(n8483)
         );
  NAND2_X1 U9928 ( .A1(n8483), .A2(n9441), .ZN(n8486) );
  AOI22_X1 U9929 ( .A1(n8584), .A2(n8484), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n4305), .ZN(n8485) );
  OAI211_X1 U9930 ( .C1(n8587), .C2(n8487), .A(n8486), .B(n8485), .ZN(P2_U3277) );
  XOR2_X1 U9931 ( .A(n8489), .B(n8488), .Z(n8592) );
  XNOR2_X1 U9932 ( .A(n8467), .B(n8489), .ZN(n8491) );
  AOI222_X1 U9933 ( .A1(n8608), .A2(n8491), .B1(n8490), .B2(n8603), .C1(n8604), 
        .C2(n8605), .ZN(n8591) );
  INV_X1 U9934 ( .A(n8591), .ZN(n8500) );
  INV_X1 U9935 ( .A(n8505), .ZN(n8493) );
  AOI21_X1 U9936 ( .B1(n8588), .B2(n8493), .A(n8492), .ZN(n8589) );
  NAND2_X1 U9937 ( .A1(n8589), .A2(n8494), .ZN(n8497) );
  AOI22_X1 U9938 ( .A1(n4305), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8495), .B2(
        n9435), .ZN(n8496) );
  OAI211_X1 U9939 ( .C1(n8498), .C2(n9438), .A(n8497), .B(n8496), .ZN(n8499)
         );
  AOI21_X1 U9940 ( .B1(n8500), .B2(n9441), .A(n8499), .ZN(n8501) );
  OAI21_X1 U9941 ( .B1(n8592), .B2(n9444), .A(n8501), .ZN(P2_U3278) );
  OAI21_X1 U9942 ( .B1(n8503), .B2(n8514), .A(n8502), .ZN(n8504) );
  INV_X1 U9943 ( .A(n8504), .ZN(n8597) );
  AOI211_X1 U9944 ( .C1(n8594), .C2(n8609), .A(n9996), .B(n8505), .ZN(n8593)
         );
  AOI22_X1 U9945 ( .A1(n4305), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8506), .B2(
        n9435), .ZN(n8507) );
  OAI21_X1 U9946 ( .B1(n8285), .B2(n9438), .A(n8507), .ZN(n8518) );
  NAND2_X1 U9947 ( .A1(n8508), .A2(n8509), .ZN(n8513) );
  INV_X1 U9948 ( .A(n8510), .ZN(n8511) );
  AOI211_X1 U9949 ( .C1(n8514), .C2(n8513), .A(n8512), .B(n8511), .ZN(n8516)
         );
  NOR2_X1 U9950 ( .A1(n8516), .A2(n8515), .ZN(n8596) );
  NOR2_X1 U9951 ( .A1(n8596), .A2(n4305), .ZN(n8517) );
  AOI211_X1 U9952 ( .C1(n8593), .C2(n8519), .A(n8518), .B(n8517), .ZN(n8520)
         );
  OAI21_X1 U9953 ( .B1(n8597), .B2(n9444), .A(n8520), .ZN(P2_U3279) );
  AOI21_X1 U9954 ( .B1(n8522), .B2(n9930), .A(n8521), .ZN(n8523) );
  OAI21_X1 U9955 ( .B1(n8524), .B2(n9996), .A(n8523), .ZN(n8615) );
  NAND2_X1 U9956 ( .A1(n8526), .A2(n8525), .ZN(n8528) );
  MUX2_X1 U9957 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8615), .S(n10023), .Z(
        P2_U3551) );
  AND2_X1 U9958 ( .A1(n6109), .A2(n8530), .ZN(n8532) );
  NAND2_X1 U9959 ( .A1(n8532), .A2(n8531), .ZN(n9471) );
  AOI22_X1 U9960 ( .A1(n8538), .A2(n9456), .B1(n9930), .B2(n8537), .ZN(n8539)
         );
  OAI211_X1 U9961 ( .C1(n8541), .C2(n9924), .A(n8540), .B(n8539), .ZN(n8617)
         );
  MUX2_X1 U9962 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8617), .S(n10023), .Z(
        P2_U3548) );
  AOI22_X1 U9963 ( .A1(n8543), .A2(n9456), .B1(n9930), .B2(n8542), .ZN(n8544)
         );
  OAI211_X1 U9964 ( .C1(n8546), .C2(n9924), .A(n8545), .B(n8544), .ZN(n8618)
         );
  MUX2_X1 U9965 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8618), .S(n10023), .Z(
        P2_U3547) );
  AOI21_X1 U9966 ( .B1(n9930), .B2(n8548), .A(n8547), .ZN(n8549) );
  OAI211_X1 U9967 ( .C1(n8551), .C2(n9924), .A(n8550), .B(n8549), .ZN(n8619)
         );
  MUX2_X1 U9968 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8619), .S(n10023), .Z(
        P2_U3546) );
  AOI211_X1 U9969 ( .C1(n9930), .C2(n8554), .A(n8553), .B(n8552), .ZN(n8555)
         );
  OAI21_X1 U9970 ( .B1(n8556), .B2(n9924), .A(n8555), .ZN(n8620) );
  MUX2_X1 U9971 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8620), .S(n10023), .Z(
        P2_U3545) );
  AOI21_X1 U9972 ( .B1(n9930), .B2(n8558), .A(n8557), .ZN(n8559) );
  OAI211_X1 U9973 ( .C1(n8561), .C2(n9924), .A(n8560), .B(n8559), .ZN(n8621)
         );
  MUX2_X1 U9974 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8621), .S(n10023), .Z(
        P2_U3544) );
  AOI22_X1 U9975 ( .A1(n8563), .A2(n9456), .B1(n9930), .B2(n8562), .ZN(n8564)
         );
  OAI211_X1 U9976 ( .C1(n8566), .C2(n9924), .A(n8565), .B(n8564), .ZN(n8622)
         );
  MUX2_X1 U9977 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8622), .S(n10023), .Z(
        P2_U3543) );
  AOI22_X1 U9978 ( .A1(n8568), .A2(n9456), .B1(n9930), .B2(n8567), .ZN(n8569)
         );
  OAI211_X1 U9979 ( .C1(n8571), .C2(n9924), .A(n8570), .B(n8569), .ZN(n8811)
         );
  MUX2_X1 U9980 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8811), .S(n10023), .Z(
        P2_U3542) );
  INV_X1 U9981 ( .A(n8572), .ZN(n8574) );
  AOI22_X1 U9982 ( .A1(n8574), .A2(n9456), .B1(n9930), .B2(n8573), .ZN(n8575)
         );
  OAI211_X1 U9983 ( .C1(n8577), .C2(n9924), .A(n8576), .B(n8575), .ZN(n8812)
         );
  MUX2_X1 U9984 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8812), .S(n10023), .Z(
        P2_U3541) );
  AOI22_X1 U9985 ( .A1(n8579), .A2(n9456), .B1(n9930), .B2(n8578), .ZN(n8580)
         );
  OAI211_X1 U9986 ( .C1(n8582), .C2(n9924), .A(n8581), .B(n8580), .ZN(n8813)
         );
  MUX2_X1 U9987 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8813), .S(n10023), .Z(
        P2_U3540) );
  AOI21_X1 U9988 ( .B1(n9930), .B2(n8584), .A(n8583), .ZN(n8585) );
  OAI211_X1 U9989 ( .C1(n8587), .C2(n9924), .A(n8586), .B(n8585), .ZN(n8814)
         );
  MUX2_X1 U9990 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8814), .S(n10023), .Z(
        P2_U3539) );
  AOI22_X1 U9991 ( .A1(n8589), .A2(n9456), .B1(n9930), .B2(n8588), .ZN(n8590)
         );
  OAI211_X1 U9992 ( .C1(n8592), .C2(n9924), .A(n8591), .B(n8590), .ZN(n8815)
         );
  MUX2_X1 U9993 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8815), .S(n10023), .Z(
        P2_U3538) );
  AOI21_X1 U9994 ( .B1(n9930), .B2(n8594), .A(n8593), .ZN(n8595) );
  OAI211_X1 U9995 ( .C1(n8597), .C2(n9924), .A(n8596), .B(n8595), .ZN(n8816)
         );
  MUX2_X1 U9996 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8816), .S(n10023), .Z(
        P2_U3537) );
  NAND2_X1 U9997 ( .A1(n8598), .A2(n8599), .ZN(n9443) );
  NAND2_X1 U9998 ( .A1(n9443), .A2(n10001), .ZN(n8612) );
  NAND3_X1 U9999 ( .A1(n8601), .A2(n8600), .A3(n4710), .ZN(n8602) );
  NAND2_X1 U10000 ( .A1(n8508), .A2(n8602), .ZN(n8607) );
  AOI222_X1 U10001 ( .A1(n8608), .A2(n8607), .B1(n8606), .B2(n8605), .C1(n8604), .C2(n8603), .ZN(n9434) );
  AOI211_X1 U10002 ( .C1(n8610), .C2(n4336), .A(n9996), .B(n4532), .ZN(n9449)
         );
  AOI21_X1 U10003 ( .B1(n9930), .B2(n8610), .A(n9449), .ZN(n8611) );
  OAI211_X1 U10004 ( .C1(n9446), .C2(n8612), .A(n9434), .B(n8611), .ZN(n8817)
         );
  MUX2_X1 U10005 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8817), .S(n10023), .Z(
        P2_U3536) );
  MUX2_X1 U10006 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8615), .S(n10004), .Z(
        P2_U3519) );
  MUX2_X1 U10007 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8616), .S(n10004), .Z(
        P2_U3517) );
  MUX2_X1 U10008 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8617), .S(n10004), .Z(
        P2_U3516) );
  MUX2_X1 U10009 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8618), .S(n10004), .Z(
        P2_U3515) );
  MUX2_X1 U10010 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8619), .S(n10004), .Z(
        P2_U3514) );
  MUX2_X1 U10011 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8620), .S(n10004), .Z(
        P2_U3513) );
  MUX2_X1 U10012 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8621), .S(n10004), .Z(
        P2_U3512) );
  MUX2_X1 U10013 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8622), .S(n10004), .Z(
        n8810) );
  INV_X1 U10014 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9918) );
  AOI22_X1 U10015 ( .A1(n8624), .A2(keyinput1), .B1(keyinput9), .B2(n9918), 
        .ZN(n8623) );
  OAI221_X1 U10016 ( .B1(n8624), .B2(keyinput1), .C1(n9918), .C2(keyinput9), 
        .A(n8623), .ZN(n8633) );
  AOI22_X1 U10017 ( .A1(n9877), .A2(keyinput36), .B1(keyinput34), .B2(n8626), 
        .ZN(n8625) );
  OAI221_X1 U10018 ( .B1(n9877), .B2(keyinput36), .C1(n8626), .C2(keyinput34), 
        .A(n8625), .ZN(n8632) );
  INV_X1 U10019 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n8725) );
  AOI22_X1 U10020 ( .A1(n8725), .A2(keyinput13), .B1(n8628), .B2(keyinput14), 
        .ZN(n8627) );
  OAI221_X1 U10021 ( .B1(n8725), .B2(keyinput13), .C1(n8628), .C2(keyinput14), 
        .A(n8627), .ZN(n8631) );
  AOI22_X1 U10022 ( .A1(n8712), .A2(keyinput43), .B1(keyinput10), .B2(n8713), 
        .ZN(n8629) );
  OAI221_X1 U10023 ( .B1(n8712), .B2(keyinput43), .C1(n8713), .C2(keyinput10), 
        .A(n8629), .ZN(n8630) );
  NOR4_X1 U10024 ( .A1(n8633), .A2(n8632), .A3(n8631), .A4(n8630), .ZN(n8678)
         );
  AOI22_X1 U10025 ( .A1(P2_REG1_REG_19__SCAN_IN), .A2(keyinput45), .B1(
        P2_REG1_REG_27__SCAN_IN), .B2(keyinput59), .ZN(n8634) );
  OAI221_X1 U10026 ( .B1(P2_REG1_REG_19__SCAN_IN), .B2(keyinput45), .C1(
        P2_REG1_REG_27__SCAN_IN), .C2(keyinput59), .A(n8634), .ZN(n8641) );
  AOI22_X1 U10027 ( .A1(P2_D_REG_29__SCAN_IN), .A2(keyinput25), .B1(
        P1_IR_REG_13__SCAN_IN), .B2(keyinput63), .ZN(n8635) );
  OAI221_X1 U10028 ( .B1(P2_D_REG_29__SCAN_IN), .B2(keyinput25), .C1(
        P1_IR_REG_13__SCAN_IN), .C2(keyinput63), .A(n8635), .ZN(n8640) );
  AOI22_X1 U10029 ( .A1(P2_REG0_REG_20__SCAN_IN), .A2(keyinput2), .B1(
        P2_IR_REG_30__SCAN_IN), .B2(keyinput15), .ZN(n8636) );
  OAI221_X1 U10030 ( .B1(P2_REG0_REG_20__SCAN_IN), .B2(keyinput2), .C1(
        P2_IR_REG_30__SCAN_IN), .C2(keyinput15), .A(n8636), .ZN(n8639) );
  AOI22_X1 U10031 ( .A1(P1_REG0_REG_1__SCAN_IN), .A2(keyinput47), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(keyinput41), .ZN(n8637) );
  OAI221_X1 U10032 ( .B1(P1_REG0_REG_1__SCAN_IN), .B2(keyinput47), .C1(
        P2_DATAO_REG_7__SCAN_IN), .C2(keyinput41), .A(n8637), .ZN(n8638) );
  NOR4_X1 U10033 ( .A1(n8641), .A2(n8640), .A3(n8639), .A4(n8638), .ZN(n8677)
         );
  INV_X1 U10034 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8643) );
  INV_X1 U10035 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9519) );
  AOI22_X1 U10036 ( .A1(n8643), .A2(keyinput55), .B1(keyinput27), .B2(n9519), 
        .ZN(n8642) );
  OAI221_X1 U10037 ( .B1(n8643), .B2(keyinput55), .C1(n9519), .C2(keyinput27), 
        .A(n8642), .ZN(n8649) );
  INV_X1 U10038 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8645) );
  AOI22_X1 U10039 ( .A1(n6837), .A2(keyinput50), .B1(keyinput37), .B2(n8645), 
        .ZN(n8644) );
  OAI221_X1 U10040 ( .B1(n6837), .B2(keyinput50), .C1(n8645), .C2(keyinput37), 
        .A(n8644), .ZN(n8648) );
  INV_X1 U10041 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9037) );
  AOI22_X1 U10042 ( .A1(n6659), .A2(keyinput49), .B1(n9037), .B2(keyinput46), 
        .ZN(n8646) );
  OAI221_X1 U10043 ( .B1(n6659), .B2(keyinput49), .C1(n9037), .C2(keyinput46), 
        .A(n8646), .ZN(n8647) );
  NOR3_X1 U10044 ( .A1(n8649), .A2(n8648), .A3(n8647), .ZN(n8676) );
  INV_X1 U10045 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9978) );
  AOI22_X1 U10046 ( .A1(n9978), .A2(keyinput44), .B1(keyinput52), .B2(n6273), 
        .ZN(n8650) );
  OAI221_X1 U10047 ( .B1(n9978), .B2(keyinput44), .C1(n6273), .C2(keyinput52), 
        .A(n8650), .ZN(n8651) );
  INV_X1 U10048 ( .A(n8651), .ZN(n8674) );
  INV_X1 U10049 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9641) );
  AOI22_X1 U10050 ( .A1(n9641), .A2(keyinput57), .B1(n8779), .B2(keyinput54), 
        .ZN(n8652) );
  OAI221_X1 U10051 ( .B1(n9641), .B2(keyinput57), .C1(n8779), .C2(keyinput54), 
        .A(n8652), .ZN(n8655) );
  AOI22_X1 U10052 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(keyinput4), .B1(
        P1_IR_REG_29__SCAN_IN), .B2(keyinput32), .ZN(n8653) );
  OAI221_X1 U10053 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(keyinput4), .C1(
        P1_IR_REG_29__SCAN_IN), .C2(keyinput32), .A(n8653), .ZN(n8654) );
  NOR2_X1 U10054 ( .A1(n8655), .A2(n8654), .ZN(n8673) );
  AOI22_X1 U10055 ( .A1(P2_D_REG_4__SCAN_IN), .A2(keyinput60), .B1(
        P1_REG0_REG_27__SCAN_IN), .B2(keyinput7), .ZN(n8656) );
  OAI221_X1 U10056 ( .B1(P2_D_REG_4__SCAN_IN), .B2(keyinput60), .C1(
        P1_REG0_REG_27__SCAN_IN), .C2(keyinput7), .A(n8656), .ZN(n8660) );
  XNOR2_X1 U10057 ( .A(keyinput35), .B(P2_REG2_REG_0__SCAN_IN), .ZN(n8658) );
  XNOR2_X1 U10058 ( .A(keyinput33), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n8657) );
  NAND2_X1 U10059 ( .A1(n8658), .A2(n8657), .ZN(n8659) );
  NOR2_X1 U10060 ( .A1(n8660), .A2(n8659), .ZN(n8672) );
  XNOR2_X1 U10061 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput12), .ZN(n8664) );
  XNOR2_X1 U10062 ( .A(SI_19_), .B(keyinput42), .ZN(n8663) );
  XNOR2_X1 U10063 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput23), .ZN(n8662) );
  XNOR2_X1 U10064 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput20), .ZN(n8661) );
  NAND4_X1 U10065 ( .A1(n8664), .A2(n8663), .A3(n8662), .A4(n8661), .ZN(n8670)
         );
  XNOR2_X1 U10066 ( .A(P1_REG1_REG_31__SCAN_IN), .B(keyinput28), .ZN(n8668) );
  XNOR2_X1 U10067 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput17), .ZN(n8667) );
  XNOR2_X1 U10068 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput24), .ZN(n8666) );
  XNOR2_X1 U10069 ( .A(keyinput21), .B(P2_REG2_REG_31__SCAN_IN), .ZN(n8665) );
  NAND4_X1 U10070 ( .A1(n8668), .A2(n8667), .A3(n8666), .A4(n8665), .ZN(n8669)
         );
  NOR2_X1 U10071 ( .A1(n8670), .A2(n8669), .ZN(n8671) );
  AND4_X1 U10072 ( .A1(n8674), .A2(n8673), .A3(n8672), .A4(n8671), .ZN(n8675)
         );
  AND4_X1 U10073 ( .A1(n8678), .A2(n8677), .A3(n8676), .A4(n8675), .ZN(n8808)
         );
  AOI22_X1 U10074 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(keyinput61), .B1(
        P2_D_REG_0__SCAN_IN), .B2(keyinput11), .ZN(n8679) );
  OAI221_X1 U10075 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(keyinput61), .C1(
        P2_D_REG_0__SCAN_IN), .C2(keyinput11), .A(n8679), .ZN(n8686) );
  AOI22_X1 U10076 ( .A1(P2_D_REG_16__SCAN_IN), .A2(keyinput5), .B1(
        P1_REG3_REG_7__SCAN_IN), .B2(keyinput53), .ZN(n8680) );
  OAI221_X1 U10077 ( .B1(P2_D_REG_16__SCAN_IN), .B2(keyinput5), .C1(
        P1_REG3_REG_7__SCAN_IN), .C2(keyinput53), .A(n8680), .ZN(n8685) );
  AOI22_X1 U10078 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(keyinput30), .B1(
        P1_REG0_REG_26__SCAN_IN), .B2(keyinput3), .ZN(n8681) );
  OAI221_X1 U10079 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(keyinput30), .C1(
        P1_REG0_REG_26__SCAN_IN), .C2(keyinput3), .A(n8681), .ZN(n8684) );
  AOI22_X1 U10080 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(keyinput26), .B1(
        P1_D_REG_10__SCAN_IN), .B2(keyinput40), .ZN(n8682) );
  OAI221_X1 U10081 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(keyinput26), .C1(
        P1_D_REG_10__SCAN_IN), .C2(keyinput40), .A(n8682), .ZN(n8683) );
  NOR4_X1 U10082 ( .A1(n8686), .A2(n8685), .A3(n8684), .A4(n8683), .ZN(n8696)
         );
  AOI22_X1 U10083 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(keyinput0), .B1(
        P1_IR_REG_14__SCAN_IN), .B2(keyinput19), .ZN(n8687) );
  OAI221_X1 U10084 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(keyinput0), .C1(
        P1_IR_REG_14__SCAN_IN), .C2(keyinput19), .A(n8687), .ZN(n8694) );
  AOI22_X1 U10085 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(keyinput8), .B1(
        P2_REG1_REG_6__SCAN_IN), .B2(keyinput29), .ZN(n8688) );
  OAI221_X1 U10086 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(keyinput8), .C1(
        P2_REG1_REG_6__SCAN_IN), .C2(keyinput29), .A(n8688), .ZN(n8693) );
  AOI22_X1 U10087 ( .A1(P2_REG1_REG_22__SCAN_IN), .A2(keyinput56), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(keyinput6), .ZN(n8689) );
  OAI221_X1 U10088 ( .B1(P2_REG1_REG_22__SCAN_IN), .B2(keyinput56), .C1(
        P2_DATAO_REG_17__SCAN_IN), .C2(keyinput6), .A(n8689), .ZN(n8692) );
  AOI22_X1 U10089 ( .A1(P2_D_REG_7__SCAN_IN), .A2(keyinput38), .B1(
        P2_IR_REG_8__SCAN_IN), .B2(keyinput18), .ZN(n8690) );
  OAI221_X1 U10090 ( .B1(P2_D_REG_7__SCAN_IN), .B2(keyinput38), .C1(
        P2_IR_REG_8__SCAN_IN), .C2(keyinput18), .A(n8690), .ZN(n8691) );
  NOR4_X1 U10091 ( .A1(n8694), .A2(n8693), .A3(n8692), .A4(n8691), .ZN(n8695)
         );
  AND2_X1 U10092 ( .A1(n8696), .A2(n8695), .ZN(n8807) );
  INV_X1 U10093 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9786) );
  AOI22_X1 U10094 ( .A1(n9786), .A2(keyinput51), .B1(keyinput39), .B2(n8698), 
        .ZN(n8697) );
  OAI221_X1 U10095 ( .B1(n9786), .B2(keyinput51), .C1(n8698), .C2(keyinput39), 
        .A(n8697), .ZN(n8708) );
  AOI22_X1 U10096 ( .A1(n8722), .A2(keyinput31), .B1(n8700), .B2(keyinput48), 
        .ZN(n8699) );
  OAI221_X1 U10097 ( .B1(n8722), .B2(keyinput31), .C1(n8700), .C2(keyinput48), 
        .A(n8699), .ZN(n8707) );
  AOI22_X1 U10098 ( .A1(n8710), .A2(keyinput22), .B1(n8702), .B2(keyinput62), 
        .ZN(n8701) );
  OAI221_X1 U10099 ( .B1(n8710), .B2(keyinput22), .C1(n8702), .C2(keyinput62), 
        .A(n8701), .ZN(n8706) );
  INV_X1 U10100 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9835) );
  AOI22_X1 U10101 ( .A1(n8704), .A2(keyinput16), .B1(keyinput58), .B2(n9835), 
        .ZN(n8703) );
  OAI221_X1 U10102 ( .B1(n8704), .B2(keyinput16), .C1(n9835), .C2(keyinput58), 
        .A(n8703), .ZN(n8705) );
  NOR4_X1 U10103 ( .A1(n8708), .A2(n8707), .A3(n8706), .A4(n8705), .ZN(n8806)
         );
  INV_X1 U10104 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n9787) );
  AOI22_X1 U10105 ( .A1(n9787), .A2(keyinput104), .B1(keyinput86), .B2(n8710), 
        .ZN(n8709) );
  OAI221_X1 U10106 ( .B1(n9787), .B2(keyinput104), .C1(n8710), .C2(keyinput86), 
        .A(n8709), .ZN(n8720) );
  AOI22_X1 U10107 ( .A1(n8713), .A2(keyinput74), .B1(n8712), .B2(keyinput107), 
        .ZN(n8711) );
  OAI221_X1 U10108 ( .B1(n8713), .B2(keyinput74), .C1(n8712), .C2(keyinput107), 
        .A(n8711), .ZN(n8719) );
  INV_X1 U10109 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9678) );
  AOI22_X1 U10110 ( .A1(n9678), .A2(keyinput64), .B1(n5025), .B2(keyinput117), 
        .ZN(n8714) );
  OAI221_X1 U10111 ( .B1(n9678), .B2(keyinput64), .C1(n5025), .C2(keyinput117), 
        .A(n8714), .ZN(n8718) );
  INV_X1 U10112 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n9905) );
  INV_X1 U10113 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8716) );
  AOI22_X1 U10114 ( .A1(n9905), .A2(keyinput102), .B1(keyinput66), .B2(n8716), 
        .ZN(n8715) );
  OAI221_X1 U10115 ( .B1(n9905), .B2(keyinput102), .C1(n8716), .C2(keyinput66), 
        .A(n8715), .ZN(n8717) );
  NOR4_X1 U10116 ( .A1(n8720), .A2(n8719), .A3(n8718), .A4(n8717), .ZN(n8804)
         );
  AOI22_X1 U10117 ( .A1(n8723), .A2(keyinput71), .B1(keyinput95), .B2(n8722), 
        .ZN(n8721) );
  OAI221_X1 U10118 ( .B1(n8723), .B2(keyinput71), .C1(n8722), .C2(keyinput95), 
        .A(n8721), .ZN(n8728) );
  AOI22_X1 U10119 ( .A1(n8726), .A2(keyinput83), .B1(keyinput77), .B2(n8725), 
        .ZN(n8724) );
  OAI221_X1 U10120 ( .B1(n8726), .B2(keyinput83), .C1(n8725), .C2(keyinput77), 
        .A(n8724), .ZN(n8727) );
  NOR2_X1 U10121 ( .A1(n8728), .A2(n8727), .ZN(n8741) );
  INV_X1 U10122 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8730) );
  AOI22_X1 U10123 ( .A1(n8730), .A2(keyinput120), .B1(n9519), .B2(keyinput91), 
        .ZN(n8729) );
  OAI221_X1 U10124 ( .B1(n8730), .B2(keyinput120), .C1(n9519), .C2(keyinput91), 
        .A(n8729), .ZN(n8731) );
  INV_X1 U10125 ( .A(n8731), .ZN(n8740) );
  AOI22_X1 U10126 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(keyinput72), .B1(
        P2_IR_REG_13__SCAN_IN), .B2(keyinput88), .ZN(n8732) );
  OAI221_X1 U10127 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(keyinput72), .C1(
        P2_IR_REG_13__SCAN_IN), .C2(keyinput88), .A(n8732), .ZN(n8735) );
  AOI22_X1 U10128 ( .A1(P2_REG0_REG_0__SCAN_IN), .A2(keyinput73), .B1(
        P1_REG1_REG_15__SCAN_IN), .B2(keyinput94), .ZN(n8733) );
  OAI221_X1 U10129 ( .B1(P2_REG0_REG_0__SCAN_IN), .B2(keyinput73), .C1(
        P1_REG1_REG_15__SCAN_IN), .C2(keyinput94), .A(n8733), .ZN(n8734) );
  NOR2_X1 U10130 ( .A1(n8735), .A2(n8734), .ZN(n8739) );
  AOI22_X1 U10131 ( .A1(n9896), .A2(keyinput99), .B1(n6307), .B2(keyinput93), 
        .ZN(n8736) );
  OAI221_X1 U10132 ( .B1(n9896), .B2(keyinput99), .C1(n6307), .C2(keyinput93), 
        .A(n8736), .ZN(n8737) );
  INV_X1 U10133 ( .A(n8737), .ZN(n8738) );
  NAND4_X1 U10134 ( .A1(n8741), .A2(n8740), .A3(n8739), .A4(n8738), .ZN(n8751)
         );
  OAI22_X1 U10135 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(keyinput76), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(keyinput125), .ZN(n8742) );
  AOI221_X1 U10136 ( .B1(P1_DATAO_REG_2__SCAN_IN), .B2(keyinput76), .C1(
        keyinput125), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n8742), .ZN(n8749) );
  OAI22_X1 U10137 ( .A1(SI_9_), .A2(keyinput65), .B1(keyinput110), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n8743) );
  AOI221_X1 U10138 ( .B1(SI_9_), .B2(keyinput65), .C1(P1_REG2_REG_19__SCAN_IN), 
        .C2(keyinput110), .A(n8743), .ZN(n8748) );
  OAI22_X1 U10139 ( .A1(P1_REG0_REG_26__SCAN_IN), .A2(keyinput67), .B1(
        keyinput113), .B2(P2_REG2_REG_7__SCAN_IN), .ZN(n8744) );
  AOI221_X1 U10140 ( .B1(P1_REG0_REG_26__SCAN_IN), .B2(keyinput67), .C1(
        P2_REG2_REG_7__SCAN_IN), .C2(keyinput113), .A(n8744), .ZN(n8747) );
  OAI22_X1 U10141 ( .A1(P1_REG1_REG_20__SCAN_IN), .A2(keyinput119), .B1(
        P2_REG0_REG_9__SCAN_IN), .B2(keyinput108), .ZN(n8745) );
  AOI221_X1 U10142 ( .B1(P1_REG1_REG_20__SCAN_IN), .B2(keyinput119), .C1(
        keyinput108), .C2(P2_REG0_REG_9__SCAN_IN), .A(n8745), .ZN(n8746) );
  NAND4_X1 U10143 ( .A1(n8749), .A2(n8748), .A3(n8747), .A4(n8746), .ZN(n8750)
         );
  NOR2_X1 U10144 ( .A1(n8751), .A2(n8750), .ZN(n8803) );
  OAI22_X1 U10145 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(keyinput116), .B1(
        P1_ADDR_REG_3__SCAN_IN), .B2(keyinput98), .ZN(n8752) );
  AOI221_X1 U10146 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(keyinput116), .C1(
        keyinput98), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n8752), .ZN(n8759) );
  OAI22_X1 U10147 ( .A1(P2_REG2_REG_27__SCAN_IN), .A2(keyinput101), .B1(
        P1_REG1_REG_31__SCAN_IN), .B2(keyinput92), .ZN(n8753) );
  AOI221_X1 U10148 ( .B1(P2_REG2_REG_27__SCAN_IN), .B2(keyinput101), .C1(
        keyinput92), .C2(P1_REG1_REG_31__SCAN_IN), .A(n8753), .ZN(n8758) );
  OAI22_X1 U10149 ( .A1(P1_D_REG_27__SCAN_IN), .A2(keyinput115), .B1(SI_16_), 
        .B2(keyinput78), .ZN(n8754) );
  AOI221_X1 U10150 ( .B1(P1_D_REG_27__SCAN_IN), .B2(keyinput115), .C1(
        keyinput78), .C2(SI_16_), .A(n8754), .ZN(n8757) );
  OAI22_X1 U10151 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(keyinput82), .B1(
        P2_D_REG_0__SCAN_IN), .B2(keyinput75), .ZN(n8755) );
  AOI221_X1 U10152 ( .B1(P2_IR_REG_8__SCAN_IN), .B2(keyinput82), .C1(
        keyinput75), .C2(P2_D_REG_0__SCAN_IN), .A(n8755), .ZN(n8756) );
  NAND4_X1 U10153 ( .A1(n8759), .A2(n8758), .A3(n8757), .A4(n8756), .ZN(n8769)
         );
  OAI22_X1 U10154 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(keyinput96), .B1(
        keyinput122), .B2(P1_REG0_REG_6__SCAN_IN), .ZN(n8760) );
  AOI221_X1 U10155 ( .B1(P1_IR_REG_29__SCAN_IN), .B2(keyinput96), .C1(
        P1_REG0_REG_6__SCAN_IN), .C2(keyinput122), .A(n8760), .ZN(n8767) );
  OAI22_X1 U10156 ( .A1(P2_D_REG_4__SCAN_IN), .A2(keyinput124), .B1(
        P2_ADDR_REG_15__SCAN_IN), .B2(keyinput90), .ZN(n8761) );
  AOI221_X1 U10157 ( .B1(P2_D_REG_4__SCAN_IN), .B2(keyinput124), .C1(
        keyinput90), .C2(P2_ADDR_REG_15__SCAN_IN), .A(n8761), .ZN(n8766) );
  OAI22_X1 U10158 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(keyinput97), .B1(
        P2_D_REG_29__SCAN_IN), .B2(keyinput89), .ZN(n8762) );
  AOI221_X1 U10159 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(keyinput97), .C1(
        keyinput89), .C2(P2_D_REG_29__SCAN_IN), .A(n8762), .ZN(n8765) );
  OAI22_X1 U10160 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(keyinput80), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(keyinput112), .ZN(n8763) );
  AOI221_X1 U10161 ( .B1(P1_DATAO_REG_18__SCAN_IN), .B2(keyinput80), .C1(
        keyinput112), .C2(P2_DATAO_REG_18__SCAN_IN), .A(n8763), .ZN(n8764) );
  NAND4_X1 U10162 ( .A1(n8767), .A2(n8766), .A3(n8765), .A4(n8764), .ZN(n8768)
         );
  NOR2_X1 U10163 ( .A1(n8769), .A2(n8768), .ZN(n8802) );
  OAI22_X1 U10164 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(keyinput100), .B1(
        keyinput121), .B2(P1_ADDR_REG_13__SCAN_IN), .ZN(n8770) );
  AOI221_X1 U10165 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(keyinput100), .C1(
        P1_ADDR_REG_13__SCAN_IN), .C2(keyinput121), .A(n8770), .ZN(n8777) );
  OAI22_X1 U10166 ( .A1(SI_19_), .A2(keyinput106), .B1(P1_REG2_REG_6__SCAN_IN), 
        .B2(keyinput114), .ZN(n8771) );
  AOI221_X1 U10167 ( .B1(SI_19_), .B2(keyinput106), .C1(keyinput114), .C2(
        P1_REG2_REG_6__SCAN_IN), .A(n8771), .ZN(n8776) );
  OAI22_X1 U10168 ( .A1(P2_D_REG_16__SCAN_IN), .A2(keyinput69), .B1(keyinput79), .B2(P2_IR_REG_30__SCAN_IN), .ZN(n8772) );
  AOI221_X1 U10169 ( .B1(P2_D_REG_16__SCAN_IN), .B2(keyinput69), .C1(
        P2_IR_REG_30__SCAN_IN), .C2(keyinput79), .A(n8772), .ZN(n8775) );
  OAI22_X1 U10170 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(keyinput126), .B1(
        keyinput85), .B2(P2_REG2_REG_31__SCAN_IN), .ZN(n8773) );
  AOI221_X1 U10171 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(keyinput126), .C1(
        P2_REG2_REG_31__SCAN_IN), .C2(keyinput85), .A(n8773), .ZN(n8774) );
  NAND4_X1 U10172 ( .A1(n8777), .A2(n8776), .A3(n8775), .A4(n8774), .ZN(n8800)
         );
  INV_X1 U10173 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8780) );
  AOI22_X1 U10174 ( .A1(n8780), .A2(keyinput68), .B1(n8779), .B2(keyinput118), 
        .ZN(n8778) );
  OAI221_X1 U10175 ( .B1(n8780), .B2(keyinput68), .C1(n8779), .C2(keyinput118), 
        .A(n8778), .ZN(n8781) );
  INV_X1 U10176 ( .A(n8781), .ZN(n8798) );
  INV_X1 U10177 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8783) );
  AOI22_X1 U10178 ( .A1(n8784), .A2(keyinput105), .B1(keyinput109), .B2(n8783), 
        .ZN(n8782) );
  OAI221_X1 U10179 ( .B1(n8784), .B2(keyinput105), .C1(n8783), .C2(keyinput109), .A(n8782), .ZN(n8785) );
  INV_X1 U10180 ( .A(n8785), .ZN(n8797) );
  XNOR2_X1 U10181 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput81), .ZN(n8789) );
  XNOR2_X1 U10182 ( .A(P2_REG1_REG_27__SCAN_IN), .B(keyinput123), .ZN(n8788)
         );
  XNOR2_X1 U10183 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput87), .ZN(n8787) );
  XNOR2_X1 U10184 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput70), .ZN(n8786)
         );
  NAND4_X1 U10185 ( .A1(n8789), .A2(n8788), .A3(n8787), .A4(n8786), .ZN(n8795)
         );
  XNOR2_X1 U10186 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput103), .ZN(n8793)
         );
  XNOR2_X1 U10187 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput84), .ZN(n8792) );
  XNOR2_X1 U10188 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput127), .ZN(n8791) );
  XNOR2_X1 U10189 ( .A(keyinput111), .B(P1_REG0_REG_1__SCAN_IN), .ZN(n8790) );
  NAND4_X1 U10190 ( .A1(n8793), .A2(n8792), .A3(n8791), .A4(n8790), .ZN(n8794)
         );
  NOR2_X1 U10191 ( .A1(n8795), .A2(n8794), .ZN(n8796) );
  NAND3_X1 U10192 ( .A1(n8798), .A2(n8797), .A3(n8796), .ZN(n8799) );
  NOR2_X1 U10193 ( .A1(n8800), .A2(n8799), .ZN(n8801) );
  NAND4_X1 U10194 ( .A1(n8804), .A2(n8803), .A3(n8802), .A4(n8801), .ZN(n8805)
         );
  NAND4_X1 U10195 ( .A1(n8808), .A2(n8807), .A3(n8806), .A4(n8805), .ZN(n8809)
         );
  XNOR2_X1 U10196 ( .A(n8810), .B(n8809), .ZN(P2_U3511) );
  MUX2_X1 U10197 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8811), .S(n10004), .Z(
        P2_U3510) );
  MUX2_X1 U10198 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8812), .S(n10004), .Z(
        P2_U3509) );
  MUX2_X1 U10199 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8813), .S(n10004), .Z(
        P2_U3508) );
  MUX2_X1 U10200 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8814), .S(n10004), .Z(
        P2_U3507) );
  MUX2_X1 U10201 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8815), .S(n10004), .Z(
        P2_U3505) );
  MUX2_X1 U10202 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8816), .S(n10004), .Z(
        P2_U3502) );
  MUX2_X1 U10203 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8817), .S(n10004), .Z(
        P2_U3499) );
  INV_X1 U10204 ( .A(n8818), .ZN(n9383) );
  INV_X1 U10205 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8819) );
  NAND3_X1 U10206 ( .A1(n8819), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8821) );
  OAI22_X1 U10207 ( .A1(n5922), .A2(n8821), .B1(n8820), .B2(n8827), .ZN(n8822)
         );
  INV_X1 U10208 ( .A(n8822), .ZN(n8823) );
  OAI21_X1 U10209 ( .B1(n9383), .B2(n8840), .A(n8823), .ZN(P2_U3327) );
  OAI222_X1 U10210 ( .A1(n8827), .A2(n8826), .B1(n8840), .B2(n8825), .C1(
        P2_U3152), .C2(n8824), .ZN(P2_U3328) );
  INV_X1 U10211 ( .A(n8828), .ZN(n9386) );
  OAI222_X1 U10212 ( .A1(n8827), .A2(n8830), .B1(n8840), .B2(n9386), .C1(n8829), .C2(P2_U3152), .ZN(P2_U3329) );
  INV_X1 U10213 ( .A(n8831), .ZN(n9393) );
  OAI222_X1 U10214 ( .A1(n8827), .A2(n8832), .B1(n8840), .B2(n9393), .C1(n6264), .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U10215 ( .A(n8833), .ZN(n9396) );
  OAI222_X1 U10216 ( .A1(n8836), .A2(P2_U3152), .B1(n8835), .B2(n9396), .C1(
        n8834), .C2(n8827), .ZN(P2_U3332) );
  INV_X1 U10217 ( .A(n8837), .ZN(n9399) );
  OAI222_X1 U10218 ( .A1(n8827), .A2(n8841), .B1(n8840), .B2(n9399), .C1(n8839), .C2(P2_U3152), .ZN(P2_U3333) );
  MUX2_X1 U10219 ( .A(n8842), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10220 ( .A(n8845), .B(n8844), .ZN(n8846) );
  XNOR2_X1 U10221 ( .A(n8843), .B(n8846), .ZN(n8855) );
  NOR2_X1 U10222 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8847), .ZN(n9645) );
  AOI21_X1 U10223 ( .B1(n8992), .B2(n9262), .A(n9645), .ZN(n8853) );
  NAND2_X1 U10224 ( .A1(n8965), .A2(n8848), .ZN(n8852) );
  NAND2_X1 U10225 ( .A1(n8997), .A2(n8849), .ZN(n8851) );
  NAND2_X1 U10226 ( .A1(n8966), .A2(n9491), .ZN(n8850) );
  NAND4_X1 U10227 ( .A1(n8853), .A2(n8852), .A3(n8851), .A4(n8850), .ZN(n8854)
         );
  AOI21_X1 U10228 ( .B1(n8855), .B2(n8977), .A(n8854), .ZN(n8856) );
  INV_X1 U10229 ( .A(n8856), .ZN(P1_U3213) );
  INV_X1 U10230 ( .A(n8857), .ZN(n8859) );
  NOR2_X1 U10231 ( .A1(n8859), .A2(n8858), .ZN(n8861) );
  XNOR2_X1 U10232 ( .A(n8861), .B(n8860), .ZN(n8866) );
  AOI22_X1 U10233 ( .A1(n8992), .A2(n9154), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8863) );
  NAND2_X1 U10234 ( .A1(n8997), .A2(n9145), .ZN(n8862) );
  OAI211_X1 U10235 ( .C1(n8882), .C2(n8994), .A(n8863), .B(n8862), .ZN(n8864)
         );
  AOI21_X1 U10236 ( .B1(n9327), .B2(n8965), .A(n8864), .ZN(n8865) );
  OAI21_X1 U10237 ( .B1(n8866), .B2(n8988), .A(n8865), .ZN(P1_U3214) );
  INV_X1 U10238 ( .A(n8870), .ZN(n8868) );
  NAND2_X1 U10239 ( .A1(n8868), .A2(n8867), .ZN(n8976) );
  NAND2_X1 U10240 ( .A1(n8976), .A2(n8974), .ZN(n8973) );
  NAND2_X1 U10241 ( .A1(n8870), .A2(n8869), .ZN(n8975) );
  OR2_X1 U10242 ( .A1(n5694), .A2(n8925), .ZN(n8872) );
  AOI21_X1 U10243 ( .B1(n8973), .B2(n8975), .A(n8872), .ZN(n8926) );
  AND3_X1 U10244 ( .A1(n8973), .A2(n8975), .A3(n8872), .ZN(n8873) );
  OAI21_X1 U10245 ( .B1(n8926), .B2(n8873), .A(n8977), .ZN(n8877) );
  NAND2_X1 U10246 ( .A1(n8992), .A2(n9216), .ZN(n8874) );
  NAND2_X1 U10247 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9058) );
  OAI211_X1 U10248 ( .C1(n8911), .C2(n8994), .A(n8874), .B(n9058), .ZN(n8875)
         );
  AOI21_X1 U10249 ( .B1(n9210), .B2(n8997), .A(n8875), .ZN(n8876) );
  OAI211_X1 U10250 ( .C1(n9212), .C2(n9000), .A(n8877), .B(n8876), .ZN(
        P1_U3217) );
  AOI21_X1 U10251 ( .B1(n8879), .B2(n8878), .A(n4366), .ZN(n8885) );
  AOI22_X1 U10252 ( .A1(n8966), .A2(n9216), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8881) );
  NAND2_X1 U10253 ( .A1(n8997), .A2(n9188), .ZN(n8880) );
  OAI211_X1 U10254 ( .C1(n8882), .C2(n8953), .A(n8881), .B(n8880), .ZN(n8883)
         );
  AOI21_X1 U10255 ( .B1(n9185), .B2(n8965), .A(n8883), .ZN(n8884) );
  OAI21_X1 U10256 ( .B1(n8885), .B2(n8988), .A(n8884), .ZN(P1_U3221) );
  OAI21_X1 U10257 ( .B1(n8887), .B2(n8886), .A(n5747), .ZN(n8888) );
  NAND2_X1 U10258 ( .A1(n8888), .A2(n8977), .ZN(n8893) );
  AOI22_X1 U10259 ( .A1(n9122), .A2(n8992), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8889) );
  OAI21_X1 U10260 ( .B1(n8890), .B2(n8994), .A(n8889), .ZN(n8891) );
  AOI21_X1 U10261 ( .B1(n9117), .B2(n8997), .A(n8891), .ZN(n8892) );
  OAI211_X1 U10262 ( .C1(n9119), .C2(n9000), .A(n8893), .B(n8892), .ZN(
        P1_U3223) );
  INV_X1 U10263 ( .A(n8895), .ZN(n8899) );
  AOI21_X1 U10264 ( .B1(n8896), .B2(n8987), .A(n8897), .ZN(n8898) );
  OAI21_X1 U10265 ( .B1(n8899), .B2(n8898), .A(n8977), .ZN(n8905) );
  NOR2_X1 U10266 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8900), .ZN(n9670) );
  AOI21_X1 U10267 ( .B1(n8992), .B2(n9261), .A(n9670), .ZN(n8901) );
  OAI21_X1 U10268 ( .B1(n8902), .B2(n8994), .A(n8901), .ZN(n8903) );
  AOI21_X1 U10269 ( .B1(n9265), .B2(n8997), .A(n8903), .ZN(n8904) );
  OAI211_X1 U10270 ( .C1(n4499), .C2(n9000), .A(n8905), .B(n8904), .ZN(
        P1_U3224) );
  INV_X1 U10271 ( .A(n9359), .ZN(n9246) );
  OAI21_X1 U10272 ( .B1(n8908), .B2(n8907), .A(n8906), .ZN(n8909) );
  NAND2_X1 U10273 ( .A1(n8909), .A2(n8977), .ZN(n8914) );
  NAND2_X1 U10274 ( .A1(n8966), .A2(n9276), .ZN(n8910) );
  NAND2_X1 U10275 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9683) );
  OAI211_X1 U10276 ( .C1(n8911), .C2(n8953), .A(n8910), .B(n9683), .ZN(n8912)
         );
  AOI21_X1 U10277 ( .B1(n9244), .B2(n8997), .A(n8912), .ZN(n8913) );
  OAI211_X1 U10278 ( .C1(n9246), .C2(n9000), .A(n8914), .B(n8913), .ZN(
        P1_U3226) );
  OAI21_X1 U10279 ( .B1(n8917), .B2(n8916), .A(n8915), .ZN(n8918) );
  NAND2_X1 U10280 ( .A1(n8918), .A2(n8977), .ZN(n8922) );
  AOI22_X1 U10281 ( .A1(n8992), .A2(n9131), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8919) );
  OAI21_X1 U10282 ( .B1(n8952), .B2(n8994), .A(n8919), .ZN(n8920) );
  AOI21_X1 U10283 ( .B1(n9135), .B2(n8997), .A(n8920), .ZN(n8921) );
  OAI211_X1 U10284 ( .C1(n9128), .C2(n9000), .A(n8922), .B(n8921), .ZN(
        P1_U3227) );
  INV_X1 U10285 ( .A(n8923), .ZN(n8924) );
  NOR3_X1 U10286 ( .A1(n8926), .A2(n8925), .A3(n8924), .ZN(n8928) );
  OAI21_X1 U10287 ( .B1(n8928), .B2(n8927), .A(n8977), .ZN(n8933) );
  INV_X1 U10288 ( .A(n8955), .ZN(n9201) );
  AOI22_X1 U10289 ( .A1(n8992), .A2(n9201), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8929) );
  OAI21_X1 U10290 ( .B1(n8930), .B2(n8994), .A(n8929), .ZN(n8931) );
  AOI21_X1 U10291 ( .B1(n9196), .B2(n8997), .A(n8931), .ZN(n8932) );
  OAI211_X1 U10292 ( .C1(n9198), .C2(n9000), .A(n8933), .B(n8932), .ZN(
        P1_U3231) );
  XNOR2_X1 U10293 ( .A(n8936), .B(n8935), .ZN(n8937) );
  XNOR2_X1 U10294 ( .A(n8934), .B(n8937), .ZN(n8945) );
  AND2_X1 U10295 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9633) );
  AOI21_X1 U10296 ( .B1(n8992), .B2(n9275), .A(n9633), .ZN(n8943) );
  NAND2_X1 U10297 ( .A1(n8965), .A2(n8938), .ZN(n8942) );
  NAND2_X1 U10298 ( .A1(n8997), .A2(n8939), .ZN(n8941) );
  NAND2_X1 U10299 ( .A1(n8966), .A2(n9004), .ZN(n8940) );
  NAND4_X1 U10300 ( .A1(n8943), .A2(n8942), .A3(n8941), .A4(n8940), .ZN(n8944)
         );
  AOI21_X1 U10301 ( .B1(n8945), .B2(n8977), .A(n8944), .ZN(n8946) );
  INV_X1 U10302 ( .A(n8946), .ZN(P1_U3232) );
  NAND2_X1 U10303 ( .A1(n8948), .A2(n8947), .ZN(n8950) );
  XNOR2_X1 U10304 ( .A(n8950), .B(n8949), .ZN(n8951) );
  NAND2_X1 U10305 ( .A1(n8951), .A2(n8977), .ZN(n8959) );
  NOR2_X1 U10306 ( .A1(n8953), .A2(n8952), .ZN(n8957) );
  OAI22_X1 U10307 ( .A1(n8994), .A2(n8955), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8954), .ZN(n8956) );
  AOI211_X1 U10308 ( .C1(n9162), .C2(n8997), .A(n8957), .B(n8956), .ZN(n8958)
         );
  OAI211_X1 U10309 ( .C1(n9164), .C2(n9000), .A(n8959), .B(n8958), .ZN(
        P1_U3233) );
  OAI21_X1 U10310 ( .B1(n8962), .B2(n8960), .A(n8961), .ZN(n8963) );
  NAND2_X1 U10311 ( .A1(n8963), .A2(n8977), .ZN(n8971) );
  AOI22_X1 U10312 ( .A1(n8966), .A2(n5562), .B1(n8965), .B2(n8964), .ZN(n8970)
         );
  AOI22_X1 U10313 ( .A1(n8992), .A2(n8967), .B1(n8968), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n8969) );
  NAND3_X1 U10314 ( .A1(n8971), .A2(n8970), .A3(n8969), .ZN(P1_U3235) );
  INV_X1 U10315 ( .A(n8975), .ZN(n8972) );
  NOR2_X1 U10316 ( .A1(n8973), .A2(n8972), .ZN(n8979) );
  AOI21_X1 U10317 ( .B1(n8976), .B2(n8975), .A(n8974), .ZN(n8978) );
  OAI21_X1 U10318 ( .B1(n8979), .B2(n8978), .A(n8977), .ZN(n8984) );
  NAND2_X1 U10319 ( .A1(n8992), .A2(n9230), .ZN(n8980) );
  NAND2_X1 U10320 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9699) );
  OAI211_X1 U10321 ( .C1(n8981), .C2(n8994), .A(n8980), .B(n9699), .ZN(n8982)
         );
  AOI21_X1 U10322 ( .B1(n9236), .B2(n8997), .A(n8982), .ZN(n8983) );
  OAI211_X1 U10323 ( .C1(n9239), .C2(n9000), .A(n8984), .B(n8983), .ZN(
        P1_U3236) );
  INV_X1 U10324 ( .A(n8987), .ZN(n8991) );
  AOI21_X1 U10325 ( .B1(n8987), .B2(n8986), .A(n8985), .ZN(n8989) );
  NOR2_X1 U10326 ( .A1(n8989), .A2(n8988), .ZN(n8990) );
  OAI21_X1 U10327 ( .B1(n8991), .B2(n8896), .A(n8990), .ZN(n8999) );
  AND2_X1 U10328 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9658) );
  AOI21_X1 U10329 ( .B1(n8992), .B2(n9276), .A(n9658), .ZN(n8993) );
  OAI21_X1 U10330 ( .B1(n8995), .B2(n8994), .A(n8993), .ZN(n8996) );
  AOI21_X1 U10331 ( .B1(n9282), .B2(n8997), .A(n8996), .ZN(n8998) );
  OAI211_X1 U10332 ( .C1(n9520), .C2(n9000), .A(n8999), .B(n8998), .ZN(
        P1_U3239) );
  MUX2_X1 U10333 ( .A(n9061), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9011), .Z(
        P1_U3586) );
  MUX2_X1 U10334 ( .A(n9001), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9011), .Z(
        P1_U3585) );
  MUX2_X1 U10335 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9080), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10336 ( .A(n9002), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9011), .Z(
        P1_U3583) );
  INV_X1 U10337 ( .A(n9003), .ZN(n9110) );
  MUX2_X1 U10338 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9110), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10339 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9122), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10340 ( .A(n9131), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9011), .Z(
        P1_U3580) );
  MUX2_X1 U10341 ( .A(n9154), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9011), .Z(
        P1_U3579) );
  MUX2_X1 U10342 ( .A(n9167), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9011), .Z(
        P1_U3578) );
  MUX2_X1 U10343 ( .A(n9182), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9011), .Z(
        P1_U3577) );
  MUX2_X1 U10344 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9201), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10345 ( .A(n9216), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9011), .Z(
        P1_U3575) );
  MUX2_X1 U10346 ( .A(n9230), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9011), .Z(
        P1_U3574) );
  MUX2_X1 U10347 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9248), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10348 ( .A(n9261), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9011), .Z(
        P1_U3572) );
  MUX2_X1 U10349 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9276), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10350 ( .A(n9262), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9011), .Z(
        P1_U3570) );
  MUX2_X1 U10351 ( .A(n9275), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9011), .Z(
        P1_U3569) );
  MUX2_X1 U10352 ( .A(n9491), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9011), .Z(
        P1_U3568) );
  MUX2_X1 U10353 ( .A(n9004), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9011), .Z(
        P1_U3567) );
  MUX2_X1 U10354 ( .A(n9490), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9011), .Z(
        P1_U3566) );
  MUX2_X1 U10355 ( .A(n9005), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9011), .Z(
        P1_U3565) );
  MUX2_X1 U10356 ( .A(n9006), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9011), .Z(
        P1_U3564) );
  MUX2_X1 U10357 ( .A(n9007), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9011), .Z(
        P1_U3563) );
  MUX2_X1 U10358 ( .A(n9008), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9011), .Z(
        P1_U3562) );
  MUX2_X1 U10359 ( .A(n9743), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9011), .Z(
        P1_U3561) );
  MUX2_X1 U10360 ( .A(n9009), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9011), .Z(
        P1_U3560) );
  MUX2_X1 U10361 ( .A(n9010), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9011), .Z(
        P1_U3559) );
  MUX2_X1 U10362 ( .A(n8967), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9011), .Z(
        P1_U3558) );
  MUX2_X1 U10363 ( .A(n4932), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9011), .Z(
        P1_U3557) );
  MUX2_X1 U10364 ( .A(n5562), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9011), .Z(
        P1_U3556) );
  MUX2_X1 U10365 ( .A(n5553), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9011), .Z(
        P1_U3555) );
  OAI21_X1 U10366 ( .B1(n9014), .B2(n9013), .A(n9012), .ZN(n9016) );
  INV_X1 U10367 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9015) );
  OAI22_X1 U10368 ( .A1(n9708), .A2(n9016), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9015), .ZN(n9017) );
  AOI21_X1 U10369 ( .B1(n9671), .B2(n9018), .A(n9017), .ZN(n9027) );
  NAND2_X1 U10370 ( .A1(n9603), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n9026) );
  INV_X1 U10371 ( .A(n9019), .ZN(n9022) );
  INV_X1 U10372 ( .A(n9020), .ZN(n9021) );
  NAND2_X1 U10373 ( .A1(n9022), .A2(n9021), .ZN(n9023) );
  NAND3_X1 U10374 ( .A1(n9698), .A2(n9024), .A3(n9023), .ZN(n9025) );
  NAND4_X1 U10375 ( .A1(n9028), .A2(n9027), .A3(n9026), .A4(n9025), .ZN(
        P1_U3243) );
  XNOR2_X1 U10376 ( .A(n9634), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n9630) );
  NOR2_X1 U10377 ( .A1(n9031), .A2(n9043), .ZN(n9032) );
  NOR2_X1 U10378 ( .A1(n7214), .A2(n9643), .ZN(n9642) );
  INV_X1 U10379 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9655) );
  NAND2_X1 U10380 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9672), .ZN(n9034) );
  OAI21_X1 U10381 ( .B1(n9672), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9034), .ZN(
        n9667) );
  NOR2_X1 U10382 ( .A1(n9668), .A2(n9667), .ZN(n9666) );
  AOI21_X1 U10383 ( .B1(n9672), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9666), .ZN(
        n9680) );
  NAND2_X1 U10384 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9039), .ZN(n9035) );
  OAI21_X1 U10385 ( .B1(n9039), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9035), .ZN(
        n9681) );
  NOR2_X1 U10386 ( .A1(n9680), .A2(n9681), .ZN(n9679) );
  INV_X1 U10387 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9036) );
  MUX2_X1 U10388 ( .A(n9036), .B(P1_REG2_REG_18__SCAN_IN), .S(n9038), .Z(n9696) );
  INV_X1 U10389 ( .A(n9055), .ZN(n9053) );
  INV_X1 U10390 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9049) );
  XNOR2_X1 U10391 ( .A(n9038), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9706) );
  INV_X1 U10392 ( .A(n9039), .ZN(n9685) );
  INV_X1 U10393 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9048) );
  XNOR2_X1 U10394 ( .A(n9685), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9690) );
  INV_X1 U10395 ( .A(n9672), .ZN(n9047) );
  MUX2_X1 U10396 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9519), .S(n9672), .Z(n9674) );
  INV_X1 U10397 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9531) );
  INV_X1 U10398 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9538) );
  INV_X1 U10399 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9544) );
  AOI21_X1 U10400 ( .B1(n9544), .B2(n9041), .A(n9040), .ZN(n9637) );
  MUX2_X1 U10401 ( .A(n9538), .B(P1_REG1_REG_13__SCAN_IN), .S(n9634), .Z(n9636) );
  NOR2_X1 U10402 ( .A1(n9637), .A2(n9636), .ZN(n9635) );
  AOI21_X1 U10403 ( .B1(n9538), .B2(n9042), .A(n9635), .ZN(n9649) );
  MUX2_X1 U10404 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9531), .S(n9043), .Z(n9648) );
  NOR2_X1 U10405 ( .A1(n9649), .A2(n9648), .ZN(n9647) );
  AOI21_X1 U10406 ( .B1(n9043), .B2(n9531), .A(n9647), .ZN(n9044) );
  NAND2_X1 U10407 ( .A1(n9659), .A2(n9044), .ZN(n9046) );
  XNOR2_X1 U10408 ( .A(n9045), .B(n9044), .ZN(n9661) );
  NAND2_X1 U10409 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9661), .ZN(n9660) );
  NAND2_X1 U10410 ( .A1(n9046), .A2(n9660), .ZN(n9675) );
  NAND2_X1 U10411 ( .A1(n9674), .A2(n9675), .ZN(n9673) );
  OAI21_X1 U10412 ( .B1(n9047), .B2(n9519), .A(n9673), .ZN(n9689) );
  NAND2_X1 U10413 ( .A1(n9690), .A2(n9689), .ZN(n9687) );
  OAI21_X1 U10414 ( .B1(n9685), .B2(n9048), .A(n9687), .ZN(n9705) );
  NOR2_X1 U10415 ( .A1(n9706), .A2(n9705), .ZN(n9704) );
  AOI21_X1 U10416 ( .B1(n9701), .B2(n9049), .A(n9704), .ZN(n9050) );
  XOR2_X1 U10417 ( .A(n9050), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9054) );
  OAI21_X1 U10418 ( .B1(n9054), .B2(n9708), .A(n9702), .ZN(n9051) );
  AOI21_X1 U10419 ( .B1(n9053), .B2(n9052), .A(n9051), .ZN(n9057) );
  AOI22_X1 U10420 ( .A1(n9055), .A2(n9698), .B1(n9688), .B2(n9054), .ZN(n9056)
         );
  MUX2_X1 U10421 ( .A(n9057), .B(n9056), .S(n9136), .Z(n9059) );
  OAI211_X1 U10422 ( .C1(n4891), .C2(n9711), .A(n9059), .B(n9058), .ZN(
        P1_U3260) );
  XNOR2_X1 U10423 ( .A(n9064), .B(n9293), .ZN(n9292) );
  NAND2_X1 U10424 ( .A1(n9292), .A2(n9720), .ZN(n9063) );
  NAND2_X1 U10425 ( .A1(n9061), .A2(n9060), .ZN(n9508) );
  NOR2_X1 U10426 ( .A1(n9755), .A2(n9508), .ZN(n9068) );
  AOI21_X1 U10427 ( .B1(n9755), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9068), .ZN(
        n9062) );
  OAI211_X1 U10428 ( .C1(n9293), .C2(n9765), .A(n9063), .B(n9062), .ZN(
        P1_U3261) );
  OAI21_X1 U10429 ( .B1(n9065), .B2(n9066), .A(n9064), .ZN(n9509) );
  NOR2_X1 U10430 ( .A1(n9066), .A2(n9765), .ZN(n9067) );
  AOI211_X1 U10431 ( .C1(n9755), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9068), .B(
        n9067), .ZN(n9069) );
  OAI21_X1 U10432 ( .B1(n9509), .B2(n9762), .A(n9069), .ZN(P1_U3262) );
  OAI21_X1 U10433 ( .B1(n9072), .B2(n9071), .A(n9070), .ZN(n9306) );
  INV_X1 U10434 ( .A(n9073), .ZN(n9074) );
  AOI21_X1 U10435 ( .B1(n9302), .B2(n9084), .A(n9074), .ZN(n9303) );
  AOI22_X1 U10436 ( .A1(n9075), .A2(n9783), .B1(n9755), .B2(
        P1_REG2_REG_28__SCAN_IN), .ZN(n9076) );
  OAI21_X1 U10437 ( .B1(n4511), .B2(n9765), .A(n9076), .ZN(n9082) );
  OAI21_X1 U10438 ( .B1(n9079), .B2(n9078), .A(n9077), .ZN(n9081) );
  XOR2_X1 U10439 ( .A(n9092), .B(n9083), .Z(n9311) );
  INV_X1 U10440 ( .A(n9100), .ZN(n9086) );
  INV_X1 U10441 ( .A(n9084), .ZN(n9085) );
  AOI21_X1 U10442 ( .B1(n9307), .B2(n9086), .A(n9085), .ZN(n9308) );
  AOI22_X1 U10443 ( .A1(n9087), .A2(n9783), .B1(n9755), .B2(
        P1_REG2_REG_27__SCAN_IN), .ZN(n9088) );
  OAI21_X1 U10444 ( .B1(n9089), .B2(n9765), .A(n9088), .ZN(n9096) );
  NOR2_X1 U10445 ( .A1(n9090), .A2(n9772), .ZN(n9094) );
  AOI211_X1 U10446 ( .C1(n9092), .C2(n9091), .A(n9749), .B(n4354), .ZN(n9093)
         );
  NOR2_X1 U10447 ( .A1(n9310), .A2(n9755), .ZN(n9095) );
  AOI211_X1 U10448 ( .C1(n9720), .C2(n9308), .A(n9096), .B(n9095), .ZN(n9097)
         );
  OAI21_X1 U10449 ( .B1(n9311), .B2(n9290), .A(n9097), .ZN(P1_U3264) );
  XNOR2_X1 U10450 ( .A(n9099), .B(n9098), .ZN(n9316) );
  INV_X1 U10451 ( .A(n9116), .ZN(n9101) );
  AOI211_X1 U10452 ( .C1(n9313), .C2(n9101), .A(n9851), .B(n9100), .ZN(n9312)
         );
  AOI22_X1 U10453 ( .A1(n9755), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9102), .B2(
        n9783), .ZN(n9103) );
  OAI21_X1 U10454 ( .B1(n9104), .B2(n9765), .A(n9103), .ZN(n9113) );
  INV_X1 U10455 ( .A(n9105), .ZN(n9106) );
  NOR2_X1 U10456 ( .A1(n9107), .A2(n9106), .ZN(n9109) );
  XNOR2_X1 U10457 ( .A(n9109), .B(n9108), .ZN(n9111) );
  AOI222_X1 U10458 ( .A1(n9770), .A2(n9111), .B1(n9110), .B2(n9742), .C1(n9131), .C2(n9489), .ZN(n9315) );
  NOR2_X1 U10459 ( .A1(n9315), .A2(n9755), .ZN(n9112) );
  AOI211_X1 U10460 ( .C1(n9312), .C2(n9235), .A(n9113), .B(n9112), .ZN(n9114)
         );
  OAI21_X1 U10461 ( .B1(n9316), .B2(n9290), .A(n9114), .ZN(P1_U3265) );
  XOR2_X1 U10462 ( .A(n9121), .B(n9115), .Z(n9321) );
  AOI21_X1 U10463 ( .B1(n9317), .B2(n9133), .A(n9116), .ZN(n9318) );
  AOI22_X1 U10464 ( .A1(n9755), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9117), .B2(
        n9783), .ZN(n9118) );
  OAI21_X1 U10465 ( .B1(n9119), .B2(n9765), .A(n9118), .ZN(n9125) );
  XOR2_X1 U10466 ( .A(n9120), .B(n9121), .Z(n9123) );
  AOI222_X1 U10467 ( .A1(n9770), .A2(n9123), .B1(n9122), .B2(n9742), .C1(n9154), .C2(n9489), .ZN(n9320) );
  NOR2_X1 U10468 ( .A1(n9320), .A2(n9755), .ZN(n9124) );
  AOI211_X1 U10469 ( .C1(n9318), .C2(n9720), .A(n9125), .B(n9124), .ZN(n9126)
         );
  OAI21_X1 U10470 ( .B1(n9321), .B2(n9290), .A(n9126), .ZN(P1_U3266) );
  XNOR2_X1 U10471 ( .A(n9127), .B(n9129), .ZN(n9326) );
  NOR2_X1 U10472 ( .A1(n9128), .A2(n9765), .ZN(n9139) );
  XNOR2_X1 U10473 ( .A(n9130), .B(n9129), .ZN(n9132) );
  AOI222_X1 U10474 ( .A1(n9770), .A2(n9132), .B1(n9131), .B2(n9742), .C1(n9167), .C2(n9489), .ZN(n9325) );
  INV_X1 U10475 ( .A(n9133), .ZN(n9134) );
  AOI211_X1 U10476 ( .C1(n9323), .C2(n9142), .A(n9851), .B(n9134), .ZN(n9322)
         );
  AOI22_X1 U10477 ( .A1(n9322), .A2(n9136), .B1(n9783), .B2(n9135), .ZN(n9137)
         );
  AOI21_X1 U10478 ( .B1(n9325), .B2(n9137), .A(n9755), .ZN(n9138) );
  AOI211_X1 U10479 ( .C1(n9755), .C2(P1_REG2_REG_24__SCAN_IN), .A(n9139), .B(
        n9138), .ZN(n9140) );
  OAI21_X1 U10480 ( .B1(n9326), .B2(n9290), .A(n9140), .ZN(P1_U3267) );
  XNOR2_X1 U10481 ( .A(n9141), .B(n9149), .ZN(n9331) );
  INV_X1 U10482 ( .A(n9161), .ZN(n9144) );
  INV_X1 U10483 ( .A(n9142), .ZN(n9143) );
  AOI21_X1 U10484 ( .B1(n9327), .B2(n9144), .A(n9143), .ZN(n9328) );
  AOI22_X1 U10485 ( .A1(n9755), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9145), .B2(
        n9783), .ZN(n9146) );
  OAI21_X1 U10486 ( .B1(n9147), .B2(n9765), .A(n9146), .ZN(n9158) );
  INV_X1 U10487 ( .A(n9148), .ZN(n9151) );
  OAI21_X1 U10488 ( .B1(n9151), .B2(n9150), .A(n9149), .ZN(n9153) );
  NAND3_X1 U10489 ( .A1(n9153), .A2(n9770), .A3(n9152), .ZN(n9156) );
  AOI22_X1 U10490 ( .A1(n9489), .A2(n9182), .B1(n9154), .B2(n9742), .ZN(n9155)
         );
  AND2_X1 U10491 ( .A1(n9156), .A2(n9155), .ZN(n9330) );
  NOR2_X1 U10492 ( .A1(n9330), .A2(n9755), .ZN(n9157) );
  AOI211_X1 U10493 ( .C1(n9328), .C2(n9720), .A(n9158), .B(n9157), .ZN(n9159)
         );
  OAI21_X1 U10494 ( .B1(n9331), .B2(n9290), .A(n9159), .ZN(P1_U3268) );
  XOR2_X1 U10495 ( .A(n9160), .B(n9166), .Z(n9336) );
  AOI21_X1 U10496 ( .B1(n9332), .B2(n9186), .A(n9161), .ZN(n9333) );
  AOI22_X1 U10497 ( .A1(n9755), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9162), .B2(
        n9783), .ZN(n9163) );
  OAI21_X1 U10498 ( .B1(n9164), .B2(n9765), .A(n9163), .ZN(n9170) );
  OAI21_X1 U10499 ( .B1(n9166), .B2(n9165), .A(n9148), .ZN(n9168) );
  AOI222_X1 U10500 ( .A1(n9770), .A2(n9168), .B1(n9167), .B2(n9742), .C1(n9201), .C2(n9489), .ZN(n9335) );
  NOR2_X1 U10501 ( .A1(n9335), .A2(n9755), .ZN(n9169) );
  AOI211_X1 U10502 ( .C1(n9333), .C2(n9720), .A(n9170), .B(n9169), .ZN(n9171)
         );
  OAI21_X1 U10503 ( .B1(n9336), .B2(n9290), .A(n9171), .ZN(P1_U3269) );
  NAND2_X1 U10504 ( .A1(n9174), .A2(n9173), .ZN(n9175) );
  NAND2_X1 U10505 ( .A1(n9172), .A2(n9175), .ZN(n9337) );
  NAND2_X1 U10506 ( .A1(n9177), .A2(n9176), .ZN(n9178) );
  NAND2_X1 U10507 ( .A1(n9178), .A2(n5325), .ZN(n9180) );
  NAND2_X1 U10508 ( .A1(n9180), .A2(n9179), .ZN(n9181) );
  NAND2_X1 U10509 ( .A1(n9181), .A2(n9770), .ZN(n9184) );
  AOI22_X1 U10510 ( .A1(n9742), .A2(n9182), .B1(n9216), .B2(n9489), .ZN(n9183)
         );
  NAND2_X1 U10511 ( .A1(n9184), .A2(n9183), .ZN(n9341) );
  AOI21_X1 U10512 ( .B1(n9194), .B2(n9185), .A(n9851), .ZN(n9187) );
  NAND2_X1 U10513 ( .A1(n9187), .A2(n9186), .ZN(n9338) );
  NOR2_X1 U10514 ( .A1(n9338), .A2(n9500), .ZN(n9191) );
  AOI22_X1 U10515 ( .A1(n9755), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9188), .B2(
        n9783), .ZN(n9189) );
  OAI21_X1 U10516 ( .B1(n9339), .B2(n9765), .A(n9189), .ZN(n9190) );
  AOI211_X1 U10517 ( .C1(n9341), .C2(n9779), .A(n9191), .B(n9190), .ZN(n9192)
         );
  OAI21_X1 U10518 ( .B1(n9337), .B2(n9290), .A(n9192), .ZN(P1_U3270) );
  XNOR2_X1 U10519 ( .A(n9193), .B(n9199), .ZN(n9348) );
  INV_X1 U10520 ( .A(n9194), .ZN(n9195) );
  AOI21_X1 U10521 ( .B1(n9344), .B2(n9207), .A(n9195), .ZN(n9345) );
  AOI22_X1 U10522 ( .A1(n9755), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9196), .B2(
        n9783), .ZN(n9197) );
  OAI21_X1 U10523 ( .B1(n9198), .B2(n9765), .A(n9197), .ZN(n9204) );
  XOR2_X1 U10524 ( .A(n9200), .B(n9199), .Z(n9202) );
  AOI222_X1 U10525 ( .A1(n9770), .A2(n9202), .B1(n9230), .B2(n9489), .C1(n9201), .C2(n9742), .ZN(n9347) );
  NOR2_X1 U10526 ( .A1(n9347), .A2(n9755), .ZN(n9203) );
  AOI211_X1 U10527 ( .C1(n9345), .C2(n9720), .A(n9204), .B(n9203), .ZN(n9205)
         );
  OAI21_X1 U10528 ( .B1(n9290), .B2(n9348), .A(n9205), .ZN(P1_U3271) );
  XOR2_X1 U10529 ( .A(n9206), .B(n9215), .Z(n9353) );
  INV_X1 U10530 ( .A(n9233), .ZN(n9209) );
  INV_X1 U10531 ( .A(n9207), .ZN(n9208) );
  AOI211_X1 U10532 ( .C1(n9350), .C2(n9209), .A(n9851), .B(n9208), .ZN(n9349)
         );
  AOI22_X1 U10533 ( .A1(n9755), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9210), .B2(
        n9783), .ZN(n9211) );
  OAI21_X1 U10534 ( .B1(n9212), .B2(n9765), .A(n9211), .ZN(n9219) );
  OAI21_X1 U10535 ( .B1(n9215), .B2(n9214), .A(n9213), .ZN(n9217) );
  AOI222_X1 U10536 ( .A1(n9770), .A2(n9217), .B1(n9248), .B2(n9489), .C1(n9216), .C2(n9742), .ZN(n9352) );
  NOR2_X1 U10537 ( .A1(n9352), .A2(n9755), .ZN(n9218) );
  AOI211_X1 U10538 ( .C1(n9349), .C2(n9235), .A(n9219), .B(n9218), .ZN(n9220)
         );
  OAI21_X1 U10539 ( .B1(n9353), .B2(n9290), .A(n9220), .ZN(P1_U3272) );
  INV_X1 U10540 ( .A(n9221), .ZN(n9224) );
  INV_X1 U10541 ( .A(n9222), .ZN(n9227) );
  OAI21_X1 U10542 ( .B1(n9224), .B2(n9227), .A(n9223), .ZN(n9358) );
  NAND2_X1 U10543 ( .A1(n9226), .A2(n9225), .ZN(n9228) );
  XNOR2_X1 U10544 ( .A(n9228), .B(n9227), .ZN(n9229) );
  NAND2_X1 U10545 ( .A1(n9229), .A2(n9770), .ZN(n9232) );
  AOI22_X1 U10546 ( .A1(n9742), .A2(n9230), .B1(n9261), .B2(n9489), .ZN(n9231)
         );
  NAND2_X1 U10547 ( .A1(n9232), .A2(n9231), .ZN(n9355) );
  INV_X1 U10548 ( .A(n9243), .ZN(n9234) );
  AOI211_X1 U10549 ( .C1(n9356), .C2(n9234), .A(n9851), .B(n9233), .ZN(n9354)
         );
  NAND2_X1 U10550 ( .A1(n9354), .A2(n9235), .ZN(n9238) );
  AOI22_X1 U10551 ( .A1(n9755), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9236), .B2(
        n9783), .ZN(n9237) );
  OAI211_X1 U10552 ( .C1(n9239), .C2(n9765), .A(n9238), .B(n9237), .ZN(n9240)
         );
  AOI21_X1 U10553 ( .B1(n9779), .B2(n9355), .A(n9240), .ZN(n9241) );
  OAI21_X1 U10554 ( .B1(n9358), .B2(n9290), .A(n9241), .ZN(P1_U3273) );
  XOR2_X1 U10555 ( .A(n9242), .B(n9247), .Z(n9363) );
  AOI21_X1 U10556 ( .B1(n9359), .B2(n4315), .A(n9243), .ZN(n9360) );
  AOI22_X1 U10557 ( .A1(n9755), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9244), .B2(
        n9783), .ZN(n9245) );
  OAI21_X1 U10558 ( .B1(n9246), .B2(n9765), .A(n9245), .ZN(n9251) );
  XOR2_X1 U10559 ( .A(n4397), .B(n9247), .Z(n9249) );
  AOI222_X1 U10560 ( .A1(n9770), .A2(n9249), .B1(n9248), .B2(n9742), .C1(n9276), .C2(n9489), .ZN(n9362) );
  NOR2_X1 U10561 ( .A1(n9362), .A2(n9755), .ZN(n9250) );
  AOI211_X1 U10562 ( .C1(n9360), .C2(n9720), .A(n9251), .B(n9250), .ZN(n9252)
         );
  OAI21_X1 U10563 ( .B1(n9290), .B2(n9363), .A(n9252), .ZN(P1_U3274) );
  XNOR2_X1 U10564 ( .A(n9254), .B(n9253), .ZN(n9518) );
  INV_X1 U10565 ( .A(n9518), .ZN(n9270) );
  NAND2_X1 U10566 ( .A1(n9257), .A2(n9256), .ZN(n9258) );
  NAND2_X1 U10567 ( .A1(n9259), .A2(n9258), .ZN(n9260) );
  NAND2_X1 U10568 ( .A1(n9260), .A2(n9770), .ZN(n9264) );
  AOI22_X1 U10569 ( .A1(n9489), .A2(n9262), .B1(n9261), .B2(n9742), .ZN(n9263)
         );
  NAND2_X1 U10570 ( .A1(n9264), .A2(n9263), .ZN(n9517) );
  AOI22_X1 U10571 ( .A1(n9755), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9265), .B2(
        n9783), .ZN(n9266) );
  OAI21_X1 U10572 ( .B1(n4499), .B2(n9765), .A(n9266), .ZN(n9268) );
  OAI211_X1 U10573 ( .C1(n4500), .C2(n4499), .A(n9828), .B(n4315), .ZN(n9515)
         );
  NOR2_X1 U10574 ( .A1(n9515), .A2(n9500), .ZN(n9267) );
  AOI211_X1 U10575 ( .C1(n9779), .C2(n9517), .A(n9268), .B(n9267), .ZN(n9269)
         );
  OAI21_X1 U10576 ( .B1(n9270), .B2(n9290), .A(n9269), .ZN(P1_U3275) );
  XNOR2_X1 U10577 ( .A(n9271), .B(n9272), .ZN(n9524) );
  INV_X1 U10578 ( .A(n9524), .ZN(n9291) );
  XNOR2_X1 U10579 ( .A(n9273), .B(n9272), .ZN(n9274) );
  NAND2_X1 U10580 ( .A1(n9274), .A2(n9770), .ZN(n9278) );
  AOI22_X1 U10581 ( .A1(n9276), .A2(n9742), .B1(n9489), .B2(n9275), .ZN(n9277)
         );
  NAND2_X1 U10582 ( .A1(n9278), .A2(n9277), .ZN(n9523) );
  OR2_X1 U10583 ( .A1(n9279), .A2(n9520), .ZN(n9280) );
  NAND2_X1 U10584 ( .A1(n9281), .A2(n9280), .ZN(n9521) );
  INV_X1 U10585 ( .A(n9282), .ZN(n9284) );
  OAI22_X1 U10586 ( .A1(n9779), .A2(n9655), .B1(n9284), .B2(n9283), .ZN(n9285)
         );
  AOI21_X1 U10587 ( .B1(n9286), .B2(n9494), .A(n9285), .ZN(n9287) );
  OAI21_X1 U10588 ( .B1(n9521), .B2(n9762), .A(n9287), .ZN(n9288) );
  AOI21_X1 U10589 ( .B1(n9523), .B2(n9779), .A(n9288), .ZN(n9289) );
  OAI21_X1 U10590 ( .B1(n9291), .B2(n9290), .A(n9289), .ZN(P1_U3276) );
  MUX2_X1 U10591 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9364), .S(n9879), .Z(
        P1_U3554) );
  AOI22_X1 U10592 ( .A1(n9298), .A2(n9828), .B1(n9827), .B2(n9297), .ZN(n9299)
         );
  OAI211_X1 U10593 ( .C1(n9301), .C2(n9514), .A(n9300), .B(n9299), .ZN(n9365)
         );
  MUX2_X1 U10594 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9365), .S(n9879), .Z(
        P1_U3552) );
  AOI22_X1 U10595 ( .A1(n9303), .A2(n9828), .B1(n9827), .B2(n9302), .ZN(n9304)
         );
  OAI211_X1 U10596 ( .C1(n9306), .C2(n9514), .A(n9305), .B(n9304), .ZN(n9366)
         );
  MUX2_X1 U10597 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9366), .S(n9879), .Z(
        P1_U3551) );
  AOI22_X1 U10598 ( .A1(n9308), .A2(n9828), .B1(n9827), .B2(n9307), .ZN(n9309)
         );
  OAI211_X1 U10599 ( .C1(n9311), .C2(n9514), .A(n9310), .B(n9309), .ZN(n9367)
         );
  MUX2_X1 U10600 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9367), .S(n9879), .Z(
        P1_U3550) );
  AOI21_X1 U10601 ( .B1(n9827), .B2(n9313), .A(n9312), .ZN(n9314) );
  OAI211_X1 U10602 ( .C1(n9316), .C2(n9514), .A(n9315), .B(n9314), .ZN(n9368)
         );
  MUX2_X1 U10603 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9368), .S(n9879), .Z(
        P1_U3549) );
  AOI22_X1 U10604 ( .A1(n9318), .A2(n9828), .B1(n9827), .B2(n9317), .ZN(n9319)
         );
  OAI211_X1 U10605 ( .C1(n9321), .C2(n9514), .A(n9320), .B(n9319), .ZN(n9369)
         );
  MUX2_X1 U10606 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9369), .S(n9879), .Z(
        P1_U3548) );
  AOI21_X1 U10607 ( .B1(n9827), .B2(n9323), .A(n9322), .ZN(n9324) );
  OAI211_X1 U10608 ( .C1(n9326), .C2(n9514), .A(n9325), .B(n9324), .ZN(n9370)
         );
  MUX2_X1 U10609 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9370), .S(n9879), .Z(
        P1_U3547) );
  AOI22_X1 U10610 ( .A1(n9328), .A2(n9828), .B1(n9827), .B2(n9327), .ZN(n9329)
         );
  OAI211_X1 U10611 ( .C1(n9331), .C2(n9514), .A(n9330), .B(n9329), .ZN(n9371)
         );
  MUX2_X1 U10612 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9371), .S(n9879), .Z(
        P1_U3546) );
  AOI22_X1 U10613 ( .A1(n9333), .A2(n9828), .B1(n9827), .B2(n9332), .ZN(n9334)
         );
  OAI211_X1 U10614 ( .C1(n9336), .C2(n9514), .A(n9335), .B(n9334), .ZN(n9372)
         );
  MUX2_X1 U10615 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9372), .S(n9879), .Z(
        P1_U3545) );
  OR2_X1 U10616 ( .A1(n9337), .A2(n9514), .ZN(n9343) );
  OAI21_X1 U10617 ( .B1(n9339), .B2(n9849), .A(n9338), .ZN(n9340) );
  NOR2_X1 U10618 ( .A1(n9341), .A2(n9340), .ZN(n9342) );
  NAND2_X1 U10619 ( .A1(n9343), .A2(n9342), .ZN(n9373) );
  MUX2_X1 U10620 ( .A(n9373), .B(P1_REG1_REG_21__SCAN_IN), .S(n9876), .Z(
        P1_U3544) );
  AOI22_X1 U10621 ( .A1(n9345), .A2(n9828), .B1(n9827), .B2(n9344), .ZN(n9346)
         );
  OAI211_X1 U10622 ( .C1(n9348), .C2(n9514), .A(n9347), .B(n9346), .ZN(n9374)
         );
  MUX2_X1 U10623 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9374), .S(n9879), .Z(
        P1_U3543) );
  AOI21_X1 U10624 ( .B1(n9827), .B2(n9350), .A(n9349), .ZN(n9351) );
  OAI211_X1 U10625 ( .C1(n9353), .C2(n9514), .A(n9352), .B(n9351), .ZN(n9375)
         );
  MUX2_X1 U10626 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9375), .S(n9879), .Z(
        P1_U3542) );
  AOI211_X1 U10627 ( .C1(n9827), .C2(n9356), .A(n9355), .B(n9354), .ZN(n9357)
         );
  OAI21_X1 U10628 ( .B1(n9358), .B2(n9514), .A(n9357), .ZN(n9376) );
  MUX2_X1 U10629 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9376), .S(n9879), .Z(
        P1_U3541) );
  AOI22_X1 U10630 ( .A1(n9360), .A2(n9828), .B1(n9827), .B2(n9359), .ZN(n9361)
         );
  OAI211_X1 U10631 ( .C1(n9363), .C2(n9514), .A(n9362), .B(n9361), .ZN(n9377)
         );
  MUX2_X1 U10632 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9377), .S(n9879), .Z(
        P1_U3540) );
  MUX2_X1 U10633 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9364), .S(n9859), .Z(
        P1_U3522) );
  MUX2_X1 U10634 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9365), .S(n9859), .Z(
        P1_U3520) );
  MUX2_X1 U10635 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9366), .S(n9859), .Z(
        P1_U3519) );
  MUX2_X1 U10636 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9367), .S(n9859), .Z(
        P1_U3518) );
  MUX2_X1 U10637 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9368), .S(n9859), .Z(
        P1_U3517) );
  MUX2_X1 U10638 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9369), .S(n9859), .Z(
        P1_U3516) );
  MUX2_X1 U10639 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9370), .S(n9859), .Z(
        P1_U3515) );
  MUX2_X1 U10640 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9371), .S(n9859), .Z(
        P1_U3514) );
  MUX2_X1 U10641 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9372), .S(n9859), .Z(
        P1_U3513) );
  MUX2_X1 U10642 ( .A(n9373), .B(P1_REG0_REG_21__SCAN_IN), .S(n9857), .Z(
        P1_U3512) );
  MUX2_X1 U10643 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9374), .S(n9859), .Z(
        P1_U3511) );
  MUX2_X1 U10644 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9375), .S(n9859), .Z(
        P1_U3510) );
  MUX2_X1 U10645 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9376), .S(n9859), .Z(
        P1_U3508) );
  MUX2_X1 U10646 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9377), .S(n9859), .Z(
        P1_U3505) );
  INV_X1 U10647 ( .A(n9378), .ZN(n9379) );
  MUX2_X1 U10648 ( .A(n9380), .B(P1_D_REG_0__SCAN_IN), .S(n9789), .Z(P1_U3440)
         );
  NOR4_X1 U10649 ( .A1(n4882), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n4878), .ZN(n9381) );
  AOI21_X1 U10650 ( .B1(n9390), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9381), .ZN(
        n9382) );
  OAI21_X1 U10651 ( .B1(n9383), .B2(n9397), .A(n9382), .ZN(P1_U3322) );
  OAI222_X1 U10652 ( .A1(n9397), .A2(n9386), .B1(n9385), .B2(P1_U3084), .C1(
        n9384), .C2(n9401), .ZN(P1_U3324) );
  AOI21_X1 U10653 ( .B1(n9390), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n9387), .ZN(
        n9388) );
  OAI21_X1 U10654 ( .B1(n9389), .B2(n9397), .A(n9388), .ZN(P1_U3325) );
  NAND2_X1 U10655 ( .A1(n9390), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9391) );
  OAI211_X1 U10656 ( .C1(n9393), .C2(n9397), .A(n9392), .B(n9391), .ZN(
        P1_U3326) );
  OAI222_X1 U10657 ( .A1(n9397), .A2(n9396), .B1(P1_U3084), .B2(n9395), .C1(
        n9394), .C2(n9401), .ZN(P1_U3327) );
  OAI222_X1 U10658 ( .A1(n9401), .A2(n9400), .B1(n9397), .B2(n9399), .C1(n9398), .C2(P1_U3084), .ZN(P1_U3328) );
  MUX2_X1 U10659 ( .A(n9402), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10660 ( .A1(n9898), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n9413) );
  NAND2_X1 U10661 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9405) );
  AOI211_X1 U10662 ( .C1(n9405), .C2(n9404), .A(n9403), .B(n9414), .ZN(n9406)
         );
  AOI21_X1 U10663 ( .B1(n9895), .B2(n9407), .A(n9406), .ZN(n9412) );
  INV_X1 U10664 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10005) );
  NOR2_X1 U10665 ( .A1(n9901), .A2(n10005), .ZN(n9410) );
  OAI211_X1 U10666 ( .C1(n9410), .C2(n9409), .A(n9892), .B(n9408), .ZN(n9411)
         );
  NAND3_X1 U10667 ( .A1(n9413), .A2(n9412), .A3(n9411), .ZN(P2_U3246) );
  AOI22_X1 U10668 ( .A1(n9898), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9425) );
  AOI211_X1 U10669 ( .C1(n9417), .C2(n9416), .A(n9415), .B(n9414), .ZN(n9418)
         );
  AOI21_X1 U10670 ( .B1(n9895), .B2(n9419), .A(n9418), .ZN(n9424) );
  OAI211_X1 U10671 ( .C1(n9422), .C2(n9421), .A(n9892), .B(n9420), .ZN(n9423)
         );
  NAND3_X1 U10672 ( .A1(n9425), .A2(n9424), .A3(n9423), .ZN(P2_U3247) );
  INV_X1 U10673 ( .A(n9832), .ZN(n9847) );
  OAI21_X1 U10674 ( .B1(n9427), .B2(n9849), .A(n9426), .ZN(n9429) );
  AOI211_X1 U10675 ( .C1(n9847), .C2(n9430), .A(n9429), .B(n9428), .ZN(n9433)
         );
  INV_X1 U10676 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9431) );
  AOI22_X1 U10677 ( .A1(n9859), .A2(n9433), .B1(n9431), .B2(n9857), .ZN(
        P1_U3484) );
  AOI22_X1 U10678 ( .A1(n9879), .A2(n9433), .B1(n9432), .B2(n9876), .ZN(
        P1_U3533) );
  INV_X1 U10679 ( .A(n9434), .ZN(n9442) );
  AOI22_X1 U10680 ( .A1(n4305), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n9436), .B2(
        n9435), .ZN(n9437) );
  OAI21_X1 U10681 ( .B1(n9439), .B2(n9438), .A(n9437), .ZN(n9440) );
  AOI21_X1 U10682 ( .B1(n9442), .B2(n9441), .A(n9440), .ZN(n9451) );
  INV_X1 U10683 ( .A(n9443), .ZN(n9445) );
  NOR3_X1 U10684 ( .A1(n9446), .A2(n9445), .A3(n9444), .ZN(n9447) );
  AOI21_X1 U10685 ( .B1(n9449), .B2(n9448), .A(n9447), .ZN(n9450) );
  NAND2_X1 U10686 ( .A1(n9451), .A2(n9450), .ZN(P2_U3280) );
  OAI21_X1 U10687 ( .B1(n9453), .B2(n9994), .A(n9452), .ZN(n9454) );
  AOI21_X1 U10688 ( .B1(n9456), .B2(n9455), .A(n9454), .ZN(n9479) );
  INV_X1 U10689 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9457) );
  AOI22_X1 U10690 ( .A1(n10023), .A2(n9479), .B1(n9457), .B2(n10021), .ZN(
        P2_U3550) );
  OAI22_X1 U10691 ( .A1(n9459), .A2(n9996), .B1(n9458), .B2(n9994), .ZN(n9460)
         );
  AOI211_X1 U10692 ( .C1(n9462), .C2(n10001), .A(n9461), .B(n9460), .ZN(n9481)
         );
  INV_X1 U10693 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9463) );
  AOI22_X1 U10694 ( .A1(n10023), .A2(n9481), .B1(n9463), .B2(n10021), .ZN(
        P2_U3535) );
  INV_X1 U10695 ( .A(n9464), .ZN(n9469) );
  OAI22_X1 U10696 ( .A1(n9466), .A2(n9996), .B1(n9465), .B2(n9994), .ZN(n9467)
         );
  AOI211_X1 U10697 ( .C1(n9469), .C2(n10001), .A(n9468), .B(n9467), .ZN(n9483)
         );
  AOI22_X1 U10698 ( .A1(n10023), .A2(n9483), .B1(n9470), .B2(n10021), .ZN(
        P2_U3534) );
  INV_X1 U10699 ( .A(n9471), .ZN(n9985) );
  INV_X1 U10700 ( .A(n9472), .ZN(n9476) );
  OAI22_X1 U10701 ( .A1(n9473), .A2(n9996), .B1(n4535), .B2(n9994), .ZN(n9475)
         );
  AOI211_X1 U10702 ( .C1(n9985), .C2(n9476), .A(n9475), .B(n9474), .ZN(n9485)
         );
  AOI22_X1 U10703 ( .A1(n10023), .A2(n9485), .B1(n9477), .B2(n10021), .ZN(
        P2_U3533) );
  INV_X1 U10704 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9478) );
  AOI22_X1 U10705 ( .A1(n10004), .A2(n9479), .B1(n9478), .B2(n10002), .ZN(
        P2_U3518) );
  INV_X1 U10706 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9480) );
  AOI22_X1 U10707 ( .A1(n10004), .A2(n9481), .B1(n9480), .B2(n10002), .ZN(
        P2_U3496) );
  INV_X1 U10708 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9482) );
  AOI22_X1 U10709 ( .A1(n10004), .A2(n9483), .B1(n9482), .B2(n10002), .ZN(
        P2_U3493) );
  INV_X1 U10710 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9484) );
  AOI22_X1 U10711 ( .A1(n10004), .A2(n9485), .B1(n9484), .B2(n10002), .ZN(
        P2_U3490) );
  NAND2_X1 U10712 ( .A1(n9487), .A2(n9486), .ZN(n9488) );
  XNOR2_X1 U10713 ( .A(n9488), .B(n9499), .ZN(n9492) );
  AOI222_X1 U10714 ( .A1(n9770), .A2(n9492), .B1(n9491), .B2(n9742), .C1(n9490), .C2(n9489), .ZN(n9540) );
  AOI222_X1 U10715 ( .A1(n9495), .A2(n9494), .B1(n9493), .B2(n9783), .C1(
        P1_REG2_REG_12__SCAN_IN), .C2(n9755), .ZN(n9507) );
  INV_X1 U10716 ( .A(n9497), .ZN(n9498) );
  AOI21_X1 U10717 ( .B1(n9499), .B2(n9496), .A(n9498), .ZN(n9543) );
  INV_X1 U10718 ( .A(n9501), .ZN(n9503) );
  OAI211_X1 U10719 ( .C1(n9503), .C2(n9541), .A(n9828), .B(n9502), .ZN(n9539)
         );
  INV_X1 U10720 ( .A(n9539), .ZN(n9504) );
  AOI22_X1 U10721 ( .A1(n9543), .A2(n9505), .B1(n9235), .B2(n9504), .ZN(n9506)
         );
  OAI211_X1 U10722 ( .C1(n9755), .C2(n9540), .A(n9507), .B(n9506), .ZN(
        P1_U3279) );
  INV_X1 U10723 ( .A(n9508), .ZN(n9511) );
  NOR2_X1 U10724 ( .A1(n9509), .A2(n9851), .ZN(n9510) );
  INV_X1 U10725 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9513) );
  AOI22_X1 U10726 ( .A1(n9879), .A2(n9552), .B1(n9513), .B2(n9876), .ZN(
        P1_U3553) );
  OAI21_X1 U10727 ( .B1(n4499), .B2(n9849), .A(n9515), .ZN(n9516) );
  AOI211_X1 U10728 ( .C1(n9518), .C2(n9855), .A(n9517), .B(n9516), .ZN(n9554)
         );
  AOI22_X1 U10729 ( .A1(n9879), .A2(n9554), .B1(n9519), .B2(n9876), .ZN(
        P1_U3539) );
  OAI22_X1 U10730 ( .A1(n9521), .A2(n9851), .B1(n9520), .B2(n9849), .ZN(n9522)
         );
  AOI211_X1 U10731 ( .C1(n9524), .C2(n9855), .A(n9523), .B(n9522), .ZN(n9556)
         );
  INV_X1 U10732 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9525) );
  AOI22_X1 U10733 ( .A1(n9879), .A2(n9556), .B1(n9525), .B2(n9876), .ZN(
        P1_U3538) );
  OAI21_X1 U10734 ( .B1(n9527), .B2(n9849), .A(n9526), .ZN(n9528) );
  AOI211_X1 U10735 ( .C1(n9530), .C2(n9855), .A(n9529), .B(n9528), .ZN(n9558)
         );
  AOI22_X1 U10736 ( .A1(n9879), .A2(n9558), .B1(n9531), .B2(n9876), .ZN(
        P1_U3537) );
  OAI22_X1 U10737 ( .A1(n9533), .A2(n9851), .B1(n9532), .B2(n9849), .ZN(n9534)
         );
  AOI21_X1 U10738 ( .B1(n9535), .B2(n9847), .A(n9534), .ZN(n9536) );
  AND2_X1 U10739 ( .A1(n9537), .A2(n9536), .ZN(n9560) );
  AOI22_X1 U10740 ( .A1(n9879), .A2(n9560), .B1(n9538), .B2(n9876), .ZN(
        P1_U3536) );
  OAI211_X1 U10741 ( .C1(n9541), .C2(n9849), .A(n9540), .B(n9539), .ZN(n9542)
         );
  AOI21_X1 U10742 ( .B1(n9543), .B2(n9855), .A(n9542), .ZN(n9562) );
  AOI22_X1 U10743 ( .A1(n9879), .A2(n9562), .B1(n9544), .B2(n9876), .ZN(
        P1_U3535) );
  OAI22_X1 U10744 ( .A1(n9546), .A2(n9851), .B1(n9545), .B2(n9849), .ZN(n9548)
         );
  AOI211_X1 U10745 ( .C1(n9847), .C2(n9549), .A(n9548), .B(n9547), .ZN(n9564)
         );
  AOI22_X1 U10746 ( .A1(n9879), .A2(n9564), .B1(n9550), .B2(n9876), .ZN(
        P1_U3534) );
  INV_X1 U10747 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9551) );
  AOI22_X1 U10748 ( .A1(n9859), .A2(n9552), .B1(n9551), .B2(n9857), .ZN(
        P1_U3521) );
  INV_X1 U10749 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9553) );
  AOI22_X1 U10750 ( .A1(n9859), .A2(n9554), .B1(n9553), .B2(n9857), .ZN(
        P1_U3502) );
  INV_X1 U10751 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9555) );
  AOI22_X1 U10752 ( .A1(n9859), .A2(n9556), .B1(n9555), .B2(n9857), .ZN(
        P1_U3499) );
  INV_X1 U10753 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9557) );
  AOI22_X1 U10754 ( .A1(n9859), .A2(n9558), .B1(n9557), .B2(n9857), .ZN(
        P1_U3496) );
  INV_X1 U10755 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9559) );
  AOI22_X1 U10756 ( .A1(n9859), .A2(n9560), .B1(n9559), .B2(n9857), .ZN(
        P1_U3493) );
  INV_X1 U10757 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9561) );
  AOI22_X1 U10758 ( .A1(n9859), .A2(n9562), .B1(n9561), .B2(n9857), .ZN(
        P1_U3490) );
  INV_X1 U10759 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9563) );
  AOI22_X1 U10760 ( .A1(n9859), .A2(n9564), .B1(n9563), .B2(n9857), .ZN(
        P1_U3487) );
  XNOR2_X1 U10761 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10762 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10763 ( .A(n9565), .ZN(n9572) );
  OAI21_X1 U10764 ( .B1(n9567), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9566), .ZN(
        n9571) );
  INV_X1 U10765 ( .A(n9568), .ZN(n9570) );
  AOI211_X1 U10766 ( .C1(n9572), .C2(n9571), .A(n9570), .B(n9569), .ZN(n9573)
         );
  AOI22_X1 U10767 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9573), .B1(n9603), .B2(
        P1_ADDR_REG_0__SCAN_IN), .ZN(n9576) );
  NAND3_X1 U10768 ( .A1(n9688), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9574), .ZN(
        n9575) );
  OAI211_X1 U10769 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n6563), .A(n9576), .B(
        n9575), .ZN(P1_U3241) );
  AOI22_X1 U10770 ( .A1(n9603), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(n9671), .B2(
        n9577), .ZN(n9589) );
  INV_X1 U10771 ( .A(n9578), .ZN(n9581) );
  INV_X1 U10772 ( .A(n9579), .ZN(n9580) );
  AOI211_X1 U10773 ( .C1(n9582), .C2(n9581), .A(n9580), .B(n9708), .ZN(n9587)
         );
  AOI211_X1 U10774 ( .C1(n9585), .C2(n9584), .A(n9583), .B(n9665), .ZN(n9586)
         );
  AOI211_X1 U10775 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(P1_U3084), .A(n9587), 
        .B(n9586), .ZN(n9588) );
  NAND2_X1 U10776 ( .A1(n9589), .A2(n9588), .ZN(P1_U3242) );
  AOI211_X1 U10777 ( .C1(n9592), .C2(n9591), .A(n9590), .B(n9708), .ZN(n9593)
         );
  AOI211_X1 U10778 ( .C1(P1_ADDR_REG_5__SCAN_IN), .C2(n9603), .A(n9594), .B(
        n9593), .ZN(n9601) );
  OAI21_X1 U10779 ( .B1(n9597), .B2(n9596), .A(n9595), .ZN(n9598) );
  AOI22_X1 U10780 ( .A1(n9671), .A2(n9599), .B1(n9698), .B2(n9598), .ZN(n9600)
         );
  NAND2_X1 U10781 ( .A1(n9601), .A2(n9600), .ZN(P1_U3246) );
  AOI22_X1 U10782 ( .A1(n9603), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n9671), .B2(
        n9602), .ZN(n9614) );
  OAI21_X1 U10783 ( .B1(n9606), .B2(n9605), .A(n9604), .ZN(n9612) );
  AOI211_X1 U10784 ( .C1(n9609), .C2(n9608), .A(n9607), .B(n9665), .ZN(n9610)
         );
  AOI211_X1 U10785 ( .C1(n9688), .C2(n9612), .A(n9611), .B(n9610), .ZN(n9613)
         );
  NAND2_X1 U10786 ( .A1(n9614), .A2(n9613), .ZN(P1_U3247) );
  OAI21_X1 U10787 ( .B1(n9617), .B2(n9616), .A(n9615), .ZN(n9622) );
  AOI211_X1 U10788 ( .C1(n9619), .C2(n9623), .A(n9618), .B(n9708), .ZN(n9620)
         );
  AOI211_X1 U10789 ( .C1(n9698), .C2(n9622), .A(n9621), .B(n9620), .ZN(n9627)
         );
  INV_X1 U10790 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9874) );
  NOR3_X1 U10791 ( .A1(n9708), .A2(n9874), .A3(n9623), .ZN(n9625) );
  OAI21_X1 U10792 ( .B1(n9671), .B2(n9625), .A(n9624), .ZN(n9626) );
  OAI211_X1 U10793 ( .C1(n9711), .C2(n9628), .A(n9627), .B(n9626), .ZN(
        P1_U3249) );
  AOI211_X1 U10794 ( .C1(n9631), .C2(n9630), .A(n9665), .B(n9629), .ZN(n9632)
         );
  AOI211_X1 U10795 ( .C1(n9671), .C2(n9634), .A(n9633), .B(n9632), .ZN(n9640)
         );
  AOI21_X1 U10796 ( .B1(n9637), .B2(n9636), .A(n9635), .ZN(n9638) );
  OR2_X1 U10797 ( .A1(n9638), .A2(n9708), .ZN(n9639) );
  OAI211_X1 U10798 ( .C1(n9711), .C2(n9641), .A(n9640), .B(n9639), .ZN(
        P1_U3254) );
  INV_X1 U10799 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9653) );
  AOI211_X1 U10800 ( .C1(n9643), .C2(n7214), .A(n9642), .B(n9665), .ZN(n9644)
         );
  AOI211_X1 U10801 ( .C1(n9671), .C2(n9646), .A(n9645), .B(n9644), .ZN(n9652)
         );
  AOI21_X1 U10802 ( .B1(n9649), .B2(n9648), .A(n9647), .ZN(n9650) );
  OR2_X1 U10803 ( .A1(n9650), .A2(n9708), .ZN(n9651) );
  OAI211_X1 U10804 ( .C1(n9653), .C2(n9711), .A(n9652), .B(n9651), .ZN(
        P1_U3255) );
  INV_X1 U10805 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9664) );
  AOI211_X1 U10806 ( .C1(n9656), .C2(n9655), .A(n9654), .B(n9665), .ZN(n9657)
         );
  AOI211_X1 U10807 ( .C1(n9659), .C2(n9671), .A(n9658), .B(n9657), .ZN(n9663)
         );
  OAI211_X1 U10808 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9661), .A(n9688), .B(
        n9660), .ZN(n9662) );
  OAI211_X1 U10809 ( .C1(n9664), .C2(n9711), .A(n9663), .B(n9662), .ZN(
        P1_U3256) );
  AOI211_X1 U10810 ( .C1(n9668), .C2(n9667), .A(n9666), .B(n9665), .ZN(n9669)
         );
  AOI211_X1 U10811 ( .C1(n9672), .C2(n9671), .A(n9670), .B(n9669), .ZN(n9677)
         );
  OAI211_X1 U10812 ( .C1(n9675), .C2(n9674), .A(n9688), .B(n9673), .ZN(n9676)
         );
  OAI211_X1 U10813 ( .C1(n9711), .C2(n9678), .A(n9677), .B(n9676), .ZN(
        P1_U3257) );
  INV_X1 U10814 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9693) );
  AOI21_X1 U10815 ( .B1(n9681), .B2(n9680), .A(n9679), .ZN(n9682) );
  NAND2_X1 U10816 ( .A1(n9698), .A2(n9682), .ZN(n9684) );
  OAI211_X1 U10817 ( .C1(n9702), .C2(n9685), .A(n9684), .B(n9683), .ZN(n9686)
         );
  INV_X1 U10818 ( .A(n9686), .ZN(n9692) );
  OAI211_X1 U10819 ( .C1(n9690), .C2(n9689), .A(n9688), .B(n9687), .ZN(n9691)
         );
  OAI211_X1 U10820 ( .C1(n9711), .C2(n9693), .A(n9692), .B(n9691), .ZN(
        P1_U3258) );
  INV_X1 U10821 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10063) );
  AOI21_X1 U10822 ( .B1(n9696), .B2(n9695), .A(n9694), .ZN(n9697) );
  NAND2_X1 U10823 ( .A1(n9698), .A2(n9697), .ZN(n9700) );
  OAI211_X1 U10824 ( .C1(n9702), .C2(n9701), .A(n9700), .B(n9699), .ZN(n9703)
         );
  INV_X1 U10825 ( .A(n9703), .ZN(n9710) );
  AOI21_X1 U10826 ( .B1(n9706), .B2(n9705), .A(n9704), .ZN(n9707) );
  OR2_X1 U10827 ( .A1(n9708), .A2(n9707), .ZN(n9709) );
  OAI211_X1 U10828 ( .C1(n10063), .C2(n9711), .A(n9710), .B(n9709), .ZN(
        P1_U3259) );
  NAND2_X1 U10829 ( .A1(n9713), .A2(n9714), .ZN(n9715) );
  NAND2_X1 U10830 ( .A1(n9712), .A2(n9715), .ZN(n9731) );
  INV_X1 U10831 ( .A(n9731), .ZN(n9846) );
  INV_X1 U10832 ( .A(n9716), .ZN(n9718) );
  OAI21_X1 U10833 ( .B1(n9718), .B2(n9842), .A(n9717), .ZN(n9843) );
  INV_X1 U10834 ( .A(n9843), .ZN(n9719) );
  AOI22_X1 U10835 ( .A1(n9846), .A2(n9764), .B1(n9720), .B2(n9719), .ZN(n9736)
         );
  OAI22_X1 U10836 ( .A1(n9722), .A2(n9774), .B1(n9721), .B2(n9772), .ZN(n9723)
         );
  INV_X1 U10837 ( .A(n9723), .ZN(n9729) );
  OAI21_X1 U10838 ( .B1(n9725), .B2(n9724), .A(n5064), .ZN(n9727) );
  NAND3_X1 U10839 ( .A1(n9727), .A2(n9770), .A3(n9726), .ZN(n9728) );
  OAI211_X1 U10840 ( .C1(n9731), .C2(n9730), .A(n9729), .B(n9728), .ZN(n9844)
         );
  AOI22_X1 U10841 ( .A1(n9755), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n9732), .B2(
        n9783), .ZN(n9733) );
  OAI21_X1 U10842 ( .B1(n9842), .B2(n9765), .A(n9733), .ZN(n9734) );
  AOI21_X1 U10843 ( .B1(n9844), .B2(n9779), .A(n9734), .ZN(n9735) );
  NAND2_X1 U10844 ( .A1(n9736), .A2(n9735), .ZN(P1_U3283) );
  INV_X1 U10845 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9754) );
  XOR2_X1 U10846 ( .A(n9737), .B(n9747), .Z(n9824) );
  XNOR2_X1 U10847 ( .A(n9761), .B(n9821), .ZN(n9738) );
  NAND2_X1 U10848 ( .A1(n9738), .A2(n9828), .ZN(n9820) );
  AOI22_X1 U10849 ( .A1(n9783), .A2(n9741), .B1(n9740), .B2(n9739), .ZN(n9744)
         );
  NAND2_X1 U10850 ( .A1(n9743), .A2(n9742), .ZN(n9819) );
  OAI211_X1 U10851 ( .C1(n9820), .C2(n9745), .A(n9744), .B(n9819), .ZN(n9751)
         );
  XOR2_X1 U10852 ( .A(n9747), .B(n9746), .Z(n9750) );
  OAI22_X1 U10853 ( .A1(n9750), .A2(n9749), .B1(n9748), .B2(n9774), .ZN(n9822)
         );
  AOI211_X1 U10854 ( .C1(n9752), .C2(n9824), .A(n9751), .B(n9822), .ZN(n9753)
         );
  AOI22_X1 U10855 ( .A1(n9755), .A2(n9754), .B1(n9753), .B2(n9779), .ZN(
        P1_U3286) );
  XNOR2_X1 U10856 ( .A(n9756), .B(n9757), .ZN(n9812) );
  NAND2_X1 U10857 ( .A1(n9759), .A2(n9758), .ZN(n9760) );
  NAND2_X1 U10858 ( .A1(n9761), .A2(n9760), .ZN(n9814) );
  NOR2_X1 U10859 ( .A1(n9814), .A2(n9762), .ZN(n9763) );
  AOI21_X1 U10860 ( .B1(n9812), .B2(n9764), .A(n9763), .ZN(n9785) );
  NOR2_X1 U10861 ( .A1(n9765), .A2(n9813), .ZN(n9781) );
  INV_X1 U10862 ( .A(n9766), .ZN(n9768) );
  INV_X1 U10863 ( .A(n9756), .ZN(n9767) );
  OAI22_X1 U10864 ( .A1(n9769), .A2(n9768), .B1(n9767), .B2(n7587), .ZN(n9771)
         );
  NAND2_X1 U10865 ( .A1(n9771), .A2(n9770), .ZN(n9778) );
  OAI22_X1 U10866 ( .A1(n4956), .A2(n9774), .B1(n9773), .B2(n9772), .ZN(n9775)
         );
  AOI21_X1 U10867 ( .B1(n9812), .B2(n9776), .A(n9775), .ZN(n9777) );
  NAND2_X1 U10868 ( .A1(n9778), .A2(n9777), .ZN(n9817) );
  MUX2_X1 U10869 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9817), .S(n9779), .Z(n9780)
         );
  AOI211_X1 U10870 ( .C1(n9783), .C2(n9782), .A(n9781), .B(n9780), .ZN(n9784)
         );
  NAND2_X1 U10871 ( .A1(n9785), .A2(n9784), .ZN(P1_U3287) );
  AND2_X1 U10872 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9789), .ZN(P1_U3292) );
  AND2_X1 U10873 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9789), .ZN(P1_U3293) );
  AND2_X1 U10874 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9789), .ZN(P1_U3294) );
  AND2_X1 U10875 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9789), .ZN(P1_U3295) );
  INV_X1 U10876 ( .A(n9789), .ZN(n9788) );
  NOR2_X1 U10877 ( .A1(n9788), .A2(n9786), .ZN(P1_U3296) );
  AND2_X1 U10878 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9789), .ZN(P1_U3297) );
  AND2_X1 U10879 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9789), .ZN(P1_U3298) );
  AND2_X1 U10880 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9789), .ZN(P1_U3299) );
  AND2_X1 U10881 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9789), .ZN(P1_U3300) );
  AND2_X1 U10882 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9789), .ZN(P1_U3301) );
  AND2_X1 U10883 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9789), .ZN(P1_U3302) );
  AND2_X1 U10884 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9789), .ZN(P1_U3303) );
  AND2_X1 U10885 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9789), .ZN(P1_U3304) );
  AND2_X1 U10886 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9789), .ZN(P1_U3305) );
  AND2_X1 U10887 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9789), .ZN(P1_U3306) );
  AND2_X1 U10888 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9789), .ZN(P1_U3307) );
  AND2_X1 U10889 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9789), .ZN(P1_U3308) );
  AND2_X1 U10890 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9789), .ZN(P1_U3309) );
  AND2_X1 U10891 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9789), .ZN(P1_U3310) );
  AND2_X1 U10892 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9789), .ZN(P1_U3311) );
  AND2_X1 U10893 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9789), .ZN(P1_U3312) );
  NOR2_X1 U10894 ( .A1(n9788), .A2(n9787), .ZN(P1_U3313) );
  AND2_X1 U10895 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9789), .ZN(P1_U3314) );
  AND2_X1 U10896 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9789), .ZN(P1_U3315) );
  AND2_X1 U10897 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9789), .ZN(P1_U3316) );
  AND2_X1 U10898 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9789), .ZN(P1_U3317) );
  AND2_X1 U10899 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9789), .ZN(P1_U3318) );
  AND2_X1 U10900 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9789), .ZN(P1_U3319) );
  AND2_X1 U10901 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9789), .ZN(P1_U3320) );
  AND2_X1 U10902 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9789), .ZN(P1_U3321) );
  AOI21_X1 U10903 ( .B1(P1_D_REG_1__SCAN_IN), .B2(n9791), .A(n9790), .ZN(n9792) );
  INV_X1 U10904 ( .A(n9792), .ZN(P1_U3441) );
  INV_X1 U10905 ( .A(n9793), .ZN(n9798) );
  OAI21_X1 U10906 ( .B1(n9795), .B2(n9849), .A(n9794), .ZN(n9797) );
  AOI211_X1 U10907 ( .C1(n9847), .C2(n9798), .A(n9797), .B(n9796), .ZN(n9861)
         );
  INV_X1 U10908 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9799) );
  AOI22_X1 U10909 ( .A1(n9859), .A2(n9861), .B1(n9799), .B2(n9857), .ZN(
        P1_U3457) );
  OAI22_X1 U10910 ( .A1(n9800), .A2(n9851), .B1(n4931), .B2(n9849), .ZN(n9802)
         );
  AOI211_X1 U10911 ( .C1(n9847), .C2(n9803), .A(n9802), .B(n9801), .ZN(n9863)
         );
  INV_X1 U10912 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9804) );
  AOI22_X1 U10913 ( .A1(n9859), .A2(n9863), .B1(n9804), .B2(n9857), .ZN(
        P1_U3460) );
  OAI22_X1 U10914 ( .A1(n9806), .A2(n9851), .B1(n9805), .B2(n9849), .ZN(n9807)
         );
  AOI21_X1 U10915 ( .B1(n9808), .B2(n9847), .A(n9807), .ZN(n9809) );
  AND2_X1 U10916 ( .A1(n9810), .A2(n9809), .ZN(n9865) );
  INV_X1 U10917 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9811) );
  AOI22_X1 U10918 ( .A1(n9859), .A2(n9865), .B1(n9811), .B2(n9857), .ZN(
        P1_U3463) );
  AND2_X1 U10919 ( .A1(n9812), .A2(n9847), .ZN(n9816) );
  OAI22_X1 U10920 ( .A1(n9814), .A2(n9851), .B1(n9813), .B2(n9849), .ZN(n9815)
         );
  NOR3_X1 U10921 ( .A1(n9817), .A2(n9816), .A3(n9815), .ZN(n9867) );
  INV_X1 U10922 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9818) );
  AOI22_X1 U10923 ( .A1(n9859), .A2(n9867), .B1(n9818), .B2(n9857), .ZN(
        P1_U3466) );
  OAI211_X1 U10924 ( .C1(n9821), .C2(n9849), .A(n9820), .B(n9819), .ZN(n9823)
         );
  AOI211_X1 U10925 ( .C1(n9855), .C2(n9824), .A(n9823), .B(n9822), .ZN(n9869)
         );
  INV_X1 U10926 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9825) );
  AOI22_X1 U10927 ( .A1(n9859), .A2(n9869), .B1(n9825), .B2(n9857), .ZN(
        P1_U3469) );
  AOI22_X1 U10928 ( .A1(n9829), .A2(n9828), .B1(n9827), .B2(n9826), .ZN(n9830)
         );
  OAI211_X1 U10929 ( .C1(n9833), .C2(n9832), .A(n9831), .B(n9830), .ZN(n9834)
         );
  INV_X1 U10930 ( .A(n9834), .ZN(n9871) );
  AOI22_X1 U10931 ( .A1(n9859), .A2(n9871), .B1(n9835), .B2(n9857), .ZN(
        P1_U3472) );
  OAI21_X1 U10932 ( .B1(n9837), .B2(n9849), .A(n9836), .ZN(n9839) );
  AOI211_X1 U10933 ( .C1(n9855), .C2(n9840), .A(n9839), .B(n9838), .ZN(n9873)
         );
  INV_X1 U10934 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9841) );
  AOI22_X1 U10935 ( .A1(n9859), .A2(n9873), .B1(n9841), .B2(n9857), .ZN(
        P1_U3475) );
  OAI22_X1 U10936 ( .A1(n9843), .A2(n9851), .B1(n9842), .B2(n9849), .ZN(n9845)
         );
  AOI211_X1 U10937 ( .C1(n9847), .C2(n9846), .A(n9845), .B(n9844), .ZN(n9875)
         );
  INV_X1 U10938 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9848) );
  AOI22_X1 U10939 ( .A1(n9859), .A2(n9875), .B1(n9848), .B2(n9857), .ZN(
        P1_U3478) );
  OAI22_X1 U10940 ( .A1(n9852), .A2(n9851), .B1(n9850), .B2(n9849), .ZN(n9854)
         );
  AOI211_X1 U10941 ( .C1(n9856), .C2(n9855), .A(n9854), .B(n9853), .ZN(n9878)
         );
  INV_X1 U10942 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9858) );
  AOI22_X1 U10943 ( .A1(n9859), .A2(n9878), .B1(n9858), .B2(n9857), .ZN(
        P1_U3481) );
  AOI22_X1 U10944 ( .A1(n9879), .A2(n9861), .B1(n9860), .B2(n9876), .ZN(
        P1_U3524) );
  AOI22_X1 U10945 ( .A1(n9879), .A2(n9863), .B1(n9862), .B2(n9876), .ZN(
        P1_U3525) );
  AOI22_X1 U10946 ( .A1(n9879), .A2(n9865), .B1(n9864), .B2(n9876), .ZN(
        P1_U3526) );
  AOI22_X1 U10947 ( .A1(n9879), .A2(n9867), .B1(n9866), .B2(n9876), .ZN(
        P1_U3527) );
  INV_X1 U10948 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9868) );
  AOI22_X1 U10949 ( .A1(n9879), .A2(n9869), .B1(n9868), .B2(n9876), .ZN(
        P1_U3528) );
  INV_X1 U10950 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9870) );
  AOI22_X1 U10951 ( .A1(n9879), .A2(n9871), .B1(n9870), .B2(n9876), .ZN(
        P1_U3529) );
  INV_X1 U10952 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9872) );
  AOI22_X1 U10953 ( .A1(n9879), .A2(n9873), .B1(n9872), .B2(n9876), .ZN(
        P1_U3530) );
  AOI22_X1 U10954 ( .A1(n9879), .A2(n9875), .B1(n9874), .B2(n9876), .ZN(
        P1_U3531) );
  AOI22_X1 U10955 ( .A1(n9879), .A2(n9878), .B1(n9877), .B2(n9876), .ZN(
        P1_U3532) );
  AOI22_X1 U10956 ( .A1(n9881), .A2(n9880), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3152), .ZN(n9890) );
  AOI21_X1 U10957 ( .B1(n9884), .B2(n9883), .A(n9882), .ZN(n9888) );
  AOI22_X1 U10958 ( .A1(n9888), .A2(n9887), .B1(n9886), .B2(n9885), .ZN(n9889)
         );
  OAI211_X1 U10959 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n9891), .A(n9890), .B(
        n9889), .ZN(P2_U3220) );
  AOI22_X1 U10960 ( .A1(n9897), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9892), .ZN(n9902) );
  NOR2_X1 U10961 ( .A1(n9893), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9894) );
  AOI211_X1 U10962 ( .C1(n9897), .C2(n9896), .A(n9895), .B(n9894), .ZN(n9900)
         );
  AOI22_X1 U10963 ( .A1(n9898), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9899) );
  OAI221_X1 U10964 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9902), .C1(n9901), .C2(
        n9900), .A(n9899), .ZN(P2_U3245) );
  AND2_X1 U10965 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9909), .ZN(P2_U3297) );
  AND2_X1 U10966 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9909), .ZN(P2_U3298) );
  AND2_X1 U10967 ( .A1(n9909), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3299) );
  AND2_X1 U10968 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9909), .ZN(P2_U3300) );
  AND2_X1 U10969 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9909), .ZN(P2_U3301) );
  AND2_X1 U10970 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9909), .ZN(P2_U3302) );
  AND2_X1 U10971 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9909), .ZN(P2_U3303) );
  AND2_X1 U10972 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9909), .ZN(P2_U3304) );
  AND2_X1 U10973 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9909), .ZN(P2_U3305) );
  AND2_X1 U10974 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9909), .ZN(P2_U3306) );
  AND2_X1 U10975 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9909), .ZN(P2_U3307) );
  AND2_X1 U10976 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9909), .ZN(P2_U3308) );
  AND2_X1 U10977 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9909), .ZN(P2_U3309) );
  AND2_X1 U10978 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9909), .ZN(P2_U3310) );
  AND2_X1 U10979 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9909), .ZN(P2_U3311) );
  AND2_X1 U10980 ( .A1(n9909), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3312) );
  AND2_X1 U10981 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9909), .ZN(P2_U3313) );
  AND2_X1 U10982 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9909), .ZN(P2_U3314) );
  AND2_X1 U10983 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9909), .ZN(P2_U3315) );
  AND2_X1 U10984 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9909), .ZN(P2_U3316) );
  AND2_X1 U10985 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9909), .ZN(P2_U3317) );
  AND2_X1 U10986 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9909), .ZN(P2_U3318) );
  AND2_X1 U10987 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9909), .ZN(P2_U3319) );
  AND2_X1 U10988 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9909), .ZN(P2_U3320) );
  NOR2_X1 U10989 ( .A1(n9906), .A2(n9905), .ZN(P2_U3321) );
  AND2_X1 U10990 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9909), .ZN(P2_U3322) );
  AND2_X1 U10991 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9909), .ZN(P2_U3323) );
  AND2_X1 U10992 ( .A1(n9909), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3324) );
  AND2_X1 U10993 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9909), .ZN(P2_U3325) );
  AND2_X1 U10994 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9909), .ZN(P2_U3326) );
  AOI22_X1 U10995 ( .A1(n9912), .A2(n9908), .B1(n9907), .B2(n9909), .ZN(
        P2_U3437) );
  AOI22_X1 U10996 ( .A1(n9912), .A2(n9911), .B1(n9910), .B2(n9909), .ZN(
        P2_U3438) );
  AOI22_X1 U10997 ( .A1(n9915), .A2(n10001), .B1(n9914), .B2(n9913), .ZN(n9916) );
  AND2_X1 U10998 ( .A1(n9917), .A2(n9916), .ZN(n10006) );
  AOI22_X1 U10999 ( .A1(n10004), .A2(n10006), .B1(n9918), .B2(n10002), .ZN(
        P2_U3451) );
  AOI21_X1 U11000 ( .B1(n9930), .B2(n9920), .A(n9919), .ZN(n9921) );
  OAI211_X1 U11001 ( .C1(n9924), .C2(n9923), .A(n9922), .B(n9921), .ZN(n9925)
         );
  INV_X1 U11002 ( .A(n9925), .ZN(n10008) );
  INV_X1 U11003 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9926) );
  AOI22_X1 U11004 ( .A1(n10004), .A2(n10008), .B1(n9926), .B2(n10002), .ZN(
        P2_U3454) );
  AOI211_X1 U11005 ( .C1(n9930), .C2(n9929), .A(n9928), .B(n9927), .ZN(n9931)
         );
  INV_X1 U11006 ( .A(n9931), .ZN(n9932) );
  AOI21_X1 U11007 ( .B1(n10001), .B2(n9933), .A(n9932), .ZN(n10009) );
  INV_X1 U11008 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9934) );
  AOI22_X1 U11009 ( .A1(n10004), .A2(n10009), .B1(n9934), .B2(n10002), .ZN(
        P2_U3457) );
  OAI21_X1 U11010 ( .B1(n9936), .B2(n9994), .A(n9935), .ZN(n9937) );
  AOI21_X1 U11011 ( .B1(n9938), .B2(n9985), .A(n9937), .ZN(n9939) );
  AND2_X1 U11012 ( .A1(n9940), .A2(n9939), .ZN(n10011) );
  INV_X1 U11013 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9941) );
  AOI22_X1 U11014 ( .A1(n10004), .A2(n10011), .B1(n9941), .B2(n10002), .ZN(
        P2_U3460) );
  OAI22_X1 U11015 ( .A1(n9943), .A2(n9996), .B1(n9942), .B2(n9994), .ZN(n9945)
         );
  AOI211_X1 U11016 ( .C1(n10001), .C2(n9946), .A(n9945), .B(n9944), .ZN(n10012) );
  INV_X1 U11017 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9947) );
  AOI22_X1 U11018 ( .A1(n10004), .A2(n10012), .B1(n9947), .B2(n10002), .ZN(
        P2_U3463) );
  OAI211_X1 U11019 ( .C1(n9950), .C2(n9994), .A(n9949), .B(n9948), .ZN(n9951)
         );
  AOI21_X1 U11020 ( .B1(n10001), .B2(n9952), .A(n9951), .ZN(n10013) );
  INV_X1 U11021 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9953) );
  AOI22_X1 U11022 ( .A1(n10004), .A2(n10013), .B1(n9953), .B2(n10002), .ZN(
        P2_U3466) );
  OAI211_X1 U11023 ( .C1(n9956), .C2(n9994), .A(n9955), .B(n9954), .ZN(n9957)
         );
  AOI21_X1 U11024 ( .B1(n10001), .B2(n9958), .A(n9957), .ZN(n10014) );
  INV_X1 U11025 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9959) );
  AOI22_X1 U11026 ( .A1(n10004), .A2(n10014), .B1(n9959), .B2(n10002), .ZN(
        P2_U3469) );
  OAI22_X1 U11027 ( .A1(n9961), .A2(n9996), .B1(n9960), .B2(n9994), .ZN(n9963)
         );
  AOI211_X1 U11028 ( .C1(n10001), .C2(n9964), .A(n9963), .B(n9962), .ZN(n10015) );
  INV_X1 U11029 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9965) );
  AOI22_X1 U11030 ( .A1(n10004), .A2(n10015), .B1(n9965), .B2(n10002), .ZN(
        P2_U3472) );
  OAI22_X1 U11031 ( .A1(n9967), .A2(n9996), .B1(n9966), .B2(n9994), .ZN(n9969)
         );
  AOI211_X1 U11032 ( .C1(n9985), .C2(n9970), .A(n9969), .B(n9968), .ZN(n10017)
         );
  INV_X1 U11033 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9971) );
  AOI22_X1 U11034 ( .A1(n10004), .A2(n10017), .B1(n9971), .B2(n10002), .ZN(
        P2_U3475) );
  INV_X1 U11035 ( .A(n9972), .ZN(n9977) );
  OAI22_X1 U11036 ( .A1(n9974), .A2(n9996), .B1(n9973), .B2(n9994), .ZN(n9976)
         );
  AOI211_X1 U11037 ( .C1(n9985), .C2(n9977), .A(n9976), .B(n9975), .ZN(n10018)
         );
  AOI22_X1 U11038 ( .A1(n10004), .A2(n10018), .B1(n9978), .B2(n10002), .ZN(
        P2_U3478) );
  INV_X1 U11039 ( .A(n9979), .ZN(n9984) );
  OAI22_X1 U11040 ( .A1(n9981), .A2(n9996), .B1(n9980), .B2(n9994), .ZN(n9983)
         );
  AOI211_X1 U11041 ( .C1(n9985), .C2(n9984), .A(n9983), .B(n9982), .ZN(n10019)
         );
  INV_X1 U11042 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9986) );
  AOI22_X1 U11043 ( .A1(n10004), .A2(n10019), .B1(n9986), .B2(n10002), .ZN(
        P2_U3481) );
  INV_X1 U11044 ( .A(n9987), .ZN(n9992) );
  OAI22_X1 U11045 ( .A1(n9989), .A2(n9996), .B1(n9988), .B2(n9994), .ZN(n9991)
         );
  AOI211_X1 U11046 ( .C1(n9992), .C2(n10001), .A(n9991), .B(n9990), .ZN(n10020) );
  INV_X1 U11047 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9993) );
  AOI22_X1 U11048 ( .A1(n10004), .A2(n10020), .B1(n9993), .B2(n10002), .ZN(
        P2_U3484) );
  OAI22_X1 U11049 ( .A1(n9997), .A2(n9996), .B1(n9995), .B2(n9994), .ZN(n9999)
         );
  AOI211_X1 U11050 ( .C1(n10001), .C2(n10000), .A(n9999), .B(n9998), .ZN(
        n10022) );
  INV_X1 U11051 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10003) );
  AOI22_X1 U11052 ( .A1(n10004), .A2(n10022), .B1(n10003), .B2(n10002), .ZN(
        P2_U3487) );
  AOI22_X1 U11053 ( .A1(n10023), .A2(n10006), .B1(n10005), .B2(n10021), .ZN(
        P2_U3520) );
  AOI22_X1 U11054 ( .A1(n10023), .A2(n10008), .B1(n10007), .B2(n10021), .ZN(
        P2_U3521) );
  AOI22_X1 U11055 ( .A1(n10023), .A2(n10009), .B1(n6270), .B2(n10021), .ZN(
        P2_U3522) );
  AOI22_X1 U11056 ( .A1(n10023), .A2(n10011), .B1(n10010), .B2(n10021), .ZN(
        P2_U3523) );
  AOI22_X1 U11057 ( .A1(n10023), .A2(n10012), .B1(n6273), .B2(n10021), .ZN(
        P2_U3524) );
  AOI22_X1 U11058 ( .A1(n10023), .A2(n10013), .B1(n6288), .B2(n10021), .ZN(
        P2_U3525) );
  AOI22_X1 U11059 ( .A1(n10023), .A2(n10014), .B1(n6307), .B2(n10021), .ZN(
        P2_U3526) );
  AOI22_X1 U11060 ( .A1(n10023), .A2(n10015), .B1(n6319), .B2(n10021), .ZN(
        P2_U3527) );
  AOI22_X1 U11061 ( .A1(n10023), .A2(n10017), .B1(n10016), .B2(n10021), .ZN(
        P2_U3528) );
  AOI22_X1 U11062 ( .A1(n10023), .A2(n10018), .B1(n6348), .B2(n10021), .ZN(
        P2_U3529) );
  AOI22_X1 U11063 ( .A1(n10023), .A2(n10019), .B1(n6362), .B2(n10021), .ZN(
        P2_U3530) );
  AOI22_X1 U11064 ( .A1(n10023), .A2(n10020), .B1(n6734), .B2(n10021), .ZN(
        P2_U3531) );
  AOI22_X1 U11065 ( .A1(n10023), .A2(n10022), .B1(n6733), .B2(n10021), .ZN(
        P2_U3532) );
  INV_X1 U11066 ( .A(n10024), .ZN(n10025) );
  NAND2_X1 U11067 ( .A1(n10026), .A2(n10025), .ZN(n10027) );
  XOR2_X1 U11068 ( .A(n10028), .B(n10027), .Z(ADD_1071_U5) );
  XOR2_X1 U11069 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11070 ( .B1(n10031), .B2(n10030), .A(n10029), .ZN(ADD_1071_U56) );
  OAI21_X1 U11071 ( .B1(n10034), .B2(n10033), .A(n10032), .ZN(ADD_1071_U57) );
  OAI21_X1 U11072 ( .B1(n10037), .B2(n10036), .A(n10035), .ZN(ADD_1071_U58) );
  OAI21_X1 U11073 ( .B1(n10040), .B2(n10039), .A(n10038), .ZN(ADD_1071_U59) );
  OAI21_X1 U11074 ( .B1(n10043), .B2(n10042), .A(n10041), .ZN(ADD_1071_U60) );
  OAI21_X1 U11075 ( .B1(n10046), .B2(n10045), .A(n10044), .ZN(ADD_1071_U61) );
  AOI21_X1 U11076 ( .B1(n10049), .B2(n10048), .A(n10047), .ZN(ADD_1071_U62) );
  AOI21_X1 U11077 ( .B1(n10052), .B2(n10051), .A(n10050), .ZN(ADD_1071_U63) );
  XOR2_X1 U11078 ( .A(n10053), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11079 ( .A1(n10055), .A2(n10054), .ZN(n10056) );
  XOR2_X1 U11080 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10056), .Z(ADD_1071_U51) );
  AOI21_X1 U11081 ( .B1(n10059), .B2(n10058), .A(n10057), .ZN(ADD_1071_U47) );
  OAI21_X1 U11082 ( .B1(n10062), .B2(n10061), .A(n10060), .ZN(n10064) );
  XOR2_X1 U11083 ( .A(n10064), .B(n10063), .Z(ADD_1071_U55) );
  XOR2_X1 U11084 ( .A(n10066), .B(n10065), .Z(ADD_1071_U54) );
  XOR2_X1 U11085 ( .A(n10067), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11086 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10068), .Z(ADD_1071_U48) );
  XOR2_X1 U11087 ( .A(n10070), .B(n10069), .Z(ADD_1071_U53) );
  XNOR2_X1 U11088 ( .A(n10072), .B(n10071), .ZN(ADD_1071_U52) );
  AND2_X1 U4911 ( .A1(n8531), .A2(n7836), .ZN(n9913) );
  AND2_X1 U4826 ( .A1(n6110), .A2(n7845), .ZN(n7390) );
  CLKBUF_X1 U4836 ( .A(n5625), .Z(n4308) );
  NAND2_X1 U4905 ( .A1(n6697), .A2(n6696), .ZN(n6702) );
  CLKBUF_X1 U6000 ( .A(n4960), .Z(n5535) );
endmodule

