

module b22_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n7448, n7449, n7451, n7452, n7454, n7455, n7456, n7457, n7458, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587;

  INV_X4 U7549 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7550 ( .A(n12707), .ZN(n15371) );
  NAND2_X1 U7551 ( .A1(n9766), .A2(n9765), .ZN(n15382) );
  INV_X4 U7553 ( .A(n14594), .ZN(n7458) );
  INV_X1 U7555 ( .A(n8592), .ZN(n16402) );
  INV_X2 U7556 ( .A(n9027), .ZN(n12997) );
  OAI211_X1 U7557 ( .C1(n8616), .C2(SI_2_), .A(n8557), .B(n8556), .ZN(n8592)
         );
  NAND2_X2 U7558 ( .A1(n10725), .A2(n10724), .ZN(n14044) );
  AND2_X1 U7559 ( .A1(n13071), .A2(n8540), .ZN(n8950) );
  CLKBUF_X2 U7560 ( .A(n9338), .Z(n9857) );
  INV_X1 U7561 ( .A(n10053), .ZN(n10051) );
  NAND2_X1 U7562 ( .A1(n10042), .A2(n10171), .ZN(n14185) );
  CLKBUF_X2 U7563 ( .A(n9283), .Z(n7719) );
  CLKBUF_X1 U7564 ( .A(n9303), .Z(n9758) );
  NAND2_X2 U7565 ( .A1(n9165), .A2(n9164), .ZN(n9724) );
  NAND2_X1 U7566 ( .A1(n9265), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9264) );
  NAND2_X1 U7567 ( .A1(n7891), .A2(n7892), .ZN(n9265) );
  INV_X1 U7568 ( .A(n14634), .ZN(n7448) );
  INV_X1 U7569 ( .A(n7448), .ZN(n7449) );
  OAI21_X1 U7570 ( .B1(n14282), .B2(n14287), .A(n10090), .ZN(n14634) );
  XNOR2_X1 U7571 ( .A(n13291), .B(n13292), .ZN(n13270) );
  NAND2_X1 U7572 ( .A1(n9253), .A2(n9730), .ZN(n9256) );
  NAND2_X1 U7573 ( .A1(n9247), .A2(n9246), .ZN(n9249) );
  NAND2_X1 U7576 ( .A1(n11422), .A2(n11839), .ZN(n11421) );
  INV_X1 U7577 ( .A(n10986), .ZN(n14181) );
  XNOR2_X1 U7578 ( .A(n9889), .B(n14939), .ZN(n15110) );
  INV_X1 U7579 ( .A(n10927), .ZN(n7613) );
  NAND2_X1 U7580 ( .A1(n9008), .A2(n9007), .ZN(n13412) );
  BUF_X1 U7581 ( .A(n13992), .Z(n11656) );
  NAND2_X1 U7582 ( .A1(n7856), .A2(n13826), .ZN(n14760) );
  NOR2_X1 U7583 ( .A1(n8164), .A2(n8163), .ZN(n8162) );
  INV_X1 U7584 ( .A(n9842), .ZN(n9808) );
  NAND2_X1 U7585 ( .A1(n15902), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9160) );
  NAND2_X1 U7586 ( .A1(n8162), .A2(n8165), .ZN(n14807) );
  NAND4_X2 U7587 ( .A1(n9308), .A2(n9307), .A3(n9306), .A4(n9305), .ZN(n9332)
         );
  NOR2_X4 U7589 ( .A1(n14578), .A2(n14564), .ZN(n7996) );
  NOR2_X2 U7590 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n7896) );
  INV_X1 U7591 ( .A(n10838), .ZN(n7692) );
  AND3_X1 U7592 ( .A1(n9330), .A2(n9328), .A3(n9329), .ZN(n7506) );
  OR2_X2 U7593 ( .A1(n12282), .A2(n8248), .ZN(n8247) );
  OAI21_X2 U7594 ( .B1(n9658), .B2(n9243), .A(n9242), .ZN(n9678) );
  AND3_X2 U7597 ( .A1(n9295), .A2(n9296), .A3(n9294), .ZN(n10439) );
  OR2_X2 U7598 ( .A1(n14041), .A2(n14040), .ZN(n7539) );
  NOR2_X2 U7599 ( .A1(n15171), .A2(n15395), .ZN(n8012) );
  XNOR2_X2 U7602 ( .A(n9254), .B(n15705), .ZN(n9253) );
  NAND2_X1 U7603 ( .A1(n9283), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9287) );
  XNOR2_X2 U7604 ( .A(n15928), .B(n7981), .ZN(n15991) );
  NAND2_X2 U7605 ( .A1(n15926), .A2(n15927), .ZN(n15928) );
  INV_X1 U7606 ( .A(n15342), .ZN(n10642) );
  CLKBUF_X1 U7607 ( .A(n7457), .Z(n7451) );
  CLKBUF_X3 U7608 ( .A(n7457), .Z(n7452) );
  AND2_X4 U7609 ( .A1(n8541), .A2(n8540), .ZN(n8718) );
  INV_X1 U7610 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7454) );
  XNOR2_X2 U7611 ( .A(n13798), .B(n13796), .ZN(n13959) );
  INV_X2 U7612 ( .A(n9165), .ZN(n15909) );
  XNOR2_X2 U7613 ( .A(n9162), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9165) );
  OAI211_X2 U7614 ( .C1(n9256), .C2(n8232), .A(n9262), .B(n8231), .ZN(n9782)
         );
  OAI21_X2 U7615 ( .B1(n8673), .B2(n8672), .A(n8674), .ZN(n8677) );
  NAND2_X2 U7616 ( .A1(n8038), .A2(n8037), .ZN(n8673) );
  OAI22_X2 U7617 ( .A1(n15935), .A2(n16000), .B1(n15936), .B2(
        P3_ADDR_REG_6__SCAN_IN), .ZN(n15937) );
  AOI21_X2 U7618 ( .B1(n14418), .B2(n7449), .A(n14417), .ZN(n14666) );
  NAND2_X4 U7619 ( .A1(n10020), .A2(n10019), .ZN(n10059) );
  AND2_X2 U7620 ( .A1(n7652), .A2(n7655), .ZN(n10019) );
  NAND4_X4 U7621 ( .A1(n10075), .A2(n10074), .A3(n10073), .A4(n10072), .ZN(
        n14318) );
  AOI21_X2 U7622 ( .B1(n16184), .B2(n16013), .A(n16297), .ZN(n16016) );
  NOR2_X2 U7623 ( .A1(n16298), .A2(n16299), .ZN(n16297) );
  AND2_X1 U7624 ( .A1(n10491), .A2(n11549), .ZN(n7455) );
  AND2_X1 U7625 ( .A1(n10491), .A2(n11549), .ZN(n15471) );
  XNOR2_X2 U7626 ( .A(n7775), .B(n7774), .ZN(n13303) );
  AOI21_X2 U7627 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n12006), .A(n12005), .ZN(
        n12195) );
  XNOR2_X2 U7628 ( .A(n9249), .B(SI_22_), .ZN(n11957) );
  XNOR2_X2 U7629 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n15982) );
  NAND2_X2 U7630 ( .A1(n11777), .A2(n11776), .ZN(n14084) );
  XNOR2_X2 U7631 ( .A(n10085), .B(P2_IR_REG_21__SCAN_IN), .ZN(n10125) );
  AOI22_X1 U7632 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n7464), .B1(n10048), .B2(
        n16107), .ZN(n8292) );
  AOI21_X2 U7633 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n16107), .A(n16102), .ZN(
        n16112) );
  NOR2_X2 U7634 ( .A1(n16009), .A2(n16010), .ZN(n16290) );
  NOR2_X2 U7635 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n16286), .ZN(n16009) );
  AOI21_X2 U7636 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n13268), .A(n13267), .ZN(
        n13291) );
  OAI21_X1 U7637 ( .B1(n14154), .B2(n7963), .A(n7960), .ZN(n14160) );
  OR2_X1 U7638 ( .A1(n14149), .A2(n14148), .ZN(n14154) );
  NAND2_X2 U7639 ( .A1(n12844), .A2(n12848), .ZN(n13413) );
  NAND2_X1 U7640 ( .A1(n13871), .A2(n7596), .ZN(n13872) );
  XNOR2_X1 U7641 ( .A(n13800), .B(n7920), .ZN(n13871) );
  NAND2_X1 U7643 ( .A1(n7909), .A2(n7910), .ZN(n12739) );
  AND2_X1 U7644 ( .A1(n7977), .A2(n7976), .ZN(n16293) );
  OAI22_X1 U7645 ( .A1(n14035), .A2(n7972), .B1(n14033), .B2(n14034), .ZN(
        n14041) );
  NOR2_X1 U7646 ( .A1(n11080), .A2(n7531), .ZN(n11083) );
  INV_X4 U7647 ( .A(n9857), .ZN(n9837) );
  AND2_X2 U7648 ( .A1(n8290), .A2(n8289), .ZN(n9338) );
  INV_X1 U7649 ( .A(n8573), .ZN(n13227) );
  CLKBUF_X2 U7650 ( .A(n14964), .Z(P1_U4016) );
  INV_X4 U7651 ( .A(n7468), .ZN(n7456) );
  NAND2_X1 U7652 ( .A1(n10441), .A2(n10437), .ZN(n10644) );
  CLKBUF_X2 U7653 ( .A(P3_U3897), .Z(n16079) );
  INV_X2 U7654 ( .A(n14206), .ZN(n14176) );
  CLKBUF_X3 U7655 ( .A(n13771), .Z(n7463) );
  BUF_X2 U7656 ( .A(n11900), .Z(n14201) );
  INV_X1 U7657 ( .A(n14206), .ZN(n7457) );
  NAND2_X2 U7660 ( .A1(n12592), .A2(n9838), .ZN(n9976) );
  INV_X2 U7661 ( .A(n12285), .ZN(n13357) );
  BUF_X2 U7662 ( .A(n10057), .Z(n10986) );
  NAND3_X1 U7663 ( .A1(n8138), .A2(n13986), .A3(n8137), .ZN(n13771) );
  INV_X4 U7664 ( .A(n14191), .ZN(n13902) );
  NAND2_X2 U7665 ( .A1(n10927), .A2(n10171), .ZN(n8616) );
  CLKBUF_X2 U7666 ( .A(n9724), .Z(n9847) );
  BUF_X2 U7667 ( .A(n8950), .Z(n9009) );
  INV_X2 U7668 ( .A(n15185), .ZN(n12592) );
  AND2_X1 U7669 ( .A1(n10008), .A2(n10009), .ZN(n7670) );
  INV_X1 U7670 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n10087) );
  NOR2_X1 U7671 ( .A1(n9049), .A2(n9048), .ZN(n13040) );
  AND2_X1 U7672 ( .A1(n8155), .A2(n8154), .ZN(n13978) );
  AOI21_X1 U7673 ( .B1(n13451), .B2(n7504), .A(n8082), .ZN(n13401) );
  NAND2_X1 U7674 ( .A1(n13811), .A2(n13801), .ZN(n7919) );
  NAND2_X1 U7675 ( .A1(n12843), .A2(n12847), .ZN(n13425) );
  NAND2_X1 U7676 ( .A1(n7991), .A2(n7990), .ZN(n14460) );
  NAND2_X1 U7677 ( .A1(n7675), .A2(n9831), .ZN(n14186) );
  NAND2_X1 U7678 ( .A1(n8999), .A2(n8998), .ZN(n9005) );
  OR2_X1 U7679 ( .A1(n11990), .A2(n7613), .ZN(n13687) );
  NAND2_X1 U7680 ( .A1(n8979), .A2(n8978), .ZN(n8996) );
  OAI21_X1 U7681 ( .B1(n9854), .B2(n9853), .A(n9789), .ZN(n9824) );
  NAND2_X1 U7682 ( .A1(n9752), .A2(n9751), .ZN(n15388) );
  NAND2_X1 U7683 ( .A1(n9785), .A2(n9784), .ZN(n9854) );
  CLKBUF_X1 U7684 ( .A(n12220), .Z(n7723) );
  NAND2_X1 U7685 ( .A1(n9733), .A2(n9732), .ZN(n15395) );
  NOR2_X1 U7686 ( .A1(n13257), .A2(n8028), .ZN(n13276) );
  NAND2_X1 U7687 ( .A1(n8975), .A2(n8963), .ZN(n8964) );
  NAND2_X1 U7688 ( .A1(n9715), .A2(n9714), .ZN(n15183) );
  OR2_X1 U7689 ( .A1(n8962), .A2(n13813), .ZN(n8975) );
  OAI21_X1 U7690 ( .B1(n8960), .B2(n8959), .A(n8961), .ZN(n8962) );
  NAND2_X1 U7691 ( .A1(n12335), .A2(n12334), .ZN(n12553) );
  NAND2_X1 U7692 ( .A1(n8947), .A2(n8946), .ZN(n8960) );
  AOI21_X1 U7693 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n12276), .A(n16190), .ZN(
        n14346) );
  OR2_X1 U7694 ( .A1(n8899), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8900) );
  NAND2_X1 U7695 ( .A1(n8899), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8913) );
  XNOR2_X1 U7696 ( .A(n9240), .B(n10656), .ZN(n9658) );
  NAND2_X2 U7697 ( .A1(n11903), .A2(n11902), .ZN(n14089) );
  NAND2_X1 U7698 ( .A1(n9490), .A2(n9489), .ZN(n12153) );
  NAND2_X2 U7699 ( .A1(n11605), .A2(n11604), .ZN(n14075) );
  OAI21_X1 U7700 ( .B1(n8821), .B2(n8045), .A(n8042), .ZN(n8846) );
  OAI21_X1 U7701 ( .B1(n8068), .B2(n8765), .A(n8067), .ZN(n8807) );
  NAND2_X1 U7702 ( .A1(n9206), .A2(n9205), .ZN(n9487) );
  OR2_X1 U7703 ( .A1(n11045), .A2(n11046), .ZN(n11265) );
  NAND2_X1 U7704 ( .A1(n8781), .A2(n8764), .ZN(n8765) );
  CLKBUF_X1 U7705 ( .A(n15295), .Z(n15333) );
  NAND2_X1 U7706 ( .A1(n8763), .A2(n10341), .ZN(n8781) );
  OR2_X1 U7707 ( .A1(n8763), .A2(n10341), .ZN(n8764) );
  XNOR2_X1 U7708 ( .A(n15941), .B(P3_ADDR_REG_8__SCAN_IN), .ZN(n15975) );
  NAND2_X1 U7709 ( .A1(n8058), .A2(n8059), .ZN(n8763) );
  NAND2_X1 U7710 ( .A1(n15939), .A2(n15940), .ZN(n15941) );
  NAND2_X1 U7711 ( .A1(n15099), .A2(n15312), .ZN(n15338) );
  AND2_X2 U7712 ( .A1(n10131), .A2(n14641), .ZN(n14571) );
  NAND2_X1 U7713 ( .A1(n7918), .A2(n7917), .ZN(n10765) );
  NAND2_X1 U7714 ( .A1(n8726), .A2(n8725), .ZN(n8729) );
  NAND2_X1 U7715 ( .A1(n8019), .A2(n11406), .ZN(n11411) );
  AND4_X1 U7716 ( .A1(n8561), .A2(n8560), .A3(n8559), .A4(n8558), .ZN(n8573)
         );
  OR2_X2 U7717 ( .A1(n10438), .A2(n10644), .ZN(n12377) );
  INV_X1 U7718 ( .A(n10851), .ZN(n16446) );
  AND3_X1 U7719 ( .A1(n9325), .A2(n9324), .A3(n9323), .ZN(n16429) );
  INV_X2 U7720 ( .A(n10644), .ZN(n12687) );
  AND2_X1 U7721 ( .A1(n9355), .A2(n9354), .ZN(n10851) );
  NAND3_X1 U7722 ( .A1(n8294), .A2(n10045), .A3(n10046), .ZN(n14320) );
  XNOR2_X1 U7723 ( .A(n7462), .B(n13995), .ZN(n10763) );
  AND3_X1 U7724 ( .A1(n7986), .A2(n10055), .A3(n8187), .ZN(n10542) );
  XNOR2_X1 U7725 ( .A(n8809), .B(P3_IR_REG_15__SCAN_IN), .ZN(n13292) );
  NAND2_X2 U7726 ( .A1(n10440), .A2(n10441), .ZN(n7468) );
  AND2_X1 U7727 ( .A1(n10437), .A2(n9976), .ZN(n7593) );
  AND4_X2 U7728 ( .A1(n9347), .A2(n9346), .A3(n9345), .A4(n9344), .ZN(n10915)
         );
  BUF_X2 U7729 ( .A(n13771), .Z(n7462) );
  AND2_X1 U7731 ( .A1(n10023), .A2(n10024), .ZN(n7949) );
  NAND2_X2 U7732 ( .A1(n12783), .A2(n9060), .ZN(n10927) );
  AND2_X1 U7733 ( .A1(n11549), .A2(n9841), .ZN(n10440) );
  CLKBUF_X1 U7734 ( .A(n12783), .Z(n7728) );
  INV_X1 U7735 ( .A(n9060), .ZN(n12285) );
  OR2_X1 U7736 ( .A1(n10057), .A2(n10017), .ZN(n10023) );
  CLKBUF_X1 U7737 ( .A(n9842), .Z(n7717) );
  INV_X1 U7738 ( .A(n10056), .ZN(n14191) );
  AND2_X2 U7739 ( .A1(n7707), .A2(n7704), .ZN(n15185) );
  NAND2_X1 U7740 ( .A1(n14800), .A2(n10020), .ZN(n13846) );
  OAI21_X1 U7741 ( .B1(n9310), .B2(n8196), .A(n9179), .ZN(n9319) );
  AND2_X1 U7742 ( .A1(n12593), .A2(n10019), .ZN(n10056) );
  AOI21_X1 U7743 ( .B1(n9177), .B2(n9176), .A(n9175), .ZN(n9310) );
  INV_X1 U7744 ( .A(n13369), .ZN(n10592) );
  NAND2_X1 U7745 ( .A1(n9099), .A2(n7499), .ZN(n8538) );
  BUF_X1 U7746 ( .A(n10018), .Z(n12593) );
  XNOR2_X1 U7747 ( .A(n8884), .B(P3_IR_REG_19__SCAN_IN), .ZN(n13369) );
  XNOR2_X1 U7748 ( .A(n10014), .B(n14793), .ZN(n10018) );
  OAI21_X1 U7749 ( .B1(n10171), .B2(n10225), .A(n7716), .ZN(n9189) );
  XNOR2_X1 U7750 ( .A(n10088), .B(n10087), .ZN(n11958) );
  NAND2_X1 U7751 ( .A1(n9207), .A2(n10208), .ZN(n9210) );
  AND2_X1 U7752 ( .A1(n8604), .A2(n8603), .ZN(n11015) );
  NAND2_X1 U7753 ( .A1(n10171), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7716) );
  OR2_X1 U7754 ( .A1(n15988), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n15926) );
  NAND2_X1 U7755 ( .A1(n10028), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10026) );
  NAND2_X2 U7756 ( .A1(n10197), .A2(P1_U3086), .ZN(n15916) );
  NAND2_X1 U7757 ( .A1(n7787), .A2(n7788), .ZN(n9058) );
  NAND2_X2 U7758 ( .A1(n10196), .A2(P2_U3088), .ZN(n14818) );
  NOR2_X1 U7759 ( .A1(n8317), .A2(n9156), .ZN(n7892) );
  NOR2_X1 U7760 ( .A1(n10027), .A2(n10015), .ZN(n7947) );
  OR2_X1 U7761 ( .A1(n10082), .A2(n10335), .ZN(n10085) );
  INV_X1 U7762 ( .A(n9574), .ZN(n7891) );
  NAND2_X1 U7763 ( .A1(n10027), .A2(n7683), .ZN(n8165) );
  NAND2_X2 U7764 ( .A1(n10196), .A2(P1_U3086), .ZN(n15919) );
  NOR2_X2 U7765 ( .A1(n8866), .A2(n7491), .ZN(n9054) );
  OAI21_X1 U7766 ( .B1(n10029), .B2(n7732), .A(n7731), .ZN(n9173) );
  AND4_X1 U7767 ( .A1(n7789), .A2(n7792), .A3(n7791), .A4(n7790), .ZN(n7788)
         );
  AND2_X1 U7768 ( .A1(n8411), .A2(n8526), .ZN(n7789) );
  OR2_X1 U7769 ( .A1(n7777), .A2(n8415), .ZN(n11228) );
  AND3_X2 U7770 ( .A1(n7928), .A2(n9952), .A3(n9951), .ZN(n8304) );
  NAND4_X1 U7771 ( .A1(n7928), .A2(n8136), .A3(n9952), .A4(n9951), .ZN(n10696)
         );
  XNOR2_X1 U7772 ( .A(n10050), .B(P2_IR_REG_2__SCAN_IN), .ZN(n16107) );
  AND2_X2 U7773 ( .A1(n8193), .A2(n8191), .ZN(n10029) );
  NAND4_X1 U7774 ( .A1(n9155), .A2(n9154), .A3(n8135), .A4(n9926), .ZN(n9933)
         );
  NAND4_X1 U7775 ( .A1(n15862), .A2(n7998), .A3(n7999), .A4(n7997), .ZN(n9352)
         );
  AND3_X1 U7776 ( .A1(n8731), .A2(n8529), .A3(n8669), .ZN(n7791) );
  AND2_X1 U7777 ( .A1(n8527), .A2(n8528), .ZN(n7792) );
  AND2_X1 U7778 ( .A1(n8412), .A2(n8530), .ZN(n8411) );
  INV_X1 U7779 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7997) );
  INV_X4 U7780 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7781 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7999) );
  NOR2_X1 U7782 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n9147) );
  INV_X1 U7783 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9926) );
  NOR2_X1 U7784 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n9150) );
  NOR2_X1 U7785 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n9148) );
  INV_X1 U7786 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8135) );
  INV_X1 U7787 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n15867) );
  NOR2_X1 U7788 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n8315) );
  NOR2_X1 U7789 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n8314) );
  NOR2_X1 U7790 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n9155) );
  INV_X1 U7791 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n15862) );
  NOR2_X1 U7792 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7898) );
  INV_X1 U7793 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n10010) );
  INV_X1 U7794 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8669) );
  INV_X1 U7795 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n10011) );
  INV_X1 U7796 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8412) );
  INV_X1 U7797 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8530) );
  NOR2_X1 U7798 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n8553) );
  INV_X1 U7799 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n10012) );
  INV_X1 U7800 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n11390) );
  NOR2_X1 U7801 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n8527) );
  NOR2_X1 U7802 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8528) );
  NOR2_X1 U7803 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n8526) );
  INV_X1 U7804 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9953) );
  NOR2_X1 U7805 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n7897) );
  INV_X1 U7806 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n10025) );
  INV_X1 U7807 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U7808 ( .A1(n9099), .A2(n7526), .ZN(n8547) );
  OR2_X1 U7809 ( .A1(n9724), .A2(n11123), .ZN(n9291) );
  NOR2_X1 U7810 ( .A1(n10696), .A2(n9954), .ZN(n10082) );
  OAI21_X1 U7811 ( .B1(n10696), .B2(n10078), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n10089) );
  NOR2_X2 U7812 ( .A1(n7733), .A2(n16315), .ZN(n16319) );
  NOR2_X2 U7813 ( .A1(n14548), .A2(n14688), .ZN(n7994) );
  NAND4_X2 U7814 ( .A1(n9371), .A2(n9370), .A3(n9369), .A4(n9368), .ZN(n14971)
         );
  OR2_X1 U7815 ( .A1(n14125), .A2(n14126), .ZN(n14127) );
  XNOR2_X2 U7816 ( .A(n16032), .B(n7982), .ZN(n16320) );
  NAND2_X2 U7817 ( .A1(n7983), .A2(n16030), .ZN(n16032) );
  OAI21_X2 U7818 ( .B1(n9265), .B2(P1_IR_REG_28__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9162) );
  NOR4_X2 U7819 ( .A1(n9919), .A2(n9918), .A3(n9917), .A4(n9916), .ZN(n9920)
         );
  NOR2_X2 U7820 ( .A1(n11817), .A2(n11818), .ZN(n11864) );
  NAND2_X1 U7821 ( .A1(n10927), .A2(n10171), .ZN(n7461) );
  INV_X1 U7822 ( .A(n10516), .ZN(n16394) );
  XNOR2_X2 U7823 ( .A(n15980), .B(n16363), .ZN(n15981) );
  XNOR2_X2 U7824 ( .A(n15930), .B(n15931), .ZN(n15980) );
  XNOR2_X2 U7825 ( .A(n16007), .B(n16008), .ZN(n16286) );
  NOR2_X2 U7826 ( .A1(n11683), .A2(n14075), .ZN(n11796) );
  NOR2_X2 U7827 ( .A1(n10516), .A2(n11126), .ZN(n10528) );
  NOR2_X2 U7828 ( .A1(n16027), .A2(n16028), .ZN(n16315) );
  NOR2_X2 U7829 ( .A1(n11247), .A2(n14060), .ZN(n7989) );
  XNOR2_X2 U7830 ( .A(n9264), .B(n9161), .ZN(n9943) );
  NAND2_X2 U7831 ( .A1(n14597), .A2(n14577), .ZN(n14578) );
  INV_X4 U7832 ( .A(n14004), .ZN(n14238) );
  AND2_X4 U7833 ( .A1(n13982), .A2(n10130), .ZN(n14004) );
  INV_X8 U7834 ( .A(n14238), .ZN(n14206) );
  INV_X1 U7835 ( .A(n10053), .ZN(n7464) );
  INV_X1 U7836 ( .A(n10053), .ZN(n7465) );
  BUF_X2 U7837 ( .A(n10042), .Z(n8296) );
  AND2_X2 U7838 ( .A1(n14282), .A2(n10125), .ZN(n10126) );
  NAND2_X2 U7839 ( .A1(n10083), .A2(n10084), .ZN(n14282) );
  INV_X1 U7840 ( .A(n8648), .ZN(n8078) );
  OR2_X1 U7841 ( .A1(n11515), .A2(n13015), .ZN(n11806) );
  NOR2_X1 U7842 ( .A1(n14430), .A2(n7953), .ZN(n7952) );
  INV_X1 U7843 ( .A(n14429), .ZN(n7953) );
  INV_X1 U7844 ( .A(n12551), .ZN(n9164) );
  NOR2_X1 U7845 ( .A1(n15327), .A2(n8436), .ZN(n8434) );
  AND2_X1 U7846 ( .A1(n8287), .A2(n9341), .ZN(n8285) );
  INV_X1 U7847 ( .A(n14118), .ZN(n8506) );
  AND2_X1 U7848 ( .A1(n8270), .A2(n9718), .ZN(n8269) );
  NAND2_X1 U7849 ( .A1(n8272), .A2(n8271), .ZN(n8270) );
  AND2_X1 U7850 ( .A1(n14152), .A2(n14153), .ZN(n7968) );
  INV_X1 U7851 ( .A(n14165), .ZN(n8489) );
  INV_X1 U7852 ( .A(n8405), .ZN(n8403) );
  OAI21_X1 U7853 ( .B1(n7849), .B2(n7852), .A(n9232), .ZN(n9637) );
  INV_X1 U7854 ( .A(n9228), .ZN(n7849) );
  INV_X1 U7855 ( .A(n8072), .ZN(n8071) );
  NAND2_X1 U7856 ( .A1(n12976), .A2(n12961), .ZN(n8075) );
  AOI211_X1 U7857 ( .C1(n12973), .C2(n12974), .A(n12972), .B(n12961), .ZN(
        n8072) );
  AND2_X1 U7858 ( .A1(n11411), .A2(n7565), .ZN(n7761) );
  INV_X1 U7859 ( .A(n7799), .ZN(n7798) );
  OAI21_X1 U7860 ( .B1(n8876), .B2(n7800), .A(n8894), .ZN(n7799) );
  OR2_X1 U7861 ( .A1(n13085), .A2(n13540), .ZN(n13012) );
  OR2_X1 U7862 ( .A1(n12855), .A2(n9138), .ZN(n10593) );
  NAND3_X1 U7863 ( .A1(n7867), .A2(n7868), .A3(n8547), .ZN(n9060) );
  NAND2_X1 U7864 ( .A1(n8638), .A2(n7869), .ZN(n7868) );
  NAND2_X1 U7865 ( .A1(n9053), .A2(n9091), .ZN(n8355) );
  INV_X1 U7866 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9052) );
  INV_X1 U7867 ( .A(n13926), .ZN(n8161) );
  NAND2_X1 U7868 ( .A1(n12593), .A2(n14800), .ZN(n10057) );
  NOR2_X1 U7869 ( .A1(n11677), .A2(n8184), .ZN(n8183) );
  INV_X1 U7870 ( .A(n11502), .ZN(n8184) );
  NAND2_X1 U7871 ( .A1(n7948), .A2(n11656), .ZN(n10043) );
  OR2_X1 U7872 ( .A1(n10086), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n9963) );
  AND2_X1 U7873 ( .A1(n14857), .A2(n14858), .ZN(n12650) );
  NAND2_X1 U7874 ( .A1(n12650), .A2(n14851), .ZN(n8122) );
  INV_X1 U7875 ( .A(n9843), .ZN(n9326) );
  NAND2_X1 U7876 ( .A1(n10442), .A2(n7817), .ZN(n10445) );
  INV_X1 U7877 ( .A(n7818), .ZN(n7817) );
  OR2_X1 U7878 ( .A1(n12377), .A2(n10439), .ZN(n10442) );
  NAND2_X1 U7879 ( .A1(n7815), .A2(n7814), .ZN(n10486) );
  OR2_X1 U7880 ( .A1(n7468), .A2(n10439), .ZN(n7814) );
  INV_X1 U7881 ( .A(n7816), .ZN(n7815) );
  OAI21_X1 U7882 ( .B1(n10644), .B2(n11207), .A(n10444), .ZN(n7816) );
  NAND2_X1 U7883 ( .A1(n15382), .A2(n15147), .ZN(n8473) );
  NAND2_X1 U7884 ( .A1(n8441), .A2(n8438), .ZN(n15157) );
  INV_X1 U7885 ( .A(n8439), .ZN(n8438) );
  OAI21_X1 U7886 ( .B1(n8440), .B2(n8445), .A(n15161), .ZN(n8439) );
  NOR2_X1 U7887 ( .A1(n7487), .A2(n8480), .ZN(n8479) );
  AND2_X1 U7888 ( .A1(n15237), .A2(n12561), .ZN(n8342) );
  NOR2_X1 U7889 ( .A1(n8009), .A2(n15446), .ZN(n8008) );
  INV_X1 U7890 ( .A(n8010), .ZN(n8009) );
  NAND2_X1 U7891 ( .A1(n10888), .A2(n10887), .ZN(n10890) );
  NAND2_X1 U7892 ( .A1(n7627), .A2(n12567), .ZN(n8325) );
  INV_X1 U7893 ( .A(n8233), .ZN(n8232) );
  INV_X1 U7894 ( .A(n9677), .ZN(n9244) );
  XNOR2_X1 U7895 ( .A(n9226), .B(n15520), .ZN(n9572) );
  OAI21_X1 U7896 ( .B1(n9487), .B2(n7859), .A(n7857), .ZN(n9573) );
  INV_X1 U7897 ( .A(n7860), .ZN(n7859) );
  AOI21_X1 U7898 ( .B1(n7860), .B2(n7866), .A(n7858), .ZN(n7857) );
  NOR2_X1 U7899 ( .A1(n7861), .A2(n8221), .ZN(n7860) );
  AND2_X1 U7900 ( .A1(n9224), .A2(n9223), .ZN(n9557) );
  AOI21_X1 U7901 ( .B1(n8200), .B2(n8202), .A(n7549), .ZN(n8198) );
  NOR2_X1 U7902 ( .A1(n15972), .A2(n15971), .ZN(n15949) );
  NOR2_X1 U7903 ( .A1(n11471), .A2(n8392), .ZN(n8391) );
  INV_X1 U7904 ( .A(n8393), .ZN(n8392) );
  INV_X1 U7905 ( .A(n13220), .ZN(n12124) );
  NAND2_X1 U7906 ( .A1(n12480), .A2(n7744), .ZN(n12491) );
  OR2_X1 U7907 ( .A1(n12481), .A2(n12482), .ZN(n7744) );
  NAND2_X1 U7908 ( .A1(n7757), .A2(n11042), .ZN(n7760) );
  NAND2_X1 U7909 ( .A1(n11411), .A2(n11035), .ZN(n7757) );
  OAI21_X1 U7910 ( .B1(n13270), .B2(n8243), .A(n7752), .ZN(n13315) );
  NAND2_X1 U7911 ( .A1(n8246), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8243) );
  NAND2_X1 U7912 ( .A1(n13294), .A2(n8246), .ZN(n7752) );
  INV_X1 U7913 ( .A(n13297), .ZN(n8246) );
  OAI21_X1 U7914 ( .B1(n12978), .B2(n13404), .A(n9037), .ZN(n13387) );
  NAND2_X1 U7915 ( .A1(n13427), .A2(n8400), .ZN(n13416) );
  NOR2_X1 U7916 ( .A1(n13413), .A2(n12846), .ZN(n8400) );
  OR2_X1 U7917 ( .A1(n13486), .A2(n13100), .ZN(n13462) );
  NAND2_X1 U7918 ( .A1(n8841), .A2(n8840), .ZN(n13566) );
  NOR2_X1 U7919 ( .A1(n12888), .A2(n8077), .ZN(n8076) );
  NOR2_X1 U7920 ( .A1(n8647), .A2(n8078), .ZN(n8077) );
  AOI21_X1 U7921 ( .B1(n8398), .B2(n12888), .A(n7534), .ZN(n8397) );
  NOR2_X1 U7922 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8610) );
  NAND2_X1 U7923 ( .A1(n13401), .A2(n13413), .ZN(n13403) );
  OR2_X1 U7924 ( .A1(n13064), .A2(n12855), .ZN(n16558) );
  XNOR2_X1 U7925 ( .A(n8539), .B(P3_IR_REG_29__SCAN_IN), .ZN(n8540) );
  XNOR2_X1 U7926 ( .A(n8081), .B(n8546), .ZN(n12783) );
  NAND2_X1 U7927 ( .A1(n8547), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8081) );
  INV_X1 U7928 ( .A(n8056), .ZN(n8055) );
  OAI21_X1 U7929 ( .B1(n8863), .B2(n8057), .A(n8881), .ZN(n8056) );
  INV_X1 U7930 ( .A(n8062), .ZN(n8061) );
  OAI21_X1 U7931 ( .B1(n8728), .B2(n8063), .A(n8743), .ZN(n8062) );
  INV_X1 U7932 ( .A(n8050), .ZN(n8049) );
  OAI21_X1 U7933 ( .B1(n8676), .B2(n8051), .A(n8693), .ZN(n8050) );
  AOI21_X1 U7934 ( .B1(n8039), .B2(n8041), .A(n7554), .ZN(n8037) );
  NAND2_X1 U7935 ( .A1(n8415), .A2(n8523), .ZN(n8554) );
  INV_X1 U7936 ( .A(n12524), .ZN(n12522) );
  NOR2_X1 U7937 ( .A1(n7924), .A2(n8151), .ZN(n7921) );
  INV_X1 U7938 ( .A(n12368), .ZN(n8151) );
  NOR2_X2 U7939 ( .A1(n14460), .A2(n14664), .ZN(n14419) );
  NAND2_X1 U7940 ( .A1(n8297), .A2(n8298), .ZN(n14459) );
  AOI21_X1 U7941 ( .B1(n8299), .B2(n14445), .A(n7474), .ZN(n8298) );
  NAND2_X1 U7942 ( .A1(n8302), .A2(n14444), .ZN(n8301) );
  NAND2_X1 U7943 ( .A1(n14409), .A2(n14408), .ZN(n14470) );
  AND2_X1 U7944 ( .A1(n7505), .A2(n14406), .ZN(n8188) );
  NOR2_X1 U7945 ( .A1(n14502), .A2(n8190), .ZN(n8189) );
  INV_X1 U7946 ( .A(n14405), .ZN(n8190) );
  AOI21_X1 U7947 ( .B1(n7952), .B2(n14610), .A(n7550), .ZN(n7951) );
  OAI21_X2 U7948 ( .B1(n11772), .B2(n7490), .A(n11773), .ZN(n11940) );
  CLKBUF_X1 U7949 ( .A(n10053), .Z(n14202) );
  INV_X2 U7950 ( .A(n8296), .ZN(n10048) );
  NAND2_X1 U7951 ( .A1(n11665), .A2(n11664), .ZN(n7827) );
  AND4_X1 U7952 ( .A1(n9852), .A2(n9851), .A3(n9850), .A4(n9849), .ZN(n15112)
         );
  NAND2_X1 U7953 ( .A1(n12551), .A2(n15909), .ZN(n9303) );
  OR2_X1 U7954 ( .A1(n9843), .A2(n10315), .ZN(n9280) );
  OR2_X1 U7955 ( .A1(n9467), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n9501) );
  OR2_X1 U7956 ( .A1(n15371), .A2(n15112), .ZN(n15089) );
  NAND2_X1 U7957 ( .A1(n9889), .A2(n14939), .ZN(n8338) );
  OAI21_X1 U7958 ( .B1(n15142), .B2(n8464), .A(n8465), .ZN(n15107) );
  NAND2_X1 U7959 ( .A1(n8468), .A2(n8472), .ZN(n8464) );
  AOI21_X1 U7960 ( .B1(n8468), .B2(n8467), .A(n8466), .ZN(n8465) );
  INV_X1 U7961 ( .A(n15110), .ZN(n8466) );
  INV_X1 U7962 ( .A(n15142), .ZN(n8463) );
  NAND2_X1 U7963 ( .A1(n15306), .A2(n7698), .ZN(n15281) );
  OR2_X1 U7964 ( .A1(n15446), .A2(n15330), .ZN(n7698) );
  AOI21_X1 U7965 ( .B1(n8434), .B2(n12552), .A(n7535), .ZN(n8432) );
  INV_X1 U7966 ( .A(n8434), .ZN(n8433) );
  INV_X1 U7967 ( .A(n8328), .ZN(n8327) );
  OAI21_X1 U7968 ( .B1(n8329), .B2(n12554), .A(n12556), .ZN(n8328) );
  CLKBUF_X2 U7969 ( .A(n9350), .Z(n9679) );
  INV_X1 U7970 ( .A(n9796), .ZN(n9350) );
  INV_X1 U7971 ( .A(n16258), .ZN(n10495) );
  NAND2_X1 U7972 ( .A1(n7540), .A2(n9153), .ZN(n9156) );
  INV_X1 U7973 ( .A(n9574), .ZN(n9158) );
  AND2_X1 U7974 ( .A1(n8134), .A2(n9154), .ZN(n8133) );
  INV_X4 U7975 ( .A(n10196), .ZN(n10171) );
  AND2_X1 U7976 ( .A1(n13370), .A2(n8018), .ZN(n8017) );
  INV_X1 U7977 ( .A(n7806), .ZN(n7803) );
  NAND2_X1 U7978 ( .A1(n12521), .A2(n12534), .ZN(n13776) );
  NAND2_X1 U7979 ( .A1(n9273), .A2(n7633), .ZN(n7707) );
  NOR2_X1 U7980 ( .A1(n7706), .A2(n7705), .ZN(n7704) );
  NOR2_X1 U7981 ( .A1(n15692), .A2(n9361), .ZN(n7633) );
  NAND2_X1 U7982 ( .A1(n9301), .A2(n7710), .ZN(n7709) );
  NAND2_X1 U7983 ( .A1(n9300), .A2(n9338), .ZN(n7708) );
  NAND2_X1 U7984 ( .A1(n9357), .A2(n9356), .ZN(n8287) );
  NAND2_X1 U7985 ( .A1(n7644), .A2(n7643), .ZN(n9356) );
  NAND2_X1 U7986 ( .A1(n9372), .A2(n14972), .ZN(n7643) );
  NAND2_X1 U7987 ( .A1(n9413), .A2(n16446), .ZN(n7644) );
  CLKBUF_X1 U7988 ( .A(n9338), .Z(n9413) );
  NAND2_X1 U7989 ( .A1(n9377), .A2(n9376), .ZN(n9393) );
  INV_X1 U7990 ( .A(n14020), .ZN(n7672) );
  NOR2_X1 U7991 ( .A1(n9432), .A2(n9431), .ZN(n7666) );
  INV_X1 U7992 ( .A(n14047), .ZN(n8495) );
  INV_X1 U7993 ( .A(n14063), .ZN(n8499) );
  INV_X1 U7994 ( .A(n14086), .ZN(n8486) );
  INV_X1 U7995 ( .A(n14103), .ZN(n7638) );
  INV_X1 U7996 ( .A(n14105), .ZN(n7636) );
  OAI21_X1 U7997 ( .B1(n7492), .B2(n7674), .A(n7959), .ZN(n14136) );
  NAND2_X1 U7998 ( .A1(n7548), .A2(n14131), .ZN(n7959) );
  INV_X1 U7999 ( .A(n14142), .ZN(n8487) );
  NAND2_X1 U8000 ( .A1(n9698), .A2(n9701), .ZN(n8271) );
  NAND2_X1 U8001 ( .A1(n9689), .A2(n9688), .ZN(n9699) );
  NOR2_X1 U8002 ( .A1(n9701), .A2(n9698), .ZN(n8272) );
  NAND2_X1 U8003 ( .A1(n7967), .A2(n7966), .ZN(n7965) );
  INV_X1 U8004 ( .A(n14152), .ZN(n7966) );
  INV_X1 U8005 ( .A(n14153), .ZN(n7967) );
  NAND2_X1 U8006 ( .A1(n14161), .A2(n7964), .ZN(n7963) );
  AND2_X1 U8007 ( .A1(n7961), .A2(n14159), .ZN(n7960) );
  INV_X1 U8008 ( .A(n7968), .ZN(n7964) );
  AOI21_X1 U8009 ( .B1(n7852), .B2(n9232), .A(n9234), .ZN(n7850) );
  NAND2_X1 U8010 ( .A1(n7850), .A2(n7851), .ZN(n7848) );
  INV_X1 U8011 ( .A(n9232), .ZN(n7851) );
  NAND2_X1 U8012 ( .A1(n7853), .A2(n9227), .ZN(n7852) );
  INV_X1 U8013 ( .A(n9594), .ZN(n7853) );
  NOR2_X1 U8014 ( .A1(n9083), .A2(n8086), .ZN(n8085) );
  INV_X1 U8015 ( .A(n8974), .ZN(n8086) );
  NAND2_X1 U8016 ( .A1(n9003), .A2(n8084), .ZN(n8083) );
  INV_X1 U8017 ( .A(n8990), .ZN(n8084) );
  INV_X1 U8018 ( .A(n12944), .ZN(n8351) );
  INV_X1 U8019 ( .A(n12921), .ZN(n8402) );
  NAND2_X1 U8020 ( .A1(n12597), .A2(n12596), .ZN(n8130) );
  NAND3_X1 U8021 ( .A1(n9903), .A2(n9918), .A3(n9916), .ZN(n9872) );
  INV_X1 U8022 ( .A(n12563), .ZN(n7880) );
  NAND2_X1 U8023 ( .A1(n9229), .A2(n15717), .ZN(n9232) );
  AND2_X1 U8024 ( .A1(n7864), .A2(n9216), .ZN(n7863) );
  AND2_X1 U8025 ( .A1(n8229), .A2(n8517), .ZN(n8228) );
  NAND2_X1 U8026 ( .A1(n9486), .A2(n9210), .ZN(n8229) );
  OAI21_X1 U8027 ( .B1(n9106), .B2(P3_D_REG_0__SCAN_IN), .A(n10378), .ZN(
        n10591) );
  NAND2_X1 U8028 ( .A1(n8022), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8021) );
  OAI21_X1 U8029 ( .B1(n10970), .B2(n8241), .A(n8240), .ZN(n11012) );
  INV_X1 U8030 ( .A(n8237), .ZN(n8240) );
  OAI21_X1 U8031 ( .B1(n11284), .B2(n8238), .A(n7482), .ZN(n8237) );
  NAND2_X1 U8032 ( .A1(n11433), .A2(n11432), .ZN(n7756) );
  NAND2_X1 U8033 ( .A1(n11420), .A2(n11419), .ZN(n11422) );
  NOR2_X1 U8034 ( .A1(n13260), .A2(n13261), .ZN(n13282) );
  NAND2_X1 U8035 ( .A1(n13451), .A2(n8085), .ZN(n13435) );
  NAND2_X1 U8036 ( .A1(n8938), .A2(n15585), .ZN(n8952) );
  AND2_X1 U8037 ( .A1(n7798), .A2(n8912), .ZN(n7796) );
  INV_X1 U8038 ( .A(n8095), .ZN(n8094) );
  OAI21_X1 U8039 ( .B1(n8097), .B2(n8096), .A(n12808), .ZN(n8095) );
  NAND2_X1 U8040 ( .A1(n7796), .A2(n7800), .ZN(n7795) );
  INV_X1 U8041 ( .A(n8877), .ZN(n7800) );
  NOR2_X1 U8042 ( .A1(n13512), .A2(n8098), .ZN(n8097) );
  INV_X1 U8043 ( .A(n8895), .ZN(n8098) );
  AND2_X1 U8044 ( .A1(n13564), .A2(n8410), .ZN(n8409) );
  NAND2_X1 U8045 ( .A1(n13575), .A2(n12929), .ZN(n8410) );
  NOR2_X1 U8046 ( .A1(n13557), .A2(n12935), .ZN(n8080) );
  NAND2_X1 U8047 ( .A1(n12034), .A2(n8698), .ZN(n8093) );
  NOR2_X1 U8048 ( .A1(n8362), .A2(n8358), .ZN(n8357) );
  INV_X1 U8049 ( .A(n13018), .ZN(n8358) );
  INV_X1 U8050 ( .A(n12871), .ZN(n8361) );
  AOI21_X1 U8051 ( .B1(n8349), .B2(n8350), .A(n8348), .ZN(n8347) );
  INV_X1 U8052 ( .A(n13012), .ZN(n8348) );
  NAND2_X1 U8053 ( .A1(n13226), .A2(n8592), .ZN(n12865) );
  NAND2_X1 U8054 ( .A1(n16402), .A2(n16373), .ZN(n12867) );
  INV_X1 U8055 ( .A(n8355), .ZN(n8353) );
  NAND2_X1 U8056 ( .A1(n8052), .A2(n8053), .ZN(n8899) );
  AOI21_X1 U8057 ( .B1(n8055), .B2(n8057), .A(n8054), .ZN(n8053) );
  INV_X1 U8058 ( .A(n8897), .ZN(n8054) );
  NAND2_X1 U8059 ( .A1(n8913), .A2(n8036), .ZN(n7623) );
  INV_X1 U8060 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8829) );
  INV_X1 U8061 ( .A(n8820), .ZN(n8044) );
  INV_X1 U8062 ( .A(n8641), .ZN(n8041) );
  NOR2_X1 U8063 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8419) );
  OR2_X1 U8064 ( .A1(n10734), .A2(n10751), .ZN(n10743) );
  INV_X1 U8065 ( .A(n10018), .ZN(n10020) );
  OR2_X1 U8066 ( .A1(n13827), .A2(n13930), .ZN(n13829) );
  NAND2_X1 U8067 ( .A1(n14270), .A2(n12450), .ZN(n7934) );
  INV_X1 U8068 ( .A(n14630), .ZN(n8173) );
  INV_X1 U8069 ( .A(n8177), .ZN(n8176) );
  OAI21_X1 U8070 ( .B1(n14264), .B2(n8178), .A(n14265), .ZN(n8177) );
  OR2_X1 U8071 ( .A1(n10743), .A2(n10997), .ZN(n10989) );
  INV_X1 U8072 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8136) );
  NOR2_X1 U8073 ( .A1(n10333), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n10338) );
  OR2_X1 U8074 ( .A1(n10288), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n10333) );
  OR2_X1 U8075 ( .A1(n10067), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n10201) );
  AND2_X1 U8076 ( .A1(n12383), .A2(n12384), .ZN(n8132) );
  AOI21_X1 U8077 ( .B1(n8131), .B2(n8130), .A(n12599), .ZN(n12602) );
  NOR2_X1 U8078 ( .A1(n15371), .A2(n9889), .ZN(n8003) );
  OR2_X1 U8079 ( .A1(n15440), .A2(n14880), .ZN(n12558) );
  NOR2_X1 U8080 ( .A1(n8329), .A2(n12339), .ZN(n8326) );
  NAND2_X1 U8081 ( .A1(n8327), .A2(n8430), .ZN(n7887) );
  INV_X1 U8082 ( .A(n10440), .ZN(n10437) );
  NOR2_X1 U8083 ( .A1(n8322), .A2(n12157), .ZN(n8321) );
  NOR2_X1 U8084 ( .A1(n12151), .A2(n8323), .ZN(n8322) );
  INV_X1 U8085 ( .A(n12154), .ZN(n8323) );
  OR2_X2 U8086 ( .A1(n10890), .A2(n10889), .ZN(n11539) );
  OR2_X1 U8087 ( .A1(n16429), .A2(n14973), .ZN(n10857) );
  XNOR2_X1 U8088 ( .A(n14973), .B(n14843), .ZN(n11113) );
  NAND2_X1 U8089 ( .A1(n15179), .A2(n7501), .ZN(n15160) );
  INV_X1 U8090 ( .A(n9749), .ZN(n8236) );
  NAND2_X1 U8091 ( .A1(n9241), .A2(SI_20_), .ZN(n9242) );
  AND2_X1 U8092 ( .A1(n8288), .A2(n7840), .ZN(n9598) );
  OR2_X1 U8093 ( .A1(n9573), .A2(n9225), .ZN(n9228) );
  INV_X1 U8094 ( .A(n8228), .ZN(n8227) );
  AOI21_X1 U8095 ( .B1(n8228), .B2(n8226), .A(n8225), .ZN(n8224) );
  INV_X1 U8096 ( .A(n9214), .ZN(n8225) );
  INV_X1 U8097 ( .A(n9210), .ZN(n8226) );
  NAND2_X1 U8098 ( .A1(n9197), .A2(n9196), .ZN(n9425) );
  INV_X1 U8099 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n15977) );
  OR2_X1 U8100 ( .A1(n15938), .A2(n15937), .ZN(n15940) );
  OR2_X1 U8101 ( .A1(n16006), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n15939) );
  NOR2_X1 U8102 ( .A1(n15961), .A2(n15960), .ZN(n15962) );
  AND2_X1 U8103 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n16025), .ZN(n15960) );
  NAND2_X1 U8104 ( .A1(n12818), .A2(n13454), .ZN(n8414) );
  AOI21_X1 U8105 ( .B1(n13073), .B2(n12830), .A(n12833), .ZN(n8385) );
  AND2_X1 U8106 ( .A1(n12828), .A2(n12826), .ZN(n13108) );
  AND2_X1 U8107 ( .A1(n13107), .A2(n12821), .ZN(n13134) );
  OR2_X1 U8108 ( .A1(n8952), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8968) );
  NOR2_X1 U8109 ( .A1(n8508), .A2(n12489), .ZN(n12490) );
  NOR2_X1 U8110 ( .A1(n8753), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8772) );
  AOI21_X1 U8111 ( .B1(n8388), .B2(n8390), .A(n8387), .ZN(n8386) );
  INV_X1 U8112 ( .A(n11645), .ZN(n8387) );
  INV_X1 U8113 ( .A(n8377), .ZN(n8376) );
  OAI21_X1 U8114 ( .B1(n12490), .B2(n8378), .A(n12787), .ZN(n8377) );
  INV_X1 U8115 ( .A(n12494), .ZN(n8378) );
  NAND2_X1 U8116 ( .A1(n7621), .A2(n7511), .ZN(n7620) );
  NAND2_X1 U8117 ( .A1(n8421), .A2(n8422), .ZN(n7621) );
  AND2_X1 U8118 ( .A1(n13054), .A2(n13055), .ZN(n8420) );
  XNOR2_X1 U8119 ( .A(n7736), .B(n10592), .ZN(n13045) );
  NAND2_X1 U8120 ( .A1(n7497), .A2(n7737), .ZN(n7736) );
  NOR2_X1 U8121 ( .A1(n13043), .A2(n13050), .ZN(n7737) );
  XNOR2_X1 U8122 ( .A(n10921), .B(n11228), .ZN(n11222) );
  OAI21_X1 U8123 ( .B1(n11228), .B2(n16335), .A(n7776), .ZN(n11212) );
  NAND2_X1 U8124 ( .A1(n8415), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7776) );
  OAI211_X1 U8125 ( .C1(n10959), .C2(n8025), .A(n8024), .B(n11288), .ZN(n11293) );
  NAND2_X1 U8126 ( .A1(n11289), .A2(n16426), .ZN(n8024) );
  INV_X1 U8127 ( .A(n11289), .ZN(n8025) );
  NAND2_X1 U8128 ( .A1(n11293), .A2(n7769), .ZN(n8022) );
  NOR2_X1 U8129 ( .A1(n7770), .A2(n11017), .ZN(n7769) );
  INV_X1 U8130 ( .A(n11016), .ZN(n7770) );
  NAND2_X1 U8131 ( .A1(n11018), .A2(n11017), .ZN(n11407) );
  NAND2_X1 U8132 ( .A1(n11293), .A2(n11016), .ZN(n11018) );
  OR2_X1 U8133 ( .A1(n8021), .A2(n8020), .ZN(n11409) );
  INV_X1 U8134 ( .A(n11407), .ZN(n8020) );
  INV_X1 U8135 ( .A(n7761), .ZN(n7758) );
  NAND2_X1 U8136 ( .A1(n7760), .A2(n7759), .ZN(n11274) );
  NAND2_X1 U8137 ( .A1(n7762), .A2(n11042), .ZN(n11272) );
  NAND2_X1 U8138 ( .A1(n11411), .A2(n11035), .ZN(n7762) );
  NAND2_X1 U8139 ( .A1(n7729), .A2(n11439), .ZN(n7767) );
  INV_X1 U8140 ( .A(n11422), .ZN(n7729) );
  NOR2_X1 U8141 ( .A1(n11992), .A2(n8027), .ZN(n12183) );
  AND2_X1 U8142 ( .A1(n12006), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8027) );
  AND2_X1 U8143 ( .A1(n12185), .A2(n7872), .ZN(n12191) );
  NAND2_X1 U8144 ( .A1(n12186), .A2(n12196), .ZN(n7872) );
  NAND2_X1 U8145 ( .A1(n12191), .A2(n12190), .ZN(n12288) );
  XNOR2_X1 U8146 ( .A(n13229), .B(n8029), .ZN(n12295) );
  NOR2_X1 U8147 ( .A1(n12293), .A2(n8030), .ZN(n13229) );
  AND2_X1 U8148 ( .A1(n12294), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8030) );
  NOR2_X1 U8149 ( .A1(n13238), .A2(n13239), .ZN(n13260) );
  INV_X1 U8150 ( .A(n8247), .ZN(n13245) );
  OAI21_X1 U8151 ( .B1(n12284), .B2(n7784), .A(n7783), .ZN(n13267) );
  NAND2_X1 U8152 ( .A1(n7785), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7784) );
  NAND2_X1 U8153 ( .A1(n13247), .A2(n7785), .ZN(n7783) );
  INV_X1 U8154 ( .A(n13249), .ZN(n7785) );
  NOR2_X1 U8155 ( .A1(n13291), .A2(n13292), .ZN(n13294) );
  OR2_X1 U8156 ( .A1(n13270), .A2(n13269), .ZN(n8245) );
  OR2_X1 U8157 ( .A1(n8826), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n8827) );
  NOR2_X1 U8158 ( .A1(n13254), .A2(n13655), .ZN(n8028) );
  OR2_X1 U8159 ( .A1(n13329), .A2(n13330), .ZN(n7781) );
  NAND2_X1 U8160 ( .A1(n7781), .A2(n7780), .ZN(n8259) );
  INV_X1 U8161 ( .A(n13332), .ZN(n7780) );
  NAND2_X1 U8162 ( .A1(n13434), .A2(n9085), .ZN(n13427) );
  NAND2_X1 U8163 ( .A1(n7514), .A2(n9083), .ZN(n13434) );
  AND4_X1 U8164 ( .A1(n8994), .A2(n8993), .A3(n8992), .A4(n8991), .ZN(n13438)
         );
  AOI21_X1 U8165 ( .B1(n8945), .B2(n7594), .A(n7472), .ZN(n13465) );
  AND4_X1 U8166 ( .A1(n8924), .A2(n8923), .A3(n8922), .A4(n8921), .ZN(n13514)
         );
  NAND2_X1 U8167 ( .A1(n7797), .A2(n7798), .ZN(n8896) );
  OR2_X1 U8168 ( .A1(n13534), .A2(n7800), .ZN(n7797) );
  NAND2_X1 U8169 ( .A1(n8896), .A2(n8097), .ZN(n13516) );
  NAND2_X1 U8170 ( .A1(n8904), .A2(n8903), .ZN(n13142) );
  NAND2_X1 U8171 ( .A1(n13534), .A2(n8876), .ZN(n13537) );
  AND2_X1 U8172 ( .A1(n13575), .A2(n8802), .ZN(n7812) );
  NAND2_X1 U8173 ( .A1(n12465), .A2(n12464), .ZN(n7813) );
  INV_X1 U8174 ( .A(n13034), .ZN(n12464) );
  AND2_X1 U8175 ( .A1(n7567), .A2(n12895), .ZN(n8405) );
  AND2_X1 U8176 ( .A1(n12905), .A2(n12246), .ZN(n9073) );
  AND2_X1 U8177 ( .A1(n12921), .A2(n12917), .ZN(n13027) );
  INV_X1 U8178 ( .A(n13219), .ZN(n12323) );
  NOR2_X1 U8179 ( .A1(n13022), .A2(n7802), .ZN(n7801) );
  INV_X1 U8180 ( .A(n8662), .ZN(n7802) );
  INV_X1 U8181 ( .A(n13221), .ZN(n12892) );
  NAND2_X1 U8182 ( .A1(n11806), .A2(n8647), .ZN(n11809) );
  INV_X1 U8183 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n15774) );
  AND4_X1 U8184 ( .A1(n8615), .A2(n8614), .A3(n8613), .A4(n8612), .ZN(n11805)
         );
  NAND2_X1 U8185 ( .A1(n11303), .A2(n13018), .ZN(n11302) );
  AND4_X1 U8186 ( .A1(n8598), .A2(n8597), .A3(n8596), .A4(n8595), .ZN(n11650)
         );
  AND2_X1 U8187 ( .A1(n12871), .A2(n12870), .ZN(n13018) );
  NAND2_X1 U8188 ( .A1(n10609), .A2(n13737), .ZN(n10924) );
  AND2_X1 U8189 ( .A1(n10655), .A2(n13369), .ZN(n13060) );
  INV_X1 U8190 ( .A(n9047), .ZN(n13380) );
  NAND2_X1 U8191 ( .A1(n7496), .A2(n13452), .ZN(n13451) );
  OAI21_X1 U8192 ( .B1(n13483), .B2(n9079), .A(n9081), .ZN(n13448) );
  NOR2_X1 U8193 ( .A1(n8511), .A2(n8510), .ZN(n9081) );
  INV_X1 U8194 ( .A(n16374), .ZN(n13500) );
  NAND2_X1 U8195 ( .A1(n8887), .A2(n8886), .ZN(n13085) );
  INV_X1 U8196 ( .A(n12326), .ZN(n16513) );
  NAND2_X1 U8197 ( .A1(n11804), .A2(n13023), .ZN(n11803) );
  OR2_X1 U8198 ( .A1(n10617), .A2(n12975), .ZN(n16374) );
  INV_X1 U8199 ( .A(n13582), .ZN(n16377) );
  INV_X1 U8200 ( .A(n16558), .ZN(n16471) );
  NAND2_X1 U8201 ( .A1(n10617), .A2(n12961), .ZN(n16372) );
  NAND2_X1 U8202 ( .A1(n8996), .A2(n8995), .ZN(n8999) );
  INV_X1 U8203 ( .A(n9102), .ZN(n7617) );
  NOR2_X1 U8204 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), .ZN(
        n7616) );
  NOR2_X1 U8205 ( .A1(n8355), .A2(P3_IR_REG_23__SCAN_IN), .ZN(n8354) );
  XNOR2_X1 U8206 ( .A(n9057), .B(P3_IR_REG_21__SCAN_IN), .ZN(n12855) );
  NAND2_X1 U8207 ( .A1(n8900), .A2(n8035), .ZN(n8914) );
  INV_X1 U8208 ( .A(n7623), .ZN(n8035) );
  XNOR2_X1 U8209 ( .A(n9059), .B(P3_IR_REG_20__SCAN_IN), .ZN(n9138) );
  AND2_X1 U8210 ( .A1(n8897), .A2(n8880), .ZN(n8881) );
  INV_X1 U8211 ( .A(n8878), .ZN(n8057) );
  AND2_X1 U8212 ( .A1(n8878), .A2(n8862), .ZN(n8863) );
  NAND2_X1 U8213 ( .A1(n8864), .A2(n8863), .ZN(n8879) );
  AND2_X1 U8214 ( .A1(n8842), .A2(n8822), .ZN(n8823) );
  INV_X1 U8215 ( .A(n8065), .ZN(n8067) );
  OAI21_X1 U8216 ( .B1(n8781), .B2(n8070), .A(n8803), .ZN(n8065) );
  AND2_X1 U8217 ( .A1(n8820), .A2(n8805), .ZN(n8806) );
  OR2_X1 U8218 ( .A1(n8765), .A2(n10340), .ZN(n8782) );
  AND2_X1 U8219 ( .A1(n8761), .A2(n8742), .ZN(n8743) );
  INV_X1 U8220 ( .A(n8740), .ZN(n8063) );
  AND2_X1 U8221 ( .A1(n8740), .A2(n8727), .ZN(n8728) );
  NAND2_X1 U8222 ( .A1(n8729), .A2(n8728), .ZN(n8741) );
  AND2_X1 U8223 ( .A1(n8706), .A2(n8692), .ZN(n8693) );
  INV_X1 U8224 ( .A(n8690), .ZN(n8051) );
  AND2_X1 U8225 ( .A1(n8690), .A2(n8675), .ZN(n8676) );
  NAND2_X1 U8226 ( .A1(n8677), .A2(n8676), .ZN(n8691) );
  NAND2_X1 U8227 ( .A1(n8419), .A2(n8523), .ZN(n8418) );
  NAND2_X1 U8228 ( .A1(n8524), .A2(n8415), .ZN(n8416) );
  AND2_X1 U8229 ( .A1(n8641), .A2(n8621), .ZN(n8622) );
  NAND2_X1 U8230 ( .A1(n8623), .A2(n8622), .ZN(n8642) );
  INV_X1 U8231 ( .A(n11916), .ZN(n7915) );
  AOI21_X1 U8232 ( .B1(n11916), .B2(n7914), .A(n7545), .ZN(n7913) );
  INV_X1 U8233 ( .A(n11899), .ZN(n7914) );
  NAND2_X1 U8234 ( .A1(n7648), .A2(n7647), .ZN(n12770) );
  INV_X1 U8235 ( .A(n10160), .ZN(n7647) );
  INV_X1 U8236 ( .A(n10159), .ZN(n7648) );
  AOI21_X1 U8237 ( .B1(n10740), .B2(n7907), .A(n7547), .ZN(n7903) );
  INV_X1 U8238 ( .A(n10729), .ZN(n7907) );
  OAI21_X1 U8239 ( .B1(n10042), .B2(n10041), .A(n10040), .ZN(n13983) );
  AND2_X1 U8240 ( .A1(n8149), .A2(n12429), .ZN(n8148) );
  NAND2_X1 U8241 ( .A1(n12368), .A2(n8150), .ZN(n8149) );
  NAND2_X1 U8242 ( .A1(n13940), .A2(n8157), .ZN(n8155) );
  OAI21_X1 U8243 ( .B1(n10986), .B2(n10044), .A(n10047), .ZN(n8295) );
  INV_X1 U8244 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n10217) );
  INV_X1 U8245 ( .A(n7991), .ZN(n14481) );
  INV_X1 U8246 ( .A(n14446), .ZN(n8300) );
  NAND2_X1 U8247 ( .A1(n14513), .A2(n14443), .ZN(n14497) );
  XNOR2_X1 U8248 ( .A(n14760), .B(n7855), .ZN(n14502) );
  NOR2_X2 U8249 ( .A1(n14532), .A2(n14760), .ZN(n14516) );
  NAND2_X1 U8250 ( .A1(n14525), .A2(n8308), .ZN(n14513) );
  NOR2_X1 U8251 ( .A1(n14510), .A2(n8309), .ZN(n8308) );
  INV_X1 U8252 ( .A(n14441), .ZN(n8309) );
  INV_X1 U8253 ( .A(n14502), .ZN(n14510) );
  OR2_X1 U8254 ( .A1(n13803), .A2(n13757), .ZN(n13817) );
  NAND2_X1 U8255 ( .A1(n14541), .A2(n14540), .ZN(n14439) );
  NAND2_X1 U8256 ( .A1(n14439), .A2(n8310), .ZN(n14525) );
  AND2_X1 U8257 ( .A1(n14526), .A2(n14438), .ZN(n8310) );
  NAND2_X1 U8258 ( .A1(n7730), .A2(n14440), .ZN(n14529) );
  NAND2_X1 U8259 ( .A1(n7996), .A2(n7995), .ZN(n14548) );
  AND2_X1 U8260 ( .A1(n14395), .A2(n14396), .ZN(n14574) );
  OAI21_X1 U8261 ( .B1(n14425), .B2(n14424), .A(n14427), .ZN(n14606) );
  OR2_X1 U8262 ( .A1(n14606), .A2(n14610), .ZN(n14608) );
  AND2_X1 U8263 ( .A1(n8171), .A2(n14638), .ZN(n8170) );
  NAND2_X1 U8264 ( .A1(n8172), .A2(n14630), .ZN(n8171) );
  INV_X1 U8265 ( .A(n14270), .ZN(n8172) );
  OR2_X1 U8266 ( .A1(n7723), .A2(n8173), .ZN(n8167) );
  NAND2_X1 U8267 ( .A1(n12210), .A2(n12209), .ZN(n12216) );
  OR2_X1 U8268 ( .A1(n12216), .A2(n14270), .ZN(n12451) );
  NAND2_X1 U8269 ( .A1(n7723), .A2(n14270), .ZN(n14632) );
  NAND2_X1 U8270 ( .A1(n7469), .A2(n14268), .ZN(n12219) );
  AOI21_X1 U8271 ( .B1(n7942), .B2(n11939), .A(n7529), .ZN(n7941) );
  NAND2_X1 U8272 ( .A1(n7936), .A2(n7938), .ZN(n12133) );
  AOI21_X1 U8273 ( .B1(n7941), .B2(n7940), .A(n7939), .ZN(n7938) );
  OR2_X1 U8274 ( .A1(n11940), .A2(n7935), .ZN(n7936) );
  INV_X1 U8275 ( .A(n7942), .ZN(n7940) );
  XNOR2_X1 U8276 ( .A(n14089), .B(n14309), .ZN(n14265) );
  NAND2_X1 U8277 ( .A1(n11676), .A2(n11675), .ZN(n11772) );
  INV_X1 U8278 ( .A(n14310), .ZN(n11938) );
  AOI21_X1 U8279 ( .B1(n8183), .B2(n11500), .A(n7551), .ZN(n8182) );
  NAND2_X1 U8280 ( .A1(n11053), .A2(n14257), .ZN(n8307) );
  NAND2_X1 U8281 ( .A1(n8307), .A2(n8305), .ZN(n11237) );
  NOR2_X1 U8282 ( .A1(n11055), .A2(n8306), .ZN(n8305) );
  INV_X1 U8283 ( .A(n11054), .ZN(n8306) );
  INV_X1 U8284 ( .A(n10821), .ZN(n8179) );
  NOR2_X2 U8285 ( .A1(n10540), .A2(n14026), .ZN(n10837) );
  INV_X1 U8286 ( .A(n10542), .ZN(n14019) );
  NAND2_X1 U8287 ( .A1(n11328), .A2(n10052), .ZN(n10543) );
  INV_X1 U8288 ( .A(n7449), .ZN(n14591) );
  XNOR2_X1 U8289 ( .A(n14319), .B(n10542), .ZN(n14250) );
  OAI22_X1 U8290 ( .A1(n10119), .A2(n14249), .B1(n11656), .B2(n14321), .ZN(
        n11327) );
  XNOR2_X1 U8291 ( .A(n14320), .B(n14005), .ZN(n14247) );
  AND2_X1 U8292 ( .A1(n11958), .A2(n14287), .ZN(n10513) );
  NAND2_X1 U8293 ( .A1(n14204), .A2(n14203), .ZN(n14664) );
  NAND2_X1 U8294 ( .A1(n13756), .A2(n13755), .ZN(n14677) );
  NAND2_X1 U8295 ( .A1(n13815), .A2(n13814), .ZN(n14688) );
  NAND2_X1 U8296 ( .A1(n12511), .A2(n12510), .ZN(n14593) );
  AND2_X1 U8297 ( .A1(n8139), .A2(n14691), .ZN(n14735) );
  OR2_X1 U8298 ( .A1(n10042), .A2(n8493), .ZN(n10031) );
  AND2_X1 U8299 ( .A1(n10513), .A2(n14290), .ZN(n14709) );
  OR2_X1 U8300 ( .A1(n7947), .A2(n7946), .ZN(n7655) );
  NOR2_X1 U8301 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n7653) );
  NOR2_X1 U8302 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n8163) );
  NAND2_X1 U8303 ( .A1(n10013), .A2(n8304), .ZN(n10027) );
  NAND2_X1 U8304 ( .A1(n9956), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9958) );
  NAND2_X1 U8305 ( .A1(n10011), .A2(n9958), .ZN(n9960) );
  NOR2_X1 U8306 ( .A1(n10201), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n10204) );
  NAND2_X1 U8307 ( .A1(n12382), .A2(n8132), .ZN(n8131) );
  NAND2_X1 U8308 ( .A1(n8120), .A2(n7533), .ZN(n7835) );
  NAND2_X1 U8309 ( .A1(n8121), .A2(n12650), .ZN(n8120) );
  NAND2_X1 U8310 ( .A1(n14925), .A2(n14926), .ZN(n7836) );
  INV_X1 U8311 ( .A(n9722), .ZN(n9743) );
  AND2_X1 U8312 ( .A1(n14869), .A2(n8102), .ZN(n8101) );
  OR2_X1 U8313 ( .A1(n14898), .A2(n12677), .ZN(n8102) );
  NAND2_X1 U8314 ( .A1(n14897), .A2(n14898), .ZN(n14896) );
  NAND2_X1 U8315 ( .A1(n7827), .A2(n7825), .ZN(n11722) );
  AND2_X1 U8316 ( .A1(n12640), .A2(n8124), .ZN(n8123) );
  NAND2_X1 U8317 ( .A1(n14851), .A2(n8125), .ZN(n8124) );
  INV_X1 U8318 ( .A(n12631), .ZN(n8125) );
  OAI21_X1 U8319 ( .B1(n14927), .B2(n14926), .A(n14925), .ZN(n14924) );
  NAND2_X1 U8320 ( .A1(n11143), .A2(n11142), .ZN(n8113) );
  NAND2_X1 U8321 ( .A1(n9326), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9295) );
  AND2_X1 U8322 ( .A1(n9292), .A2(n9291), .ZN(n9296) );
  OAI22_X1 U8323 ( .A1(n15050), .A2(n15049), .B1(n15055), .B2(n15048), .ZN(
        n15051) );
  NAND2_X1 U8324 ( .A1(n9798), .A2(n9797), .ZN(n15081) );
  NAND2_X1 U8325 ( .A1(n15089), .A2(n9890), .ZN(n15090) );
  XNOR2_X1 U8326 ( .A(n15094), .B(n14960), .ZN(n15092) );
  INV_X1 U8327 ( .A(n15090), .ZN(n12580) );
  AOI22_X1 U8328 ( .A1(n15131), .A2(n12568), .B1(n15111), .B2(n15382), .ZN(
        n15109) );
  NOR2_X2 U8329 ( .A1(n15382), .A2(n15145), .ZN(n15124) );
  NAND2_X1 U8330 ( .A1(n8463), .A2(n8472), .ZN(n15140) );
  NAND2_X1 U8331 ( .A1(n8437), .A2(n8442), .ZN(n15158) );
  OR2_X1 U8332 ( .A1(n15216), .A2(n8444), .ZN(n8437) );
  NOR2_X1 U8333 ( .A1(n12575), .A2(n8448), .ZN(n8447) );
  INV_X1 U8334 ( .A(n8452), .ZN(n8448) );
  NAND2_X1 U8335 ( .A1(n8453), .A2(n15233), .ZN(n8452) );
  OAI211_X1 U8336 ( .C1(n15921), .C2(n7885), .A(n7523), .B(n7881), .ZN(n15194)
         );
  NAND2_X1 U8337 ( .A1(n15921), .A2(n7882), .ZN(n7881) );
  NOR2_X1 U8338 ( .A1(n14961), .A2(n7883), .ZN(n7882) );
  AND2_X1 U8339 ( .A1(n8340), .A2(n15212), .ZN(n8339) );
  OR2_X1 U8340 ( .A1(n8342), .A2(n8341), .ZN(n8340) );
  NAND2_X1 U8341 ( .A1(n15218), .A2(n15217), .ZN(n15216) );
  NAND2_X1 U8342 ( .A1(n15251), .A2(n8342), .ZN(n15235) );
  OR2_X1 U8343 ( .A1(n15250), .A2(n15248), .ZN(n15251) );
  NOR2_X1 U8344 ( .A1(n7495), .A2(n8483), .ZN(n8480) );
  AND2_X1 U8345 ( .A1(n15440), .A2(n15304), .ZN(n8483) );
  NAND2_X1 U8346 ( .A1(n8431), .A2(n8429), .ZN(n15306) );
  AOI21_X1 U8347 ( .B1(n8432), .B2(n8433), .A(n8430), .ZN(n8429) );
  NAND2_X1 U8348 ( .A1(n12553), .A2(n8326), .ZN(n7889) );
  AOI21_X1 U8349 ( .B1(n12338), .B2(n15462), .A(n12337), .ZN(n12340) );
  NAND2_X1 U8350 ( .A1(n12340), .A2(n12339), .ZN(n12572) );
  NAND2_X1 U8351 ( .A1(n9529), .A2(n9528), .ZN(n12333) );
  NAND2_X1 U8352 ( .A1(n12152), .A2(n12151), .ZN(n8320) );
  NAND2_X1 U8353 ( .A1(n9450), .A2(n9449), .ZN(n11818) );
  INV_X1 U8354 ( .A(n11528), .ZN(n11540) );
  NAND2_X1 U8355 ( .A1(n11529), .A2(n11540), .ZN(n11733) );
  NAND2_X1 U8356 ( .A1(n7878), .A2(n7877), .ZN(n10888) );
  INV_X1 U8357 ( .A(n10862), .ZN(n7877) );
  INV_X1 U8358 ( .A(n15361), .ZN(n15166) );
  INV_X1 U8359 ( .A(n15230), .ZN(n15331) );
  NAND2_X1 U8360 ( .A1(n9660), .A2(n9659), .ZN(n15421) );
  NAND2_X1 U8361 ( .A1(n9577), .A2(n9576), .ZN(n15446) );
  NAND2_X1 U8362 ( .A1(n9564), .A2(n9563), .ZN(n15451) );
  NAND2_X1 U8363 ( .A1(n9503), .A2(n9502), .ZN(n15470) );
  AND2_X1 U8364 ( .A1(n10493), .A2(n10492), .ZN(n16542) );
  NAND2_X1 U8365 ( .A1(n9941), .A2(n9940), .ZN(n10441) );
  AND2_X1 U8366 ( .A1(n12317), .A2(n9982), .ZN(n9941) );
  XNOR2_X1 U8367 ( .A(n9834), .B(n9833), .ZN(n14792) );
  NAND2_X1 U8368 ( .A1(n9824), .A2(n9823), .ZN(n8217) );
  XNOR2_X1 U8369 ( .A(n9782), .B(n9263), .ZN(n14806) );
  NAND2_X1 U8370 ( .A1(n8288), .A2(n8134), .ZN(n9929) );
  XNOR2_X1 U8371 ( .A(n9275), .B(n9926), .ZN(n9998) );
  OR2_X1 U8372 ( .A1(n9927), .A2(n9361), .ZN(n9275) );
  AND2_X1 U8373 ( .A1(n9468), .A2(n9501), .ZN(n10425) );
  NAND2_X1 U8374 ( .A1(n16004), .A2(n16159), .ZN(n7640) );
  AOI21_X1 U8375 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n15946), .A(n15945), .ZN(
        n16012) );
  NOR2_X1 U8376 ( .A1(n15974), .A2(n15973), .ZN(n15945) );
  OAI21_X1 U8377 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n15952), .A(n15951), .ZN(
        n15969) );
  NOR2_X1 U8378 ( .A1(n8366), .A2(n8364), .ZN(n8363) );
  INV_X1 U8379 ( .A(n12322), .ZN(n8364) );
  AND3_X1 U8380 ( .A1(n8911), .A2(n8910), .A3(n8909), .ZN(n13527) );
  AOI21_X1 U8381 ( .B1(n10846), .B2(n12834), .A(n10598), .ZN(n10601) );
  AND2_X1 U8382 ( .A1(n8750), .A2(n8749), .ZN(n12546) );
  AND4_X1 U8383 ( .A1(n8973), .A2(n8972), .A3(n8971), .A4(n8970), .ZN(n13439)
         );
  AND4_X1 U8384 ( .A1(n8875), .A2(n8874), .A3(n8873), .A4(n8872), .ZN(n13548)
         );
  NAND2_X1 U8385 ( .A1(n11468), .A2(n13225), .ZN(n8393) );
  NAND2_X1 U8386 ( .A1(n11083), .A2(n11082), .ZN(n11469) );
  AND2_X1 U8387 ( .A1(n11469), .A2(n8391), .ZN(n11647) );
  AND4_X1 U8388 ( .A1(n8893), .A2(n8892), .A3(n8891), .A4(n8890), .ZN(n13540)
         );
  OR2_X1 U8389 ( .A1(n12810), .A2(n12809), .ZN(n12811) );
  AND4_X1 U8390 ( .A1(n8858), .A2(n8857), .A3(n8856), .A4(n8855), .ZN(n13569)
         );
  OR2_X1 U8391 ( .A1(n11086), .A2(n11085), .ZN(n13202) );
  NOR2_X1 U8392 ( .A1(n11834), .A2(n11833), .ZN(n11992) );
  XNOR2_X1 U8393 ( .A(n12183), .B(n12196), .ZN(n11993) );
  NOR2_X1 U8394 ( .A1(n12184), .A2(n12188), .ZN(n12293) );
  NOR2_X1 U8395 ( .A1(n12284), .A2(n12283), .ZN(n13246) );
  NOR2_X1 U8396 ( .A1(n13258), .A2(n13651), .ZN(n13277) );
  XNOR2_X1 U8397 ( .A(n8257), .B(n13365), .ZN(n8256) );
  NAND2_X1 U8398 ( .A1(n8259), .A2(n8258), .ZN(n8257) );
  NAND2_X1 U8399 ( .A1(n13364), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8258) );
  NAND2_X1 U8400 ( .A1(n13366), .A2(n13367), .ZN(n8255) );
  AOI21_X1 U8401 ( .B1(P3_REG1_REG_18__SCAN_IN), .B2(n13364), .A(n13350), .ZN(
        n13351) );
  NAND2_X1 U8402 ( .A1(n8852), .A2(n8851), .ZN(n13644) );
  AND3_X1 U8403 ( .A1(n8661), .A2(n8660), .A3(n8659), .ZN(n11924) );
  AND3_X1 U8404 ( .A1(n8591), .A2(n8590), .A3(n8589), .ZN(n16422) );
  OR2_X1 U8405 ( .A1(n8616), .A2(SI_3_), .ZN(n8591) );
  NOR2_X1 U8406 ( .A1(n8519), .A2(n9066), .ZN(n8089) );
  NOR2_X1 U8407 ( .A1(n13380), .A2(n13657), .ZN(n9135) );
  OAI22_X1 U8408 ( .A1(n13673), .A2(n13657), .B1(n16565), .B2(n13597), .ZN(
        n7811) );
  INV_X1 U8409 ( .A(n13040), .ZN(n9050) );
  NOR2_X1 U8410 ( .A1(n16569), .A2(n9146), .ZN(n8091) );
  INV_X1 U8411 ( .A(n8089), .ZN(n8088) );
  INV_X1 U8412 ( .A(n12978), .ZN(n13673) );
  NOR2_X1 U8413 ( .A1(n7498), .A2(n7807), .ZN(n7806) );
  INV_X1 U8414 ( .A(n13394), .ZN(n7807) );
  NAND2_X1 U8415 ( .A1(n8917), .A2(n8916), .ZN(n13702) );
  NAND2_X1 U8416 ( .A1(n16569), .A2(n16471), .ZN(n13731) );
  OAI21_X1 U8417 ( .B1(n8415), .B2(n8252), .A(n8251), .ZN(n8250) );
  INV_X1 U8418 ( .A(n8554), .ZN(n8555) );
  NAND2_X1 U8419 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n8252) );
  INV_X1 U8420 ( .A(n8154), .ZN(n8153) );
  AOI21_X1 U8421 ( .B1(n8158), .B2(n8154), .A(n8160), .ZN(n8152) );
  NAND2_X1 U8422 ( .A1(n12503), .A2(n12502), .ZN(n14621) );
  NAND2_X1 U8423 ( .A1(n7922), .A2(n7923), .ZN(n12753) );
  NAND2_X1 U8424 ( .A1(n12356), .A2(n12355), .ZN(n14728) );
  AND2_X1 U8425 ( .A1(n13887), .A2(n12504), .ZN(n7646) );
  NOR2_X1 U8426 ( .A1(n14285), .A2(n14294), .ZN(n8207) );
  NAND2_X1 U8427 ( .A1(n13849), .A2(n13848), .ZN(n14447) );
  NAND2_X1 U8428 ( .A1(n14189), .A2(n14188), .ZN(n14382) );
  OR2_X1 U8429 ( .A1(n14186), .A2(n14185), .ZN(n14189) );
  XNOR2_X1 U8430 ( .A(n7927), .B(n8313), .ZN(n14667) );
  NAND2_X1 U8431 ( .A1(n14457), .A2(n14448), .ZN(n7927) );
  NAND2_X1 U8432 ( .A1(n14644), .A2(n10129), .ZN(n14604) );
  NAND2_X1 U8433 ( .A1(n16076), .A2(n10117), .ZN(n14641) );
  OAI21_X1 U8434 ( .B1(n10904), .B2(n8109), .A(n8107), .ZN(n11665) );
  INV_X1 U8435 ( .A(n8108), .ZN(n8107) );
  NAND2_X1 U8436 ( .A1(n8114), .A2(n8110), .ZN(n8109) );
  OAI22_X1 U8437 ( .A1(n8113), .A2(n11457), .B1(n11455), .B2(n11456), .ZN(
        n8108) );
  AND2_X1 U8438 ( .A1(n7586), .A2(n8118), .ZN(n8116) );
  INV_X1 U8439 ( .A(n8119), .ZN(n8118) );
  OAI21_X1 U8440 ( .B1(n12710), .B2(n12704), .A(n14947), .ZN(n8119) );
  INV_X1 U8441 ( .A(n14963), .ZN(n12312) );
  AND2_X1 U8442 ( .A1(n7631), .A2(n9886), .ZN(n7630) );
  NAND2_X1 U8443 ( .A1(n12551), .A2(n7528), .ZN(n9308) );
  OR2_X1 U8444 ( .A1(n9724), .A2(n10458), .ZN(n9305) );
  OR2_X1 U8445 ( .A1(n9724), .A2(n10503), .ZN(n9279) );
  NAND2_X1 U8446 ( .A1(n10306), .A2(n10305), .ZN(n14996) );
  AND2_X1 U8447 ( .A1(n9856), .A2(n9855), .ZN(n12707) );
  OAI21_X1 U8448 ( .B1(n8463), .B2(n8467), .A(n7541), .ZN(n15108) );
  NAND2_X1 U8449 ( .A1(n8469), .A2(n15143), .ZN(n8462) );
  AND2_X1 U8450 ( .A1(n7895), .A2(n7893), .ZN(n15381) );
  NAND2_X1 U8451 ( .A1(n7894), .A2(n15431), .ZN(n7893) );
  AOI21_X1 U8452 ( .B1(n15379), .B2(n15166), .A(n15113), .ZN(n7895) );
  XNOR2_X1 U8453 ( .A(n15109), .B(n15110), .ZN(n7894) );
  NOR2_X1 U8454 ( .A1(n12155), .A2(n8461), .ZN(n12158) );
  OAI21_X1 U8455 ( .B1(n11862), .B2(n8461), .A(n8457), .ZN(n8460) );
  OR2_X1 U8456 ( .A1(n9351), .A2(n10229), .ZN(n9313) );
  NAND2_X1 U8457 ( .A1(n7883), .A2(n10461), .ZN(n9314) );
  NAND2_X1 U8458 ( .A1(n10495), .A2(n9999), .ZN(n15312) );
  NOR3_X1 U8459 ( .A1(n8317), .A2(n9156), .A3(n7542), .ZN(n7890) );
  NAND2_X1 U8460 ( .A1(n9936), .A2(n7642), .ZN(n7702) );
  NOR2_X1 U8461 ( .A1(n7703), .A2(n9361), .ZN(n7642) );
  NAND2_X1 U8462 ( .A1(n14003), .A2(n14002), .ZN(n14011) );
  INV_X1 U8463 ( .A(n14022), .ZN(n7651) );
  INV_X1 U8464 ( .A(n14021), .ZN(n7650) );
  INV_X1 U8465 ( .A(n7587), .ZN(n8504) );
  NAND2_X1 U8466 ( .A1(n8260), .A2(n8261), .ZN(n9432) );
  NAND2_X1 U8467 ( .A1(n9414), .A2(n9416), .ZN(n8261) );
  NAND2_X1 U8468 ( .A1(n9451), .A2(n8275), .ZN(n8274) );
  NAND2_X1 U8469 ( .A1(n7682), .A2(n7681), .ZN(n7625) );
  INV_X1 U8470 ( .A(n14039), .ZN(n7681) );
  NAND2_X1 U8471 ( .A1(n9491), .A2(n9493), .ZN(n8265) );
  NOR2_X1 U8472 ( .A1(n14063), .A2(n14065), .ZN(n8500) );
  NAND2_X1 U8473 ( .A1(n8281), .A2(n9530), .ZN(n8280) );
  INV_X1 U8474 ( .A(n14069), .ZN(n7677) );
  NAND2_X1 U8475 ( .A1(n9565), .A2(n9567), .ZN(n8267) );
  NAND2_X1 U8476 ( .A1(n8486), .A2(n8485), .ZN(n8484) );
  INV_X1 U8477 ( .A(n14085), .ZN(n8485) );
  NAND2_X1 U8478 ( .A1(n9602), .A2(n9604), .ZN(n8263) );
  NAND2_X1 U8479 ( .A1(n9647), .A2(n8278), .ZN(n8277) );
  INV_X1 U8480 ( .A(n14104), .ZN(n7635) );
  OAI21_X1 U8481 ( .B1(n14137), .B2(n7649), .A(n7555), .ZN(n14147) );
  NAND2_X1 U8482 ( .A1(n9721), .A2(n9720), .ZN(n9736) );
  AND2_X1 U8483 ( .A1(n8271), .A2(n9719), .ZN(n7750) );
  NAND2_X1 U8484 ( .A1(n14161), .A2(n7962), .ZN(n7961) );
  INV_X1 U8485 ( .A(n7965), .ZN(n7962) );
  NAND2_X1 U8486 ( .A1(n8284), .A2(n9753), .ZN(n8283) );
  NOR2_X1 U8487 ( .A1(n9712), .A2(n8206), .ZN(n8204) );
  INV_X1 U8488 ( .A(n11956), .ZN(n8206) );
  INV_X1 U8489 ( .A(SI_17_), .ZN(n15717) );
  AND2_X1 U8490 ( .A1(n8223), .A2(n9557), .ZN(n8222) );
  NAND2_X1 U8491 ( .A1(n9539), .A2(n9220), .ZN(n8223) );
  INV_X1 U8492 ( .A(SI_15_), .ZN(n15521) );
  NAND2_X1 U8493 ( .A1(n8074), .A2(n8073), .ZN(n12970) );
  NAND2_X1 U8494 ( .A1(n8489), .A2(n7512), .ZN(n8488) );
  INV_X1 U8495 ( .A(n14178), .ZN(n8490) );
  NAND2_X1 U8496 ( .A1(n9811), .A2(n9841), .ZN(n8290) );
  NAND2_X1 U8497 ( .A1(n10443), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n7819) );
  INV_X1 U8498 ( .A(n8442), .ZN(n8440) );
  AND2_X1 U8499 ( .A1(n9763), .A2(n9260), .ZN(n8233) );
  NAND2_X1 U8500 ( .A1(n7844), .A2(n7843), .ZN(n9254) );
  INV_X1 U8501 ( .A(n8203), .ZN(n7843) );
  NAND2_X1 U8502 ( .A1(n9248), .A2(n8204), .ZN(n7844) );
  OAI21_X1 U8503 ( .B1(n9250), .B2(n9712), .A(n9252), .ZN(n8203) );
  NAND2_X1 U8504 ( .A1(n7676), .A2(n7517), .ZN(n9240) );
  NAND2_X1 U8505 ( .A1(n9228), .A2(n7850), .ZN(n7676) );
  INV_X1 U8506 ( .A(n7863), .ZN(n7861) );
  INV_X1 U8507 ( .A(n8222), .ZN(n8221) );
  INV_X1 U8508 ( .A(n8218), .ZN(n7858) );
  AOI21_X1 U8509 ( .B1(n8222), .B2(n8220), .A(n8219), .ZN(n8218) );
  INV_X1 U8510 ( .A(n9220), .ZN(n8220) );
  INV_X1 U8511 ( .A(n9224), .ZN(n8219) );
  INV_X1 U8512 ( .A(n8201), .ZN(n8200) );
  OAI21_X1 U8513 ( .B1(n9198), .B2(n8202), .A(n9201), .ZN(n8201) );
  INV_X1 U8514 ( .A(n9200), .ZN(n8202) );
  OAI21_X1 U8515 ( .B1(n10196), .B2(n10179), .A(n7854), .ZN(n9181) );
  NAND2_X1 U8516 ( .A1(n10029), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7724) );
  OAI21_X1 U8517 ( .B1(P3_ADDR_REG_15__SCAN_IN), .B2(n15958), .A(n15957), .ZN(
        n15959) );
  OR2_X1 U8518 ( .A1(n13702), .A2(n13514), .ZN(n12852) );
  AOI21_X1 U8519 ( .B1(n8391), .B2(n8389), .A(n11646), .ZN(n8388) );
  INV_X1 U8520 ( .A(n11082), .ZN(n8389) );
  INV_X1 U8521 ( .A(n8391), .ZN(n8390) );
  NOR2_X1 U8522 ( .A1(n13049), .A2(n13050), .ZN(n8421) );
  NAND2_X1 U8523 ( .A1(n13052), .A2(n13051), .ZN(n8422) );
  NOR4_X1 U8524 ( .A1(n13390), .A2(n9080), .A3(n13452), .A4(n13038), .ZN(
        n13041) );
  NAND2_X1 U8525 ( .A1(n13009), .A2(n13008), .ZN(n13043) );
  NOR2_X1 U8526 ( .A1(n13315), .A2(n7605), .ZN(n13327) );
  NOR2_X1 U8527 ( .A1(n13335), .A2(n13336), .ZN(n13352) );
  AND2_X1 U8528 ( .A1(n8525), .A2(n8829), .ZN(n7790) );
  INV_X1 U8529 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8525) );
  OR2_X1 U8530 ( .A1(n9013), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9031) );
  NOR2_X1 U8531 ( .A1(n8399), .A2(n8396), .ZN(n8395) );
  INV_X1 U8532 ( .A(n13023), .ZN(n8396) );
  INV_X1 U8533 ( .A(n9069), .ZN(n8398) );
  NAND2_X1 U8534 ( .A1(n7558), .A2(n8083), .ZN(n8082) );
  AND2_X1 U8535 ( .A1(n12852), .A2(n12853), .ZN(n13494) );
  NAND2_X1 U8536 ( .A1(n8345), .A2(n7515), .ZN(n13511) );
  INV_X1 U8537 ( .A(n9075), .ZN(n8404) );
  AOI21_X1 U8538 ( .B1(n9075), .B2(n8403), .A(n8402), .ZN(n8401) );
  AND2_X1 U8539 ( .A1(n13027), .A2(n12396), .ZN(n9075) );
  AOI21_X1 U8540 ( .B1(n8061), .B2(n8063), .A(n8060), .ZN(n8059) );
  INV_X1 U8541 ( .A(n8761), .ZN(n8060) );
  NOR2_X1 U8542 ( .A1(n8712), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n8732) );
  INV_X1 U8543 ( .A(n8040), .ZN(n8039) );
  OAI21_X1 U8544 ( .B1(n8622), .B2(n8041), .A(n8655), .ZN(n8040) );
  INV_X1 U8545 ( .A(n12353), .ZN(n8150) );
  INV_X1 U8546 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10578) );
  OR2_X1 U8547 ( .A1(n10579), .A2(n10578), .ZN(n10734) );
  INV_X1 U8548 ( .A(n7941), .ZN(n7935) );
  NAND2_X1 U8549 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), 
        .ZN(n7946) );
  INV_X1 U8550 ( .A(n10016), .ZN(n7654) );
  INV_X1 U8551 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9949) );
  OR2_X1 U8552 ( .A1(n10238), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n10245) );
  INV_X1 U8553 ( .A(n9952), .ZN(n10067) );
  INV_X1 U8554 ( .A(n8123), .ZN(n8121) );
  NOR2_X1 U8555 ( .A1(n7826), .A2(n8103), .ZN(n7824) );
  NAND2_X1 U8556 ( .A1(n11968), .A2(n7466), .ZN(n8103) );
  INV_X1 U8557 ( .A(n11664), .ZN(n7822) );
  NAND2_X1 U8558 ( .A1(n7560), .A2(n7466), .ZN(n7828) );
  OR2_X1 U8559 ( .A1(n8105), .A2(n11967), .ZN(n8104) );
  AOI21_X1 U8560 ( .B1(n8445), .B2(n8443), .A(n8449), .ZN(n8442) );
  NOR2_X1 U8561 ( .A1(n15183), .A2(n15198), .ZN(n8449) );
  INV_X1 U8562 ( .A(n8447), .ZN(n8443) );
  INV_X1 U8563 ( .A(n12562), .ZN(n8341) );
  INV_X1 U8564 ( .A(n15327), .ZN(n8329) );
  NOR2_X1 U8565 ( .A1(n15456), .A2(n15451), .ZN(n8010) );
  INV_X1 U8566 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9532) );
  NOR2_X1 U8567 ( .A1(n9533), .A2(n9532), .ZN(n9553) );
  NAND2_X1 U8568 ( .A1(n12311), .A2(n12312), .ZN(n8459) );
  INV_X1 U8569 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9479) );
  NOR2_X1 U8570 ( .A1(n9480), .A2(n9479), .ZN(n9494) );
  INV_X1 U8571 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9436) );
  AND2_X1 U8572 ( .A1(n11528), .A2(n11538), .ZN(n8334) );
  NOR2_X1 U8573 ( .A1(n11531), .A2(n16478), .ZN(n8005) );
  OR2_X1 U8574 ( .A1(n9332), .A2(n15342), .ZN(n10847) );
  NOR2_X1 U8575 ( .A1(n15194), .A2(n7880), .ZN(n7879) );
  NOR2_X1 U8576 ( .A1(n8000), .A2(n16446), .ZN(n11159) );
  INV_X1 U8577 ( .A(n15915), .ZN(n9982) );
  AOI21_X1 U8578 ( .B1(n8213), .B2(n8214), .A(n8212), .ZN(n8211) );
  INV_X1 U8579 ( .A(n9830), .ZN(n8212) );
  INV_X1 U8580 ( .A(n9823), .ZN(n8213) );
  INV_X1 U8581 ( .A(n9794), .ZN(n8216) );
  AND2_X1 U8582 ( .A1(n7481), .A2(n9926), .ZN(n8134) );
  INV_X1 U8583 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n15684) );
  NAND2_X1 U8584 ( .A1(n9217), .A2(n15525), .ZN(n9220) );
  NAND2_X1 U8585 ( .A1(n7862), .A2(n7863), .ZN(n9540) );
  NAND2_X1 U8586 ( .A1(n9487), .A2(n7865), .ZN(n7862) );
  NAND2_X1 U8587 ( .A1(n7841), .A2(n9193), .ZN(n9409) );
  NAND2_X1 U8588 ( .A1(n10029), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7731) );
  NAND2_X1 U8589 ( .A1(n15924), .A2(n7984), .ZN(n15925) );
  NAND2_X1 U8590 ( .A1(n7985), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7984) );
  NAND2_X1 U8591 ( .A1(n15984), .A2(n15982), .ZN(n15924) );
  INV_X1 U8592 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7985) );
  INV_X1 U8593 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7981) );
  INV_X1 U8594 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n11267) );
  NAND2_X2 U8595 ( .A1(n10597), .A2(n10596), .ZN(n12834) );
  AND2_X1 U8596 ( .A1(n8834), .A2(n15773), .ZN(n8853) );
  INV_X1 U8597 ( .A(n8968), .ZN(n8967) );
  AND2_X1 U8598 ( .A1(n8369), .A2(n8372), .ZN(n8368) );
  INV_X1 U8599 ( .A(n12123), .ZN(n8369) );
  OR2_X1 U8600 ( .A1(n12119), .A2(n12124), .ZN(n8372) );
  NAND2_X1 U8601 ( .A1(n8371), .A2(n8373), .ZN(n8370) );
  INV_X1 U8602 ( .A(n12121), .ZN(n8371) );
  NAND2_X1 U8603 ( .A1(n8772), .A2(n8771), .ZN(n8796) );
  NAND2_X1 U8604 ( .A1(n12812), .A2(n13100), .ZN(n13162) );
  OR2_X1 U8605 ( .A1(n8700), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8719) );
  OR2_X1 U8606 ( .A1(n8719), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8753) );
  NAND2_X1 U8607 ( .A1(n8631), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8577) );
  AND2_X1 U8608 ( .A1(n10619), .A2(n10618), .ZN(n13185) );
  OR2_X1 U8609 ( .A1(n8983), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9011) );
  NOR2_X1 U8610 ( .A1(n8813), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8834) );
  INV_X1 U8611 ( .A(n13043), .ZN(n13042) );
  AND4_X1 U8612 ( .A1(n8705), .A2(n8704), .A3(n8703), .A4(n8702), .ZN(n12416)
         );
  AND4_X1 U8613 ( .A1(n8567), .A2(n8566), .A3(n8565), .A4(n8564), .ZN(n16375)
         );
  NAND2_X1 U8614 ( .A1(n8631), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U8615 ( .A1(n7753), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n11215) );
  MUX2_X1 U8616 ( .A(P3_REG2_REG_2__SCAN_IN), .B(n16413), .S(n8249), .Z(n10942) );
  NAND2_X1 U8617 ( .A1(n11215), .A2(n10931), .ZN(n10932) );
  OAI21_X1 U8618 ( .B1(n8249), .B2(n10928), .A(n8013), .ZN(n10933) );
  NAND2_X1 U8619 ( .A1(n10933), .A2(n10932), .ZN(n10957) );
  NAND2_X1 U8620 ( .A1(n10959), .A2(n11289), .ZN(n10961) );
  NAND2_X1 U8621 ( .A1(n8026), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n11291) );
  INV_X1 U8622 ( .A(n11015), .ZN(n11296) );
  OR2_X1 U8623 ( .A1(n11012), .A2(n11017), .ZN(n7763) );
  OR2_X1 U8624 ( .A1(n11014), .A2(n11523), .ZN(n11403) );
  NAND2_X1 U8625 ( .A1(n11270), .A2(n11271), .ZN(n11433) );
  NAND2_X1 U8626 ( .A1(n11434), .A2(n7754), .ZN(n11435) );
  NAND2_X1 U8627 ( .A1(n7755), .A2(n11439), .ZN(n7754) );
  INV_X1 U8628 ( .A(n7756), .ZN(n7755) );
  INV_X1 U8629 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n15946) );
  NAND2_X1 U8630 ( .A1(n7756), .A2(n11839), .ZN(n11434) );
  NOR2_X1 U8631 ( .A1(n11435), .A2(n16503), .ZN(n11831) );
  NAND2_X1 U8632 ( .A1(n8253), .A2(n7768), .ZN(n7765) );
  NAND2_X1 U8633 ( .A1(n7767), .A2(n7606), .ZN(n7766) );
  AND2_X1 U8634 ( .A1(n12294), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8248) );
  AND2_X1 U8635 ( .A1(n12288), .A2(n12287), .ZN(n12290) );
  XNOR2_X1 U8636 ( .A(n13282), .B(n7871), .ZN(n13263) );
  XNOR2_X1 U8637 ( .A(n13352), .B(n13364), .ZN(n13339) );
  NAND2_X1 U8638 ( .A1(n13339), .A2(n13338), .ZN(n13355) );
  NAND2_X1 U8639 ( .A1(n7786), .A2(n7787), .ZN(n8866) );
  AND4_X1 U8640 ( .A1(n7792), .A2(n7791), .A3(n7790), .A4(n8526), .ZN(n7786)
         );
  NAND2_X1 U8641 ( .A1(n13386), .A2(n12977), .ZN(n13052) );
  NAND2_X1 U8642 ( .A1(n13388), .A2(n13387), .ZN(n13386) );
  NAND2_X1 U8643 ( .A1(n13435), .A2(n8990), .ZN(n13420) );
  NAND2_X1 U8644 ( .A1(n13465), .A2(n9080), .ZN(n13464) );
  AND2_X1 U8645 ( .A1(n8094), .A2(n7795), .ZN(n7794) );
  NAND2_X1 U8646 ( .A1(n15761), .A2(n8918), .ZN(n8939) );
  AOI21_X1 U8647 ( .B1(n8409), .B2(n8407), .A(n7475), .ZN(n8406) );
  INV_X1 U8648 ( .A(n8409), .ZN(n8408) );
  AND2_X1 U8649 ( .A1(n12926), .A2(n12927), .ZN(n13034) );
  OR2_X1 U8650 ( .A1(n9072), .A2(n9071), .ZN(n12246) );
  NAND2_X1 U8651 ( .A1(n8093), .A2(n8699), .ZN(n12072) );
  AND2_X1 U8652 ( .A1(n13024), .A2(n8699), .ZN(n8092) );
  NAND2_X1 U8653 ( .A1(n11977), .A2(n12895), .ZN(n12245) );
  NAND2_X1 U8654 ( .A1(n8682), .A2(n15782), .ZN(n8700) );
  INV_X1 U8655 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n15782) );
  AND2_X1 U8656 ( .A1(n8663), .A2(n11267), .ZN(n8682) );
  NAND2_X1 U8657 ( .A1(n11979), .A2(n8681), .ZN(n12034) );
  AND2_X1 U8658 ( .A1(n12899), .A2(n12900), .ZN(n13014) );
  NOR2_X1 U8659 ( .A1(n8649), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8663) );
  OR2_X1 U8660 ( .A1(n8629), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8649) );
  NAND2_X1 U8661 ( .A1(n8356), .A2(n8359), .ZN(n11512) );
  AOI21_X1 U8662 ( .B1(n13016), .B2(n8361), .A(n8360), .ZN(n8359) );
  INV_X1 U8663 ( .A(n12877), .ZN(n8360) );
  AND4_X1 U8664 ( .A1(n8545), .A2(n8544), .A3(n8543), .A4(n8542), .ZN(n16373)
         );
  OR2_X1 U8665 ( .A1(n16375), .A2(n10846), .ZN(n16371) );
  NAND2_X1 U8666 ( .A1(n10689), .A2(n10688), .ZN(n10690) );
  NAND2_X1 U8667 ( .A1(n12999), .A2(n12998), .ZN(n13054) );
  NAND2_X1 U8668 ( .A1(n8982), .A2(n8981), .ZN(n13104) );
  AND4_X1 U8669 ( .A1(n8988), .A2(n8987), .A3(n8986), .A4(n8985), .ZN(n13453)
         );
  NAND2_X1 U8670 ( .A1(n13516), .A2(n8912), .ZN(n13497) );
  OAI21_X1 U8671 ( .B1(n16367), .B2(n16370), .A(n12857), .ZN(n11130) );
  NAND2_X1 U8672 ( .A1(n13017), .A2(n11130), .ZN(n12863) );
  AND2_X1 U8673 ( .A1(n12865), .A2(n12867), .ZN(n13017) );
  NAND2_X1 U8674 ( .A1(n9090), .A2(n9124), .ZN(n13661) );
  NAND2_X1 U8675 ( .A1(n12985), .A2(n12984), .ZN(n12991) );
  NAND2_X1 U8676 ( .A1(n9005), .A2(n9004), .ZN(n9021) );
  XNOR2_X1 U8677 ( .A(n9094), .B(n9093), .ZN(n9105) );
  NAND2_X1 U8678 ( .A1(n9095), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9094) );
  INV_X1 U8679 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8031) );
  XNOR2_X1 U8680 ( .A(n9121), .B(n9120), .ZN(n10925) );
  NAND2_X1 U8681 ( .A1(n8913), .A2(n7623), .ZN(n7622) );
  AOI21_X1 U8682 ( .B1(n8823), .B2(n8044), .A(n8043), .ZN(n8042) );
  INV_X1 U8683 ( .A(n8823), .ZN(n8045) );
  INV_X1 U8684 ( .A(n8842), .ZN(n8043) );
  AND2_X1 U8685 ( .A1(n8860), .A2(n8844), .ZN(n8845) );
  AND2_X1 U8686 ( .A1(n8788), .A2(n8787), .ZN(n8792) );
  NAND2_X1 U8687 ( .A1(n8782), .A2(n8781), .ZN(n8785) );
  NOR2_X1 U8688 ( .A1(n8767), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n8788) );
  OR2_X1 U8689 ( .A1(n8746), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n8767) );
  AOI21_X1 U8690 ( .B1(n8049), .B2(n8051), .A(n8048), .ZN(n8047) );
  INV_X1 U8691 ( .A(n8706), .ZN(n8048) );
  OR2_X1 U8692 ( .A1(n8688), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8712) );
  OR2_X1 U8693 ( .A1(n8639), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8688) );
  AND2_X1 U8694 ( .A1(n8674), .A2(n8657), .ZN(n8671) );
  AND2_X1 U8695 ( .A1(n8619), .A2(n8601), .ZN(n8617) );
  INV_X1 U8696 ( .A(n8418), .ZN(n8417) );
  AND2_X1 U8697 ( .A1(n8599), .A2(n8584), .ZN(n8585) );
  NAND2_X1 U8698 ( .A1(n8638), .A2(n8523), .ZN(n8251) );
  AND2_X1 U8699 ( .A1(n8549), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8568) );
  AND2_X1 U8700 ( .A1(n13842), .A2(n13841), .ZN(n8160) );
  OR2_X1 U8701 ( .A1(n11785), .A2(n11784), .ZN(n11905) );
  NAND2_X1 U8702 ( .A1(n11606), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n11785) );
  INV_X1 U8703 ( .A(n11608), .ZN(n11606) );
  OR2_X1 U8704 ( .A1(n12104), .A2(n7502), .ZN(n7925) );
  INV_X1 U8705 ( .A(n12513), .ZN(n12512) );
  AND2_X1 U8706 ( .A1(n11617), .A2(n8143), .ZN(n8142) );
  OR2_X1 U8707 ( .A1(n11345), .A2(n7470), .ZN(n8143) );
  NAND2_X1 U8708 ( .A1(n10987), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n11355) );
  OR2_X1 U8709 ( .A1(n11355), .A2(n11354), .ZN(n11608) );
  INV_X1 U8710 ( .A(n12223), .ZN(n12221) );
  AND2_X1 U8711 ( .A1(n8156), .A2(n7569), .ZN(n8154) );
  NAND2_X1 U8712 ( .A1(n8161), .A2(n13825), .ZN(n8156) );
  OR2_X1 U8713 ( .A1(n11905), .A2(n11904), .ZN(n12020) );
  AND2_X1 U8714 ( .A1(n8210), .A2(n14237), .ZN(n8209) );
  NAND2_X1 U8715 ( .A1(n14225), .A2(n7527), .ZN(n8210) );
  INV_X1 U8716 ( .A(n10059), .ZN(n13843) );
  OR2_X1 U8717 ( .A1(n10057), .A2(n10034), .ZN(n10037) );
  OR2_X1 U8718 ( .A1(n10059), .A2(n10878), .ZN(n10035) );
  NAND2_X1 U8719 ( .A1(n10270), .A2(n8296), .ZN(n10271) );
  NOR2_X1 U8720 ( .A1(n16151), .A2(n7694), .ZN(n14326) );
  AND2_X1 U8721 ( .A1(n16156), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7694) );
  OR2_X1 U8722 ( .A1(n10234), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n10238) );
  NOR2_X1 U8723 ( .A1(n16166), .A2(n16165), .ZN(n16164) );
  NOR2_X1 U8724 ( .A1(n16164), .A2(n7695), .ZN(n16243) );
  AND2_X1 U8725 ( .A1(n16169), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7695) );
  NOR2_X1 U8726 ( .A1(n10245), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n10252) );
  NOR2_X1 U8727 ( .A1(n16176), .A2(n7696), .ZN(n11196) );
  AND2_X1 U8728 ( .A1(n16181), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7696) );
  NOR2_X1 U8729 ( .A1(n14348), .A2(n14347), .ZN(n16204) );
  NOR2_X1 U8730 ( .A1(n16204), .A2(n16203), .ZN(n16202) );
  AOI21_X1 U8731 ( .B1(n16207), .B2(P2_REG1_REG_16__SCAN_IN), .A(n16202), .ZN(
        n16212) );
  AOI21_X1 U8732 ( .B1(n16218), .B2(P2_REG1_REG_17__SCAN_IN), .A(n16210), .ZN(
        n14355) );
  NAND2_X1 U8733 ( .A1(n7990), .A2(n14412), .ZN(n7846) );
  NAND2_X1 U8734 ( .A1(n14459), .A2(n14458), .ZN(n14457) );
  NAND2_X1 U8735 ( .A1(n14529), .A2(n14405), .ZN(n14503) );
  NAND2_X1 U8736 ( .A1(n13758), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n13827) );
  OR2_X1 U8737 ( .A1(n12357), .A2(n12445), .ZN(n12439) );
  AOI21_X1 U8738 ( .B1(n7932), .B2(n7931), .A(n7508), .ZN(n7930) );
  OR2_X1 U8739 ( .A1(n12216), .A2(n7933), .ZN(n7929) );
  INV_X1 U8740 ( .A(n12450), .ZN(n7931) );
  AOI21_X1 U8741 ( .B1(n8170), .B2(n8173), .A(n7537), .ZN(n8168) );
  INV_X1 U8742 ( .A(n7993), .ZN(n14648) );
  OR2_X1 U8743 ( .A1(n12096), .A2(n12741), .ZN(n12223) );
  NAND2_X1 U8744 ( .A1(n12018), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n12096) );
  INV_X1 U8745 ( .A(n12020), .ZN(n12018) );
  NAND2_X1 U8746 ( .A1(n7740), .A2(n7739), .ZN(n12142) );
  AOI21_X1 U8747 ( .B1(n8176), .B2(n8178), .A(n7477), .ZN(n8175) );
  OAI21_X1 U8748 ( .B1(n7721), .B2(n8178), .A(n8176), .ZN(n12013) );
  NAND2_X1 U8749 ( .A1(n11796), .A2(n16572), .ZN(n11949) );
  AND2_X1 U8750 ( .A1(n11943), .A2(n11778), .ZN(n14264) );
  CLKBUF_X1 U8751 ( .A(n11782), .Z(n7721) );
  NAND2_X1 U8752 ( .A1(n7721), .A2(n14264), .ZN(n11944) );
  NAND2_X1 U8753 ( .A1(n11499), .A2(n11498), .ZN(n11674) );
  NAND2_X1 U8754 ( .A1(n7989), .A2(n7988), .ZN(n11683) );
  NAND2_X1 U8755 ( .A1(n8185), .A2(n11502), .ZN(n11678) );
  OR2_X1 U8756 ( .A1(n11501), .A2(n11500), .ZN(n8185) );
  NAND2_X1 U8757 ( .A1(n11237), .A2(n11236), .ZN(n11238) );
  NAND2_X1 U8758 ( .A1(n11238), .A2(n14259), .ZN(n11499) );
  NOR2_X2 U8759 ( .A1(n10828), .A2(n14044), .ZN(n11062) );
  NAND2_X1 U8760 ( .A1(n10801), .A2(n10800), .ZN(n10833) );
  INV_X1 U8761 ( .A(n14374), .ZN(n14614) );
  AND2_X2 U8762 ( .A1(n10043), .A2(n10033), .ZN(n14249) );
  OR2_X1 U8763 ( .A1(n7458), .A2(n14366), .ZN(n10505) );
  NAND2_X1 U8764 ( .A1(n13789), .A2(n13788), .ZN(n14564) );
  AND2_X1 U8765 ( .A1(n10143), .A2(n16082), .ZN(n16076) );
  OR2_X1 U8766 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n10015) );
  NAND2_X1 U8767 ( .A1(n10016), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10014) );
  OAI21_X1 U8768 ( .B1(n9963), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9961) );
  INV_X1 U8769 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n9955) );
  XNOR2_X1 U8770 ( .A(n10401), .B(P2_IR_REG_14__SCAN_IN), .ZN(n12276) );
  AND2_X1 U8771 ( .A1(n10339), .A2(n10468), .ZN(n12275) );
  AND2_X1 U8772 ( .A1(n10204), .A2(n10203), .ZN(n10218) );
  INV_X1 U8773 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9400) );
  NOR2_X1 U8774 ( .A1(n9401), .A2(n9400), .ZN(n9417) );
  NOR2_X1 U8775 ( .A1(n8112), .A2(n11457), .ZN(n8110) );
  NAND2_X1 U8776 ( .A1(n14924), .A2(n12631), .ZN(n14850) );
  NOR2_X1 U8777 ( .A1(n9606), .A2(n9605), .ZN(n9626) );
  AND2_X1 U8778 ( .A1(n10487), .A2(n7593), .ZN(n10488) );
  INV_X1 U8779 ( .A(n9703), .ZN(n9723) );
  NAND2_X1 U8780 ( .A1(n9723), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9722) );
  NAND2_X1 U8781 ( .A1(n14850), .A2(n14851), .ZN(n14906) );
  NAND2_X1 U8782 ( .A1(n9494), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9514) );
  NOR2_X1 U8783 ( .A1(n7835), .A2(n8514), .ZN(n7833) );
  NOR2_X1 U8784 ( .A1(n8122), .A2(n7838), .ZN(n7837) );
  INV_X1 U8785 ( .A(n14925), .ZN(n7838) );
  OAI21_X1 U8786 ( .B1(n11665), .B2(n7823), .A(n7820), .ZN(n12062) );
  INV_X1 U8787 ( .A(n7824), .ZN(n7823) );
  AND2_X1 U8788 ( .A1(n7828), .A2(n7821), .ZN(n7820) );
  NAND2_X1 U8789 ( .A1(n7824), .A2(n7822), .ZN(n7821) );
  NAND2_X1 U8790 ( .A1(n8100), .A2(n8099), .ZN(n14935) );
  AOI21_X1 U8791 ( .B1(n8101), .B2(n12677), .A(n12686), .ZN(n8099) );
  OAI21_X1 U8792 ( .B1(n12258), .B2(n8129), .A(n8127), .ZN(n12600) );
  INV_X1 U8793 ( .A(n9931), .ZN(n7631) );
  OR2_X1 U8794 ( .A1(n9884), .A2(n9883), .ZN(n8513) );
  OR2_X1 U8795 ( .A1(n9843), .A2(n15340), .ZN(n9306) );
  INV_X1 U8796 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n15992) );
  AOI21_X1 U8797 ( .B1(n10351), .B2(P1_REG1_REG_6__SCAN_IN), .A(n10350), .ZN(
        n10353) );
  AOI21_X1 U8798 ( .B1(n10425), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10420), .ZN(
        n15034) );
  NAND2_X1 U8799 ( .A1(n10706), .A2(n10707), .ZN(n10705) );
  INV_X1 U8800 ( .A(n9274), .ZN(n7706) );
  NOR2_X1 U8801 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7705) );
  NOR2_X1 U8802 ( .A1(n15094), .A2(n8002), .ZN(n8001) );
  INV_X1 U8803 ( .A(n8003), .ZN(n8002) );
  INV_X1 U8804 ( .A(n12577), .ZN(n8470) );
  INV_X1 U8805 ( .A(n8473), .ZN(n8471) );
  NAND2_X1 U8806 ( .A1(n9166), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9845) );
  OAI21_X1 U8807 ( .B1(n8011), .B2(n15132), .A(n15137), .ZN(n15131) );
  NAND2_X1 U8808 ( .A1(n8012), .A2(n8011), .ZN(n15145) );
  OR2_X1 U8809 ( .A1(n15395), .A2(n15146), .ZN(n12576) );
  AND2_X1 U8810 ( .A1(n8325), .A2(n8324), .ZN(n15138) );
  NAND2_X1 U8811 ( .A1(n15173), .A2(n15146), .ZN(n8324) );
  NAND2_X1 U8812 ( .A1(n8478), .A2(n15282), .ZN(n8474) );
  AOI21_X1 U8813 ( .B1(n8478), .B2(n7487), .A(n7467), .ZN(n8476) );
  NAND2_X1 U8814 ( .A1(n15251), .A2(n12561), .ZN(n15229) );
  NOR2_X1 U8815 ( .A1(n15440), .A2(n8007), .ZN(n8006) );
  INV_X1 U8816 ( .A(n8008), .ZN(n8007) );
  OAI21_X1 U8817 ( .B1(n12553), .B2(n7887), .A(n7619), .ZN(n15287) );
  AND2_X1 U8818 ( .A1(n7886), .A2(n12557), .ZN(n7619) );
  NAND2_X1 U8819 ( .A1(n7553), .A2(n8327), .ZN(n7886) );
  AND2_X1 U8820 ( .A1(n9553), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9568) );
  NAND2_X1 U8821 ( .A1(n7889), .A2(n7888), .ZN(n15302) );
  NAND2_X1 U8822 ( .A1(n12343), .A2(n12574), .ZN(n15321) );
  NAND2_X1 U8823 ( .A1(n12343), .A2(n8010), .ZN(n15319) );
  OAI22_X1 U8824 ( .A1(n11862), .A2(n8455), .B1(n8457), .B2(n8454), .ZN(n12313) );
  NAND2_X1 U8825 ( .A1(n8459), .A2(n8456), .ZN(n8455) );
  INV_X1 U8826 ( .A(n8459), .ZN(n8454) );
  INV_X1 U8827 ( .A(n8461), .ZN(n8456) );
  AND2_X1 U8828 ( .A1(n15462), .A2(n12305), .ZN(n12343) );
  AOI21_X1 U8829 ( .B1(n8321), .B2(n8323), .A(n7538), .ZN(n8319) );
  NOR2_X1 U8830 ( .A1(n8458), .A2(n12303), .ZN(n8457) );
  NOR2_X1 U8831 ( .A1(n8461), .A2(n12150), .ZN(n8458) );
  NOR2_X1 U8832 ( .A1(n12153), .A2(n14965), .ZN(n8461) );
  NOR2_X1 U8833 ( .A1(n12162), .A2(n15470), .ZN(n12305) );
  OR2_X1 U8834 ( .A1(n11865), .A2(n12153), .ZN(n12162) );
  AND2_X1 U8835 ( .A1(n11862), .A2(n12150), .ZN(n12155) );
  OR2_X1 U8836 ( .A1(n9437), .A2(n9436), .ZN(n9454) );
  OR2_X1 U8837 ( .A1(n9454), .A2(n9453), .ZN(n9480) );
  AOI21_X1 U8838 ( .B1(n11734), .B2(n8426), .A(n7493), .ZN(n8425) );
  INV_X1 U8839 ( .A(n11732), .ZN(n8426) );
  OAI21_X1 U8840 ( .B1(n11539), .B2(n8333), .A(n8331), .ZN(n11758) );
  INV_X1 U8841 ( .A(n8332), .ZN(n8331) );
  OAI21_X1 U8842 ( .B1(n8334), .B2(n8333), .A(n11745), .ZN(n8332) );
  INV_X1 U8843 ( .A(n11743), .ZN(n8333) );
  NAND2_X1 U8844 ( .A1(n11744), .A2(n11743), .ZN(n11746) );
  NAND2_X1 U8845 ( .A1(n8005), .A2(n8004), .ZN(n11817) );
  NAND2_X1 U8846 ( .A1(n11539), .A2(n8334), .ZN(n11744) );
  NAND2_X1 U8847 ( .A1(n11539), .A2(n11538), .ZN(n11541) );
  INV_X1 U8848 ( .A(n8005), .ZN(n11737) );
  AND2_X1 U8849 ( .A1(n11159), .A2(n16463), .ZN(n10897) );
  AND3_X1 U8850 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n9378) );
  NAND2_X1 U8851 ( .A1(n10859), .A2(n10858), .ZN(n10861) );
  NAND2_X1 U8852 ( .A1(n11112), .A2(n10857), .ZN(n11157) );
  INV_X1 U8853 ( .A(n10524), .ZN(n10520) );
  AND2_X1 U8854 ( .A1(n7876), .A2(n7875), .ZN(n10523) );
  OAI21_X1 U8855 ( .B1(n10522), .B2(n10517), .A(n16394), .ZN(n7876) );
  NOR2_X1 U8856 ( .A1(n10439), .A2(n11207), .ZN(n9975) );
  AND2_X1 U8857 ( .A1(n7455), .A2(n12592), .ZN(n10438) );
  OR2_X1 U8858 ( .A1(n10266), .A2(n9285), .ZN(n9286) );
  CLKBUF_X1 U8859 ( .A(n9970), .Z(n9974) );
  INV_X1 U8860 ( .A(n15367), .ZN(n8335) );
  INV_X1 U8861 ( .A(n8325), .ZN(n15159) );
  AND2_X1 U8862 ( .A1(n15921), .A2(n10266), .ZN(n15408) );
  NAND2_X1 U8863 ( .A1(n9617), .A2(n9616), .ZN(n15435) );
  INV_X1 U8864 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n15688) );
  NAND2_X1 U8865 ( .A1(n11110), .A2(n8000), .ZN(n16430) );
  INV_X1 U8866 ( .A(n16542), .ZN(n16445) );
  AND2_X1 U8867 ( .A1(n11731), .A2(n9998), .ZN(n10491) );
  AND2_X1 U8868 ( .A1(n10264), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9948) );
  XNOR2_X1 U8869 ( .A(n9824), .B(n9823), .ZN(n14798) );
  NAND2_X1 U8870 ( .A1(n9782), .A2(n9781), .ZN(n9785) );
  INV_X1 U8871 ( .A(n9265), .ZN(n7701) );
  NOR2_X1 U8872 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n7700) );
  NOR2_X1 U8873 ( .A1(n9156), .A2(n9933), .ZN(n9157) );
  NAND2_X1 U8874 ( .A1(n8230), .A2(n9260), .ZN(n9764) );
  NAND2_X1 U8875 ( .A1(n9256), .A2(n8234), .ZN(n8230) );
  INV_X1 U8876 ( .A(n8235), .ZN(n8234) );
  NAND2_X1 U8877 ( .A1(n9598), .A2(n7839), .ZN(n9274) );
  AND2_X1 U8878 ( .A1(n15684), .A2(n15692), .ZN(n7839) );
  XNOR2_X1 U8879 ( .A(n9644), .B(n9643), .ZN(n12590) );
  INV_X1 U8880 ( .A(n8288), .ZN(n9596) );
  NAND2_X1 U8881 ( .A1(n9228), .A2(n9227), .ZN(n9595) );
  XNOR2_X1 U8882 ( .A(n9522), .B(n9521), .ZN(n11901) );
  AND2_X1 U8883 ( .A1(n9541), .A2(n9527), .ZN(n10675) );
  NAND2_X1 U8884 ( .A1(n8199), .A2(n9200), .ZN(n9445) );
  NAND2_X1 U8885 ( .A1(n9425), .A2(n9198), .ZN(n8199) );
  OR2_X1 U8886 ( .A1(n9560), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9446) );
  OR2_X1 U8887 ( .A1(n9387), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n9560) );
  XNOR2_X1 U8888 ( .A(n15984), .B(n15982), .ZN(n15983) );
  AOI21_X1 U8889 ( .B1(n15990), .B2(n15989), .A(n16273), .ZN(n15993) );
  OAI21_X1 U8890 ( .B1(n15934), .B2(n15978), .A(n15976), .ZN(n16003) );
  XNOR2_X1 U8891 ( .A(n15937), .B(n15938), .ZN(n16006) );
  NOR2_X1 U8892 ( .A1(n15943), .A2(n15942), .ZN(n15974) );
  NOR2_X1 U8893 ( .A1(n15975), .A2(n15005), .ZN(n15942) );
  OAI21_X1 U8894 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(n15948), .A(n15947), .ZN(
        n15971) );
  AOI22_X1 U8895 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n15954), .B1(n15969), 
        .B2(n15953), .ZN(n16019) );
  OR2_X1 U8896 ( .A1(n15964), .A2(n15963), .ZN(n16035) );
  NAND2_X1 U8897 ( .A1(n13152), .A2(n12494), .ZN(n12788) );
  INV_X1 U8898 ( .A(n8414), .ZN(n8413) );
  NAND2_X1 U8899 ( .A1(n8949), .A2(n8948), .ZN(n13469) );
  AND3_X1 U8900 ( .A1(n8716), .A2(n8715), .A3(n8714), .ZN(n12326) );
  AND4_X1 U8901 ( .A1(n13004), .A2(n9046), .A3(n9045), .A4(n9044), .ZN(n12838)
         );
  OR2_X1 U8902 ( .A1(n13180), .A2(n8384), .ZN(n7686) );
  AND2_X1 U8903 ( .A1(n8381), .A2(n13183), .ZN(n7687) );
  NAND2_X1 U8904 ( .A1(n9029), .A2(n9028), .ZN(n12978) );
  OR2_X1 U8905 ( .A1(n7461), .A2(n15498), .ZN(n9028) );
  CLKBUF_X1 U8906 ( .A(n13110), .Z(n13111) );
  CLKBUF_X1 U8907 ( .A(n13105), .Z(n13106) );
  AND2_X1 U8908 ( .A1(n8370), .A2(n8368), .ZN(n12320) );
  NAND2_X1 U8909 ( .A1(n8370), .A2(n8372), .ZN(n12122) );
  AND2_X1 U8910 ( .A1(n8757), .A2(n8756), .ZN(n13157) );
  NAND2_X1 U8911 ( .A1(n12491), .A2(n12490), .ZN(n13152) );
  NAND2_X1 U8912 ( .A1(n8937), .A2(n8936), .ZN(n13486) );
  AND3_X1 U8913 ( .A1(n8736), .A2(n8735), .A3(n8734), .ZN(n12919) );
  AND2_X1 U8914 ( .A1(n11697), .A2(n11694), .ZN(n11695) );
  AND4_X1 U8915 ( .A1(n9018), .A2(n9017), .A3(n9016), .A4(n9015), .ZN(n13421)
         );
  AOI21_X1 U8916 ( .B1(n8376), .B2(n8378), .A(n7520), .ZN(n8374) );
  NOR2_X1 U8917 ( .A1(n13045), .A2(n13044), .ZN(n7715) );
  XNOR2_X1 U8918 ( .A(n7620), .B(n10592), .ZN(n13057) );
  INV_X1 U8919 ( .A(n13421), .ZN(n13392) );
  INV_X1 U8920 ( .A(n13438), .ZN(n13207) );
  NAND2_X1 U8921 ( .A1(n8631), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8954) );
  INV_X1 U8922 ( .A(n13514), .ZN(n13479) );
  INV_X1 U8923 ( .A(n13569), .ZN(n13211) );
  INV_X1 U8924 ( .A(n13157), .ZN(n13216) );
  OAI21_X1 U8925 ( .B1(P3_IR_REG_31__SCAN_IN), .B2(P3_IR_REG_1__SCAN_IN), .A(
        n7778), .ZN(n7777) );
  NAND2_X1 U8926 ( .A1(n7559), .A2(P3_IR_REG_1__SCAN_IN), .ZN(n7778) );
  OR2_X1 U8927 ( .A1(n11212), .A2(n16392), .ZN(n11213) );
  OR2_X1 U8928 ( .A1(n10970), .A2(n10969), .ZN(n11285) );
  NAND2_X1 U8929 ( .A1(n8022), .A2(n11407), .ZN(n11019) );
  NAND2_X1 U8930 ( .A1(n7760), .A2(n7758), .ZN(n11037) );
  INV_X1 U8931 ( .A(n7766), .ZN(n11836) );
  NOR2_X1 U8932 ( .A1(n11831), .A2(n8023), .ZN(n11834) );
  INV_X1 U8933 ( .A(n11434), .ZN(n8023) );
  NOR2_X1 U8934 ( .A1(n7782), .A2(n7532), .ZN(n12184) );
  NOR2_X1 U8935 ( .A1(n7521), .A2(n7779), .ZN(n13231) );
  NOR2_X1 U8936 ( .A1(n13246), .A2(n13247), .ZN(n13250) );
  INV_X1 U8937 ( .A(n8245), .ZN(n13293) );
  INV_X1 U8938 ( .A(n13294), .ZN(n8244) );
  AND2_X1 U8939 ( .A1(n8831), .A2(n8848), .ZN(n13296) );
  NOR2_X1 U8940 ( .A1(n13277), .A2(n13278), .ZN(n13280) );
  INV_X1 U8941 ( .A(n13328), .ZN(n7774) );
  NOR2_X1 U8942 ( .A1(n13303), .A2(n13304), .ZN(n13324) );
  INV_X1 U8943 ( .A(n7781), .ZN(n13333) );
  OAI21_X1 U8944 ( .B1(n13303), .B2(n7772), .A(n7771), .ZN(n13350) );
  NAND2_X1 U8945 ( .A1(n7773), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n7772) );
  NAND2_X1 U8946 ( .A1(n13325), .A2(n7773), .ZN(n7771) );
  INV_X1 U8947 ( .A(n13326), .ZN(n7773) );
  NAND2_X1 U8948 ( .A1(n7808), .A2(n13394), .ZN(n13595) );
  NAND2_X1 U8949 ( .A1(n13427), .A2(n12843), .ZN(n13414) );
  NAND2_X1 U8950 ( .A1(n13451), .A2(n8974), .ZN(n13437) );
  NAND2_X1 U8951 ( .A1(n8896), .A2(n8895), .ZN(n13513) );
  NAND2_X1 U8952 ( .A1(n8352), .A2(n12944), .ZN(n13523) );
  NAND2_X1 U8953 ( .A1(n13533), .A2(n13535), .ZN(n8352) );
  NAND2_X1 U8954 ( .A1(n13537), .A2(n8877), .ZN(n13524) );
  NAND2_X1 U8955 ( .A1(n13566), .A2(n12934), .ZN(n13547) );
  NAND2_X1 U8956 ( .A1(n7813), .A2(n8802), .ZN(n13579) );
  NAND2_X1 U8957 ( .A1(n8770), .A2(n8769), .ZN(n13659) );
  INV_X1 U8958 ( .A(n12546), .ZN(n16559) );
  NAND2_X1 U8959 ( .A1(n11977), .A2(n8405), .ZN(n12397) );
  OR2_X1 U8960 ( .A1(n10690), .A2(n16400), .ZN(n13587) );
  NAND2_X1 U8961 ( .A1(n8079), .A2(n8662), .ZN(n11981) );
  NAND2_X1 U8962 ( .A1(n11809), .A2(n8648), .ZN(n11874) );
  AND3_X1 U8963 ( .A1(n8628), .A2(n8627), .A3(n8626), .ZN(n16456) );
  NAND2_X1 U8964 ( .A1(n11594), .A2(n13016), .ZN(n11593) );
  NAND2_X1 U8965 ( .A1(n11302), .A2(n12871), .ZN(n11594) );
  OR2_X1 U8966 ( .A1(n10924), .A2(n10621), .ZN(n16405) );
  OR2_X1 U8967 ( .A1(n9027), .A2(n10176), .ZN(n8572) );
  NAND2_X1 U8968 ( .A1(n7613), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n7612) );
  INV_X1 U8969 ( .A(n16405), .ZN(n16388) );
  NAND2_X1 U8970 ( .A1(n16565), .A2(n16471), .ZN(n13657) );
  INV_X1 U8971 ( .A(n13054), .ZN(n13667) );
  NAND2_X1 U8972 ( .A1(n7483), .A2(n7809), .ZN(n7808) );
  INV_X1 U8973 ( .A(n13395), .ZN(n7809) );
  INV_X1 U8974 ( .A(n13104), .ZN(n13685) );
  NAND2_X1 U8975 ( .A1(n8812), .A2(n8811), .ZN(n13726) );
  NAND2_X1 U8976 ( .A1(n8795), .A2(n8794), .ZN(n13730) );
  NAND2_X1 U8977 ( .A1(n11873), .A2(n12888), .ZN(n11872) );
  NAND2_X1 U8978 ( .A1(n11803), .A2(n9069), .ZN(n11873) );
  AND2_X1 U8979 ( .A1(n10925), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13737) );
  INV_X1 U8980 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8535) );
  XNOR2_X1 U8981 ( .A(n8537), .B(n8536), .ZN(n13071) );
  INV_X1 U8982 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n8536) );
  NAND2_X1 U8983 ( .A1(n13742), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8537) );
  INV_X1 U8984 ( .A(n8540), .ZN(n13748) );
  OAI21_X1 U8985 ( .B1(n9026), .B2(n9025), .A(n9039), .ZN(n12784) );
  OR2_X1 U8986 ( .A1(n8999), .A2(n8998), .ZN(n9000) );
  NAND2_X1 U8987 ( .A1(n7618), .A2(n7615), .ZN(n12042) );
  OR2_X1 U8988 ( .A1(n9101), .A2(n8534), .ZN(n7618) );
  NOR2_X1 U8989 ( .A1(n7617), .A2(n7616), .ZN(n7615) );
  INV_X1 U8990 ( .A(SI_25_), .ZN(n15704) );
  XNOR2_X1 U8991 ( .A(n9097), .B(n9096), .ZN(n11922) );
  OAI21_X1 U8992 ( .B1(n9095), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9097) );
  XNOR2_X1 U8993 ( .A(n9055), .B(P3_IR_REG_22__SCAN_IN), .ZN(n13064) );
  NAND2_X1 U8994 ( .A1(n9054), .A2(n9053), .ZN(n9092) );
  NAND2_X1 U8995 ( .A1(n8914), .A2(n8913), .ZN(n8927) );
  NAND2_X1 U8996 ( .A1(n8900), .A2(n8913), .ZN(n8901) );
  INV_X1 U8997 ( .A(SI_20_), .ZN(n10656) );
  OAI21_X1 U8998 ( .B1(n8864), .B2(n8057), .A(n8055), .ZN(n8898) );
  NAND2_X1 U8999 ( .A1(n8879), .A2(n8878), .ZN(n8882) );
  NAND2_X1 U9000 ( .A1(n8824), .A2(n8823), .ZN(n8843) );
  NAND2_X1 U9001 ( .A1(n8821), .A2(n8820), .ZN(n8824) );
  INV_X1 U9002 ( .A(SI_16_), .ZN(n15520) );
  INV_X1 U9003 ( .A(SI_14_), .ZN(n15525) );
  INV_X1 U9004 ( .A(SI_13_), .ZN(n15724) );
  OAI21_X1 U9005 ( .B1(n8729), .B2(n8063), .A(n8061), .ZN(n8762) );
  NAND2_X1 U9006 ( .A1(n8741), .A2(n8740), .ZN(n8744) );
  INV_X1 U9007 ( .A(SI_11_), .ZN(n10208) );
  OAI21_X1 U9008 ( .B1(n8677), .B2(n8051), .A(n8049), .ZN(n8707) );
  NAND2_X1 U9009 ( .A1(n8691), .A2(n8690), .ZN(n8694) );
  NAND2_X1 U9010 ( .A1(n8642), .A2(n8641), .ZN(n8656) );
  OR2_X1 U9011 ( .A1(n8640), .A2(n7787), .ZN(n11418) );
  NOR2_X1 U9012 ( .A1(n8418), .A2(n8416), .ZN(n8636) );
  NAND2_X1 U9013 ( .A1(n8554), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U9014 ( .A1(n13739), .A2(n10184), .ZN(n8016) );
  OR2_X1 U9015 ( .A1(n10143), .A2(n12070), .ZN(n10272) );
  AND2_X1 U9016 ( .A1(n7911), .A2(n12733), .ZN(n7910) );
  NAND2_X1 U9017 ( .A1(n7913), .A2(n7915), .ZN(n7911) );
  NAND2_X1 U9018 ( .A1(n10048), .A2(n11184), .ZN(n8187) );
  NAND2_X1 U9019 ( .A1(n10051), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U9020 ( .A1(n7906), .A2(n10740), .ZN(n10984) );
  NAND2_X1 U9021 ( .A1(n12767), .A2(n10729), .ZN(n7906) );
  NAND2_X1 U9022 ( .A1(n13940), .A2(n13939), .ZN(n13938) );
  NOR2_X1 U9023 ( .A1(n7908), .A2(n7603), .ZN(n7904) );
  NOR2_X1 U9024 ( .A1(n7603), .A2(n7903), .ZN(n7902) );
  INV_X1 U9025 ( .A(n13983), .ZN(n13987) );
  INV_X1 U9026 ( .A(n13967), .ZN(n13957) );
  NAND2_X1 U9027 ( .A1(n7912), .A2(n11916), .ZN(n12731) );
  NAND2_X1 U9028 ( .A1(n12728), .A2(n11899), .ZN(n7912) );
  OR2_X1 U9029 ( .A1(n10163), .A2(n14290), .ZN(n13975) );
  OAI21_X1 U9030 ( .B1(n11344), .B2(n7470), .A(n8142), .ZN(n12720) );
  NAND2_X1 U9031 ( .A1(n10765), .A2(n10151), .ZN(n7916) );
  NOR2_X1 U9032 ( .A1(n12435), .A2(n8145), .ZN(n8144) );
  INV_X1 U9033 ( .A(n8148), .ZN(n8145) );
  NAND2_X1 U9034 ( .A1(n8146), .A2(n8148), .ZN(n12436) );
  AND2_X1 U9035 ( .A1(n10660), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13972) );
  NAND2_X1 U9036 ( .A1(n8155), .A2(n8156), .ZN(n13970) );
  NAND2_X1 U9037 ( .A1(n12095), .A2(n12104), .ZN(n12750) );
  NAND2_X1 U9038 ( .A1(n12094), .A2(n12093), .ZN(n14108) );
  OAI22_X1 U9039 ( .A1(n8296), .A2(n14345), .B1(n14202), .B2(n12091), .ZN(
        n12092) );
  AND2_X1 U9040 ( .A1(n14299), .A2(n14288), .ZN(n7667) );
  INV_X1 U9041 ( .A(n8295), .ZN(n8294) );
  CLKBUF_X1 U9042 ( .A(n13984), .Z(n14323) );
  NOR2_X1 U9043 ( .A1(n16124), .A2(n16123), .ZN(n16122) );
  NOR2_X1 U9044 ( .A1(n16122), .A2(n7693), .ZN(n16136) );
  AND2_X1 U9045 ( .A1(n11186), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7693) );
  NOR2_X1 U9046 ( .A1(n16153), .A2(n16152), .ZN(n16151) );
  NOR2_X1 U9047 ( .A1(n16178), .A2(n16177), .ZN(n16176) );
  NOR2_X1 U9048 ( .A1(n12410), .A2(n12272), .ZN(n14347) );
  AND2_X1 U9049 ( .A1(n14456), .A2(n14455), .ZN(n14669) );
  NAND2_X1 U9050 ( .A1(n8301), .A2(n8299), .ZN(n14476) );
  NAND2_X1 U9051 ( .A1(n8301), .A2(n14446), .ZN(n14474) );
  NAND2_X1 U9052 ( .A1(n13754), .A2(n13753), .ZN(n14672) );
  NAND2_X1 U9053 ( .A1(n14505), .A2(n14406), .ZN(n14487) );
  NAND2_X1 U9054 ( .A1(n14525), .A2(n14441), .ZN(n14511) );
  NAND2_X1 U9055 ( .A1(n13780), .A2(n13779), .ZN(n14708) );
  NAND2_X1 U9056 ( .A1(n7950), .A2(n7951), .ZN(n14572) );
  NAND2_X1 U9057 ( .A1(n14608), .A2(n14429), .ZN(n14587) );
  NAND2_X1 U9058 ( .A1(n12451), .A2(n12450), .ZN(n14639) );
  NAND2_X1 U9059 ( .A1(n8167), .A2(n8170), .ZN(n14635) );
  NAND2_X1 U9060 ( .A1(n7937), .A2(n7941), .ZN(n12027) );
  NAND2_X1 U9061 ( .A1(n11940), .A2(n7942), .ZN(n7937) );
  NAND2_X1 U9062 ( .A1(n7943), .A2(n7944), .ZN(n11941) );
  OR2_X1 U9063 ( .A1(n11940), .A2(n11939), .ZN(n7943) );
  NAND2_X1 U9064 ( .A1(n8181), .A2(n8182), .ZN(n11680) );
  NAND2_X1 U9065 ( .A1(n8307), .A2(n11054), .ZN(n11056) );
  NAND2_X1 U9066 ( .A1(n10822), .A2(n10821), .ZN(n10823) );
  OR2_X1 U9067 ( .A1(n10131), .A2(n10130), .ZN(n14553) );
  NAND2_X1 U9068 ( .A1(n11900), .A2(n10180), .ZN(n8293) );
  INV_X1 U9069 ( .A(n14622), .ZN(n14646) );
  INV_X1 U9070 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n7662) );
  NOR2_X1 U9071 ( .A1(n7990), .A2(n14734), .ZN(n7663) );
  INV_X1 U9072 ( .A(n14382), .ZN(n14753) );
  INV_X1 U9073 ( .A(n7690), .ZN(n7689) );
  INV_X1 U9074 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n7658) );
  NAND2_X1 U9075 ( .A1(n14813), .A2(n14201), .ZN(n7856) );
  NAND2_X1 U9076 ( .A1(n12213), .A2(n12212), .ZN(n14789) );
  INV_X1 U9077 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n14793) );
  NOR2_X1 U9078 ( .A1(n8166), .A2(n10335), .ZN(n7683) );
  XNOR2_X1 U9079 ( .A(n9957), .B(P2_IR_REG_26__SCAN_IN), .ZN(n14809) );
  AND2_X1 U9080 ( .A1(n9960), .A2(n9959), .ZN(n14814) );
  NOR2_X1 U9081 ( .A1(n10335), .A2(n9953), .ZN(n10080) );
  INV_X1 U9082 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10698) );
  INV_X1 U9083 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n12091) );
  INV_X1 U9084 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10402) );
  INV_X1 U9085 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10291) );
  INV_X1 U9086 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10255) );
  INV_X1 U9087 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10247) );
  INV_X1 U9088 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10240) );
  INV_X1 U9089 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10237) );
  INV_X1 U9090 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10220) );
  INV_X1 U9091 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10215) );
  INV_X1 U9092 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10206) );
  INV_X1 U9093 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10193) );
  INV_X1 U9094 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10181) );
  INV_X1 U9095 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10172) );
  INV_X1 U9096 ( .A(n8131), .ZN(n12595) );
  NAND2_X1 U9097 ( .A1(n11969), .A2(n11968), .ZN(n12061) );
  AND2_X1 U9098 ( .A1(n7827), .A2(n7494), .ZN(n11666) );
  NAND2_X1 U9099 ( .A1(n7834), .A2(n7832), .ZN(n14860) );
  INV_X1 U9100 ( .A(n7835), .ZN(n7832) );
  OAI21_X1 U9101 ( .B1(n14897), .B2(n12677), .A(n8101), .ZN(n14867) );
  NAND2_X1 U9102 ( .A1(n14896), .A2(n12678), .ZN(n14868) );
  INV_X1 U9103 ( .A(n14966), .ZN(n11961) );
  NAND2_X1 U9104 ( .A1(n11722), .A2(n8105), .ZN(n11969) );
  OAI21_X1 U9105 ( .B1(n14924), .B2(n8126), .A(n8123), .ZN(n14907) );
  NAND2_X1 U9106 ( .A1(n7834), .A2(n7829), .ZN(n14916) );
  NOR2_X1 U9107 ( .A1(n7831), .A2(n7830), .ZN(n7829) );
  INV_X1 U9108 ( .A(n14917), .ZN(n7830) );
  INV_X1 U9109 ( .A(n7833), .ZN(n7831) );
  AND2_X1 U9110 ( .A1(n7834), .A2(n7833), .ZN(n14918) );
  NOR2_X1 U9111 ( .A1(n10499), .A2(n10498), .ZN(n14915) );
  AOI21_X1 U9112 ( .B1(n7608), .B2(n8111), .A(n8106), .ZN(n11458) );
  INV_X1 U9113 ( .A(n8113), .ZN(n8106) );
  INV_X1 U9114 ( .A(n14844), .ZN(n14958) );
  INV_X1 U9115 ( .A(n11466), .ZN(n14947) );
  AND2_X1 U9116 ( .A1(n10481), .A2(n15331), .ZN(n14955) );
  OR2_X1 U9117 ( .A1(n9808), .A2(n10307), .ZN(n9327) );
  AOI21_X1 U9118 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n16341), .A(n16348), .ZN(
        n10364) );
  AND2_X1 U9119 ( .A1(n15002), .A2(n15001), .ZN(n15018) );
  AND2_X1 U9120 ( .A1(n15034), .A2(n15033), .ZN(n15035) );
  NOR2_X1 U9121 ( .A1(n10423), .A2(n10422), .ZN(n10671) );
  XNOR2_X1 U9122 ( .A(n11569), .B(n11382), .ZN(n11377) );
  NOR2_X1 U9123 ( .A1(n11377), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11574) );
  XNOR2_X1 U9124 ( .A(n7632), .B(n9630), .ZN(n15063) );
  NAND2_X1 U9125 ( .A1(n16259), .A2(n15052), .ZN(n7632) );
  NAND2_X1 U9126 ( .A1(n9836), .A2(n9835), .ZN(n15351) );
  INV_X1 U9127 ( .A(n15092), .ZN(n8336) );
  AND2_X1 U9128 ( .A1(n12571), .A2(n12570), .ZN(n15374) );
  NAND2_X1 U9129 ( .A1(n15140), .A2(n12577), .ZN(n15123) );
  INV_X1 U9130 ( .A(n15183), .ZN(n15402) );
  NAND2_X1 U9131 ( .A1(n8446), .A2(n8450), .ZN(n15178) );
  NAND2_X1 U9132 ( .A1(n15216), .A2(n8447), .ZN(n8446) );
  INV_X1 U9133 ( .A(n15408), .ZN(n15206) );
  NAND2_X1 U9134 ( .A1(n15216), .A2(n8452), .ZN(n15195) );
  NAND2_X1 U9135 ( .A1(n7884), .A2(n12563), .ZN(n15193) );
  NAND2_X1 U9136 ( .A1(n15235), .A2(n12562), .ZN(n15213) );
  AOI21_X1 U9137 ( .B1(n8481), .B2(n8480), .A(n7487), .ZN(n15249) );
  INV_X1 U9138 ( .A(n15280), .ZN(n8481) );
  NOR2_X1 U9139 ( .A1(n15280), .A2(n8483), .ZN(n15276) );
  NAND2_X1 U9140 ( .A1(n8428), .A2(n8432), .ZN(n15308) );
  OR2_X1 U9141 ( .A1(n12340), .A2(n8433), .ZN(n8428) );
  NAND2_X1 U9142 ( .A1(n8330), .A2(n12554), .ZN(n15326) );
  NAND2_X1 U9143 ( .A1(n12553), .A2(n12552), .ZN(n8330) );
  NAND2_X1 U9144 ( .A1(n12572), .A2(n8435), .ZN(n15318) );
  NAND2_X1 U9145 ( .A1(n8320), .A2(n12154), .ZN(n12304) );
  NAND2_X1 U9146 ( .A1(n9470), .A2(n9469), .ZN(n11963) );
  NAND2_X1 U9147 ( .A1(n11735), .A2(n11734), .ZN(n11753) );
  NAND2_X1 U9148 ( .A1(n11733), .A2(n11732), .ZN(n11735) );
  INV_X1 U9149 ( .A(n16429), .ZN(n14843) );
  NAND2_X1 U9150 ( .A1(n15338), .A2(n10438), .ZN(n15221) );
  INV_X1 U9151 ( .A(n15221), .ZN(n15347) );
  NAND2_X1 U9152 ( .A1(n15380), .A2(n15381), .ZN(n15483) );
  NAND2_X1 U9153 ( .A1(n8217), .A2(n8214), .ZN(n9831) );
  NAND2_X1 U9154 ( .A1(n8217), .A2(n9792), .ZN(n9795) );
  INV_X1 U9155 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9159) );
  XNOR2_X1 U9156 ( .A(n9854), .B(n9853), .ZN(n14802) );
  XNOR2_X1 U9157 ( .A(n9939), .B(n9938), .ZN(n15920) );
  OAI21_X1 U9158 ( .B1(n7486), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9939) );
  XNOR2_X1 U9159 ( .A(n9932), .B(P1_IR_REG_24__SCAN_IN), .ZN(n12317) );
  NAND2_X1 U9160 ( .A1(n8205), .A2(n9250), .ZN(n9713) );
  NAND2_X1 U9161 ( .A1(n9248), .A2(n11956), .ZN(n8205) );
  INV_X1 U9162 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10632) );
  INV_X1 U9163 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10467) );
  INV_X1 U9164 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10403) );
  XNOR2_X1 U9165 ( .A(n9542), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11378) );
  INV_X1 U9166 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10341) );
  INV_X1 U9167 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10250) );
  INV_X1 U9168 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10248) );
  INV_X1 U9169 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10241) );
  INV_X1 U9170 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10232) );
  INV_X1 U9171 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10222) );
  INV_X1 U9172 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10211) );
  INV_X1 U9173 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10223) );
  INV_X1 U9174 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10198) );
  NOR2_X1 U9175 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n8427) );
  NOR2_X1 U9176 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9311) );
  INV_X1 U9177 ( .A(P2_RD_REG_SCAN_IN), .ZN(n8548) );
  XNOR2_X1 U9178 ( .A(n15983), .B(n7748), .ZN(n16326) );
  INV_X1 U9179 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7748) );
  XNOR2_X1 U9180 ( .A(n15981), .B(n7979), .ZN(n16280) );
  AND2_X1 U9181 ( .A1(n7747), .A2(n7746), .ZN(n16323) );
  OR2_X1 U9182 ( .A1(n16282), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n7747) );
  NOR2_X1 U9183 ( .A1(n16323), .A2(n16322), .ZN(n16321) );
  XNOR2_X1 U9184 ( .A(n16005), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n16285) );
  NOR2_X1 U9185 ( .A1(n16290), .A2(n16289), .ZN(n16288) );
  OAI21_X1 U9186 ( .B1(n16293), .B2(n16294), .A(P2_ADDR_REG_10__SCAN_IN), .ZN(
        n7975) );
  XNOR2_X1 U9187 ( .A(n16017), .B(n16016), .ZN(n16301) );
  NOR2_X1 U9188 ( .A1(n16304), .A2(n16303), .ZN(n16302) );
  INV_X1 U9189 ( .A(n16028), .ZN(n7734) );
  INV_X1 U9190 ( .A(n16031), .ZN(n7982) );
  NOR2_X1 U9191 ( .A1(n10609), .A2(n10614), .ZN(P3_U3897) );
  INV_X1 U9192 ( .A(n7742), .ZN(n7741) );
  OAI21_X1 U9193 ( .B1(n13677), .B2(n13199), .A(n13078), .ZN(n7742) );
  NAND2_X1 U9194 ( .A1(n11469), .A2(n8393), .ZN(n11472) );
  NOR2_X1 U9195 ( .A1(n10950), .A2(n8017), .ZN(n10951) );
  AOI21_X1 U9196 ( .B1(n13370), .B2(n13369), .A(n8255), .ZN(n8254) );
  NAND2_X1 U9197 ( .A1(n8256), .A2(n16336), .ZN(n7874) );
  NOR2_X1 U9198 ( .A1(n9135), .A2(n9134), .ZN(n9136) );
  OAI21_X1 U9199 ( .B1(n7804), .B2(n7805), .A(n7810), .ZN(P3_U3487) );
  INV_X1 U9200 ( .A(n7811), .ZN(n7810) );
  AND2_X1 U9201 ( .A1(n13395), .A2(n7806), .ZN(n7805) );
  AOI21_X1 U9202 ( .B1(n8088), .B2(n16569), .A(n7480), .ZN(n8087) );
  AOI21_X1 U9203 ( .B1(n10360), .B2(SI_2_), .A(n8014), .ZN(n10185) );
  NAND2_X1 U9204 ( .A1(n8016), .A2(n8015), .ZN(n8014) );
  NAND2_X1 U9205 ( .A1(n8147), .A2(n12368), .ZN(n12430) );
  NAND2_X1 U9206 ( .A1(n12753), .A2(n12353), .ZN(n8147) );
  NAND2_X1 U9207 ( .A1(n8208), .A2(n8207), .ZN(n14303) );
  INV_X1 U9208 ( .A(n8311), .ZN(n14451) );
  OAI21_X1 U9209 ( .B1(n14667), .B2(n14604), .A(n8312), .ZN(n8311) );
  AOI21_X1 U9210 ( .B1(n14663), .B2(n14650), .A(n14450), .ZN(n8312) );
  NAND2_X1 U9211 ( .A1(n7664), .A2(n7660), .ZN(P2_U3527) );
  NOR2_X1 U9212 ( .A1(n7663), .A2(n7661), .ZN(n7660) );
  NAND2_X1 U9213 ( .A1(n14755), .A2(n14740), .ZN(n7664) );
  NOR2_X1 U9214 ( .A1(n14740), .A2(n7662), .ZN(n7661) );
  NAND2_X1 U9215 ( .A1(n14240), .A2(n14790), .ZN(n7738) );
  NAND2_X1 U9216 ( .A1(n7659), .A2(n7656), .ZN(P2_U3495) );
  NOR2_X1 U9217 ( .A1(n7657), .A2(n7600), .ZN(n7656) );
  NAND2_X1 U9218 ( .A1(n14755), .A2(n16534), .ZN(n7659) );
  NOR2_X1 U9219 ( .A1(n16534), .A2(n7658), .ZN(n7657) );
  NAND2_X1 U9220 ( .A1(n8118), .A2(n12710), .ZN(n8117) );
  NAND2_X1 U9221 ( .A1(n7629), .A2(n12047), .ZN(n9947) );
  INV_X1 U9222 ( .A(n10130), .ZN(n14366) );
  NAND2_X1 U9223 ( .A1(n12059), .A2(n12058), .ZN(n7466) );
  AND2_X1 U9224 ( .A1(n8482), .A2(n15231), .ZN(n7467) );
  NAND2_X1 U9225 ( .A1(n11343), .A2(n11342), .ZN(n14068) );
  INV_X1 U9226 ( .A(n14068), .ZN(n7988) );
  NAND2_X1 U9227 ( .A1(n12016), .A2(n12015), .ZN(n14102) );
  INV_X1 U9228 ( .A(n14102), .ZN(n7739) );
  NOR2_X1 U9229 ( .A1(n7945), .A2(n14265), .ZN(n7942) );
  AND2_X1 U9230 ( .A1(n12138), .A2(n12137), .ZN(n7469) );
  AND2_X1 U9231 ( .A1(n11602), .A2(n11601), .ZN(n7470) );
  AND2_X1 U9232 ( .A1(n8413), .A2(n13133), .ZN(n7471) );
  NOR2_X1 U9233 ( .A1(n13486), .A2(n13499), .ZN(n7472) );
  NAND2_X1 U9234 ( .A1(n9681), .A2(n9680), .ZN(n12645) );
  INV_X1 U9235 ( .A(n15388), .ZN(n8011) );
  NOR2_X1 U9236 ( .A1(n8471), .A2(n8470), .ZN(n8469) );
  INV_X1 U9237 ( .A(n8469), .ZN(n8467) );
  INV_X1 U9238 ( .A(n8068), .ZN(n8069) );
  OR2_X1 U9239 ( .A1(n14047), .A2(n14049), .ZN(n7473) );
  AND2_X1 U9240 ( .A1(n14672), .A2(n14447), .ZN(n7474) );
  AND4_X1 U9241 ( .A1(n8579), .A2(n8578), .A3(n8577), .A4(n8576), .ZN(n11590)
         );
  AND2_X1 U9242 ( .A1(n13118), .A2(n13584), .ZN(n7475) );
  OR2_X1 U9243 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n16005), .ZN(n7476) );
  AND2_X1 U9244 ( .A1(n14089), .A2(n14091), .ZN(n7477) );
  OR2_X1 U9245 ( .A1(n14136), .A2(n14135), .ZN(n7478) );
  OR2_X1 U9246 ( .A1(n14172), .A2(n14171), .ZN(n7479) );
  OR2_X1 U9247 ( .A1(n8091), .A2(n7516), .ZN(n7480) );
  AND2_X1 U9248 ( .A1(n7540), .A2(n8135), .ZN(n7481) );
  AND2_X1 U9249 ( .A1(n9267), .A2(n9266), .ZN(n15376) );
  INV_X1 U9250 ( .A(n15376), .ZN(n9889) );
  NAND2_X1 U9251 ( .A1(n11296), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7482) );
  AND2_X1 U9252 ( .A1(n13389), .A2(n16377), .ZN(n7483) );
  INV_X1 U9253 ( .A(n7887), .ZN(n7888) );
  INV_X1 U9254 ( .A(n14240), .ZN(n14749) );
  NAND2_X1 U9255 ( .A1(n14180), .A2(n14179), .ZN(n14240) );
  AND2_X1 U9256 ( .A1(n7768), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7484) );
  INV_X1 U9257 ( .A(n10740), .ZN(n7908) );
  NOR2_X1 U9258 ( .A1(n10783), .A2(n10782), .ZN(n10904) );
  INV_X1 U9259 ( .A(n10904), .ZN(n8111) );
  AND2_X1 U9260 ( .A1(n11421), .A2(n7766), .ZN(n7485) );
  NAND2_X1 U9261 ( .A1(n10513), .A2(n14282), .ZN(n10148) );
  INV_X1 U9262 ( .A(n10148), .ZN(n14594) );
  INV_X1 U9263 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n10335) );
  NAND2_X1 U9264 ( .A1(n8288), .A2(n8133), .ZN(n7486) );
  INV_X1 U9265 ( .A(n12888), .ZN(n8399) );
  NOR2_X1 U9266 ( .A1(n15281), .A2(n15282), .ZN(n15280) );
  AND2_X1 U9267 ( .A1(n15274), .A2(n14891), .ZN(n7487) );
  NAND2_X1 U9268 ( .A1(n14927), .A2(n7837), .ZN(n7834) );
  NAND2_X1 U9269 ( .A1(n8861), .A2(n8860), .ZN(n8864) );
  AND2_X1 U9270 ( .A1(n10445), .A2(n10486), .ZN(n7488) );
  INV_X1 U9271 ( .A(n10196), .ZN(n10197) );
  INV_X1 U9272 ( .A(n14449), .ZN(n8313) );
  OR2_X1 U9273 ( .A1(n14708), .A2(n14431), .ZN(n7489) );
  AND2_X1 U9274 ( .A1(n9826), .A2(n9825), .ZN(n15366) );
  INV_X1 U9275 ( .A(n15366), .ZN(n15094) );
  AND2_X1 U9276 ( .A1(n14075), .A2(n14311), .ZN(n7490) );
  NAND2_X1 U9277 ( .A1(n8411), .A2(n9052), .ZN(n7491) );
  AND2_X1 U9278 ( .A1(n14124), .A2(n14123), .ZN(n7492) );
  NAND2_X1 U9279 ( .A1(n10691), .A2(n16375), .ZN(n16367) );
  INV_X1 U9280 ( .A(n14442), .ZN(n7855) );
  NOR2_X1 U9281 ( .A1(n11756), .A2(n14968), .ZN(n7493) );
  INV_X1 U9282 ( .A(n9338), .ZN(n7710) );
  INV_X1 U9283 ( .A(n14961), .ZN(n7885) );
  AND2_X1 U9284 ( .A1(n10126), .A2(n11958), .ZN(n13982) );
  XNOR2_X1 U9285 ( .A(n10030), .B(P2_IR_REG_1__SCAN_IN), .ZN(n16094) );
  INV_X1 U9286 ( .A(n16094), .ZN(n8493) );
  NAND2_X1 U9287 ( .A1(n11662), .A2(n11663), .ZN(n7494) );
  XNOR2_X1 U9288 ( .A(n9215), .B(n15724), .ZN(n9521) );
  AND2_X1 U9289 ( .A1(n15435), .A2(n15289), .ZN(n7495) );
  INV_X1 U9290 ( .A(n15143), .ZN(n8472) );
  AND2_X1 U9291 ( .A1(n13464), .A2(n8958), .ZN(n7496) );
  AND4_X1 U9292 ( .A1(n13041), .A2(n13040), .A3(n13039), .A4(n13047), .ZN(
        n7497) );
  INV_X1 U9293 ( .A(n14851), .ZN(n8126) );
  AND2_X1 U9294 ( .A1(n13596), .A2(n16561), .ZN(n7498) );
  AND3_X1 U9295 ( .A1(n8534), .A2(n7869), .A3(n8546), .ZN(n7499) );
  NAND2_X1 U9296 ( .A1(n13897), .A2(n13896), .ZN(n14465) );
  INV_X1 U9297 ( .A(n14465), .ZN(n7990) );
  INV_X1 U9298 ( .A(n13222), .ZN(n12884) );
  INV_X1 U9299 ( .A(n13215), .ZN(n12543) );
  NAND2_X1 U9300 ( .A1(n10266), .A2(n10171), .ZN(n9351) );
  NOR4_X1 U9301 ( .A1(n14526), .A2(n14540), .A3(n14562), .A4(n14274), .ZN(
        n7500) );
  INV_X1 U9302 ( .A(n14268), .ZN(n12139) );
  OR2_X1 U9303 ( .A1(n15402), .A2(n15198), .ZN(n7501) );
  NAND2_X1 U9304 ( .A1(n12818), .A2(n13133), .ZN(n13079) );
  AND2_X1 U9305 ( .A1(n12747), .A2(n12350), .ZN(n7502) );
  INV_X1 U9306 ( .A(n9452), .ZN(n8275) );
  INV_X1 U9307 ( .A(n9648), .ZN(n8278) );
  INV_X1 U9308 ( .A(n12567), .ZN(n15161) );
  OR2_X1 U9309 ( .A1(n13181), .A2(n13182), .ZN(n7503) );
  AOI21_X1 U9310 ( .B1(n13392), .B2(n12832), .A(n12833), .ZN(n13073) );
  AND2_X1 U9311 ( .A1(n8085), .A2(n9003), .ZN(n7504) );
  OR2_X1 U9312 ( .A1(n14677), .A2(n14407), .ZN(n7505) );
  NAND2_X1 U9313 ( .A1(n9601), .A2(n9600), .ZN(n15440) );
  AND2_X1 U9314 ( .A1(n12877), .A2(n12876), .ZN(n13016) );
  INV_X1 U9315 ( .A(n13016), .ZN(n8362) );
  NAND2_X1 U9316 ( .A1(n8427), .A2(n15862), .ZN(n9321) );
  OR2_X1 U9317 ( .A1(n9356), .A2(n9357), .ZN(n7507) );
  OR2_X1 U9318 ( .A1(n13179), .A2(n13438), .ZN(n12843) );
  INV_X1 U9319 ( .A(n15456), .ZN(n12574) );
  NAND2_X1 U9320 ( .A1(n9544), .A2(n9543), .ZN(n15456) );
  AND2_X1 U9321 ( .A1(n14728), .A2(n14305), .ZN(n7508) );
  NOR2_X1 U9322 ( .A1(n14257), .A2(n8179), .ZN(n7509) );
  NOR2_X1 U9323 ( .A1(n13324), .A2(n13325), .ZN(n7510) );
  NOR2_X1 U9324 ( .A1(n8420), .A2(n13053), .ZN(n7511) );
  AND2_X1 U9325 ( .A1(n14164), .A2(n14163), .ZN(n7512) );
  AND2_X1 U9326 ( .A1(n8186), .A2(n8182), .ZN(n7513) );
  AND2_X1 U9327 ( .A1(n9082), .A2(n12971), .ZN(n7514) );
  AND2_X1 U9328 ( .A1(n13512), .A2(n8347), .ZN(n7515) );
  NOR2_X1 U9329 ( .A1(n13380), .A2(n13731), .ZN(n7516) );
  AND2_X1 U9330 ( .A1(n7848), .A2(n9239), .ZN(n7517) );
  INV_X1 U9331 ( .A(n9754), .ZN(n8284) );
  AND2_X1 U9332 ( .A1(n14668), .A2(n7749), .ZN(n7518) );
  AND2_X1 U9333 ( .A1(n14439), .A2(n14438), .ZN(n7519) );
  INV_X1 U9334 ( .A(n9531), .ZN(n8281) );
  AND2_X1 U9335 ( .A1(n12790), .A2(n13214), .ZN(n7520) );
  NOR2_X1 U9336 ( .A1(n8029), .A2(n13229), .ZN(n7521) );
  INV_X1 U9337 ( .A(n7866), .ZN(n7865) );
  NAND2_X1 U9338 ( .A1(n8224), .A2(n9521), .ZN(n7866) );
  INV_X1 U9339 ( .A(n7996), .ZN(n14563) );
  INV_X1 U9340 ( .A(n8012), .ZN(n15170) );
  OR2_X1 U9341 ( .A1(n14071), .A2(n14070), .ZN(n7522) );
  OR2_X1 U9342 ( .A1(n7885), .A2(n10266), .ZN(n7523) );
  AND2_X1 U9343 ( .A1(n8245), .A2(n8244), .ZN(n7524) );
  AND2_X1 U9344 ( .A1(n8417), .A2(n8415), .ZN(n7525) );
  INV_X1 U9345 ( .A(n8436), .ZN(n8435) );
  AND2_X1 U9346 ( .A1(n8534), .A2(n7869), .ZN(n7526) );
  INV_X1 U9347 ( .A(n7945), .ZN(n7944) );
  NOR2_X1 U9348 ( .A1(n16572), .A2(n11938), .ZN(n7945) );
  AND2_X1 U9349 ( .A1(n14223), .A2(n14224), .ZN(n7527) );
  AND2_X1 U9350 ( .A1(n15909), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n7528) );
  INV_X1 U9351 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8523) );
  NOR2_X1 U9352 ( .A1(n14089), .A2(n14309), .ZN(n7529) );
  AND2_X1 U9353 ( .A1(n8090), .A2(n9067), .ZN(n7530) );
  AND2_X1 U9354 ( .A1(n11081), .A2(n16373), .ZN(n7531) );
  NOR2_X1 U9355 ( .A1(n12196), .A2(n12183), .ZN(n7532) );
  INV_X1 U9356 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n15692) );
  OR2_X1 U9357 ( .A1(n8122), .A2(n7836), .ZN(n7533) );
  AND2_X1 U9358 ( .A1(n12892), .A2(n11924), .ZN(n7534) );
  NOR2_X1 U9359 ( .A1(n15451), .A2(n15303), .ZN(n7535) );
  OR2_X1 U9360 ( .A1(n16327), .A2(n13362), .ZN(n7536) );
  NOR2_X1 U9361 ( .A1(n14728), .A2(n12452), .ZN(n7537) );
  NOR2_X1 U9362 ( .A1(n15470), .A2(n12312), .ZN(n7538) );
  INV_X1 U9363 ( .A(n13413), .ZN(n8074) );
  INV_X1 U9364 ( .A(n7924), .ZN(n7923) );
  NAND2_X1 U9365 ( .A1(n7925), .A2(n12745), .ZN(n7924) );
  XNOR2_X1 U9366 ( .A(n15382), .B(n15147), .ZN(n15130) );
  INV_X1 U9367 ( .A(n7826), .ZN(n7825) );
  NAND2_X1 U9368 ( .A1(n11667), .A2(n7494), .ZN(n7826) );
  AND2_X1 U9369 ( .A1(n8315), .A2(n8314), .ZN(n7540) );
  INV_X1 U9370 ( .A(n8445), .ZN(n8444) );
  NOR2_X1 U9371 ( .A1(n15180), .A2(n8451), .ZN(n8445) );
  INV_X1 U9372 ( .A(n11144), .ZN(n8112) );
  AND2_X1 U9373 ( .A1(n8468), .A2(n8462), .ZN(n7541) );
  INV_X1 U9374 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9361) );
  OR2_X1 U9375 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n7542) );
  INV_X1 U9376 ( .A(n8451), .ZN(n8450) );
  NOR2_X1 U9377 ( .A1(n15206), .A2(n7885), .ZN(n8451) );
  OR2_X1 U9378 ( .A1(n8866), .A2(P3_IR_REG_18__SCAN_IN), .ZN(n7543) );
  OR2_X1 U9379 ( .A1(n15248), .A2(n8341), .ZN(n7544) );
  AND2_X1 U9380 ( .A1(n12086), .A2(n12085), .ZN(n7545) );
  AND2_X1 U9381 ( .A1(n11895), .A2(n11894), .ZN(n7546) );
  AND2_X1 U9382 ( .A1(n10977), .A2(n10976), .ZN(n7547) );
  AND2_X1 U9383 ( .A1(n14129), .A2(n14128), .ZN(n7548) );
  AND2_X1 U9384 ( .A1(n9202), .A2(SI_9_), .ZN(n7549) );
  NOR2_X1 U9385 ( .A1(n14593), .A2(n14615), .ZN(n7550) );
  NOR2_X1 U9386 ( .A1(n14068), .A2(n11682), .ZN(n7551) );
  OR2_X1 U9387 ( .A1(n15363), .A2(n16544), .ZN(n7552) );
  INV_X1 U9388 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10225) );
  INV_X1 U9389 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10229) );
  INV_X1 U9390 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10179) );
  INV_X1 U9391 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9120) );
  NOR2_X1 U9392 ( .A1(n8326), .A2(n15307), .ZN(n7553) );
  AND2_X1 U9393 ( .A1(n10215), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7554) );
  OR2_X1 U9394 ( .A1(n8487), .A2(n14140), .ZN(n7555) );
  AND2_X1 U9395 ( .A1(n12321), .A2(n12323), .ZN(n7556) );
  INV_X1 U9396 ( .A(n8478), .ZN(n8477) );
  NOR2_X1 U9397 ( .A1(n8479), .A2(n15252), .ZN(n8478) );
  INV_X1 U9398 ( .A(n8158), .ZN(n8157) );
  NAND2_X1 U9399 ( .A1(n8161), .A2(n13939), .ZN(n8158) );
  AND2_X1 U9400 ( .A1(n8571), .A2(n7612), .ZN(n7557) );
  NAND2_X1 U9401 ( .A1(n13179), .A2(n13207), .ZN(n7558) );
  AND2_X1 U9402 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7559) );
  NAND2_X1 U9403 ( .A1(n15130), .A2(n8473), .ZN(n8468) );
  NAND2_X1 U9404 ( .A1(n8104), .A2(n12060), .ZN(n7560) );
  OR2_X1 U9405 ( .A1(n16016), .A2(n16017), .ZN(n7561) );
  OR2_X1 U9406 ( .A1(n7548), .A2(n14131), .ZN(n7562) );
  OR2_X1 U9407 ( .A1(n9414), .A2(n9416), .ZN(n7563) );
  OR2_X1 U9408 ( .A1(n14142), .A2(n14139), .ZN(n7564) );
  AND2_X1 U9409 ( .A1(n12946), .A2(n12944), .ZN(n13535) );
  INV_X1 U9410 ( .A(n13535), .ZN(n8349) );
  AND2_X1 U9411 ( .A1(n11035), .A2(n11258), .ZN(n7565) );
  INV_X1 U9412 ( .A(n13575), .ZN(n13580) );
  AND2_X1 U9413 ( .A1(n7951), .A2(n7489), .ZN(n7566) );
  NOR2_X1 U9414 ( .A1(n12244), .A2(n9074), .ZN(n7567) );
  AND2_X1 U9415 ( .A1(n7808), .A2(n7806), .ZN(n7568) );
  NOR2_X1 U9416 ( .A1(n13971), .A2(n13840), .ZN(n7569) );
  NOR2_X1 U9417 ( .A1(n14473), .A2(n8300), .ZN(n8299) );
  INV_X1 U9418 ( .A(n8912), .ZN(n8096) );
  AND2_X1 U9419 ( .A1(n8090), .A2(n8089), .ZN(n7570) );
  AND2_X1 U9420 ( .A1(n14301), .A2(n14302), .ZN(n7571) );
  AND2_X1 U9421 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), .ZN(
        n7572) );
  NOR2_X1 U9422 ( .A1(n12941), .A2(n8351), .ZN(n8350) );
  OR2_X1 U9423 ( .A1(n14177), .A2(n14178), .ZN(n7573) );
  OR2_X1 U9424 ( .A1(n14118), .A2(n8507), .ZN(n7574) );
  AND2_X1 U9425 ( .A1(n7552), .A2(n8335), .ZN(n7575) );
  OR2_X1 U9426 ( .A1(n8490), .A2(n8492), .ZN(n7576) );
  OR2_X1 U9427 ( .A1(n8281), .A2(n9530), .ZN(n7577) );
  OR2_X1 U9428 ( .A1(n9567), .A2(n9565), .ZN(n7578) );
  OR2_X1 U9429 ( .A1(n8284), .A2(n9753), .ZN(n7579) );
  OR2_X1 U9430 ( .A1(n8495), .A2(n14048), .ZN(n7580) );
  OR2_X1 U9431 ( .A1(n8499), .A2(n14064), .ZN(n7581) );
  OR2_X1 U9432 ( .A1(n9604), .A2(n9602), .ZN(n7582) );
  OR2_X1 U9433 ( .A1(n9493), .A2(n9491), .ZN(n7583) );
  OR2_X1 U9434 ( .A1(n9451), .A2(n8275), .ZN(n7584) );
  OR2_X1 U9435 ( .A1(n8278), .A2(n9647), .ZN(n7585) );
  NAND2_X1 U9436 ( .A1(n12710), .A2(n12704), .ZN(n7586) );
  AND2_X1 U9437 ( .A1(n14025), .A2(n14024), .ZN(n7587) );
  AND2_X1 U9438 ( .A1(n7499), .A2(n8535), .ZN(n7588) );
  NAND2_X1 U9439 ( .A1(n14085), .A2(n14086), .ZN(n7589) );
  NAND2_X1 U9440 ( .A1(n12599), .A2(n8130), .ZN(n7590) );
  INV_X1 U9441 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9154) );
  OR2_X1 U9442 ( .A1(n8554), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n7591) );
  OR2_X1 U9443 ( .A1(n8489), .A2(n7512), .ZN(n7592) );
  INV_X1 U9444 ( .A(n7933), .ZN(n7932) );
  NAND2_X1 U9445 ( .A1(n14631), .A2(n7934), .ZN(n7933) );
  INV_X1 U9446 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8534) );
  INV_X1 U9447 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7703) );
  INV_X1 U9448 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7869) );
  INV_X1 U9449 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8166) );
  NAND2_X1 U9450 ( .A1(n13770), .A2(n13769), .ZN(n14693) );
  INV_X1 U9451 ( .A(n14693), .ZN(n7995) );
  NAND2_X1 U9452 ( .A1(n12258), .A2(n12257), .ZN(n12382) );
  NAND2_X1 U9453 ( .A1(n11896), .A2(n12722), .ZN(n12728) );
  NAND2_X1 U9454 ( .A1(n13486), .A2(n13499), .ZN(n7594) );
  INV_X1 U9455 ( .A(n13801), .ZN(n7920) );
  AND2_X1 U9456 ( .A1(n12343), .A2(n8008), .ZN(n7595) );
  AND2_X1 U9457 ( .A1(n14437), .A2(n7458), .ZN(n7596) );
  INV_X1 U9458 ( .A(n14939), .ZN(n15133) );
  AND4_X1 U9459 ( .A1(n9171), .A2(n9170), .A3(n9169), .A4(n9168), .ZN(n14939)
         );
  AND2_X1 U9460 ( .A1(n8345), .A2(n8347), .ZN(n7597) );
  OR2_X1 U9461 ( .A1(n13726), .A2(n13213), .ZN(n12929) );
  INV_X1 U9462 ( .A(n12929), .ZN(n8407) );
  AND2_X1 U9463 ( .A1(n7889), .A2(n8327), .ZN(n7598) );
  AND2_X1 U9464 ( .A1(n7943), .A2(n7942), .ZN(n7599) );
  INV_X1 U9465 ( .A(n11837), .ZN(n7768) );
  NOR2_X1 U9466 ( .A1(n7990), .A2(n14785), .ZN(n7600) );
  NAND2_X1 U9467 ( .A1(n12294), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7601) );
  NOR2_X1 U9468 ( .A1(n12295), .A2(n12296), .ZN(n7779) );
  INV_X1 U9469 ( .A(n8784), .ZN(n8070) );
  AND2_X1 U9470 ( .A1(n8803), .A2(n8783), .ZN(n8784) );
  INV_X2 U9471 ( .A(n14571), .ZN(n14644) );
  NAND2_X1 U9472 ( .A1(n12425), .A2(n12424), .ZN(n14426) );
  INV_X1 U9473 ( .A(n14426), .ZN(n7992) );
  INV_X1 U9474 ( .A(n13234), .ZN(n8029) );
  INV_X1 U9475 ( .A(n15307), .ZN(n8430) );
  NAND2_X1 U9476 ( .A1(n9646), .A2(n9645), .ZN(n15257) );
  INV_X1 U9477 ( .A(n15257), .ZN(n8482) );
  NAND2_X1 U9478 ( .A1(n9269), .A2(n9934), .ZN(n11549) );
  INV_X1 U9479 ( .A(n11549), .ZN(n8291) );
  INV_X1 U9480 ( .A(n14267), .ZN(n7939) );
  AND2_X1 U9481 ( .A1(n11344), .A2(n11345), .ZN(n7602) );
  NOR2_X1 U9482 ( .A1(n11949), .A2(n14089), .ZN(n7740) );
  XOR2_X1 U9483 ( .A(n11346), .B(n11338), .Z(n7603) );
  INV_X1 U9484 ( .A(n11943), .ZN(n8178) );
  AND2_X2 U9485 ( .A1(n9145), .A2(n10603), .ZN(n16569) );
  NAND2_X1 U9486 ( .A1(n9054), .A2(n8353), .ZN(n7604) );
  AND2_X1 U9487 ( .A1(n13316), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7605) );
  AND2_X1 U9488 ( .A1(n11421), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7606) );
  OR2_X1 U9489 ( .A1(n16566), .A2(n13582), .ZN(n7607) );
  AND2_X1 U9490 ( .A1(n8114), .A2(n11144), .ZN(n7608) );
  INV_X1 U9491 ( .A(n11421), .ZN(n8253) );
  AND2_X1 U9492 ( .A1(n8114), .A2(n8111), .ZN(n7609) );
  INV_X1 U9493 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7840) );
  INV_X1 U9494 ( .A(n8367), .ZN(n8366) );
  AOI21_X1 U9495 ( .B1(n12120), .B2(n8368), .A(n7556), .ZN(n8367) );
  AND2_X1 U9496 ( .A1(n8365), .A2(n8367), .ZN(n7610) );
  NOR2_X1 U9497 ( .A1(n11993), .A2(n16539), .ZN(n7782) );
  INV_X1 U9498 ( .A(n8215), .ZN(n8214) );
  NAND2_X1 U9499 ( .A1(n9792), .A2(n8216), .ZN(n8215) );
  INV_X1 U9500 ( .A(n8139), .ZN(n10128) );
  INV_X1 U9501 ( .A(n11756), .ZN(n8004) );
  INV_X1 U9502 ( .A(n14321), .ZN(n7948) );
  NAND2_X1 U9503 ( .A1(n10604), .A2(n10603), .ZN(n13204) );
  INV_X1 U9504 ( .A(n13204), .ZN(n13183) );
  INV_X1 U9505 ( .A(n15431), .ZN(n16449) );
  NAND2_X1 U9506 ( .A1(n9969), .A2(n9968), .ZN(n15431) );
  AND2_X1 U9507 ( .A1(n8000), .A2(n16446), .ZN(n7611) );
  INV_X1 U9508 ( .A(n11283), .ZN(n8238) );
  INV_X1 U9509 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7732) );
  INV_X1 U9510 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7979) );
  INV_X1 U9511 ( .A(n13292), .ZN(n7871) );
  XNOR2_X1 U9512 ( .A(n13276), .B(n13292), .ZN(n13258) );
  INV_X1 U9513 ( .A(n10125), .ZN(n14287) );
  NAND2_X1 U9514 ( .A1(n7557), .A2(n8572), .ZN(n10691) );
  AOI22_X2 U9515 ( .A1(n11932), .A2(n11931), .B1(n11930), .B2(n13221), .ZN(
        n12121) );
  OAI21_X1 U9516 ( .B1(n13097), .B2(n13095), .A(n13093), .ZN(n12810) );
  NOR2_X1 U9517 ( .A1(n10601), .A2(n8344), .ZN(n10715) );
  INV_X1 U9518 ( .A(n10591), .ZN(n10597) );
  NAND2_X1 U9519 ( .A1(n8365), .A2(n8363), .ZN(n12480) );
  NAND2_X1 U9520 ( .A1(n13128), .A2(n13127), .ZN(n13126) );
  NAND2_X1 U9521 ( .A1(n13088), .A2(n13087), .ZN(n13086) );
  NAND2_X1 U9522 ( .A1(n11696), .A2(n11695), .ZN(n11880) );
  XNOR2_X1 U9523 ( .A(n16368), .B(n12834), .ZN(n10599) );
  NAND2_X2 U9524 ( .A1(n13181), .A2(n13182), .ZN(n13180) );
  NAND2_X1 U9525 ( .A1(n13174), .A2(n13173), .ZN(n13172) );
  NAND2_X1 U9526 ( .A1(n13145), .A2(n13144), .ZN(n13143) );
  NAND2_X1 U9527 ( .A1(n13121), .A2(n13120), .ZN(n13119) );
  NOR2_X1 U9528 ( .A1(n10716), .A2(n10717), .ZN(n11080) );
  OAI21_X2 U9529 ( .B1(n15250), .B2(n7544), .A(n8339), .ZN(n7884) );
  INV_X1 U9530 ( .A(n15160), .ZN(n7627) );
  NAND2_X1 U9531 ( .A1(n15368), .A2(n15431), .ZN(n7628) );
  NAND2_X1 U9532 ( .A1(n10523), .A2(n10524), .ZN(n10856) );
  NAND2_X1 U9533 ( .A1(n11758), .A2(n11757), .ZN(n11821) );
  NAND2_X1 U9534 ( .A1(n11856), .A2(n11855), .ZN(n12152) );
  NAND4_X1 U9535 ( .A1(n15072), .A2(n8195), .A3(n8194), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n8193) );
  NAND3_X1 U9536 ( .A1(n14173), .A2(n7479), .A3(n7576), .ZN(n7626) );
  NAND2_X1 U9537 ( .A1(n7636), .A2(n7635), .ZN(n7634) );
  NAND2_X1 U9538 ( .A1(n7970), .A2(n14243), .ZN(n8208) );
  NAND2_X1 U9539 ( .A1(n14289), .A2(n7667), .ZN(n7624) );
  NOR2_X1 U9540 ( .A1(n14056), .A2(n8500), .ZN(n8497) );
  OAI211_X1 U9541 ( .C1(n14162), .C2(n14161), .A(n14160), .B(n7592), .ZN(n7680) );
  NAND2_X1 U9542 ( .A1(n8033), .A2(n7622), .ZN(n8929) );
  NAND3_X1 U9543 ( .A1(n7624), .A2(n14303), .A3(n7571), .ZN(P2_U3328) );
  NAND3_X1 U9544 ( .A1(n7539), .A2(n7473), .A3(n7625), .ZN(n8494) );
  NAND2_X1 U9545 ( .A1(n7626), .A2(n7573), .ZN(n8491) );
  INV_X1 U9546 ( .A(n13988), .ZN(n7720) );
  NAND2_X1 U9547 ( .A1(n13984), .A2(n13985), .ZN(n13988) );
  AND2_X1 U9548 ( .A1(n7714), .A2(n7711), .ZN(n13067) );
  INV_X1 U9549 ( .A(n13006), .ZN(n13670) );
  NAND2_X1 U9550 ( .A1(n9026), .A2(n9025), .ZN(n9039) );
  NAND2_X1 U9551 ( .A1(n8600), .A2(n8599), .ZN(n8618) );
  NAND2_X1 U9552 ( .A1(n8620), .A2(n8619), .ZN(n8623) );
  NAND2_X1 U9553 ( .A1(n14016), .A2(n14015), .ZN(n14022) );
  OAI22_X1 U9554 ( .A1(n14112), .A2(n7973), .B1(n14119), .B2(n8506), .ZN(
        n14125) );
  INV_X1 U9555 ( .A(n9351), .ZN(n9283) );
  NOR2_X1 U9556 ( .A1(n7701), .A2(n7700), .ZN(n7699) );
  XNOR2_X1 U9557 ( .A(n8337), .B(n8336), .ZN(n15368) );
  NAND3_X1 U9558 ( .A1(n15369), .A2(n7628), .A3(n7575), .ZN(n15481) );
  OAI21_X1 U9559 ( .B1(n15091), .B2(n15090), .A(n15089), .ZN(n8337) );
  NAND2_X1 U9560 ( .A1(n12560), .A2(n12559), .ZN(n15250) );
  NAND2_X1 U9561 ( .A1(n7884), .A2(n7879), .ZN(n12565) );
  NAND2_X1 U9562 ( .A1(n15181), .A2(n15180), .ZN(n15179) );
  INV_X1 U9563 ( .A(n10861), .ZN(n7878) );
  NAND2_X1 U9564 ( .A1(n12793), .A2(n13192), .ZN(n13121) );
  NAND2_X1 U9565 ( .A1(n11880), .A2(n11879), .ZN(n11932) );
  NAND4_X1 U9566 ( .A1(n9149), .A2(n9147), .A3(n9150), .A4(n9148), .ZN(n9559)
         );
  NAND3_X1 U9567 ( .A1(n9888), .A2(n9887), .A3(n7630), .ZN(n7629) );
  NAND2_X1 U9568 ( .A1(n8346), .A2(n8350), .ZN(n8345) );
  NAND2_X1 U9569 ( .A1(n13511), .A2(n12953), .ZN(n13495) );
  NAND2_X1 U9570 ( .A1(n8286), .A2(n7507), .ZN(n7751) );
  NAND2_X1 U9571 ( .A1(n13493), .A2(n12853), .ZN(n13483) );
  NAND2_X1 U9572 ( .A1(n13448), .A2(n13447), .ZN(n9082) );
  NAND2_X1 U9573 ( .A1(n9076), .A2(n12925), .ZN(n12463) );
  OAI21_X1 U9574 ( .B1(n11977), .B2(n8404), .A(n8401), .ZN(n12472) );
  NOR2_X1 U9575 ( .A1(n13058), .A2(n7715), .ZN(n7714) );
  INV_X1 U9576 ( .A(n9304), .ZN(n9842) );
  NAND2_X2 U9577 ( .A1(n9327), .A2(n7506), .ZN(n14973) );
  XNOR2_X1 U9578 ( .A(n9312), .B(P1_IR_REG_2__SCAN_IN), .ZN(n10461) );
  NOR2_X2 U9579 ( .A1(n7974), .A2(n16302), .ZN(n16308) );
  INV_X1 U9580 ( .A(n7727), .ZN(n16007) );
  NAND2_X1 U9581 ( .A1(n8375), .A2(n8374), .ZN(n13193) );
  INV_X1 U9582 ( .A(n11332), .ZN(n7987) );
  NAND2_X1 U9583 ( .A1(n16418), .A2(n11333), .ZN(n11332) );
  NAND2_X1 U9584 ( .A1(n14666), .A2(n7689), .ZN(n14754) );
  OAI21_X1 U9585 ( .B1(n14735), .B2(n14667), .A(n14665), .ZN(n7690) );
  NAND2_X1 U9586 ( .A1(n7639), .A2(n7638), .ZN(n7637) );
  NAND2_X1 U9587 ( .A1(n7637), .A2(n7634), .ZN(n14111) );
  NAND2_X1 U9588 ( .A1(n14105), .A2(n14104), .ZN(n7639) );
  NOR2_X2 U9589 ( .A1(n15985), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n15984) );
  NAND2_X1 U9590 ( .A1(n16293), .A2(n16294), .ZN(n16292) );
  AND2_X2 U9591 ( .A1(n7641), .A2(n7640), .ZN(n16005) );
  INV_X1 U9592 ( .A(n16321), .ZN(n7641) );
  OAI21_X1 U9593 ( .B1(n16285), .B2(n16284), .A(n7476), .ZN(n7727) );
  NAND2_X1 U9594 ( .A1(n16023), .A2(n16024), .ZN(n7725) );
  NOR2_X2 U9595 ( .A1(n7735), .A2(n7734), .ZN(n16314) );
  AOI21_X1 U9596 ( .B1(n16304), .B2(n16303), .A(P2_ADDR_REG_13__SCAN_IN), .ZN(
        n7974) );
  NAND2_X1 U9597 ( .A1(n7975), .A2(n16292), .ZN(n16298) );
  INV_X1 U9598 ( .A(n7697), .ZN(n16304) );
  AOI21_X2 U9599 ( .B1(n16198), .B2(n16020), .A(n16306), .ZN(n16311) );
  NAND2_X1 U9600 ( .A1(n7725), .A2(n7726), .ZN(n7735) );
  NAND2_X1 U9601 ( .A1(n7645), .A2(n16255), .ZN(n7976) );
  NAND2_X1 U9602 ( .A1(n16290), .A2(n16289), .ZN(n7645) );
  NOR2_X1 U9603 ( .A1(n16311), .A2(n16312), .ZN(n16310) );
  OAI21_X1 U9604 ( .B1(n16301), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7561), .ZN(
        n7697) );
  INV_X4 U9605 ( .A(n10266), .ZN(n7883) );
  NAND2_X2 U9606 ( .A1(n13882), .A2(n7646), .ZN(n13881) );
  NAND2_X2 U9607 ( .A1(n8146), .A2(n8144), .ZN(n13882) );
  NAND2_X1 U9608 ( .A1(n13982), .A2(n14366), .ZN(n8137) );
  NAND2_X1 U9609 ( .A1(n7478), .A2(n7564), .ZN(n7649) );
  INV_X1 U9610 ( .A(n10028), .ZN(n8164) );
  NAND2_X1 U9611 ( .A1(n7680), .A2(n8488), .ZN(n14172) );
  AND4_X2 U9612 ( .A1(n10087), .A2(n10012), .A3(n10011), .A4(n10010), .ZN(
        n7669) );
  AOI21_X1 U9613 ( .B1(n14147), .B2(n14146), .A(n14145), .ZN(n14149) );
  NAND2_X1 U9614 ( .A1(n7651), .A2(n7650), .ZN(n14023) );
  NAND3_X1 U9615 ( .A1(n7671), .A2(n14023), .A3(n8503), .ZN(n8502) );
  NOR2_X1 U9616 ( .A1(n7654), .A2(n7653), .ZN(n7652) );
  NAND2_X1 U9617 ( .A1(n14099), .A2(n14098), .ZN(n14105) );
  NAND2_X1 U9618 ( .A1(n7720), .A2(n14004), .ZN(n13991) );
  NAND2_X1 U9619 ( .A1(n14436), .A2(n14435), .ZN(n14541) );
  OR2_X1 U9620 ( .A1(n14670), .A2(n14735), .ZN(n7749) );
  NAND3_X2 U9621 ( .A1(n7949), .A2(n10021), .A3(n10022), .ZN(n14321) );
  NAND2_X1 U9622 ( .A1(n8197), .A2(n8198), .ZN(n9462) );
  NAND2_X1 U9623 ( .A1(n7926), .A2(n10799), .ZN(n10817) );
  INV_X1 U9624 ( .A(n14247), .ZN(n10120) );
  NAND2_X1 U9625 ( .A1(n10797), .A2(n10796), .ZN(n10832) );
  OAI21_X1 U9626 ( .B1(n9487), .B2(n8227), .A(n8224), .ZN(n9522) );
  NAND2_X1 U9627 ( .A1(n7751), .A2(n9375), .ZN(n9376) );
  NAND2_X1 U9628 ( .A1(n7709), .A2(n7708), .ZN(n9302) );
  NAND2_X4 U9629 ( .A1(n15909), .A2(n9164), .ZN(n9843) );
  NAND3_X1 U9630 ( .A1(n7665), .A2(n9336), .A3(n9337), .ZN(n9342) );
  NAND3_X1 U9631 ( .A1(n9318), .A2(n9317), .A3(n10524), .ZN(n7665) );
  INV_X1 U9632 ( .A(n7666), .ZN(n9433) );
  NAND2_X1 U9633 ( .A1(n7684), .A2(n13227), .ZN(n10600) );
  NAND4_X1 U9634 ( .A1(n10035), .A2(n10036), .A3(n10037), .A4(n10038), .ZN(
        n13984) );
  NAND2_X1 U9635 ( .A1(n7969), .A2(n8304), .ZN(n10016) );
  NAND2_X1 U9636 ( .A1(n14022), .A2(n14021), .ZN(n7673) );
  NAND2_X1 U9637 ( .A1(n7673), .A2(n7672), .ZN(n7671) );
  AND3_X2 U9638 ( .A1(n7670), .A2(n7669), .A3(n7668), .ZN(n10013) );
  AND2_X1 U9639 ( .A1(n10007), .A2(n10006), .ZN(n7668) );
  NAND2_X1 U9640 ( .A1(n13997), .A2(n13993), .ZN(n7679) );
  NAND2_X1 U9641 ( .A1(n14127), .A2(n7562), .ZN(n7674) );
  NAND2_X1 U9642 ( .A1(n7678), .A2(n7677), .ZN(n14072) );
  INV_X1 U9643 ( .A(n10599), .ZN(n7684) );
  XNOR2_X1 U9644 ( .A(n9173), .B(SI_1_), .ZN(n9282) );
  INV_X1 U9645 ( .A(n9282), .ZN(n9177) );
  NAND4_X1 U9646 ( .A1(n8548), .A2(n8192), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n8191) );
  NAND2_X1 U9647 ( .A1(n9795), .A2(n9794), .ZN(n7675) );
  MUX2_X2 U9648 ( .A(n9813), .B(n15081), .S(n9837), .Z(n9861) );
  NAND2_X1 U9649 ( .A1(n9255), .A2(n8236), .ZN(n8235) );
  NAND2_X1 U9650 ( .A1(n9678), .A2(n9244), .ZN(n9247) );
  NOR2_X1 U9651 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n10007) );
  NAND2_X1 U9652 ( .A1(n14071), .A2(n14070), .ZN(n7678) );
  NAND2_X1 U9653 ( .A1(n7679), .A2(n13996), .ZN(n14003) );
  NAND2_X1 U9654 ( .A1(n14041), .A2(n14040), .ZN(n7682) );
  NAND2_X1 U9655 ( .A1(n9054), .A2(n8354), .ZN(n9095) );
  NAND2_X1 U9656 ( .A1(n7685), .A2(n12840), .ZN(P3_U3160) );
  NAND3_X1 U9657 ( .A1(n7686), .A2(n7687), .A3(n8379), .ZN(n7685) );
  INV_X1 U9658 ( .A(n9054), .ZN(n9056) );
  NAND2_X1 U9659 ( .A1(n7718), .A2(n8386), .ZN(n11696) );
  NAND2_X1 U9660 ( .A1(n7688), .A2(n9373), .ZN(n9377) );
  NAND3_X1 U9661 ( .A1(n8286), .A2(n7507), .A3(n9374), .ZN(n7688) );
  NAND2_X1 U9662 ( .A1(n10820), .A2(n14255), .ZN(n10822) );
  NAND2_X1 U9663 ( .A1(n11244), .A2(n11243), .ZN(n11501) );
  OAI21_X1 U9664 ( .B1(n12136), .B2(n14102), .A(n12135), .ZN(n12138) );
  OAI21_X2 U9665 ( .B1(n14609), .B2(n14389), .A(n14391), .ZN(n14588) );
  OAI21_X1 U9666 ( .B1(n14543), .B2(n14401), .A(n14403), .ZN(n14527) );
  NAND2_X1 U9667 ( .A1(n14249), .A2(n11320), .ZN(n11319) );
  NAND2_X1 U9668 ( .A1(n8174), .A2(n8175), .ZN(n12136) );
  NAND2_X1 U9669 ( .A1(n11781), .A2(n11780), .ZN(n11782) );
  NAND2_X1 U9670 ( .A1(n13180), .A2(n7503), .ZN(n13184) );
  MUX2_X2 U9671 ( .A(n14657), .B(n14746), .S(n14740), .Z(n14658) );
  NAND2_X1 U9672 ( .A1(n8303), .A2(n8304), .ZN(n10028) );
  NAND2_X1 U9673 ( .A1(n7692), .A2(n7691), .ZN(n10828) );
  INV_X1 U9674 ( .A(n14038), .ZN(n7691) );
  NOR2_X1 U9675 ( .A1(n16103), .A2(n16104), .ZN(n16102) );
  OR2_X1 U9676 ( .A1(n13371), .A2(n16328), .ZN(n7873) );
  NAND2_X1 U9677 ( .A1(n10957), .A2(n10956), .ZN(n10958) );
  INV_X1 U9678 ( .A(n7735), .ZN(n16027) );
  NOR2_X1 U9679 ( .A1(n7761), .A2(n11038), .ZN(n7759) );
  INV_X1 U9680 ( .A(n11217), .ZN(n7753) );
  OAI211_X1 U9681 ( .C1(n8477), .C2(n8475), .A(n8474), .B(n8476), .ZN(n15238)
         );
  NAND2_X2 U9682 ( .A1(n7702), .A2(n7699), .ZN(n15912) );
  OR2_X1 U9683 ( .A1(n10642), .A2(n9332), .ZN(n10855) );
  NAND2_X1 U9684 ( .A1(n8933), .A2(n8932), .ZN(n8947) );
  NOR2_X1 U9685 ( .A1(n12970), .A2(n12967), .ZN(n12972) );
  NAND2_X1 U9686 ( .A1(n8075), .A2(n8071), .ZN(n12981) );
  NAND2_X1 U9687 ( .A1(n8976), .A2(n8975), .ZN(n8979) );
  XNOR2_X1 U9688 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8562) );
  INV_X1 U9689 ( .A(n7712), .ZN(n7711) );
  OAI21_X1 U9690 ( .B1(n13059), .B2(n13046), .A(n7713), .ZN(n7712) );
  NAND2_X1 U9691 ( .A1(n13059), .A2(n13060), .ZN(n7713) );
  NAND2_X1 U9692 ( .A1(n15197), .A2(n15402), .ZN(n15171) );
  NAND2_X1 U9693 ( .A1(n11864), .A2(n16521), .ZN(n11865) );
  NOR2_X2 U9694 ( .A1(n15254), .A2(n15421), .ZN(n15240) );
  NAND2_X1 U9695 ( .A1(n12569), .A2(n15431), .ZN(n12571) );
  NAND2_X1 U9696 ( .A1(n7842), .A2(n9190), .ZN(n9385) );
  XNOR2_X1 U9697 ( .A(n9409), .B(n9408), .ZN(n10723) );
  NAND3_X1 U9698 ( .A1(n15375), .A2(n15373), .A3(n15374), .ZN(n15482) );
  NOR2_X2 U9699 ( .A1(n9559), .A2(n9151), .ZN(n9152) );
  NAND2_X1 U9700 ( .A1(n9342), .A2(n8285), .ZN(n8286) );
  NAND2_X1 U9701 ( .A1(n9102), .A2(n7572), .ZN(n7867) );
  XNOR2_X1 U9702 ( .A(n13072), .B(n13073), .ZN(n13074) );
  NAND2_X1 U9703 ( .A1(n13126), .A2(n12798), .ZN(n13174) );
  NOR2_X1 U9704 ( .A1(n10715), .A2(n10714), .ZN(n10716) );
  NAND2_X1 U9705 ( .A1(n13172), .A2(n12800), .ZN(n13088) );
  INV_X1 U9706 ( .A(n8639), .ZN(n7787) );
  NAND2_X1 U9707 ( .A1(n11083), .A2(n8388), .ZN(n7718) );
  NAND2_X1 U9708 ( .A1(n9104), .A2(n9103), .ZN(n9106) );
  INV_X1 U9709 ( .A(n9303), .ZN(n9290) );
  NAND2_X1 U9710 ( .A1(n9290), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9292) );
  NAND3_X1 U9711 ( .A1(n7955), .A2(n7957), .A3(n7589), .ZN(n7954) );
  OAI21_X1 U9712 ( .B1(n14111), .B2(n14110), .A(n7574), .ZN(n7973) );
  NAND2_X1 U9713 ( .A1(n8494), .A2(n7580), .ZN(n14055) );
  NAND2_X1 U9714 ( .A1(n8491), .A2(n8520), .ZN(n7971) );
  NAND2_X1 U9715 ( .A1(n7958), .A2(n14081), .ZN(n7957) );
  NAND2_X1 U9716 ( .A1(n7971), .A2(n8209), .ZN(n7970) );
  INV_X1 U9717 ( .A(n8208), .ZN(n14289) );
  NAND2_X1 U9718 ( .A1(n7954), .A2(n8484), .ZN(n14094) );
  OAI21_X1 U9719 ( .B1(n14154), .B2(n7968), .A(n7965), .ZN(n14162) );
  NAND2_X1 U9720 ( .A1(n8169), .A2(n8168), .ZN(n14385) );
  INV_X1 U9721 ( .A(n8304), .ZN(n10628) );
  INV_X1 U9722 ( .A(n10019), .ZN(n14800) );
  XNOR2_X1 U9723 ( .A(n7845), .B(n8313), .ZN(n14418) );
  NAND2_X1 U9724 ( .A1(n12219), .A2(n12218), .ZN(n12220) );
  INV_X1 U9725 ( .A(n14454), .ZN(n7722) );
  INV_X2 U9726 ( .A(n9338), .ZN(n9372) );
  MUX2_X1 U9727 ( .A(n10851), .B(n10915), .S(n9338), .Z(n9357) );
  NOR2_X4 U9728 ( .A1(n9574), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n8288) );
  NAND2_X1 U9729 ( .A1(n7722), .A2(n7847), .ZN(n14456) );
  NAND2_X1 U9730 ( .A1(n14453), .A2(n14452), .ZN(n7847) );
  OAI21_X1 U9731 ( .B1(n10029), .B2(n10229), .A(n7724), .ZN(n9178) );
  NAND2_X1 U9732 ( .A1(n14669), .A2(n7518), .ZN(n14755) );
  INV_X1 U9733 ( .A(n14261), .ZN(n8186) );
  XNOR2_X1 U9734 ( .A(n15925), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n15988) );
  NAND2_X2 U9735 ( .A1(n7980), .A2(n15929), .ZN(n15930) );
  INV_X1 U9736 ( .A(n16310), .ZN(n7726) );
  NOR2_X4 U9737 ( .A1(n9058), .A2(n8533), .ZN(n9099) );
  AOI21_X1 U9738 ( .B1(n11284), .B2(n10969), .A(n8238), .ZN(n8242) );
  NOR2_X1 U9739 ( .A1(n13317), .A2(n13553), .ZN(n13329) );
  NAND2_X1 U9740 ( .A1(n7763), .A2(n11401), .ZN(n11014) );
  NOR2_X1 U9741 ( .A1(n12200), .A2(n12199), .ZN(n12282) );
  CLKBUF_X3 U9742 ( .A(n8553), .Z(n8415) );
  NAND2_X1 U9743 ( .A1(n14388), .A2(n14387), .ZN(n14609) );
  NAND2_X1 U9744 ( .A1(n7847), .A2(n7846), .ZN(n7845) );
  NAND2_X1 U9745 ( .A1(n9319), .A2(n9180), .ZN(n9183) );
  INV_X1 U9746 ( .A(n14527), .ZN(n7730) );
  NOR2_X1 U9747 ( .A1(n16314), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n7733) );
  NAND2_X1 U9748 ( .A1(n15933), .A2(n15932), .ZN(n15978) );
  NAND2_X1 U9749 ( .A1(n15991), .A2(n15992), .ZN(n7980) );
  INV_X1 U9750 ( .A(n16281), .ZN(n7746) );
  INV_X1 U9751 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15985) );
  NAND2_X1 U9752 ( .A1(n7978), .A2(n15997), .ZN(n15999) );
  INV_X1 U9753 ( .A(n16288), .ZN(n7977) );
  NAND3_X2 U9754 ( .A1(n12757), .A2(n12762), .A3(n10726), .ZN(n12767) );
  NAND2_X1 U9755 ( .A1(n13776), .A2(n13775), .ZN(n13921) );
  NAND2_X1 U9756 ( .A1(n10770), .A2(n10155), .ZN(n10159) );
  AOI21_X2 U9757 ( .B1(n7905), .B2(n7904), .A(n7902), .ZN(n11350) );
  INV_X1 U9758 ( .A(n10664), .ZN(n7918) );
  NAND2_X1 U9759 ( .A1(n8032), .A2(n8031), .ZN(n8976) );
  NAND2_X1 U9760 ( .A1(n8929), .A2(n8928), .ZN(n8933) );
  NAND2_X1 U9761 ( .A1(n7993), .A2(n7992), .ZN(n14620) );
  NAND2_X1 U9762 ( .A1(n12232), .A2(n12235), .ZN(n14647) );
  NAND2_X1 U9763 ( .A1(n14419), .A2(n14753), .ZN(n14378) );
  INV_X1 U9764 ( .A(n7994), .ZN(n14532) );
  NAND2_X1 U9765 ( .A1(n14748), .A2(n7738), .ZN(P2_U3498) );
  NAND2_X1 U9766 ( .A1(n7743), .A2(n7741), .ZN(P3_U3154) );
  NAND2_X1 U9767 ( .A1(n13074), .A2(n13183), .ZN(n7743) );
  XNOR2_X1 U9768 ( .A(n7745), .B(n16042), .ZN(SUB_1596_U4) );
  NAND2_X1 U9769 ( .A1(n16033), .A2(n16034), .ZN(n7745) );
  NAND2_X1 U9770 ( .A1(n16319), .A2(n16318), .ZN(n7983) );
  NAND2_X1 U9771 ( .A1(n16280), .A2(n16279), .ZN(n7978) );
  NAND2_X1 U9772 ( .A1(n8180), .A2(n14400), .ZN(n14543) );
  AND4_X2 U9773 ( .A1(n7898), .A2(n7900), .A3(n7901), .A4(n7899), .ZN(n7928)
         );
  AOI21_X1 U9774 ( .B1(n14470), .B2(n14473), .A(n14411), .ZN(n14453) );
  NAND2_X1 U9775 ( .A1(n11059), .A2(n11058), .ZN(n11241) );
  NAND2_X1 U9776 ( .A1(n8181), .A2(n7513), .ZN(n11781) );
  NAND2_X1 U9777 ( .A1(n14558), .A2(n14398), .ZN(n8180) );
  NAND2_X1 U9778 ( .A1(n14588), .A2(n14589), .ZN(n14394) );
  OAI21_X1 U9779 ( .B1(n9699), .B2(n8272), .A(n7750), .ZN(n9720) );
  OAI21_X1 U9780 ( .B1(n9777), .B2(n9776), .A(n9775), .ZN(n9778) );
  NAND2_X2 U9781 ( .A1(n9152), .A2(n9360), .ZN(n9574) );
  NAND2_X1 U9782 ( .A1(n8846), .A2(n8845), .ZN(n8861) );
  INV_X1 U9783 ( .A(n8964), .ZN(n8032) );
  NAND2_X1 U9784 ( .A1(n8710), .A2(n8709), .ZN(n8726) );
  NAND2_X1 U9785 ( .A1(n8064), .A2(n8784), .ZN(n8068) );
  NAND2_X1 U9786 ( .A1(n8807), .A2(n8806), .ZN(n8821) );
  NAND2_X1 U9787 ( .A1(n11012), .A2(n11017), .ZN(n11401) );
  NAND2_X1 U9788 ( .A1(n11403), .A2(n11401), .ZN(n11040) );
  NAND2_X1 U9789 ( .A1(n7765), .A2(n7764), .ZN(n12005) );
  NAND3_X1 U9790 ( .A1(n7767), .A2(n11421), .A3(n7484), .ZN(n7764) );
  NAND2_X1 U9791 ( .A1(n11421), .A2(n7767), .ZN(n11423) );
  INV_X1 U9792 ( .A(n13323), .ZN(n7775) );
  INV_X1 U9793 ( .A(n8259), .ZN(n13363) );
  XNOR2_X2 U9794 ( .A(n8247), .B(n13234), .ZN(n12284) );
  NAND4_X1 U9795 ( .A1(n8419), .A2(n7870), .A3(n8553), .A4(n8524), .ZN(n8639)
         );
  NAND2_X1 U9796 ( .A1(n7793), .A2(n7794), .ZN(n8925) );
  NAND2_X1 U9797 ( .A1(n13534), .A2(n7796), .ZN(n7793) );
  NAND2_X1 U9798 ( .A1(n8079), .A2(n7801), .ZN(n11979) );
  OAI21_X1 U9799 ( .B1(n7483), .B2(n7803), .A(n16565), .ZN(n7804) );
  NAND2_X1 U9800 ( .A1(n7813), .A2(n7812), .ZN(n13577) );
  NAND2_X1 U9801 ( .A1(n9099), .A2(n7588), .ZN(n13742) );
  NAND2_X1 U9802 ( .A1(n9099), .A2(n8534), .ZN(n9102) );
  OAI21_X1 U9803 ( .B1(n7468), .B2(n11207), .A(n7819), .ZN(n7818) );
  NAND2_X1 U9804 ( .A1(n12062), .A2(n12063), .ZN(n12173) );
  NAND2_X1 U9805 ( .A1(n9385), .A2(n9191), .ZN(n7841) );
  NAND2_X1 U9806 ( .A1(n9359), .A2(n9188), .ZN(n7842) );
  INV_X1 U9807 ( .A(n9253), .ZN(n9731) );
  NAND2_X1 U9808 ( .A1(n10196), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7854) );
  AND2_X1 U9809 ( .A1(n10196), .A2(P3_U3151), .ZN(n13739) );
  MUX2_X1 U9810 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n10196), .Z(n9185) );
  MUX2_X1 U9811 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n10196), .Z(n9832) );
  NAND3_X1 U9812 ( .A1(n8224), .A2(n8227), .A3(n9521), .ZN(n7864) );
  NOR2_X1 U9813 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n7870) );
  NOR2_X1 U9814 ( .A1(n11221), .A2(n11222), .ZN(n11220) );
  MUX2_X1 U9815 ( .A(P3_REG1_REG_1__SCAN_IN), .B(P3_REG2_REG_1__SCAN_IN), .S(
        n12285), .Z(n10921) );
  NAND4_X1 U9816 ( .A1(n7874), .A2(n8254), .A3(n7873), .A4(n7536), .ZN(
        P3_U3201) );
  NAND2_X1 U9817 ( .A1(n10856), .A2(n10855), .ZN(n11114) );
  NAND2_X1 U9818 ( .A1(n10522), .A2(n10517), .ZN(n7875) );
  XNOR2_X2 U9819 ( .A(n9160), .B(n9159), .ZN(n12551) );
  NAND2_X1 U9820 ( .A1(n9158), .A2(n7890), .ZN(n15902) );
  AND2_X2 U9821 ( .A1(n10049), .A2(n9949), .ZN(n9952) );
  NOR2_X2 U9822 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7899) );
  NOR2_X2 U9823 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7900) );
  NOR2_X2 U9824 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n7901) );
  INV_X1 U9825 ( .A(n12767), .ZN(n7905) );
  NAND2_X1 U9826 ( .A1(n12728), .A2(n7913), .ZN(n7909) );
  NAND2_X1 U9827 ( .A1(n7916), .A2(n10764), .ZN(n10770) );
  NOR2_X1 U9828 ( .A1(n10658), .A2(n10149), .ZN(n7917) );
  OAI21_X2 U9829 ( .B1(n13940), .B2(n8153), .A(n8152), .ZN(n8159) );
  NAND2_X2 U9830 ( .A1(n13872), .A2(n7919), .ZN(n13940) );
  NAND2_X2 U9831 ( .A1(n7922), .A2(n7921), .ZN(n8146) );
  OR2_X2 U9832 ( .A1(n12095), .A2(n7502), .ZN(n7922) );
  OR2_X2 U9833 ( .A1(n13921), .A2(n13922), .ZN(n13919) );
  NAND2_X1 U9834 ( .A1(n10817), .A2(n10816), .ZN(n10819) );
  NAND2_X1 U9835 ( .A1(n10832), .A2(n10798), .ZN(n7926) );
  NAND2_X1 U9836 ( .A1(n7929), .A2(n7930), .ZN(n14425) );
  INV_X1 U9837 ( .A(n13992), .ZN(n13995) );
  NAND2_X1 U9838 ( .A1(n14606), .A2(n7952), .ZN(n7950) );
  NAND2_X1 U9839 ( .A1(n7950), .A2(n7566), .ZN(n14433) );
  NOR2_X2 U9840 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n10049) );
  NAND2_X1 U9841 ( .A1(n7956), .A2(n14078), .ZN(n7955) );
  NAND2_X1 U9842 ( .A1(n14079), .A2(n14080), .ZN(n7956) );
  INV_X1 U9843 ( .A(n14079), .ZN(n7958) );
  AND2_X1 U9844 ( .A1(n10013), .A2(n8516), .ZN(n7969) );
  AND2_X1 U9845 ( .A1(n14033), .A2(n14034), .ZN(n7972) );
  AND2_X1 U9846 ( .A1(n15999), .A2(n15998), .ZN(n16282) );
  NAND2_X1 U9847 ( .A1(n7987), .A2(n10542), .ZN(n10540) );
  INV_X2 U9848 ( .A(n14005), .ZN(n16418) );
  NAND2_X2 U9849 ( .A1(n8292), .A2(n8293), .ZN(n14005) );
  NOR2_X2 U9850 ( .A1(n14491), .A2(n14672), .ZN(n7991) );
  NOR2_X2 U9851 ( .A1(n14647), .A2(n14728), .ZN(n7993) );
  NOR2_X2 U9852 ( .A1(n12142), .A2(n14108), .ZN(n12232) );
  INV_X2 U9853 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7998) );
  OR2_X1 U9854 ( .A1(n11109), .A2(n14843), .ZN(n8000) );
  NAND2_X1 U9855 ( .A1(n15124), .A2(n8003), .ZN(n15093) );
  AND2_X1 U9856 ( .A1(n15124), .A2(n15376), .ZN(n15114) );
  NAND2_X1 U9857 ( .A1(n15124), .A2(n8001), .ZN(n15080) );
  NAND2_X1 U9858 ( .A1(n12343), .A2(n8006), .ZN(n15293) );
  NOR2_X2 U9859 ( .A1(n15220), .A2(n15408), .ZN(n15197) );
  NAND2_X1 U9860 ( .A1(n8249), .A2(n10928), .ZN(n8013) );
  NAND2_X1 U9861 ( .A1(n8249), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10956) );
  NAND2_X1 U9862 ( .A1(n8249), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10964) );
  OR2_X1 U9863 ( .A1(n8249), .A2(P3_U3151), .ZN(n8015) );
  NAND2_X1 U9864 ( .A1(n7613), .A2(n8249), .ZN(n8556) );
  XNOR2_X1 U9865 ( .A(n10953), .B(n8249), .ZN(n10954) );
  INV_X1 U9866 ( .A(n8249), .ZN(n8018) );
  NAND2_X1 U9867 ( .A1(n8021), .A2(n11407), .ZN(n8019) );
  INV_X1 U9868 ( .A(n10961), .ZN(n8026) );
  INV_X1 U9869 ( .A(n8900), .ZN(n8034) );
  AOI21_X1 U9870 ( .B1(n8034), .B2(n8913), .A(n8926), .ZN(n8033) );
  INV_X1 U9871 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8036) );
  NAND2_X1 U9872 ( .A1(n8623), .A2(n8039), .ZN(n8038) );
  NAND2_X1 U9873 ( .A1(n8677), .A2(n8049), .ZN(n8046) );
  NAND2_X1 U9874 ( .A1(n8046), .A2(n8047), .ZN(n8710) );
  NAND2_X1 U9875 ( .A1(n8864), .A2(n8055), .ZN(n8052) );
  NAND2_X1 U9876 ( .A1(n8729), .A2(n8061), .ZN(n8058) );
  NAND2_X1 U9877 ( .A1(n8781), .A2(n10340), .ZN(n8064) );
  NAND2_X1 U9878 ( .A1(n8066), .A2(n8069), .ZN(n8804) );
  NAND2_X1 U9879 ( .A1(n8765), .A2(n8781), .ZN(n8066) );
  NOR2_X1 U9880 ( .A1(n13425), .A2(n12841), .ZN(n8073) );
  OAI21_X1 U9881 ( .B1(n11806), .B2(n8078), .A(n8076), .ZN(n8079) );
  NAND2_X1 U9882 ( .A1(n13566), .A2(n8080), .ZN(n13534) );
  OAI21_X1 U9883 ( .B1(n9068), .B2(n7607), .A(n8087), .ZN(P3_U3456) );
  OR2_X1 U9884 ( .A1(n9068), .A2(n13582), .ZN(n8090) );
  NAND2_X1 U9885 ( .A1(n8093), .A2(n8092), .ZN(n12074) );
  NAND2_X1 U9886 ( .A1(n14897), .A2(n8101), .ZN(n8100) );
  AND2_X1 U9887 ( .A1(n11723), .A2(n11721), .ZN(n8105) );
  NAND2_X1 U9888 ( .A1(n10783), .A2(n10782), .ZN(n10905) );
  NAND2_X1 U9889 ( .A1(n10905), .A2(n10906), .ZN(n8114) );
  NAND2_X1 U9890 ( .A1(n14820), .A2(n8116), .ZN(n8115) );
  OAI211_X1 U9891 ( .C1(n14820), .C2(n8117), .A(n12716), .B(n8115), .ZN(
        P1_U3220) );
  AOI21_X1 U9892 ( .B1(n8132), .B2(n8128), .A(n7590), .ZN(n8127) );
  INV_X1 U9893 ( .A(n12257), .ZN(n8128) );
  INV_X1 U9894 ( .A(n8132), .ZN(n8129) );
  AND2_X1 U9895 ( .A1(n8288), .A2(n7481), .ZN(n9927) );
  NAND2_X1 U9896 ( .A1(n8288), .A2(n7540), .ZN(n9934) );
  NAND2_X1 U9897 ( .A1(n8760), .A2(n8759), .ZN(n12473) );
  NAND2_X1 U9898 ( .A1(n8739), .A2(n8738), .ZN(n12392) );
  NAND2_X1 U9899 ( .A1(n12074), .A2(n8717), .ZN(n12240) );
  NAND2_X1 U9900 ( .A1(n8780), .A2(n8779), .ZN(n12465) );
  OR2_X1 U9901 ( .A1(n10053), .A2(n10172), .ZN(n10032) );
  NOR2_X1 U9902 ( .A1(n13992), .A2(n13951), .ZN(n11333) );
  NOR2_X2 U9903 ( .A1(n14371), .A2(n7458), .ZN(n14656) );
  NOR2_X4 U9904 ( .A1(n14618), .A2(n14593), .ZN(n14597) );
  NAND3_X1 U9905 ( .A1(n14916), .A2(n14830), .A3(n14831), .ZN(n14829) );
  NAND2_X2 U9906 ( .A1(n13919), .A2(n13785), .ZN(n13798) );
  NAND2_X1 U9907 ( .A1(n10127), .A2(n14366), .ZN(n8138) );
  OAI21_X1 U9908 ( .B1(n10127), .B2(n13982), .A(n14366), .ZN(n8139) );
  NAND2_X1 U9909 ( .A1(n11344), .A2(n8142), .ZN(n8140) );
  NAND2_X1 U9910 ( .A1(n8140), .A2(n8141), .ZN(n11896) );
  AOI21_X1 U9911 ( .B1(n8142), .B2(n7470), .A(n7546), .ZN(n8141) );
  INV_X1 U9912 ( .A(n8159), .ZN(n13853) );
  NAND2_X2 U9913 ( .A1(n10042), .A2(n10196), .ZN(n10053) );
  NAND2_X2 U9914 ( .A1(n10278), .A2(n14807), .ZN(n10042) );
  NAND2_X1 U9915 ( .A1(n12220), .A2(n8170), .ZN(n8169) );
  NAND2_X1 U9916 ( .A1(n11782), .A2(n8176), .ZN(n8174) );
  NAND2_X1 U9917 ( .A1(n10822), .A2(n7509), .ZN(n11059) );
  NAND2_X1 U9918 ( .A1(n11241), .A2(n11240), .ZN(n11244) );
  NAND2_X1 U9919 ( .A1(n11501), .A2(n8183), .ZN(n8181) );
  NAND2_X1 U9920 ( .A1(n14505), .A2(n8188), .ZN(n14409) );
  INV_X1 U9921 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n15072) );
  INV_X1 U9922 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n8192) );
  INV_X1 U9923 ( .A(P1_RD_REG_SCAN_IN), .ZN(n8194) );
  INV_X1 U9924 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8195) );
  INV_X1 U9925 ( .A(n9309), .ZN(n8196) );
  NAND2_X1 U9926 ( .A1(n9425), .A2(n8200), .ZN(n8197) );
  OAI21_X1 U9927 ( .B1(n9824), .B2(n8215), .A(n8211), .ZN(n9834) );
  OAI21_X1 U9928 ( .B1(n9540), .B2(n9539), .A(n9220), .ZN(n9558) );
  OAI21_X1 U9929 ( .B1(n9487), .B2(n9486), .A(n9210), .ZN(n9500) );
  NAND2_X1 U9930 ( .A1(n8235), .A2(n8233), .ZN(n8231) );
  NAND2_X1 U9931 ( .A1(n9256), .A2(n9255), .ZN(n9750) );
  NAND2_X1 U9932 ( .A1(n8239), .A2(n8242), .ZN(n11287) );
  NAND2_X1 U9933 ( .A1(n10970), .A2(n11284), .ZN(n8239) );
  INV_X1 U9934 ( .A(n8242), .ZN(n8241) );
  OR2_X2 U9935 ( .A1(n8555), .A2(n8250), .ZN(n8249) );
  NAND3_X1 U9936 ( .A1(n9398), .A2(n7563), .A3(n9397), .ZN(n8260) );
  NAND2_X1 U9937 ( .A1(n8262), .A2(n8263), .ZN(n9620) );
  NAND3_X1 U9938 ( .A1(n9585), .A2(n7582), .A3(n9584), .ZN(n8262) );
  NAND2_X1 U9939 ( .A1(n8264), .A2(n8265), .ZN(n9506) );
  NAND3_X1 U9940 ( .A1(n9478), .A2(n7583), .A3(n9477), .ZN(n8264) );
  NAND2_X1 U9941 ( .A1(n8266), .A2(n8267), .ZN(n9580) );
  NAND3_X1 U9942 ( .A1(n9552), .A2(n7578), .A3(n9551), .ZN(n8266) );
  NAND2_X1 U9943 ( .A1(n8268), .A2(n8269), .ZN(n9717) );
  NAND2_X1 U9944 ( .A1(n9699), .A2(n8271), .ZN(n8268) );
  NAND2_X1 U9945 ( .A1(n8273), .A2(n8274), .ZN(n9473) );
  NAND3_X1 U9946 ( .A1(n9433), .A2(n9434), .A3(n7584), .ZN(n8273) );
  NAND2_X1 U9947 ( .A1(n8276), .A2(n8277), .ZN(n9663) );
  NAND3_X1 U9948 ( .A1(n9625), .A2(n7585), .A3(n9624), .ZN(n8276) );
  NAND2_X1 U9949 ( .A1(n8279), .A2(n8280), .ZN(n9547) );
  NAND3_X1 U9950 ( .A1(n9511), .A2(n7577), .A3(n9510), .ZN(n8279) );
  NAND2_X1 U9951 ( .A1(n8282), .A2(n8283), .ZN(n9769) );
  NAND3_X1 U9952 ( .A1(n9741), .A2(n7579), .A3(n9740), .ZN(n8282) );
  NAND2_X1 U9953 ( .A1(n9976), .A2(n10413), .ZN(n9811) );
  NAND2_X1 U9954 ( .A1(n9998), .A2(n15185), .ZN(n10413) );
  NAND3_X1 U9955 ( .A1(n11549), .A2(n10413), .A3(n9976), .ZN(n8289) );
  INV_X1 U9956 ( .A(n14497), .ZN(n8302) );
  NAND2_X1 U9957 ( .A1(n8299), .A2(n14497), .ZN(n8297) );
  AND2_X1 U9958 ( .A1(n10013), .A2(n8166), .ZN(n8303) );
  INV_X2 U9959 ( .A(n9303), .ZN(n9804) );
  INV_X1 U9960 ( .A(n9933), .ZN(n8316) );
  NAND2_X1 U9961 ( .A1(n8316), .A2(n7703), .ZN(n8317) );
  NAND2_X1 U9962 ( .A1(n12152), .A2(n8321), .ZN(n8318) );
  NAND2_X1 U9963 ( .A1(n8318), .A2(n8319), .ZN(n12332) );
  NAND2_X1 U9964 ( .A1(n10847), .A2(n9316), .ZN(n10524) );
  OAI21_X2 U9965 ( .B1(n15109), .B2(n15110), .A(n8338), .ZN(n15091) );
  NOR2_X1 U9966 ( .A1(n10715), .A2(n8343), .ZN(n10627) );
  AND2_X1 U9967 ( .A1(n8344), .A2(n10601), .ZN(n8343) );
  NAND2_X1 U9968 ( .A1(n10600), .A2(n10713), .ZN(n8344) );
  INV_X1 U9969 ( .A(n13533), .ZN(n8346) );
  NAND2_X1 U9970 ( .A1(n11303), .A2(n8357), .ZN(n8356) );
  NAND2_X1 U9971 ( .A1(n12121), .A2(n8368), .ZN(n8365) );
  INV_X1 U9972 ( .A(n12120), .ZN(n8373) );
  NAND2_X1 U9973 ( .A1(n12491), .A2(n8376), .ZN(n8375) );
  NAND2_X1 U9974 ( .A1(n13180), .A2(n12831), .ZN(n13072) );
  NAND2_X1 U9975 ( .A1(n13180), .A2(n8380), .ZN(n8379) );
  NOR2_X1 U9976 ( .A1(n8383), .A2(n12835), .ZN(n8380) );
  OAI22_X1 U9977 ( .A1(n8383), .A2(n8382), .B1(n12835), .B2(n8385), .ZN(n8381)
         );
  NOR2_X1 U9978 ( .A1(n12835), .A2(n13073), .ZN(n8382) );
  INV_X1 U9979 ( .A(n8385), .ZN(n8383) );
  NAND2_X1 U9980 ( .A1(n13073), .A2(n12835), .ZN(n8384) );
  NAND2_X1 U9981 ( .A1(n11804), .A2(n8395), .ZN(n8394) );
  NAND2_X1 U9982 ( .A1(n8394), .A2(n8397), .ZN(n11978) );
  OAI21_X1 U9983 ( .B1(n13576), .B2(n8408), .A(n8406), .ZN(n13558) );
  OAI21_X1 U9984 ( .B1(n13576), .B2(n13575), .A(n12929), .ZN(n13562) );
  NAND2_X1 U9985 ( .A1(n8414), .A2(n13133), .ZN(n12822) );
  NAND2_X1 U9986 ( .A1(n12858), .A2(n12857), .ZN(n16370) );
  NAND2_X1 U9987 ( .A1(n11733), .A2(n8425), .ZN(n8424) );
  OAI21_X1 U9988 ( .B1(n11733), .B2(n11745), .A(n8425), .ZN(n11827) );
  NAND3_X1 U9989 ( .A1(n8424), .A2(n11826), .A3(n8423), .ZN(n11825) );
  NAND2_X1 U9990 ( .A1(n8425), .A2(n11745), .ZN(n8423) );
  NAND2_X1 U9991 ( .A1(n9158), .A2(n9157), .ZN(n9936) );
  NAND2_X1 U9992 ( .A1(n12340), .A2(n8432), .ZN(n8431) );
  NOR2_X1 U9993 ( .A1(n12574), .A2(n12573), .ZN(n8436) );
  NAND2_X1 U9994 ( .A1(n15216), .A2(n8442), .ZN(n8441) );
  INV_X1 U9995 ( .A(n12645), .ZN(n8453) );
  INV_X1 U9996 ( .A(n8460), .ZN(n12310) );
  INV_X1 U9997 ( .A(n15281), .ZN(n8475) );
  INV_X1 U9998 ( .A(n14177), .ZN(n8492) );
  XNOR2_X2 U9999 ( .A(n10026), .B(n10025), .ZN(n10278) );
  NAND2_X1 U10000 ( .A1(n8496), .A2(n7581), .ZN(n14071) );
  NAND2_X1 U10001 ( .A1(n8498), .A2(n8497), .ZN(n8496) );
  INV_X1 U10002 ( .A(n14057), .ZN(n8498) );
  NAND2_X1 U10003 ( .A1(n8502), .A2(n8501), .ZN(n14035) );
  NAND2_X1 U10004 ( .A1(n14029), .A2(n7587), .ZN(n8501) );
  NAND2_X1 U10005 ( .A1(n8505), .A2(n8504), .ZN(n8503) );
  INV_X1 U10006 ( .A(n14029), .ZN(n8505) );
  INV_X1 U10007 ( .A(n14119), .ZN(n8507) );
  NAND2_X1 U10008 ( .A1(n10441), .A2(n9948), .ZN(n16258) );
  OR2_X1 U10009 ( .A1(n7461), .A2(n11315), .ZN(n8948) );
  OR2_X1 U10010 ( .A1(n12784), .A2(n9027), .ZN(n9029) );
  OR2_X1 U10011 ( .A1(n12043), .A2(n9027), .ZN(n9002) );
  OR2_X1 U10012 ( .A1(n11923), .A2(n9027), .ZN(n8982) );
  OR2_X1 U10013 ( .A1(n11104), .A2(n9027), .ZN(n8937) );
  OR2_X1 U10014 ( .A1(n10657), .A2(n9027), .ZN(n8904) );
  INV_X1 U10015 ( .A(n9598), .ZN(n9614) );
  NOR2_X2 U10016 ( .A1(n12602), .A2(n12601), .ZN(n14945) );
  CLKBUF_X1 U10017 ( .A(n10591), .Z(n9141) );
  NAND2_X1 U10018 ( .A1(n9868), .A2(n8521), .ZN(n9887) );
  AND2_X1 U10019 ( .A1(n15087), .A2(n12582), .ZN(n15370) );
  AOI22_X1 U10020 ( .A1(n10777), .A2(n10776), .B1(n10775), .B2(n10774), .ZN(
        n14842) );
  NAND2_X1 U10021 ( .A1(n10599), .A2(n8573), .ZN(n10713) );
  NAND2_X1 U10022 ( .A1(n12551), .A2(n9165), .ZN(n9304) );
  XNOR2_X1 U10023 ( .A(n14026), .B(n14318), .ZN(n14252) );
  OAI21_X1 U10024 ( .B1(n12463), .B2(n9077), .A(n12927), .ZN(n13576) );
  INV_X1 U10025 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10041) );
  NAND2_X1 U10026 ( .A1(n10162), .A2(n14641), .ZN(n13952) );
  CLKBUF_X2 U10027 ( .A(P2_U3947), .Z(n14322) );
  OR2_X1 U10028 ( .A1(n12485), .A2(n12484), .ZN(n8508) );
  INV_X1 U10029 ( .A(n13557), .ZN(n8859) );
  AND2_X1 U10030 ( .A1(n8753), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8509) );
  NOR2_X1 U10031 ( .A1(n9080), .A2(n13462), .ZN(n8510) );
  NOR2_X1 U10032 ( .A1(n13469), .A2(n13454), .ZN(n8511) );
  AND2_X1 U10033 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8512) );
  AND2_X1 U10034 ( .A1(n12653), .A2(n12652), .ZN(n8514) );
  OR2_X1 U10035 ( .A1(n10494), .A2(n10450), .ZN(n15232) );
  NOR2_X1 U10036 ( .A1(n13064), .A2(n16386), .ZN(n8515) );
  INV_X1 U10037 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n9091) );
  NOR2_X1 U10038 ( .A1(n10015), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n8516) );
  AND2_X1 U10039 ( .A1(n9214), .A2(n9213), .ZN(n8517) );
  AND2_X2 U10040 ( .A1(n10689), .A2(n9132), .ZN(n16565) );
  AND2_X1 U10041 ( .A1(n9480), .A2(n9479), .ZN(n8518) );
  AND2_X1 U10042 ( .A1(n13383), .A2(n16561), .ZN(n8519) );
  AND2_X1 U10043 ( .A1(n14225), .A2(n14220), .ZN(n8520) );
  AND2_X1 U10044 ( .A1(n9882), .A2(n9869), .ZN(n8521) );
  AND2_X1 U10045 ( .A1(n9880), .A2(n9883), .ZN(n8522) );
  INV_X1 U10046 ( .A(n16411), .ZN(n13492) );
  MUX2_X1 U10047 ( .A(n9289), .B(n9288), .S(n10516), .Z(n9318) );
  OAI21_X1 U10048 ( .B1(n13995), .B2(n14238), .A(n13994), .ZN(n13996) );
  INV_X1 U10049 ( .A(n9374), .ZN(n9375) );
  INV_X1 U10050 ( .A(n14080), .ZN(n14081) );
  INV_X1 U10051 ( .A(n14095), .ZN(n14096) );
  INV_X1 U10052 ( .A(n14122), .ZN(n14123) );
  INV_X1 U10053 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9950) );
  INV_X1 U10054 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8529) );
  INV_X1 U10055 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n15868) );
  INV_X1 U10056 ( .A(n8939), .ZN(n8938) );
  INV_X1 U10057 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8524) );
  INV_X1 U10058 ( .A(n12816), .ZN(n12814) );
  NAND2_X1 U10059 ( .A1(n8575), .A2(n8574), .ZN(n11131) );
  INV_X1 U10060 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9053) );
  INV_X1 U10061 ( .A(n13817), .ZN(n13758) );
  INV_X1 U10062 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n11354) );
  NOR2_X1 U10063 ( .A1(n11966), .A2(n11965), .ZN(n11967) );
  INV_X1 U10064 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9513) );
  INV_X1 U10065 ( .A(n9755), .ZN(n9166) );
  INV_X1 U10066 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9453) );
  INV_X1 U10067 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n15885) );
  NAND2_X1 U10068 ( .A1(n9598), .A2(n15684), .ZN(n9273) );
  NOR2_X1 U10069 ( .A1(n10595), .A2(n10594), .ZN(n10596) );
  NAND2_X1 U10070 ( .A1(n12488), .A2(n13153), .ZN(n12489) );
  INV_X1 U10071 ( .A(n12841), .ZN(n9083) );
  AND2_X1 U10072 ( .A1(n12880), .A2(n12881), .ZN(n13015) );
  OAI22_X1 U10073 ( .A1(n13076), .A2(n16374), .B1(n13373), .B2(n13007), .ZN(
        n9066) );
  OR2_X1 U10074 ( .A1(n13604), .A2(n13603), .ZN(n13605) );
  INV_X1 U10075 ( .A(n12961), .ZN(n12975) );
  AND2_X1 U10076 ( .A1(n13064), .A2(n12855), .ZN(n12961) );
  AND2_X1 U10077 ( .A1(n8725), .A2(n8708), .ZN(n8709) );
  INV_X1 U10078 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10751) );
  INV_X1 U10079 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10997) );
  NAND2_X1 U10080 ( .A1(n10042), .A2(n14819), .ZN(n10040) );
  OR2_X1 U10081 ( .A1(n13829), .A2(n13759), .ZN(n13857) );
  NAND2_X1 U10082 ( .A1(n12221), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n12357) );
  INV_X1 U10083 ( .A(n14313), .ZN(n14062) );
  INV_X1 U10084 ( .A(n11967), .ZN(n11968) );
  AND2_X1 U10085 ( .A1(n12259), .A2(n12256), .ZN(n12257) );
  NAND2_X1 U10086 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n9743), .ZN(n9755) );
  OR2_X1 U10087 ( .A1(n9649), .A2(n14910), .ZN(n9669) );
  OR2_X1 U10088 ( .A1(n9514), .A2(n9513), .ZN(n9533) );
  INV_X1 U10089 ( .A(n10497), .ZN(n10475) );
  INV_X1 U10090 ( .A(n15920), .ZN(n9940) );
  NAND2_X1 U10091 ( .A1(n9221), .A2(n15521), .ZN(n9224) );
  NOR2_X1 U10092 ( .A1(P3_ADDR_REG_8__SCAN_IN), .A2(n15941), .ZN(n15943) );
  NAND2_X1 U10093 ( .A1(n11878), .A2(n13222), .ZN(n11879) );
  OR2_X1 U10094 ( .A1(n8796), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8813) );
  NOR2_X1 U10095 ( .A1(n8888), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8907) );
  NAND2_X1 U10096 ( .A1(n8853), .A2(n15575), .ZN(n8870) );
  NAND2_X1 U10097 ( .A1(n8967), .A2(n15576), .ZN(n8983) );
  OR2_X1 U10098 ( .A1(n8870), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8888) );
  NAND2_X1 U10099 ( .A1(n10619), .A2(n10617), .ZN(n13187) );
  AND2_X1 U10100 ( .A1(n10946), .A2(n10944), .ZN(n10938) );
  OR2_X1 U10101 ( .A1(n8616), .A2(n15700), .ZN(n9007) );
  AND2_X1 U10102 ( .A1(n12925), .A2(n12471), .ZN(n13029) );
  AND2_X1 U10103 ( .A1(n9139), .A2(n13056), .ZN(n13582) );
  AND2_X1 U10104 ( .A1(n14814), .A2(n12401), .ZN(n9962) );
  NAND2_X1 U10105 ( .A1(n12512), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n12524) );
  NAND2_X1 U10106 ( .A1(n12522), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n13803) );
  INV_X1 U10107 ( .A(n13972), .ZN(n13943) );
  AND2_X1 U10108 ( .A1(n14278), .A2(n14277), .ZN(n14279) );
  AND2_X1 U10109 ( .A1(n13857), .A2(n13760), .ZN(n14494) );
  OR2_X1 U10110 ( .A1(n12439), .A2(n12438), .ZN(n12513) );
  INV_X1 U10111 ( .A(n14272), .ZN(n14424) );
  AND2_X1 U10112 ( .A1(n14630), .A2(n12215), .ZN(n14270) );
  INV_X1 U10113 ( .A(n10505), .ZN(n10117) );
  NAND2_X2 U10114 ( .A1(n10070), .A2(n10069), .ZN(n14026) );
  OR3_X1 U10115 ( .A1(n14739), .A2(n14738), .A3(n14737), .ZN(n14787) );
  INV_X1 U10116 ( .A(n14084), .ZN(n16572) );
  AND2_X1 U10117 ( .A1(n10103), .A2(n14809), .ZN(n16074) );
  NAND2_X1 U10118 ( .A1(n9960), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9957) );
  INV_X1 U10119 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n10203) );
  INV_X1 U10120 ( .A(n14965), .ZN(n12156) );
  OR2_X1 U10121 ( .A1(n9669), .A2(n14862), .ZN(n9690) );
  OR2_X1 U10122 ( .A1(n9587), .A2(n9586), .ZN(n9606) );
  AND2_X1 U10123 ( .A1(n14908), .A2(n14905), .ZN(n12640) );
  OR2_X1 U10124 ( .A1(n14836), .A2(n15232), .ZN(n14951) );
  NAND2_X1 U10125 ( .A1(n9860), .A2(n8522), .ZN(n9888) );
  NOR2_X1 U10126 ( .A1(n9690), .A2(n14919), .ZN(n9702) );
  NAND2_X1 U10127 ( .A1(n9568), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9587) );
  XNOR2_X1 U10128 ( .A(n15388), .B(n15132), .ZN(n15143) );
  INV_X1 U10129 ( .A(n12566), .ZN(n15180) );
  NAND2_X1 U10130 ( .A1(n15287), .A2(n12558), .ZN(n15268) );
  OR2_X1 U10131 ( .A1(n10407), .A2(n10406), .ZN(n10499) );
  INV_X1 U10132 ( .A(n12552), .ZN(n12339) );
  NAND2_X1 U10133 ( .A1(n10265), .A2(n10450), .ZN(n15230) );
  OR2_X1 U10134 ( .A1(n11163), .A2(n15185), .ZN(n15361) );
  NAND2_X1 U10135 ( .A1(n9997), .A2(n10257), .ZN(n10497) );
  INV_X1 U10136 ( .A(n13187), .ZN(n13196) );
  NAND2_X1 U10137 ( .A1(n12811), .A2(n12813), .ZN(n13164) );
  NAND2_X1 U10138 ( .A1(n10622), .A2(n16405), .ZN(n13168) );
  AND4_X1 U10139 ( .A1(n13004), .A2(n9065), .A3(n9064), .A4(n9063), .ZN(n13007) );
  AND4_X1 U10140 ( .A1(n8944), .A2(n8943), .A3(n8942), .A4(n8941), .ZN(n13100)
         );
  INV_X1 U10141 ( .A(n16327), .ZN(n13342) );
  MUX2_X1 U10142 ( .A(n10938), .B(n16079), .S(n13061), .Z(n13370) );
  INV_X1 U10143 ( .A(n16372), .ZN(n13498) );
  AOI21_X1 U10144 ( .B1(n16380), .B2(n11595), .A(n13492), .ZN(n13559) );
  INV_X1 U10145 ( .A(n13587), .ZN(n13555) );
  AND2_X1 U10146 ( .A1(n9123), .A2(n9122), .ZN(n10689) );
  OR2_X1 U10147 ( .A1(n13661), .A2(n8515), .ZN(n16561) );
  OR2_X1 U10148 ( .A1(n9106), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9108) );
  INV_X1 U10149 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8546) );
  AND2_X1 U10150 ( .A1(n14295), .A2(n10125), .ZN(n10269) );
  INV_X1 U10151 ( .A(n13915), .ZN(n13977) );
  INV_X1 U10152 ( .A(n16234), .ZN(n16189) );
  AND2_X1 U10153 ( .A1(n16237), .A2(P2_STATE_REG_SCAN_IN), .ZN(n16234) );
  AND2_X1 U10154 ( .A1(n10283), .A2(n10274), .ZN(n10275) );
  NAND2_X1 U10155 ( .A1(n14416), .A2(n14415), .ZN(n14417) );
  INV_X1 U10156 ( .A(n14553), .ZN(n14650) );
  INV_X1 U10157 ( .A(n16585), .ZN(n12115) );
  OR2_X1 U10158 ( .A1(n10508), .A2(n10507), .ZN(n10639) );
  NAND2_X1 U10159 ( .A1(n10081), .A2(n10080), .ZN(n10084) );
  OR2_X1 U10160 ( .A1(n10702), .A2(n10701), .ZN(n10703) );
  INV_X1 U10161 ( .A(n16266), .ZN(n16354) );
  INV_X1 U10162 ( .A(n15130), .ZN(n15122) );
  INV_X1 U10163 ( .A(n15232), .ZN(n15329) );
  INV_X1 U10164 ( .A(n15337), .ZN(n15309) );
  NAND3_X2 U10165 ( .A1(n9315), .A2(n9314), .A3(n9313), .ZN(n15342) );
  AND2_X1 U10166 ( .A1(n15338), .A2(n10001), .ZN(n15345) );
  NOR2_X1 U10167 ( .A1(n10499), .A2(n10409), .ZN(n10476) );
  NOR2_X1 U10168 ( .A1(n15238), .A2(n15237), .ZN(n15426) );
  INV_X1 U10169 ( .A(n16547), .ZN(n15463) );
  NAND2_X1 U10170 ( .A1(n15361), .A2(n15475), .ZN(n16547) );
  AND2_X1 U10171 ( .A1(n10497), .A2(n10474), .ZN(n10534) );
  NAND2_X1 U10172 ( .A1(n9981), .A2(n9982), .ZN(n10256) );
  INV_X1 U10173 ( .A(n9998), .ZN(n9838) );
  OR3_X1 U10174 ( .A1(n11922), .A2(n9105), .A3(n12042), .ZN(n10609) );
  INV_X1 U10175 ( .A(n13168), .ZN(n13199) );
  INV_X1 U10176 ( .A(n13100), .ZN(n13499) );
  INV_X1 U10177 ( .A(n16373), .ZN(n13226) );
  INV_X1 U10178 ( .A(n16336), .ZN(n13368) );
  OR2_X1 U10179 ( .A1(n10935), .A2(n12285), .ZN(n16328) );
  INV_X1 U10180 ( .A(n13559), .ZN(n13590) );
  NAND2_X2 U10181 ( .A1(n10690), .A2(n16405), .ZN(n16411) );
  INV_X1 U10182 ( .A(n16565), .ZN(n16563) );
  INV_X1 U10183 ( .A(n13179), .ZN(n13681) );
  INV_X1 U10184 ( .A(n16569), .ZN(n16566) );
  NAND2_X1 U10185 ( .A1(n9106), .A2(n13737), .ZN(n10377) );
  AND2_X1 U10186 ( .A1(n9108), .A2(n9107), .ZN(n13738) );
  INV_X1 U10187 ( .A(n9138), .ZN(n10655) );
  INV_X1 U10188 ( .A(SI_18_), .ZN(n15716) );
  INV_X1 U10189 ( .A(SI_12_), .ZN(n15728) );
  INV_X1 U10190 ( .A(n13952), .ZN(n13966) );
  NAND2_X1 U10191 ( .A1(n13863), .A2(n13862), .ZN(n14412) );
  INV_X1 U10192 ( .A(n16097), .ZN(n16254) );
  NAND2_X1 U10193 ( .A1(n14644), .A2(n10135), .ZN(n14622) );
  NAND2_X1 U10194 ( .A1(n14740), .A2(n14709), .ZN(n14734) );
  INV_X1 U10195 ( .A(n14740), .ZN(n16584) );
  INV_X1 U10196 ( .A(n14564), .ZN(n14769) );
  NAND2_X1 U10197 ( .A1(n12115), .A2(n14709), .ZN(n14785) );
  INV_X1 U10198 ( .A(n16534), .ZN(n16585) );
  NAND2_X1 U10199 ( .A1(n16076), .A2(n16075), .ZN(n16080) );
  INV_X1 U10200 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n14817) );
  INV_X1 U10201 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10340) );
  INV_X1 U10202 ( .A(n16364), .ZN(n14978) );
  INV_X1 U10203 ( .A(n12333), .ZN(n15462) );
  INV_X1 U10204 ( .A(n15435), .ZN(n15274) );
  INV_X1 U10205 ( .A(n12713), .ZN(n14960) );
  NOR2_X1 U10206 ( .A1(n10441), .A2(n10258), .ZN(n14964) );
  INV_X1 U10207 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n16363) );
  INV_X1 U10208 ( .A(n15065), .ZN(n16358) );
  NAND2_X1 U10209 ( .A1(n15338), .A2(n10478), .ZN(n15310) );
  INV_X1 U10210 ( .A(n15338), .ZN(n15295) );
  INV_X1 U10211 ( .A(n15345), .ZN(n15177) );
  AND2_X2 U10212 ( .A1(n10476), .A2(n10534), .ZN(n16553) );
  AND2_X1 U10213 ( .A1(n16550), .A2(n16549), .ZN(n16555) );
  INV_X1 U10214 ( .A(n16556), .ZN(n16554) );
  AND2_X2 U10215 ( .A1(n10535), .A2(n10534), .ZN(n16556) );
  INV_X1 U10216 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10700) );
  INV_X1 U10217 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10287) );
  NOR2_X1 U10218 ( .A1(n10272), .A2(P2_U3088), .ZN(P2_U3947) );
  NOR2_X1 U10219 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), 
        .ZN(n8532) );
  NOR2_X1 U10220 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), 
        .ZN(n8531) );
  NAND4_X1 U10221 ( .A1(n8532), .A2(n8531), .A3(n9053), .A4(n9091), .ZN(n8533)
         );
  NAND2_X1 U10222 ( .A1(n8538), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8539) );
  NAND2_X1 U10223 ( .A1(n8950), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8545) );
  AND2_X2 U10224 ( .A1(n13071), .A2(n13748), .ZN(n8951) );
  NAND2_X1 U10225 ( .A1(n8951), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8544) );
  INV_X1 U10226 ( .A(n13071), .ZN(n8541) );
  AND2_X2 U10227 ( .A1(n8541), .A2(n13748), .ZN(n8631) );
  NAND2_X1 U10228 ( .A1(n8631), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8543) );
  NAND2_X1 U10229 ( .A1(n8718), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8542) );
  INV_X2 U10230 ( .A(n10029), .ZN(n10196) );
  INV_X1 U10231 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U10232 ( .A1(n8562), .A2(n8568), .ZN(n8551) );
  NAND2_X1 U10233 ( .A1(n10172), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8550) );
  NAND2_X1 U10234 ( .A1(n8551), .A2(n8550), .ZN(n8581) );
  NAND2_X1 U10235 ( .A1(n10181), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8582) );
  NAND2_X1 U10236 ( .A1(n10229), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8552) );
  AND2_X1 U10237 ( .A1(n8582), .A2(n8552), .ZN(n8580) );
  XNOR2_X1 U10238 ( .A(n8581), .B(n8580), .ZN(n10184) );
  OR2_X1 U10239 ( .A1(n9027), .A2(n10184), .ZN(n8557) );
  INV_X1 U10241 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8638) );
  INV_X1 U10242 ( .A(n13017), .ZN(n8575) );
  NAND2_X1 U10243 ( .A1(n8950), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U10244 ( .A1(n8951), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8560) );
  NAND2_X1 U10245 ( .A1(n8631), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8559) );
  NAND2_X1 U10246 ( .A1(n8718), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8558) );
  INV_X1 U10247 ( .A(n11228), .ZN(n13751) );
  XNOR2_X1 U10248 ( .A(n8562), .B(n8568), .ZN(n8563) );
  MUX2_X1 U10249 ( .A(n8563), .B(SI_1_), .S(n10171), .Z(n13752) );
  MUX2_X1 U10250 ( .A(n13751), .B(n13752), .S(n10927), .Z(n10623) );
  NAND2_X1 U10251 ( .A1(n8573), .A2(n10623), .ZN(n12857) );
  INV_X1 U10252 ( .A(n10623), .ZN(n16368) );
  NAND2_X1 U10253 ( .A1(n13227), .A2(n16368), .ZN(n12858) );
  NAND2_X1 U10254 ( .A1(n8951), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8567) );
  NAND2_X1 U10255 ( .A1(n8950), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U10256 ( .A1(n8718), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8564) );
  INV_X1 U10257 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10177) );
  INV_X1 U10258 ( .A(n8568), .ZN(n8570) );
  INV_X1 U10259 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9297) );
  NAND2_X1 U10260 ( .A1(n9297), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8569) );
  AND2_X1 U10261 ( .A1(n8570), .A2(n8569), .ZN(n10176) );
  INV_X1 U10262 ( .A(SI_0_), .ZN(n10175) );
  OR2_X1 U10263 ( .A1(n7461), .A2(n10175), .ZN(n8571) );
  INV_X1 U10264 ( .A(n10691), .ZN(n10846) );
  NAND2_X1 U10265 ( .A1(n16370), .A2(n16371), .ZN(n16369) );
  NAND2_X1 U10266 ( .A1(n8573), .A2(n16368), .ZN(n11132) );
  NAND2_X1 U10267 ( .A1(n16369), .A2(n11132), .ZN(n8574) );
  NAND2_X1 U10268 ( .A1(n8950), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8579) );
  NAND2_X1 U10269 ( .A1(n8951), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8578) );
  INV_X1 U10270 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15756) );
  NAND2_X1 U10271 ( .A1(n8718), .A2(n15756), .ZN(n8576) );
  NAND2_X1 U10272 ( .A1(n8581), .A2(n8580), .ZN(n8583) );
  NAND2_X1 U10273 ( .A1(n8583), .A2(n8582), .ZN(n8586) );
  NAND2_X1 U10274 ( .A1(n10179), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8599) );
  NAND2_X1 U10275 ( .A1(n10198), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8584) );
  NAND2_X1 U10276 ( .A1(n8586), .A2(n8585), .ZN(n8600) );
  OR2_X1 U10277 ( .A1(n8586), .A2(n8585), .ZN(n8587) );
  NAND2_X1 U10278 ( .A1(n8600), .A2(n8587), .ZN(n10186) );
  OR2_X1 U10279 ( .A1(n9027), .A2(n10186), .ZN(n8590) );
  XNOR2_X1 U10280 ( .A(n8588), .B(P3_IR_REG_3__SCAN_IN), .ZN(n11008) );
  OR2_X1 U10281 ( .A1(n10927), .A2(n11008), .ZN(n8589) );
  NAND2_X1 U10282 ( .A1(n11590), .A2(n16422), .ZN(n12871) );
  INV_X1 U10283 ( .A(n11590), .ZN(n13225) );
  INV_X1 U10284 ( .A(n16422), .ZN(n11084) );
  NAND2_X1 U10285 ( .A1(n13225), .A2(n11084), .ZN(n12870) );
  AND2_X1 U10286 ( .A1(n16373), .A2(n8592), .ZN(n11304) );
  NOR2_X1 U10287 ( .A1(n13018), .A2(n11304), .ZN(n8593) );
  NAND2_X1 U10288 ( .A1(n11131), .A2(n8593), .ZN(n11307) );
  OR2_X1 U10289 ( .A1(n11590), .A2(n11084), .ZN(n8594) );
  NAND2_X1 U10290 ( .A1(n11307), .A2(n8594), .ZN(n11589) );
  NAND2_X1 U10291 ( .A1(n8950), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8598) );
  NAND2_X1 U10292 ( .A1(n8951), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8597) );
  OR2_X1 U10293 ( .A1(n8512), .A2(n8610), .ZN(n11596) );
  NAND2_X1 U10294 ( .A1(n8718), .A2(n11596), .ZN(n8596) );
  NAND2_X1 U10295 ( .A1(n8631), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8595) );
  OR2_X1 U10296 ( .A1(n8616), .A2(SI_4_), .ZN(n8607) );
  NAND2_X1 U10297 ( .A1(n10193), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8619) );
  NAND2_X1 U10298 ( .A1(n10223), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8601) );
  XNOR2_X1 U10299 ( .A(n8618), .B(n8617), .ZN(n10190) );
  OR2_X1 U10300 ( .A1(n9027), .A2(n10190), .ZN(n8606) );
  NAND2_X1 U10301 ( .A1(n7591), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8602) );
  MUX2_X1 U10302 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8602), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n8604) );
  INV_X1 U10303 ( .A(n7525), .ZN(n8603) );
  OR2_X1 U10304 ( .A1(n10927), .A2(n11015), .ZN(n8605) );
  NAND2_X1 U10306 ( .A1(n11650), .A2(n16437), .ZN(n12877) );
  INV_X1 U10307 ( .A(n11650), .ZN(n13224) );
  INV_X1 U10308 ( .A(n16437), .ZN(n11475) );
  NAND2_X1 U10309 ( .A1(n13224), .A2(n11475), .ZN(n12876) );
  NAND2_X1 U10310 ( .A1(n11589), .A2(n8362), .ZN(n8609) );
  OR2_X1 U10311 ( .A1(n11650), .A2(n11475), .ZN(n8608) );
  NAND2_X1 U10312 ( .A1(n8609), .A2(n8608), .ZN(n11515) );
  NAND2_X1 U10313 ( .A1(n8950), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U10314 ( .A1(n8951), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8614) );
  NAND2_X1 U10315 ( .A1(n8610), .A2(n15774), .ZN(n8629) );
  OR2_X1 U10316 ( .A1(n8610), .A2(n15774), .ZN(n8611) );
  NAND2_X1 U10317 ( .A1(n8629), .A2(n8611), .ZN(n11643) );
  NAND2_X1 U10318 ( .A1(n8718), .A2(n11643), .ZN(n8613) );
  NAND2_X1 U10319 ( .A1(n8631), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8612) );
  OR2_X1 U10320 ( .A1(n8616), .A2(SI_5_), .ZN(n8628) );
  NAND2_X1 U10321 ( .A1(n8618), .A2(n8617), .ZN(n8620) );
  NAND2_X1 U10322 ( .A1(n10206), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8641) );
  NAND2_X1 U10323 ( .A1(n10225), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8621) );
  OR2_X1 U10324 ( .A1(n8623), .A2(n8622), .ZN(n8624) );
  NAND2_X1 U10325 ( .A1(n8642), .A2(n8624), .ZN(n10188) );
  OR2_X1 U10326 ( .A1(n9027), .A2(n10188), .ZN(n8627) );
  OR2_X1 U10327 ( .A1(n7525), .A2(n8638), .ZN(n8625) );
  XNOR2_X1 U10328 ( .A(n8625), .B(P3_IR_REG_5__SCAN_IN), .ZN(n11029) );
  OR2_X1 U10329 ( .A1(n10927), .A2(n11029), .ZN(n8626) );
  NAND2_X1 U10330 ( .A1(n11805), .A2(n16456), .ZN(n12880) );
  INV_X1 U10331 ( .A(n11805), .ZN(n13223) );
  INV_X1 U10332 ( .A(n16456), .ZN(n8646) );
  NAND2_X1 U10333 ( .A1(n13223), .A2(n8646), .ZN(n12881) );
  NAND2_X1 U10334 ( .A1(n8950), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8635) );
  NAND2_X1 U10335 ( .A1(n8951), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8634) );
  NAND2_X1 U10336 ( .A1(n8629), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8630) );
  NAND2_X1 U10337 ( .A1(n8649), .A2(n8630), .ZN(n11813) );
  NAND2_X1 U10338 ( .A1(n8718), .A2(n11813), .ZN(n8633) );
  NAND2_X1 U10339 ( .A1(n8631), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8632) );
  NAND4_X1 U10340 ( .A1(n8635), .A2(n8634), .A3(n8633), .A4(n8632), .ZN(n13222) );
  NOR2_X1 U10341 ( .A1(n8636), .A2(n8638), .ZN(n8637) );
  MUX2_X1 U10342 ( .A(n8638), .B(n8637), .S(P3_IR_REG_6__SCAN_IN), .Z(n8640)
         );
  INV_X1 U10343 ( .A(SI_6_), .ZN(n10169) );
  OR2_X1 U10344 ( .A1(n8616), .A2(n10169), .ZN(n8645) );
  XNOR2_X1 U10345 ( .A(n10215), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8643) );
  XNOR2_X1 U10346 ( .A(n8656), .B(n8643), .ZN(n10170) );
  OR2_X1 U10347 ( .A1(n9027), .A2(n10170), .ZN(n8644) );
  OAI211_X1 U10348 ( .C1(n10927), .C2(n11418), .A(n8645), .B(n8644), .ZN(
        n16470) );
  XNOR2_X1 U10349 ( .A(n13222), .B(n16470), .ZN(n13023) );
  AND2_X1 U10350 ( .A1(n11805), .A2(n8646), .ZN(n11807) );
  NOR2_X1 U10351 ( .A1(n13023), .A2(n11807), .ZN(n8647) );
  NAND2_X1 U10352 ( .A1(n13222), .A2(n16470), .ZN(n8648) );
  NAND2_X1 U10353 ( .A1(n8950), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8654) );
  NAND2_X1 U10354 ( .A1(n8951), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8653) );
  AND2_X1 U10355 ( .A1(n8649), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8650) );
  OR2_X1 U10356 ( .A1(n8650), .A2(n8663), .ZN(n11883) );
  NAND2_X1 U10357 ( .A1(n8718), .A2(n11883), .ZN(n8652) );
  NAND2_X1 U10358 ( .A1(n8631), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8651) );
  NAND4_X1 U10359 ( .A1(n8654), .A2(n8653), .A3(n8652), .A4(n8651), .ZN(n13221) );
  OR2_X1 U10360 ( .A1(n8616), .A2(SI_7_), .ZN(n8661) );
  NAND2_X1 U10361 ( .A1(n10211), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8655) );
  NAND2_X1 U10362 ( .A1(n10222), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8674) );
  NAND2_X1 U10363 ( .A1(n10220), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8657) );
  XNOR2_X1 U10364 ( .A(n8673), .B(n8671), .ZN(n10182) );
  OR2_X1 U10365 ( .A1(n9027), .A2(n10182), .ZN(n8660) );
  NAND2_X1 U10366 ( .A1(n8639), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8658) );
  XNOR2_X1 U10367 ( .A(n8658), .B(P3_IR_REG_7__SCAN_IN), .ZN(n11258) );
  OR2_X1 U10368 ( .A1(n10927), .A2(n11258), .ZN(n8659) );
  XNOR2_X1 U10369 ( .A(n13221), .B(n11924), .ZN(n12888) );
  NAND2_X1 U10370 ( .A1(n13221), .A2(n11924), .ZN(n8662) );
  NAND2_X1 U10371 ( .A1(n8951), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8668) );
  NAND2_X1 U10372 ( .A1(n8950), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8667) );
  NOR2_X1 U10373 ( .A1(n8663), .A2(n11267), .ZN(n8664) );
  OR2_X1 U10374 ( .A1(n8682), .A2(n8664), .ZN(n11983) );
  NAND2_X1 U10375 ( .A1(n8718), .A2(n11983), .ZN(n8666) );
  NAND2_X1 U10376 ( .A1(n13000), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8665) );
  NAND4_X1 U10377 ( .A1(n8668), .A2(n8667), .A3(n8666), .A4(n8665), .ZN(n13220) );
  NAND2_X1 U10378 ( .A1(n8688), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8670) );
  XNOR2_X1 U10379 ( .A(n8670), .B(n8669), .ZN(n11431) );
  INV_X1 U10380 ( .A(SI_8_), .ZN(n10173) );
  OR2_X1 U10381 ( .A1(n7461), .A2(n10173), .ZN(n8680) );
  INV_X1 U10382 ( .A(n8671), .ZN(n8672) );
  NAND2_X1 U10383 ( .A1(n10232), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8690) );
  NAND2_X1 U10384 ( .A1(n10237), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8675) );
  OR2_X1 U10385 ( .A1(n8677), .A2(n8676), .ZN(n8678) );
  NAND2_X1 U10386 ( .A1(n8691), .A2(n8678), .ZN(n10174) );
  OR2_X1 U10387 ( .A1(n9027), .A2(n10174), .ZN(n8679) );
  OAI211_X1 U10388 ( .C1(n10927), .C2(n11431), .A(n8680), .B(n8679), .ZN(
        n11984) );
  XNOR2_X1 U10389 ( .A(n13220), .B(n11984), .ZN(n13022) );
  INV_X1 U10390 ( .A(n11984), .ZN(n16485) );
  NAND2_X1 U10391 ( .A1(n12124), .A2(n16485), .ZN(n8681) );
  NAND2_X1 U10392 ( .A1(n8951), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8687) );
  NAND2_X1 U10393 ( .A1(n13000), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8686) );
  OR2_X1 U10394 ( .A1(n8682), .A2(n15782), .ZN(n8683) );
  NAND2_X1 U10395 ( .A1(n8700), .A2(n8683), .ZN(n12128) );
  NAND2_X1 U10396 ( .A1(n8718), .A2(n12128), .ZN(n8685) );
  NAND2_X1 U10397 ( .A1(n8950), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8684) );
  NAND4_X1 U10398 ( .A1(n8687), .A2(n8686), .A3(n8685), .A4(n8684), .ZN(n13219) );
  NAND2_X1 U10399 ( .A1(n8712), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8689) );
  XNOR2_X1 U10400 ( .A(n8689), .B(P3_IR_REG_9__SCAN_IN), .ZN(n11439) );
  OR2_X1 U10401 ( .A1(n8616), .A2(SI_9_), .ZN(n8697) );
  NAND2_X1 U10402 ( .A1(n10241), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8706) );
  NAND2_X1 U10403 ( .A1(n10240), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8692) );
  OR2_X1 U10404 ( .A1(n8694), .A2(n8693), .ZN(n8695) );
  AND2_X1 U10405 ( .A1(n8707), .A2(n8695), .ZN(n10194) );
  OR2_X1 U10406 ( .A1(n9027), .A2(n10194), .ZN(n8696) );
  OAI211_X1 U10407 ( .C1(n11439), .C2(n10927), .A(n8697), .B(n8696), .ZN(
        n16498) );
  INV_X1 U10408 ( .A(n16498), .ZN(n12127) );
  NAND2_X1 U10409 ( .A1(n13219), .A2(n12127), .ZN(n8698) );
  NAND2_X1 U10410 ( .A1(n12323), .A2(n16498), .ZN(n8699) );
  NAND2_X1 U10411 ( .A1(n8951), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8705) );
  NAND2_X1 U10412 ( .A1(n8631), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U10413 ( .A1(n8700), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8701) );
  NAND2_X1 U10414 ( .A1(n8719), .A2(n8701), .ZN(n12080) );
  NAND2_X1 U10415 ( .A1(n8718), .A2(n12080), .ZN(n8703) );
  NAND2_X1 U10416 ( .A1(n8950), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8702) );
  NAND2_X1 U10417 ( .A1(n10248), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8725) );
  NAND2_X1 U10418 ( .A1(n10247), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8708) );
  OR2_X1 U10419 ( .A1(n8710), .A2(n8709), .ZN(n8711) );
  AND2_X1 U10420 ( .A1(n8726), .A2(n8711), .ZN(n10209) );
  OR2_X1 U10421 ( .A1(n9027), .A2(n10209), .ZN(n8716) );
  OR2_X1 U10422 ( .A1(n8616), .A2(SI_10_), .ZN(n8715) );
  OR2_X1 U10423 ( .A1(n8732), .A2(n8638), .ZN(n8713) );
  XNOR2_X1 U10424 ( .A(n8731), .B(n8713), .ZN(n12006) );
  INV_X1 U10425 ( .A(n12006), .ZN(n11850) );
  OR2_X1 U10426 ( .A1(n10927), .A2(n11850), .ZN(n8714) );
  NAND2_X1 U10427 ( .A1(n12416), .A2(n12326), .ZN(n12904) );
  INV_X1 U10428 ( .A(n12416), .ZN(n13218) );
  NAND2_X1 U10429 ( .A1(n13218), .A2(n16513), .ZN(n12903) );
  NAND2_X1 U10430 ( .A1(n12904), .A2(n12903), .ZN(n13024) );
  OR2_X1 U10431 ( .A1(n12416), .A2(n16513), .ZN(n8717) );
  NAND2_X1 U10432 ( .A1(n8951), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8724) );
  NAND2_X1 U10433 ( .A1(n8950), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U10434 ( .A1(n8719), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8720) );
  NAND2_X1 U10435 ( .A1(n8753), .A2(n8720), .ZN(n12419) );
  NAND2_X1 U10436 ( .A1(n8718), .A2(n12419), .ZN(n8722) );
  NAND2_X1 U10437 ( .A1(n8631), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8721) );
  NAND4_X1 U10438 ( .A1(n8724), .A2(n8723), .A3(n8722), .A4(n8721), .ZN(n13217) );
  INV_X1 U10439 ( .A(n13217), .ZN(n12920) );
  NAND2_X1 U10440 ( .A1(n10250), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8740) );
  NAND2_X1 U10441 ( .A1(n10255), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8727) );
  OR2_X1 U10442 ( .A1(n8729), .A2(n8728), .ZN(n8730) );
  NAND2_X1 U10443 ( .A1(n8741), .A2(n8730), .ZN(n10207) );
  NAND2_X1 U10444 ( .A1(n12997), .A2(n10207), .ZN(n8736) );
  OR2_X1 U10445 ( .A1(n8616), .A2(SI_11_), .ZN(n8735) );
  NAND2_X1 U10446 ( .A1(n8732), .A2(n8731), .ZN(n8746) );
  NAND2_X1 U10447 ( .A1(n8746), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8733) );
  XNOR2_X1 U10448 ( .A(n8733), .B(P3_IR_REG_11__SCAN_IN), .ZN(n12196) );
  OR2_X1 U10449 ( .A1(n10927), .A2(n12196), .ZN(n8734) );
  INV_X1 U10450 ( .A(n12919), .ZN(n16536) );
  NAND2_X1 U10451 ( .A1(n12920), .A2(n16536), .ZN(n8737) );
  NAND2_X1 U10452 ( .A1(n12240), .A2(n8737), .ZN(n8739) );
  NAND2_X1 U10453 ( .A1(n13217), .A2(n12919), .ZN(n8738) );
  NAND2_X1 U10454 ( .A1(n10287), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8761) );
  NAND2_X1 U10455 ( .A1(n10291), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8742) );
  OR2_X1 U10456 ( .A1(n8744), .A2(n8743), .ZN(n8745) );
  NAND2_X1 U10457 ( .A1(n8762), .A2(n8745), .ZN(n10216) );
  NAND2_X1 U10458 ( .A1(n10216), .A2(n12997), .ZN(n8750) );
  INV_X1 U10459 ( .A(n8616), .ZN(n8885) );
  NAND2_X1 U10460 ( .A1(n8767), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8748) );
  INV_X1 U10461 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8747) );
  XNOR2_X1 U10462 ( .A(n8748), .B(n8747), .ZN(n12294) );
  AOI22_X1 U10463 ( .A1(n8885), .A2(n15728), .B1(n7613), .B2(n12294), .ZN(
        n8749) );
  NAND2_X1 U10464 ( .A1(n9010), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U10465 ( .A1(n13000), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8751) );
  AND2_X1 U10466 ( .A1(n8752), .A2(n8751), .ZN(n8757) );
  OR2_X1 U10467 ( .A1(n8509), .A2(n8772), .ZN(n12547) );
  NAND2_X1 U10468 ( .A1(n8718), .A2(n12547), .ZN(n8755) );
  NAND2_X1 U10469 ( .A1(n9009), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8754) );
  AND2_X1 U10470 ( .A1(n8755), .A2(n8754), .ZN(n8756) );
  NAND2_X1 U10471 ( .A1(n16559), .A2(n13157), .ZN(n8758) );
  NAND2_X1 U10472 ( .A1(n12392), .A2(n8758), .ZN(n8760) );
  NAND2_X1 U10473 ( .A1(n13216), .A2(n12546), .ZN(n8759) );
  NAND2_X1 U10474 ( .A1(n8765), .A2(n10340), .ZN(n8766) );
  NAND2_X1 U10475 ( .A1(n8782), .A2(n8766), .ZN(n10244) );
  NAND2_X1 U10476 ( .A1(n10244), .A2(n12997), .ZN(n8770) );
  OR2_X1 U10477 ( .A1(n8788), .A2(n8638), .ZN(n8768) );
  INV_X1 U10478 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8787) );
  XNOR2_X1 U10479 ( .A(n8768), .B(n8787), .ZN(n13234) );
  AOI22_X1 U10480 ( .A1(n8885), .A2(n15724), .B1(n7613), .B2(n13234), .ZN(
        n8769) );
  NAND2_X1 U10481 ( .A1(n9009), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U10482 ( .A1(n9010), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8776) );
  INV_X1 U10483 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8771) );
  OR2_X1 U10484 ( .A1(n8772), .A2(n8771), .ZN(n8773) );
  NAND2_X1 U10485 ( .A1(n8796), .A2(n8773), .ZN(n13159) );
  NAND2_X1 U10486 ( .A1(n8718), .A2(n13159), .ZN(n8775) );
  NAND2_X1 U10487 ( .A1(n13000), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8774) );
  NAND4_X1 U10488 ( .A1(n8777), .A2(n8776), .A3(n8775), .A4(n8774), .ZN(n13215) );
  NAND2_X1 U10489 ( .A1(n13659), .A2(n12543), .ZN(n8778) );
  NAND2_X1 U10490 ( .A1(n12473), .A2(n8778), .ZN(n8780) );
  OR2_X1 U10491 ( .A1(n13659), .A2(n12543), .ZN(n8779) );
  NAND2_X1 U10492 ( .A1(n10403), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8803) );
  NAND2_X1 U10493 ( .A1(n10402), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8783) );
  OR2_X1 U10494 ( .A1(n8785), .A2(n8784), .ZN(n8786) );
  NAND2_X1 U10495 ( .A1(n8804), .A2(n8786), .ZN(n10260) );
  NAND2_X1 U10496 ( .A1(n10260), .A2(n12997), .ZN(n8795) );
  NOR2_X1 U10497 ( .A1(n8792), .A2(n8638), .ZN(n8789) );
  MUX2_X1 U10498 ( .A(n8638), .B(n8789), .S(P3_IR_REG_14__SCAN_IN), .Z(n8790)
         );
  INV_X1 U10499 ( .A(n8790), .ZN(n8793) );
  INV_X1 U10500 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8791) );
  NAND2_X1 U10501 ( .A1(n8792), .A2(n8791), .ZN(n8826) );
  NAND2_X1 U10502 ( .A1(n8793), .A2(n8826), .ZN(n13268) );
  AOI22_X1 U10503 ( .A1(n13268), .A2(n7613), .B1(n8885), .B2(n15525), .ZN(
        n8794) );
  NAND2_X1 U10504 ( .A1(n9009), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8801) );
  NAND2_X1 U10505 ( .A1(n9010), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8800) );
  NAND2_X1 U10506 ( .A1(n8796), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8797) );
  NAND2_X1 U10507 ( .A1(n8813), .A2(n8797), .ZN(n12499) );
  NAND2_X1 U10508 ( .A1(n8718), .A2(n12499), .ZN(n8799) );
  NAND2_X1 U10509 ( .A1(n13000), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8798) );
  NAND4_X1 U10510 ( .A1(n8801), .A2(n8800), .A3(n8799), .A4(n8798), .ZN(n13214) );
  NOR2_X1 U10511 ( .A1(n13730), .A2(n13214), .ZN(n9077) );
  INV_X1 U10512 ( .A(n9077), .ZN(n12926) );
  NAND2_X1 U10513 ( .A1(n13730), .A2(n13214), .ZN(n12927) );
  INV_X1 U10514 ( .A(n13214), .ZN(n13583) );
  OR2_X1 U10515 ( .A1(n13730), .A2(n13583), .ZN(n8802) );
  NAND2_X1 U10516 ( .A1(n10467), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8820) );
  NAND2_X1 U10517 ( .A1(n12091), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8805) );
  OR2_X1 U10518 ( .A1(n8807), .A2(n8806), .ZN(n8808) );
  NAND2_X1 U10519 ( .A1(n8821), .A2(n8808), .ZN(n10262) );
  NAND2_X1 U10520 ( .A1(n10262), .A2(n12997), .ZN(n8812) );
  NAND2_X1 U10521 ( .A1(n8826), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8809) );
  OAI22_X1 U10522 ( .A1(n13292), .A2(n10927), .B1(n8616), .B2(SI_15_), .ZN(
        n8810) );
  INV_X1 U10523 ( .A(n8810), .ZN(n8811) );
  NAND2_X1 U10524 ( .A1(n9010), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8818) );
  NAND2_X1 U10525 ( .A1(n9009), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8817) );
  AND2_X1 U10526 ( .A1(n8813), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8814) );
  OR2_X1 U10527 ( .A1(n8814), .A2(n8834), .ZN(n13585) );
  NAND2_X1 U10528 ( .A1(n8718), .A2(n13585), .ZN(n8816) );
  NAND2_X1 U10529 ( .A1(n13000), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8815) );
  NAND4_X1 U10530 ( .A1(n8818), .A2(n8817), .A3(n8816), .A4(n8815), .ZN(n13213) );
  NAND2_X1 U10531 ( .A1(n13726), .A2(n13213), .ZN(n8819) );
  NAND2_X1 U10532 ( .A1(n12929), .A2(n8819), .ZN(n13575) );
  INV_X1 U10533 ( .A(n13213), .ZN(n13568) );
  NAND2_X1 U10534 ( .A1(n13726), .A2(n13568), .ZN(n13563) );
  NAND2_X1 U10535 ( .A1(n13577), .A2(n13563), .ZN(n8841) );
  NAND2_X1 U10536 ( .A1(n10632), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8842) );
  INV_X1 U10537 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10631) );
  NAND2_X1 U10538 ( .A1(n10631), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8822) );
  OR2_X1 U10539 ( .A1(n8824), .A2(n8823), .ZN(n8825) );
  NAND2_X1 U10540 ( .A1(n8843), .A2(n8825), .ZN(n10301) );
  OR2_X1 U10541 ( .A1(n10301), .A2(n9027), .ZN(n8833) );
  NAND2_X1 U10542 ( .A1(n8827), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8830) );
  INV_X1 U10543 ( .A(n8830), .ZN(n8828) );
  NAND2_X1 U10544 ( .A1(n8828), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n8831) );
  NAND2_X1 U10545 ( .A1(n8830), .A2(n8829), .ZN(n8848) );
  AOI22_X1 U10546 ( .A1(n13296), .A2(n7613), .B1(SI_16_), .B2(n8885), .ZN(
        n8832) );
  NAND2_X1 U10547 ( .A1(n8833), .A2(n8832), .ZN(n13118) );
  NAND2_X1 U10548 ( .A1(n9009), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8839) );
  NAND2_X1 U10549 ( .A1(n9010), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8838) );
  INV_X1 U10550 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n15773) );
  NOR2_X1 U10551 ( .A1(n8834), .A2(n15773), .ZN(n8835) );
  OR2_X1 U10552 ( .A1(n8853), .A2(n8835), .ZN(n13570) );
  NAND2_X1 U10553 ( .A1(n8718), .A2(n13570), .ZN(n8837) );
  NAND2_X1 U10554 ( .A1(n13000), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8836) );
  NAND4_X1 U10555 ( .A1(n8839), .A2(n8838), .A3(n8837), .A4(n8836), .ZN(n13212) );
  OR2_X1 U10556 ( .A1(n13118), .A2(n13212), .ZN(n12934) );
  NAND2_X1 U10557 ( .A1(n13118), .A2(n13212), .ZN(n12933) );
  NAND2_X1 U10558 ( .A1(n12934), .A2(n12933), .ZN(n13564) );
  INV_X1 U10559 ( .A(n13564), .ZN(n8840) );
  NAND2_X1 U10560 ( .A1(n10700), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8860) );
  NAND2_X1 U10561 ( .A1(n10698), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8844) );
  OR2_X1 U10562 ( .A1(n8846), .A2(n8845), .ZN(n8847) );
  NAND2_X1 U10563 ( .A1(n8861), .A2(n8847), .ZN(n10362) );
  NAND2_X1 U10564 ( .A1(n10362), .A2(n12997), .ZN(n8852) );
  NAND2_X1 U10565 ( .A1(n8848), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8849) );
  XNOR2_X1 U10566 ( .A(n8849), .B(P3_IR_REG_17__SCAN_IN), .ZN(n13328) );
  OAI22_X1 U10567 ( .A1(n13328), .A2(n10927), .B1(SI_17_), .B2(n7461), .ZN(
        n8850) );
  INV_X1 U10568 ( .A(n8850), .ZN(n8851) );
  NAND2_X1 U10569 ( .A1(n9010), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8858) );
  NAND2_X1 U10570 ( .A1(n9009), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8857) );
  INV_X1 U10571 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n15575) );
  OR2_X1 U10572 ( .A1(n8853), .A2(n15575), .ZN(n8854) );
  NAND2_X1 U10573 ( .A1(n8870), .A2(n8854), .ZN(n13551) );
  NAND2_X1 U10574 ( .A1(n8718), .A2(n13551), .ZN(n8856) );
  NAND2_X1 U10575 ( .A1(n13000), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8855) );
  XNOR2_X1 U10576 ( .A(n13644), .B(n13569), .ZN(n13557) );
  INV_X1 U10577 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11395) );
  NAND2_X1 U10578 ( .A1(n11395), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8878) );
  INV_X1 U10579 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11394) );
  NAND2_X1 U10580 ( .A1(n11394), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8862) );
  OR2_X1 U10581 ( .A1(n8864), .A2(n8863), .ZN(n8865) );
  NAND2_X1 U10582 ( .A1(n8879), .A2(n8865), .ZN(n10419) );
  OR2_X1 U10583 ( .A1(n10419), .A2(n9027), .ZN(n8869) );
  NAND2_X1 U10584 ( .A1(n8866), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8867) );
  XNOR2_X1 U10585 ( .A(n8867), .B(P3_IR_REG_18__SCAN_IN), .ZN(n13353) );
  AOI22_X1 U10586 ( .A1(n8885), .A2(SI_18_), .B1(n7613), .B2(n13353), .ZN(
        n8868) );
  NAND2_X1 U10587 ( .A1(n8869), .A2(n8868), .ZN(n13171) );
  NAND2_X1 U10588 ( .A1(n9009), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8875) );
  NAND2_X1 U10589 ( .A1(n9010), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8874) );
  NAND2_X1 U10590 ( .A1(n8870), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8871) );
  NAND2_X1 U10591 ( .A1(n8888), .A2(n8871), .ZN(n13541) );
  NAND2_X1 U10592 ( .A1(n8718), .A2(n13541), .ZN(n8873) );
  NAND2_X1 U10593 ( .A1(n13000), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8872) );
  OR2_X1 U10594 ( .A1(n13171), .A2(n13548), .ZN(n12946) );
  NAND2_X1 U10595 ( .A1(n13171), .A2(n13548), .ZN(n12944) );
  NOR2_X1 U10596 ( .A1(n13644), .A2(n13569), .ZN(n13536) );
  NOR2_X1 U10597 ( .A1(n13535), .A2(n13536), .ZN(n8876) );
  INV_X1 U10598 ( .A(n13548), .ZN(n13210) );
  OR2_X1 U10599 ( .A1(n13171), .A2(n13210), .ZN(n8877) );
  INV_X1 U10600 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n12591) );
  NAND2_X1 U10601 ( .A1(n12591), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8897) );
  INV_X1 U10602 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12786) );
  NAND2_X1 U10603 ( .A1(n12786), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8880) );
  OR2_X1 U10604 ( .A1(n8882), .A2(n8881), .ZN(n8883) );
  NAND2_X1 U10605 ( .A1(n8898), .A2(n8883), .ZN(n10466) );
  OR2_X1 U10606 ( .A1(n10466), .A2(n9027), .ZN(n8887) );
  NAND2_X1 U10607 ( .A1(n7543), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8884) );
  AOI22_X1 U10608 ( .A1(n8885), .A2(SI_19_), .B1(n7613), .B2(n13369), .ZN(
        n8886) );
  AND2_X1 U10609 ( .A1(n8888), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8889) );
  OR2_X1 U10610 ( .A1(n8889), .A2(n8907), .ZN(n13528) );
  NAND2_X1 U10611 ( .A1(n13528), .A2(n8718), .ZN(n8893) );
  NAND2_X1 U10612 ( .A1(n9009), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U10613 ( .A1(n9010), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8891) );
  NAND2_X1 U10614 ( .A1(n13000), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8890) );
  INV_X1 U10615 ( .A(n13540), .ZN(n13209) );
  NAND2_X1 U10616 ( .A1(n13085), .A2(n13209), .ZN(n8894) );
  OR2_X1 U10617 ( .A1(n13085), .A2(n13209), .ZN(n8895) );
  NAND2_X1 U10618 ( .A1(n8901), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8902) );
  NAND2_X1 U10619 ( .A1(n8914), .A2(n8902), .ZN(n10657) );
  OR2_X1 U10620 ( .A1(n8616), .A2(n10656), .ZN(n8903) );
  NAND2_X1 U10621 ( .A1(n9009), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8906) );
  NAND2_X1 U10622 ( .A1(n9010), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8905) );
  AND2_X1 U10623 ( .A1(n8906), .A2(n8905), .ZN(n8911) );
  INV_X1 U10624 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n15788) );
  OR2_X1 U10625 ( .A1(n8907), .A2(n15788), .ZN(n8908) );
  NAND2_X1 U10626 ( .A1(n15788), .A2(n8907), .ZN(n8919) );
  NAND2_X1 U10627 ( .A1(n8908), .A2(n8919), .ZN(n13518) );
  NAND2_X1 U10628 ( .A1(n13518), .A2(n8718), .ZN(n8910) );
  NAND2_X1 U10629 ( .A1(n13000), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8909) );
  OR2_X1 U10630 ( .A1(n13142), .A2(n13527), .ZN(n12952) );
  NAND2_X1 U10631 ( .A1(n13142), .A2(n13527), .ZN(n12953) );
  NAND2_X1 U10632 ( .A1(n12952), .A2(n12953), .ZN(n13037) );
  INV_X1 U10633 ( .A(n13037), .ZN(n13512) );
  INV_X1 U10634 ( .A(n13527), .ZN(n13501) );
  NAND2_X1 U10635 ( .A1(n13142), .A2(n13501), .ZN(n8912) );
  INV_X1 U10636 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11729) );
  NAND2_X1 U10637 ( .A1(n11729), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8928) );
  INV_X1 U10638 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n13778) );
  NAND2_X1 U10639 ( .A1(n13778), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8915) );
  NAND2_X1 U10640 ( .A1(n8928), .A2(n8915), .ZN(n8926) );
  XNOR2_X1 U10641 ( .A(n8927), .B(n8926), .ZN(n11067) );
  NAND2_X1 U10642 ( .A1(n11067), .A2(n12997), .ZN(n8917) );
  INV_X1 U10643 ( .A(SI_21_), .ZN(n11068) );
  OR2_X1 U10644 ( .A1(n7461), .A2(n11068), .ZN(n8916) );
  NAND2_X1 U10645 ( .A1(n9009), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8924) );
  NAND2_X1 U10646 ( .A1(n9010), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8923) );
  INV_X1 U10647 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n15761) );
  INV_X1 U10648 ( .A(n8919), .ZN(n8918) );
  NAND2_X1 U10649 ( .A1(P3_REG3_REG_21__SCAN_IN), .A2(n8919), .ZN(n8920) );
  NAND2_X1 U10650 ( .A1(n8939), .A2(n8920), .ZN(n13507) );
  NAND2_X1 U10651 ( .A1(n8718), .A2(n13507), .ZN(n8922) );
  NAND2_X1 U10652 ( .A1(n13000), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8921) );
  OR2_X1 U10653 ( .A1(n13702), .A2(n13479), .ZN(n12808) );
  NAND2_X1 U10654 ( .A1(n13702), .A2(n13479), .ZN(n12805) );
  NAND2_X1 U10655 ( .A1(n8925), .A2(n12805), .ZN(n13476) );
  INV_X1 U10656 ( .A(n13476), .ZN(n8945) );
  INV_X1 U10657 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8930) );
  NAND2_X1 U10658 ( .A1(n8930), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8946) );
  INV_X1 U10659 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n13787) );
  NAND2_X1 U10660 ( .A1(n13787), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8931) );
  AND2_X1 U10661 ( .A1(n8946), .A2(n8931), .ZN(n8932) );
  OR2_X1 U10662 ( .A1(n8933), .A2(n8932), .ZN(n8934) );
  NAND2_X1 U10663 ( .A1(n8947), .A2(n8934), .ZN(n11104) );
  INV_X1 U10664 ( .A(SI_22_), .ZN(n8935) );
  OR2_X1 U10665 ( .A1(n8616), .A2(n8935), .ZN(n8936) );
  NAND2_X1 U10666 ( .A1(n9009), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8944) );
  NAND2_X1 U10667 ( .A1(n9010), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8943) );
  INV_X1 U10668 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n15585) );
  NAND2_X1 U10669 ( .A1(n8939), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8940) );
  NAND2_X1 U10670 ( .A1(n8952), .A2(n8940), .ZN(n13487) );
  NAND2_X1 U10671 ( .A1(n8718), .A2(n13487), .ZN(n8942) );
  NAND2_X1 U10672 ( .A1(n8631), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8941) );
  INV_X1 U10673 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n13768) );
  XNOR2_X1 U10674 ( .A(n13768), .B(P2_DATAO_REG_23__SCAN_IN), .ZN(n8959) );
  XNOR2_X1 U10675 ( .A(n8960), .B(n8959), .ZN(n11313) );
  NAND2_X1 U10676 ( .A1(n11313), .A2(n12997), .ZN(n8949) );
  INV_X1 U10677 ( .A(SI_23_), .ZN(n11315) );
  NAND2_X1 U10678 ( .A1(n9009), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8957) );
  NAND2_X1 U10679 ( .A1(n9010), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8956) );
  NAND2_X1 U10680 ( .A1(n8952), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8953) );
  NAND2_X1 U10681 ( .A1(n8968), .A2(n8953), .ZN(n13470) );
  NAND2_X1 U10682 ( .A1(n8718), .A2(n13470), .ZN(n8955) );
  NAND4_X1 U10683 ( .A1(n8957), .A2(n8956), .A3(n8955), .A4(n8954), .ZN(n13478) );
  XNOR2_X1 U10684 ( .A(n13469), .B(n13478), .ZN(n12960) );
  NAND2_X1 U10685 ( .A1(n13469), .A2(n13478), .ZN(n8958) );
  INV_X1 U10686 ( .A(SI_24_), .ZN(n15705) );
  NAND2_X1 U10687 ( .A1(n13768), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8961) );
  INV_X1 U10688 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13813) );
  NAND2_X1 U10689 ( .A1(n8962), .A2(n13813), .ZN(n8963) );
  NAND2_X1 U10690 ( .A1(n8964), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8965) );
  NAND2_X1 U10691 ( .A1(n8976), .A2(n8965), .ZN(n8966) );
  MUX2_X1 U10692 ( .A(n15705), .B(n8966), .S(n10196), .Z(n11990) );
  NAND2_X1 U10693 ( .A1(n9009), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8973) );
  NAND2_X1 U10694 ( .A1(n9010), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8972) );
  INV_X1 U10695 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n15576) );
  NAND2_X1 U10696 ( .A1(n8968), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8969) );
  NAND2_X1 U10697 ( .A1(n8983), .A2(n8969), .ZN(n13449) );
  NAND2_X1 U10698 ( .A1(n8718), .A2(n13449), .ZN(n8971) );
  NAND2_X1 U10699 ( .A1(n13000), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8970) );
  XNOR2_X1 U10700 ( .A(n13687), .B(n13439), .ZN(n13447) );
  INV_X1 U10701 ( .A(n13447), .ZN(n13452) );
  NAND2_X1 U10702 ( .A1(n13687), .A2(n13439), .ZN(n8974) );
  INV_X1 U10703 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15917) );
  NAND2_X1 U10704 ( .A1(n15917), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8995) );
  NAND2_X1 U10705 ( .A1(n14817), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8977) );
  AND2_X1 U10706 ( .A1(n8995), .A2(n8977), .ZN(n8978) );
  OR2_X1 U10707 ( .A1(n8979), .A2(n8978), .ZN(n8980) );
  NAND2_X1 U10708 ( .A1(n8996), .A2(n8980), .ZN(n11923) );
  OR2_X1 U10709 ( .A1(n7461), .A2(n15704), .ZN(n8981) );
  NAND2_X1 U10710 ( .A1(n9009), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8988) );
  NAND2_X1 U10711 ( .A1(n9010), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8987) );
  NAND2_X1 U10712 ( .A1(n8983), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8984) );
  NAND2_X1 U10713 ( .A1(n9011), .A2(n8984), .ZN(n13442) );
  NAND2_X1 U10714 ( .A1(n8718), .A2(n13442), .ZN(n8986) );
  NAND2_X1 U10715 ( .A1(n13000), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8985) );
  NAND2_X1 U10716 ( .A1(n13104), .A2(n13453), .ZN(n13424) );
  OR2_X1 U10717 ( .A1(n13104), .A2(n13453), .ZN(n8989) );
  NAND2_X1 U10718 ( .A1(n13424), .A2(n8989), .ZN(n12841) );
  INV_X1 U10719 ( .A(n13453), .ZN(n13208) );
  NAND2_X1 U10720 ( .A1(n13104), .A2(n13208), .ZN(n8990) );
  NAND2_X1 U10721 ( .A1(n9009), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8994) );
  NAND2_X1 U10722 ( .A1(n9010), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8993) );
  XNOR2_X1 U10723 ( .A(n9011), .B(P3_REG3_REG_26__SCAN_IN), .ZN(n13429) );
  NAND2_X1 U10724 ( .A1(n8718), .A2(n13429), .ZN(n8992) );
  NAND2_X1 U10725 ( .A1(n13000), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8991) );
  INV_X1 U10726 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15913) );
  NAND2_X1 U10727 ( .A1(n15913), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9004) );
  INV_X1 U10728 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14811) );
  NAND2_X1 U10729 ( .A1(n14811), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8997) );
  AND2_X1 U10730 ( .A1(n9004), .A2(n8997), .ZN(n8998) );
  NAND2_X1 U10731 ( .A1(n9005), .A2(n9000), .ZN(n12043) );
  INV_X1 U10732 ( .A(SI_26_), .ZN(n15502) );
  OR2_X1 U10733 ( .A1(n8616), .A2(n15502), .ZN(n9001) );
  NAND2_X2 U10734 ( .A1(n9002), .A2(n9001), .ZN(n13179) );
  OR2_X1 U10735 ( .A1(n13207), .A2(n13179), .ZN(n9003) );
  INV_X1 U10736 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15910) );
  NAND2_X1 U10737 ( .A1(n15910), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9022) );
  INV_X1 U10738 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n14808) );
  NAND2_X1 U10739 ( .A1(n14808), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9006) );
  NAND2_X1 U10740 ( .A1(n9022), .A2(n9006), .ZN(n9019) );
  XNOR2_X1 U10741 ( .A(n9021), .B(n9019), .ZN(n12207) );
  NAND2_X1 U10742 ( .A1(n12207), .A2(n12997), .ZN(n9008) );
  INV_X1 U10743 ( .A(SI_27_), .ZN(n15700) );
  NAND2_X1 U10744 ( .A1(n9009), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9018) );
  NAND2_X1 U10745 ( .A1(n9010), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9017) );
  INV_X1 U10746 ( .A(n9011), .ZN(n9012) );
  INV_X1 U10747 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n15795) );
  NAND2_X1 U10748 ( .A1(n9012), .A2(n15795), .ZN(n9013) );
  NAND2_X1 U10749 ( .A1(n9013), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9014) );
  NAND2_X1 U10750 ( .A1(n9031), .A2(n9014), .ZN(n13408) );
  NAND2_X1 U10751 ( .A1(n8718), .A2(n13408), .ZN(n9016) );
  NAND2_X1 U10752 ( .A1(n8631), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9015) );
  OR2_X1 U10753 ( .A1(n13412), .A2(n13421), .ZN(n12844) );
  NAND2_X1 U10754 ( .A1(n13412), .A2(n13421), .ZN(n12848) );
  INV_X1 U10755 ( .A(n9019), .ZN(n9020) );
  NAND2_X1 U10756 ( .A1(n9021), .A2(n9020), .ZN(n9023) );
  NAND2_X1 U10757 ( .A1(n9023), .A2(n9022), .ZN(n9026) );
  INV_X1 U10758 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n12781) );
  NAND2_X1 U10759 ( .A1(n12781), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9038) );
  INV_X1 U10760 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14805) );
  NAND2_X1 U10761 ( .A1(n14805), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9024) );
  AND2_X1 U10762 ( .A1(n9038), .A2(n9024), .ZN(n9025) );
  INV_X1 U10763 ( .A(SI_28_), .ZN(n15498) );
  NAND2_X1 U10764 ( .A1(n9009), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9036) );
  NAND2_X1 U10765 ( .A1(n9010), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9035) );
  INV_X1 U10766 ( .A(n9031), .ZN(n9030) );
  INV_X1 U10767 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n15762) );
  NAND2_X1 U10768 ( .A1(n9030), .A2(n15762), .ZN(n13372) );
  NAND2_X1 U10769 ( .A1(n9031), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9032) );
  NAND2_X1 U10770 ( .A1(n13372), .A2(n9032), .ZN(n13396) );
  NAND2_X1 U10771 ( .A1(n8718), .A2(n13396), .ZN(n9034) );
  NAND2_X1 U10772 ( .A1(n8631), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9033) );
  NAND4_X1 U10773 ( .A1(n9036), .A2(n9035), .A3(n9034), .A4(n9033), .ZN(n13404) );
  NAND2_X1 U10774 ( .A1(n12978), .A2(n13404), .ZN(n9037) );
  INV_X1 U10775 ( .A(n13387), .ZN(n13390) );
  OR2_X1 U10776 ( .A1(n13412), .A2(n13392), .ZN(n13391) );
  NAND3_X1 U10777 ( .A1(n13403), .A2(n13390), .A3(n13391), .ZN(n13389) );
  NAND2_X1 U10778 ( .A1(n13389), .A2(n9037), .ZN(n9051) );
  NAND2_X1 U10779 ( .A1(n9039), .A2(n9038), .ZN(n12983) );
  XNOR2_X1 U10780 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n12982) );
  INV_X1 U10781 ( .A(n12982), .ZN(n9040) );
  XNOR2_X1 U10782 ( .A(n12983), .B(n9040), .ZN(n13747) );
  NAND2_X1 U10783 ( .A1(n13747), .A2(n12997), .ZN(n9042) );
  INV_X1 U10784 ( .A(SI_29_), .ZN(n15696) );
  OR2_X1 U10785 ( .A1(n8616), .A2(n15696), .ZN(n9041) );
  NAND2_X1 U10786 ( .A1(n9042), .A2(n9041), .ZN(n9047) );
  INV_X1 U10787 ( .A(n13372), .ZN(n9043) );
  NAND2_X1 U10788 ( .A1(n8718), .A2(n9043), .ZN(n13004) );
  NAND2_X1 U10789 ( .A1(n9010), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9046) );
  NAND2_X1 U10790 ( .A1(n8631), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9045) );
  NAND2_X1 U10791 ( .A1(n9009), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9044) );
  NAND2_X1 U10792 ( .A1(n9047), .A2(n12838), .ZN(n13048) );
  INV_X1 U10793 ( .A(n13048), .ZN(n9049) );
  INV_X1 U10794 ( .A(n12838), .ZN(n13393) );
  NAND2_X1 U10795 ( .A1(n13380), .A2(n13393), .ZN(n13051) );
  INV_X1 U10796 ( .A(n13051), .ZN(n9048) );
  XNOR2_X1 U10797 ( .A(n9051), .B(n9050), .ZN(n9068) );
  NAND2_X1 U10798 ( .A1(n9092), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9055) );
  NAND2_X1 U10799 ( .A1(n13064), .A2(n13369), .ZN(n9139) );
  NAND2_X1 U10800 ( .A1(n9056), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9057) );
  NAND2_X1 U10801 ( .A1(n9058), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9059) );
  NAND2_X1 U10802 ( .A1(n12855), .A2(n9138), .ZN(n13056) );
  INV_X1 U10803 ( .A(n13404), .ZN(n13076) );
  OR2_X1 U10804 ( .A1(n7728), .A2(n13357), .ZN(n10936) );
  NAND2_X1 U10805 ( .A1(n10927), .A2(n10936), .ZN(n10617) );
  INV_X1 U10806 ( .A(P3_B_REG_SCAN_IN), .ZN(n9061) );
  NOR2_X1 U10807 ( .A1(n7728), .A2(n9061), .ZN(n9062) );
  OR2_X1 U10808 ( .A1(n16372), .A2(n9062), .ZN(n13373) );
  NAND2_X1 U10809 ( .A1(n9009), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9065) );
  NAND2_X1 U10810 ( .A1(n9010), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9064) );
  NAND2_X1 U10811 ( .A1(n13000), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9063) );
  INV_X1 U10812 ( .A(n9066), .ZN(n9067) );
  NAND2_X1 U10813 ( .A1(n12863), .A2(n12867), .ZN(n11303) );
  NAND2_X1 U10814 ( .A1(n11512), .A2(n13015), .ZN(n11514) );
  NAND2_X1 U10815 ( .A1(n11514), .A2(n12880), .ZN(n11804) );
  NAND2_X1 U10816 ( .A1(n12884), .A2(n16470), .ZN(n9069) );
  NAND2_X1 U10817 ( .A1(n11978), .A2(n13022), .ZN(n11977) );
  NAND2_X1 U10818 ( .A1(n12124), .A2(n11984), .ZN(n12895) );
  NOR2_X1 U10819 ( .A1(n13219), .A2(n16498), .ZN(n12077) );
  INV_X1 U10820 ( .A(n12904), .ZN(n9072) );
  OR2_X1 U10821 ( .A1(n12077), .A2(n9072), .ZN(n12244) );
  NAND2_X1 U10822 ( .A1(n12920), .A2(n12919), .ZN(n12909) );
  INV_X1 U10823 ( .A(n12909), .ZN(n9074) );
  NAND2_X1 U10824 ( .A1(n13157), .A2(n12546), .ZN(n12921) );
  NAND2_X1 U10825 ( .A1(n13216), .A2(n16559), .ZN(n12917) );
  XNOR2_X1 U10826 ( .A(n13217), .B(n12919), .ZN(n12905) );
  INV_X1 U10827 ( .A(n13024), .ZN(n9070) );
  NAND2_X1 U10828 ( .A1(n13219), .A2(n16498), .ZN(n12900) );
  AND2_X1 U10829 ( .A1(n9070), .A2(n12900), .ZN(n9071) );
  OR2_X1 U10830 ( .A1(n9074), .A2(n9073), .ZN(n12396) );
  NAND2_X1 U10831 ( .A1(n13659), .A2(n13215), .ZN(n12471) );
  NAND2_X1 U10832 ( .A1(n12472), .A2(n12471), .ZN(n9076) );
  OR2_X1 U10833 ( .A1(n13659), .A2(n13215), .ZN(n12925) );
  INV_X1 U10834 ( .A(n13212), .ZN(n13584) );
  NAND2_X1 U10835 ( .A1(n13558), .A2(n13557), .ZN(n9078) );
  OR2_X1 U10836 ( .A1(n13644), .A2(n13211), .ZN(n12942) );
  NAND2_X1 U10837 ( .A1(n9078), .A2(n12942), .ZN(n13533) );
  AND2_X1 U10838 ( .A1(n13085), .A2(n13540), .ZN(n12941) );
  NAND2_X1 U10839 ( .A1(n13702), .A2(n13514), .ZN(n12853) );
  NAND2_X1 U10840 ( .A1(n13495), .A2(n13494), .ZN(n13493) );
  NAND2_X1 U10841 ( .A1(n13486), .A2(n13100), .ZN(n12851) );
  NAND2_X1 U10842 ( .A1(n13462), .A2(n12851), .ZN(n13482) );
  INV_X1 U10843 ( .A(n12960), .ZN(n9080) );
  OR2_X1 U10844 ( .A1(n13482), .A2(n9080), .ZN(n9079) );
  INV_X1 U10845 ( .A(n13478), .ZN(n13454) );
  INV_X1 U10846 ( .A(n13439), .ZN(n13466) );
  NAND2_X1 U10847 ( .A1(n13687), .A2(n13466), .ZN(n12971) );
  NAND2_X1 U10848 ( .A1(n13179), .A2(n13438), .ZN(n12847) );
  INV_X1 U10849 ( .A(n13424), .ZN(n9084) );
  NOR2_X1 U10850 ( .A1(n13425), .A2(n9084), .ZN(n9085) );
  NAND2_X1 U10851 ( .A1(n13416), .A2(n12848), .ZN(n13388) );
  NAND2_X1 U10852 ( .A1(n12978), .A2(n13076), .ZN(n12977) );
  XNOR2_X1 U10853 ( .A(n13052), .B(n13040), .ZN(n13383) );
  XNOR2_X1 U10854 ( .A(n13064), .B(n10593), .ZN(n9087) );
  OR2_X1 U10855 ( .A1(n12855), .A2(n13369), .ZN(n9086) );
  NAND2_X1 U10856 ( .A1(n9087), .A2(n9086), .ZN(n10605) );
  NAND2_X1 U10857 ( .A1(n10655), .A2(n10592), .ZN(n13046) );
  INV_X1 U10858 ( .A(n13046), .ZN(n9088) );
  AND2_X1 U10859 ( .A1(n16558), .A2(n9088), .ZN(n9089) );
  NAND2_X1 U10860 ( .A1(n10605), .A2(n9089), .ZN(n9090) );
  NAND2_X1 U10861 ( .A1(n9139), .A2(n13046), .ZN(n9126) );
  INV_X1 U10862 ( .A(n13064), .ZN(n9125) );
  OR2_X1 U10863 ( .A1(n9126), .A2(n9125), .ZN(n9124) );
  INV_X1 U10864 ( .A(n13060), .ZN(n16386) );
  INV_X1 U10865 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9093) );
  XNOR2_X1 U10866 ( .A(n9105), .B(P3_B_REG_SCAN_IN), .ZN(n9098) );
  INV_X1 U10867 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9096) );
  NAND2_X1 U10868 ( .A1(n9098), .A2(n11922), .ZN(n9104) );
  INV_X1 U10869 ( .A(n9099), .ZN(n9100) );
  NAND2_X1 U10870 ( .A1(n9100), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9101) );
  INV_X1 U10871 ( .A(n12042), .ZN(n9103) );
  NAND2_X1 U10872 ( .A1(n9105), .A2(n12042), .ZN(n10378) );
  NAND2_X1 U10873 ( .A1(n11922), .A2(n12042), .ZN(n9107) );
  XNOR2_X1 U10874 ( .A(n9141), .B(n13738), .ZN(n9123) );
  NOR2_X1 U10875 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .ZN(
        n9112) );
  NOR4_X1 U10876 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n9111) );
  NOR4_X1 U10877 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9110) );
  NOR4_X1 U10878 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9109) );
  NAND4_X1 U10879 ( .A1(n9112), .A2(n9111), .A3(n9110), .A4(n9109), .ZN(n9118)
         );
  NOR4_X1 U10880 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n9116) );
  NOR4_X1 U10881 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n9115) );
  NOR4_X1 U10882 ( .A1(P3_D_REG_7__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_2__SCAN_IN), .ZN(n9114) );
  NOR4_X1 U10883 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_8__SCAN_IN), .ZN(n9113) );
  NAND4_X1 U10884 ( .A1(n9116), .A2(n9115), .A3(n9114), .A4(n9113), .ZN(n9117)
         );
  NOR2_X1 U10885 ( .A1(n9118), .A2(n9117), .ZN(n9119) );
  OR2_X1 U10886 ( .A1(n9106), .A2(n9119), .ZN(n9140) );
  NAND2_X1 U10887 ( .A1(n7604), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9121) );
  INV_X1 U10888 ( .A(n10924), .ZN(n10603) );
  AND2_X1 U10889 ( .A1(n9140), .A2(n10603), .ZN(n9122) );
  INV_X1 U10890 ( .A(n13738), .ZN(n9130) );
  NAND2_X1 U10891 ( .A1(n9124), .A2(n12975), .ZN(n10686) );
  NAND2_X1 U10892 ( .A1(n12961), .A2(n13046), .ZN(n10684) );
  AND2_X1 U10893 ( .A1(n10686), .A2(n10684), .ZN(n9129) );
  INV_X1 U10894 ( .A(n12855), .ZN(n11070) );
  AOI22_X1 U10895 ( .A1(n9126), .A2(n11070), .B1(n10593), .B2(n9125), .ZN(
        n9127) );
  NAND2_X1 U10896 ( .A1(n9130), .A2(n9127), .ZN(n9128) );
  OAI21_X1 U10897 ( .B1(n9130), .B2(n9129), .A(n9128), .ZN(n9131) );
  INV_X1 U10898 ( .A(n9131), .ZN(n9132) );
  INV_X1 U10899 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9133) );
  NOR2_X1 U10900 ( .A1(n16565), .A2(n9133), .ZN(n9134) );
  OAI21_X1 U10901 ( .B1(n7570), .B2(n16563), .A(n9136), .ZN(P3_U3488) );
  INV_X1 U10902 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9146) );
  INV_X1 U10903 ( .A(n9141), .ZN(n9137) );
  NAND3_X1 U10904 ( .A1(n9137), .A2(n13738), .A3(n9140), .ZN(n10620) );
  OR2_X1 U10905 ( .A1(n12975), .A2(n13046), .ZN(n10692) );
  NAND2_X1 U10906 ( .A1(n11070), .A2(n9138), .ZN(n13044) );
  OR2_X1 U10907 ( .A1(n9139), .A2(n13044), .ZN(n10606) );
  AND2_X1 U10908 ( .A1(n10692), .A2(n10606), .ZN(n9144) );
  NAND2_X1 U10909 ( .A1(n9141), .A2(n9140), .ZN(n9142) );
  OR2_X1 U10910 ( .A1(n9142), .A2(n13738), .ZN(n10616) );
  INV_X1 U10911 ( .A(n10605), .ZN(n9143) );
  OAI22_X1 U10912 ( .A1(n10620), .A2(n9144), .B1(n10616), .B2(n9143), .ZN(
        n9145) );
  NOR2_X2 U10913 ( .A1(n9352), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9360) );
  NOR2_X1 U10914 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n9149) );
  NAND3_X1 U10915 ( .A1(n15867), .A2(n15885), .A3(n15868), .ZN(n9151) );
  NOR2_X1 U10916 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n9153) );
  INV_X1 U10917 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9161) );
  NAND2_X1 U10918 ( .A1(n9803), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9171) );
  INV_X1 U10919 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9163) );
  OR2_X1 U10920 ( .A1(n9808), .A2(n9163), .ZN(n9170) );
  NAND2_X1 U10921 ( .A1(n9378), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9401) );
  NAND2_X1 U10922 ( .A1(n9417), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9437) );
  INV_X1 U10923 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9586) );
  INV_X1 U10924 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9605) );
  NAND2_X1 U10925 ( .A1(n9626), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9649) );
  INV_X1 U10926 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14910) );
  INV_X1 U10927 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14862) );
  INV_X1 U10928 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14919) );
  NAND2_X1 U10929 ( .A1(n9702), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9703) );
  INV_X1 U10930 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n14824) );
  XNOR2_X1 U10931 ( .A(n9845), .B(n14824), .ZN(n15116) );
  OR2_X1 U10932 ( .A1(n9724), .A2(n15116), .ZN(n9169) );
  INV_X1 U10933 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9167) );
  OR2_X1 U10934 ( .A1(n9758), .A2(n9167), .ZN(n9168) );
  MUX2_X1 U10935 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(P1_DATAO_REG_0__SCAN_IN), 
        .S(n10029), .Z(n9172) );
  NAND2_X1 U10936 ( .A1(n9172), .A2(SI_0_), .ZN(n9281) );
  INV_X1 U10937 ( .A(n9281), .ZN(n9176) );
  INV_X1 U10938 ( .A(n9173), .ZN(n9174) );
  INV_X1 U10939 ( .A(SI_1_), .ZN(n15545) );
  NOR2_X1 U10940 ( .A1(n9174), .A2(n15545), .ZN(n9175) );
  INV_X1 U10941 ( .A(SI_2_), .ZN(n15544) );
  XNOR2_X1 U10942 ( .A(n9178), .B(n15544), .ZN(n9309) );
  NAND2_X1 U10943 ( .A1(n9178), .A2(SI_2_), .ZN(n9179) );
  XNOR2_X1 U10944 ( .A(n9181), .B(SI_3_), .ZN(n9320) );
  INV_X1 U10945 ( .A(n9320), .ZN(n9180) );
  NAND2_X1 U10946 ( .A1(n9181), .A2(SI_3_), .ZN(n9182) );
  NAND2_X1 U10947 ( .A1(n9183), .A2(n9182), .ZN(n9349) );
  XNOR2_X1 U10948 ( .A(n9185), .B(SI_4_), .ZN(n9348) );
  INV_X1 U10949 ( .A(n9348), .ZN(n9184) );
  NAND2_X1 U10950 ( .A1(n9349), .A2(n9184), .ZN(n9187) );
  NAND2_X1 U10951 ( .A1(n9185), .A2(SI_4_), .ZN(n9186) );
  NAND2_X1 U10952 ( .A1(n9187), .A2(n9186), .ZN(n9359) );
  XNOR2_X1 U10953 ( .A(n9189), .B(SI_5_), .ZN(n9358) );
  INV_X1 U10954 ( .A(n9358), .ZN(n9188) );
  NAND2_X1 U10955 ( .A1(n9189), .A2(SI_5_), .ZN(n9190) );
  MUX2_X1 U10956 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n10171), .Z(n9192) );
  XNOR2_X1 U10957 ( .A(n9192), .B(SI_6_), .ZN(n9384) );
  INV_X1 U10958 ( .A(n9384), .ZN(n9191) );
  NAND2_X1 U10959 ( .A1(n9192), .A2(SI_6_), .ZN(n9193) );
  MUX2_X1 U10960 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n10171), .Z(n9195) );
  XNOR2_X1 U10961 ( .A(n9195), .B(SI_7_), .ZN(n9408) );
  INV_X1 U10962 ( .A(n9408), .ZN(n9194) );
  NAND2_X1 U10963 ( .A1(n9409), .A2(n9194), .ZN(n9197) );
  NAND2_X1 U10964 ( .A1(n9195), .A2(SI_7_), .ZN(n9196) );
  MUX2_X1 U10965 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n10171), .Z(n9199) );
  XNOR2_X1 U10966 ( .A(n9199), .B(SI_8_), .ZN(n9424) );
  INV_X1 U10967 ( .A(n9424), .ZN(n9198) );
  NAND2_X1 U10968 ( .A1(n9199), .A2(SI_8_), .ZN(n9200) );
  MUX2_X1 U10969 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n10171), .Z(n9202) );
  XNOR2_X1 U10970 ( .A(n9202), .B(SI_9_), .ZN(n9444) );
  INV_X1 U10971 ( .A(n9444), .ZN(n9201) );
  MUX2_X1 U10972 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n10171), .Z(n9204) );
  XNOR2_X1 U10973 ( .A(n9204), .B(SI_10_), .ZN(n9461) );
  INV_X1 U10974 ( .A(n9461), .ZN(n9203) );
  NAND2_X1 U10975 ( .A1(n9462), .A2(n9203), .ZN(n9206) );
  NAND2_X1 U10976 ( .A1(n9204), .A2(SI_10_), .ZN(n9205) );
  MUX2_X1 U10977 ( .A(n10250), .B(n10255), .S(n10171), .Z(n9207) );
  INV_X1 U10978 ( .A(n9207), .ZN(n9208) );
  NAND2_X1 U10979 ( .A1(n9208), .A2(SI_11_), .ZN(n9209) );
  NAND2_X1 U10980 ( .A1(n9210), .A2(n9209), .ZN(n9486) );
  MUX2_X1 U10981 ( .A(n10287), .B(n10291), .S(n10171), .Z(n9211) );
  NAND2_X1 U10982 ( .A1(n9211), .A2(n15728), .ZN(n9214) );
  INV_X1 U10983 ( .A(n9211), .ZN(n9212) );
  NAND2_X1 U10984 ( .A1(n9212), .A2(SI_12_), .ZN(n9213) );
  MUX2_X1 U10985 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n10171), .Z(n9215) );
  NAND2_X1 U10986 ( .A1(n9215), .A2(SI_13_), .ZN(n9216) );
  MUX2_X1 U10987 ( .A(n10403), .B(n10402), .S(n10171), .Z(n9217) );
  INV_X1 U10988 ( .A(n9217), .ZN(n9218) );
  NAND2_X1 U10989 ( .A1(n9218), .A2(SI_14_), .ZN(n9219) );
  NAND2_X1 U10990 ( .A1(n9220), .A2(n9219), .ZN(n9539) );
  MUX2_X1 U10991 ( .A(n10467), .B(n12091), .S(n10171), .Z(n9221) );
  INV_X1 U10992 ( .A(n9221), .ZN(n9222) );
  NAND2_X1 U10993 ( .A1(n9222), .A2(SI_15_), .ZN(n9223) );
  MUX2_X1 U10994 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(P1_DATAO_REG_16__SCAN_IN), 
        .S(n10171), .Z(n9226) );
  INV_X1 U10995 ( .A(n9572), .ZN(n9225) );
  NAND2_X1 U10996 ( .A1(n9226), .A2(SI_16_), .ZN(n9227) );
  MUX2_X1 U10997 ( .A(n10700), .B(n10698), .S(n10171), .Z(n9229) );
  INV_X1 U10998 ( .A(n9229), .ZN(n9230) );
  NAND2_X1 U10999 ( .A1(n9230), .A2(SI_17_), .ZN(n9231) );
  NAND2_X1 U11000 ( .A1(n9232), .A2(n9231), .ZN(n9594) );
  MUX2_X1 U11001 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n10171), .Z(n9635) );
  INV_X1 U11002 ( .A(n9635), .ZN(n9233) );
  MUX2_X1 U11003 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n10171), .Z(n9235) );
  NAND2_X1 U11004 ( .A1(n9235), .A2(SI_19_), .ZN(n9642) );
  OAI21_X1 U11005 ( .B1(n15716), .B2(n9233), .A(n9642), .ZN(n9234) );
  NOR2_X1 U11006 ( .A1(n9635), .A2(SI_18_), .ZN(n9238) );
  INV_X1 U11007 ( .A(n9235), .ZN(n9236) );
  INV_X1 U11008 ( .A(SI_19_), .ZN(n15512) );
  NAND2_X1 U11009 ( .A1(n9236), .A2(n15512), .ZN(n9641) );
  INV_X1 U11010 ( .A(n9641), .ZN(n9237) );
  AOI21_X1 U11011 ( .B1(n9238), .B2(n9642), .A(n9237), .ZN(n9239) );
  MUX2_X1 U11012 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n10171), .Z(n9657) );
  INV_X1 U11013 ( .A(n9657), .ZN(n9243) );
  INV_X1 U11014 ( .A(n9240), .ZN(n9241) );
  MUX2_X1 U11015 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n10171), .Z(n9245) );
  XNOR2_X1 U11016 ( .A(n9245), .B(SI_21_), .ZN(n9677) );
  NAND2_X1 U11017 ( .A1(n9245), .A2(SI_21_), .ZN(n9246) );
  INV_X1 U11018 ( .A(n11957), .ZN(n9248) );
  MUX2_X1 U11019 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n10197), .Z(n11956) );
  NAND2_X1 U11020 ( .A1(n9249), .A2(SI_22_), .ZN(n9250) );
  MUX2_X1 U11021 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n10171), .Z(n9251) );
  XNOR2_X1 U11022 ( .A(n9251), .B(SI_23_), .ZN(n9712) );
  NAND2_X1 U11023 ( .A1(n9251), .A2(SI_23_), .ZN(n9252) );
  MUX2_X1 U11024 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n10197), .Z(n9730) );
  NAND2_X1 U11025 ( .A1(n9254), .A2(SI_24_), .ZN(n9255) );
  MUX2_X1 U11026 ( .A(n15917), .B(n14817), .S(n10171), .Z(n9257) );
  NAND2_X1 U11027 ( .A1(n9257), .A2(n15704), .ZN(n9260) );
  INV_X1 U11028 ( .A(n9257), .ZN(n9258) );
  NAND2_X1 U11029 ( .A1(n9258), .A2(SI_25_), .ZN(n9259) );
  NAND2_X1 U11030 ( .A1(n9260), .A2(n9259), .ZN(n9749) );
  MUX2_X1 U11031 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n10197), .Z(n9261) );
  XNOR2_X1 U11032 ( .A(n9261), .B(n15502), .ZN(n9763) );
  NAND2_X1 U11033 ( .A1(n9261), .A2(SI_26_), .ZN(n9262) );
  MUX2_X1 U11034 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n10171), .Z(n9783) );
  XNOR2_X1 U11035 ( .A(n9783), .B(n15700), .ZN(n9781) );
  INV_X1 U11036 ( .A(n9781), .ZN(n9263) );
  NAND2_X2 U11037 ( .A1(n9943), .A2(n15912), .ZN(n10266) );
  NAND2_X1 U11038 ( .A1(n10266), .A2(n10196), .ZN(n9796) );
  NAND2_X1 U11039 ( .A1(n14806), .A2(n9679), .ZN(n9267) );
  NAND2_X1 U11040 ( .A1(n7719), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9266) );
  NAND2_X1 U11041 ( .A1(n9274), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9268) );
  MUX2_X1 U11042 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9268), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n9269) );
  NAND2_X1 U11043 ( .A1(n9934), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9270) );
  MUX2_X1 U11044 ( .A(n9270), .B(P1_IR_REG_31__SCAN_IN), .S(n8135), .Z(n9271)
         );
  INV_X1 U11045 ( .A(n9271), .ZN(n9272) );
  NOR2_X2 U11046 ( .A1(n9272), .A2(n9927), .ZN(n9841) );
  MUX2_X1 U11047 ( .A(n14939), .B(n15376), .S(n9857), .Z(n9776) );
  INV_X1 U11048 ( .A(n9776), .ZN(n9780) );
  INV_X1 U11049 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10315) );
  INV_X1 U11050 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10503) );
  INV_X1 U11051 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9276) );
  OR2_X1 U11052 ( .A1(n9303), .A2(n9276), .ZN(n9278) );
  NAND2_X1 U11053 ( .A1(n9842), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9277) );
  NAND4_X2 U11054 ( .A1(n9280), .A2(n9279), .A3(n9278), .A4(n9277), .ZN(n10517) );
  NAND2_X1 U11055 ( .A1(n9372), .A2(n10517), .ZN(n9289) );
  INV_X1 U11056 ( .A(n10517), .ZN(n10651) );
  NAND2_X1 U11057 ( .A1(n9338), .A2(n10651), .ZN(n9288) );
  XNOR2_X1 U11058 ( .A(n9282), .B(n9281), .ZN(n10228) );
  NAND2_X1 U11059 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9284) );
  XNOR2_X1 U11060 ( .A(n9284), .B(P1_IR_REG_1__SCAN_IN), .ZN(n14982) );
  INV_X1 U11061 ( .A(n14982), .ZN(n9285) );
  OAI211_X2 U11062 ( .C1(n9796), .C2(n10228), .A(n9287), .B(n9286), .ZN(n10516) );
  INV_X1 U11063 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11123) );
  INV_X1 U11064 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9293) );
  OR2_X1 U11065 ( .A1(n9304), .A2(n9293), .ZN(n9294) );
  NOR2_X1 U11066 ( .A1(n10171), .A2(n10175), .ZN(n9298) );
  XNOR2_X1 U11067 ( .A(n9298), .B(n9297), .ZN(n15922) );
  MUX2_X1 U11068 ( .A(P1_IR_REG_0__SCAN_IN), .B(n15922), .S(n10266), .Z(n11126) );
  NAND2_X1 U11069 ( .A1(n10522), .A2(n10437), .ZN(n9299) );
  INV_X1 U11070 ( .A(n10439), .ZN(n14974) );
  INV_X1 U11071 ( .A(n11126), .ZN(n11207) );
  NAND2_X1 U11072 ( .A1(n14974), .A2(n11207), .ZN(n9892) );
  NAND2_X1 U11073 ( .A1(n9299), .A2(n9892), .ZN(n9301) );
  INV_X1 U11074 ( .A(n10522), .ZN(n9300) );
  XNOR2_X1 U11075 ( .A(n10517), .B(n10516), .ZN(n9970) );
  NAND2_X1 U11076 ( .A1(n9302), .A2(n9974), .ZN(n9317) );
  INV_X1 U11077 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10303) );
  OR2_X1 U11078 ( .A1(n9304), .A2(n10303), .ZN(n9307) );
  INV_X1 U11079 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n15340) );
  INV_X1 U11080 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10458) );
  XNOR2_X1 U11081 ( .A(n9310), .B(n9309), .ZN(n10180) );
  NAND2_X1 U11082 ( .A1(n9350), .A2(n10180), .ZN(n9315) );
  OR2_X1 U11083 ( .A1(n9311), .A2(n9361), .ZN(n9312) );
  NAND2_X1 U11084 ( .A1(n9332), .A2(n15342), .ZN(n9316) );
  XNOR2_X1 U11085 ( .A(n9319), .B(n9320), .ZN(n10178) );
  NAND2_X1 U11086 ( .A1(n10178), .A2(n9350), .ZN(n9325) );
  NAND2_X1 U11087 ( .A1(n9321), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9322) );
  XNOR2_X1 U11088 ( .A(n9322), .B(P1_IR_REG_3__SCAN_IN), .ZN(n14993) );
  NAND2_X1 U11089 ( .A1(n7883), .A2(n14993), .ZN(n9324) );
  NAND2_X1 U11090 ( .A1(n9283), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9323) );
  NAND2_X1 U11091 ( .A1(n9326), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9330) );
  NAND2_X1 U11092 ( .A1(n9804), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9329) );
  OR2_X1 U11093 ( .A1(n9724), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9328) );
  INV_X1 U11094 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10307) );
  AND2_X1 U11095 ( .A1(n16429), .A2(n14973), .ZN(n9340) );
  NAND2_X1 U11096 ( .A1(n9372), .A2(n10857), .ZN(n9331) );
  OAI21_X1 U11097 ( .B1(n9372), .B2(n9340), .A(n9331), .ZN(n9337) );
  AND2_X1 U11098 ( .A1(n10642), .A2(n9332), .ZN(n9333) );
  NAND2_X1 U11099 ( .A1(n9338), .A2(n9333), .ZN(n9334) );
  OAI21_X1 U11100 ( .B1(n9338), .B2(n10855), .A(n9334), .ZN(n9335) );
  INV_X1 U11101 ( .A(n9335), .ZN(n9336) );
  NAND2_X1 U11102 ( .A1(n9338), .A2(n10857), .ZN(n9339) );
  OAI21_X1 U11103 ( .B1(n9413), .B2(n9340), .A(n9339), .ZN(n9341) );
  NAND2_X1 U11104 ( .A1(n9804), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9347) );
  INV_X1 U11105 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9343) );
  OR2_X1 U11106 ( .A1(n9304), .A2(n9343), .ZN(n9346) );
  INV_X1 U11107 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10321) );
  OR2_X1 U11108 ( .A1(n9843), .A2(n10321), .ZN(n9345) );
  XNOR2_X1 U11109 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n11160) );
  OR2_X1 U11110 ( .A1(n9724), .A2(n11160), .ZN(n9344) );
  XNOR2_X1 U11111 ( .A(n9349), .B(n9348), .ZN(n10192) );
  NAND2_X1 U11112 ( .A1(n10192), .A2(n9350), .ZN(n9355) );
  NAND2_X1 U11113 ( .A1(n9352), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9353) );
  XNOR2_X1 U11114 ( .A(n9353), .B(P1_IR_REG_4__SCAN_IN), .ZN(n16341) );
  AOI22_X1 U11115 ( .A1(n9283), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n7883), .B2(
        n16341), .ZN(n9354) );
  INV_X1 U11116 ( .A(n10915), .ZN(n14972) );
  XNOR2_X1 U11117 ( .A(n9359), .B(n9358), .ZN(n10552) );
  NAND2_X1 U11118 ( .A1(n10552), .A2(n9679), .ZN(n9364) );
  OR2_X1 U11119 ( .A1(n9360), .A2(n9361), .ZN(n9362) );
  XNOR2_X1 U11120 ( .A(n9362), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10370) );
  AOI22_X1 U11121 ( .A1(n7719), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7883), .B2(
        n10370), .ZN(n9363) );
  NAND2_X1 U11122 ( .A1(n9364), .A2(n9363), .ZN(n10909) );
  INV_X1 U11123 ( .A(n9847), .ZN(n9705) );
  AOI21_X1 U11124 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9365) );
  NOR2_X1 U11125 ( .A1(n9365), .A2(n9378), .ZN(n10918) );
  NAND2_X1 U11126 ( .A1(n9705), .A2(n10918), .ZN(n9371) );
  INV_X1 U11127 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10865) );
  OR2_X1 U11128 ( .A1(n9843), .A2(n10865), .ZN(n9370) );
  INV_X1 U11129 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9366) );
  OR2_X1 U11130 ( .A1(n9758), .A2(n9366), .ZN(n9369) );
  INV_X1 U11131 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9367) );
  OR2_X1 U11132 ( .A1(n9808), .A2(n9367), .ZN(n9368) );
  MUX2_X1 U11133 ( .A(n10909), .B(n14971), .S(n9372), .Z(n9374) );
  MUX2_X1 U11134 ( .A(n14971), .B(n10909), .S(n9372), .Z(n9373) );
  NAND2_X1 U11135 ( .A1(n7717), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9383) );
  INV_X1 U11136 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11072) );
  OR2_X1 U11137 ( .A1(n9843), .A2(n11072), .ZN(n9382) );
  OAI21_X1 U11138 ( .B1(n9378), .B2(P1_REG3_REG_6__SCAN_IN), .A(n9401), .ZN(
        n11152) );
  OR2_X1 U11139 ( .A1(n9847), .A2(n11152), .ZN(n9381) );
  INV_X1 U11140 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9379) );
  OR2_X1 U11141 ( .A1(n9758), .A2(n9379), .ZN(n9380) );
  NAND4_X1 U11142 ( .A1(n9383), .A2(n9382), .A3(n9381), .A4(n9380), .ZN(n14970) );
  XNOR2_X1 U11143 ( .A(n9385), .B(n9384), .ZN(n10560) );
  NAND2_X1 U11144 ( .A1(n10560), .A2(n9679), .ZN(n9390) );
  NAND2_X1 U11145 ( .A1(n9360), .A2(n15867), .ZN(n9387) );
  NAND2_X1 U11146 ( .A1(n9387), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9386) );
  MUX2_X1 U11147 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9386), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n9388) );
  AND2_X1 U11148 ( .A1(n9388), .A2(n9560), .ZN(n10351) );
  AOI22_X1 U11149 ( .A1(n7719), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7883), .B2(
        n10351), .ZN(n9389) );
  NAND2_X1 U11150 ( .A1(n9390), .A2(n9389), .ZN(n11537) );
  MUX2_X1 U11151 ( .A(n14970), .B(n11537), .S(n7710), .Z(n9394) );
  NAND2_X1 U11152 ( .A1(n9393), .A2(n9394), .ZN(n9392) );
  MUX2_X1 U11153 ( .A(n14970), .B(n11537), .S(n9413), .Z(n9391) );
  NAND2_X1 U11154 ( .A1(n9392), .A2(n9391), .ZN(n9398) );
  INV_X1 U11155 ( .A(n9393), .ZN(n9396) );
  INV_X1 U11156 ( .A(n9394), .ZN(n9395) );
  NAND2_X1 U11157 ( .A1(n9396), .A2(n9395), .ZN(n9397) );
  NAND2_X1 U11158 ( .A1(n9803), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9407) );
  INV_X1 U11159 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9399) );
  OR2_X1 U11160 ( .A1(n9808), .A2(n9399), .ZN(n9406) );
  AND2_X1 U11161 ( .A1(n9401), .A2(n9400), .ZN(n9402) );
  OR2_X1 U11162 ( .A1(n9402), .A2(n9417), .ZN(n11533) );
  OR2_X1 U11163 ( .A1(n9847), .A2(n11533), .ZN(n9405) );
  INV_X1 U11164 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9403) );
  OR2_X1 U11165 ( .A1(n9758), .A2(n9403), .ZN(n9404) );
  NAND4_X1 U11166 ( .A1(n9407), .A2(n9406), .A3(n9405), .A4(n9404), .ZN(n14969) );
  NAND2_X1 U11167 ( .A1(n10723), .A2(n9679), .ZN(n9412) );
  NAND2_X1 U11168 ( .A1(n9560), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9410) );
  XNOR2_X1 U11169 ( .A(n9410), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10384) );
  AOI22_X1 U11170 ( .A1(n7719), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7883), .B2(
        n10384), .ZN(n9411) );
  NAND2_X1 U11171 ( .A1(n9412), .A2(n9411), .ZN(n16478) );
  MUX2_X1 U11172 ( .A(n14969), .B(n16478), .S(n9413), .Z(n9415) );
  MUX2_X1 U11173 ( .A(n14969), .B(n16478), .S(n7710), .Z(n9414) );
  INV_X1 U11174 ( .A(n9415), .ZN(n9416) );
  NAND2_X1 U11175 ( .A1(n7717), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9423) );
  INV_X1 U11176 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10385) );
  OR2_X1 U11177 ( .A1(n9843), .A2(n10385), .ZN(n9422) );
  OR2_X1 U11178 ( .A1(n9417), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9418) );
  NAND2_X1 U11179 ( .A1(n9437), .A2(n9418), .ZN(n11739) );
  OR2_X1 U11180 ( .A1(n9847), .A2(n11739), .ZN(n9421) );
  INV_X1 U11181 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9419) );
  OR2_X1 U11182 ( .A1(n9758), .A2(n9419), .ZN(n9420) );
  NAND4_X1 U11183 ( .A1(n9423), .A2(n9422), .A3(n9421), .A4(n9420), .ZN(n14968) );
  XNOR2_X1 U11184 ( .A(n9425), .B(n9424), .ZN(n10730) );
  NAND2_X1 U11185 ( .A1(n10730), .A2(n9679), .ZN(n9428) );
  NAND2_X1 U11186 ( .A1(n9446), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9426) );
  XNOR2_X1 U11187 ( .A(n9426), .B(P1_IR_REG_8__SCAN_IN), .ZN(n15007) );
  AOI22_X1 U11188 ( .A1(n7719), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7883), .B2(
        n15007), .ZN(n9427) );
  NAND2_X1 U11189 ( .A1(n9428), .A2(n9427), .ZN(n11756) );
  MUX2_X1 U11190 ( .A(n14968), .B(n11756), .S(n9837), .Z(n9431) );
  NAND2_X1 U11191 ( .A1(n9432), .A2(n9431), .ZN(n9430) );
  MUX2_X1 U11192 ( .A(n14968), .B(n11756), .S(n9857), .Z(n9429) );
  NAND2_X1 U11193 ( .A1(n9430), .A2(n9429), .ZN(n9434) );
  NAND2_X1 U11194 ( .A1(n9803), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9443) );
  INV_X1 U11195 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9435) );
  OR2_X1 U11196 ( .A1(n9808), .A2(n9435), .ZN(n9442) );
  NAND2_X1 U11197 ( .A1(n9437), .A2(n9436), .ZN(n9438) );
  NAND2_X1 U11198 ( .A1(n9454), .A2(n9438), .ZN(n11819) );
  OR2_X1 U11199 ( .A1(n9847), .A2(n11819), .ZN(n9441) );
  INV_X1 U11200 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9439) );
  OR2_X1 U11201 ( .A1(n9758), .A2(n9439), .ZN(n9440) );
  NAND4_X1 U11202 ( .A1(n9443), .A2(n9442), .A3(n9441), .A4(n9440), .ZN(n14967) );
  XNOR2_X1 U11203 ( .A(n9445), .B(n9444), .ZN(n10978) );
  NAND2_X1 U11204 ( .A1(n10978), .A2(n9679), .ZN(n9450) );
  INV_X1 U11205 ( .A(n9446), .ZN(n9447) );
  INV_X1 U11206 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n15874) );
  NAND2_X1 U11207 ( .A1(n9447), .A2(n15874), .ZN(n9463) );
  NAND2_X1 U11208 ( .A1(n9463), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9448) );
  XNOR2_X1 U11209 ( .A(n9448), .B(P1_IR_REG_9__SCAN_IN), .ZN(n15024) );
  AOI22_X1 U11210 ( .A1(n7719), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7883), .B2(
        n15024), .ZN(n9449) );
  MUX2_X1 U11211 ( .A(n14967), .B(n11818), .S(n9857), .Z(n9452) );
  MUX2_X1 U11212 ( .A(n14967), .B(n11818), .S(n9837), .Z(n9451) );
  NAND2_X1 U11213 ( .A1(n7717), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9460) );
  INV_X1 U11214 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11767) );
  OR2_X1 U11215 ( .A1(n9843), .A2(n11767), .ZN(n9459) );
  NAND2_X1 U11216 ( .A1(n9454), .A2(n9453), .ZN(n9455) );
  NAND2_X1 U11217 ( .A1(n9480), .A2(n9455), .ZN(n11972) );
  OR2_X1 U11218 ( .A1(n9847), .A2(n11972), .ZN(n9458) );
  INV_X1 U11219 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9456) );
  OR2_X1 U11220 ( .A1(n9758), .A2(n9456), .ZN(n9457) );
  NAND4_X1 U11221 ( .A1(n9460), .A2(n9459), .A3(n9458), .A4(n9457), .ZN(n14966) );
  XNOR2_X1 U11222 ( .A(n9462), .B(n9461), .ZN(n11341) );
  NAND2_X1 U11223 ( .A1(n11341), .A2(n9679), .ZN(n9470) );
  INV_X1 U11224 ( .A(n9463), .ZN(n9465) );
  INV_X1 U11225 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9464) );
  NAND2_X1 U11226 ( .A1(n9465), .A2(n9464), .ZN(n9467) );
  NAND2_X1 U11227 ( .A1(n9467), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9466) );
  MUX2_X1 U11228 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9466), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n9468) );
  AOI22_X1 U11229 ( .A1(n10425), .A2(n7883), .B1(n7719), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n9469) );
  MUX2_X1 U11230 ( .A(n14966), .B(n11963), .S(n9837), .Z(n9474) );
  NAND2_X1 U11231 ( .A1(n9473), .A2(n9474), .ZN(n9472) );
  MUX2_X1 U11232 ( .A(n14966), .B(n11963), .S(n9857), .Z(n9471) );
  NAND2_X1 U11233 ( .A1(n9472), .A2(n9471), .ZN(n9478) );
  INV_X1 U11234 ( .A(n9473), .ZN(n9476) );
  INV_X1 U11235 ( .A(n9474), .ZN(n9475) );
  NAND2_X1 U11236 ( .A1(n9476), .A2(n9475), .ZN(n9477) );
  NAND2_X1 U11237 ( .A1(n7717), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9485) );
  INV_X1 U11238 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11867) );
  OR2_X1 U11239 ( .A1(n9843), .A2(n11867), .ZN(n9484) );
  OR2_X1 U11240 ( .A1(n8518), .A2(n9494), .ZN(n12065) );
  OR2_X1 U11241 ( .A1(n9724), .A2(n12065), .ZN(n9483) );
  INV_X1 U11242 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9481) );
  OR2_X1 U11243 ( .A1(n9758), .A2(n9481), .ZN(n9482) );
  NAND4_X1 U11244 ( .A1(n9485), .A2(n9484), .A3(n9483), .A4(n9482), .ZN(n14965) );
  XNOR2_X1 U11245 ( .A(n9487), .B(n9486), .ZN(n11603) );
  NAND2_X1 U11246 ( .A1(n11603), .A2(n9679), .ZN(n9490) );
  NAND2_X1 U11247 ( .A1(n9501), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9488) );
  XNOR2_X1 U11248 ( .A(n9488), .B(P1_IR_REG_11__SCAN_IN), .ZN(n15039) );
  AOI22_X1 U11249 ( .A1(n15039), .A2(n7883), .B1(n7719), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n9489) );
  MUX2_X1 U11250 ( .A(n14965), .B(n12153), .S(n9857), .Z(n9492) );
  MUX2_X1 U11251 ( .A(n14965), .B(n12153), .S(n9837), .Z(n9491) );
  INV_X1 U11252 ( .A(n9492), .ZN(n9493) );
  NAND2_X1 U11253 ( .A1(n9804), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9499) );
  INV_X1 U11254 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10429) );
  OR2_X1 U11255 ( .A1(n9843), .A2(n10429), .ZN(n9498) );
  OR2_X1 U11256 ( .A1(n9494), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9495) );
  NAND2_X1 U11257 ( .A1(n9514), .A2(n9495), .ZN(n12178) );
  OR2_X1 U11258 ( .A1(n9847), .A2(n12178), .ZN(n9497) );
  INV_X1 U11259 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10672) );
  OR2_X1 U11260 ( .A1(n9808), .A2(n10672), .ZN(n9496) );
  NAND4_X1 U11261 ( .A1(n9499), .A2(n9498), .A3(n9497), .A4(n9496), .ZN(n14963) );
  XNOR2_X1 U11262 ( .A(n9500), .B(n8517), .ZN(n11774) );
  NAND2_X1 U11263 ( .A1(n11774), .A2(n9679), .ZN(n9503) );
  OAI21_X1 U11264 ( .B1(n9501), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9524) );
  XNOR2_X1 U11265 ( .A(n9524), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10666) );
  AOI22_X1 U11266 ( .A1(n10666), .A2(n7883), .B1(n7719), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n9502) );
  MUX2_X1 U11267 ( .A(n14963), .B(n15470), .S(n9837), .Z(n9507) );
  NAND2_X1 U11268 ( .A1(n9506), .A2(n9507), .ZN(n9505) );
  MUX2_X1 U11269 ( .A(n14963), .B(n15470), .S(n9857), .Z(n9504) );
  NAND2_X1 U11270 ( .A1(n9505), .A2(n9504), .ZN(n9511) );
  INV_X1 U11271 ( .A(n9506), .ZN(n9509) );
  INV_X1 U11272 ( .A(n9507), .ZN(n9508) );
  NAND2_X1 U11273 ( .A1(n9509), .A2(n9508), .ZN(n9510) );
  NAND2_X1 U11274 ( .A1(n9803), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9520) );
  INV_X1 U11275 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9512) );
  OR2_X1 U11276 ( .A1(n9758), .A2(n9512), .ZN(n9519) );
  NAND2_X1 U11277 ( .A1(n9514), .A2(n9513), .ZN(n9515) );
  NAND2_X1 U11278 ( .A1(n9533), .A2(n9515), .ZN(n12307) );
  OR2_X1 U11279 ( .A1(n9847), .A2(n12307), .ZN(n9518) );
  INV_X1 U11280 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9516) );
  OR2_X1 U11281 ( .A1(n9808), .A2(n9516), .ZN(n9517) );
  NAND4_X1 U11282 ( .A1(n9520), .A2(n9519), .A3(n9518), .A4(n9517), .ZN(n14962) );
  NAND2_X1 U11283 ( .A1(n11901), .A2(n9679), .ZN(n9529) );
  INV_X1 U11284 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9523) );
  NAND2_X1 U11285 ( .A1(n9524), .A2(n9523), .ZN(n9525) );
  NAND2_X1 U11286 ( .A1(n9525), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9526) );
  INV_X1 U11287 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n15675) );
  NAND2_X1 U11288 ( .A1(n9526), .A2(n15675), .ZN(n9541) );
  OR2_X1 U11289 ( .A1(n9526), .A2(n15675), .ZN(n9527) );
  AOI22_X1 U11290 ( .A1(n10675), .A2(n7883), .B1(n7719), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n9528) );
  MUX2_X1 U11291 ( .A(n14962), .B(n12333), .S(n9857), .Z(n9531) );
  MUX2_X1 U11292 ( .A(n14962), .B(n12333), .S(n9837), .Z(n9530) );
  AND2_X1 U11293 ( .A1(n9533), .A2(n9532), .ZN(n9534) );
  OR2_X1 U11294 ( .A1(n9534), .A2(n9553), .ZN(n12387) );
  INV_X1 U11295 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10674) );
  OR2_X1 U11296 ( .A1(n9808), .A2(n10674), .ZN(n9536) );
  INV_X1 U11297 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n12341) );
  OR2_X1 U11298 ( .A1(n9843), .A2(n12341), .ZN(n9535) );
  AND2_X1 U11299 ( .A1(n9536), .A2(n9535), .ZN(n9538) );
  NAND2_X1 U11300 ( .A1(n9804), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9537) );
  OAI211_X1 U11301 ( .C1(n9847), .C2(n12387), .A(n9538), .B(n9537), .ZN(n15332) );
  XNOR2_X1 U11302 ( .A(n9540), .B(n9539), .ZN(n12014) );
  NAND2_X1 U11303 ( .A1(n12014), .A2(n9679), .ZN(n9544) );
  NAND2_X1 U11304 ( .A1(n9541), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9542) );
  AOI22_X1 U11305 ( .A1(n11378), .A2(n7883), .B1(n7719), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9543) );
  MUX2_X1 U11306 ( .A(n15332), .B(n15456), .S(n9837), .Z(n9548) );
  NAND2_X1 U11307 ( .A1(n9547), .A2(n9548), .ZN(n9546) );
  MUX2_X1 U11308 ( .A(n15332), .B(n15456), .S(n9857), .Z(n9545) );
  NAND2_X1 U11309 ( .A1(n9546), .A2(n9545), .ZN(n9552) );
  INV_X1 U11310 ( .A(n9547), .ZN(n9550) );
  INV_X1 U11311 ( .A(n9548), .ZN(n9549) );
  NAND2_X1 U11312 ( .A1(n9550), .A2(n9549), .ZN(n9551) );
  NOR2_X1 U11313 ( .A1(n9553), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9554) );
  OR2_X1 U11314 ( .A1(n9568), .A2(n9554), .ZN(n15322) );
  AOI22_X1 U11315 ( .A1(n7717), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n9803), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n9556) );
  NAND2_X1 U11316 ( .A1(n9804), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n9555) );
  OAI211_X1 U11317 ( .C1(n15322), .C2(n9847), .A(n9556), .B(n9555), .ZN(n15303) );
  XNOR2_X1 U11318 ( .A(n9558), .B(n9557), .ZN(n12090) );
  NAND2_X1 U11319 ( .A1(n12090), .A2(n9679), .ZN(n9564) );
  OAI21_X1 U11320 ( .B1(n9560), .B2(n9559), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9561) );
  MUX2_X1 U11321 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9561), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n9562) );
  AND2_X1 U11322 ( .A1(n9574), .A2(n9562), .ZN(n11570) );
  AOI22_X1 U11323 ( .A1(n7719), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7883), 
        .B2(n11570), .ZN(n9563) );
  MUX2_X1 U11324 ( .A(n15303), .B(n15451), .S(n9857), .Z(n9566) );
  MUX2_X1 U11325 ( .A(n15303), .B(n15451), .S(n9837), .Z(n9565) );
  INV_X1 U11326 ( .A(n9566), .ZN(n9567) );
  OR2_X1 U11327 ( .A1(n9568), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9569) );
  NAND2_X1 U11328 ( .A1(n9587), .A2(n9569), .ZN(n15313) );
  AOI22_X1 U11329 ( .A1(n7717), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9803), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n9571) );
  NAND2_X1 U11330 ( .A1(n9804), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9570) );
  OAI211_X1 U11331 ( .C1(n15313), .C2(n9847), .A(n9571), .B(n9570), .ZN(n15330) );
  XNOR2_X1 U11332 ( .A(n9573), .B(n9572), .ZN(n12211) );
  NAND2_X1 U11333 ( .A1(n12211), .A2(n9679), .ZN(n9577) );
  NAND2_X1 U11334 ( .A1(n9574), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9575) );
  XNOR2_X1 U11335 ( .A(n9575), .B(P1_IR_REG_16__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U11336 ( .A1(n7719), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7883), 
        .B2(n11705), .ZN(n9576) );
  MUX2_X1 U11337 ( .A(n15330), .B(n15446), .S(n9837), .Z(n9581) );
  NAND2_X1 U11338 ( .A1(n9580), .A2(n9581), .ZN(n9579) );
  MUX2_X1 U11339 ( .A(n15330), .B(n15446), .S(n9857), .Z(n9578) );
  NAND2_X1 U11340 ( .A1(n9579), .A2(n9578), .ZN(n9585) );
  INV_X1 U11341 ( .A(n9580), .ZN(n9583) );
  INV_X1 U11342 ( .A(n9581), .ZN(n9582) );
  NAND2_X1 U11343 ( .A1(n9583), .A2(n9582), .ZN(n9584) );
  NAND2_X1 U11344 ( .A1(n9587), .A2(n9586), .ZN(n9588) );
  AND2_X1 U11345 ( .A1(n9606), .A2(n9588), .ZN(n15294) );
  NAND2_X1 U11346 ( .A1(n15294), .A2(n9705), .ZN(n9593) );
  INV_X1 U11347 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n15048) );
  NAND2_X1 U11348 ( .A1(n9804), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9590) );
  NAND2_X1 U11349 ( .A1(n9803), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9589) );
  OAI211_X1 U11350 ( .C1(n9808), .C2(n15048), .A(n9590), .B(n9589), .ZN(n9591)
         );
  INV_X1 U11351 ( .A(n9591), .ZN(n9592) );
  NAND2_X1 U11352 ( .A1(n9593), .A2(n9592), .ZN(n15304) );
  XNOR2_X1 U11353 ( .A(n9595), .B(n9594), .ZN(n12354) );
  NAND2_X1 U11354 ( .A1(n12354), .A2(n9679), .ZN(n9601) );
  NAND2_X1 U11355 ( .A1(n9596), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9597) );
  MUX2_X1 U11356 ( .A(n9597), .B(P1_IR_REG_31__SCAN_IN), .S(n7840), .Z(n9599)
         );
  AND2_X1 U11357 ( .A1(n9599), .A2(n9614), .ZN(n11708) );
  AOI22_X1 U11358 ( .A1(n7719), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7883), 
        .B2(n11708), .ZN(n9600) );
  MUX2_X1 U11359 ( .A(n15304), .B(n15440), .S(n9857), .Z(n9603) );
  MUX2_X1 U11360 ( .A(n15304), .B(n15440), .S(n9837), .Z(n9602) );
  INV_X1 U11361 ( .A(n9603), .ZN(n9604) );
  AND2_X1 U11362 ( .A1(n9606), .A2(n9605), .ZN(n9607) );
  OR2_X1 U11363 ( .A1(n9607), .A2(n9626), .ZN(n15271) );
  INV_X1 U11364 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9611) );
  NAND2_X1 U11365 ( .A1(n9804), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9610) );
  INV_X1 U11366 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9608) );
  OR2_X1 U11367 ( .A1(n9843), .A2(n9608), .ZN(n9609) );
  OAI211_X1 U11368 ( .C1(n9808), .C2(n9611), .A(n9610), .B(n9609), .ZN(n9612)
         );
  INV_X1 U11369 ( .A(n9612), .ZN(n9613) );
  OAI21_X1 U11370 ( .B1(n15271), .B2(n9847), .A(n9613), .ZN(n15289) );
  XNOR2_X1 U11371 ( .A(n9637), .B(n15716), .ZN(n9634) );
  XNOR2_X1 U11372 ( .A(n9634), .B(n9635), .ZN(n12423) );
  NAND2_X1 U11373 ( .A1(n12423), .A2(n9679), .ZN(n9617) );
  NAND2_X1 U11374 ( .A1(n9614), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9615) );
  XNOR2_X1 U11375 ( .A(n9615), .B(P1_IR_REG_18__SCAN_IN), .ZN(n15059) );
  AOI22_X1 U11376 ( .A1(n7719), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7883), 
        .B2(n15059), .ZN(n9616) );
  MUX2_X1 U11377 ( .A(n15289), .B(n15435), .S(n9837), .Z(n9621) );
  NAND2_X1 U11378 ( .A1(n9620), .A2(n9621), .ZN(n9619) );
  MUX2_X1 U11379 ( .A(n15289), .B(n15435), .S(n9857), .Z(n9618) );
  NAND2_X1 U11380 ( .A1(n9619), .A2(n9618), .ZN(n9625) );
  INV_X1 U11381 ( .A(n9620), .ZN(n9623) );
  INV_X1 U11382 ( .A(n9621), .ZN(n9622) );
  NAND2_X1 U11383 ( .A1(n9623), .A2(n9622), .ZN(n9624) );
  OR2_X1 U11384 ( .A1(n9626), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9627) );
  AND2_X1 U11385 ( .A1(n9649), .A2(n9627), .ZN(n15259) );
  NAND2_X1 U11386 ( .A1(n15259), .A2(n9705), .ZN(n9633) );
  INV_X1 U11387 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9630) );
  NAND2_X1 U11388 ( .A1(n9804), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9629) );
  NAND2_X1 U11389 ( .A1(n9803), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9628) );
  OAI211_X1 U11390 ( .C1(n9808), .C2(n9630), .A(n9629), .B(n9628), .ZN(n9631)
         );
  INV_X1 U11391 ( .A(n9631), .ZN(n9632) );
  NAND2_X1 U11392 ( .A1(n9633), .A2(n9632), .ZN(n15270) );
  INV_X1 U11393 ( .A(n9634), .ZN(n9636) );
  NAND2_X1 U11394 ( .A1(n9636), .A2(n9635), .ZN(n9640) );
  INV_X1 U11395 ( .A(n9637), .ZN(n9638) );
  NAND2_X1 U11396 ( .A1(n9638), .A2(SI_18_), .ZN(n9639) );
  NAND2_X1 U11397 ( .A1(n9640), .A2(n9639), .ZN(n9644) );
  NAND2_X1 U11398 ( .A1(n9642), .A2(n9641), .ZN(n9643) );
  NAND2_X1 U11399 ( .A1(n12590), .A2(n9679), .ZN(n9646) );
  AOI22_X1 U11400 ( .A1(n7719), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n15185), 
        .B2(n7883), .ZN(n9645) );
  MUX2_X1 U11401 ( .A(n15270), .B(n15257), .S(n9857), .Z(n9648) );
  MUX2_X1 U11402 ( .A(n15270), .B(n15257), .S(n9837), .Z(n9647) );
  NAND2_X1 U11403 ( .A1(n9649), .A2(n14910), .ZN(n9650) );
  NAND2_X1 U11404 ( .A1(n9669), .A2(n9650), .ZN(n15241) );
  OR2_X1 U11405 ( .A1(n15241), .A2(n9724), .ZN(n9656) );
  INV_X1 U11406 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9653) );
  NAND2_X1 U11407 ( .A1(n9803), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9652) );
  NAND2_X1 U11408 ( .A1(n9804), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9651) );
  OAI211_X1 U11409 ( .C1(n9808), .C2(n9653), .A(n9652), .B(n9651), .ZN(n9654)
         );
  INV_X1 U11410 ( .A(n9654), .ZN(n9655) );
  NAND2_X1 U11411 ( .A1(n9656), .A2(n9655), .ZN(n15258) );
  XNOR2_X1 U11412 ( .A(n9658), .B(n9657), .ZN(n12508) );
  NAND2_X1 U11413 ( .A1(n12508), .A2(n9679), .ZN(n9660) );
  NAND2_X1 U11414 ( .A1(n7719), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9659) );
  MUX2_X1 U11415 ( .A(n15258), .B(n15421), .S(n9837), .Z(n9664) );
  NAND2_X1 U11416 ( .A1(n9663), .A2(n9664), .ZN(n9662) );
  MUX2_X1 U11417 ( .A(n15258), .B(n15421), .S(n9857), .Z(n9661) );
  NAND2_X1 U11418 ( .A1(n9662), .A2(n9661), .ZN(n9668) );
  INV_X1 U11419 ( .A(n9663), .ZN(n9666) );
  INV_X1 U11420 ( .A(n9664), .ZN(n9665) );
  NAND2_X1 U11421 ( .A1(n9666), .A2(n9665), .ZN(n9667) );
  NAND2_X1 U11422 ( .A1(n9668), .A2(n9667), .ZN(n9684) );
  NAND2_X1 U11423 ( .A1(n9669), .A2(n14862), .ZN(n9670) );
  AND2_X1 U11424 ( .A1(n9690), .A2(n9670), .ZN(n15222) );
  NAND2_X1 U11425 ( .A1(n15222), .A2(n9705), .ZN(n9676) );
  INV_X1 U11426 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9673) );
  NAND2_X1 U11427 ( .A1(n9803), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9672) );
  NAND2_X1 U11428 ( .A1(n9804), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9671) );
  OAI211_X1 U11429 ( .C1(n9673), .C2(n9808), .A(n9672), .B(n9671), .ZN(n9674)
         );
  INV_X1 U11430 ( .A(n9674), .ZN(n9675) );
  NAND2_X1 U11431 ( .A1(n9676), .A2(n9675), .ZN(n15199) );
  XNOR2_X1 U11432 ( .A(n9678), .B(n9677), .ZN(n13777) );
  NAND2_X1 U11433 ( .A1(n13777), .A2(n9679), .ZN(n9681) );
  NAND2_X1 U11434 ( .A1(n7719), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9680) );
  MUX2_X1 U11435 ( .A(n15199), .B(n12645), .S(n9857), .Z(n9685) );
  NAND2_X1 U11436 ( .A1(n9684), .A2(n9685), .ZN(n9683) );
  MUX2_X1 U11437 ( .A(n15199), .B(n12645), .S(n9837), .Z(n9682) );
  NAND2_X1 U11438 ( .A1(n9683), .A2(n9682), .ZN(n9689) );
  INV_X1 U11439 ( .A(n9684), .ZN(n9687) );
  INV_X1 U11440 ( .A(n9685), .ZN(n9686) );
  NAND2_X1 U11441 ( .A1(n9687), .A2(n9686), .ZN(n9688) );
  AND2_X1 U11442 ( .A1(n9690), .A2(n14919), .ZN(n9691) );
  OR2_X1 U11443 ( .A1(n9691), .A2(n9702), .ZN(n15202) );
  INV_X1 U11444 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9694) );
  NAND2_X1 U11445 ( .A1(n9804), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9693) );
  NAND2_X1 U11446 ( .A1(n9803), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9692) );
  OAI211_X1 U11447 ( .C1(n9808), .C2(n9694), .A(n9693), .B(n9692), .ZN(n9695)
         );
  INV_X1 U11448 ( .A(n9695), .ZN(n9696) );
  OAI21_X1 U11449 ( .B1(n15202), .B2(n9847), .A(n9696), .ZN(n14961) );
  OR2_X1 U11450 ( .A1(n11957), .A2(n10171), .ZN(n9697) );
  XNOR2_X1 U11451 ( .A(n9697), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15921) );
  MUX2_X1 U11452 ( .A(n14961), .B(n15408), .S(n9837), .Z(n9700) );
  MUX2_X1 U11453 ( .A(n15408), .B(n14961), .S(n9837), .Z(n9698) );
  INV_X1 U11454 ( .A(n9700), .ZN(n9701) );
  OR2_X1 U11455 ( .A1(n9702), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9704) );
  AND2_X1 U11456 ( .A1(n9704), .A2(n9703), .ZN(n15187) );
  NAND2_X1 U11457 ( .A1(n15187), .A2(n9705), .ZN(n9711) );
  INV_X1 U11458 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9708) );
  NAND2_X1 U11459 ( .A1(n9803), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9707) );
  NAND2_X1 U11460 ( .A1(n9804), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9706) );
  OAI211_X1 U11461 ( .C1(n9708), .C2(n9808), .A(n9707), .B(n9706), .ZN(n9709)
         );
  INV_X1 U11462 ( .A(n9709), .ZN(n9710) );
  NAND2_X1 U11463 ( .A1(n9711), .A2(n9710), .ZN(n15198) );
  XNOR2_X1 U11464 ( .A(n9713), .B(n9712), .ZN(n13767) );
  NAND2_X1 U11465 ( .A1(n13767), .A2(n9679), .ZN(n9715) );
  NAND2_X1 U11466 ( .A1(n7719), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9714) );
  MUX2_X1 U11467 ( .A(n15198), .B(n15183), .S(n9857), .Z(n9718) );
  MUX2_X1 U11468 ( .A(n15198), .B(n15183), .S(n9837), .Z(n9716) );
  NAND2_X1 U11469 ( .A1(n9717), .A2(n9716), .ZN(n9721) );
  INV_X1 U11470 ( .A(n9718), .ZN(n9719) );
  NAND2_X1 U11471 ( .A1(n7717), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9729) );
  INV_X1 U11472 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n15172) );
  OR2_X1 U11473 ( .A1(n9843), .A2(n15172), .ZN(n9728) );
  OAI21_X1 U11474 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n9723), .A(n9722), .ZN(
        n15168) );
  OR2_X1 U11475 ( .A1(n9724), .A2(n15168), .ZN(n9727) );
  INV_X1 U11476 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9725) );
  OR2_X1 U11477 ( .A1(n9758), .A2(n9725), .ZN(n9726) );
  NAND4_X1 U11478 ( .A1(n9729), .A2(n9728), .A3(n9727), .A4(n9726), .ZN(n15146) );
  XNOR2_X1 U11479 ( .A(n9731), .B(n9730), .ZN(n13812) );
  NAND2_X1 U11480 ( .A1(n13812), .A2(n9679), .ZN(n9733) );
  NAND2_X1 U11481 ( .A1(n7719), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9732) );
  MUX2_X1 U11482 ( .A(n15146), .B(n15395), .S(n9837), .Z(n9737) );
  NAND2_X1 U11483 ( .A1(n9736), .A2(n9737), .ZN(n9735) );
  MUX2_X1 U11484 ( .A(n15146), .B(n15395), .S(n9857), .Z(n9734) );
  NAND2_X1 U11485 ( .A1(n9735), .A2(n9734), .ZN(n9741) );
  INV_X1 U11486 ( .A(n9736), .ZN(n9739) );
  INV_X1 U11487 ( .A(n9737), .ZN(n9738) );
  NAND2_X1 U11488 ( .A1(n9739), .A2(n9738), .ZN(n9740) );
  NAND2_X1 U11489 ( .A1(n7717), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9748) );
  INV_X1 U11490 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9742) );
  OR2_X1 U11491 ( .A1(n9843), .A2(n9742), .ZN(n9747) );
  OAI21_X1 U11492 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n9743), .A(n9755), .ZN(
        n15150) );
  OR2_X1 U11493 ( .A1(n9847), .A2(n15150), .ZN(n9746) );
  INV_X1 U11494 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9744) );
  OR2_X1 U11495 ( .A1(n9758), .A2(n9744), .ZN(n9745) );
  NAND4_X1 U11496 ( .A1(n9748), .A2(n9747), .A3(n9746), .A4(n9745), .ZN(n15132) );
  XNOR2_X1 U11497 ( .A(n9750), .B(n9749), .ZN(n14813) );
  NAND2_X1 U11498 ( .A1(n14813), .A2(n9679), .ZN(n9752) );
  NAND2_X1 U11499 ( .A1(n7719), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9751) );
  MUX2_X1 U11500 ( .A(n15132), .B(n15388), .S(n9857), .Z(n9754) );
  MUX2_X1 U11501 ( .A(n15132), .B(n15388), .S(n9837), .Z(n9753) );
  NAND2_X1 U11502 ( .A1(n7717), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9762) );
  INV_X1 U11503 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n15127) );
  OR2_X1 U11504 ( .A1(n9843), .A2(n15127), .ZN(n9761) );
  INV_X1 U11505 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n14938) );
  NAND2_X1 U11506 ( .A1(n9755), .A2(n14938), .ZN(n9756) );
  NAND2_X1 U11507 ( .A1(n9845), .A2(n9756), .ZN(n15126) );
  OR2_X1 U11508 ( .A1(n9847), .A2(n15126), .ZN(n9760) );
  INV_X1 U11509 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9757) );
  OR2_X1 U11510 ( .A1(n9758), .A2(n9757), .ZN(n9759) );
  NAND4_X1 U11511 ( .A1(n9762), .A2(n9761), .A3(n9760), .A4(n9759), .ZN(n15147) );
  XNOR2_X1 U11512 ( .A(n9764), .B(n9763), .ZN(n14810) );
  NAND2_X1 U11513 ( .A1(n14810), .A2(n9679), .ZN(n9766) );
  NAND2_X1 U11514 ( .A1(n7719), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9765) );
  MUX2_X1 U11515 ( .A(n15147), .B(n15382), .S(n9837), .Z(n9770) );
  NAND2_X1 U11516 ( .A1(n9769), .A2(n9770), .ZN(n9768) );
  MUX2_X1 U11517 ( .A(n15147), .B(n15382), .S(n9857), .Z(n9767) );
  NAND2_X1 U11518 ( .A1(n9768), .A2(n9767), .ZN(n9774) );
  INV_X1 U11519 ( .A(n9769), .ZN(n9772) );
  INV_X1 U11520 ( .A(n9770), .ZN(n9771) );
  NAND2_X1 U11521 ( .A1(n9772), .A2(n9771), .ZN(n9773) );
  NAND2_X1 U11522 ( .A1(n9774), .A2(n9773), .ZN(n9779) );
  INV_X1 U11523 ( .A(n9779), .ZN(n9777) );
  MUX2_X1 U11524 ( .A(n9889), .B(n15133), .S(n9857), .Z(n9775) );
  OAI21_X1 U11525 ( .B1(n9780), .B2(n9779), .A(n9778), .ZN(n9868) );
  INV_X1 U11526 ( .A(n9868), .ZN(n9860) );
  NAND2_X1 U11527 ( .A1(n9783), .A2(SI_27_), .ZN(n9784) );
  MUX2_X1 U11528 ( .A(n12781), .B(n14805), .S(n10197), .Z(n9786) );
  NAND2_X1 U11529 ( .A1(n9786), .A2(n15498), .ZN(n9789) );
  INV_X1 U11530 ( .A(n9786), .ZN(n9787) );
  NAND2_X1 U11531 ( .A1(n9787), .A2(SI_28_), .ZN(n9788) );
  NAND2_X1 U11532 ( .A1(n9789), .A2(n9788), .ZN(n9853) );
  MUX2_X1 U11533 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n10171), .Z(n9790) );
  XNOR2_X1 U11534 ( .A(n9790), .B(n15696), .ZN(n9823) );
  INV_X1 U11535 ( .A(n9790), .ZN(n9791) );
  NAND2_X1 U11536 ( .A1(n9791), .A2(n15696), .ZN(n9792) );
  MUX2_X1 U11537 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n10197), .Z(n9793) );
  NAND2_X1 U11538 ( .A1(n9793), .A2(SI_30_), .ZN(n9830) );
  OAI21_X1 U11539 ( .B1(SI_30_), .B2(n9793), .A(n9830), .ZN(n9794) );
  OR2_X1 U11540 ( .A1(n14186), .A2(n9796), .ZN(n9798) );
  NAND2_X1 U11541 ( .A1(n7719), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9797) );
  INV_X1 U11542 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n15355) );
  NOR2_X1 U11543 ( .A1(n9808), .A2(n15355), .ZN(n9802) );
  INV_X1 U11544 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9799) );
  NOR2_X1 U11545 ( .A1(n9843), .A2(n9799), .ZN(n9801) );
  INV_X1 U11546 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n15478) );
  NOR2_X1 U11547 ( .A1(n9758), .A2(n15478), .ZN(n9800) );
  OR3_X1 U11548 ( .A1(n9802), .A2(n9801), .A3(n9800), .ZN(n14959) );
  NAND2_X1 U11549 ( .A1(n8291), .A2(n9841), .ZN(n9969) );
  INV_X1 U11550 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9807) );
  NAND2_X1 U11551 ( .A1(n9803), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9806) );
  NAND2_X1 U11552 ( .A1(n9804), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n9805) );
  OAI211_X1 U11553 ( .C1(n9808), .C2(n9807), .A(n9806), .B(n9805), .ZN(n15095)
         );
  OAI21_X1 U11554 ( .B1(n14959), .B2(n9969), .A(n15095), .ZN(n9809) );
  INV_X1 U11555 ( .A(n9809), .ZN(n9810) );
  MUX2_X1 U11556 ( .A(n15081), .B(n9810), .S(n9837), .Z(n9862) );
  INV_X1 U11557 ( .A(n9862), .ZN(n9814) );
  OAI21_X1 U11558 ( .B1(n14959), .B2(n9811), .A(n15095), .ZN(n9812) );
  INV_X1 U11559 ( .A(n9812), .ZN(n9813) );
  NAND2_X1 U11560 ( .A1(n9814), .A2(n9861), .ZN(n9873) );
  NAND2_X1 U11561 ( .A1(n7717), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9822) );
  INV_X1 U11562 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9815) );
  OR2_X1 U11563 ( .A1(n9843), .A2(n9815), .ZN(n9821) );
  INV_X1 U11564 ( .A(n9845), .ZN(n9817) );
  AND2_X1 U11565 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n9816) );
  NAND2_X1 U11566 ( .A1(n9817), .A2(n9816), .ZN(n15098) );
  OR2_X1 U11567 ( .A1(n9847), .A2(n15098), .ZN(n9820) );
  INV_X1 U11568 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9818) );
  OR2_X1 U11569 ( .A1(n9758), .A2(n9818), .ZN(n9819) );
  AND4_X1 U11570 ( .A1(n9822), .A2(n9821), .A3(n9820), .A4(n9819), .ZN(n12713)
         );
  NAND2_X1 U11571 ( .A1(n14798), .A2(n9679), .ZN(n9826) );
  NAND2_X1 U11572 ( .A1(n7719), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9825) );
  MUX2_X1 U11573 ( .A(n14960), .B(n15094), .S(n9857), .Z(n9864) );
  INV_X1 U11574 ( .A(n9864), .ZN(n9828) );
  MUX2_X1 U11575 ( .A(n12713), .B(n15366), .S(n9837), .Z(n9865) );
  INV_X1 U11576 ( .A(n9865), .ZN(n9827) );
  NAND2_X1 U11577 ( .A1(n9828), .A2(n9827), .ZN(n9829) );
  NAND2_X1 U11578 ( .A1(n9873), .A2(n9829), .ZN(n9870) );
  XNOR2_X1 U11579 ( .A(n9832), .B(SI_31_), .ZN(n9833) );
  NAND2_X1 U11580 ( .A1(n14792), .A2(n9679), .ZN(n9836) );
  NAND2_X1 U11581 ( .A1(n7719), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n9835) );
  NAND2_X1 U11582 ( .A1(n9837), .A2(n14959), .ZN(n9909) );
  OR2_X1 U11583 ( .A1(n15351), .A2(n9909), .ZN(n9914) );
  INV_X1 U11584 ( .A(n14959), .ZN(n15075) );
  AND2_X1 U11585 ( .A1(n9857), .A2(n15075), .ZN(n9906) );
  NAND2_X1 U11586 ( .A1(n15351), .A2(n9906), .ZN(n9915) );
  NAND2_X1 U11587 ( .A1(n10440), .A2(n15185), .ZN(n10000) );
  NAND2_X1 U11588 ( .A1(n11549), .A2(n9998), .ZN(n9839) );
  NAND2_X1 U11589 ( .A1(n9838), .A2(n9841), .ZN(n10494) );
  NAND2_X1 U11590 ( .A1(n9839), .A2(n10494), .ZN(n9840) );
  AND2_X1 U11591 ( .A1(n10000), .A2(n9840), .ZN(n9916) );
  INV_X1 U11592 ( .A(n9916), .ZN(n9911) );
  INV_X1 U11593 ( .A(n9841), .ZN(n11731) );
  NAND2_X1 U11594 ( .A1(n8291), .A2(n11731), .ZN(n9912) );
  NAND4_X1 U11595 ( .A1(n9914), .A2(n9915), .A3(n9911), .A4(n9912), .ZN(n9876)
         );
  NOR2_X1 U11596 ( .A1(n9870), .A2(n9876), .ZN(n9880) );
  NAND2_X1 U11597 ( .A1(n7717), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9852) );
  INV_X1 U11598 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n12584) );
  OR2_X1 U11599 ( .A1(n9843), .A2(n12584), .ZN(n9851) );
  INV_X1 U11600 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9844) );
  OAI21_X1 U11601 ( .B1(n9845), .B2(n14824), .A(n9844), .ZN(n9846) );
  NAND2_X1 U11602 ( .A1(n9846), .A2(n15098), .ZN(n12711) );
  OR2_X1 U11603 ( .A1(n9847), .A2(n12711), .ZN(n9850) );
  INV_X1 U11604 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9848) );
  OR2_X1 U11605 ( .A1(n9758), .A2(n9848), .ZN(n9849) );
  INV_X1 U11606 ( .A(n15112), .ZN(n15085) );
  NAND2_X1 U11607 ( .A1(n14802), .A2(n9679), .ZN(n9856) );
  NAND2_X1 U11608 ( .A1(n7719), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9855) );
  MUX2_X1 U11609 ( .A(n15085), .B(n15371), .S(n9857), .Z(n9866) );
  INV_X1 U11610 ( .A(n9866), .ZN(n9859) );
  MUX2_X1 U11611 ( .A(n15112), .B(n12707), .S(n9837), .Z(n9867) );
  INV_X1 U11612 ( .A(n9867), .ZN(n9858) );
  NAND2_X1 U11613 ( .A1(n9859), .A2(n9858), .ZN(n9883) );
  XNOR2_X1 U11614 ( .A(n15351), .B(n14959), .ZN(n9903) );
  INV_X1 U11615 ( .A(n9861), .ZN(n9863) );
  NAND2_X1 U11616 ( .A1(n9863), .A2(n9862), .ZN(n9918) );
  AND2_X1 U11617 ( .A1(n9865), .A2(n9864), .ZN(n9874) );
  NOR2_X2 U11618 ( .A1(n9872), .A2(n9874), .ZN(n9882) );
  NAND2_X1 U11619 ( .A1(n9867), .A2(n9866), .ZN(n9869) );
  INV_X1 U11620 ( .A(n9869), .ZN(n9881) );
  INV_X1 U11621 ( .A(n9870), .ZN(n9871) );
  NOR2_X1 U11622 ( .A1(n9872), .A2(n9871), .ZN(n9879) );
  INV_X1 U11623 ( .A(n9873), .ZN(n9877) );
  INV_X1 U11624 ( .A(n9874), .ZN(n9875) );
  NOR3_X1 U11625 ( .A1(n9877), .A2(n9876), .A3(n9875), .ZN(n9878) );
  AOI211_X1 U11626 ( .C1(n9881), .C2(n9880), .A(n9879), .B(n9878), .ZN(n9885)
         );
  INV_X1 U11627 ( .A(n9882), .ZN(n9884) );
  AND2_X1 U11628 ( .A1(n9885), .A2(n8513), .ZN(n9886) );
  INV_X1 U11629 ( .A(n9912), .ZN(n9925) );
  XOR2_X1 U11630 ( .A(n15081), .B(n15095), .Z(n9902) );
  NAND2_X1 U11631 ( .A1(n15371), .A2(n15112), .ZN(n9890) );
  INV_X1 U11632 ( .A(n15198), .ZN(n15163) );
  XNOR2_X1 U11633 ( .A(n15183), .B(n15163), .ZN(n12566) );
  XNOR2_X1 U11634 ( .A(n12645), .B(n15199), .ZN(n15212) );
  INV_X1 U11635 ( .A(n15289), .ZN(n14891) );
  XNOR2_X1 U11636 ( .A(n15435), .B(n14891), .ZN(n15267) );
  INV_X1 U11637 ( .A(n15330), .ZN(n14950) );
  XNOR2_X1 U11638 ( .A(n15446), .B(n14950), .ZN(n15307) );
  INV_X1 U11639 ( .A(n15304), .ZN(n14880) );
  NAND2_X1 U11640 ( .A1(n15440), .A2(n14880), .ZN(n9891) );
  NAND2_X1 U11641 ( .A1(n12558), .A2(n9891), .ZN(n15284) );
  XNOR2_X1 U11642 ( .A(n15451), .B(n15303), .ZN(n15327) );
  XNOR2_X1 U11643 ( .A(n15470), .B(n12312), .ZN(n12157) );
  XNOR2_X1 U11644 ( .A(n12153), .B(n12156), .ZN(n12150) );
  XNOR2_X1 U11645 ( .A(n11963), .B(n11961), .ZN(n11762) );
  XNOR2_X1 U11646 ( .A(n11818), .B(n14967), .ZN(n11820) );
  INV_X1 U11647 ( .A(n14970), .ZN(n11536) );
  XNOR2_X1 U11648 ( .A(n11537), .B(n11536), .ZN(n10889) );
  INV_X1 U11649 ( .A(n14971), .ZN(n10886) );
  XNOR2_X1 U11650 ( .A(n10909), .B(n10886), .ZN(n10862) );
  AND2_X1 U11651 ( .A1(n10522), .A2(n9892), .ZN(n11129) );
  NAND4_X1 U11652 ( .A1(n10524), .A2(n11129), .A3(n11113), .A4(n9974), .ZN(
        n9893) );
  XNOR2_X1 U11653 ( .A(n16446), .B(n10915), .ZN(n11166) );
  NOR4_X1 U11654 ( .A1(n10889), .A2(n10862), .A3(n9893), .A4(n11166), .ZN(
        n9894) );
  XNOR2_X1 U11655 ( .A(n11756), .B(n14968), .ZN(n11745) );
  XNOR2_X1 U11656 ( .A(n16478), .B(n14969), .ZN(n11528) );
  NAND4_X1 U11657 ( .A1(n11820), .A2(n9894), .A3(n11745), .A4(n11528), .ZN(
        n9895) );
  NOR4_X1 U11658 ( .A1(n12157), .A2(n12150), .A3(n11762), .A4(n9895), .ZN(
        n9896) );
  XNOR2_X1 U11659 ( .A(n15456), .B(n15332), .ZN(n12552) );
  XNOR2_X1 U11660 ( .A(n12333), .B(n14962), .ZN(n12331) );
  NAND4_X1 U11661 ( .A1(n15327), .A2(n9896), .A3(n12552), .A4(n12331), .ZN(
        n9897) );
  NOR4_X1 U11662 ( .A1(n15267), .A2(n15307), .A3(n15284), .A4(n9897), .ZN(
        n9898) );
  XNOR2_X1 U11663 ( .A(n15421), .B(n15258), .ZN(n15237) );
  XNOR2_X1 U11664 ( .A(n15257), .B(n15270), .ZN(n15252) );
  NAND4_X1 U11665 ( .A1(n15212), .A2(n9898), .A3(n15237), .A4(n15252), .ZN(
        n9899) );
  NOR3_X1 U11666 ( .A1(n12566), .A2(n15194), .A3(n9899), .ZN(n9900) );
  XNOR2_X1 U11667 ( .A(n15395), .B(n15146), .ZN(n12567) );
  NAND4_X1 U11668 ( .A1(n15130), .A2(n9900), .A3(n15143), .A4(n12567), .ZN(
        n9901) );
  NOR4_X1 U11669 ( .A1(n9902), .A2(n15110), .A3(n15090), .A4(n9901), .ZN(n9904) );
  NAND3_X1 U11670 ( .A1(n9904), .A2(n9903), .A3(n15092), .ZN(n9905) );
  XNOR2_X1 U11671 ( .A(n9905), .B(n12592), .ZN(n9924) );
  INV_X1 U11672 ( .A(n9906), .ZN(n9908) );
  NAND3_X1 U11673 ( .A1(n9908), .A2(n15075), .A3(n9911), .ZN(n9907) );
  OAI21_X1 U11674 ( .B1(n9908), .B2(n9911), .A(n9907), .ZN(n9922) );
  NAND2_X1 U11675 ( .A1(n9911), .A2(n14959), .ZN(n9910) );
  MUX2_X1 U11676 ( .A(n9911), .B(n9910), .S(n9909), .Z(n9913) );
  OAI21_X1 U11677 ( .B1(n15351), .B2(n9913), .A(n9912), .ZN(n9921) );
  INV_X1 U11678 ( .A(n9914), .ZN(n9919) );
  INV_X1 U11679 ( .A(n9915), .ZN(n9917) );
  AOI211_X1 U11680 ( .C1(n15351), .C2(n9922), .A(n9921), .B(n9920), .ZN(n9923)
         );
  AOI21_X1 U11681 ( .B1(n9925), .B2(n9924), .A(n9923), .ZN(n9931) );
  NAND2_X1 U11682 ( .A1(n9929), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9928) );
  MUX2_X1 U11683 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9928), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n9930) );
  NAND2_X1 U11684 ( .A1(n9930), .A2(n7486), .ZN(n10264) );
  NOR2_X1 U11685 ( .A1(n10264), .A2(P1_U3086), .ZN(n12047) );
  NAND2_X1 U11686 ( .A1(n7486), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9932) );
  OAI21_X1 U11687 ( .B1(n9934), .B2(n9933), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9935) );
  MUX2_X1 U11688 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9935), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n9937) );
  NAND2_X1 U11689 ( .A1(n9937), .A2(n9936), .ZN(n15915) );
  INV_X1 U11690 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U11691 ( .A1(n11549), .A2(n12592), .ZN(n9942) );
  INV_X1 U11692 ( .A(n10494), .ZN(n10265) );
  AND2_X1 U11693 ( .A1(n9942), .A2(n10265), .ZN(n10473) );
  INV_X1 U11694 ( .A(n9943), .ZN(n10450) );
  NOR4_X1 U11695 ( .A1(n16258), .A2(n10473), .A3(n15912), .A4(n15230), .ZN(
        n9945) );
  INV_X1 U11696 ( .A(n12047), .ZN(n10263) );
  OAI21_X1 U11697 ( .B1(n10263), .B2(n9838), .A(P1_B_REG_SCAN_IN), .ZN(n9944)
         );
  OR2_X1 U11698 ( .A1(n9945), .A2(n9944), .ZN(n9946) );
  NAND2_X1 U11699 ( .A1(n9947), .A2(n9946), .ZN(P1_U3242) );
  INV_X1 U11700 ( .A(n9948), .ZN(n10258) );
  NOR2_X2 U11701 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n10009) );
  NAND3_X1 U11702 ( .A1(n10009), .A2(n11390), .A3(n9953), .ZN(n9954) );
  NAND2_X1 U11703 ( .A1(n10082), .A2(n9955), .ZN(n10086) );
  NAND2_X1 U11704 ( .A1(n9961), .A2(n10010), .ZN(n9956) );
  OR2_X1 U11705 ( .A1(n9958), .A2(n10011), .ZN(n9959) );
  XNOR2_X1 U11706 ( .A(n9961), .B(P2_IR_REG_24__SCAN_IN), .ZN(n12401) );
  NAND2_X1 U11707 ( .A1(n14809), .A2(n9962), .ZN(n10143) );
  NAND2_X1 U11708 ( .A1(n9963), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9964) );
  XNOR2_X1 U11709 ( .A(n9964), .B(n10012), .ZN(n10268) );
  INV_X1 U11710 ( .A(n10268), .ZN(n12070) );
  INV_X1 U11711 ( .A(n13737), .ZN(n10614) );
  INV_X2 U11712 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  AND2_X1 U11713 ( .A1(n10516), .A2(n11126), .ZN(n9965) );
  OR2_X1 U11714 ( .A1(n9965), .A2(n10528), .ZN(n16395) );
  INV_X1 U11715 ( .A(n16395), .ZN(n9966) );
  XNOR2_X1 U11716 ( .A(n9966), .B(n10517), .ZN(n9967) );
  MUX2_X1 U11717 ( .A(n9967), .B(n9974), .S(n14974), .Z(n9979) );
  NAND2_X1 U11718 ( .A1(n9838), .A2(n15185), .ZN(n9968) );
  AOI22_X1 U11719 ( .A1(n14974), .A2(n15331), .B1(n15329), .B2(n9332), .ZN(
        n9978) );
  INV_X1 U11720 ( .A(n9975), .ZN(n9972) );
  INV_X1 U11721 ( .A(n9970), .ZN(n9971) );
  NAND2_X1 U11722 ( .A1(n9972), .A2(n9971), .ZN(n10519) );
  INV_X1 U11723 ( .A(n10519), .ZN(n9973) );
  AOI21_X1 U11724 ( .B1(n9975), .B2(n9974), .A(n9973), .ZN(n10002) );
  INV_X1 U11725 ( .A(n10002), .ZN(n16398) );
  OAI21_X1 U11726 ( .B1(n10437), .B2(n9976), .A(n12705), .ZN(n11163) );
  NAND2_X1 U11727 ( .A1(n16398), .A2(n15166), .ZN(n9977) );
  OAI211_X1 U11728 ( .C1(n9979), .C2(n16449), .A(n9978), .B(n9977), .ZN(n16396) );
  NAND2_X1 U11729 ( .A1(n15920), .A2(P1_B_REG_SCAN_IN), .ZN(n9980) );
  MUX2_X1 U11730 ( .A(n9980), .B(P1_B_REG_SCAN_IN), .S(n12317), .Z(n9981) );
  OAI22_X1 U11731 ( .A1(n10256), .A2(P1_D_REG_0__SCAN_IN), .B1(n12317), .B2(
        n9982), .ZN(n10407) );
  AND2_X1 U11732 ( .A1(n10407), .A2(n10495), .ZN(n16256) );
  NOR4_X1 U11733 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n9986) );
  NOR4_X1 U11734 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n9985) );
  NOR4_X1 U11735 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n9984) );
  NOR4_X1 U11736 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n9983) );
  NAND4_X1 U11737 ( .A1(n9986), .A2(n9985), .A3(n9984), .A4(n9983), .ZN(n9992)
         );
  NOR2_X1 U11738 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n9990) );
  NOR4_X1 U11739 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n9989) );
  NOR4_X1 U11740 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n9988) );
  NOR4_X1 U11741 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n9987) );
  NAND4_X1 U11742 ( .A1(n9990), .A2(n9989), .A3(n9988), .A4(n9987), .ZN(n9991)
         );
  NOR2_X1 U11743 ( .A1(n9992), .A2(n9991), .ZN(n9993) );
  NOR2_X1 U11744 ( .A1(n10256), .A2(n9993), .ZN(n10406) );
  NOR2_X1 U11745 ( .A1(n10406), .A2(n10473), .ZN(n9994) );
  AND2_X1 U11746 ( .A1(n16256), .A2(n9994), .ZN(n10535) );
  INV_X1 U11747 ( .A(n10256), .ZN(n9996) );
  INV_X1 U11748 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9995) );
  NAND2_X1 U11749 ( .A1(n9996), .A2(n9995), .ZN(n9997) );
  NAND2_X1 U11750 ( .A1(n15920), .A2(n15915), .ZN(n10257) );
  NAND2_X1 U11751 ( .A1(n10535), .A2(n10475), .ZN(n15099) );
  NAND2_X1 U11752 ( .A1(n15471), .A2(n15185), .ZN(n10474) );
  INV_X1 U11753 ( .A(n10474), .ZN(n9999) );
  MUX2_X1 U11754 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n16396), .S(n15338), .Z(
        n10005) );
  INV_X1 U11755 ( .A(n10000), .ZN(n10001) );
  NAND2_X1 U11756 ( .A1(n10491), .A2(n8291), .ZN(n10493) );
  INV_X1 U11757 ( .A(n10493), .ZN(n10478) );
  OAI22_X1 U11758 ( .A1(n15177), .A2(n10002), .B1(n16394), .B2(n15310), .ZN(
        n10004) );
  OAI22_X1 U11759 ( .A1(n15221), .A2(n16395), .B1(n10503), .B2(n15312), .ZN(
        n10003) );
  OR3_X1 U11760 ( .A1(n10005), .A2(n10004), .A3(n10003), .ZN(P1_U3292) );
  NOR2_X1 U11761 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), 
        .ZN(n10008) );
  INV_X1 U11762 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n10006) );
  NAND2_X1 U11763 ( .A1(n10056), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10024) );
  INV_X1 U11764 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10017) );
  INV_X1 U11765 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n11449) );
  OR2_X1 U11766 ( .A1(n13846), .A2(n11449), .ZN(n10022) );
  INV_X1 U11767 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11444) );
  OR2_X1 U11768 ( .A1(n10059), .A2(n11444), .ZN(n10021) );
  NAND2_X1 U11769 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n10030) );
  OAI211_X2 U11770 ( .C1(n14185), .C2(n10228), .A(n10032), .B(n10031), .ZN(
        n13992) );
  NAND2_X1 U11771 ( .A1(n14321), .A2(n13995), .ZN(n10033) );
  INV_X1 U11772 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10276) );
  OR2_X1 U11773 ( .A1(n13846), .A2(n10276), .ZN(n10038) );
  INV_X1 U11774 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10034) );
  NAND2_X1 U11775 ( .A1(n10056), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10036) );
  INV_X1 U11776 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10878) );
  NAND2_X1 U11777 ( .A1(n10197), .A2(SI_0_), .ZN(n10039) );
  XNOR2_X1 U11778 ( .A(n10039), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n14819) );
  NOR2_X1 U11779 ( .A1(n14323), .A2(n13987), .ZN(n11320) );
  NAND2_X1 U11780 ( .A1(n11319), .A2(n10043), .ZN(n11329) );
  NAND2_X1 U11781 ( .A1(n10056), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10047) );
  INV_X1 U11782 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10044) );
  INV_X1 U11783 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n11331) );
  OR2_X1 U11784 ( .A1(n13846), .A2(n11331), .ZN(n10046) );
  INV_X1 U11785 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11334) );
  OR2_X1 U11786 ( .A1(n10059), .A2(n11334), .ZN(n10045) );
  OR2_X1 U11787 ( .A1(n10049), .A2(n7454), .ZN(n10050) );
  INV_X2 U11788 ( .A(n14185), .ZN(n11900) );
  NAND2_X1 U11789 ( .A1(n11329), .A2(n14247), .ZN(n11328) );
  OR2_X1 U11790 ( .A1(n14320), .A2(n16418), .ZN(n10052) );
  NAND2_X1 U11791 ( .A1(n10178), .A2(n11900), .ZN(n10055) );
  NAND2_X1 U11792 ( .A1(n10067), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10054) );
  XNOR2_X1 U11793 ( .A(n10054), .B(P2_IR_REG_3__SCAN_IN), .ZN(n11184) );
  NAND2_X1 U11794 ( .A1(n10056), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10063) );
  INV_X1 U11795 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10058) );
  OR2_X1 U11796 ( .A1(n10986), .A2(n10058), .ZN(n10062) );
  INV_X1 U11797 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n11171) );
  OR2_X1 U11798 ( .A1(n13846), .A2(n11171), .ZN(n10061) );
  OR2_X1 U11799 ( .A1(n10059), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n10060) );
  NAND4_X1 U11800 ( .A1(n10063), .A2(n10062), .A3(n10061), .A4(n10060), .ZN(
        n14319) );
  INV_X1 U11801 ( .A(n14250), .ZN(n10064) );
  NAND2_X1 U11802 ( .A1(n10543), .A2(n10064), .ZN(n10066) );
  INV_X1 U11803 ( .A(n14319), .ZN(n10760) );
  NAND2_X1 U11804 ( .A1(n10760), .A2(n14019), .ZN(n10065) );
  NAND2_X1 U11805 ( .A1(n10066), .A2(n10065), .ZN(n10076) );
  NAND2_X1 U11806 ( .A1(n10192), .A2(n14201), .ZN(n10070) );
  NAND2_X1 U11807 ( .A1(n10201), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10068) );
  XNOR2_X1 U11808 ( .A(n10068), .B(P2_IR_REG_4__SCAN_IN), .ZN(n11186) );
  AOI22_X1 U11809 ( .A1(n7465), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n10048), 
        .B2(n11186), .ZN(n10069) );
  NAND2_X1 U11810 ( .A1(n13902), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10075) );
  INV_X1 U11811 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10071) );
  OR2_X1 U11812 ( .A1(n10986), .A2(n10071), .ZN(n10074) );
  NAND2_X1 U11813 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n10094) );
  OAI21_X1 U11814 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n10094), .ZN(n12775) );
  OR2_X1 U11815 ( .A1(n10059), .A2(n12775), .ZN(n10073) );
  INV_X2 U11816 ( .A(n12022), .ZN(n14192) );
  INV_X1 U11817 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11172) );
  OR2_X1 U11818 ( .A1(n14192), .A2(n11172), .ZN(n10072) );
  NAND2_X1 U11819 ( .A1(n10076), .A2(n14252), .ZN(n10801) );
  OAI21_X1 U11820 ( .B1(n10076), .B2(n14252), .A(n10801), .ZN(n10101) );
  INV_X1 U11821 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n10077) );
  NAND2_X1 U11822 ( .A1(n11390), .A2(n10077), .ZN(n10078) );
  INV_X1 U11823 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n10079) );
  NAND2_X1 U11824 ( .A1(n10089), .A2(n10079), .ZN(n10081) );
  NAND2_X1 U11825 ( .A1(n10085), .A2(n9953), .ZN(n10083) );
  NAND2_X1 U11826 ( .A1(n10086), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10088) );
  XNOR2_X1 U11827 ( .A(n10089), .B(P2_IR_REG_19__SCAN_IN), .ZN(n10130) );
  OR2_X1 U11828 ( .A1(n11958), .A2(n14366), .ZN(n10090) );
  NAND2_X1 U11829 ( .A1(n13902), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10099) );
  INV_X1 U11830 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10091) );
  OR2_X1 U11831 ( .A1(n10986), .A2(n10091), .ZN(n10098) );
  INV_X1 U11832 ( .A(n10094), .ZN(n10092) );
  NAND2_X1 U11833 ( .A1(n10092), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10566) );
  INV_X1 U11834 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10093) );
  NAND2_X1 U11835 ( .A1(n10094), .A2(n10093), .ZN(n10095) );
  NAND2_X1 U11836 ( .A1(n10566), .A2(n10095), .ZN(n11479) );
  OR2_X1 U11837 ( .A1(n10059), .A2(n11479), .ZN(n10097) );
  INV_X1 U11838 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11480) );
  OR2_X1 U11839 ( .A1(n13846), .A2(n11480), .ZN(n10096) );
  NAND4_X1 U11840 ( .A1(n10099), .A2(n10098), .A3(n10097), .A4(n10096), .ZN(
        n14317) );
  INV_X1 U11841 ( .A(n14317), .ZN(n10803) );
  INV_X1 U11842 ( .A(n11958), .ZN(n14295) );
  NAND2_X1 U11843 ( .A1(n10269), .A2(n10278), .ZN(n14374) );
  INV_X1 U11844 ( .A(n10278), .ZN(n10100) );
  AND2_X2 U11845 ( .A1(n10269), .A2(n10100), .ZN(n14613) );
  INV_X1 U11846 ( .A(n14613), .ZN(n13941) );
  OAI22_X1 U11847 ( .A1(n10803), .A2(n14374), .B1(n10760), .B2(n13941), .ZN(
        n12772) );
  AOI21_X1 U11848 ( .B1(n10101), .B2(n7449), .A(n12772), .ZN(n10813) );
  INV_X1 U11849 ( .A(n10813), .ZN(n10118) );
  AND2_X1 U11850 ( .A1(n10268), .A2(P2_STATE_REG_SCAN_IN), .ZN(n16082) );
  NAND2_X1 U11851 ( .A1(n14282), .A2(n14366), .ZN(n14290) );
  NAND2_X1 U11852 ( .A1(n10269), .A2(n14290), .ZN(n10142) );
  NAND2_X1 U11853 ( .A1(n16076), .A2(n10142), .ZN(n10636) );
  INV_X1 U11854 ( .A(n10636), .ZN(n10509) );
  NOR2_X1 U11855 ( .A1(n14809), .A2(n12401), .ZN(n16083) );
  INV_X1 U11856 ( .A(n16083), .ZN(n10105) );
  INV_X1 U11857 ( .A(P2_B_REG_SCAN_IN), .ZN(n14372) );
  XOR2_X1 U11858 ( .A(n14372), .B(n12401), .Z(n10102) );
  OR2_X1 U11859 ( .A1(n14814), .A2(n10102), .ZN(n10103) );
  INV_X1 U11860 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n16081) );
  NAND2_X1 U11861 ( .A1(n16074), .A2(n16081), .ZN(n10104) );
  NAND2_X1 U11862 ( .A1(n10105), .A2(n10104), .ZN(n10637) );
  INV_X1 U11863 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n16077) );
  NOR2_X1 U11864 ( .A1(n14814), .A2(n14809), .ZN(n16078) );
  AOI21_X1 U11865 ( .B1(n16077), .B2(n16074), .A(n16078), .ZN(n10507) );
  NOR4_X1 U11866 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n10109) );
  NOR4_X1 U11867 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n10108) );
  NOR4_X1 U11868 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n10107) );
  NOR4_X1 U11869 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n10106) );
  NAND4_X1 U11870 ( .A1(n10109), .A2(n10108), .A3(n10107), .A4(n10106), .ZN(
        n10115) );
  NOR2_X1 U11871 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n10113) );
  NOR4_X1 U11872 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n10112) );
  NOR4_X1 U11873 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n10111) );
  NOR4_X1 U11874 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n10110) );
  NAND4_X1 U11875 ( .A1(n10113), .A2(n10112), .A3(n10111), .A4(n10110), .ZN(
        n10114) );
  OAI21_X1 U11876 ( .B1(n10115), .B2(n10114), .A(n16074), .ZN(n10506) );
  NAND2_X1 U11877 ( .A1(n10507), .A2(n10506), .ZN(n10141) );
  INV_X1 U11878 ( .A(n10141), .ZN(n10116) );
  NAND3_X1 U11879 ( .A1(n10509), .A2(n10637), .A3(n10116), .ZN(n10131) );
  MUX2_X1 U11880 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10118), .S(n14644), .Z(
        n10140) );
  NAND2_X1 U11881 ( .A1(n14323), .A2(n13951), .ZN(n11316) );
  INV_X1 U11882 ( .A(n11316), .ZN(n10119) );
  NAND2_X1 U11883 ( .A1(n11327), .A2(n10120), .ZN(n10122) );
  OR2_X1 U11884 ( .A1(n14320), .A2(n14005), .ZN(n10121) );
  NAND2_X1 U11885 ( .A1(n10122), .A2(n10121), .ZN(n10539) );
  NAND2_X1 U11886 ( .A1(n10539), .A2(n14250), .ZN(n10124) );
  OR2_X1 U11887 ( .A1(n14319), .A2(n14019), .ZN(n10123) );
  NAND2_X1 U11888 ( .A1(n10124), .A2(n10123), .ZN(n10795) );
  XNOR2_X1 U11889 ( .A(n10795), .B(n14252), .ZN(n10814) );
  NOR2_X1 U11890 ( .A1(n10126), .A2(n11958), .ZN(n10127) );
  AND2_X1 U11891 ( .A1(n14282), .A2(n10130), .ZN(n14296) );
  NAND2_X1 U11892 ( .A1(n14296), .A2(n10125), .ZN(n10873) );
  NAND2_X1 U11893 ( .A1(n8139), .A2(n10873), .ZN(n10129) );
  NOR2_X1 U11894 ( .A1(n10814), .A2(n14604), .ZN(n10139) );
  NAND2_X1 U11895 ( .A1(n10540), .A2(n14026), .ZN(n10132) );
  NAND2_X1 U11896 ( .A1(n10132), .A2(n14594), .ZN(n10133) );
  NOR2_X1 U11897 ( .A1(n10837), .A2(n10133), .ZN(n10811) );
  INV_X1 U11898 ( .A(n10811), .ZN(n10134) );
  NOR2_X1 U11899 ( .A1(n14553), .A2(n10134), .ZN(n10138) );
  INV_X1 U11900 ( .A(n14282), .ZN(n14248) );
  NAND2_X1 U11901 ( .A1(n10513), .A2(n14248), .ZN(n10161) );
  INV_X1 U11902 ( .A(n10161), .ZN(n10135) );
  INV_X1 U11903 ( .A(n14026), .ZN(n10136) );
  OAI22_X1 U11904 ( .A1(n14622), .A2(n10136), .B1(n14641), .B2(n12775), .ZN(
        n10137) );
  OR4_X1 U11905 ( .A1(n10140), .A2(n10139), .A3(n10138), .A4(n10137), .ZN(
        P2_U3261) );
  OR2_X1 U11906 ( .A1(n10637), .A2(n10141), .ZN(n10156) );
  NAND2_X1 U11907 ( .A1(n10156), .A2(n10505), .ZN(n10145) );
  AND3_X1 U11908 ( .A1(n10143), .A2(n10268), .A3(n10142), .ZN(n10144) );
  NAND2_X1 U11909 ( .A1(n10145), .A2(n10144), .ZN(n10660) );
  MUX2_X1 U11910 ( .A(n13972), .B(P2_U3088), .S(P2_REG3_REG_3__SCAN_IN), .Z(
        n10166) );
  INV_X1 U11911 ( .A(n10126), .ZN(n13986) );
  XNOR2_X1 U11912 ( .A(n7463), .B(n14019), .ZN(n12768) );
  AND2_X1 U11913 ( .A1(n14319), .A2(n7458), .ZN(n10146) );
  NAND2_X1 U11914 ( .A1(n12768), .A2(n10146), .ZN(n10548) );
  OR2_X1 U11915 ( .A1(n12768), .A2(n10146), .ZN(n10147) );
  NAND2_X1 U11916 ( .A1(n10548), .A2(n10147), .ZN(n10160) );
  NAND2_X1 U11917 ( .A1(n14321), .A2(n10148), .ZN(n10150) );
  XNOR2_X1 U11918 ( .A(n10763), .B(n10150), .ZN(n10664) );
  INV_X1 U11919 ( .A(n7462), .ZN(n13816) );
  AND2_X1 U11920 ( .A1(n13816), .A2(n13987), .ZN(n10658) );
  NOR2_X1 U11921 ( .A1(n11316), .A2(n14594), .ZN(n10149) );
  NAND2_X1 U11922 ( .A1(n10763), .A2(n10150), .ZN(n10151) );
  XNOR2_X1 U11923 ( .A(n7463), .B(n14005), .ZN(n10152) );
  NAND2_X1 U11924 ( .A1(n14320), .A2(n10148), .ZN(n10153) );
  XNOR2_X1 U11925 ( .A(n10152), .B(n10153), .ZN(n10764) );
  INV_X1 U11926 ( .A(n10152), .ZN(n10154) );
  NAND2_X1 U11927 ( .A1(n10154), .A2(n10153), .ZN(n10155) );
  INV_X1 U11928 ( .A(n10156), .ZN(n10157) );
  NAND2_X1 U11929 ( .A1(n10157), .A2(n16076), .ZN(n10163) );
  OR3_X2 U11930 ( .A1(n10163), .A2(n10269), .A3(n14709), .ZN(n13915) );
  INV_X1 U11931 ( .A(n12770), .ZN(n10158) );
  AOI211_X1 U11932 ( .C1(n10160), .C2(n10159), .A(n13915), .B(n10158), .ZN(
        n10165) );
  OR2_X1 U11933 ( .A1(n10163), .A2(n10161), .ZN(n10162) );
  AOI22_X1 U11934 ( .A1(n14614), .A2(n14318), .B1(n14320), .B2(n14613), .ZN(
        n10544) );
  OAI22_X1 U11935 ( .A1(n13966), .A2(n10542), .B1(n10544), .B2(n13975), .ZN(
        n10164) );
  OR3_X1 U11936 ( .A1(n10166), .A2(n10165), .A3(n10164), .ZN(P2_U3190) );
  MUX2_X1 U11937 ( .A(P2_RD_REG_SCAN_IN), .B(n8548), .S(P1_RD_REG_SCAN_IN), 
        .Z(n10168) );
  INV_X1 U11938 ( .A(P3_RD_REG_SCAN_IN), .ZN(n10167) );
  NAND2_X1 U11939 ( .A1(n10168), .A2(n10167), .ZN(U29) );
  INV_X1 U11940 ( .A(n13739), .ZN(n13750) );
  NAND2_X1 U11941 ( .A1(n10197), .A2(P3_U3151), .ZN(n13745) );
  OAI222_X1 U11942 ( .A1(P3_U3151), .A2(n11418), .B1(n13750), .B2(n10170), 
        .C1(n10169), .C2(n13745), .ZN(P3_U3289) );
  NAND2_X2 U11943 ( .A1(n10171), .A2(P2_U3088), .ZN(n14816) );
  OAI222_X1 U11944 ( .A1(n14818), .A2(n10172), .B1(n14816), .B2(n10228), .C1(
        n8493), .C2(P2_U3088), .ZN(P2_U3326) );
  OAI222_X1 U11945 ( .A1(n13750), .A2(n10174), .B1(n13745), .B2(n10173), .C1(
        P3_U3151), .C2(n11431), .ZN(P3_U3287) );
  OAI222_X1 U11946 ( .A1(P3_U3151), .A2(n10177), .B1(n13750), .B2(n10176), 
        .C1(n10175), .C2(n13745), .ZN(P3_U3295) );
  INV_X1 U11947 ( .A(n10178), .ZN(n10199) );
  INV_X1 U11948 ( .A(n11184), .ZN(n16117) );
  OAI222_X1 U11949 ( .A1(n14818), .A2(n10179), .B1(n14816), .B2(n10199), .C1(
        P2_U3088), .C2(n16117), .ZN(P2_U3324) );
  INV_X1 U11950 ( .A(n10180), .ZN(n10230) );
  INV_X1 U11951 ( .A(n16107), .ZN(n11170) );
  OAI222_X1 U11952 ( .A1(n14818), .A2(n10181), .B1(n14816), .B2(n10230), .C1(
        P2_U3088), .C2(n11170), .ZN(P2_U3325) );
  INV_X1 U11953 ( .A(n13745), .ZN(n10360) );
  AOI222_X1 U11954 ( .A1(n10182), .A2(n13739), .B1(SI_7_), .B2(n10360), .C1(
        n11258), .C2(P3_STATE_REG_SCAN_IN), .ZN(n10183) );
  INV_X1 U11955 ( .A(n10183), .ZN(P3_U3288) );
  INV_X1 U11956 ( .A(n10185), .ZN(P3_U3293) );
  AOI222_X1 U11957 ( .A1(n10186), .A2(n13739), .B1(n11008), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_3_), .C2(n10360), .ZN(n10187) );
  INV_X1 U11958 ( .A(n10187), .ZN(P3_U3292) );
  AOI222_X1 U11959 ( .A1(n10188), .A2(n13739), .B1(n11029), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_5_), .C2(n10360), .ZN(n10189) );
  INV_X1 U11960 ( .A(n10189), .ZN(P3_U3290) );
  AOI222_X1 U11961 ( .A1(n10190), .A2(n13739), .B1(n11015), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_4_), .C2(n10360), .ZN(n10191) );
  INV_X1 U11962 ( .A(n10191), .ZN(P3_U3291) );
  INV_X1 U11963 ( .A(n10192), .ZN(n10224) );
  INV_X1 U11964 ( .A(n11186), .ZN(n16129) );
  OAI222_X1 U11965 ( .A1(n14818), .A2(n10193), .B1(n14816), .B2(n10224), .C1(
        P2_U3088), .C2(n16129), .ZN(P2_U3323) );
  AOI222_X1 U11966 ( .A1(n10194), .A2(n13739), .B1(SI_9_), .B2(n10360), .C1(
        n11439), .C2(P3_STATE_REG_SCAN_IN), .ZN(n10195) );
  INV_X1 U11967 ( .A(n10195), .ZN(P3_U3286) );
  INV_X1 U11968 ( .A(n14993), .ZN(n10200) );
  OAI222_X1 U11969 ( .A1(n10200), .A2(P1_U3086), .B1(n15919), .B2(n10199), 
        .C1(n10198), .C2(n15916), .ZN(P1_U3352) );
  INV_X1 U11970 ( .A(n10552), .ZN(n10226) );
  NOR2_X1 U11971 ( .A1(n10204), .A2(n10335), .ZN(n10202) );
  MUX2_X1 U11972 ( .A(n10335), .B(n10202), .S(P2_IR_REG_5__SCAN_IN), .Z(n10205) );
  OR2_X1 U11973 ( .A1(n10205), .A2(n10218), .ZN(n16141) );
  OAI222_X1 U11974 ( .A1(n14818), .A2(n10206), .B1(n14816), .B2(n10226), .C1(
        P2_U3088), .C2(n16141), .ZN(P2_U3322) );
  INV_X1 U11975 ( .A(n12196), .ZN(n11995) );
  OAI222_X1 U11976 ( .A1(P3_U3151), .A2(n11995), .B1(n13745), .B2(n10208), 
        .C1(n13750), .C2(n10207), .ZN(P3_U3284) );
  AOI222_X1 U11977 ( .A1(n10209), .A2(n13739), .B1(SI_10_), .B2(n10360), .C1(
        n11850), .C2(P3_STATE_REG_SCAN_IN), .ZN(n10210) );
  INV_X1 U11978 ( .A(n10210), .ZN(P3_U3285) );
  INV_X1 U11979 ( .A(n10351), .ZN(n10212) );
  INV_X1 U11980 ( .A(n10560), .ZN(n10214) );
  OAI222_X1 U11981 ( .A1(n10212), .A2(P1_U3086), .B1(n15919), .B2(n10214), 
        .C1(n10211), .C2(n15916), .ZN(P1_U3349) );
  OR2_X1 U11982 ( .A1(n10218), .A2(n10335), .ZN(n10213) );
  XNOR2_X1 U11983 ( .A(n10213), .B(P2_IR_REG_6__SCAN_IN), .ZN(n16156) );
  INV_X1 U11984 ( .A(n16156), .ZN(n11173) );
  OAI222_X1 U11985 ( .A1(n14818), .A2(n10215), .B1(n14816), .B2(n10214), .C1(
        P2_U3088), .C2(n11173), .ZN(P2_U3321) );
  OAI222_X1 U11986 ( .A1(P3_U3151), .A2(n12294), .B1(n13745), .B2(n15728), 
        .C1(n13750), .C2(n10216), .ZN(P3_U3283) );
  INV_X1 U11987 ( .A(n10723), .ZN(n10221) );
  NAND2_X1 U11988 ( .A1(n10218), .A2(n10217), .ZN(n10234) );
  NAND2_X1 U11989 ( .A1(n10234), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10219) );
  XNOR2_X1 U11990 ( .A(n10219), .B(P2_IR_REG_7__SCAN_IN), .ZN(n14331) );
  INV_X1 U11991 ( .A(n14331), .ZN(n11175) );
  OAI222_X1 U11992 ( .A1(n14818), .A2(n10220), .B1(n14816), .B2(n10221), .C1(
        P2_U3088), .C2(n11175), .ZN(P2_U3320) );
  INV_X1 U11993 ( .A(n10384), .ZN(n10359) );
  OAI222_X1 U11994 ( .A1(n15916), .A2(n10222), .B1(n15919), .B2(n10221), .C1(
        n10359), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U11995 ( .A(n16341), .ZN(n16357) );
  OAI222_X1 U11996 ( .A1(n16357), .A2(P1_U3086), .B1(n15919), .B2(n10224), 
        .C1(n10223), .C2(n15916), .ZN(P1_U3351) );
  INV_X1 U11997 ( .A(n10370), .ZN(n10227) );
  OAI222_X1 U11998 ( .A1(n10227), .A2(P1_U3086), .B1(n15919), .B2(n10226), 
        .C1(n10225), .C2(n15916), .ZN(P1_U3350) );
  OAI222_X1 U11999 ( .A1(P1_U3086), .A2(n9285), .B1(n15919), .B2(n10228), .C1(
        n7732), .C2(n15916), .ZN(P1_U3354) );
  INV_X1 U12000 ( .A(n10461), .ZN(n10231) );
  OAI222_X1 U12001 ( .A1(n10231), .A2(P1_U3086), .B1(n15919), .B2(n10230), 
        .C1(n10229), .C2(n15916), .ZN(P1_U3353) );
  INV_X1 U12002 ( .A(n15007), .ZN(n10233) );
  INV_X1 U12003 ( .A(n10730), .ZN(n10236) );
  OAI222_X1 U12004 ( .A1(n10233), .A2(P1_U3086), .B1(n15919), .B2(n10236), 
        .C1(n10232), .C2(n15916), .ZN(P1_U3347) );
  NAND2_X1 U12005 ( .A1(n10238), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10235) );
  XNOR2_X1 U12006 ( .A(n10235), .B(P2_IR_REG_8__SCAN_IN), .ZN(n16169) );
  INV_X1 U12007 ( .A(n16169), .ZN(n11176) );
  OAI222_X1 U12008 ( .A1(n14818), .A2(n10237), .B1(n14816), .B2(n10236), .C1(
        P2_U3088), .C2(n11176), .ZN(P2_U3319) );
  INV_X1 U12009 ( .A(n10978), .ZN(n10242) );
  NAND2_X1 U12010 ( .A1(n10245), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10239) );
  XNOR2_X1 U12011 ( .A(n10239), .B(P2_IR_REG_9__SCAN_IN), .ZN(n11192) );
  INV_X1 U12012 ( .A(n11192), .ZN(n16238) );
  OAI222_X1 U12013 ( .A1(n14818), .A2(n10240), .B1(n14816), .B2(n10242), .C1(
        P2_U3088), .C2(n16238), .ZN(P2_U3318) );
  INV_X1 U12014 ( .A(n15024), .ZN(n10243) );
  OAI222_X1 U12015 ( .A1(n10243), .A2(P1_U3086), .B1(n15919), .B2(n10242), 
        .C1(n10241), .C2(n15916), .ZN(P1_U3346) );
  OAI222_X1 U12016 ( .A1(P3_U3151), .A2(n13234), .B1(n13745), .B2(n15724), 
        .C1(n13750), .C2(n10244), .ZN(P3_U3282) );
  INV_X1 U12017 ( .A(n11341), .ZN(n10249) );
  OR2_X1 U12018 ( .A1(n10252), .A2(n10335), .ZN(n10246) );
  XNOR2_X1 U12019 ( .A(n10246), .B(P2_IR_REG_10__SCAN_IN), .ZN(n16233) );
  INV_X1 U12020 ( .A(n16233), .ZN(n11179) );
  OAI222_X1 U12021 ( .A1(n14818), .A2(n10247), .B1(n14816), .B2(n10249), .C1(
        P2_U3088), .C2(n11179), .ZN(P2_U3317) );
  INV_X1 U12022 ( .A(n10425), .ZN(n10397) );
  OAI222_X1 U12023 ( .A1(n10397), .A2(P1_U3086), .B1(n15919), .B2(n10249), 
        .C1(n10248), .C2(n15916), .ZN(P1_U3345) );
  AND2_X1 U12024 ( .A1(n10377), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12025 ( .A1(n10377), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12026 ( .A1(n10377), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12027 ( .A1(n10377), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12028 ( .A1(n10377), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12029 ( .A1(n10377), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12030 ( .A1(n10377), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12031 ( .A1(n10377), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12032 ( .A1(n10377), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12033 ( .A1(n10377), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U12034 ( .A1(n10377), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  INV_X1 U12035 ( .A(n15039), .ZN(n10421) );
  INV_X1 U12036 ( .A(n11603), .ZN(n10254) );
  OAI222_X1 U12037 ( .A1(n10421), .A2(P1_U3086), .B1(n15919), .B2(n10254), 
        .C1(n10250), .C2(n15916), .ZN(P1_U3344) );
  INV_X1 U12038 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n10251) );
  NAND2_X1 U12039 ( .A1(n10252), .A2(n10251), .ZN(n10288) );
  NAND2_X1 U12040 ( .A1(n10288), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10253) );
  XNOR2_X1 U12041 ( .A(n10253), .B(P2_IR_REG_11__SCAN_IN), .ZN(n16181) );
  INV_X1 U12042 ( .A(n16181), .ZN(n11180) );
  OAI222_X1 U12043 ( .A1(n14818), .A2(n10255), .B1(n14816), .B2(n10254), .C1(
        P2_U3088), .C2(n11180), .ZN(P2_U3316) );
  AND2_X2 U12044 ( .A1(n10256), .A2(n10495), .ZN(n16073) );
  OAI22_X1 U12045 ( .A1(n16073), .A2(P1_D_REG_1__SCAN_IN), .B1(n10258), .B2(
        n10257), .ZN(n10259) );
  INV_X1 U12046 ( .A(n10259), .ZN(P1_U3446) );
  OAI222_X1 U12047 ( .A1(P3_U3151), .A2(n13268), .B1(n13745), .B2(n15525), 
        .C1(n13750), .C2(n10260), .ZN(P3_U3281) );
  AOI22_X1 U12048 ( .A1(n13292), .A2(P3_STATE_REG_SCAN_IN), .B1(SI_15_), .B2(
        n10360), .ZN(n10261) );
  OAI21_X1 U12049 ( .B1(n10262), .B2(n13750), .A(n10261), .ZN(P3_U3280) );
  NAND2_X1 U12050 ( .A1(n16258), .A2(n10263), .ZN(n10294) );
  NAND2_X1 U12051 ( .A1(n10265), .A2(n10264), .ZN(n10267) );
  NAND2_X1 U12052 ( .A1(n10267), .A2(n10266), .ZN(n10292) );
  NAND2_X1 U12053 ( .A1(n10294), .A2(n10292), .ZN(n16364) );
  NOR2_X1 U12054 ( .A1(n14978), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12055 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10277) );
  NAND2_X1 U12056 ( .A1(n10269), .A2(n10268), .ZN(n10270) );
  NAND2_X1 U12057 ( .A1(n10272), .A2(n10271), .ZN(n10283) );
  OR2_X1 U12058 ( .A1(n10278), .A2(P2_U3088), .ZN(n14803) );
  INV_X1 U12059 ( .A(n14803), .ZN(n10274) );
  NAND2_X1 U12060 ( .A1(n10275), .A2(n14807), .ZN(n16228) );
  INV_X1 U12061 ( .A(n14807), .ZN(n14292) );
  NAND2_X1 U12062 ( .A1(n10275), .A2(n14292), .ZN(n16247) );
  OAI22_X1 U12063 ( .A1(n10277), .A2(n16228), .B1(n16247), .B2(n10276), .ZN(
        n10282) );
  INV_X1 U12064 ( .A(n16247), .ZN(n16222) );
  NAND2_X1 U12065 ( .A1(n16222), .A2(n10276), .ZN(n10280) );
  INV_X1 U12066 ( .A(n16228), .ZN(n16250) );
  NAND2_X1 U12067 ( .A1(n16250), .A2(n10277), .ZN(n10279) );
  AND2_X1 U12068 ( .A1(n10278), .A2(n10283), .ZN(n16237) );
  NAND3_X1 U12069 ( .A1(n10280), .A2(n10279), .A3(n16189), .ZN(n10281) );
  MUX2_X1 U12070 ( .A(n10282), .B(n10281), .S(P2_IR_REG_0__SCAN_IN), .Z(n10286) );
  NOR2_X1 U12071 ( .A1(n10283), .A2(P2_U3088), .ZN(n16097) );
  INV_X1 U12072 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10284) );
  OAI22_X1 U12073 ( .A1(n16254), .A2(n10284), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10878), .ZN(n10285) );
  OR2_X1 U12074 ( .A1(n10286), .A2(n10285), .ZN(P2_U3214) );
  INV_X1 U12075 ( .A(n10666), .ZN(n10673) );
  INV_X1 U12076 ( .A(n11774), .ZN(n10290) );
  OAI222_X1 U12077 ( .A1(P1_U3086), .A2(n10673), .B1(n15919), .B2(n10290), 
        .C1(n10287), .C2(n15916), .ZN(P1_U3343) );
  NAND2_X1 U12078 ( .A1(n10333), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10289) );
  XNOR2_X1 U12079 ( .A(n10289), .B(P2_IR_REG_12__SCAN_IN), .ZN(n11775) );
  INV_X1 U12080 ( .A(n11775), .ZN(n11198) );
  OAI222_X1 U12081 ( .A1(n14818), .A2(n10291), .B1(n14816), .B2(n10290), .C1(
        n11198), .C2(P2_U3088), .ZN(P2_U3315) );
  INV_X1 U12082 ( .A(n10292), .ZN(n10293) );
  AND2_X1 U12083 ( .A1(n10294), .A2(n10293), .ZN(n10302) );
  INV_X1 U12084 ( .A(n10302), .ZN(n10314) );
  NOR2_X1 U12085 ( .A1(n15912), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10295) );
  NOR2_X1 U12086 ( .A1(n9943), .A2(n10295), .ZN(n10448) );
  INV_X1 U12087 ( .A(n15912), .ZN(n15073) );
  OAI21_X1 U12088 ( .B1(n15073), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10448), .ZN(
        n10296) );
  MUX2_X1 U12089 ( .A(n10448), .B(n10296), .S(n7998), .Z(n10297) );
  OAI22_X1 U12090 ( .A1(n10314), .A2(n10297), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11123), .ZN(n10299) );
  NAND2_X1 U12091 ( .A1(n10302), .A2(n15912), .ZN(n16266) );
  NOR3_X1 U12092 ( .A1(n16266), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n7998), .ZN(
        n10298) );
  AOI211_X1 U12093 ( .C1(n14978), .C2(P1_ADDR_REG_0__SCAN_IN), .A(n10299), .B(
        n10298), .ZN(n10300) );
  INV_X1 U12094 ( .A(n10300), .ZN(P1_U3243) );
  INV_X1 U12095 ( .A(n13296), .ZN(n13316) );
  OAI222_X1 U12096 ( .A1(P3_U3151), .A2(n13316), .B1(n13745), .B2(n15520), 
        .C1(n13750), .C2(n10301), .ZN(P3_U3279) );
  AND2_X1 U12097 ( .A1(n10302), .A2(n9943), .ZN(n15065) );
  INV_X1 U12098 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n15936) );
  NAND2_X1 U12099 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n11150) );
  OAI21_X1 U12100 ( .B1(n16364), .B2(n15936), .A(n11150), .ZN(n10313) );
  MUX2_X1 U12101 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10303), .S(n10461), .Z(
        n10306) );
  INV_X1 U12102 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10304) );
  MUX2_X1 U12103 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n10304), .S(n14982), .Z(
        n14980) );
  AND2_X1 U12104 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14981) );
  NAND2_X1 U12105 ( .A1(n14980), .A2(n14981), .ZN(n14979) );
  NAND2_X1 U12106 ( .A1(n14982), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10452) );
  NAND2_X1 U12107 ( .A1(n14979), .A2(n10452), .ZN(n10305) );
  NAND2_X1 U12108 ( .A1(n10461), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14994) );
  NAND2_X1 U12109 ( .A1(n14996), .A2(n14994), .ZN(n10309) );
  MUX2_X1 U12110 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10307), .S(n14993), .Z(
        n10308) );
  NAND2_X1 U12111 ( .A1(n10309), .A2(n10308), .ZN(n16351) );
  NAND2_X1 U12112 ( .A1(n14993), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n16350) );
  MUX2_X1 U12113 ( .A(n9343), .B(P1_REG1_REG_4__SCAN_IN), .S(n16341), .Z(
        n16349) );
  AOI21_X1 U12114 ( .B1(n16351), .B2(n16350), .A(n16349), .ZN(n16348) );
  MUX2_X1 U12115 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9367), .S(n10370), .Z(
        n10365) );
  NAND2_X1 U12116 ( .A1(n10364), .A2(n10365), .ZN(n10363) );
  OAI21_X1 U12117 ( .B1(n10370), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10363), .ZN(
        n10311) );
  INV_X1 U12118 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10901) );
  MUX2_X1 U12119 ( .A(n10901), .B(P1_REG1_REG_6__SCAN_IN), .S(n10351), .Z(
        n10310) );
  NOR2_X1 U12120 ( .A1(n10311), .A2(n10310), .ZN(n10350) );
  AOI211_X1 U12121 ( .C1(n10311), .C2(n10310), .A(n10350), .B(n16266), .ZN(
        n10312) );
  AOI211_X1 U12122 ( .C1(n15065), .C2(n10351), .A(n10313), .B(n10312), .ZN(
        n10332) );
  NOR2_X1 U12123 ( .A1(n10314), .A2(n15912), .ZN(n15067) );
  AND2_X1 U12124 ( .A1(n15067), .A2(n10450), .ZN(n16347) );
  MUX2_X1 U12125 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n15340), .S(n10461), .Z(
        n10318) );
  MUX2_X1 U12126 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n10315), .S(n14982), .Z(
        n14977) );
  AND2_X1 U12127 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10316) );
  NAND2_X1 U12128 ( .A1(n14977), .A2(n10316), .ZN(n14976) );
  NAND2_X1 U12129 ( .A1(n14982), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10455) );
  NAND2_X1 U12130 ( .A1(n14976), .A2(n10455), .ZN(n10317) );
  NAND2_X1 U12131 ( .A1(n10318), .A2(n10317), .ZN(n14989) );
  NAND2_X1 U12132 ( .A1(n10461), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14987) );
  NAND2_X1 U12133 ( .A1(n14989), .A2(n14987), .ZN(n10320) );
  INV_X1 U12134 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n11119) );
  MUX2_X1 U12135 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n11119), .S(n14993), .Z(
        n10319) );
  NAND2_X1 U12136 ( .A1(n10320), .A2(n10319), .ZN(n16344) );
  NAND2_X1 U12137 ( .A1(n14993), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n16343) );
  NAND2_X1 U12138 ( .A1(n16344), .A2(n16343), .ZN(n10323) );
  MUX2_X1 U12139 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10321), .S(n16341), .Z(
        n10322) );
  NAND2_X1 U12140 ( .A1(n10323), .A2(n10322), .ZN(n16346) );
  NAND2_X1 U12141 ( .A1(n16341), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10372) );
  NAND2_X1 U12142 ( .A1(n16346), .A2(n10372), .ZN(n10325) );
  MUX2_X1 U12143 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10865), .S(n10370), .Z(
        n10324) );
  NAND2_X1 U12144 ( .A1(n10325), .A2(n10324), .ZN(n10374) );
  NAND2_X1 U12145 ( .A1(n10370), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10329) );
  NAND2_X1 U12146 ( .A1(n10374), .A2(n10329), .ZN(n10327) );
  MUX2_X1 U12147 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11072), .S(n10351), .Z(
        n10326) );
  NAND2_X1 U12148 ( .A1(n10327), .A2(n10326), .ZN(n10348) );
  MUX2_X1 U12149 ( .A(n11072), .B(P1_REG2_REG_6__SCAN_IN), .S(n10351), .Z(
        n10328) );
  NAND3_X1 U12150 ( .A1(n10374), .A2(n10329), .A3(n10328), .ZN(n10330) );
  NAND3_X1 U12151 ( .A1(n16347), .A2(n10348), .A3(n10330), .ZN(n10331) );
  NAND2_X1 U12152 ( .A1(n10332), .A2(n10331), .ZN(P1_U3249) );
  INV_X1 U12153 ( .A(n11901), .ZN(n10342) );
  NOR2_X1 U12154 ( .A1(n10338), .A2(n10335), .ZN(n10334) );
  MUX2_X1 U12155 ( .A(n10335), .B(n10334), .S(P2_IR_REG_13__SCAN_IN), .Z(
        n10336) );
  INV_X1 U12156 ( .A(n10336), .ZN(n10339) );
  INV_X1 U12157 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n10337) );
  NAND2_X1 U12158 ( .A1(n10338), .A2(n10337), .ZN(n10468) );
  INV_X1 U12159 ( .A(n12275), .ZN(n11631) );
  OAI222_X1 U12160 ( .A1(n14818), .A2(n10340), .B1(n14816), .B2(n10342), .C1(
        n11631), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U12161 ( .A(n10675), .ZN(n10712) );
  OAI222_X1 U12162 ( .A1(P1_U3086), .A2(n10712), .B1(n15919), .B2(n10342), 
        .C1(n10341), .C2(n15916), .ZN(P1_U3342) );
  NAND2_X1 U12163 ( .A1(n10351), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10347) );
  NAND2_X1 U12164 ( .A1(n10348), .A2(n10347), .ZN(n10345) );
  INV_X1 U12165 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10343) );
  MUX2_X1 U12166 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10343), .S(n10384), .Z(
        n10344) );
  NAND2_X1 U12167 ( .A1(n10345), .A2(n10344), .ZN(n15010) );
  MUX2_X1 U12168 ( .A(n10343), .B(P1_REG2_REG_7__SCAN_IN), .S(n10384), .Z(
        n10346) );
  NAND3_X1 U12169 ( .A1(n10348), .A2(n10347), .A3(n10346), .ZN(n10349) );
  NAND3_X1 U12170 ( .A1(n16347), .A2(n15010), .A3(n10349), .ZN(n10358) );
  NAND2_X1 U12171 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11461) );
  MUX2_X1 U12172 ( .A(n9399), .B(P1_REG1_REG_7__SCAN_IN), .S(n10384), .Z(
        n10352) );
  NOR2_X1 U12173 ( .A1(n10353), .A2(n10352), .ZN(n10381) );
  AOI211_X1 U12174 ( .C1(n10353), .C2(n10352), .A(n10381), .B(n16266), .ZN(
        n10354) );
  INV_X1 U12175 ( .A(n10354), .ZN(n10355) );
  NAND2_X1 U12176 ( .A1(n11461), .A2(n10355), .ZN(n10356) );
  AOI21_X1 U12177 ( .B1(n14978), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n10356), .ZN(
        n10357) );
  OAI211_X1 U12178 ( .C1(n16358), .C2(n10359), .A(n10358), .B(n10357), .ZN(
        P1_U3250) );
  AOI22_X1 U12179 ( .A1(n13328), .A2(P3_STATE_REG_SCAN_IN), .B1(SI_17_), .B2(
        n10360), .ZN(n10361) );
  OAI21_X1 U12180 ( .B1(n10362), .B2(n13750), .A(n10361), .ZN(P3_U3278) );
  OAI21_X1 U12181 ( .B1(n10365), .B2(n10364), .A(n10363), .ZN(n10369) );
  INV_X1 U12182 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10367) );
  NAND2_X1 U12183 ( .A1(n15065), .A2(n10370), .ZN(n10366) );
  NAND2_X1 U12184 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n10914) );
  OAI211_X1 U12185 ( .C1(n10367), .C2(n16364), .A(n10366), .B(n10914), .ZN(
        n10368) );
  AOI21_X1 U12186 ( .B1(n16354), .B2(n10369), .A(n10368), .ZN(n10376) );
  MUX2_X1 U12187 ( .A(n10865), .B(P1_REG2_REG_5__SCAN_IN), .S(n10370), .Z(
        n10371) );
  NAND3_X1 U12188 ( .A1(n16346), .A2(n10372), .A3(n10371), .ZN(n10373) );
  NAND3_X1 U12189 ( .A1(n16347), .A2(n10374), .A3(n10373), .ZN(n10375) );
  NAND2_X1 U12190 ( .A1(n10376), .A2(n10375), .ZN(P1_U3248) );
  INV_X1 U12191 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n10380) );
  INV_X1 U12192 ( .A(n10378), .ZN(n10379) );
  AOI22_X1 U12193 ( .A1(n10377), .A2(n10380), .B1(n10379), .B2(n13737), .ZN(
        P3_U3376) );
  AOI21_X1 U12194 ( .B1(n10384), .B2(P1_REG1_REG_7__SCAN_IN), .A(n10381), .ZN(
        n15002) );
  INV_X1 U12195 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n16496) );
  MUX2_X1 U12196 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n16496), .S(n15007), .Z(
        n15001) );
  NOR2_X1 U12197 ( .A1(n15007), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n15016) );
  MUX2_X1 U12198 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9435), .S(n15024), .Z(
        n15017) );
  OAI21_X1 U12199 ( .B1(n15018), .B2(n15016), .A(n15017), .ZN(n15015) );
  OAI21_X1 U12200 ( .B1(n15024), .B2(P1_REG1_REG_9__SCAN_IN), .A(n15015), .ZN(
        n10383) );
  INV_X1 U12201 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n16525) );
  MUX2_X1 U12202 ( .A(n16525), .B(P1_REG1_REG_10__SCAN_IN), .S(n10425), .Z(
        n10382) );
  NOR2_X1 U12203 ( .A1(n10383), .A2(n10382), .ZN(n10420) );
  AOI211_X1 U12204 ( .C1(n10383), .C2(n10382), .A(n16266), .B(n10420), .ZN(
        n10400) );
  NAND2_X1 U12205 ( .A1(n10384), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n15009) );
  NAND2_X1 U12206 ( .A1(n15010), .A2(n15009), .ZN(n10387) );
  MUX2_X1 U12207 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10385), .S(n15007), .Z(
        n10386) );
  NAND2_X1 U12208 ( .A1(n10387), .A2(n10386), .ZN(n15027) );
  NAND2_X1 U12209 ( .A1(n15007), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n15026) );
  NAND2_X1 U12210 ( .A1(n15027), .A2(n15026), .ZN(n10390) );
  INV_X1 U12211 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10388) );
  MUX2_X1 U12212 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10388), .S(n15024), .Z(
        n10389) );
  NAND2_X1 U12213 ( .A1(n10390), .A2(n10389), .ZN(n15029) );
  NAND2_X1 U12214 ( .A1(n15024), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10394) );
  NAND2_X1 U12215 ( .A1(n15029), .A2(n10394), .ZN(n10392) );
  MUX2_X1 U12216 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11767), .S(n10425), .Z(
        n10391) );
  NAND2_X1 U12217 ( .A1(n10392), .A2(n10391), .ZN(n15042) );
  MUX2_X1 U12218 ( .A(n11767), .B(P1_REG2_REG_10__SCAN_IN), .S(n10425), .Z(
        n10393) );
  NAND3_X1 U12219 ( .A1(n15029), .A2(n10394), .A3(n10393), .ZN(n10395) );
  AND3_X1 U12220 ( .A1(n16347), .A2(n15042), .A3(n10395), .ZN(n10399) );
  NAND2_X1 U12221 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11971)
         );
  NAND2_X1 U12222 ( .A1(n14978), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n10396) );
  OAI211_X1 U12223 ( .C1(n16358), .C2(n10397), .A(n11971), .B(n10396), .ZN(
        n10398) );
  OR3_X1 U12224 ( .A1(n10400), .A2(n10399), .A3(n10398), .ZN(P1_U3253) );
  AND2_X1 U12225 ( .A1(n10377), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12226 ( .A1(n10377), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12227 ( .A1(n10377), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12228 ( .A1(n10377), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12229 ( .A1(n10377), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12230 ( .A1(n10377), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12231 ( .A1(n10377), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12232 ( .A1(n10377), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12233 ( .A1(n10377), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12234 ( .A1(n10377), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12235 ( .A1(n10377), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12236 ( .A1(n10377), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12237 ( .A1(n10377), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12238 ( .A1(n10377), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12239 ( .A1(n10377), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12240 ( .A1(n10377), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12241 ( .A1(n10377), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12242 ( .A1(n10377), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12243 ( .A1(n10377), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  INV_X1 U12244 ( .A(n12014), .ZN(n10404) );
  NAND2_X1 U12245 ( .A1(n10468), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10401) );
  INV_X1 U12246 ( .A(n12276), .ZN(n16188) );
  OAI222_X1 U12247 ( .A1(n14818), .A2(n10402), .B1(n14816), .B2(n10404), .C1(
        P2_U3088), .C2(n16188), .ZN(P2_U3313) );
  INV_X1 U12248 ( .A(n11378), .ZN(n10405) );
  OAI222_X1 U12249 ( .A1(n10405), .A2(P1_U3086), .B1(n15919), .B2(n10404), 
        .C1(n10403), .C2(n15916), .ZN(P1_U3341) );
  INV_X1 U12250 ( .A(n10473), .ZN(n10408) );
  NAND2_X1 U12251 ( .A1(n10495), .A2(n10408), .ZN(n10409) );
  INV_X1 U12252 ( .A(n16553), .ZN(n16551) );
  INV_X1 U12253 ( .A(n11129), .ZN(n10412) );
  NAND2_X1 U12254 ( .A1(n15361), .A2(n16449), .ZN(n10411) );
  AND2_X1 U12255 ( .A1(n10517), .A2(n15329), .ZN(n10410) );
  AOI21_X1 U12256 ( .B1(n10412), .B2(n10411), .A(n10410), .ZN(n11124) );
  INV_X1 U12257 ( .A(n10413), .ZN(n10414) );
  NAND2_X1 U12258 ( .A1(n10414), .A2(n11549), .ZN(n15475) );
  INV_X1 U12259 ( .A(n10491), .ZN(n10415) );
  OAI22_X1 U12260 ( .A1(n11129), .A2(n15475), .B1(n11207), .B2(n10415), .ZN(
        n10416) );
  INV_X1 U12261 ( .A(n10416), .ZN(n10417) );
  AND2_X1 U12262 ( .A1(n11124), .A2(n10417), .ZN(n16366) );
  NAND2_X1 U12263 ( .A1(n16551), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10418) );
  OAI21_X1 U12264 ( .B1(n16551), .B2(n16366), .A(n10418), .ZN(P1_U3528) );
  INV_X1 U12265 ( .A(n13353), .ZN(n13364) );
  OAI222_X1 U12266 ( .A1(P3_U3151), .A2(n13364), .B1(n13745), .B2(n15716), 
        .C1(n13750), .C2(n10419), .ZN(P3_U3277) );
  INV_X1 U12267 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n16552) );
  MUX2_X1 U12268 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n16552), .S(n15039), .Z(
        n15033) );
  AOI21_X1 U12269 ( .B1(n16552), .B2(n10421), .A(n15035), .ZN(n10423) );
  XNOR2_X1 U12270 ( .A(n10666), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n10422) );
  AOI21_X1 U12271 ( .B1(n10423), .B2(n10422), .A(n10671), .ZN(n10436) );
  INV_X1 U12272 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10424) );
  NAND2_X1 U12273 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n12177)
         );
  OAI21_X1 U12274 ( .B1(n16364), .B2(n10424), .A(n12177), .ZN(n10434) );
  NAND2_X1 U12275 ( .A1(n10425), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n15041) );
  NAND2_X1 U12276 ( .A1(n15042), .A2(n15041), .ZN(n10427) );
  MUX2_X1 U12277 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n11867), .S(n15039), .Z(
        n10426) );
  NAND2_X1 U12278 ( .A1(n10427), .A2(n10426), .ZN(n15044) );
  NAND2_X1 U12279 ( .A1(n15039), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10428) );
  NAND2_X1 U12280 ( .A1(n15044), .A2(n10428), .ZN(n10431) );
  MUX2_X1 U12281 ( .A(n10429), .B(P1_REG2_REG_12__SCAN_IN), .S(n10666), .Z(
        n10430) );
  OR2_X1 U12282 ( .A1(n10431), .A2(n10430), .ZN(n10668) );
  NAND2_X1 U12283 ( .A1(n10431), .A2(n10430), .ZN(n10432) );
  INV_X1 U12284 ( .A(n16347), .ZN(n16264) );
  AOI21_X1 U12285 ( .B1(n10668), .B2(n10432), .A(n16264), .ZN(n10433) );
  AOI211_X1 U12286 ( .C1(n15065), .C2(n10666), .A(n10434), .B(n10433), .ZN(
        n10435) );
  OAI21_X1 U12287 ( .B1(n10436), .B2(n16266), .A(n10435), .ZN(P1_U3255) );
  NAND2_X1 U12288 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14975) );
  INV_X1 U12289 ( .A(n10441), .ZN(n10443) );
  NAND2_X1 U12290 ( .A1(n10443), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10444) );
  NOR2_X1 U12291 ( .A1(n10445), .A2(n10486), .ZN(n10446) );
  NOR2_X1 U12292 ( .A1(n7488), .A2(n10446), .ZN(n11204) );
  MUX2_X1 U12293 ( .A(n14975), .B(n11204), .S(n15912), .Z(n10447) );
  INV_X1 U12294 ( .A(n10447), .ZN(n10451) );
  OAI21_X1 U12295 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n10448), .A(P1_U4016), .ZN(
        n10449) );
  AOI21_X1 U12296 ( .B1(n10451), .B2(n10450), .A(n10449), .ZN(n16360) );
  MUX2_X1 U12297 ( .A(n10303), .B(P1_REG1_REG_2__SCAN_IN), .S(n10461), .Z(
        n10453) );
  NAND3_X1 U12298 ( .A1(n10453), .A2(n14979), .A3(n10452), .ZN(n10454) );
  NAND2_X1 U12299 ( .A1(n10454), .A2(n14996), .ZN(n10464) );
  MUX2_X1 U12300 ( .A(n15340), .B(P1_REG2_REG_2__SCAN_IN), .S(n10461), .Z(
        n10456) );
  NAND3_X1 U12301 ( .A1(n10456), .A2(n14976), .A3(n10455), .ZN(n10457) );
  NAND3_X1 U12302 ( .A1(n16347), .A2(n14989), .A3(n10457), .ZN(n10463) );
  INV_X1 U12303 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10459) );
  OAI22_X1 U12304 ( .A1(n16364), .A2(n10459), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10458), .ZN(n10460) );
  AOI21_X1 U12305 ( .B1(n10461), .B2(n15065), .A(n10460), .ZN(n10462) );
  OAI211_X1 U12306 ( .C1(n16266), .C2(n10464), .A(n10463), .B(n10462), .ZN(
        n10465) );
  OR2_X1 U12307 ( .A1(n16360), .A2(n10465), .ZN(P1_U3245) );
  OAI222_X1 U12308 ( .A1(n13750), .A2(n10466), .B1(n13745), .B2(n15512), .C1(
        P3_U3151), .C2(n10592), .ZN(P3_U3276) );
  INV_X1 U12309 ( .A(n12090), .ZN(n10471) );
  INV_X1 U12310 ( .A(n11570), .ZN(n11382) );
  OAI222_X1 U12311 ( .A1(n15916), .A2(n10467), .B1(n15919), .B2(n10471), .C1(
        P1_U3086), .C2(n11382), .ZN(P1_U3340) );
  OAI21_X1 U12312 ( .B1(n10468), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n10470) );
  INV_X1 U12313 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n10469) );
  XNOR2_X1 U12314 ( .A(n10470), .B(n10469), .ZN(n14345) );
  OAI222_X1 U12315 ( .A1(n14818), .A2(n12091), .B1(n14816), .B2(n10471), .C1(
        n14345), .C2(P2_U3088), .ZN(P2_U3312) );
  INV_X1 U12316 ( .A(n10499), .ZN(n10472) );
  NAND2_X1 U12317 ( .A1(n10472), .A2(n10475), .ZN(n10477) );
  AOI21_X1 U12318 ( .B1(n10477), .B2(n10474), .A(n10473), .ZN(n10788) );
  NAND2_X1 U12319 ( .A1(n10788), .A2(n10495), .ZN(n11203) );
  INV_X1 U12320 ( .A(n11203), .ZN(n10504) );
  AND2_X1 U12321 ( .A1(n10476), .A2(n10475), .ZN(n10481) );
  INV_X1 U12322 ( .A(n10477), .ZN(n10479) );
  NAND3_X1 U12323 ( .A1(n10479), .A2(n10495), .A3(n10478), .ZN(n10480) );
  NAND2_X1 U12324 ( .A1(n10480), .A2(n15312), .ZN(n14844) );
  INV_X1 U12325 ( .A(n10481), .ZN(n14836) );
  INV_X1 U12326 ( .A(n9332), .ZN(n10482) );
  OAI22_X1 U12327 ( .A1(n14958), .A2(n16394), .B1(n14951), .B2(n10482), .ZN(
        n10483) );
  AOI21_X1 U12328 ( .B1(n14955), .B2(n14974), .A(n10483), .ZN(n10502) );
  OAI22_X1 U12329 ( .A1(n10651), .A2(n7468), .B1(n10644), .B2(n16394), .ZN(
        n10484) );
  XNOR2_X1 U12330 ( .A(n10484), .B(n12705), .ZN(n10648) );
  INV_X4 U12331 ( .A(n12377), .ZN(n12698) );
  NOR2_X1 U12332 ( .A1(n7468), .A2(n16394), .ZN(n10485) );
  AOI21_X1 U12333 ( .B1(n12698), .B2(n10517), .A(n10485), .ZN(n10646) );
  XNOR2_X1 U12334 ( .A(n10648), .B(n10646), .ZN(n10490) );
  INV_X1 U12335 ( .A(n10486), .ZN(n10487) );
  NOR2_X1 U12336 ( .A1(n7488), .A2(n10488), .ZN(n10489) );
  NAND2_X1 U12337 ( .A1(n10489), .A2(n10490), .ZN(n10647) );
  OAI21_X1 U12338 ( .B1(n10490), .B2(n10489), .A(n10647), .ZN(n10500) );
  NAND2_X1 U12339 ( .A1(n10491), .A2(n15185), .ZN(n10492) );
  NAND3_X1 U12340 ( .A1(n10495), .A2(n16542), .A3(n10494), .ZN(n10496) );
  OR2_X1 U12341 ( .A1(n10497), .A2(n10496), .ZN(n10498) );
  NAND2_X1 U12342 ( .A1(n10500), .A2(n14915), .ZN(n10501) );
  OAI211_X1 U12343 ( .C1(n10504), .C2(n10503), .A(n10502), .B(n10501), .ZN(
        P1_U3222) );
  NAND2_X1 U12344 ( .A1(n10506), .A2(n10505), .ZN(n10508) );
  NAND2_X1 U12345 ( .A1(n10509), .A2(n10637), .ZN(n10510) );
  NOR2_X4 U12346 ( .A1(n10639), .A2(n10510), .ZN(n16534) );
  NAND2_X1 U12347 ( .A1(n14296), .A2(n11958), .ZN(n14691) );
  OR2_X1 U12348 ( .A1(n14323), .A2(n13951), .ZN(n10511) );
  NAND2_X1 U12349 ( .A1(n11316), .A2(n10511), .ZN(n14246) );
  AND2_X1 U12350 ( .A1(n8139), .A2(n14591), .ZN(n10512) );
  OAI22_X1 U12351 ( .A1(n14246), .A2(n10512), .B1(n7948), .B2(n14374), .ZN(
        n10875) );
  AND2_X1 U12352 ( .A1(n13951), .A2(n10513), .ZN(n10514) );
  NOR2_X1 U12353 ( .A1(n10875), .A2(n10514), .ZN(n10876) );
  OAI21_X1 U12354 ( .B1(n14691), .B2(n14246), .A(n10876), .ZN(n11210) );
  NAND2_X1 U12355 ( .A1(n16534), .A2(n11210), .ZN(n10515) );
  OAI21_X1 U12356 ( .B1(n16534), .B2(n10034), .A(n10515), .ZN(P2_U3430) );
  OR2_X1 U12357 ( .A1(n10517), .A2(n10516), .ZN(n10518) );
  NAND2_X1 U12358 ( .A1(n10519), .A2(n10518), .ZN(n10521) );
  NAND2_X1 U12359 ( .A1(n10521), .A2(n10520), .ZN(n10848) );
  OAI21_X1 U12360 ( .B1(n10521), .B2(n10520), .A(n10848), .ZN(n15344) );
  INV_X1 U12361 ( .A(n15344), .ZN(n10532) );
  OAI21_X1 U12362 ( .B1(n10524), .B2(n10523), .A(n10856), .ZN(n10527) );
  INV_X1 U12363 ( .A(n14973), .ZN(n10849) );
  OAI22_X1 U12364 ( .A1(n10849), .A2(n15232), .B1(n10651), .B2(n15230), .ZN(
        n10526) );
  NOR2_X1 U12365 ( .A1(n10532), .A2(n15361), .ZN(n10525) );
  AOI211_X1 U12366 ( .C1(n15431), .C2(n10527), .A(n10526), .B(n10525), .ZN(
        n15339) );
  INV_X1 U12367 ( .A(n10528), .ZN(n10530) );
  NAND2_X1 U12368 ( .A1(n10528), .A2(n10642), .ZN(n11109) );
  INV_X1 U12369 ( .A(n11109), .ZN(n10529) );
  AOI21_X1 U12370 ( .B1(n15342), .B2(n10530), .A(n10529), .ZN(n15346) );
  AOI22_X1 U12371 ( .A1(n15346), .A2(n15471), .B1(n15342), .B2(n16445), .ZN(
        n10531) );
  OAI211_X1 U12372 ( .C1(n10532), .C2(n15475), .A(n15339), .B(n10531), .ZN(
        n10536) );
  NAND2_X1 U12373 ( .A1(n10536), .A2(n16553), .ZN(n10533) );
  OAI21_X1 U12374 ( .B1(n16553), .B2(n10303), .A(n10533), .ZN(P1_U3530) );
  INV_X1 U12375 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10538) );
  NAND2_X1 U12376 ( .A1(n10536), .A2(n16556), .ZN(n10537) );
  OAI21_X1 U12377 ( .B1(n16556), .B2(n10538), .A(n10537), .ZN(P1_U3465) );
  XNOR2_X1 U12378 ( .A(n10539), .B(n14250), .ZN(n11640) );
  INV_X1 U12379 ( .A(n14735), .ZN(n16583) );
  INV_X1 U12380 ( .A(n14709), .ZN(n16579) );
  AOI21_X1 U12381 ( .B1(n11332), .B2(n14019), .A(n7458), .ZN(n10541) );
  NAND2_X1 U12382 ( .A1(n10541), .A2(n10540), .ZN(n11638) );
  OAI21_X1 U12383 ( .B1(n10542), .B2(n16579), .A(n11638), .ZN(n10546) );
  XNOR2_X1 U12384 ( .A(n10543), .B(n14250), .ZN(n10545) );
  OAI21_X1 U12385 ( .B1(n10545), .B2(n14591), .A(n10544), .ZN(n11635) );
  AOI211_X1 U12386 ( .C1(n11640), .C2(n16583), .A(n10546), .B(n11635), .ZN(
        n10641) );
  OR2_X1 U12387 ( .A1(n10641), .A2(n16585), .ZN(n10547) );
  OAI21_X1 U12388 ( .B1(n16534), .B2(n10058), .A(n10547), .ZN(P2_U3439) );
  XNOR2_X1 U12389 ( .A(n14026), .B(n7463), .ZN(n11095) );
  NAND2_X1 U12390 ( .A1(n14318), .A2(n7458), .ZN(n10549) );
  XNOR2_X1 U12391 ( .A(n11095), .B(n10549), .ZN(n12771) );
  NAND3_X1 U12392 ( .A1(n12770), .A2(n12771), .A3(n10548), .ZN(n12780) );
  INV_X1 U12393 ( .A(n11095), .ZN(n10550) );
  NAND2_X1 U12394 ( .A1(n10550), .A2(n10549), .ZN(n10551) );
  NAND2_X1 U12395 ( .A1(n12780), .A2(n10551), .ZN(n10555) );
  NAND2_X1 U12396 ( .A1(n10552), .A2(n11900), .ZN(n10554) );
  INV_X1 U12397 ( .A(n16141), .ZN(n11187) );
  AOI22_X1 U12398 ( .A1(n10051), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n10048), 
        .B2(n11187), .ZN(n10553) );
  NAND2_X1 U12399 ( .A1(n10554), .A2(n10553), .ZN(n14032) );
  XNOR2_X1 U12400 ( .A(n14032), .B(n7463), .ZN(n10556) );
  NAND2_X1 U12401 ( .A1(n14317), .A2(n7458), .ZN(n10557) );
  XNOR2_X1 U12402 ( .A(n10556), .B(n10557), .ZN(n11096) );
  NAND2_X1 U12403 ( .A1(n10555), .A2(n11096), .ZN(n11102) );
  INV_X1 U12404 ( .A(n10556), .ZN(n10558) );
  NAND2_X1 U12405 ( .A1(n10558), .A2(n10557), .ZN(n10559) );
  AND2_X1 U12406 ( .A1(n11102), .A2(n10559), .ZN(n10577) );
  NAND2_X1 U12407 ( .A1(n10560), .A2(n11900), .ZN(n10562) );
  AOI22_X1 U12408 ( .A1(n10051), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n10048), 
        .B2(n16156), .ZN(n10561) );
  NAND2_X1 U12409 ( .A1(n10562), .A2(n10561), .ZN(n14038) );
  XNOR2_X1 U12410 ( .A(n14038), .B(n7463), .ZN(n10572) );
  NAND2_X1 U12411 ( .A1(n13902), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10571) );
  INV_X1 U12412 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10563) );
  OR2_X1 U12413 ( .A1(n10986), .A2(n10563), .ZN(n10570) );
  INV_X1 U12414 ( .A(n10566), .ZN(n10564) );
  NAND2_X1 U12415 ( .A1(n10564), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10579) );
  INV_X1 U12416 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10565) );
  NAND2_X1 U12417 ( .A1(n10566), .A2(n10565), .ZN(n10567) );
  NAND2_X1 U12418 ( .A1(n10579), .A2(n10567), .ZN(n11370) );
  OR2_X1 U12419 ( .A1(n10059), .A2(n11370), .ZN(n10569) );
  INV_X1 U12420 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11369) );
  OR2_X1 U12421 ( .A1(n14192), .A2(n11369), .ZN(n10568) );
  NAND4_X1 U12422 ( .A1(n10571), .A2(n10570), .A3(n10569), .A4(n10568), .ZN(
        n14316) );
  AND2_X1 U12423 ( .A1(n14316), .A2(n7458), .ZN(n10573) );
  NAND2_X1 U12424 ( .A1(n10572), .A2(n10573), .ZN(n10726) );
  INV_X1 U12425 ( .A(n10572), .ZN(n12758) );
  INV_X1 U12426 ( .A(n10573), .ZN(n10574) );
  NAND2_X1 U12427 ( .A1(n12758), .A2(n10574), .ZN(n10575) );
  AND2_X1 U12428 ( .A1(n10726), .A2(n10575), .ZN(n10576) );
  NAND2_X1 U12429 ( .A1(n10577), .A2(n10576), .ZN(n12757) );
  OAI211_X1 U12430 ( .C1(n10577), .C2(n10576), .A(n12757), .B(n13977), .ZN(
        n10590) );
  INV_X1 U12431 ( .A(n13975), .ZN(n13945) );
  NAND2_X1 U12432 ( .A1(n14317), .A2(n14613), .ZN(n10586) );
  NAND2_X1 U12433 ( .A1(n14181), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n10584) );
  INV_X1 U12434 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11174) );
  OR2_X1 U12435 ( .A1(n14192), .A2(n11174), .ZN(n10583) );
  NAND2_X1 U12436 ( .A1(n10579), .A2(n10578), .ZN(n10580) );
  NAND2_X1 U12437 ( .A1(n10734), .A2(n10580), .ZN(n11489) );
  OR2_X1 U12438 ( .A1(n10059), .A2(n11489), .ZN(n10582) );
  INV_X1 U12439 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n11189) );
  OR2_X1 U12440 ( .A1(n14191), .A2(n11189), .ZN(n10581) );
  NAND4_X1 U12441 ( .A1(n10584), .A2(n10583), .A3(n10582), .A4(n10581), .ZN(
        n14315) );
  NAND2_X1 U12442 ( .A1(n14315), .A2(n14614), .ZN(n10585) );
  NAND2_X1 U12443 ( .A1(n10586), .A2(n10585), .ZN(n10806) );
  AOI22_X1 U12444 ( .A1(n13945), .A2(n10806), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10587) );
  OAI21_X1 U12445 ( .B1(n11370), .B2(n13943), .A(n10587), .ZN(n10588) );
  AOI21_X1 U12446 ( .B1(n14038), .B2(n13952), .A(n10588), .ZN(n10589) );
  NAND2_X1 U12447 ( .A1(n10590), .A2(n10589), .ZN(P2_U3211) );
  NOR2_X1 U12448 ( .A1(n10593), .A2(n10592), .ZN(n10595) );
  INV_X1 U12449 ( .A(n13056), .ZN(n10594) );
  INV_X1 U12450 ( .A(n16367), .ZN(n10598) );
  NAND2_X1 U12451 ( .A1(n10605), .A2(n16558), .ZN(n10602) );
  OAI22_X1 U12452 ( .A1(n10620), .A2(n10602), .B1(n10616), .B2(n10606), .ZN(
        n10604) );
  NAND2_X1 U12453 ( .A1(n10620), .A2(n10605), .ZN(n10610) );
  INV_X1 U12454 ( .A(n10606), .ZN(n10607) );
  NAND2_X1 U12455 ( .A1(n10616), .A2(n10607), .ZN(n10608) );
  NAND4_X1 U12456 ( .A1(n10610), .A2(n10609), .A3(n10608), .A4(n10684), .ZN(
        n10611) );
  NAND2_X1 U12457 ( .A1(n10611), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10613) );
  NOR2_X1 U12458 ( .A1(n10924), .A2(n10692), .ZN(n13062) );
  NAND2_X1 U12459 ( .A1(n10616), .A2(n13062), .ZN(n10612) );
  NAND2_X1 U12460 ( .A1(n10613), .A2(n10612), .ZN(n11086) );
  OR2_X1 U12461 ( .A1(n11086), .A2(n10614), .ZN(n10720) );
  INV_X1 U12462 ( .A(n13062), .ZN(n10615) );
  NOR2_X1 U12463 ( .A1(n10616), .A2(n10615), .ZN(n10619) );
  INV_X1 U12464 ( .A(n10617), .ZN(n10618) );
  INV_X1 U12465 ( .A(n16375), .ZN(n13228) );
  OR3_X1 U12466 ( .A1(n10620), .A2(n10924), .A3(n16558), .ZN(n10622) );
  NAND2_X1 U12467 ( .A1(n16471), .A2(n13060), .ZN(n10621) );
  AOI22_X1 U12468 ( .A1(n13185), .A2(n13228), .B1(n10623), .B2(n13168), .ZN(
        n10624) );
  OAI21_X1 U12469 ( .B1(n16373), .B2(n13187), .A(n10624), .ZN(n10625) );
  AOI21_X1 U12470 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(n10720), .A(n10625), .ZN(
        n10626) );
  OAI21_X1 U12471 ( .B1(n10627), .B2(n13204), .A(n10626), .ZN(P3_U3162) );
  INV_X1 U12472 ( .A(n12211), .ZN(n10633) );
  NAND2_X1 U12473 ( .A1(n10628), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10629) );
  XNOR2_X1 U12474 ( .A(n10629), .B(P2_IR_REG_16__SCAN_IN), .ZN(n16207) );
  INV_X1 U12475 ( .A(n16207), .ZN(n10630) );
  OAI222_X1 U12476 ( .A1(n14818), .A2(n10631), .B1(n14816), .B2(n10633), .C1(
        n10630), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U12477 ( .A(n11705), .ZN(n11588) );
  OAI222_X1 U12478 ( .A1(P1_U3086), .A2(n11588), .B1(n15919), .B2(n10633), 
        .C1(n10632), .C2(n15916), .ZN(P1_U3339) );
  AND2_X1 U12479 ( .A1(n13228), .A2(n10846), .ZN(n12856) );
  INV_X1 U12480 ( .A(n12856), .ZN(n12854) );
  AND2_X1 U12481 ( .A1(n16367), .A2(n12854), .ZN(n13013) );
  AOI22_X1 U12482 ( .A1(n13196), .A2(n13227), .B1(n10691), .B2(n13168), .ZN(
        n10635) );
  NAND2_X1 U12483 ( .A1(n10720), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10634) );
  OAI211_X1 U12484 ( .C1(n13013), .C2(n13204), .A(n10635), .B(n10634), .ZN(
        P3_U3172) );
  OR2_X1 U12485 ( .A1(n10637), .A2(n10636), .ZN(n10638) );
  NOR2_X4 U12486 ( .A1(n10639), .A2(n10638), .ZN(n14740) );
  INV_X1 U12487 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n11183) );
  NAND2_X1 U12488 ( .A1(n16584), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10640) );
  OAI21_X1 U12489 ( .B1(n10641), .B2(n16584), .A(n10640), .ZN(P2_U3502) );
  INV_X1 U12490 ( .A(n14915), .ZN(n11466) );
  NOR2_X1 U12491 ( .A1(n7468), .A2(n10642), .ZN(n10643) );
  AOI21_X1 U12492 ( .B1(n12698), .B2(n9332), .A(n10643), .ZN(n10774) );
  AOI22_X1 U12493 ( .A1(n7456), .A2(n9332), .B1(n12687), .B2(n15342), .ZN(
        n10645) );
  XNOR2_X1 U12494 ( .A(n10645), .B(n12705), .ZN(n10775) );
  XOR2_X1 U12495 ( .A(n10774), .B(n10775), .Z(n10776) );
  INV_X1 U12496 ( .A(n10646), .ZN(n10649) );
  OAI21_X1 U12497 ( .B1(n10649), .B2(n10648), .A(n10647), .ZN(n10777) );
  XOR2_X1 U12498 ( .A(n10776), .B(n10777), .Z(n10654) );
  INV_X1 U12499 ( .A(n14955), .ZN(n14861) );
  INV_X1 U12500 ( .A(n14951), .ZN(n14845) );
  AOI22_X1 U12501 ( .A1(n14845), .A2(n14973), .B1(n15342), .B2(n14844), .ZN(
        n10650) );
  OAI21_X1 U12502 ( .B1(n10651), .B2(n14861), .A(n10650), .ZN(n10652) );
  AOI21_X1 U12503 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n11203), .A(n10652), .ZN(
        n10653) );
  OAI21_X1 U12504 ( .B1(n11466), .B2(n10654), .A(n10653), .ZN(P1_U3237) );
  OAI222_X1 U12505 ( .A1(n13750), .A2(n10657), .B1(n13745), .B2(n10656), .C1(
        P3_U3151), .C2(n10655), .ZN(P3_U3275) );
  NAND2_X1 U12506 ( .A1(n13977), .A2(n7458), .ZN(n13967) );
  INV_X1 U12507 ( .A(n10658), .ZN(n10659) );
  OAI22_X1 U12508 ( .A1(n13967), .A2(n11316), .B1(n10659), .B2(n13915), .ZN(
        n10663) );
  NOR2_X1 U12509 ( .A1(n10660), .A2(P2_U3088), .ZN(n13948) );
  AOI22_X1 U12510 ( .A1(n14614), .A2(n14320), .B1(n14323), .B2(n14613), .ZN(
        n11323) );
  OAI22_X1 U12511 ( .A1(n13948), .A2(n11444), .B1(n13975), .B2(n11323), .ZN(
        n10662) );
  NOR2_X1 U12512 ( .A1(n13966), .A2(n13995), .ZN(n10661) );
  AOI211_X1 U12513 ( .C1(n10664), .C2(n10663), .A(n10662), .B(n10661), .ZN(
        n10665) );
  OAI21_X1 U12514 ( .B1(n10765), .B2(n13915), .A(n10665), .ZN(P2_U3194) );
  OR2_X1 U12515 ( .A1(n10666), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10667) );
  NAND2_X1 U12516 ( .A1(n10668), .A2(n10667), .ZN(n10702) );
  INV_X1 U12517 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10669) );
  MUX2_X1 U12518 ( .A(n10669), .B(P1_REG2_REG_13__SCAN_IN), .S(n10675), .Z(
        n10701) );
  NAND2_X1 U12519 ( .A1(n10675), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10670) );
  NAND2_X1 U12520 ( .A1(n10703), .A2(n10670), .ZN(n11381) );
  XNOR2_X1 U12521 ( .A(n11378), .B(n12341), .ZN(n11380) );
  XNOR2_X1 U12522 ( .A(n11381), .B(n11380), .ZN(n10683) );
  AOI21_X1 U12523 ( .B1(n10673), .B2(n10672), .A(n10671), .ZN(n10706) );
  XOR2_X1 U12524 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10675), .Z(n10707) );
  XNOR2_X1 U12525 ( .A(n11378), .B(n10674), .ZN(n10676) );
  NAND2_X1 U12526 ( .A1(n10675), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n10677) );
  NAND3_X1 U12527 ( .A1(n10705), .A2(n10676), .A3(n10677), .ZN(n11376) );
  INV_X1 U12528 ( .A(n11376), .ZN(n10679) );
  AOI21_X1 U12529 ( .B1(n10705), .B2(n10677), .A(n10676), .ZN(n10678) );
  OAI21_X1 U12530 ( .B1(n10679), .B2(n10678), .A(n16354), .ZN(n10682) );
  INV_X1 U12531 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n15956) );
  NAND2_X1 U12532 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n12386)
         );
  OAI21_X1 U12533 ( .B1(n16364), .B2(n15956), .A(n12386), .ZN(n10680) );
  AOI21_X1 U12534 ( .B1(n11378), .B2(n15065), .A(n10680), .ZN(n10681) );
  OAI211_X1 U12535 ( .C1(n10683), .C2(n16264), .A(n10682), .B(n10681), .ZN(
        P1_U3257) );
  INV_X1 U12536 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10939) );
  INV_X1 U12537 ( .A(n10684), .ZN(n10685) );
  NOR2_X1 U12538 ( .A1(n13738), .A2(n10685), .ZN(n10687) );
  MUX2_X1 U12539 ( .A(n13738), .B(n10687), .S(n10686), .Z(n10688) );
  OR2_X1 U12540 ( .A1(n16558), .A2(n13060), .ZN(n16400) );
  AOI22_X1 U12541 ( .A1(n13555), .A2(n10691), .B1(n16388), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10695) );
  NAND2_X1 U12542 ( .A1(n10692), .A2(n16558), .ZN(n10693) );
  OAI22_X1 U12543 ( .A1(n13013), .A2(n10693), .B1(n8573), .B2(n16372), .ZN(
        n10844) );
  NAND2_X1 U12544 ( .A1(n16411), .A2(n10844), .ZN(n10694) );
  OAI211_X1 U12545 ( .C1(n10939), .C2(n16411), .A(n10695), .B(n10694), .ZN(
        P3_U3233) );
  INV_X1 U12546 ( .A(n12354), .ZN(n10699) );
  NAND2_X1 U12547 ( .A1(n10696), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n11391) );
  XNOR2_X1 U12548 ( .A(n11391), .B(P2_IR_REG_17__SCAN_IN), .ZN(n16218) );
  INV_X1 U12549 ( .A(n16218), .ZN(n10697) );
  OAI222_X1 U12550 ( .A1(n14818), .A2(n10698), .B1(n14816), .B2(n10699), .C1(
        P2_U3088), .C2(n10697), .ZN(P2_U3310) );
  INV_X1 U12551 ( .A(n11708), .ZN(n15055) );
  OAI222_X1 U12552 ( .A1(n15916), .A2(n10700), .B1(n15919), .B2(n10699), .C1(
        n15055), .C2(P1_U3086), .ZN(P1_U3338) );
  AOI21_X1 U12553 ( .B1(n10702), .B2(n10701), .A(n16264), .ZN(n10704) );
  NAND2_X1 U12554 ( .A1(n10704), .A2(n10703), .ZN(n10711) );
  NAND2_X1 U12555 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n12263)
         );
  OAI211_X1 U12556 ( .C1(n10707), .C2(n10706), .A(n16354), .B(n10705), .ZN(
        n10708) );
  NAND2_X1 U12557 ( .A1(n12263), .A2(n10708), .ZN(n10709) );
  AOI21_X1 U12558 ( .B1(n14978), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10709), 
        .ZN(n10710) );
  OAI211_X1 U12559 ( .C1(n16358), .C2(n10712), .A(n10711), .B(n10710), .ZN(
        P1_U3256) );
  XNOR2_X1 U12560 ( .A(n12834), .B(n16402), .ZN(n11079) );
  XNOR2_X1 U12561 ( .A(n11079), .B(n13226), .ZN(n10717) );
  INV_X1 U12562 ( .A(n10713), .ZN(n10714) );
  AOI21_X1 U12563 ( .B1(n10717), .B2(n10716), .A(n11080), .ZN(n10722) );
  AOI22_X1 U12564 ( .A1(n13185), .A2(n13227), .B1(n16402), .B2(n13168), .ZN(
        n10718) );
  OAI21_X1 U12565 ( .B1(n11590), .B2(n13187), .A(n10718), .ZN(n10719) );
  AOI21_X1 U12566 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10720), .A(n10719), .ZN(
        n10721) );
  OAI21_X1 U12567 ( .B1(n10722), .B2(n13204), .A(n10721), .ZN(P3_U3177) );
  NAND2_X1 U12568 ( .A1(n10723), .A2(n11900), .ZN(n10725) );
  AOI22_X1 U12569 ( .A1(n10051), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n10048), 
        .B2(n14331), .ZN(n10724) );
  XNOR2_X1 U12570 ( .A(n14044), .B(n7463), .ZN(n10727) );
  NAND2_X1 U12571 ( .A1(n14315), .A2(n7458), .ZN(n10728) );
  XNOR2_X1 U12572 ( .A(n10727), .B(n10728), .ZN(n12762) );
  INV_X1 U12573 ( .A(n10727), .ZN(n10741) );
  NAND2_X1 U12574 ( .A1(n10741), .A2(n10728), .ZN(n10729) );
  NAND2_X1 U12575 ( .A1(n10730), .A2(n11900), .ZN(n10732) );
  AOI22_X1 U12576 ( .A1(n10051), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n16169), 
        .B2(n10048), .ZN(n10731) );
  NAND2_X1 U12577 ( .A1(n10732), .A2(n10731), .ZN(n14052) );
  XNOR2_X1 U12578 ( .A(n14052), .B(n7463), .ZN(n10981) );
  NAND2_X1 U12579 ( .A1(n13902), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10739) );
  INV_X1 U12580 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10733) );
  OR2_X1 U12581 ( .A1(n10986), .A2(n10733), .ZN(n10738) );
  NAND2_X1 U12582 ( .A1(n10734), .A2(n10751), .ZN(n10735) );
  NAND2_X1 U12583 ( .A1(n10743), .A2(n10735), .ZN(n10754) );
  OR2_X1 U12584 ( .A1(n10059), .A2(n10754), .ZN(n10737) );
  INV_X1 U12585 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n11177) );
  OR2_X1 U12586 ( .A1(n14192), .A2(n11177), .ZN(n10736) );
  NAND4_X1 U12587 ( .A1(n10739), .A2(n10738), .A3(n10737), .A4(n10736), .ZN(
        n14314) );
  NAND2_X1 U12588 ( .A1(n14314), .A2(n7458), .ZN(n10976) );
  XNOR2_X1 U12589 ( .A(n10981), .B(n10976), .ZN(n10740) );
  INV_X1 U12590 ( .A(n14315), .ZN(n14046) );
  OAI22_X1 U12591 ( .A1(n13967), .A2(n14046), .B1(n10741), .B2(n13915), .ZN(
        n10742) );
  NAND3_X1 U12592 ( .A1(n12767), .A2(n7908), .A3(n10742), .ZN(n10758) );
  NAND2_X1 U12593 ( .A1(n14315), .A2(n14613), .ZN(n10750) );
  NAND2_X1 U12594 ( .A1(n14181), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n10748) );
  INV_X1 U12595 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11191) );
  OR2_X1 U12596 ( .A1(n14191), .A2(n11191), .ZN(n10747) );
  NAND2_X1 U12597 ( .A1(n10743), .A2(n10997), .ZN(n10744) );
  NAND2_X1 U12598 ( .A1(n10989), .A2(n10744), .ZN(n11000) );
  OR2_X1 U12599 ( .A1(n10059), .A2(n11000), .ZN(n10746) );
  INV_X1 U12600 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11178) );
  OR2_X1 U12601 ( .A1(n14192), .A2(n11178), .ZN(n10745) );
  NAND4_X1 U12602 ( .A1(n10748), .A2(n10747), .A3(n10746), .A4(n10745), .ZN(
        n14313) );
  NAND2_X1 U12603 ( .A1(n14313), .A2(n14614), .ZN(n10749) );
  NAND2_X1 U12604 ( .A1(n10750), .A2(n10749), .ZN(n11060) );
  INV_X1 U12605 ( .A(n11060), .ZN(n10752) );
  OAI22_X1 U12606 ( .A1(n13975), .A2(n10752), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10751), .ZN(n10753) );
  INV_X1 U12607 ( .A(n10753), .ZN(n10757) );
  NAND2_X1 U12608 ( .A1(n13952), .A2(n14052), .ZN(n10756) );
  INV_X1 U12609 ( .A(n10754), .ZN(n11550) );
  NAND2_X1 U12610 ( .A1(n13972), .A2(n11550), .ZN(n10755) );
  AND4_X1 U12611 ( .A1(n10758), .A2(n10757), .A3(n10756), .A4(n10755), .ZN(
        n10759) );
  OAI21_X1 U12612 ( .B1(n10984), .B2(n13915), .A(n10759), .ZN(P2_U3193) );
  OR2_X1 U12613 ( .A1(n13975), .A2(n13941), .ZN(n13932) );
  INV_X1 U12614 ( .A(n13932), .ZN(n13888) );
  OR2_X1 U12615 ( .A1(n13975), .A2(n14374), .ZN(n13933) );
  NOR2_X1 U12616 ( .A1(n13933), .A2(n10760), .ZN(n10762) );
  OAI22_X1 U12617 ( .A1(n13966), .A2(n16418), .B1(n13948), .B2(n11334), .ZN(
        n10761) );
  AOI211_X1 U12618 ( .C1(n13888), .C2(n14321), .A(n10762), .B(n10761), .ZN(
        n10769) );
  OAI22_X1 U12619 ( .A1(n13967), .A2(n7948), .B1(n10763), .B2(n13915), .ZN(
        n10767) );
  INV_X1 U12620 ( .A(n10764), .ZN(n10766) );
  NAND3_X1 U12621 ( .A1(n10767), .A2(n10766), .A3(n10765), .ZN(n10768) );
  OAI211_X1 U12622 ( .C1(n13915), .C2(n10770), .A(n10769), .B(n10768), .ZN(
        P2_U3209) );
  NOR2_X1 U12623 ( .A1(n16565), .A2(n10929), .ZN(n10771) );
  AOI21_X1 U12624 ( .B1(n16565), .B2(n10844), .A(n10771), .ZN(n10772) );
  OAI21_X1 U12625 ( .B1(n10846), .B2(n13657), .A(n10772), .ZN(P3_U3459) );
  AOI22_X1 U12626 ( .A1(n12698), .A2(n14973), .B1(n7456), .B2(n14843), .ZN(
        n10780) );
  OAI22_X1 U12627 ( .A1(n10849), .A2(n7468), .B1(n10644), .B2(n16429), .ZN(
        n10773) );
  XNOR2_X1 U12628 ( .A(n10773), .B(n12705), .ZN(n10778) );
  INV_X1 U12629 ( .A(n10778), .ZN(n10779) );
  XNOR2_X1 U12630 ( .A(n10780), .B(n10778), .ZN(n14841) );
  NAND2_X1 U12631 ( .A1(n14842), .A2(n14841), .ZN(n14840) );
  OAI21_X1 U12632 ( .B1(n10780), .B2(n10779), .A(n14840), .ZN(n10783) );
  AOI21_X1 U12633 ( .B1(n7456), .B2(n16446), .A(n12698), .ZN(n10781) );
  AOI21_X1 U12634 ( .B1(n10915), .B2(n7468), .A(n10781), .ZN(n10782) );
  NAND2_X1 U12635 ( .A1(n8111), .A2(n10905), .ZN(n10785) );
  OAI22_X1 U12636 ( .A1(n10851), .A2(n10644), .B1(n7468), .B2(n10915), .ZN(
        n10784) );
  XOR2_X1 U12637 ( .A(n12705), .B(n10784), .Z(n10906) );
  XNOR2_X1 U12638 ( .A(n10785), .B(n10906), .ZN(n10793) );
  NAND2_X1 U12639 ( .A1(n14973), .A2(n15331), .ZN(n10787) );
  NAND2_X1 U12640 ( .A1(n14971), .A2(n15329), .ZN(n10786) );
  AND2_X1 U12641 ( .A1(n10787), .A2(n10786), .ZN(n11158) );
  NAND2_X1 U12642 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n16361) );
  OAI21_X1 U12643 ( .B1(n14836), .B2(n11158), .A(n16361), .ZN(n10791) );
  AOI21_X1 U12644 ( .B1(n10788), .B2(n10441), .A(P1_U3086), .ZN(n10789) );
  NOR2_X2 U12645 ( .A1(n10789), .A2(n12047), .ZN(n14952) );
  NOR2_X1 U12646 ( .A1(n14952), .A2(n11160), .ZN(n10790) );
  AOI211_X1 U12647 ( .C1(n16446), .C2(n14844), .A(n10791), .B(n10790), .ZN(
        n10792) );
  OAI21_X1 U12648 ( .B1(n10793), .B2(n11466), .A(n10792), .ZN(P1_U3230) );
  INV_X1 U12649 ( .A(n14252), .ZN(n10794) );
  NAND2_X1 U12650 ( .A1(n10795), .A2(n10794), .ZN(n10797) );
  OR2_X1 U12651 ( .A1(n14026), .A2(n14318), .ZN(n10796) );
  XNOR2_X1 U12652 ( .A(n14032), .B(n14317), .ZN(n14253) );
  INV_X1 U12653 ( .A(n14253), .ZN(n10798) );
  OR2_X1 U12654 ( .A1(n14032), .A2(n14317), .ZN(n10799) );
  XNOR2_X1 U12655 ( .A(n14038), .B(n14316), .ZN(n14255) );
  XNOR2_X1 U12656 ( .A(n10817), .B(n14255), .ZN(n11375) );
  INV_X1 U12657 ( .A(n14318), .ZN(n14028) );
  NAND2_X1 U12658 ( .A1(n14026), .A2(n14028), .ZN(n10800) );
  OR2_X1 U12659 ( .A1(n14032), .A2(n10803), .ZN(n10802) );
  NAND2_X1 U12660 ( .A1(n10833), .A2(n10802), .ZN(n10805) );
  NAND2_X1 U12661 ( .A1(n14032), .A2(n10803), .ZN(n10804) );
  NAND2_X1 U12662 ( .A1(n10805), .A2(n10804), .ZN(n10820) );
  XNOR2_X1 U12663 ( .A(n10820), .B(n14255), .ZN(n10807) );
  AOI21_X1 U12664 ( .B1(n10807), .B2(n7449), .A(n10806), .ZN(n11368) );
  INV_X1 U12665 ( .A(n14032), .ZN(n11481) );
  NAND2_X1 U12666 ( .A1(n11481), .A2(n10837), .ZN(n10838) );
  INV_X1 U12667 ( .A(n10828), .ZN(n10808) );
  AOI211_X1 U12668 ( .C1(n14038), .C2(n10838), .A(n7458), .B(n10808), .ZN(
        n11372) );
  AOI21_X1 U12669 ( .B1(n14709), .B2(n14038), .A(n11372), .ZN(n10809) );
  OAI211_X1 U12670 ( .C1(n14735), .C2(n11375), .A(n11368), .B(n10809), .ZN(
        n14744) );
  NAND2_X1 U12671 ( .A1(n14744), .A2(n12115), .ZN(n10810) );
  OAI21_X1 U12672 ( .B1(n16534), .B2(n10563), .A(n10810), .ZN(P2_U3448) );
  AOI21_X1 U12673 ( .B1(n14709), .B2(n14026), .A(n10811), .ZN(n10812) );
  OAI211_X1 U12674 ( .C1(n14735), .C2(n10814), .A(n10813), .B(n10812), .ZN(
        n14745) );
  NAND2_X1 U12675 ( .A1(n14745), .A2(n12115), .ZN(n10815) );
  OAI21_X1 U12676 ( .B1(n16534), .B2(n10071), .A(n10815), .ZN(P2_U3442) );
  INV_X1 U12677 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10831) );
  XNOR2_X1 U12678 ( .A(n14044), .B(n14046), .ZN(n14257) );
  INV_X1 U12679 ( .A(n14255), .ZN(n10816) );
  OR2_X1 U12680 ( .A1(n14038), .A2(n14316), .ZN(n10818) );
  NAND2_X1 U12681 ( .A1(n10819), .A2(n10818), .ZN(n11053) );
  XOR2_X1 U12682 ( .A(n11053), .B(n14257), .Z(n11497) );
  INV_X1 U12683 ( .A(n14316), .ZN(n12759) );
  NAND2_X1 U12684 ( .A1(n14038), .A2(n12759), .ZN(n10821) );
  AOI21_X1 U12685 ( .B1(n10823), .B2(n14257), .A(n14591), .ZN(n10827) );
  NAND2_X1 U12686 ( .A1(n14316), .A2(n14613), .ZN(n10825) );
  NAND2_X1 U12687 ( .A1(n14314), .A2(n14614), .ZN(n10824) );
  AND2_X1 U12688 ( .A1(n10825), .A2(n10824), .ZN(n12756) );
  INV_X1 U12689 ( .A(n12756), .ZN(n10826) );
  AOI21_X1 U12690 ( .B1(n10827), .B2(n11059), .A(n10826), .ZN(n11492) );
  AOI211_X1 U12691 ( .C1(n14044), .C2(n10828), .A(n7458), .B(n11062), .ZN(
        n11495) );
  AOI21_X1 U12692 ( .B1(n14709), .B2(n14044), .A(n11495), .ZN(n10829) );
  OAI211_X1 U12693 ( .C1(n11497), .C2(n14735), .A(n11492), .B(n10829), .ZN(
        n11229) );
  NAND2_X1 U12694 ( .A1(n11229), .A2(n12115), .ZN(n10830) );
  OAI21_X1 U12695 ( .B1(n16534), .B2(n10831), .A(n10830), .ZN(P2_U3451) );
  XNOR2_X1 U12696 ( .A(n10832), .B(n14253), .ZN(n11485) );
  XNOR2_X1 U12697 ( .A(n10833), .B(n14253), .ZN(n10836) );
  NAND2_X1 U12698 ( .A1(n14318), .A2(n14613), .ZN(n10835) );
  NAND2_X1 U12699 ( .A1(n14316), .A2(n14614), .ZN(n10834) );
  NAND2_X1 U12700 ( .A1(n10835), .A2(n10834), .ZN(n11091) );
  AOI21_X1 U12701 ( .B1(n10836), .B2(n7449), .A(n11091), .ZN(n11488) );
  INV_X1 U12702 ( .A(n10837), .ZN(n10839) );
  AOI211_X1 U12703 ( .C1(n14032), .C2(n10839), .A(n7458), .B(n7692), .ZN(
        n11484) );
  AOI21_X1 U12704 ( .B1(n14709), .B2(n14032), .A(n11484), .ZN(n10840) );
  OAI211_X1 U12705 ( .C1(n14735), .C2(n11485), .A(n11488), .B(n10840), .ZN(
        n11231) );
  NAND2_X1 U12706 ( .A1(n11231), .A2(n12115), .ZN(n10841) );
  OAI21_X1 U12707 ( .B1(n16534), .B2(n10091), .A(n10841), .ZN(P2_U3445) );
  INV_X1 U12708 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10842) );
  NOR2_X1 U12709 ( .A1(n16569), .A2(n10842), .ZN(n10843) );
  AOI21_X1 U12710 ( .B1(n16569), .B2(n10844), .A(n10843), .ZN(n10845) );
  OAI21_X1 U12711 ( .B1(n10846), .B2(n13731), .A(n10845), .ZN(P3_U3390) );
  NAND2_X1 U12712 ( .A1(n10848), .A2(n10847), .ZN(n11106) );
  INV_X1 U12713 ( .A(n11113), .ZN(n11105) );
  NAND2_X1 U12714 ( .A1(n11106), .A2(n11105), .ZN(n11108) );
  NAND2_X1 U12715 ( .A1(n10849), .A2(n16429), .ZN(n10850) );
  NAND2_X1 U12716 ( .A1(n11108), .A2(n10850), .ZN(n11167) );
  NAND2_X1 U12717 ( .A1(n11167), .A2(n11166), .ZN(n11165) );
  NAND2_X1 U12718 ( .A1(n10851), .A2(n10915), .ZN(n10852) );
  NAND2_X1 U12719 ( .A1(n11165), .A2(n10852), .ZN(n10853) );
  NAND2_X1 U12720 ( .A1(n10853), .A2(n10862), .ZN(n10883) );
  OR2_X1 U12721 ( .A1(n10853), .A2(n10862), .ZN(n10854) );
  NAND2_X1 U12722 ( .A1(n10883), .A2(n10854), .ZN(n16468) );
  INV_X1 U12723 ( .A(n16468), .ZN(n10872) );
  OAI22_X1 U12724 ( .A1(n11536), .A2(n15232), .B1(n10915), .B2(n15230), .ZN(
        n10864) );
  NAND2_X1 U12725 ( .A1(n11114), .A2(n11113), .ZN(n11112) );
  OAI21_X1 U12726 ( .B1(n11157), .B2(n10915), .A(n16446), .ZN(n10859) );
  NAND2_X1 U12727 ( .A1(n11157), .A2(n10915), .ZN(n10858) );
  INV_X1 U12728 ( .A(n10888), .ZN(n10860) );
  AOI211_X1 U12729 ( .C1(n10862), .C2(n10861), .A(n16449), .B(n10860), .ZN(
        n10863) );
  AOI211_X1 U12730 ( .C1(n15166), .C2(n16468), .A(n10864), .B(n10863), .ZN(
        n16465) );
  MUX2_X1 U12731 ( .A(n10865), .B(n16465), .S(n15338), .Z(n10871) );
  INV_X1 U12732 ( .A(n10909), .ZN(n16463) );
  NOR2_X1 U12733 ( .A1(n11159), .A2(n16463), .ZN(n10866) );
  OR2_X1 U12734 ( .A1(n10897), .A2(n10866), .ZN(n16464) );
  INV_X1 U12735 ( .A(n10918), .ZN(n10867) );
  OAI22_X1 U12736 ( .A1(n15221), .A2(n16464), .B1(n10867), .B2(n15312), .ZN(
        n10869) );
  NOR2_X1 U12737 ( .A1(n15310), .A2(n16463), .ZN(n10868) );
  NOR2_X1 U12738 ( .A1(n10869), .A2(n10868), .ZN(n10870) );
  OAI211_X1 U12739 ( .C1(n10872), .C2(n15177), .A(n10871), .B(n10870), .ZN(
        P1_U3288) );
  INV_X1 U12740 ( .A(n10873), .ZN(n10874) );
  NAND2_X1 U12741 ( .A1(n14644), .A2(n10874), .ZN(n14629) );
  INV_X1 U12742 ( .A(n10875), .ZN(n10877) );
  AOI211_X1 U12743 ( .C1(n14296), .C2(n10877), .A(n10876), .B(n14571), .ZN(
        n10880) );
  OAI22_X1 U12744 ( .A1(n14644), .A2(n10276), .B1(n10878), .B2(n14641), .ZN(
        n10879) );
  NOR2_X1 U12745 ( .A1(n10880), .A2(n10879), .ZN(n10881) );
  OAI21_X1 U12746 ( .B1(n14246), .B2(n14629), .A(n10881), .ZN(P2_U3265) );
  OR2_X1 U12747 ( .A1(n10909), .A2(n14971), .ZN(n10882) );
  NAND2_X1 U12748 ( .A1(n10883), .A2(n10882), .ZN(n10884) );
  NAND2_X1 U12749 ( .A1(n10884), .A2(n10889), .ZN(n11527) );
  OR2_X1 U12750 ( .A1(n10884), .A2(n10889), .ZN(n10885) );
  NAND2_X1 U12751 ( .A1(n11527), .A2(n10885), .ZN(n10893) );
  INV_X1 U12752 ( .A(n10893), .ZN(n11078) );
  OR2_X1 U12753 ( .A1(n10909), .A2(n10886), .ZN(n10887) );
  NAND2_X1 U12754 ( .A1(n10890), .A2(n10889), .ZN(n10891) );
  NAND2_X1 U12755 ( .A1(n11539), .A2(n10891), .ZN(n10892) );
  NAND2_X1 U12756 ( .A1(n10892), .A2(n15431), .ZN(n10896) );
  AOI22_X1 U12757 ( .A1(n15331), .A2(n14971), .B1(n14969), .B2(n15329), .ZN(
        n10895) );
  NAND2_X1 U12758 ( .A1(n10893), .A2(n15166), .ZN(n10894) );
  AND3_X1 U12759 ( .A1(n10896), .A2(n10895), .A3(n10894), .ZN(n11071) );
  INV_X1 U12760 ( .A(n11537), .ZN(n11073) );
  NAND2_X1 U12761 ( .A1(n10897), .A2(n11073), .ZN(n11531) );
  OR2_X1 U12762 ( .A1(n10897), .A2(n11073), .ZN(n10898) );
  AND2_X1 U12763 ( .A1(n11531), .A2(n10898), .ZN(n11075) );
  AOI22_X1 U12764 ( .A1(n11075), .A2(n15471), .B1(n11537), .B2(n16445), .ZN(
        n10899) );
  OAI211_X1 U12765 ( .C1(n11078), .C2(n15475), .A(n11071), .B(n10899), .ZN(
        n10902) );
  NAND2_X1 U12766 ( .A1(n10902), .A2(n16553), .ZN(n10900) );
  OAI21_X1 U12767 ( .B1(n16553), .B2(n10901), .A(n10900), .ZN(P1_U3534) );
  NAND2_X1 U12768 ( .A1(n10902), .A2(n16556), .ZN(n10903) );
  OAI21_X1 U12769 ( .B1(n16556), .B2(n9379), .A(n10903), .ZN(P1_U3477) );
  NAND2_X1 U12770 ( .A1(n12698), .A2(n14971), .ZN(n10908) );
  NAND2_X1 U12771 ( .A1(n10909), .A2(n7456), .ZN(n10907) );
  AND2_X1 U12772 ( .A1(n10908), .A2(n10907), .ZN(n11140) );
  INV_X1 U12773 ( .A(n11140), .ZN(n11142) );
  NAND2_X1 U12774 ( .A1(n10909), .A2(n12687), .ZN(n10911) );
  NAND2_X1 U12775 ( .A1(n7456), .A2(n14971), .ZN(n10910) );
  NAND2_X1 U12776 ( .A1(n10911), .A2(n10910), .ZN(n10912) );
  XNOR2_X1 U12777 ( .A(n10912), .B(n7593), .ZN(n11141) );
  XNOR2_X1 U12778 ( .A(n11142), .B(n11141), .ZN(n10913) );
  XNOR2_X1 U12779 ( .A(n7609), .B(n10913), .ZN(n10920) );
  INV_X1 U12780 ( .A(n14952), .ZN(n14893) );
  OAI21_X1 U12781 ( .B1(n14958), .B2(n16463), .A(n10914), .ZN(n10917) );
  OAI22_X1 U12782 ( .A1(n14861), .A2(n10915), .B1(n11536), .B2(n14951), .ZN(
        n10916) );
  AOI211_X1 U12783 ( .C1(n10918), .C2(n14893), .A(n10917), .B(n10916), .ZN(
        n10919) );
  OAI21_X1 U12784 ( .B1(n10920), .B2(n11466), .A(n10919), .ZN(P1_U3227) );
  MUX2_X1 U12785 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n13357), .Z(n10953) );
  INV_X1 U12786 ( .A(n10921), .ZN(n10922) );
  MUX2_X1 U12787 ( .A(n10939), .B(n10929), .S(n13357), .Z(n16331) );
  NAND2_X1 U12788 ( .A1(n16331), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n11221) );
  AOI21_X1 U12789 ( .B1(n13751), .B2(n10922), .A(n11220), .ZN(n10955) );
  XOR2_X1 U12790 ( .A(n10954), .B(n10955), .Z(n10952) );
  NAND2_X1 U12791 ( .A1(n16079), .A2(n7728), .ZN(n16327) );
  INV_X1 U12792 ( .A(n10925), .ZN(n10923) );
  NAND2_X1 U12793 ( .A1(n10923), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13066) );
  NAND2_X1 U12794 ( .A1(n10924), .A2(n13066), .ZN(n10946) );
  NAND2_X1 U12795 ( .A1(n12961), .A2(n10925), .ZN(n10926) );
  AND2_X1 U12796 ( .A1(n10927), .A2(n10926), .ZN(n10944) );
  INV_X1 U12797 ( .A(n7728), .ZN(n13061) );
  INV_X1 U12798 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10928) );
  INV_X1 U12799 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10929) );
  NOR2_X1 U12800 ( .A1(n10929), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10930) );
  NAND2_X1 U12801 ( .A1(n8415), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10931) );
  OAI21_X1 U12802 ( .B1(n11228), .B2(n10930), .A(n10931), .ZN(n11217) );
  INV_X1 U12803 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n16382) );
  OAI21_X1 U12804 ( .B1(n10933), .B2(n10932), .A(n10957), .ZN(n10934) );
  INV_X1 U12805 ( .A(n10934), .ZN(n10949) );
  INV_X1 U12806 ( .A(n10938), .ZN(n10935) );
  INV_X1 U12807 ( .A(n10936), .ZN(n10937) );
  AND2_X1 U12808 ( .A1(n10938), .A2(n10937), .ZN(n16336) );
  INV_X1 U12809 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n16413) );
  NOR2_X1 U12810 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10939), .ZN(n16335) );
  INV_X1 U12811 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n16392) );
  NAND2_X1 U12812 ( .A1(n8415), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10940) );
  NAND2_X1 U12813 ( .A1(n11213), .A2(n10940), .ZN(n10941) );
  NAND2_X1 U12814 ( .A1(n10942), .A2(n10941), .ZN(n10965) );
  OAI21_X1 U12815 ( .B1(n10942), .B2(n10941), .A(n10965), .ZN(n10943) );
  NAND2_X1 U12816 ( .A1(n16336), .A2(n10943), .ZN(n10948) );
  INV_X1 U12817 ( .A(n10944), .ZN(n10945) );
  AND2_X1 U12818 ( .A1(n10946), .A2(n10945), .ZN(n16330) );
  AOI22_X1 U12819 ( .A1(n16330), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10947) );
  OAI211_X1 U12820 ( .C1(n10949), .C2(n16328), .A(n10948), .B(n10947), .ZN(
        n10950) );
  OAI21_X1 U12821 ( .B1(n10952), .B2(n16327), .A(n10951), .ZN(P3_U3184) );
  MUX2_X1 U12822 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n13357), .Z(n11006) );
  XNOR2_X1 U12823 ( .A(n11006), .B(n11008), .ZN(n11009) );
  OAI22_X1 U12824 ( .A1(n10955), .A2(n10954), .B1(n10953), .B2(n8249), .ZN(
        n11010) );
  XOR2_X1 U12825 ( .A(n11009), .B(n11010), .Z(n10975) );
  INV_X1 U12826 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n16426) );
  INV_X1 U12827 ( .A(n11008), .ZN(n10966) );
  NAND2_X1 U12828 ( .A1(n10958), .A2(n10966), .ZN(n11289) );
  OR2_X1 U12829 ( .A1(n10958), .A2(n10966), .ZN(n10959) );
  INV_X1 U12830 ( .A(n11291), .ZN(n10960) );
  AOI21_X1 U12831 ( .B1(n16426), .B2(n10961), .A(n10960), .ZN(n10963) );
  AOI22_X1 U12832 ( .A1(n16330), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n10962) );
  OAI21_X1 U12833 ( .B1(n10963), .B2(n16328), .A(n10962), .ZN(n10973) );
  NAND2_X1 U12834 ( .A1(n10965), .A2(n10964), .ZN(n10967) );
  NAND2_X1 U12835 ( .A1(n10967), .A2(n10966), .ZN(n11284) );
  OR2_X1 U12836 ( .A1(n10967), .A2(n10966), .ZN(n10968) );
  NAND2_X1 U12837 ( .A1(n11284), .A2(n10968), .ZN(n10970) );
  INV_X1 U12838 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10969) );
  NAND2_X1 U12839 ( .A1(n10970), .A2(n10969), .ZN(n10971) );
  AOI21_X1 U12840 ( .B1(n11285), .B2(n10971), .A(n13368), .ZN(n10972) );
  AOI211_X1 U12841 ( .C1(n13370), .C2(n11008), .A(n10973), .B(n10972), .ZN(
        n10974) );
  OAI21_X1 U12842 ( .B1(n10975), .B2(n16327), .A(n10974), .ZN(P3_U3185) );
  INV_X1 U12843 ( .A(n10981), .ZN(n10977) );
  NAND2_X1 U12844 ( .A1(n10978), .A2(n11900), .ZN(n10980) );
  AOI22_X1 U12845 ( .A1(n11192), .A2(n10048), .B1(n10051), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n10979) );
  NAND2_X2 U12846 ( .A1(n10980), .A2(n10979), .ZN(n14060) );
  XNOR2_X1 U12847 ( .A(n14060), .B(n7463), .ZN(n11346) );
  NAND2_X1 U12848 ( .A1(n14313), .A2(n7458), .ZN(n11338) );
  INV_X1 U12849 ( .A(n14314), .ZN(n11242) );
  NAND2_X1 U12850 ( .A1(n10981), .A2(n13977), .ZN(n10982) );
  OAI21_X1 U12851 ( .B1(n13967), .B2(n11242), .A(n10982), .ZN(n10983) );
  NAND3_X1 U12852 ( .A1(n10984), .A2(n7603), .A3(n10983), .ZN(n11004) );
  NAND2_X1 U12853 ( .A1(n13902), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10994) );
  INV_X1 U12854 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10985) );
  OR2_X1 U12855 ( .A1(n10986), .A2(n10985), .ZN(n10993) );
  INV_X1 U12856 ( .A(n10989), .ZN(n10987) );
  INV_X1 U12857 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10988) );
  NAND2_X1 U12858 ( .A1(n10989), .A2(n10988), .ZN(n10990) );
  NAND2_X1 U12859 ( .A1(n11355), .A2(n10990), .ZN(n11506) );
  OR2_X1 U12860 ( .A1(n10059), .A2(n11506), .ZN(n10992) );
  INV_X1 U12861 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11507) );
  OR2_X1 U12862 ( .A1(n14192), .A2(n11507), .ZN(n10991) );
  NAND4_X1 U12863 ( .A1(n10994), .A2(n10993), .A3(n10992), .A4(n10991), .ZN(
        n14312) );
  NAND2_X1 U12864 ( .A1(n14312), .A2(n14614), .ZN(n10996) );
  NAND2_X1 U12865 ( .A1(n14314), .A2(n14613), .ZN(n10995) );
  NAND2_X1 U12866 ( .A1(n10996), .A2(n10995), .ZN(n11245) );
  INV_X1 U12867 ( .A(n11245), .ZN(n10998) );
  OAI22_X1 U12868 ( .A1(n13975), .A2(n10998), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10997), .ZN(n10999) );
  INV_X1 U12869 ( .A(n10999), .ZN(n11003) );
  NAND2_X1 U12870 ( .A1(n14060), .A2(n13952), .ZN(n11002) );
  INV_X1 U12871 ( .A(n11000), .ZN(n11559) );
  NAND2_X1 U12872 ( .A1(n13972), .A2(n11559), .ZN(n11001) );
  AND4_X1 U12873 ( .A1(n11004), .A2(n11003), .A3(n11002), .A4(n11001), .ZN(
        n11005) );
  OAI21_X1 U12874 ( .B1(n11350), .B2(n13915), .A(n11005), .ZN(P2_U3203) );
  MUX2_X1 U12875 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n13357), .Z(n11027) );
  XNOR2_X1 U12876 ( .A(n11027), .B(n11029), .ZN(n11030) );
  INV_X1 U12877 ( .A(n11006), .ZN(n11007) );
  AOI22_X1 U12878 ( .A1(n11010), .A2(n11009), .B1(n11008), .B2(n11007), .ZN(
        n11281) );
  MUX2_X1 U12879 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13357), .Z(n11011) );
  XOR2_X1 U12880 ( .A(n11015), .B(n11011), .Z(n11282) );
  OAI22_X1 U12881 ( .A1(n11281), .A2(n11282), .B1(n11011), .B2(n11296), .ZN(
        n11031) );
  XOR2_X1 U12882 ( .A(n11030), .B(n11031), .Z(n11026) );
  INV_X1 U12883 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n11523) );
  INV_X1 U12884 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11598) );
  MUX2_X1 U12885 ( .A(n11598), .B(P3_REG2_REG_4__SCAN_IN), .S(n11015), .Z(
        n11283) );
  INV_X1 U12886 ( .A(n11029), .ZN(n11017) );
  INV_X1 U12887 ( .A(n11403), .ZN(n11013) );
  AOI21_X1 U12888 ( .B1(n11523), .B2(n11014), .A(n11013), .ZN(n11023) );
  NOR2_X1 U12889 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15774), .ZN(n11652) );
  INV_X1 U12890 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n16441) );
  MUX2_X1 U12891 ( .A(n16441), .B(P3_REG1_REG_4__SCAN_IN), .S(n11015), .Z(
        n11288) );
  NAND2_X1 U12892 ( .A1(n11296), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n11016) );
  INV_X1 U12893 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n16460) );
  NAND2_X1 U12894 ( .A1(n11019), .A2(n16460), .ZN(n11020) );
  AOI21_X1 U12895 ( .B1(n11409), .B2(n11020), .A(n16328), .ZN(n11021) );
  AOI211_X1 U12896 ( .C1(n16330), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n11652), .B(
        n11021), .ZN(n11022) );
  OAI21_X1 U12897 ( .B1(n11023), .B2(n13368), .A(n11022), .ZN(n11024) );
  AOI21_X1 U12898 ( .B1(n11029), .B2(n13370), .A(n11024), .ZN(n11025) );
  OAI21_X1 U12899 ( .B1(n11026), .B2(n16327), .A(n11025), .ZN(P3_U3187) );
  MUX2_X1 U12900 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n13357), .Z(n11256) );
  XNOR2_X1 U12901 ( .A(n11256), .B(n11258), .ZN(n11259) );
  INV_X1 U12902 ( .A(n11027), .ZN(n11028) );
  AOI22_X1 U12903 ( .A1(n11031), .A2(n11030), .B1(n11029), .B2(n11028), .ZN(
        n11398) );
  MUX2_X1 U12904 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n13357), .Z(n11032) );
  XNOR2_X1 U12905 ( .A(n11032), .B(n11418), .ZN(n11397) );
  OAI22_X1 U12906 ( .A1(n11398), .A2(n11397), .B1(n11032), .B2(n11418), .ZN(
        n11260) );
  XOR2_X1 U12907 ( .A(n11259), .B(n11260), .Z(n11052) );
  INV_X1 U12908 ( .A(n16330), .ZN(n13345) );
  INV_X1 U12909 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15938) );
  INV_X1 U12910 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n11033) );
  NOR2_X1 U12911 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11033), .ZN(n11882) );
  INV_X1 U12912 ( .A(n11882), .ZN(n11034) );
  OAI21_X1 U12913 ( .B1(n13345), .B2(n15938), .A(n11034), .ZN(n11050) );
  INV_X1 U12914 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11038) );
  INV_X1 U12915 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n16475) );
  MUX2_X1 U12916 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n16475), .S(n11418), .Z(
        n11406) );
  NAND2_X1 U12917 ( .A1(n11418), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n11035) );
  INV_X1 U12918 ( .A(n11258), .ZN(n11042) );
  INV_X1 U12919 ( .A(n11274), .ZN(n11036) );
  AOI21_X1 U12920 ( .B1(n11038), .B2(n11037), .A(n11036), .ZN(n11048) );
  INV_X1 U12921 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11046) );
  INV_X1 U12922 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11039) );
  MUX2_X1 U12923 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n11039), .S(n11418), .Z(
        n11400) );
  NAND2_X1 U12924 ( .A1(n11040), .A2(n11400), .ZN(n11405) );
  NAND2_X1 U12925 ( .A1(n11418), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n11041) );
  NAND2_X1 U12926 ( .A1(n11405), .A2(n11041), .ZN(n11043) );
  NAND2_X1 U12927 ( .A1(n11043), .A2(n11042), .ZN(n11263) );
  OAI21_X1 U12928 ( .B1(n11043), .B2(n11042), .A(n11263), .ZN(n11045) );
  INV_X1 U12929 ( .A(n11265), .ZN(n11044) );
  AOI21_X1 U12930 ( .B1(n11046), .B2(n11045), .A(n11044), .ZN(n11047) );
  OAI22_X1 U12931 ( .A1(n11048), .A2(n16328), .B1(n11047), .B2(n13368), .ZN(
        n11049) );
  AOI211_X1 U12932 ( .C1(n11258), .C2(n13370), .A(n11050), .B(n11049), .ZN(
        n11051) );
  OAI21_X1 U12933 ( .B1(n11052), .B2(n16327), .A(n11051), .ZN(P3_U3189) );
  OR2_X1 U12934 ( .A1(n14044), .A2(n14315), .ZN(n11054) );
  XNOR2_X1 U12935 ( .A(n14052), .B(n11242), .ZN(n14258) );
  INV_X1 U12936 ( .A(n14258), .ZN(n11055) );
  NAND2_X1 U12937 ( .A1(n11056), .A2(n11055), .ZN(n11057) );
  NAND2_X1 U12938 ( .A1(n11237), .A2(n11057), .ZN(n11553) );
  OR2_X1 U12939 ( .A1(n14044), .A2(n14046), .ZN(n11058) );
  XNOR2_X1 U12940 ( .A(n11241), .B(n14258), .ZN(n11061) );
  AOI21_X1 U12941 ( .B1(n11061), .B2(n7449), .A(n11060), .ZN(n11558) );
  INV_X1 U12942 ( .A(n11062), .ZN(n11064) );
  INV_X1 U12943 ( .A(n14052), .ZN(n11552) );
  NAND2_X1 U12944 ( .A1(n11552), .A2(n11062), .ZN(n11247) );
  INV_X1 U12945 ( .A(n11247), .ZN(n11063) );
  AOI211_X1 U12946 ( .C1(n14052), .C2(n11064), .A(n7458), .B(n11063), .ZN(
        n11556) );
  AOI21_X1 U12947 ( .B1(n14709), .B2(n14052), .A(n11556), .ZN(n11065) );
  OAI211_X1 U12948 ( .C1(n14735), .C2(n11553), .A(n11558), .B(n11065), .ZN(
        n11234) );
  NAND2_X1 U12949 ( .A1(n11234), .A2(n12115), .ZN(n11066) );
  OAI21_X1 U12950 ( .B1(n16534), .B2(n10733), .A(n11066), .ZN(P2_U3454) );
  INV_X1 U12951 ( .A(n11067), .ZN(n11069) );
  OAI222_X1 U12952 ( .A1(P3_U3151), .A2(n11070), .B1(n13750), .B2(n11069), 
        .C1(n11068), .C2(n13745), .ZN(P3_U3274) );
  MUX2_X1 U12953 ( .A(n11072), .B(n11071), .S(n15338), .Z(n11077) );
  OAI22_X1 U12954 ( .A1(n15310), .A2(n11073), .B1(n15312), .B2(n11152), .ZN(
        n11074) );
  AOI21_X1 U12955 ( .B1(n15347), .B2(n11075), .A(n11074), .ZN(n11076) );
  OAI211_X1 U12956 ( .C1(n11078), .C2(n15177), .A(n11077), .B(n11076), .ZN(
        P1_U3287) );
  INV_X1 U12957 ( .A(n11079), .ZN(n11081) );
  XNOR2_X1 U12958 ( .A(n12834), .B(n16422), .ZN(n11468) );
  XNOR2_X1 U12959 ( .A(n11468), .B(n11590), .ZN(n11082) );
  OAI211_X1 U12960 ( .C1(n11083), .C2(n11082), .A(n11469), .B(n13183), .ZN(
        n11090) );
  INV_X1 U12961 ( .A(n13185), .ZN(n13198) );
  OAI22_X1 U12962 ( .A1(n13198), .A2(n16373), .B1(n13199), .B2(n11084), .ZN(
        n11088) );
  INV_X1 U12963 ( .A(n13066), .ZN(n11085) );
  MUX2_X1 U12964 ( .A(n13202), .B(P3_U3151), .S(P3_REG3_REG_3__SCAN_IN), .Z(
        n11087) );
  AOI211_X1 U12965 ( .C1(n13196), .C2(n13224), .A(n11088), .B(n11087), .ZN(
        n11089) );
  NAND2_X1 U12966 ( .A1(n11090), .A2(n11089), .ZN(P3_U3158) );
  INV_X1 U12967 ( .A(n11091), .ZN(n11094) );
  INV_X1 U12968 ( .A(n11479), .ZN(n11092) );
  NAND2_X1 U12969 ( .A1(n13972), .A2(n11092), .ZN(n11093) );
  NAND2_X1 U12970 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n16144) );
  OAI211_X1 U12971 ( .C1(n13975), .C2(n11094), .A(n11093), .B(n16144), .ZN(
        n11100) );
  AOI22_X1 U12972 ( .A1(n13957), .A2(n14318), .B1(n13977), .B2(n11095), .ZN(
        n11098) );
  INV_X1 U12973 ( .A(n12780), .ZN(n11097) );
  NOR3_X1 U12974 ( .A1(n11098), .A2(n11097), .A3(n11096), .ZN(n11099) );
  AOI211_X1 U12975 ( .C1(n14032), .C2(n13952), .A(n11100), .B(n11099), .ZN(
        n11101) );
  OAI21_X1 U12976 ( .B1(n11102), .B2(n13915), .A(n11101), .ZN(P2_U3199) );
  OAI22_X1 U12977 ( .A1(n13064), .A2(P3_U3151), .B1(SI_22_), .B2(n13745), .ZN(
        n11103) );
  AOI21_X1 U12978 ( .B1(n11104), .B2(n13739), .A(n11103), .ZN(P3_U3273) );
  OR2_X1 U12979 ( .A1(n11106), .A2(n11105), .ZN(n11107) );
  NAND2_X1 U12980 ( .A1(n11108), .A2(n11107), .ZN(n16434) );
  INV_X1 U12981 ( .A(n16434), .ZN(n11122) );
  INV_X1 U12982 ( .A(n15310), .ZN(n15343) );
  NAND2_X1 U12983 ( .A1(n11109), .A2(n14843), .ZN(n11110) );
  OAI22_X1 U12984 ( .A1(n15221), .A2(n16430), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n15312), .ZN(n11111) );
  AOI21_X1 U12985 ( .B1(n15343), .B2(n14843), .A(n11111), .ZN(n11121) );
  NAND2_X1 U12986 ( .A1(n16434), .A2(n15166), .ZN(n11118) );
  OAI21_X1 U12987 ( .B1(n11114), .B2(n11113), .A(n11112), .ZN(n11115) );
  NAND2_X1 U12988 ( .A1(n11115), .A2(n15431), .ZN(n11117) );
  AOI22_X1 U12989 ( .A1(n14972), .A2(n15329), .B1(n15331), .B2(n9332), .ZN(
        n11116) );
  AND3_X1 U12990 ( .A1(n11118), .A2(n11117), .A3(n11116), .ZN(n16431) );
  MUX2_X1 U12991 ( .A(n16431), .B(n11119), .S(n15295), .Z(n11120) );
  OAI211_X1 U12992 ( .C1(n11122), .C2(n15177), .A(n11121), .B(n11120), .ZN(
        P1_U3290) );
  OAI22_X1 U12993 ( .A1(n15295), .A2(n11124), .B1(n11123), .B2(n15312), .ZN(
        n11125) );
  AOI21_X1 U12994 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n15333), .A(n11125), .ZN(
        n11128) );
  OAI21_X1 U12995 ( .B1(n15347), .B2(n15343), .A(n11126), .ZN(n11127) );
  OAI211_X1 U12996 ( .C1(n11129), .C2(n15177), .A(n11128), .B(n11127), .ZN(
        P1_U3293) );
  OAI21_X1 U12997 ( .B1(n11130), .B2(n13017), .A(n12863), .ZN(n16409) );
  NAND2_X1 U12998 ( .A1(n16409), .A2(n13661), .ZN(n11137) );
  NAND3_X1 U12999 ( .A1(n16369), .A2(n13017), .A3(n11132), .ZN(n11133) );
  NAND2_X1 U13000 ( .A1(n11131), .A2(n11133), .ZN(n11135) );
  OAI22_X1 U13001 ( .A1(n8573), .A2(n16374), .B1(n11590), .B2(n16372), .ZN(
        n11134) );
  AOI21_X1 U13002 ( .B1(n11135), .B2(n16377), .A(n11134), .ZN(n11136) );
  AND2_X1 U13003 ( .A1(n11137), .A2(n11136), .ZN(n16406) );
  NAND2_X1 U13004 ( .A1(n16569), .A2(n8515), .ZN(n13735) );
  INV_X1 U13005 ( .A(n13735), .ZN(n11927) );
  AOI22_X1 U13006 ( .A1(n11927), .A2(n16409), .B1(P3_REG0_REG_2__SCAN_IN), 
        .B2(n16566), .ZN(n11139) );
  INV_X1 U13007 ( .A(n13731), .ZN(n13701) );
  NAND2_X1 U13008 ( .A1(n13701), .A2(n16402), .ZN(n11138) );
  OAI211_X1 U13009 ( .C1(n16406), .C2(n16566), .A(n11139), .B(n11138), .ZN(
        P3_U3396) );
  NAND2_X1 U13010 ( .A1(n11141), .A2(n11140), .ZN(n11144) );
  INV_X1 U13011 ( .A(n11141), .ZN(n11143) );
  NAND2_X1 U13012 ( .A1(n11537), .A2(n12687), .ZN(n11146) );
  NAND2_X1 U13013 ( .A1(n7456), .A2(n14970), .ZN(n11145) );
  NAND2_X1 U13014 ( .A1(n11146), .A2(n11145), .ZN(n11147) );
  INV_X2 U13015 ( .A(n7593), .ZN(n12705) );
  XNOR2_X1 U13016 ( .A(n11147), .B(n12705), .ZN(n11454) );
  NAND2_X1 U13017 ( .A1(n11537), .A2(n7456), .ZN(n11149) );
  NAND2_X1 U13018 ( .A1(n12698), .A2(n14970), .ZN(n11148) );
  NAND2_X1 U13019 ( .A1(n11149), .A2(n11148), .ZN(n11453) );
  XNOR2_X1 U13020 ( .A(n11454), .B(n11453), .ZN(n11457) );
  XNOR2_X1 U13021 ( .A(n11458), .B(n11457), .ZN(n11156) );
  INV_X1 U13022 ( .A(n14969), .ZN(n11742) );
  NAND2_X1 U13023 ( .A1(n14955), .A2(n14971), .ZN(n11151) );
  OAI211_X1 U13024 ( .C1(n11742), .C2(n14951), .A(n11151), .B(n11150), .ZN(
        n11154) );
  NOR2_X1 U13025 ( .A1(n14952), .A2(n11152), .ZN(n11153) );
  AOI211_X1 U13026 ( .C1(n11537), .C2(n14844), .A(n11154), .B(n11153), .ZN(
        n11155) );
  OAI21_X1 U13027 ( .B1(n11156), .B2(n11466), .A(n11155), .ZN(P1_U3239) );
  XNOR2_X1 U13028 ( .A(n11157), .B(n11166), .ZN(n16450) );
  NOR2_X1 U13029 ( .A1(n15333), .A2(n16449), .ZN(n15265) );
  INV_X1 U13030 ( .A(n15265), .ZN(n15211) );
  INV_X1 U13031 ( .A(n11158), .ZN(n16444) );
  MUX2_X1 U13032 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n16444), .S(n15338), .Z(
        n11162) );
  OR2_X1 U13033 ( .A1(n7611), .A2(n11159), .ZN(n16448) );
  OAI22_X1 U13034 ( .A1(n15221), .A2(n16448), .B1(n11160), .B2(n15312), .ZN(
        n11161) );
  AOI211_X1 U13035 ( .C1(n15343), .C2(n16446), .A(n11162), .B(n11161), .ZN(
        n11169) );
  INV_X1 U13036 ( .A(n11163), .ZN(n11164) );
  NAND2_X1 U13037 ( .A1(n15338), .A2(n11164), .ZN(n15337) );
  OAI21_X1 U13038 ( .B1(n11167), .B2(n11166), .A(n11165), .ZN(n16453) );
  NAND2_X1 U13039 ( .A1(n15309), .A2(n16453), .ZN(n11168) );
  OAI211_X1 U13040 ( .C1(n16450), .C2(n15211), .A(n11169), .B(n11168), .ZN(
        P1_U3289) );
  XNOR2_X1 U13041 ( .A(n11775), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n11626) );
  INV_X1 U13042 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11686) );
  MUX2_X1 U13043 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n11449), .S(n16094), .Z(
        n16084) );
  NAND3_X1 U13044 ( .A1(n16084), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_REG2_REG_0__SCAN_IN), .ZN(n16085) );
  OAI21_X1 U13045 ( .B1(n8493), .B2(n11449), .A(n16085), .ZN(n16099) );
  MUX2_X1 U13046 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n11331), .S(n16107), .Z(
        n16100) );
  NAND2_X1 U13047 ( .A1(n16099), .A2(n16100), .ZN(n16098) );
  OAI21_X1 U13048 ( .B1(n11331), .B2(n11170), .A(n16098), .ZN(n16114) );
  MUX2_X1 U13049 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n11171), .S(n11184), .Z(
        n16115) );
  NAND2_X1 U13050 ( .A1(n16114), .A2(n16115), .ZN(n16113) );
  OAI21_X1 U13051 ( .B1(n16117), .B2(n11171), .A(n16113), .ZN(n16126) );
  MUX2_X1 U13052 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11172), .S(n11186), .Z(
        n16127) );
  NAND2_X1 U13053 ( .A1(n16126), .A2(n16127), .ZN(n16125) );
  OAI21_X1 U13054 ( .B1(n11172), .B2(n16129), .A(n16125), .ZN(n16138) );
  XNOR2_X1 U13055 ( .A(n16141), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n16139) );
  NAND2_X1 U13056 ( .A1(n16138), .A2(n16139), .ZN(n16137) );
  OAI21_X1 U13057 ( .B1(n16141), .B2(n11480), .A(n16137), .ZN(n16148) );
  MUX2_X1 U13058 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11369), .S(n16156), .Z(
        n16149) );
  NAND2_X1 U13059 ( .A1(n16148), .A2(n16149), .ZN(n16147) );
  OAI21_X1 U13060 ( .B1(n11369), .B2(n11173), .A(n16147), .ZN(n14333) );
  XOR2_X1 U13061 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n14331), .Z(n14334) );
  NAND2_X1 U13062 ( .A1(n14333), .A2(n14334), .ZN(n14332) );
  OAI21_X1 U13063 ( .B1(n11175), .B2(n11174), .A(n14332), .ZN(n16161) );
  MUX2_X1 U13064 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n11177), .S(n16169), .Z(
        n16162) );
  NAND2_X1 U13065 ( .A1(n16161), .A2(n16162), .ZN(n16160) );
  OAI21_X1 U13066 ( .B1(n11177), .B2(n11176), .A(n16160), .ZN(n16245) );
  MUX2_X1 U13067 ( .A(n11178), .B(P2_REG2_REG_9__SCAN_IN), .S(n11192), .Z(
        n16246) );
  NOR2_X1 U13068 ( .A1(n16245), .A2(n16246), .ZN(n16244) );
  AOI21_X1 U13069 ( .B1(n11178), .B2(n16238), .A(n16244), .ZN(n16225) );
  MUX2_X1 U13070 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n11507), .S(n16233), .Z(
        n16224) );
  NAND2_X1 U13071 ( .A1(n16225), .A2(n16224), .ZN(n16223) );
  OAI21_X1 U13072 ( .B1(n11507), .B2(n11179), .A(n16223), .ZN(n16173) );
  MUX2_X1 U13073 ( .A(n11686), .B(P2_REG2_REG_11__SCAN_IN), .S(n16181), .Z(
        n16174) );
  NOR2_X1 U13074 ( .A1(n16173), .A2(n16174), .ZN(n16172) );
  AOI21_X1 U13075 ( .B1(n11686), .B2(n11180), .A(n16172), .ZN(n11627) );
  XOR2_X1 U13076 ( .A(n11626), .B(n11627), .Z(n11202) );
  INV_X1 U13077 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n11181) );
  MUX2_X1 U13078 ( .A(n11181), .B(P2_REG1_REG_1__SCAN_IN), .S(n16094), .Z(
        n16090) );
  NOR3_X1 U13079 ( .A1(n16090), .A2(n10277), .A3(n10041), .ZN(n16089) );
  AOI21_X1 U13080 ( .B1(n16094), .B2(P2_REG1_REG_1__SCAN_IN), .A(n16089), .ZN(
        n16104) );
  INV_X1 U13081 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n11182) );
  MUX2_X1 U13082 ( .A(n11182), .B(P2_REG1_REG_2__SCAN_IN), .S(n16107), .Z(
        n16103) );
  MUX2_X1 U13083 ( .A(n11183), .B(P2_REG1_REG_3__SCAN_IN), .S(n11184), .Z(
        n16111) );
  NOR2_X1 U13084 ( .A1(n16112), .A2(n16111), .ZN(n16110) );
  AOI21_X1 U13085 ( .B1(n11184), .B2(P2_REG1_REG_3__SCAN_IN), .A(n16110), .ZN(
        n16124) );
  INV_X1 U13086 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n11185) );
  MUX2_X1 U13087 ( .A(n11185), .B(P2_REG1_REG_4__SCAN_IN), .S(n11186), .Z(
        n16123) );
  XNOR2_X1 U13088 ( .A(n11187), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n16135) );
  NOR2_X1 U13089 ( .A1(n16136), .A2(n16135), .ZN(n16134) );
  AOI21_X1 U13090 ( .B1(n11187), .B2(P2_REG1_REG_5__SCAN_IN), .A(n16134), .ZN(
        n16153) );
  INV_X1 U13091 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n11188) );
  MUX2_X1 U13092 ( .A(n11188), .B(P2_REG1_REG_6__SCAN_IN), .S(n16156), .Z(
        n16152) );
  MUX2_X1 U13093 ( .A(n11189), .B(P2_REG1_REG_7__SCAN_IN), .S(n14331), .Z(
        n14325) );
  NOR2_X1 U13094 ( .A1(n14326), .A2(n14325), .ZN(n14324) );
  AOI21_X1 U13095 ( .B1(n14331), .B2(P2_REG1_REG_7__SCAN_IN), .A(n14324), .ZN(
        n16166) );
  INV_X1 U13096 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n11190) );
  MUX2_X1 U13097 ( .A(n11190), .B(P2_REG1_REG_8__SCAN_IN), .S(n16169), .Z(
        n16165) );
  MUX2_X1 U13098 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n11191), .S(n11192), .Z(
        n16242) );
  NAND2_X1 U13099 ( .A1(n16243), .A2(n16242), .ZN(n16241) );
  OAI21_X1 U13100 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n11192), .A(n16241), .ZN(
        n16229) );
  INV_X1 U13101 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n11193) );
  MUX2_X1 U13102 ( .A(n11193), .B(P2_REG1_REG_10__SCAN_IN), .S(n16233), .Z(
        n16230) );
  NOR2_X1 U13103 ( .A1(n16229), .A2(n16230), .ZN(n16227) );
  AOI21_X1 U13104 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n16233), .A(n16227), 
        .ZN(n16178) );
  INV_X1 U13105 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11194) );
  MUX2_X1 U13106 ( .A(n11194), .B(P2_REG1_REG_11__SCAN_IN), .S(n16181), .Z(
        n16177) );
  INV_X1 U13107 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11610) );
  MUX2_X1 U13108 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n11610), .S(n11775), .Z(
        n11195) );
  NAND2_X1 U13109 ( .A1(n11196), .A2(n11195), .ZN(n11622) );
  OAI21_X1 U13110 ( .B1(n11196), .B2(n11195), .A(n11622), .ZN(n11200) );
  NAND2_X1 U13111 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n12717)
         );
  NAND2_X1 U13112 ( .A1(n16097), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n11197) );
  OAI211_X1 U13113 ( .C1(n16189), .C2(n11198), .A(n12717), .B(n11197), .ZN(
        n11199) );
  AOI21_X1 U13114 ( .B1(n11200), .B2(n16250), .A(n11199), .ZN(n11201) );
  OAI21_X1 U13115 ( .B1(n16247), .B2(n11202), .A(n11201), .ZN(P2_U3226) );
  NAND2_X1 U13116 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n11203), .ZN(n11206) );
  NAND2_X1 U13117 ( .A1(n11204), .A2(n14947), .ZN(n11205) );
  OAI211_X1 U13118 ( .C1(n14958), .C2(n11207), .A(n11206), .B(n11205), .ZN(
        n11208) );
  AOI21_X1 U13119 ( .B1(n14845), .B2(n10517), .A(n11208), .ZN(n11209) );
  INV_X1 U13120 ( .A(n11209), .ZN(P1_U3232) );
  NAND2_X1 U13121 ( .A1(n14740), .A2(n11210), .ZN(n11211) );
  OAI21_X1 U13122 ( .B1(n14740), .B2(n10277), .A(n11211), .ZN(P2_U3499) );
  INV_X1 U13123 ( .A(n13370), .ZN(n16333) );
  INV_X1 U13124 ( .A(n11212), .ZN(n11214) );
  OAI21_X1 U13125 ( .B1(n11214), .B2(P3_REG2_REG_1__SCAN_IN), .A(n11213), .ZN(
        n11226) );
  INV_X1 U13126 ( .A(n11215), .ZN(n11216) );
  AOI21_X1 U13127 ( .B1(n16382), .B2(n11217), .A(n11216), .ZN(n11219) );
  AOI22_X1 U13128 ( .A1(n16330), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n11218) );
  OAI21_X1 U13129 ( .B1(n11219), .B2(n16328), .A(n11218), .ZN(n11225) );
  AOI21_X1 U13130 ( .B1(n11222), .B2(n11221), .A(n11220), .ZN(n11223) );
  NOR2_X1 U13131 ( .A1(n11223), .A2(n16327), .ZN(n11224) );
  AOI211_X1 U13132 ( .C1(n16336), .C2(n11226), .A(n11225), .B(n11224), .ZN(
        n11227) );
  OAI21_X1 U13133 ( .B1(n11228), .B2(n16333), .A(n11227), .ZN(P3_U3183) );
  NAND2_X1 U13134 ( .A1(n11229), .A2(n14740), .ZN(n11230) );
  OAI21_X1 U13135 ( .B1(n14740), .B2(n11189), .A(n11230), .ZN(P2_U3506) );
  INV_X1 U13136 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n11233) );
  NAND2_X1 U13137 ( .A1(n11231), .A2(n14740), .ZN(n11232) );
  OAI21_X1 U13138 ( .B1(n14740), .B2(n11233), .A(n11232), .ZN(P2_U3504) );
  NAND2_X1 U13139 ( .A1(n11234), .A2(n14740), .ZN(n11235) );
  OAI21_X1 U13140 ( .B1(n14740), .B2(n11190), .A(n11235), .ZN(P2_U3507) );
  INV_X1 U13141 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11250) );
  NAND2_X1 U13142 ( .A1(n14052), .A2(n14314), .ZN(n11236) );
  XNOR2_X1 U13143 ( .A(n14060), .B(n14062), .ZN(n14259) );
  OR2_X1 U13144 ( .A1(n11238), .A2(n14259), .ZN(n11239) );
  NAND2_X1 U13145 ( .A1(n11499), .A2(n11239), .ZN(n11562) );
  NAND2_X1 U13146 ( .A1(n14052), .A2(n11242), .ZN(n11240) );
  OR2_X1 U13147 ( .A1(n14052), .A2(n11242), .ZN(n11243) );
  XNOR2_X1 U13148 ( .A(n11501), .B(n14259), .ZN(n11246) );
  AOI21_X1 U13149 ( .B1(n11246), .B2(n7449), .A(n11245), .ZN(n11567) );
  AOI211_X1 U13150 ( .C1(n14060), .C2(n11247), .A(n7458), .B(n7989), .ZN(
        n11565) );
  AOI21_X1 U13151 ( .B1(n14709), .B2(n14060), .A(n11565), .ZN(n11248) );
  OAI211_X1 U13152 ( .C1(n14735), .C2(n11562), .A(n11567), .B(n11248), .ZN(
        n11251) );
  NAND2_X1 U13153 ( .A1(n11251), .A2(n12115), .ZN(n11249) );
  OAI21_X1 U13154 ( .B1(n16534), .B2(n11250), .A(n11249), .ZN(P2_U3457) );
  NAND2_X1 U13155 ( .A1(n11251), .A2(n14740), .ZN(n11252) );
  OAI21_X1 U13156 ( .B1(n14740), .B2(n11191), .A(n11252), .ZN(P2_U3508) );
  MUX2_X1 U13157 ( .A(n10928), .B(n16406), .S(n16565), .Z(n11255) );
  INV_X1 U13158 ( .A(n13657), .ZN(n13624) );
  NAND2_X1 U13159 ( .A1(n16565), .A2(n8515), .ZN(n13664) );
  INV_X1 U13160 ( .A(n13664), .ZN(n11253) );
  AOI22_X1 U13161 ( .A1(n16402), .A2(n13624), .B1(n11253), .B2(n16409), .ZN(
        n11254) );
  NAND2_X1 U13162 ( .A1(n11255), .A2(n11254), .ZN(P3_U3461) );
  MUX2_X1 U13163 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n13357), .Z(n11424) );
  XNOR2_X1 U13164 ( .A(n11424), .B(n11431), .ZN(n11425) );
  INV_X1 U13165 ( .A(n11256), .ZN(n11257) );
  AOI22_X1 U13166 ( .A1(n11260), .A2(n11259), .B1(n11258), .B2(n11257), .ZN(
        n11426) );
  XOR2_X1 U13167 ( .A(n11425), .B(n11426), .Z(n11280) );
  NAND2_X1 U13168 ( .A1(n11265), .A2(n11263), .ZN(n11261) );
  INV_X1 U13169 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11986) );
  XNOR2_X1 U13170 ( .A(n11431), .B(n11986), .ZN(n11262) );
  NAND2_X1 U13171 ( .A1(n11261), .A2(n11262), .ZN(n11420) );
  INV_X1 U13172 ( .A(n11262), .ZN(n11264) );
  NAND3_X1 U13173 ( .A1(n11265), .A2(n11264), .A3(n11263), .ZN(n11266) );
  AOI21_X1 U13174 ( .B1(n11420), .B2(n11266), .A(n13368), .ZN(n11278) );
  NOR2_X1 U13175 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11267), .ZN(n11934) );
  AOI21_X1 U13176 ( .B1(n16330), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11934), .ZN(
        n11268) );
  OAI21_X1 U13177 ( .B1(n16333), .B2(n11431), .A(n11268), .ZN(n11277) );
  NAND2_X1 U13178 ( .A1(n11274), .A2(n11272), .ZN(n11270) );
  INV_X1 U13179 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11269) );
  XNOR2_X1 U13180 ( .A(n11431), .B(n11269), .ZN(n11271) );
  INV_X1 U13181 ( .A(n11271), .ZN(n11273) );
  NAND3_X1 U13182 ( .A1(n11274), .A2(n11273), .A3(n11272), .ZN(n11275) );
  AOI21_X1 U13183 ( .B1(n11433), .B2(n11275), .A(n16328), .ZN(n11276) );
  NOR3_X1 U13184 ( .A1(n11278), .A2(n11277), .A3(n11276), .ZN(n11279) );
  OAI21_X1 U13185 ( .B1(n11280), .B2(n16327), .A(n11279), .ZN(P3_U3190) );
  XOR2_X1 U13186 ( .A(n11282), .B(n11281), .Z(n11301) );
  NAND3_X1 U13187 ( .A1(n11285), .A2(n8238), .A3(n11284), .ZN(n11286) );
  NAND2_X1 U13188 ( .A1(n11287), .A2(n11286), .ZN(n11299) );
  INV_X1 U13189 ( .A(n11288), .ZN(n11290) );
  NAND3_X1 U13190 ( .A1(n11291), .A2(n11290), .A3(n11289), .ZN(n11292) );
  AND2_X1 U13191 ( .A1(n11293), .A2(n11292), .ZN(n11295) );
  NAND2_X1 U13192 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n11473) );
  NAND2_X1 U13193 ( .A1(n16330), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n11294) );
  OAI211_X1 U13194 ( .C1(n16328), .C2(n11295), .A(n11473), .B(n11294), .ZN(
        n11298) );
  NOR2_X1 U13195 ( .A1(n16333), .A2(n11296), .ZN(n11297) );
  AOI211_X1 U13196 ( .C1(n16336), .C2(n11299), .A(n11298), .B(n11297), .ZN(
        n11300) );
  OAI21_X1 U13197 ( .B1(n11301), .B2(n16327), .A(n11300), .ZN(P3_U3186) );
  OAI21_X1 U13198 ( .B1(n11303), .B2(n13018), .A(n11302), .ZN(n16423) );
  INV_X1 U13199 ( .A(n16423), .ZN(n11312) );
  NAND2_X1 U13200 ( .A1(n13060), .A2(n12855), .ZN(n11595) );
  INV_X1 U13201 ( .A(n11595), .ZN(n16410) );
  NAND2_X1 U13202 ( .A1(n16411), .A2(n16410), .ZN(n13510) );
  OAI22_X1 U13203 ( .A1(n16373), .A2(n16374), .B1(n11650), .B2(n16372), .ZN(
        n11309) );
  INV_X1 U13204 ( .A(n11131), .ZN(n11305) );
  OAI21_X1 U13205 ( .B1(n11305), .B2(n11304), .A(n13018), .ZN(n11306) );
  AND3_X1 U13206 ( .A1(n11307), .A2(n16377), .A3(n11306), .ZN(n11308) );
  AOI211_X1 U13207 ( .C1(n13661), .C2(n16423), .A(n11309), .B(n11308), .ZN(
        n16425) );
  MUX2_X1 U13208 ( .A(n10969), .B(n16425), .S(n16411), .Z(n11311) );
  AOI22_X1 U13209 ( .A1(n13555), .A2(n16422), .B1(n16388), .B2(n15756), .ZN(
        n11310) );
  OAI211_X1 U13210 ( .C1(n11312), .C2(n13510), .A(n11311), .B(n11310), .ZN(
        P3_U3230) );
  NAND2_X1 U13211 ( .A1(n11313), .A2(n13739), .ZN(n11314) );
  OAI211_X1 U13212 ( .C1(n11315), .C2(n13745), .A(n11314), .B(n13066), .ZN(
        P3_U3272) );
  INV_X1 U13213 ( .A(n14691), .ZN(n16532) );
  XNOR2_X1 U13214 ( .A(n14249), .B(n11316), .ZN(n11452) );
  INV_X1 U13215 ( .A(n11452), .ZN(n11324) );
  NAND2_X1 U13216 ( .A1(n11656), .A2(n13951), .ZN(n11317) );
  NAND2_X1 U13217 ( .A1(n11317), .A2(n14594), .ZN(n11318) );
  NOR2_X1 U13218 ( .A1(n11333), .A2(n11318), .ZN(n11443) );
  OAI21_X1 U13219 ( .B1(n14249), .B2(n11320), .A(n11319), .ZN(n11321) );
  NAND2_X1 U13220 ( .A1(n11321), .A2(n7449), .ZN(n11322) );
  OAI211_X1 U13221 ( .C1(n11452), .C2(n8139), .A(n11323), .B(n11322), .ZN(
        n11447) );
  AOI211_X1 U13222 ( .C1(n16532), .C2(n11324), .A(n11443), .B(n11447), .ZN(
        n11658) );
  OAI22_X1 U13223 ( .A1(n14785), .A2(n13995), .B1(n12115), .B2(n10017), .ZN(
        n11325) );
  INV_X1 U13224 ( .A(n11325), .ZN(n11326) );
  OAI21_X1 U13225 ( .B1(n11658), .B2(n16585), .A(n11326), .ZN(P2_U3433) );
  XNOR2_X1 U13226 ( .A(n11327), .B(n14247), .ZN(n16415) );
  OAI21_X1 U13227 ( .B1(n11329), .B2(n14247), .A(n11328), .ZN(n11330) );
  AOI222_X1 U13228 ( .A1(n7449), .A2(n11330), .B1(n14321), .B2(n14613), .C1(
        n14319), .C2(n14614), .ZN(n16417) );
  MUX2_X1 U13229 ( .A(n11331), .B(n16417), .S(n14644), .Z(n11337) );
  OAI211_X1 U13230 ( .C1(n11333), .C2(n16418), .A(n14594), .B(n11332), .ZN(
        n16416) );
  OAI22_X1 U13231 ( .A1(n14553), .A2(n16416), .B1(n11334), .B2(n14641), .ZN(
        n11335) );
  AOI21_X1 U13232 ( .B1(n14646), .B2(n14005), .A(n11335), .ZN(n11336) );
  OAI211_X1 U13233 ( .C1(n14604), .C2(n16415), .A(n11337), .B(n11336), .ZN(
        P2_U3263) );
  INV_X1 U13234 ( .A(n11346), .ZN(n11339) );
  NAND2_X1 U13235 ( .A1(n11339), .A2(n11338), .ZN(n11340) );
  NAND2_X1 U13236 ( .A1(n11350), .A2(n11340), .ZN(n11344) );
  NAND2_X1 U13237 ( .A1(n11341), .A2(n11900), .ZN(n11343) );
  AOI22_X1 U13238 ( .A1(n16233), .A2(n10048), .B1(n10051), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n11342) );
  XNOR2_X1 U13239 ( .A(n14068), .B(n7463), .ZN(n11616) );
  NAND2_X1 U13240 ( .A1(n14312), .A2(n7458), .ZN(n11601) );
  XNOR2_X1 U13241 ( .A(n11616), .B(n11601), .ZN(n11345) );
  INV_X1 U13242 ( .A(n11345), .ZN(n11349) );
  NAND2_X1 U13243 ( .A1(n11346), .A2(n13977), .ZN(n11347) );
  OAI21_X1 U13244 ( .B1(n14062), .B2(n13967), .A(n11347), .ZN(n11348) );
  NAND3_X1 U13245 ( .A1(n11350), .A2(n11349), .A3(n11348), .ZN(n11365) );
  INV_X1 U13246 ( .A(n11506), .ZN(n11352) );
  NAND2_X1 U13247 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n16235)
         );
  INV_X1 U13248 ( .A(n16235), .ZN(n11351) );
  AOI21_X1 U13249 ( .B1(n13972), .B2(n11352), .A(n11351), .ZN(n11364) );
  NAND2_X1 U13250 ( .A1(n13902), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n11360) );
  INV_X1 U13251 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11353) );
  OR2_X1 U13252 ( .A1(n10986), .A2(n11353), .ZN(n11359) );
  NAND2_X1 U13253 ( .A1(n11355), .A2(n11354), .ZN(n11356) );
  NAND2_X1 U13254 ( .A1(n11608), .A2(n11356), .ZN(n11685) );
  OR2_X1 U13255 ( .A1(n10059), .A2(n11685), .ZN(n11358) );
  OR2_X1 U13256 ( .A1(n14192), .A2(n11686), .ZN(n11357) );
  NAND4_X1 U13257 ( .A1(n11360), .A2(n11359), .A3(n11358), .A4(n11357), .ZN(
        n14311) );
  INV_X1 U13258 ( .A(n14311), .ZN(n14077) );
  OAI22_X1 U13259 ( .A1(n14077), .A2(n13933), .B1(n13932), .B2(n14062), .ZN(
        n11361) );
  INV_X1 U13260 ( .A(n11361), .ZN(n11363) );
  NAND2_X1 U13261 ( .A1(n14068), .A2(n13952), .ZN(n11362) );
  NAND4_X1 U13262 ( .A1(n11365), .A2(n11364), .A3(n11363), .A4(n11362), .ZN(
        n11366) );
  AOI21_X1 U13263 ( .B1(n7602), .B2(n13977), .A(n11366), .ZN(n11367) );
  INV_X1 U13264 ( .A(n11367), .ZN(P2_U3189) );
  MUX2_X1 U13265 ( .A(n11369), .B(n11368), .S(n14644), .Z(n11374) );
  OAI22_X1 U13266 ( .A1(n14622), .A2(n7691), .B1(n14641), .B2(n11370), .ZN(
        n11371) );
  AOI21_X1 U13267 ( .B1(n11372), .B2(n14650), .A(n11371), .ZN(n11373) );
  OAI211_X1 U13268 ( .C1(n14604), .C2(n11375), .A(n11374), .B(n11373), .ZN(
        P2_U3259) );
  OAI21_X1 U13269 ( .B1(n11378), .B2(P1_REG1_REG_14__SCAN_IN), .A(n11376), 
        .ZN(n11569) );
  AOI21_X1 U13270 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n11377), .A(n11574), 
        .ZN(n11389) );
  INV_X1 U13271 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15958) );
  NAND2_X1 U13272 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14949)
         );
  OAI21_X1 U13273 ( .B1(n16364), .B2(n15958), .A(n14949), .ZN(n11387) );
  AND2_X1 U13274 ( .A1(n11378), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11379) );
  AOI21_X1 U13275 ( .B1(n11381), .B2(n11380), .A(n11379), .ZN(n11383) );
  NAND2_X1 U13276 ( .A1(n11383), .A2(n11382), .ZN(n11579) );
  OAI21_X1 U13277 ( .B1(n11383), .B2(n11382), .A(n11579), .ZN(n11384) );
  NOR2_X1 U13278 ( .A1(n11384), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11581) );
  AOI21_X1 U13279 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n11384), .A(n11581), 
        .ZN(n11385) );
  NOR2_X1 U13280 ( .A1(n11385), .A2(n16264), .ZN(n11386) );
  AOI211_X1 U13281 ( .C1(n15065), .C2(n11570), .A(n11387), .B(n11386), .ZN(
        n11388) );
  OAI21_X1 U13282 ( .B1(n11389), .B2(n16266), .A(n11388), .ZN(P1_U3258) );
  NAND2_X1 U13283 ( .A1(n11391), .A2(n11390), .ZN(n11392) );
  NAND2_X1 U13284 ( .A1(n11392), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n11393) );
  XNOR2_X1 U13285 ( .A(n11393), .B(P2_IR_REG_18__SCAN_IN), .ZN(n14349) );
  INV_X1 U13286 ( .A(n14349), .ZN(n14359) );
  INV_X1 U13287 ( .A(n12423), .ZN(n11396) );
  OAI222_X1 U13288 ( .A1(P2_U3088), .A2(n14359), .B1(n14816), .B2(n11396), 
        .C1(n11394), .C2(n14818), .ZN(P2_U3309) );
  INV_X1 U13289 ( .A(n15059), .ZN(n16267) );
  OAI222_X1 U13290 ( .A1(P1_U3086), .A2(n16267), .B1(n15919), .B2(n11396), 
        .C1(n11395), .C2(n15916), .ZN(P1_U3337) );
  XNOR2_X1 U13291 ( .A(n11398), .B(n11397), .ZN(n11399) );
  NAND2_X1 U13292 ( .A1(n11399), .A2(n13342), .ZN(n11417) );
  INV_X1 U13293 ( .A(n11400), .ZN(n11402) );
  NAND3_X1 U13294 ( .A1(n11403), .A2(n11402), .A3(n11401), .ZN(n11404) );
  AOI21_X1 U13295 ( .B1(n11405), .B2(n11404), .A(n13368), .ZN(n11415) );
  INV_X1 U13296 ( .A(n11406), .ZN(n11408) );
  NAND3_X1 U13297 ( .A1(n11409), .A2(n11408), .A3(n11407), .ZN(n11410) );
  AOI21_X1 U13298 ( .B1(n11411), .B2(n11410), .A(n16328), .ZN(n11414) );
  INV_X1 U13299 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n16001) );
  NOR2_X1 U13300 ( .A1(n13345), .A2(n16001), .ZN(n11413) );
  INV_X1 U13301 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n11412) );
  NOR2_X1 U13302 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11412), .ZN(n11700) );
  NOR4_X1 U13303 ( .A1(n11415), .A2(n11414), .A3(n11413), .A4(n11700), .ZN(
        n11416) );
  OAI211_X1 U13304 ( .C1(n16333), .C2(n11418), .A(n11417), .B(n11416), .ZN(
        P3_U3188) );
  NAND2_X1 U13305 ( .A1(n11431), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n11419) );
  INV_X1 U13306 ( .A(n11439), .ZN(n11839) );
  INV_X1 U13307 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n12039) );
  AOI21_X1 U13308 ( .B1(n11423), .B2(n12039), .A(n11836), .ZN(n11442) );
  OAI22_X1 U13309 ( .A1(n11426), .A2(n11425), .B1(n11424), .B2(n11431), .ZN(
        n11428) );
  MUX2_X1 U13310 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n13357), .Z(n11840) );
  XNOR2_X1 U13311 ( .A(n11840), .B(n11439), .ZN(n11427) );
  NAND2_X1 U13312 ( .A1(n11427), .A2(n11428), .ZN(n11841) );
  OAI21_X1 U13313 ( .B1(n11428), .B2(n11427), .A(n11841), .ZN(n11429) );
  NAND2_X1 U13314 ( .A1(n11429), .A2(n13342), .ZN(n11441) );
  NOR2_X1 U13315 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15782), .ZN(n12126) );
  INV_X1 U13316 ( .A(n12126), .ZN(n11430) );
  OAI21_X1 U13317 ( .B1(n13345), .B2(n15946), .A(n11430), .ZN(n11438) );
  NAND2_X1 U13318 ( .A1(n11431), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n11432) );
  INV_X1 U13319 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n16503) );
  AOI21_X1 U13320 ( .B1(n11435), .B2(n16503), .A(n11831), .ZN(n11436) );
  NOR2_X1 U13321 ( .A1(n11436), .A2(n16328), .ZN(n11437) );
  AOI211_X1 U13322 ( .C1(n13370), .C2(n11439), .A(n11438), .B(n11437), .ZN(
        n11440) );
  OAI211_X1 U13323 ( .C1(n11442), .C2(n13368), .A(n11441), .B(n11440), .ZN(
        P3_U3191) );
  INV_X1 U13324 ( .A(n11443), .ZN(n11445) );
  OAI22_X1 U13325 ( .A1(n14553), .A2(n11445), .B1(n11444), .B2(n14641), .ZN(
        n11446) );
  AOI21_X1 U13326 ( .B1(n14646), .B2(n11656), .A(n11446), .ZN(n11451) );
  INV_X1 U13327 ( .A(n11447), .ZN(n11448) );
  MUX2_X1 U13328 ( .A(n11449), .B(n11448), .S(n14644), .Z(n11450) );
  OAI211_X1 U13329 ( .C1(n11452), .C2(n14629), .A(n11451), .B(n11450), .ZN(
        P2_U3264) );
  INV_X1 U13330 ( .A(n11453), .ZN(n11456) );
  INV_X1 U13331 ( .A(n11454), .ZN(n11455) );
  NOR2_X1 U13332 ( .A1(n12377), .A2(n11742), .ZN(n11459) );
  AOI21_X1 U13333 ( .B1(n16478), .B2(n7456), .A(n11459), .ZN(n11660) );
  AOI22_X1 U13334 ( .A1(n16478), .A2(n12687), .B1(n7456), .B2(n14969), .ZN(
        n11460) );
  XNOR2_X1 U13335 ( .A(n11460), .B(n12705), .ZN(n11661) );
  XOR2_X1 U13336 ( .A(n11660), .B(n11661), .Z(n11664) );
  XNOR2_X1 U13337 ( .A(n11665), .B(n11664), .ZN(n11467) );
  INV_X1 U13338 ( .A(n14968), .ZN(n11822) );
  OAI21_X1 U13339 ( .B1(n14951), .B2(n11822), .A(n11461), .ZN(n11462) );
  AOI21_X1 U13340 ( .B1(n14955), .B2(n14970), .A(n11462), .ZN(n11463) );
  OAI21_X1 U13341 ( .B1(n14952), .B2(n11533), .A(n11463), .ZN(n11464) );
  AOI21_X1 U13342 ( .B1(n16478), .B2(n14844), .A(n11464), .ZN(n11465) );
  OAI21_X1 U13343 ( .B1(n11467), .B2(n11466), .A(n11465), .ZN(P1_U3213) );
  XNOR2_X1 U13344 ( .A(n11475), .B(n12834), .ZN(n11470) );
  NAND2_X1 U13345 ( .A1(n11470), .A2(n11650), .ZN(n11644) );
  OAI21_X1 U13346 ( .B1(n11470), .B2(n11650), .A(n11644), .ZN(n11471) );
  AOI21_X1 U13347 ( .B1(n11472), .B2(n11471), .A(n11647), .ZN(n11478) );
  AOI22_X1 U13348 ( .A1(n13196), .A2(n13223), .B1(n13185), .B2(n13225), .ZN(
        n11474) );
  OAI211_X1 U13349 ( .C1(n13199), .C2(n11475), .A(n11474), .B(n11473), .ZN(
        n11476) );
  AOI21_X1 U13350 ( .B1(n11596), .B2(n13202), .A(n11476), .ZN(n11477) );
  OAI21_X1 U13351 ( .B1(n11478), .B2(n13204), .A(n11477), .ZN(P3_U3170) );
  OAI22_X1 U13352 ( .A1(n14644), .A2(n11480), .B1(n11479), .B2(n14641), .ZN(
        n11483) );
  NOR2_X1 U13353 ( .A1(n14622), .A2(n11481), .ZN(n11482) );
  AOI211_X1 U13354 ( .C1(n11484), .C2(n14650), .A(n11483), .B(n11482), .ZN(
        n11487) );
  OR2_X1 U13355 ( .A1(n11485), .A2(n14604), .ZN(n11486) );
  OAI211_X1 U13356 ( .C1(n11488), .C2(n14571), .A(n11487), .B(n11486), .ZN(
        P2_U3260) );
  INV_X1 U13357 ( .A(n14044), .ZN(n11491) );
  INV_X1 U13358 ( .A(n11489), .ZN(n12754) );
  INV_X1 U13359 ( .A(n14641), .ZN(n14598) );
  AOI22_X1 U13360 ( .A1(n14571), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n12754), 
        .B2(n14598), .ZN(n11490) );
  OAI21_X1 U13361 ( .B1(n11491), .B2(n14622), .A(n11490), .ZN(n11494) );
  NOR2_X1 U13362 ( .A1(n11492), .A2(n14571), .ZN(n11493) );
  AOI211_X1 U13363 ( .C1(n11495), .C2(n14650), .A(n11494), .B(n11493), .ZN(
        n11496) );
  OAI21_X1 U13364 ( .B1(n14604), .B2(n11497), .A(n11496), .ZN(P2_U3258) );
  XNOR2_X1 U13365 ( .A(n14068), .B(n14312), .ZN(n14262) );
  NAND2_X1 U13366 ( .A1(n14060), .A2(n14313), .ZN(n11498) );
  XOR2_X1 U13367 ( .A(n11674), .B(n14262), .Z(n16527) );
  NOR2_X1 U13368 ( .A1(n14060), .A2(n14062), .ZN(n11500) );
  NAND2_X1 U13369 ( .A1(n14060), .A2(n14062), .ZN(n11502) );
  XNOR2_X1 U13370 ( .A(n11678), .B(n14262), .ZN(n11504) );
  OAI22_X1 U13371 ( .A1(n14077), .A2(n14374), .B1(n14062), .B2(n13941), .ZN(
        n11503) );
  AOI21_X1 U13372 ( .B1(n11504), .B2(n7449), .A(n11503), .ZN(n11505) );
  OAI21_X1 U13373 ( .B1(n16527), .B2(n8139), .A(n11505), .ZN(n16529) );
  NAND2_X1 U13374 ( .A1(n16529), .A2(n14644), .ZN(n11511) );
  OAI22_X1 U13375 ( .A1(n14644), .A2(n11507), .B1(n11506), .B2(n14641), .ZN(
        n11509) );
  OAI211_X1 U13376 ( .C1(n7988), .C2(n7989), .A(n14594), .B(n11683), .ZN(
        n16528) );
  NOR2_X1 U13377 ( .A1(n16528), .A2(n14553), .ZN(n11508) );
  AOI211_X1 U13378 ( .C1(n14646), .C2(n14068), .A(n11509), .B(n11508), .ZN(
        n11510) );
  OAI211_X1 U13379 ( .C1(n16527), .C2(n14629), .A(n11511), .B(n11510), .ZN(
        P2_U3255) );
  OR2_X1 U13380 ( .A1(n11512), .A2(n13015), .ZN(n11513) );
  NAND2_X1 U13381 ( .A1(n11514), .A2(n11513), .ZN(n16457) );
  NAND2_X1 U13382 ( .A1(n16457), .A2(n13661), .ZN(n11521) );
  NAND2_X1 U13383 ( .A1(n11515), .A2(n13015), .ZN(n11516) );
  NAND2_X1 U13384 ( .A1(n11806), .A2(n11516), .ZN(n11519) );
  NAND2_X1 U13385 ( .A1(n13222), .A2(n13498), .ZN(n11517) );
  OAI21_X1 U13386 ( .B1(n11650), .B2(n16374), .A(n11517), .ZN(n11518) );
  AOI21_X1 U13387 ( .B1(n11519), .B2(n16377), .A(n11518), .ZN(n11520) );
  AND2_X1 U13388 ( .A1(n11521), .A2(n11520), .ZN(n16459) );
  INV_X1 U13389 ( .A(n13510), .ZN(n16390) );
  AOI22_X1 U13390 ( .A1(n13555), .A2(n16456), .B1(n16388), .B2(n11643), .ZN(
        n11522) );
  OAI21_X1 U13391 ( .B1(n11523), .B2(n16411), .A(n11522), .ZN(n11524) );
  AOI21_X1 U13392 ( .B1(n16457), .B2(n16390), .A(n11524), .ZN(n11525) );
  OAI21_X1 U13393 ( .B1(n16459), .B2(n16414), .A(n11525), .ZN(P3_U3228) );
  OR2_X1 U13394 ( .A1(n11537), .A2(n14970), .ZN(n11526) );
  NAND2_X1 U13395 ( .A1(n11527), .A2(n11526), .ZN(n11529) );
  OR2_X1 U13396 ( .A1(n11529), .A2(n11540), .ZN(n11530) );
  NAND2_X1 U13397 ( .A1(n11733), .A2(n11530), .ZN(n16483) );
  NAND2_X1 U13398 ( .A1(n11531), .A2(n16478), .ZN(n11532) );
  NAND2_X1 U13399 ( .A1(n11737), .A2(n11532), .ZN(n16480) );
  INV_X1 U13400 ( .A(n15312), .ZN(n15341) );
  INV_X1 U13401 ( .A(n11533), .ZN(n11534) );
  AOI22_X1 U13402 ( .A1(n15343), .A2(n16478), .B1(n15341), .B2(n11534), .ZN(
        n11535) );
  OAI21_X1 U13403 ( .B1(n15221), .B2(n16480), .A(n11535), .ZN(n11547) );
  NAND2_X1 U13404 ( .A1(n11537), .A2(n11536), .ZN(n11538) );
  NAND2_X1 U13405 ( .A1(n11541), .A2(n11540), .ZN(n11542) );
  NAND3_X1 U13406 ( .A1(n11744), .A2(n15431), .A3(n11542), .ZN(n11545) );
  AOI22_X1 U13407 ( .A1(n15331), .A2(n14970), .B1(n14968), .B2(n15329), .ZN(
        n11544) );
  NAND2_X1 U13408 ( .A1(n16483), .A2(n15166), .ZN(n11543) );
  NAND3_X1 U13409 ( .A1(n11545), .A2(n11544), .A3(n11543), .ZN(n16481) );
  MUX2_X1 U13410 ( .A(n16481), .B(P1_REG2_REG_7__SCAN_IN), .S(n15295), .Z(
        n11546) );
  AOI211_X1 U13411 ( .C1(n15345), .C2(n16483), .A(n11547), .B(n11546), .ZN(
        n11548) );
  INV_X1 U13412 ( .A(n11548), .ZN(P1_U3286) );
  INV_X1 U13413 ( .A(n12508), .ZN(n11568) );
  OAI222_X1 U13414 ( .A1(P1_U3086), .A2(n11549), .B1(n15919), .B2(n11568), 
        .C1(n8036), .C2(n15916), .ZN(P1_U3335) );
  AOI22_X1 U13415 ( .A1(n14571), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n11550), 
        .B2(n14598), .ZN(n11551) );
  OAI21_X1 U13416 ( .B1(n11552), .B2(n14622), .A(n11551), .ZN(n11555) );
  NOR2_X1 U13417 ( .A1(n11553), .A2(n14604), .ZN(n11554) );
  AOI211_X1 U13418 ( .C1(n11556), .C2(n14650), .A(n11555), .B(n11554), .ZN(
        n11557) );
  OAI21_X1 U13419 ( .B1(n14571), .B2(n11558), .A(n11557), .ZN(P2_U3257) );
  INV_X1 U13420 ( .A(n14060), .ZN(n11561) );
  AOI22_X1 U13421 ( .A1(n14571), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n11559), 
        .B2(n14598), .ZN(n11560) );
  OAI21_X1 U13422 ( .B1(n11561), .B2(n14622), .A(n11560), .ZN(n11564) );
  NOR2_X1 U13423 ( .A1(n11562), .A2(n14604), .ZN(n11563) );
  AOI211_X1 U13424 ( .C1(n11565), .C2(n14650), .A(n11564), .B(n11563), .ZN(
        n11566) );
  OAI21_X1 U13425 ( .B1(n14571), .B2(n11567), .A(n11566), .ZN(P2_U3256) );
  INV_X1 U13426 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n12509) );
  OAI222_X1 U13427 ( .A1(n14818), .A2(n12509), .B1(P2_U3088), .B2(n14282), 
        .C1(n14816), .C2(n11568), .ZN(P2_U3307) );
  INV_X1 U13428 ( .A(n11569), .ZN(n11571) );
  NOR2_X1 U13429 ( .A1(n11571), .A2(n11570), .ZN(n11573) );
  XNOR2_X1 U13430 ( .A(n11705), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11572) );
  NOR3_X1 U13431 ( .A1(n11574), .A2(n11573), .A3(n11572), .ZN(n11704) );
  INV_X1 U13432 ( .A(n11704), .ZN(n11576) );
  OAI21_X1 U13433 ( .B1(n11574), .B2(n11573), .A(n11572), .ZN(n11575) );
  NAND3_X1 U13434 ( .A1(n11576), .A2(n16354), .A3(n11575), .ZN(n11587) );
  NAND2_X1 U13435 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14879)
         );
  INV_X1 U13436 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11578) );
  NAND2_X1 U13437 ( .A1(n11705), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11707) );
  INV_X1 U13438 ( .A(n11707), .ZN(n11577) );
  AOI21_X1 U13439 ( .B1(n11578), .B2(n11588), .A(n11577), .ZN(n11583) );
  INV_X1 U13440 ( .A(n11579), .ZN(n11580) );
  NOR2_X1 U13441 ( .A1(n11581), .A2(n11580), .ZN(n11582) );
  NAND2_X1 U13442 ( .A1(n11582), .A2(n11583), .ZN(n11706) );
  OAI211_X1 U13443 ( .C1(n11583), .C2(n11582), .A(n16347), .B(n11706), .ZN(
        n11584) );
  NAND2_X1 U13444 ( .A1(n14879), .A2(n11584), .ZN(n11585) );
  AOI21_X1 U13445 ( .B1(n14978), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11585), 
        .ZN(n11586) );
  OAI211_X1 U13446 ( .C1(n16358), .C2(n11588), .A(n11587), .B(n11586), .ZN(
        P1_U3259) );
  XNOR2_X1 U13447 ( .A(n11589), .B(n13016), .ZN(n11592) );
  OAI22_X1 U13448 ( .A1(n11805), .A2(n16372), .B1(n11590), .B2(n16374), .ZN(
        n11591) );
  AOI21_X1 U13449 ( .B1(n11592), .B2(n16377), .A(n11591), .ZN(n16439) );
  OAI21_X1 U13450 ( .B1(n11594), .B2(n13016), .A(n11593), .ZN(n16438) );
  INV_X1 U13451 ( .A(n13661), .ZN(n16380) );
  AOI22_X1 U13452 ( .A1(n13555), .A2(n16437), .B1(n16388), .B2(n11596), .ZN(
        n11597) );
  OAI21_X1 U13453 ( .B1(n11598), .B2(n16411), .A(n11597), .ZN(n11599) );
  AOI21_X1 U13454 ( .B1(n16438), .B2(n13559), .A(n11599), .ZN(n11600) );
  OAI21_X1 U13455 ( .B1(n13492), .B2(n16439), .A(n11600), .ZN(P3_U3229) );
  INV_X1 U13456 ( .A(n11616), .ZN(n11602) );
  NAND2_X1 U13457 ( .A1(n11603), .A2(n11900), .ZN(n11605) );
  AOI22_X1 U13458 ( .A1(n16181), .A2(n10048), .B1(n7465), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n11604) );
  XNOR2_X1 U13459 ( .A(n14075), .B(n7463), .ZN(n12721) );
  NAND2_X1 U13460 ( .A1(n14311), .A2(n7458), .ZN(n11894) );
  XNOR2_X1 U13461 ( .A(n12721), .B(n11894), .ZN(n11617) );
  INV_X1 U13462 ( .A(n13933), .ZN(n13950) );
  NAND2_X1 U13463 ( .A1(n14181), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n11614) );
  INV_X1 U13464 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11797) );
  OR2_X1 U13465 ( .A1(n14192), .A2(n11797), .ZN(n11613) );
  INV_X1 U13466 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n11607) );
  NAND2_X1 U13467 ( .A1(n11608), .A2(n11607), .ZN(n11609) );
  NAND2_X1 U13468 ( .A1(n11785), .A2(n11609), .ZN(n12719) );
  OR2_X1 U13469 ( .A1(n10059), .A2(n12719), .ZN(n11612) );
  OR2_X1 U13470 ( .A1(n14191), .A2(n11610), .ZN(n11611) );
  NAND4_X1 U13471 ( .A1(n11614), .A2(n11613), .A3(n11612), .A4(n11611), .ZN(
        n14310) );
  AOI22_X1 U13472 ( .A1(n13950), .A2(n14310), .B1(n13888), .B2(n14312), .ZN(
        n11615) );
  NAND2_X1 U13473 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n16182)
         );
  OAI211_X1 U13474 ( .C1(n11685), .C2(n13943), .A(n11615), .B(n16182), .ZN(
        n11620) );
  AOI22_X1 U13475 ( .A1(n11616), .A2(n13977), .B1(n13957), .B2(n14312), .ZN(
        n11618) );
  NOR3_X1 U13476 ( .A1(n7602), .A2(n11618), .A3(n11617), .ZN(n11619) );
  AOI211_X1 U13477 ( .C1(n14075), .C2(n13952), .A(n11620), .B(n11619), .ZN(
        n11621) );
  OAI21_X1 U13478 ( .B1(n12720), .B2(n13915), .A(n11621), .ZN(P2_U3208) );
  INV_X1 U13479 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11787) );
  MUX2_X1 U13480 ( .A(n11787), .B(P2_REG1_REG_13__SCAN_IN), .S(n12275), .Z(
        n11624) );
  OAI21_X1 U13481 ( .B1(n11775), .B2(P2_REG1_REG_12__SCAN_IN), .A(n11622), 
        .ZN(n11623) );
  NOR2_X1 U13482 ( .A1(n11623), .A2(n11624), .ZN(n12270) );
  AOI211_X1 U13483 ( .C1(n11624), .C2(n11623), .A(n16228), .B(n12270), .ZN(
        n11634) );
  NAND2_X1 U13484 ( .A1(n12275), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11625) );
  OAI21_X1 U13485 ( .B1(n12275), .B2(P2_REG2_REG_13__SCAN_IN), .A(n11625), 
        .ZN(n11629) );
  OAI22_X1 U13486 ( .A1(n11627), .A2(n11626), .B1(n11775), .B2(
        P2_REG2_REG_12__SCAN_IN), .ZN(n11628) );
  NOR2_X1 U13487 ( .A1(n11628), .A2(n11629), .ZN(n12274) );
  AOI211_X1 U13488 ( .C1(n11629), .C2(n11628), .A(n16247), .B(n12274), .ZN(
        n11633) );
  NAND2_X1 U13489 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n11912)
         );
  NAND2_X1 U13490 ( .A1(n16097), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n11630) );
  OAI211_X1 U13491 ( .C1(n16189), .C2(n11631), .A(n11912), .B(n11630), .ZN(
        n11632) );
  OR3_X1 U13492 ( .A1(n11634), .A2(n11633), .A3(n11632), .ZN(P2_U3227) );
  INV_X1 U13493 ( .A(n11635), .ZN(n11642) );
  INV_X1 U13494 ( .A(n14604), .ZN(n14640) );
  OAI22_X1 U13495 ( .A1(n14644), .A2(n11171), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14641), .ZN(n11636) );
  AOI21_X1 U13496 ( .B1(n14646), .B2(n14019), .A(n11636), .ZN(n11637) );
  OAI21_X1 U13497 ( .B1(n14553), .B2(n11638), .A(n11637), .ZN(n11639) );
  AOI21_X1 U13498 ( .B1(n14640), .B2(n11640), .A(n11639), .ZN(n11641) );
  OAI21_X1 U13499 ( .B1(n14571), .B2(n11642), .A(n11641), .ZN(P2_U3262) );
  INV_X1 U13500 ( .A(n11643), .ZN(n11655) );
  INV_X1 U13501 ( .A(n13202), .ZN(n12329) );
  INV_X1 U13502 ( .A(n11644), .ZN(n11646) );
  XNOR2_X1 U13503 ( .A(n12834), .B(n16456), .ZN(n11692) );
  XNOR2_X1 U13504 ( .A(n11692), .B(n11805), .ZN(n11645) );
  INV_X1 U13505 ( .A(n11696), .ZN(n11649) );
  NOR3_X1 U13506 ( .A1(n11647), .A2(n11646), .A3(n11645), .ZN(n11648) );
  OAI21_X1 U13507 ( .B1(n11649), .B2(n11648), .A(n13183), .ZN(n11654) );
  OAI22_X1 U13508 ( .A1(n13198), .A2(n11650), .B1(n12884), .B2(n13187), .ZN(
        n11651) );
  AOI211_X1 U13509 ( .C1(n16456), .C2(n13168), .A(n11652), .B(n11651), .ZN(
        n11653) );
  OAI211_X1 U13510 ( .C1(n11655), .C2(n12329), .A(n11654), .B(n11653), .ZN(
        P3_U3167) );
  INV_X1 U13511 ( .A(n14734), .ZN(n14742) );
  AOI22_X1 U13512 ( .A1(n14742), .A2(n11656), .B1(n16584), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n11657) );
  OAI21_X1 U13513 ( .B1(n11658), .B2(n16584), .A(n11657), .ZN(P2_U3500) );
  AOI22_X1 U13514 ( .A1(n11756), .A2(n7456), .B1(n12698), .B2(n14968), .ZN(
        n11715) );
  AOI22_X1 U13515 ( .A1(n11756), .A2(n12687), .B1(n7456), .B2(n14968), .ZN(
        n11659) );
  XNOR2_X1 U13516 ( .A(n11659), .B(n12705), .ZN(n11716) );
  XOR2_X1 U13517 ( .A(n11715), .B(n11716), .Z(n11667) );
  INV_X1 U13518 ( .A(n11660), .ZN(n11663) );
  INV_X1 U13519 ( .A(n11661), .ZN(n11662) );
  OAI21_X1 U13520 ( .B1(n11667), .B2(n11666), .A(n11722), .ZN(n11668) );
  NAND2_X1 U13521 ( .A1(n11668), .A2(n14947), .ZN(n11672) );
  INV_X1 U13522 ( .A(n14967), .ZN(n11763) );
  NAND2_X1 U13523 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n15004) );
  OAI21_X1 U13524 ( .B1(n14951), .B2(n11763), .A(n15004), .ZN(n11670) );
  NOR2_X1 U13525 ( .A1(n14952), .A2(n11739), .ZN(n11669) );
  AOI211_X1 U13526 ( .C1(n14955), .C2(n14969), .A(n11670), .B(n11669), .ZN(
        n11671) );
  OAI211_X1 U13527 ( .C1(n8004), .C2(n14958), .A(n11672), .B(n11671), .ZN(
        P1_U3221) );
  NAND2_X1 U13528 ( .A1(n14075), .A2(n14077), .ZN(n11780) );
  OR2_X1 U13529 ( .A1(n14075), .A2(n14077), .ZN(n11673) );
  NAND2_X1 U13530 ( .A1(n11780), .A2(n11673), .ZN(n14261) );
  OAI21_X1 U13531 ( .B1(n11674), .B2(n14068), .A(n14312), .ZN(n11676) );
  NAND2_X1 U13532 ( .A1(n11674), .A2(n14068), .ZN(n11675) );
  XOR2_X1 U13533 ( .A(n14261), .B(n11772), .Z(n11889) );
  INV_X1 U13534 ( .A(n11889), .ZN(n11691) );
  INV_X1 U13535 ( .A(n14312), .ZN(n11682) );
  AND2_X1 U13536 ( .A1(n14068), .A2(n11682), .ZN(n11677) );
  INV_X1 U13537 ( .A(n11781), .ZN(n11679) );
  AOI21_X1 U13538 ( .B1(n14261), .B2(n11680), .A(n11679), .ZN(n11681) );
  OAI222_X1 U13539 ( .A1(n13941), .A2(n11682), .B1(n14374), .B2(n11938), .C1(
        n14591), .C2(n11681), .ZN(n11887) );
  NAND2_X1 U13540 ( .A1(n11887), .A2(n14644), .ZN(n11690) );
  AOI211_X1 U13541 ( .C1(n14075), .C2(n11683), .A(n7458), .B(n11796), .ZN(
        n11888) );
  INV_X1 U13542 ( .A(n14075), .ZN(n11684) );
  NOR2_X1 U13543 ( .A1(n11684), .A2(n14622), .ZN(n11688) );
  OAI22_X1 U13544 ( .A1(n14644), .A2(n11686), .B1(n11685), .B2(n14641), .ZN(
        n11687) );
  AOI211_X1 U13545 ( .C1(n11888), .C2(n14650), .A(n11688), .B(n11687), .ZN(
        n11689) );
  OAI211_X1 U13546 ( .C1(n14604), .C2(n11691), .A(n11690), .B(n11689), .ZN(
        P2_U3254) );
  INV_X1 U13547 ( .A(n11813), .ZN(n11703) );
  INV_X1 U13548 ( .A(n11692), .ZN(n11693) );
  NAND2_X1 U13549 ( .A1(n11693), .A2(n11805), .ZN(n11694) );
  AND2_X1 U13550 ( .A1(n11696), .A2(n11694), .ZN(n11698) );
  XNOR2_X1 U13551 ( .A(n12834), .B(n16470), .ZN(n11878) );
  XNOR2_X1 U13552 ( .A(n11878), .B(n12884), .ZN(n11697) );
  OAI211_X1 U13553 ( .C1(n11698), .C2(n11697), .A(n13183), .B(n11880), .ZN(
        n11702) );
  OAI22_X1 U13554 ( .A1(n13198), .A2(n11805), .B1(n12892), .B2(n13187), .ZN(
        n11699) );
  AOI211_X1 U13555 ( .C1(n16470), .C2(n13168), .A(n11700), .B(n11699), .ZN(
        n11701) );
  OAI211_X1 U13556 ( .C1(n11703), .C2(n12329), .A(n11702), .B(n11701), .ZN(
        P3_U3179) );
  AOI21_X1 U13557 ( .B1(n11705), .B2(P1_REG1_REG_16__SCAN_IN), .A(n11704), 
        .ZN(n15050) );
  XNOR2_X1 U13558 ( .A(n11708), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n15049) );
  XNOR2_X1 U13559 ( .A(n15050), .B(n15049), .ZN(n11714) );
  NAND2_X1 U13560 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14889)
         );
  NAND2_X1 U13561 ( .A1(n11707), .A2(n11706), .ZN(n15053) );
  XNOR2_X1 U13562 ( .A(n11708), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n15056) );
  XNOR2_X1 U13563 ( .A(n15053), .B(n15056), .ZN(n11709) );
  NAND2_X1 U13564 ( .A1(n16347), .A2(n11709), .ZN(n11710) );
  NAND2_X1 U13565 ( .A1(n14889), .A2(n11710), .ZN(n11712) );
  NOR2_X1 U13566 ( .A1(n16358), .A2(n15055), .ZN(n11711) );
  AOI211_X1 U13567 ( .C1(n14978), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n11712), 
        .B(n11711), .ZN(n11713) );
  OAI21_X1 U13568 ( .B1(n11714), .B2(n16266), .A(n11713), .ZN(P1_U3260) );
  INV_X1 U13569 ( .A(n11818), .ZN(n16508) );
  NAND2_X1 U13570 ( .A1(n11716), .A2(n11715), .ZN(n11721) );
  AND2_X1 U13571 ( .A1(n11722), .A2(n11721), .ZN(n11724) );
  NAND2_X1 U13572 ( .A1(n11818), .A2(n12687), .ZN(n11718) );
  NAND2_X1 U13573 ( .A1(n7456), .A2(n14967), .ZN(n11717) );
  NAND2_X1 U13574 ( .A1(n11718), .A2(n11717), .ZN(n11719) );
  XNOR2_X1 U13575 ( .A(n11719), .B(n12705), .ZN(n11964) );
  NOR2_X1 U13576 ( .A1(n12377), .A2(n11763), .ZN(n11720) );
  AOI21_X1 U13577 ( .B1(n11818), .B2(n7456), .A(n11720), .ZN(n11965) );
  XNOR2_X1 U13578 ( .A(n11964), .B(n11965), .ZN(n11723) );
  OAI211_X1 U13579 ( .C1(n11724), .C2(n11723), .A(n14947), .B(n11969), .ZN(
        n11728) );
  NAND2_X1 U13580 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n15021) );
  OAI21_X1 U13581 ( .B1(n14951), .B2(n11961), .A(n15021), .ZN(n11726) );
  NOR2_X1 U13582 ( .A1(n14952), .A2(n11819), .ZN(n11725) );
  AOI211_X1 U13583 ( .C1(n14955), .C2(n14968), .A(n11726), .B(n11725), .ZN(
        n11727) );
  OAI211_X1 U13584 ( .C1(n16508), .C2(n14958), .A(n11728), .B(n11727), .ZN(
        P1_U3231) );
  INV_X1 U13585 ( .A(n13777), .ZN(n11730) );
  OAI222_X1 U13586 ( .A1(n14818), .A2(n13778), .B1(n14816), .B2(n11730), .C1(
        n14287), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI222_X1 U13587 ( .A1(n11731), .A2(P1_U3086), .B1(n15919), .B2(n11730), 
        .C1(n11729), .C2(n15916), .ZN(P1_U3334) );
  OR2_X1 U13588 ( .A1(n16478), .A2(n14969), .ZN(n11732) );
  INV_X1 U13589 ( .A(n11745), .ZN(n11734) );
  OR2_X1 U13590 ( .A1(n11735), .A2(n11734), .ZN(n11736) );
  NAND2_X1 U13591 ( .A1(n11753), .A2(n11736), .ZN(n16494) );
  NAND2_X1 U13592 ( .A1(n11737), .A2(n11756), .ZN(n11738) );
  NAND2_X1 U13593 ( .A1(n11817), .A2(n11738), .ZN(n16491) );
  INV_X1 U13594 ( .A(n11739), .ZN(n11740) );
  AOI22_X1 U13595 ( .A1(n15343), .A2(n11756), .B1(n15341), .B2(n11740), .ZN(
        n11741) );
  OAI21_X1 U13596 ( .B1(n15221), .B2(n16491), .A(n11741), .ZN(n11751) );
  OR2_X1 U13597 ( .A1(n16478), .A2(n11742), .ZN(n11743) );
  OAI211_X1 U13598 ( .C1(n11746), .C2(n11745), .A(n11758), .B(n15431), .ZN(
        n11749) );
  AOI22_X1 U13599 ( .A1(n15331), .A2(n14969), .B1(n14967), .B2(n15329), .ZN(
        n11748) );
  NAND2_X1 U13600 ( .A1(n16494), .A2(n15166), .ZN(n11747) );
  NAND3_X1 U13601 ( .A1(n11749), .A2(n11748), .A3(n11747), .ZN(n16492) );
  MUX2_X1 U13602 ( .A(n16492), .B(P1_REG2_REG_8__SCAN_IN), .S(n15295), .Z(
        n11750) );
  AOI211_X1 U13603 ( .C1(n15345), .C2(n16494), .A(n11751), .B(n11750), .ZN(
        n11752) );
  INV_X1 U13604 ( .A(n11752), .ZN(P1_U3285) );
  INV_X1 U13605 ( .A(n11820), .ZN(n11826) );
  OR2_X1 U13606 ( .A1(n11818), .A2(n14967), .ZN(n11754) );
  NAND2_X1 U13607 ( .A1(n11825), .A2(n11754), .ZN(n11755) );
  NAND2_X1 U13608 ( .A1(n11755), .A2(n11762), .ZN(n11861) );
  OAI21_X1 U13609 ( .B1(n11755), .B2(n11762), .A(n11861), .ZN(n16524) );
  INV_X1 U13610 ( .A(n16524), .ZN(n11771) );
  OR2_X1 U13611 ( .A1(n11756), .A2(n11822), .ZN(n11757) );
  NAND2_X1 U13612 ( .A1(n11818), .A2(n11763), .ZN(n11759) );
  NAND2_X1 U13613 ( .A1(n11821), .A2(n11759), .ZN(n11761) );
  OR2_X1 U13614 ( .A1(n11818), .A2(n11763), .ZN(n11760) );
  NAND2_X1 U13615 ( .A1(n11761), .A2(n11760), .ZN(n11854) );
  INV_X1 U13616 ( .A(n11762), .ZN(n11853) );
  XNOR2_X1 U13617 ( .A(n11854), .B(n11853), .ZN(n11764) );
  OAI22_X1 U13618 ( .A1(n11764), .A2(n16449), .B1(n11763), .B2(n15230), .ZN(
        n16522) );
  XNOR2_X1 U13619 ( .A(n11864), .B(n11963), .ZN(n11765) );
  AOI22_X1 U13620 ( .A1(n11765), .A2(n15471), .B1(n15329), .B2(n14965), .ZN(
        n16520) );
  OAI22_X1 U13621 ( .A1(n11771), .A2(n15361), .B1(n15185), .B2(n16520), .ZN(
        n11766) );
  OAI21_X1 U13622 ( .B1(n16522), .B2(n11766), .A(n15338), .ZN(n11770) );
  OAI22_X1 U13623 ( .A1(n15338), .A2(n11767), .B1(n11972), .B2(n15312), .ZN(
        n11768) );
  AOI21_X1 U13624 ( .B1(n15343), .B2(n11963), .A(n11768), .ZN(n11769) );
  OAI211_X1 U13625 ( .C1(n11771), .C2(n15177), .A(n11770), .B(n11769), .ZN(
        P1_U3283) );
  OR2_X1 U13626 ( .A1(n14075), .A2(n14311), .ZN(n11773) );
  NAND2_X1 U13627 ( .A1(n11774), .A2(n11900), .ZN(n11777) );
  AOI22_X1 U13628 ( .A1(n11775), .A2(n10048), .B1(n10051), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n11776) );
  NAND2_X1 U13629 ( .A1(n14084), .A2(n11938), .ZN(n11943) );
  OR2_X1 U13630 ( .A1(n14084), .A2(n11938), .ZN(n11778) );
  INV_X1 U13631 ( .A(n14264), .ZN(n11779) );
  XNOR2_X1 U13632 ( .A(n11940), .B(n11779), .ZN(n16570) );
  INV_X1 U13633 ( .A(n16570), .ZN(n11802) );
  OAI21_X1 U13634 ( .B1(n14264), .B2(n7721), .A(n11944), .ZN(n11783) );
  NAND2_X1 U13635 ( .A1(n11783), .A2(n7449), .ZN(n11795) );
  INV_X1 U13636 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11784) );
  NAND2_X1 U13637 ( .A1(n11785), .A2(n11784), .ZN(n11786) );
  AND2_X1 U13638 ( .A1(n11905), .A2(n11786), .ZN(n11950) );
  NAND2_X1 U13639 ( .A1(n13843), .A2(n11950), .ZN(n11793) );
  OR2_X1 U13640 ( .A1(n14191), .A2(n11787), .ZN(n11792) );
  INV_X1 U13641 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11788) );
  OR2_X1 U13642 ( .A1(n10986), .A2(n11788), .ZN(n11791) );
  INV_X1 U13643 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11789) );
  OR2_X1 U13644 ( .A1(n14192), .A2(n11789), .ZN(n11790) );
  NAND4_X1 U13645 ( .A1(n11793), .A2(n11792), .A3(n11791), .A4(n11790), .ZN(
        n14309) );
  AOI22_X1 U13646 ( .A1(n14614), .A2(n14309), .B1(n14311), .B2(n14613), .ZN(
        n11794) );
  NAND2_X1 U13647 ( .A1(n11795), .A2(n11794), .ZN(n16575) );
  OAI211_X1 U13648 ( .C1(n16572), .C2(n11796), .A(n14594), .B(n11949), .ZN(
        n16571) );
  OAI22_X1 U13649 ( .A1(n14644), .A2(n11797), .B1(n12719), .B2(n14641), .ZN(
        n11798) );
  AOI21_X1 U13650 ( .B1(n14084), .B2(n14646), .A(n11798), .ZN(n11799) );
  OAI21_X1 U13651 ( .B1(n16571), .B2(n14553), .A(n11799), .ZN(n11800) );
  AOI21_X1 U13652 ( .B1(n16575), .B2(n14644), .A(n11800), .ZN(n11801) );
  OAI21_X1 U13653 ( .B1(n11802), .B2(n14604), .A(n11801), .ZN(P2_U3253) );
  OAI21_X1 U13654 ( .B1(n11804), .B2(n13023), .A(n11803), .ZN(n16472) );
  INV_X1 U13655 ( .A(n16472), .ZN(n11816) );
  OAI22_X1 U13656 ( .A1(n12892), .A2(n16372), .B1(n11805), .B2(n16374), .ZN(
        n11812) );
  INV_X1 U13657 ( .A(n11806), .ZN(n11808) );
  OAI21_X1 U13658 ( .B1(n11808), .B2(n11807), .A(n13023), .ZN(n11810) );
  AND3_X1 U13659 ( .A1(n11810), .A2(n16377), .A3(n11809), .ZN(n11811) );
  AOI211_X1 U13660 ( .C1(n13661), .C2(n16472), .A(n11812), .B(n11811), .ZN(
        n16474) );
  MUX2_X1 U13661 ( .A(n11039), .B(n16474), .S(n16411), .Z(n11815) );
  AOI22_X1 U13662 ( .A1(n13555), .A2(n16470), .B1(n16388), .B2(n11813), .ZN(
        n11814) );
  OAI211_X1 U13663 ( .C1(n11816), .C2(n13510), .A(n11815), .B(n11814), .ZN(
        P3_U3227) );
  INV_X1 U13664 ( .A(n15471), .ZN(n16544) );
  AOI211_X1 U13665 ( .C1(n11818), .C2(n11817), .A(n16544), .B(n11864), .ZN(
        n16506) );
  NOR2_X1 U13666 ( .A1(n15312), .A2(n11819), .ZN(n11824) );
  XNOR2_X1 U13667 ( .A(n11821), .B(n11820), .ZN(n11823) );
  OAI222_X1 U13668 ( .A1(n15232), .A2(n11961), .B1(n11823), .B2(n16449), .C1(
        n15230), .C2(n11822), .ZN(n16509) );
  AOI211_X1 U13669 ( .C1(n16506), .C2(n12592), .A(n11824), .B(n16509), .ZN(
        n11830) );
  OAI21_X1 U13670 ( .B1(n11827), .B2(n11826), .A(n11825), .ZN(n16511) );
  OAI22_X1 U13671 ( .A1(n15310), .A2(n16508), .B1(n10388), .B2(n15338), .ZN(
        n11828) );
  AOI21_X1 U13672 ( .B1(n16511), .B2(n15309), .A(n11828), .ZN(n11829) );
  OAI21_X1 U13673 ( .B1(n11830), .B2(n15333), .A(n11829), .ZN(P1_U3284) );
  NAND2_X1 U13674 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n12006), .ZN(n11832) );
  OAI21_X1 U13675 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(n12006), .A(n11832), 
        .ZN(n11833) );
  AOI21_X1 U13676 ( .B1(n11834), .B2(n11833), .A(n11992), .ZN(n11852) );
  NAND2_X1 U13677 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n12006), .ZN(n11835) );
  OAI21_X1 U13678 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n12006), .A(n11835), 
        .ZN(n11837) );
  AOI21_X1 U13679 ( .B1(n11837), .B2(n7485), .A(n12005), .ZN(n11848) );
  INV_X1 U13680 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11838) );
  NOR2_X1 U13681 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11838), .ZN(n12325) );
  AOI21_X1 U13682 ( .B1(n16330), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n12325), 
        .ZN(n11847) );
  MUX2_X1 U13683 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n13357), .Z(n11996) );
  XNOR2_X1 U13684 ( .A(n11996), .B(n11850), .ZN(n11844) );
  OR2_X1 U13685 ( .A1(n11840), .A2(n11839), .ZN(n11842) );
  NAND2_X1 U13686 ( .A1(n11842), .A2(n11841), .ZN(n11843) );
  NAND2_X1 U13687 ( .A1(n11844), .A2(n11843), .ZN(n11997) );
  OAI21_X1 U13688 ( .B1(n11844), .B2(n11843), .A(n11997), .ZN(n11845) );
  NAND2_X1 U13689 ( .A1(n13342), .A2(n11845), .ZN(n11846) );
  OAI211_X1 U13690 ( .C1(n13368), .C2(n11848), .A(n11847), .B(n11846), .ZN(
        n11849) );
  AOI21_X1 U13691 ( .B1(n11850), .B2(n13370), .A(n11849), .ZN(n11851) );
  OAI21_X1 U13692 ( .B1(n11852), .B2(n16328), .A(n11851), .ZN(P3_U3192) );
  NAND2_X1 U13693 ( .A1(n11854), .A2(n11853), .ZN(n11856) );
  OR2_X1 U13694 ( .A1(n11963), .A2(n11961), .ZN(n11855) );
  XNOR2_X1 U13695 ( .A(n12152), .B(n12150), .ZN(n11857) );
  NAND2_X1 U13696 ( .A1(n11857), .A2(n15431), .ZN(n11859) );
  AOI22_X1 U13697 ( .A1(n15331), .A2(n14966), .B1(n14963), .B2(n15329), .ZN(
        n11858) );
  AND2_X1 U13698 ( .A1(n11859), .A2(n11858), .ZN(n16550) );
  OR2_X1 U13699 ( .A1(n11963), .A2(n14966), .ZN(n11860) );
  NAND2_X1 U13700 ( .A1(n11861), .A2(n11860), .ZN(n11862) );
  NOR2_X1 U13701 ( .A1(n11862), .A2(n12150), .ZN(n11863) );
  OR2_X1 U13702 ( .A1(n12155), .A2(n11863), .ZN(n16548) );
  INV_X1 U13703 ( .A(n11963), .ZN(n16521) );
  NAND2_X1 U13704 ( .A1(n11865), .A2(n12153), .ZN(n11866) );
  NAND2_X1 U13705 ( .A1(n12162), .A2(n11866), .ZN(n16545) );
  OAI22_X1 U13706 ( .A1(n15338), .A2(n11867), .B1(n12065), .B2(n15312), .ZN(
        n11868) );
  AOI21_X1 U13707 ( .B1(n12153), .B2(n15343), .A(n11868), .ZN(n11869) );
  OAI21_X1 U13708 ( .B1(n16545), .B2(n15221), .A(n11869), .ZN(n11870) );
  AOI21_X1 U13709 ( .B1(n16548), .B2(n15309), .A(n11870), .ZN(n11871) );
  OAI21_X1 U13710 ( .B1(n16550), .B2(n15333), .A(n11871), .ZN(P1_U3282) );
  OAI21_X1 U13711 ( .B1(n11873), .B2(n12888), .A(n11872), .ZN(n11928) );
  INV_X1 U13712 ( .A(n11928), .ZN(n12046) );
  XNOR2_X1 U13713 ( .A(n11874), .B(n12888), .ZN(n11875) );
  AOI222_X1 U13714 ( .A1(n16377), .A2(n11875), .B1(n13222), .B2(n13500), .C1(
        n13220), .C2(n13498), .ZN(n11925) );
  MUX2_X1 U13715 ( .A(n11046), .B(n11925), .S(n16411), .Z(n11877) );
  AOI22_X1 U13716 ( .A1(n13555), .A2(n11924), .B1(n16388), .B2(n11883), .ZN(
        n11876) );
  OAI211_X1 U13717 ( .C1(n13590), .C2(n12046), .A(n11877), .B(n11876), .ZN(
        P3_U3226) );
  XNOR2_X1 U13718 ( .A(n7614), .B(n11924), .ZN(n11930) );
  XNOR2_X1 U13719 ( .A(n11930), .B(n12892), .ZN(n11931) );
  XNOR2_X1 U13720 ( .A(n11932), .B(n11931), .ZN(n11886) );
  OAI22_X1 U13721 ( .A1(n13198), .A2(n12884), .B1(n12124), .B2(n13187), .ZN(
        n11881) );
  AOI211_X1 U13722 ( .C1(n11924), .C2(n13168), .A(n11882), .B(n11881), .ZN(
        n11885) );
  NAND2_X1 U13723 ( .A1(n13202), .A2(n11883), .ZN(n11884) );
  OAI211_X1 U13724 ( .C1(n11886), .C2(n13204), .A(n11885), .B(n11884), .ZN(
        P3_U3153) );
  AOI211_X1 U13725 ( .C1(n11889), .C2(n16583), .A(n11888), .B(n11887), .ZN(
        n11893) );
  INV_X1 U13726 ( .A(n14785), .ZN(n14790) );
  NOR2_X1 U13727 ( .A1(n12115), .A2(n11353), .ZN(n11890) );
  AOI21_X1 U13728 ( .B1(n14075), .B2(n14790), .A(n11890), .ZN(n11891) );
  OAI21_X1 U13729 ( .B1(n11893), .B2(n16585), .A(n11891), .ZN(P2_U3463) );
  AOI22_X1 U13730 ( .A1(n14075), .A2(n14742), .B1(n16584), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11892) );
  OAI21_X1 U13731 ( .B1(n11893), .B2(n16584), .A(n11892), .ZN(P2_U3510) );
  INV_X1 U13732 ( .A(n12721), .ZN(n11895) );
  XNOR2_X1 U13733 ( .A(n14084), .B(n7463), .ZN(n11915) );
  NAND2_X1 U13734 ( .A1(n14310), .A2(n7458), .ZN(n11897) );
  XNOR2_X1 U13735 ( .A(n11915), .B(n11897), .ZN(n12722) );
  INV_X1 U13736 ( .A(n11915), .ZN(n11898) );
  NAND2_X1 U13737 ( .A1(n11898), .A2(n11897), .ZN(n11899) );
  NAND2_X1 U13738 ( .A1(n11901), .A2(n11900), .ZN(n11903) );
  AOI22_X1 U13739 ( .A1(n12275), .A2(n10048), .B1(n10051), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n11902) );
  XNOR2_X1 U13740 ( .A(n14089), .B(n7463), .ZN(n12732) );
  NAND2_X1 U13741 ( .A1(n14309), .A2(n7458), .ZN(n12085) );
  XNOR2_X1 U13742 ( .A(n12732), .B(n12085), .ZN(n11916) );
  INV_X1 U13743 ( .A(n11950), .ZN(n11914) );
  INV_X1 U13744 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11904) );
  NAND2_X1 U13745 ( .A1(n11905), .A2(n11904), .ZN(n11906) );
  NAND2_X1 U13746 ( .A1(n12020), .A2(n11906), .ZN(n12730) );
  INV_X1 U13747 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n12271) );
  OR2_X1 U13748 ( .A1(n14191), .A2(n12271), .ZN(n11909) );
  INV_X1 U13749 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n11907) );
  OR2_X1 U13750 ( .A1(n10986), .A2(n11907), .ZN(n11908) );
  AND2_X1 U13751 ( .A1(n11909), .A2(n11908), .ZN(n11911) );
  INV_X1 U13752 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n12028) );
  OR2_X1 U13753 ( .A1(n14192), .A2(n12028), .ZN(n11910) );
  OAI211_X1 U13754 ( .C1(n12730), .C2(n10059), .A(n11911), .B(n11910), .ZN(
        n14308) );
  AOI22_X1 U13755 ( .A1(n13888), .A2(n14310), .B1(n13950), .B2(n14308), .ZN(
        n11913) );
  OAI211_X1 U13756 ( .C1(n11914), .C2(n13943), .A(n11913), .B(n11912), .ZN(
        n11920) );
  INV_X1 U13757 ( .A(n12728), .ZN(n11918) );
  AOI22_X1 U13758 ( .A1(n11915), .A2(n13977), .B1(n13957), .B2(n14310), .ZN(
        n11917) );
  NOR3_X1 U13759 ( .A1(n11918), .A2(n11917), .A3(n11916), .ZN(n11919) );
  AOI211_X1 U13760 ( .C1(n14089), .C2(n13952), .A(n11920), .B(n11919), .ZN(
        n11921) );
  OAI21_X1 U13761 ( .B1(n12731), .B2(n13915), .A(n11921), .ZN(P2_U3206) );
  OAI222_X1 U13762 ( .A1(n13750), .A2(n11923), .B1(n13745), .B2(n15704), .C1(
        P3_U3151), .C2(n11922), .ZN(P3_U3270) );
  INV_X1 U13763 ( .A(n11924), .ZN(n12890) );
  OAI21_X1 U13764 ( .B1(n12890), .B2(n16558), .A(n11925), .ZN(n11926) );
  AOI21_X1 U13765 ( .B1(n13661), .B2(n11928), .A(n11926), .ZN(n12044) );
  AOI22_X1 U13766 ( .A1(n11928), .A2(n11927), .B1(P3_REG0_REG_7__SCAN_IN), 
        .B2(n16566), .ZN(n11929) );
  OAI21_X1 U13767 ( .B1(n12044), .B2(n16566), .A(n11929), .ZN(P3_U3411) );
  XNOR2_X1 U13768 ( .A(n7614), .B(n16485), .ZN(n12119) );
  XNOR2_X1 U13769 ( .A(n12119), .B(n12124), .ZN(n12120) );
  XNOR2_X1 U13770 ( .A(n12121), .B(n12120), .ZN(n11937) );
  OAI22_X1 U13771 ( .A1(n13198), .A2(n12892), .B1(n12323), .B2(n13187), .ZN(
        n11933) );
  AOI211_X1 U13772 ( .C1(n11984), .C2(n13168), .A(n11934), .B(n11933), .ZN(
        n11936) );
  NAND2_X1 U13773 ( .A1(n13202), .A2(n11983), .ZN(n11935) );
  OAI211_X1 U13774 ( .C1(n11937), .C2(n13204), .A(n11936), .B(n11935), .ZN(
        P3_U3161) );
  NOR2_X1 U13775 ( .A1(n14084), .A2(n14310), .ZN(n11939) );
  AOI21_X1 U13776 ( .B1(n14265), .B2(n11941), .A(n7599), .ZN(n12110) );
  AOI22_X1 U13777 ( .A1(n14308), .A2(n14614), .B1(n14310), .B2(n14613), .ZN(
        n11948) );
  INV_X1 U13778 ( .A(n11944), .ZN(n11942) );
  NOR3_X1 U13779 ( .A1(n11942), .A2(n8178), .A3(n14265), .ZN(n11946) );
  INV_X1 U13780 ( .A(n12013), .ZN(n11945) );
  OAI21_X1 U13781 ( .B1(n11946), .B2(n11945), .A(n7449), .ZN(n11947) );
  OAI211_X1 U13782 ( .C1(n12110), .C2(n8139), .A(n11948), .B(n11947), .ZN(
        n12111) );
  NAND2_X1 U13783 ( .A1(n12111), .A2(n14644), .ZN(n11955) );
  AOI211_X1 U13784 ( .C1(n14089), .C2(n11949), .A(n7458), .B(n7740), .ZN(
        n12112) );
  INV_X1 U13785 ( .A(n14089), .ZN(n11952) );
  AOI22_X1 U13786 ( .A1(n14571), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11950), 
        .B2(n14598), .ZN(n11951) );
  OAI21_X1 U13787 ( .B1(n11952), .B2(n14622), .A(n11951), .ZN(n11953) );
  AOI21_X1 U13788 ( .B1(n12112), .B2(n14650), .A(n11953), .ZN(n11954) );
  OAI211_X1 U13789 ( .C1(n12110), .C2(n14629), .A(n11955), .B(n11954), .ZN(
        P2_U3252) );
  XNOR2_X1 U13790 ( .A(n11957), .B(n11956), .ZN(n13786) );
  INV_X1 U13791 ( .A(n13786), .ZN(n11959) );
  OAI222_X1 U13792 ( .A1(n14818), .A2(n13787), .B1(n14816), .B2(n11959), .C1(
        n11958), .C2(P2_U3088), .ZN(P2_U3305) );
  OAI22_X1 U13793 ( .A1(n16521), .A2(n10644), .B1(n11961), .B2(n7468), .ZN(
        n11960) );
  XNOR2_X1 U13794 ( .A(n11960), .B(n12705), .ZN(n12059) );
  NOR2_X1 U13795 ( .A1(n12377), .A2(n11961), .ZN(n11962) );
  AOI21_X1 U13796 ( .B1(n11963), .B2(n7456), .A(n11962), .ZN(n12057) );
  XNOR2_X1 U13797 ( .A(n12059), .B(n12057), .ZN(n12060) );
  INV_X1 U13798 ( .A(n11964), .ZN(n11966) );
  XOR2_X1 U13799 ( .A(n12060), .B(n12061), .Z(n11970) );
  NAND2_X1 U13800 ( .A1(n11970), .A2(n14915), .ZN(n11976) );
  OAI21_X1 U13801 ( .B1(n14951), .B2(n12156), .A(n11971), .ZN(n11974) );
  NOR2_X1 U13802 ( .A1(n14952), .A2(n11972), .ZN(n11973) );
  AOI211_X1 U13803 ( .C1(n14955), .C2(n14967), .A(n11974), .B(n11973), .ZN(
        n11975) );
  OAI211_X1 U13804 ( .C1(n16521), .C2(n14958), .A(n11976), .B(n11975), .ZN(
        P1_U3217) );
  OAI21_X1 U13805 ( .B1(n11978), .B2(n13022), .A(n11977), .ZN(n16488) );
  INV_X1 U13806 ( .A(n16488), .ZN(n11989) );
  INV_X1 U13807 ( .A(n11979), .ZN(n11980) );
  AOI21_X1 U13808 ( .B1(n13022), .B2(n11981), .A(n11980), .ZN(n11982) );
  OAI222_X1 U13809 ( .A1(n16372), .A2(n12323), .B1(n16374), .B2(n12892), .C1(
        n13582), .C2(n11982), .ZN(n16486) );
  AOI22_X1 U13810 ( .A1(n13555), .A2(n11984), .B1(n16388), .B2(n11983), .ZN(
        n11985) );
  OAI21_X1 U13811 ( .B1(n11986), .B2(n16411), .A(n11985), .ZN(n11987) );
  AOI21_X1 U13812 ( .B1(n16486), .B2(n16411), .A(n11987), .ZN(n11988) );
  OAI21_X1 U13813 ( .B1(n11989), .B2(n13590), .A(n11988), .ZN(P3_U3225) );
  MUX2_X1 U13814 ( .A(n9105), .B(n11990), .S(P3_U3151), .Z(n11991) );
  INV_X1 U13815 ( .A(n11991), .ZN(P3_U3271) );
  INV_X1 U13816 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n16539) );
  AOI21_X1 U13817 ( .B1(n16539), .B2(n11993), .A(n7782), .ZN(n12012) );
  INV_X1 U13818 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11994) );
  MUX2_X1 U13819 ( .A(n11994), .B(n16539), .S(n13357), .Z(n12186) );
  XNOR2_X1 U13820 ( .A(n12186), .B(n11995), .ZN(n12000) );
  OR2_X1 U13821 ( .A1(n11996), .A2(n12006), .ZN(n11998) );
  NAND2_X1 U13822 ( .A1(n11998), .A2(n11997), .ZN(n11999) );
  NAND2_X1 U13823 ( .A1(n12000), .A2(n11999), .ZN(n12185) );
  OAI21_X1 U13824 ( .B1(n12000), .B2(n11999), .A(n12185), .ZN(n12001) );
  INV_X1 U13825 ( .A(n12001), .ZN(n12004) );
  AND2_X1 U13826 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n12418) );
  INV_X1 U13827 ( .A(n12418), .ZN(n12003) );
  NAND2_X1 U13828 ( .A1(n16330), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n12002) );
  OAI211_X1 U13829 ( .C1(n12004), .C2(n16327), .A(n12003), .B(n12002), .ZN(
        n12010) );
  XNOR2_X1 U13830 ( .A(n12195), .B(n12196), .ZN(n12007) );
  NOR2_X1 U13831 ( .A1(n11994), .A2(n12007), .ZN(n12197) );
  AOI21_X1 U13832 ( .B1(n12007), .B2(n11994), .A(n12197), .ZN(n12008) );
  NOR2_X1 U13833 ( .A1(n12008), .A2(n13368), .ZN(n12009) );
  AOI211_X1 U13834 ( .C1(n13370), .C2(n12196), .A(n12010), .B(n12009), .ZN(
        n12011) );
  OAI21_X1 U13835 ( .B1(n12012), .B2(n16328), .A(n12011), .ZN(P3_U3193) );
  INV_X1 U13836 ( .A(n14309), .ZN(n14091) );
  NAND2_X1 U13837 ( .A1(n12014), .A2(n14201), .ZN(n12016) );
  AOI22_X1 U13838 ( .A1(n12276), .A2(n10048), .B1(n10051), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n12015) );
  INV_X1 U13839 ( .A(n14308), .ZN(n12135) );
  XNOR2_X1 U13840 ( .A(n14102), .B(n12135), .ZN(n14267) );
  XNOR2_X1 U13841 ( .A(n12136), .B(n7939), .ZN(n12017) );
  NAND2_X1 U13842 ( .A1(n12017), .A2(n7449), .ZN(n12026) );
  INV_X1 U13843 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n12410) );
  INV_X1 U13844 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n12019) );
  NAND2_X1 U13845 ( .A1(n12020), .A2(n12019), .ZN(n12021) );
  NAND2_X1 U13846 ( .A1(n12096), .A2(n12021), .ZN(n12143) );
  OR2_X1 U13847 ( .A1(n12143), .A2(n10059), .ZN(n12024) );
  INV_X1 U13848 ( .A(n13846), .ZN(n12022) );
  AOI22_X1 U13849 ( .A1(n12022), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n14181), 
        .B2(P2_REG0_REG_15__SCAN_IN), .ZN(n12023) );
  OAI211_X1 U13850 ( .C1(n14191), .C2(n12410), .A(n12024), .B(n12023), .ZN(
        n14307) );
  AOI22_X1 U13851 ( .A1(n14307), .A2(n14614), .B1(n14613), .B2(n14309), .ZN(
        n12025) );
  NAND2_X1 U13852 ( .A1(n12026), .A2(n12025), .ZN(n16580) );
  INV_X1 U13853 ( .A(n16580), .ZN(n12033) );
  OAI21_X1 U13854 ( .B1(n12027), .B2(n14267), .A(n12133), .ZN(n16582) );
  OAI211_X1 U13855 ( .C1(n7739), .C2(n7740), .A(n14594), .B(n12142), .ZN(
        n16578) );
  OAI22_X1 U13856 ( .A1(n14644), .A2(n12028), .B1(n12730), .B2(n14641), .ZN(
        n12029) );
  AOI21_X1 U13857 ( .B1(n14102), .B2(n14646), .A(n12029), .ZN(n12030) );
  OAI21_X1 U13858 ( .B1(n16578), .B2(n14553), .A(n12030), .ZN(n12031) );
  AOI21_X1 U13859 ( .B1(n16582), .B2(n14640), .A(n12031), .ZN(n12032) );
  OAI21_X1 U13860 ( .B1(n12033), .B2(n14571), .A(n12032), .ZN(P2_U3251) );
  INV_X1 U13861 ( .A(n12077), .ZN(n12899) );
  XNOR2_X1 U13862 ( .A(n12245), .B(n13014), .ZN(n16500) );
  XNOR2_X1 U13863 ( .A(n12034), .B(n13014), .ZN(n12036) );
  AOI22_X1 U13864 ( .A1(n13218), .A2(n13498), .B1(n13500), .B2(n13220), .ZN(
        n12035) );
  OAI21_X1 U13865 ( .B1(n12036), .B2(n13582), .A(n12035), .ZN(n12037) );
  AOI21_X1 U13866 ( .B1(n16500), .B2(n13661), .A(n12037), .ZN(n16502) );
  AOI22_X1 U13867 ( .A1(n13555), .A2(n12127), .B1(n16388), .B2(n12128), .ZN(
        n12038) );
  OAI21_X1 U13868 ( .B1(n12039), .B2(n16411), .A(n12038), .ZN(n12040) );
  AOI21_X1 U13869 ( .B1(n16500), .B2(n16390), .A(n12040), .ZN(n12041) );
  OAI21_X1 U13870 ( .B1(n16502), .B2(n16414), .A(n12041), .ZN(P3_U3224) );
  OAI222_X1 U13871 ( .A1(n13750), .A2(n12043), .B1(n13745), .B2(n15502), .C1(
        P3_U3151), .C2(n12042), .ZN(P3_U3269) );
  MUX2_X1 U13872 ( .A(n11038), .B(n12044), .S(n16565), .Z(n12045) );
  OAI21_X1 U13873 ( .B1(n12046), .B2(n13664), .A(n12045), .ZN(P3_U3466) );
  INV_X1 U13874 ( .A(n13767), .ZN(n12049) );
  INV_X1 U13875 ( .A(n15916), .ZN(n15904) );
  AOI21_X1 U13876 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n15904), .A(n12047), 
        .ZN(n12048) );
  OAI21_X1 U13877 ( .B1(n12049), .B2(n15919), .A(n12048), .ZN(P1_U3332) );
  INV_X1 U13878 ( .A(n12153), .ZN(n16543) );
  NAND2_X1 U13879 ( .A1(n12153), .A2(n12687), .ZN(n12051) );
  NAND2_X1 U13880 ( .A1(n7456), .A2(n14965), .ZN(n12050) );
  NAND2_X1 U13881 ( .A1(n12051), .A2(n12050), .ZN(n12052) );
  XNOR2_X1 U13882 ( .A(n12052), .B(n12705), .ZN(n12056) );
  NAND2_X1 U13883 ( .A1(n12153), .A2(n7456), .ZN(n12054) );
  NAND2_X1 U13884 ( .A1(n12698), .A2(n14965), .ZN(n12053) );
  NAND2_X1 U13885 ( .A1(n12054), .A2(n12053), .ZN(n12055) );
  NOR2_X1 U13886 ( .A1(n12056), .A2(n12055), .ZN(n12171) );
  AOI21_X1 U13887 ( .B1(n12056), .B2(n12055), .A(n12171), .ZN(n12063) );
  INV_X1 U13888 ( .A(n12057), .ZN(n12058) );
  OAI21_X1 U13889 ( .B1(n12063), .B2(n12062), .A(n12173), .ZN(n12064) );
  NAND2_X1 U13890 ( .A1(n12064), .A2(n14947), .ZN(n12069) );
  NAND2_X1 U13891 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n15037)
         );
  OAI21_X1 U13892 ( .B1(n14951), .B2(n12312), .A(n15037), .ZN(n12067) );
  NOR2_X1 U13893 ( .A1(n14952), .A2(n12065), .ZN(n12066) );
  AOI211_X1 U13894 ( .C1(n14955), .C2(n14966), .A(n12067), .B(n12066), .ZN(
        n12068) );
  OAI211_X1 U13895 ( .C1(n16543), .C2(n14958), .A(n12069), .B(n12068), .ZN(
        P1_U3236) );
  INV_X1 U13896 ( .A(n14816), .ZN(n14801) );
  NAND2_X1 U13897 ( .A1(n13767), .A2(n14801), .ZN(n12071) );
  NAND2_X1 U13898 ( .A1(n12070), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14294) );
  OAI211_X1 U13899 ( .C1(n13768), .C2(n14818), .A(n12071), .B(n14294), .ZN(
        P2_U3304) );
  NAND2_X1 U13900 ( .A1(n12072), .A2(n9070), .ZN(n12073) );
  NAND3_X1 U13901 ( .A1(n12074), .A2(n16377), .A3(n12073), .ZN(n12076) );
  AOI22_X1 U13902 ( .A1(n13498), .A2(n13217), .B1(n13219), .B2(n13500), .ZN(
        n12075) );
  NAND2_X1 U13903 ( .A1(n12076), .A2(n12075), .ZN(n16514) );
  INV_X1 U13904 ( .A(n16514), .ZN(n12084) );
  OR2_X1 U13905 ( .A1(n12245), .A2(n12077), .ZN(n12078) );
  NAND2_X1 U13906 ( .A1(n12078), .A2(n12900), .ZN(n12079) );
  XNOR2_X1 U13907 ( .A(n12079), .B(n13024), .ZN(n16516) );
  NAND2_X1 U13908 ( .A1(n16516), .A2(n13559), .ZN(n12083) );
  INV_X1 U13909 ( .A(n12080), .ZN(n12330) );
  OAI22_X1 U13910 ( .A1(n13587), .A2(n16513), .B1(n12330), .B2(n16405), .ZN(
        n12081) );
  AOI21_X1 U13911 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n16414), .A(n12081), 
        .ZN(n12082) );
  OAI211_X1 U13912 ( .C1(n13492), .C2(n12084), .A(n12083), .B(n12082), .ZN(
        P3_U3223) );
  INV_X1 U13913 ( .A(n12732), .ZN(n12086) );
  XNOR2_X1 U13914 ( .A(n14102), .B(n7463), .ZN(n12103) );
  NAND2_X1 U13915 ( .A1(n14308), .A2(n7458), .ZN(n12087) );
  XNOR2_X1 U13916 ( .A(n12103), .B(n12087), .ZN(n12733) );
  INV_X1 U13917 ( .A(n12103), .ZN(n12088) );
  NAND2_X1 U13918 ( .A1(n12088), .A2(n12087), .ZN(n12089) );
  NAND2_X1 U13919 ( .A1(n12739), .A2(n12089), .ZN(n12095) );
  NAND2_X1 U13920 ( .A1(n12090), .A2(n14201), .ZN(n12094) );
  INV_X1 U13921 ( .A(n12092), .ZN(n12093) );
  XNOR2_X1 U13922 ( .A(n14108), .B(n7463), .ZN(n12349) );
  NAND2_X1 U13923 ( .A1(n14307), .A2(n7458), .ZN(n12350) );
  XNOR2_X1 U13924 ( .A(n12349), .B(n12350), .ZN(n12104) );
  INV_X1 U13925 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n12741) );
  NAND2_X1 U13926 ( .A1(n12096), .A2(n12741), .ZN(n12097) );
  NAND2_X1 U13927 ( .A1(n12223), .A2(n12097), .ZN(n12740) );
  AOI22_X1 U13928 ( .A1(n12022), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n14181), 
        .B2(P2_REG0_REG_16__SCAN_IN), .ZN(n12099) );
  NAND2_X1 U13929 ( .A1(n13902), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n12098) );
  OAI211_X1 U13930 ( .C1(n12740), .C2(n10059), .A(n12099), .B(n12098), .ZN(
        n14306) );
  AND2_X1 U13931 ( .A1(n14308), .A2(n14613), .ZN(n12100) );
  AOI21_X1 U13932 ( .B1(n14306), .B2(n14614), .A(n12100), .ZN(n12140) );
  INV_X1 U13933 ( .A(n12140), .ZN(n12101) );
  AOI22_X1 U13934 ( .A1(n13945), .A2(n12101), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12102) );
  OAI21_X1 U13935 ( .B1(n12143), .B2(n13943), .A(n12102), .ZN(n12108) );
  INV_X1 U13936 ( .A(n12739), .ZN(n12106) );
  AOI22_X1 U13937 ( .A1(n12103), .A2(n13977), .B1(n13957), .B2(n14308), .ZN(
        n12105) );
  NOR3_X1 U13938 ( .A1(n12106), .A2(n12105), .A3(n12104), .ZN(n12107) );
  AOI211_X1 U13939 ( .C1(n14108), .C2(n13952), .A(n12108), .B(n12107), .ZN(
        n12109) );
  OAI21_X1 U13940 ( .B1(n12750), .B2(n13915), .A(n12109), .ZN(P2_U3213) );
  INV_X1 U13941 ( .A(n12110), .ZN(n12113) );
  AOI211_X1 U13942 ( .C1(n16532), .C2(n12113), .A(n12112), .B(n12111), .ZN(
        n12118) );
  AOI22_X1 U13943 ( .A1(n14089), .A2(n14742), .B1(n16584), .B2(
        P2_REG1_REG_13__SCAN_IN), .ZN(n12114) );
  OAI21_X1 U13944 ( .B1(n12118), .B2(n16584), .A(n12114), .ZN(P2_U3512) );
  NOR2_X1 U13945 ( .A1(n12115), .A2(n11788), .ZN(n12116) );
  AOI21_X1 U13946 ( .B1(n14089), .B2(n14790), .A(n12116), .ZN(n12117) );
  OAI21_X1 U13947 ( .B1(n12118), .B2(n16585), .A(n12117), .ZN(P2_U3469) );
  XNOR2_X1 U13948 ( .A(n12834), .B(n12127), .ZN(n12319) );
  XNOR2_X1 U13949 ( .A(n12319), .B(n13219), .ZN(n12123) );
  AOI21_X1 U13950 ( .B1(n12123), .B2(n12122), .A(n12320), .ZN(n12131) );
  OAI22_X1 U13951 ( .A1(n13198), .A2(n12124), .B1(n12416), .B2(n13187), .ZN(
        n12125) );
  AOI211_X1 U13952 ( .C1(n12127), .C2(n13168), .A(n12126), .B(n12125), .ZN(
        n12130) );
  NAND2_X1 U13953 ( .A1(n13202), .A2(n12128), .ZN(n12129) );
  OAI211_X1 U13954 ( .C1(n12131), .C2(n13204), .A(n12130), .B(n12129), .ZN(
        P3_U3171) );
  OR2_X1 U13955 ( .A1(n14102), .A2(n14308), .ZN(n12132) );
  NAND2_X1 U13956 ( .A1(n12133), .A2(n12132), .ZN(n12134) );
  XNOR2_X1 U13957 ( .A(n14108), .B(n14307), .ZN(n14268) );
  NAND2_X1 U13958 ( .A1(n12134), .A2(n12139), .ZN(n12210) );
  OAI21_X1 U13959 ( .B1(n12134), .B2(n12139), .A(n12210), .ZN(n12406) );
  INV_X1 U13960 ( .A(n12406), .ZN(n12149) );
  NAND2_X1 U13961 ( .A1(n12136), .A2(n14102), .ZN(n12137) );
  OAI211_X1 U13962 ( .C1(n7469), .C2(n14268), .A(n7449), .B(n12219), .ZN(
        n12141) );
  NAND2_X1 U13963 ( .A1(n12141), .A2(n12140), .ZN(n12404) );
  NAND2_X1 U13964 ( .A1(n12404), .A2(n14644), .ZN(n12148) );
  AOI211_X1 U13965 ( .C1(n14108), .C2(n12142), .A(n7458), .B(n12232), .ZN(
        n12405) );
  INV_X1 U13966 ( .A(n14108), .ZN(n12412) );
  INV_X1 U13967 ( .A(n12143), .ZN(n12144) );
  AOI22_X1 U13968 ( .A1(n14571), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n12144), 
        .B2(n14598), .ZN(n12145) );
  OAI21_X1 U13969 ( .B1(n12412), .B2(n14622), .A(n12145), .ZN(n12146) );
  AOI21_X1 U13970 ( .B1(n12405), .B2(n14650), .A(n12146), .ZN(n12147) );
  OAI211_X1 U13971 ( .C1(n14604), .C2(n12149), .A(n12148), .B(n12147), .ZN(
        P2_U3250) );
  INV_X1 U13972 ( .A(n12150), .ZN(n12151) );
  OR2_X1 U13973 ( .A1(n12153), .A2(n12156), .ZN(n12154) );
  XNOR2_X1 U13974 ( .A(n12304), .B(n12157), .ZN(n12161) );
  INV_X1 U13975 ( .A(n12157), .ZN(n12303) );
  AOI21_X1 U13976 ( .B1(n12158), .B2(n12303), .A(n12310), .ZN(n15476) );
  AOI22_X1 U13977 ( .A1(n15331), .A2(n14965), .B1(n14962), .B2(n15329), .ZN(
        n12159) );
  OAI21_X1 U13978 ( .B1(n15476), .B2(n15361), .A(n12159), .ZN(n12160) );
  AOI21_X1 U13979 ( .B1(n12161), .B2(n15431), .A(n12160), .ZN(n15474) );
  AOI21_X1 U13980 ( .B1(n15470), .B2(n12162), .A(n12305), .ZN(n15472) );
  INV_X1 U13981 ( .A(n15470), .ZN(n12311) );
  INV_X1 U13982 ( .A(n12178), .ZN(n12163) );
  AOI22_X1 U13983 ( .A1(n15295), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n12163), 
        .B2(n15341), .ZN(n12164) );
  OAI21_X1 U13984 ( .B1(n12311), .B2(n15310), .A(n12164), .ZN(n12166) );
  NOR2_X1 U13985 ( .A1(n15476), .A2(n15177), .ZN(n12165) );
  AOI211_X1 U13986 ( .C1(n15472), .C2(n15347), .A(n12166), .B(n12165), .ZN(
        n12167) );
  OAI21_X1 U13987 ( .B1(n15295), .B2(n15474), .A(n12167), .ZN(P1_U3281) );
  NAND2_X1 U13988 ( .A1(n15470), .A2(n12687), .ZN(n12169) );
  NAND2_X1 U13989 ( .A1(n7456), .A2(n14963), .ZN(n12168) );
  NAND2_X1 U13990 ( .A1(n12169), .A2(n12168), .ZN(n12170) );
  XNOR2_X1 U13991 ( .A(n12170), .B(n12705), .ZN(n12251) );
  AOI22_X1 U13992 ( .A1(n15470), .A2(n7456), .B1(n12698), .B2(n14963), .ZN(
        n12252) );
  XNOR2_X1 U13993 ( .A(n12251), .B(n12252), .ZN(n12175) );
  INV_X1 U13994 ( .A(n12171), .ZN(n12172) );
  NAND2_X1 U13995 ( .A1(n12173), .A2(n12172), .ZN(n12174) );
  NAND2_X1 U13996 ( .A1(n12174), .A2(n12175), .ZN(n12258) );
  OAI21_X1 U13997 ( .B1(n12175), .B2(n12174), .A(n12258), .ZN(n12176) );
  NAND2_X1 U13998 ( .A1(n12176), .A2(n14947), .ZN(n12182) );
  INV_X1 U13999 ( .A(n14962), .ZN(n12338) );
  OAI21_X1 U14000 ( .B1(n14951), .B2(n12338), .A(n12177), .ZN(n12180) );
  NOR2_X1 U14001 ( .A1(n14952), .A2(n12178), .ZN(n12179) );
  AOI211_X1 U14002 ( .C1(n14955), .C2(n14965), .A(n12180), .B(n12179), .ZN(
        n12181) );
  OAI211_X1 U14003 ( .C1(n12311), .C2(n14958), .A(n12182), .B(n12181), .ZN(
        P1_U3224) );
  INV_X1 U14004 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n16564) );
  MUX2_X1 U14005 ( .A(n16564), .B(P3_REG1_REG_12__SCAN_IN), .S(n12294), .Z(
        n12188) );
  AOI21_X1 U14006 ( .B1(n12184), .B2(n12188), .A(n12293), .ZN(n12206) );
  INV_X1 U14007 ( .A(n12294), .ZN(n12204) );
  INV_X1 U14008 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12187) );
  MUX2_X1 U14009 ( .A(n12187), .B(P3_REG2_REG_12__SCAN_IN), .S(n12294), .Z(
        n12199) );
  MUX2_X1 U14010 ( .A(n12188), .B(n12199), .S(n12285), .Z(n12189) );
  INV_X1 U14011 ( .A(n12189), .ZN(n12190) );
  OAI211_X1 U14012 ( .C1(n12191), .C2(n12190), .A(n13342), .B(n12288), .ZN(
        n12194) );
  INV_X1 U14013 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n12192) );
  NOR2_X1 U14014 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12192), .ZN(n12545) );
  AOI21_X1 U14015 ( .B1(n16330), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12545), 
        .ZN(n12193) );
  NAND2_X1 U14016 ( .A1(n12194), .A2(n12193), .ZN(n12203) );
  NOR2_X1 U14017 ( .A1(n12196), .A2(n12195), .ZN(n12198) );
  NOR2_X1 U14018 ( .A1(n12198), .A2(n12197), .ZN(n12200) );
  AOI21_X1 U14019 ( .B1(n12200), .B2(n12199), .A(n12282), .ZN(n12201) );
  NOR2_X1 U14020 ( .A1(n12201), .A2(n13368), .ZN(n12202) );
  AOI211_X1 U14021 ( .C1(n13370), .C2(n12204), .A(n12203), .B(n12202), .ZN(
        n12205) );
  OAI21_X1 U14022 ( .B1(n12206), .B2(n16328), .A(n12205), .ZN(P3_U3194) );
  INV_X1 U14023 ( .A(n12207), .ZN(n12208) );
  OAI222_X1 U14024 ( .A1(P3_U3151), .A2(n13357), .B1(n13750), .B2(n12208), 
        .C1(n15700), .C2(n13745), .ZN(P3_U3268) );
  OR2_X1 U14025 ( .A1(n14108), .A2(n14307), .ZN(n12209) );
  NAND2_X1 U14026 ( .A1(n12211), .A2(n14201), .ZN(n12213) );
  AOI22_X1 U14027 ( .A1(n10051), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n10048), 
        .B2(n16207), .ZN(n12212) );
  INV_X1 U14028 ( .A(n14306), .ZN(n12214) );
  OR2_X1 U14029 ( .A1(n14789), .A2(n12214), .ZN(n14630) );
  NAND2_X1 U14030 ( .A1(n14789), .A2(n12214), .ZN(n12215) );
  NAND2_X1 U14031 ( .A1(n12216), .A2(n14270), .ZN(n12217) );
  NAND2_X1 U14032 ( .A1(n12451), .A2(n12217), .ZN(n14736) );
  INV_X1 U14033 ( .A(n14307), .ZN(n12746) );
  OR2_X1 U14034 ( .A1(n14108), .A2(n12746), .ZN(n12218) );
  OAI211_X1 U14035 ( .C1(n14270), .C2(n7723), .A(n14632), .B(n7449), .ZN(
        n12231) );
  INV_X1 U14036 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n12222) );
  NAND2_X1 U14037 ( .A1(n12223), .A2(n12222), .ZN(n12224) );
  NAND2_X1 U14038 ( .A1(n12357), .A2(n12224), .ZN(n14642) );
  OR2_X1 U14039 ( .A1(n14642), .A2(n10059), .ZN(n12229) );
  INV_X1 U14040 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n14643) );
  NAND2_X1 U14041 ( .A1(n14181), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n12226) );
  NAND2_X1 U14042 ( .A1(n13902), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n12225) );
  OAI211_X1 U14043 ( .C1(n14192), .C2(n14643), .A(n12226), .B(n12225), .ZN(
        n12227) );
  INV_X1 U14044 ( .A(n12227), .ZN(n12228) );
  NAND2_X1 U14045 ( .A1(n12229), .A2(n12228), .ZN(n14305) );
  AND2_X1 U14046 ( .A1(n14307), .A2(n14613), .ZN(n12230) );
  AOI21_X1 U14047 ( .B1(n14305), .B2(n14614), .A(n12230), .ZN(n12742) );
  NAND2_X1 U14048 ( .A1(n12231), .A2(n12742), .ZN(n14737) );
  NAND2_X1 U14049 ( .A1(n14737), .A2(n14644), .ZN(n12239) );
  INV_X1 U14050 ( .A(n14789), .ZN(n12235) );
  OR2_X1 U14051 ( .A1(n12235), .A2(n12232), .ZN(n12233) );
  AND3_X1 U14052 ( .A1(n14647), .A2(n12233), .A3(n14594), .ZN(n14738) );
  INV_X1 U14053 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n12234) );
  OAI22_X1 U14054 ( .A1(n14644), .A2(n12234), .B1(n12740), .B2(n14641), .ZN(
        n12237) );
  NOR2_X1 U14055 ( .A1(n12235), .A2(n14622), .ZN(n12236) );
  AOI211_X1 U14056 ( .C1(n14738), .C2(n14650), .A(n12237), .B(n12236), .ZN(
        n12238) );
  OAI211_X1 U14057 ( .C1(n14604), .C2(n14736), .A(n12239), .B(n12238), .ZN(
        P2_U3249) );
  XNOR2_X1 U14058 ( .A(n12240), .B(n12905), .ZN(n12241) );
  AOI222_X1 U14059 ( .A1(n16377), .A2(n12241), .B1(n13218), .B2(n13500), .C1(
        n13216), .C2(n13498), .ZN(n16535) );
  INV_X1 U14060 ( .A(n12419), .ZN(n12242) );
  OAI22_X1 U14061 ( .A1(n13587), .A2(n16536), .B1(n12242), .B2(n16405), .ZN(
        n12243) );
  AOI21_X1 U14062 ( .B1(n13492), .B2(P3_REG2_REG_11__SCAN_IN), .A(n12243), 
        .ZN(n12250) );
  OR2_X1 U14063 ( .A1(n12245), .A2(n12244), .ZN(n12247) );
  AND2_X1 U14064 ( .A1(n12247), .A2(n12246), .ZN(n12248) );
  XNOR2_X1 U14065 ( .A(n12248), .B(n12905), .ZN(n16538) );
  NAND2_X1 U14066 ( .A1(n16538), .A2(n13559), .ZN(n12249) );
  OAI211_X1 U14067 ( .C1(n16535), .C2(n16414), .A(n12250), .B(n12249), .ZN(
        P3_U3222) );
  INV_X1 U14068 ( .A(n12251), .ZN(n12253) );
  NAND2_X1 U14069 ( .A1(n12253), .A2(n12252), .ZN(n12256) );
  AND2_X1 U14070 ( .A1(n12258), .A2(n12256), .ZN(n12260) );
  OAI22_X1 U14071 ( .A1(n15462), .A2(n10644), .B1(n12338), .B2(n7468), .ZN(
        n12254) );
  XNOR2_X1 U14072 ( .A(n12254), .B(n12705), .ZN(n12381) );
  NOR2_X1 U14073 ( .A1(n12377), .A2(n12338), .ZN(n12255) );
  AOI21_X1 U14074 ( .B1(n12333), .B2(n7456), .A(n12255), .ZN(n12379) );
  XNOR2_X1 U14075 ( .A(n12381), .B(n12379), .ZN(n12259) );
  OAI211_X1 U14076 ( .C1(n12260), .C2(n12259), .A(n14947), .B(n12382), .ZN(
        n12267) );
  INV_X1 U14077 ( .A(n12307), .ZN(n12265) );
  NAND2_X1 U14078 ( .A1(n15332), .A2(n15329), .ZN(n12262) );
  NAND2_X1 U14079 ( .A1(n14963), .A2(n15331), .ZN(n12261) );
  AND2_X1 U14080 ( .A1(n12262), .A2(n12261), .ZN(n15461) );
  OAI21_X1 U14081 ( .B1(n14836), .B2(n15461), .A(n12263), .ZN(n12264) );
  AOI21_X1 U14082 ( .B1(n14893), .B2(n12265), .A(n12264), .ZN(n12266) );
  OAI211_X1 U14083 ( .C1(n15462), .C2(n14958), .A(n12267), .B(n12266), .ZN(
        P1_U3234) );
  NAND2_X1 U14084 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n12269)
         );
  NAND2_X1 U14085 ( .A1(n16097), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n12268) );
  OAI211_X1 U14086 ( .C1(n16189), .C2(n14345), .A(n12269), .B(n12268), .ZN(
        n12281) );
  AOI21_X1 U14087 ( .B1(n12275), .B2(P2_REG1_REG_13__SCAN_IN), .A(n12270), 
        .ZN(n16192) );
  MUX2_X1 U14088 ( .A(n12271), .B(P2_REG1_REG_14__SCAN_IN), .S(n12276), .Z(
        n16191) );
  NOR2_X1 U14089 ( .A1(n16192), .A2(n16191), .ZN(n16190) );
  XNOR2_X1 U14090 ( .A(n14345), .B(n14346), .ZN(n12272) );
  AOI211_X1 U14091 ( .C1(n12272), .C2(n12410), .A(n14347), .B(n16228), .ZN(
        n12280) );
  MUX2_X1 U14092 ( .A(n12028), .B(P2_REG2_REG_14__SCAN_IN), .S(n12276), .Z(
        n12273) );
  INV_X1 U14093 ( .A(n12273), .ZN(n16186) );
  AOI21_X1 U14094 ( .B1(n12275), .B2(P2_REG2_REG_13__SCAN_IN), .A(n12274), 
        .ZN(n16187) );
  NAND2_X1 U14095 ( .A1(n16186), .A2(n16187), .ZN(n16185) );
  OAI21_X1 U14096 ( .B1(n12276), .B2(P2_REG2_REG_14__SCAN_IN), .A(n16185), 
        .ZN(n14338) );
  XNOR2_X1 U14097 ( .A(n14345), .B(n14338), .ZN(n12278) );
  INV_X1 U14098 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n12277) );
  NOR2_X1 U14099 ( .A1(n12277), .A2(n12278), .ZN(n14339) );
  AOI211_X1 U14100 ( .C1(n12278), .C2(n12277), .A(n14339), .B(n16247), .ZN(
        n12279) );
  OR3_X1 U14101 ( .A1(n12281), .A2(n12280), .A3(n12279), .ZN(P2_U3229) );
  INV_X1 U14102 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12283) );
  AOI21_X1 U14103 ( .B1(n12284), .B2(n12283), .A(n13246), .ZN(n12302) );
  NAND2_X1 U14104 ( .A1(n12294), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12286) );
  MUX2_X1 U14105 ( .A(n7601), .B(n12286), .S(n12285), .Z(n12287) );
  MUX2_X1 U14106 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13357), .Z(n13235) );
  XNOR2_X1 U14107 ( .A(n13235), .B(n8029), .ZN(n12289) );
  NAND2_X1 U14108 ( .A1(n12290), .A2(n12289), .ZN(n13236) );
  OAI21_X1 U14109 ( .B1(n12290), .B2(n12289), .A(n13236), .ZN(n12300) );
  NAND2_X1 U14110 ( .A1(n13370), .A2(n8029), .ZN(n12292) );
  NOR2_X1 U14111 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8771), .ZN(n13155) );
  AOI21_X1 U14112 ( .B1(n16330), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n13155), 
        .ZN(n12291) );
  NAND2_X1 U14113 ( .A1(n12292), .A2(n12291), .ZN(n12299) );
  INV_X1 U14114 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12296) );
  AOI21_X1 U14115 ( .B1(n12296), .B2(n12295), .A(n7779), .ZN(n12297) );
  NOR2_X1 U14116 ( .A1(n12297), .A2(n16328), .ZN(n12298) );
  AOI211_X1 U14117 ( .C1(n13342), .C2(n12300), .A(n12299), .B(n12298), .ZN(
        n12301) );
  OAI21_X1 U14118 ( .B1(n12302), .B2(n13368), .A(n12301), .ZN(P3_U3195) );
  XNOR2_X1 U14119 ( .A(n12332), .B(n12331), .ZN(n15469) );
  NOR2_X1 U14120 ( .A1(n12305), .A2(n15462), .ZN(n12306) );
  NOR2_X1 U14121 ( .A1(n12306), .A2(n12343), .ZN(n15467) );
  OAI22_X1 U14122 ( .A1(n15295), .A2(n15461), .B1(n12307), .B2(n15312), .ZN(
        n12308) );
  AOI21_X1 U14123 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n15333), .A(n12308), 
        .ZN(n12309) );
  OAI21_X1 U14124 ( .B1(n15462), .B2(n15310), .A(n12309), .ZN(n12315) );
  NOR2_X1 U14125 ( .A1(n12313), .A2(n12331), .ZN(n12337) );
  AOI21_X1 U14126 ( .B1(n12313), .B2(n12331), .A(n12337), .ZN(n15464) );
  NOR2_X1 U14127 ( .A1(n15464), .A2(n15337), .ZN(n12314) );
  AOI211_X1 U14128 ( .C1(n15467), .C2(n15347), .A(n12315), .B(n12314), .ZN(
        n12316) );
  OAI21_X1 U14129 ( .B1(n15211), .B2(n15469), .A(n12316), .ZN(P1_U3280) );
  INV_X1 U14130 ( .A(n13812), .ZN(n12403) );
  AOI22_X1 U14131 ( .A1(n12317), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n15904), .ZN(n12318) );
  OAI21_X1 U14132 ( .B1(n12403), .B2(n15919), .A(n12318), .ZN(P1_U3331) );
  INV_X1 U14133 ( .A(n12319), .ZN(n12321) );
  XNOR2_X1 U14134 ( .A(n7614), .B(n12326), .ZN(n12413) );
  XNOR2_X1 U14135 ( .A(n12413), .B(n12416), .ZN(n12322) );
  OAI211_X1 U14136 ( .C1(n7610), .C2(n12322), .A(n12480), .B(n13183), .ZN(
        n12328) );
  OAI22_X1 U14137 ( .A1(n13198), .A2(n12323), .B1(n12920), .B2(n13187), .ZN(
        n12324) );
  AOI211_X1 U14138 ( .C1(n12326), .C2(n13168), .A(n12325), .B(n12324), .ZN(
        n12327) );
  OAI211_X1 U14139 ( .C1(n12330), .C2(n12329), .A(n12328), .B(n12327), .ZN(
        P3_U3157) );
  NAND2_X1 U14140 ( .A1(n12332), .A2(n12331), .ZN(n12335) );
  OR2_X1 U14141 ( .A1(n12333), .A2(n12338), .ZN(n12334) );
  XNOR2_X1 U14142 ( .A(n12553), .B(n12339), .ZN(n12336) );
  AOI222_X1 U14143 ( .A1(n14962), .A2(n15331), .B1(n15303), .B2(n15329), .C1(
        n15431), .C2(n12336), .ZN(n15459) );
  OAI21_X1 U14144 ( .B1(n12340), .B2(n12339), .A(n12572), .ZN(n15460) );
  OAI22_X1 U14145 ( .A1(n15338), .A2(n12341), .B1(n12387), .B2(n15312), .ZN(
        n12342) );
  AOI21_X1 U14146 ( .B1(n15456), .B2(n15343), .A(n12342), .ZN(n12346) );
  OR2_X1 U14147 ( .A1(n12574), .A2(n12343), .ZN(n12344) );
  AND2_X1 U14148 ( .A1(n15321), .A2(n12344), .ZN(n15457) );
  NAND2_X1 U14149 ( .A1(n15457), .A2(n15347), .ZN(n12345) );
  OAI211_X1 U14150 ( .C1(n15460), .C2(n15337), .A(n12346), .B(n12345), .ZN(
        n12347) );
  INV_X1 U14151 ( .A(n12347), .ZN(n12348) );
  OAI21_X1 U14152 ( .B1(n15295), .B2(n15459), .A(n12348), .ZN(P1_U3279) );
  INV_X1 U14153 ( .A(n12349), .ZN(n12747) );
  XNOR2_X1 U14154 ( .A(n14789), .B(n7463), .ZN(n12367) );
  NAND2_X1 U14155 ( .A1(n14306), .A2(n7458), .ZN(n12351) );
  XNOR2_X1 U14156 ( .A(n12367), .B(n12351), .ZN(n12745) );
  INV_X1 U14157 ( .A(n12367), .ZN(n12352) );
  NAND2_X1 U14158 ( .A1(n12352), .A2(n12351), .ZN(n12353) );
  NAND2_X1 U14159 ( .A1(n12354), .A2(n14201), .ZN(n12356) );
  AOI22_X1 U14160 ( .A1(n7465), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n10048), 
        .B2(n16218), .ZN(n12355) );
  XNOR2_X1 U14161 ( .A(n14728), .B(n7463), .ZN(n12426) );
  NAND2_X1 U14162 ( .A1(n14305), .A2(n7458), .ZN(n12427) );
  XNOR2_X1 U14163 ( .A(n12426), .B(n12427), .ZN(n12368) );
  INV_X1 U14164 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n12445) );
  NAND2_X1 U14165 ( .A1(n12357), .A2(n12445), .ZN(n12358) );
  NAND2_X1 U14166 ( .A1(n12439), .A2(n12358), .ZN(n12456) );
  OR2_X1 U14167 ( .A1(n12456), .A2(n10059), .ZN(n12363) );
  INV_X1 U14168 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n12457) );
  NAND2_X1 U14169 ( .A1(n13902), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n12360) );
  NAND2_X1 U14170 ( .A1(n14181), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n12359) );
  OAI211_X1 U14171 ( .C1(n12457), .C2(n14192), .A(n12360), .B(n12359), .ZN(
        n12361) );
  INV_X1 U14172 ( .A(n12361), .ZN(n12362) );
  NAND2_X1 U14173 ( .A1(n12363), .A2(n12362), .ZN(n14612) );
  AND2_X1 U14174 ( .A1(n14306), .A2(n14613), .ZN(n12364) );
  AOI21_X1 U14175 ( .B1(n14612), .B2(n14614), .A(n12364), .ZN(n14636) );
  INV_X1 U14176 ( .A(n14636), .ZN(n12365) );
  AOI22_X1 U14177 ( .A1(n13945), .A2(n12365), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12366) );
  OAI21_X1 U14178 ( .B1(n14642), .B2(n13943), .A(n12366), .ZN(n12372) );
  INV_X1 U14179 ( .A(n12753), .ZN(n12370) );
  AOI22_X1 U14180 ( .A1(n12367), .A2(n13977), .B1(n13957), .B2(n14306), .ZN(
        n12369) );
  NOR3_X1 U14181 ( .A1(n12370), .A2(n12369), .A3(n12368), .ZN(n12371) );
  AOI211_X1 U14182 ( .C1(n14728), .C2(n13952), .A(n12372), .B(n12371), .ZN(
        n12373) );
  OAI21_X1 U14183 ( .B1(n12430), .B2(n13915), .A(n12373), .ZN(P2_U3200) );
  NAND2_X1 U14184 ( .A1(n15456), .A2(n12687), .ZN(n12375) );
  NAND2_X1 U14185 ( .A1(n7456), .A2(n15332), .ZN(n12374) );
  NAND2_X1 U14186 ( .A1(n12375), .A2(n12374), .ZN(n12376) );
  XNOR2_X1 U14187 ( .A(n12376), .B(n12705), .ZN(n12594) );
  INV_X1 U14188 ( .A(n15332), .ZN(n12573) );
  NOR2_X1 U14189 ( .A1(n12377), .A2(n12573), .ZN(n12378) );
  AOI21_X1 U14190 ( .B1(n15456), .B2(n7456), .A(n12378), .ZN(n12596) );
  XNOR2_X1 U14191 ( .A(n12594), .B(n12596), .ZN(n12383) );
  INV_X1 U14192 ( .A(n12379), .ZN(n12380) );
  NAND2_X1 U14193 ( .A1(n12381), .A2(n12380), .ZN(n12384) );
  AOI21_X1 U14194 ( .B1(n12382), .B2(n12384), .A(n12383), .ZN(n12385) );
  OAI21_X1 U14195 ( .B1(n12595), .B2(n12385), .A(n14915), .ZN(n12391) );
  INV_X1 U14196 ( .A(n15303), .ZN(n12555) );
  OAI21_X1 U14197 ( .B1(n14951), .B2(n12555), .A(n12386), .ZN(n12389) );
  NOR2_X1 U14198 ( .A1(n14952), .A2(n12387), .ZN(n12388) );
  AOI211_X1 U14199 ( .C1(n14955), .C2(n14962), .A(n12389), .B(n12388), .ZN(
        n12390) );
  OAI211_X1 U14200 ( .C1(n12574), .C2(n14958), .A(n12391), .B(n12390), .ZN(
        P1_U3215) );
  XNOR2_X1 U14201 ( .A(n12392), .B(n13027), .ZN(n12393) );
  AOI222_X1 U14202 ( .A1(n16377), .A2(n12393), .B1(n13215), .B2(n13498), .C1(
        n13217), .C2(n13500), .ZN(n16557) );
  INV_X1 U14203 ( .A(n12547), .ZN(n12394) );
  OAI22_X1 U14204 ( .A1(n13587), .A2(n16559), .B1(n12394), .B2(n16405), .ZN(
        n12395) );
  AOI21_X1 U14205 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n16414), .A(n12395), 
        .ZN(n12400) );
  AND2_X1 U14206 ( .A1(n12397), .A2(n12396), .ZN(n12398) );
  XNOR2_X1 U14207 ( .A(n12398), .B(n13027), .ZN(n16562) );
  NAND2_X1 U14208 ( .A1(n16562), .A2(n13559), .ZN(n12399) );
  OAI211_X1 U14209 ( .C1(n16557), .C2(n16414), .A(n12400), .B(n12399), .ZN(
        P3_U3221) );
  INV_X1 U14210 ( .A(n12401), .ZN(n12402) );
  OAI222_X1 U14211 ( .A1(n14818), .A2(n13813), .B1(n14816), .B2(n12403), .C1(
        n12402), .C2(P2_U3088), .ZN(P2_U3303) );
  INV_X1 U14212 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n12407) );
  AOI211_X1 U14213 ( .C1(n16583), .C2(n12406), .A(n12405), .B(n12404), .ZN(
        n12409) );
  MUX2_X1 U14214 ( .A(n12407), .B(n12409), .S(n16534), .Z(n12408) );
  OAI21_X1 U14215 ( .B1(n12412), .B2(n14785), .A(n12408), .ZN(P2_U3475) );
  MUX2_X1 U14216 ( .A(n12410), .B(n12409), .S(n14740), .Z(n12411) );
  OAI21_X1 U14217 ( .B1(n12412), .B2(n14734), .A(n12411), .ZN(P2_U3514) );
  INV_X1 U14218 ( .A(n12413), .ZN(n12414) );
  NOR2_X1 U14219 ( .A1(n12414), .A2(n12416), .ZN(n12479) );
  INV_X1 U14220 ( .A(n12479), .ZN(n12415) );
  NAND2_X1 U14221 ( .A1(n12480), .A2(n12415), .ZN(n12541) );
  INV_X1 U14222 ( .A(n7614), .ZN(n12823) );
  XNOR2_X1 U14223 ( .A(n12905), .B(n12823), .ZN(n12540) );
  XNOR2_X1 U14224 ( .A(n12541), .B(n12540), .ZN(n12422) );
  OAI22_X1 U14225 ( .A1(n13198), .A2(n12416), .B1(n13157), .B2(n13187), .ZN(
        n12417) );
  AOI211_X1 U14226 ( .C1(n12919), .C2(n13168), .A(n12418), .B(n12417), .ZN(
        n12421) );
  NAND2_X1 U14227 ( .A1(n13202), .A2(n12419), .ZN(n12420) );
  OAI211_X1 U14228 ( .C1(n12422), .C2(n13204), .A(n12421), .B(n12420), .ZN(
        P3_U3176) );
  NAND2_X1 U14229 ( .A1(n12423), .A2(n14201), .ZN(n12425) );
  AOI22_X1 U14230 ( .A1(n10051), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n10048), 
        .B2(n14349), .ZN(n12424) );
  INV_X1 U14231 ( .A(n12426), .ZN(n12428) );
  NAND2_X1 U14232 ( .A1(n12428), .A2(n12427), .ZN(n12429) );
  XNOR2_X1 U14233 ( .A(n14426), .B(n7463), .ZN(n12431) );
  AND2_X1 U14234 ( .A1(n14612), .A2(n7458), .ZN(n12432) );
  NAND2_X1 U14235 ( .A1(n12431), .A2(n12432), .ZN(n12504) );
  INV_X1 U14236 ( .A(n12431), .ZN(n13886) );
  INV_X1 U14237 ( .A(n12432), .ZN(n12433) );
  NAND2_X1 U14238 ( .A1(n13886), .A2(n12433), .ZN(n12434) );
  NAND2_X1 U14239 ( .A1(n12504), .A2(n12434), .ZN(n12435) );
  AOI21_X1 U14240 ( .B1(n12436), .B2(n12435), .A(n13915), .ZN(n12437) );
  NAND2_X1 U14241 ( .A1(n12437), .A2(n13882), .ZN(n12449) );
  INV_X1 U14242 ( .A(n12456), .ZN(n12447) );
  INV_X1 U14243 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n12438) );
  NAND2_X1 U14244 ( .A1(n12439), .A2(n12438), .ZN(n12440) );
  NAND2_X1 U14245 ( .A1(n12513), .A2(n12440), .ZN(n14623) );
  INV_X1 U14246 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n14624) );
  NAND2_X1 U14247 ( .A1(n14181), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n12442) );
  NAND2_X1 U14248 ( .A1(n13902), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n12441) );
  OAI211_X1 U14249 ( .C1(n14192), .C2(n14624), .A(n12442), .B(n12441), .ZN(
        n12443) );
  INV_X1 U14250 ( .A(n12443), .ZN(n12444) );
  OAI21_X1 U14251 ( .B1(n14623), .B2(n10059), .A(n12444), .ZN(n14428) );
  AOI22_X1 U14252 ( .A1(n14428), .A2(n14614), .B1(n14613), .B2(n14305), .ZN(
        n12453) );
  OAI22_X1 U14253 ( .A1(n12453), .A2(n13975), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12445), .ZN(n12446) );
  AOI21_X1 U14254 ( .B1(n12447), .B2(n13972), .A(n12446), .ZN(n12448) );
  OAI211_X1 U14255 ( .C1(n7992), .C2(n13966), .A(n12449), .B(n12448), .ZN(
        P2_U3210) );
  NAND2_X1 U14256 ( .A1(n14789), .A2(n14306), .ZN(n12450) );
  XNOR2_X1 U14257 ( .A(n14728), .B(n14305), .ZN(n14638) );
  INV_X1 U14258 ( .A(n14638), .ZN(n14631) );
  INV_X1 U14259 ( .A(n14612), .ZN(n14386) );
  XNOR2_X1 U14260 ( .A(n14426), .B(n14386), .ZN(n14272) );
  XNOR2_X1 U14261 ( .A(n14425), .B(n14424), .ZN(n14725) );
  INV_X1 U14262 ( .A(n14725), .ZN(n12462) );
  INV_X1 U14263 ( .A(n14305), .ZN(n12452) );
  XNOR2_X1 U14264 ( .A(n14385), .B(n14424), .ZN(n12454) );
  OAI21_X1 U14265 ( .B1(n12454), .B2(n14591), .A(n12453), .ZN(n14723) );
  NAND2_X1 U14266 ( .A1(n14723), .A2(n14644), .ZN(n12461) );
  INV_X1 U14267 ( .A(n14620), .ZN(n12455) );
  AOI211_X1 U14268 ( .C1(n14426), .C2(n14648), .A(n7458), .B(n12455), .ZN(
        n14724) );
  NOR2_X1 U14269 ( .A1(n7992), .A2(n14622), .ZN(n12459) );
  OAI22_X1 U14270 ( .A1(n14644), .A2(n12457), .B1(n12456), .B2(n14641), .ZN(
        n12458) );
  AOI211_X1 U14271 ( .C1(n14724), .C2(n14650), .A(n12459), .B(n12458), .ZN(
        n12460) );
  OAI211_X1 U14272 ( .C1(n12462), .C2(n14604), .A(n12461), .B(n12460), .ZN(
        P2_U3247) );
  XNOR2_X1 U14273 ( .A(n12463), .B(n13034), .ZN(n13654) );
  INV_X1 U14274 ( .A(n13654), .ZN(n12470) );
  XNOR2_X1 U14275 ( .A(n12465), .B(n12464), .ZN(n12466) );
  OAI222_X1 U14276 ( .A1(n16372), .A2(n13568), .B1(n16374), .B2(n12543), .C1(
        n12466), .C2(n13582), .ZN(n13653) );
  AOI22_X1 U14277 ( .A1(n16414), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n16388), 
        .B2(n12499), .ZN(n12467) );
  OAI21_X1 U14278 ( .B1(n13730), .B2(n13587), .A(n12467), .ZN(n12468) );
  AOI21_X1 U14279 ( .B1(n13653), .B2(n16411), .A(n12468), .ZN(n12469) );
  OAI21_X1 U14280 ( .B1(n13590), .B2(n12470), .A(n12469), .ZN(P3_U3219) );
  XNOR2_X1 U14281 ( .A(n12472), .B(n13029), .ZN(n13662) );
  INV_X1 U14282 ( .A(n13662), .ZN(n13736) );
  XNOR2_X1 U14283 ( .A(n12473), .B(n13029), .ZN(n12474) );
  AOI222_X1 U14284 ( .A1(n16377), .A2(n12474), .B1(n13216), .B2(n13500), .C1(
        n13214), .C2(n13498), .ZN(n13658) );
  INV_X1 U14285 ( .A(n13658), .ZN(n12477) );
  AOI22_X1 U14286 ( .A1(n16414), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n16388), 
        .B2(n13159), .ZN(n12475) );
  OAI21_X1 U14287 ( .B1(n13659), .B2(n13587), .A(n12475), .ZN(n12476) );
  AOI21_X1 U14288 ( .B1(n12477), .B2(n16411), .A(n12476), .ZN(n12478) );
  OAI21_X1 U14289 ( .B1(n13590), .B2(n13736), .A(n12478), .ZN(P3_U3220) );
  INV_X1 U14290 ( .A(n12905), .ZN(n13031) );
  NAND2_X1 U14291 ( .A1(n13027), .A2(n12823), .ZN(n12486) );
  NOR3_X1 U14292 ( .A1(n12479), .A2(n13031), .A3(n12486), .ZN(n12482) );
  INV_X1 U14293 ( .A(n13027), .ZN(n12483) );
  NAND2_X1 U14294 ( .A1(n12483), .A2(n7614), .ZN(n12487) );
  NOR3_X1 U14295 ( .A1(n12479), .A2(n12487), .A3(n12905), .ZN(n12481) );
  NOR4_X1 U14296 ( .A1(n13031), .A2(n13027), .A3(n12823), .A4(n13217), .ZN(
        n12485) );
  NOR4_X1 U14297 ( .A1(n12483), .A2(n12905), .A3(n7614), .A4(n13217), .ZN(
        n12484) );
  NAND3_X1 U14298 ( .A1(n12487), .A2(n13157), .A3(n12486), .ZN(n12488) );
  XNOR2_X1 U14299 ( .A(n13659), .B(n7614), .ZN(n12492) );
  XNOR2_X1 U14300 ( .A(n12492), .B(n13215), .ZN(n13153) );
  INV_X1 U14301 ( .A(n12492), .ZN(n12493) );
  NAND2_X1 U14302 ( .A1(n12493), .A2(n13215), .ZN(n12494) );
  XNOR2_X1 U14303 ( .A(n13730), .B(n7614), .ZN(n12789) );
  XNOR2_X1 U14304 ( .A(n12789), .B(n13214), .ZN(n12787) );
  XNOR2_X1 U14305 ( .A(n12788), .B(n12787), .ZN(n12501) );
  NOR2_X1 U14306 ( .A1(n13199), .A2(n13730), .ZN(n12498) );
  INV_X1 U14307 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n12495) );
  NOR2_X1 U14308 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12495), .ZN(n13242) );
  AOI21_X1 U14309 ( .B1(n13185), .B2(n13215), .A(n13242), .ZN(n12496) );
  OAI21_X1 U14310 ( .B1(n13568), .B2(n13187), .A(n12496), .ZN(n12497) );
  AOI211_X1 U14311 ( .C1(n12499), .C2(n13202), .A(n12498), .B(n12497), .ZN(
        n12500) );
  OAI21_X1 U14312 ( .B1(n12501), .B2(n13204), .A(n12500), .ZN(P3_U3155) );
  NAND2_X1 U14313 ( .A1(n12590), .A2(n14201), .ZN(n12503) );
  AOI22_X1 U14314 ( .A1(n7465), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10130), 
        .B2(n10048), .ZN(n12502) );
  XNOR2_X1 U14315 ( .A(n14621), .B(n7463), .ZN(n12505) );
  NAND2_X1 U14316 ( .A1(n14428), .A2(n7458), .ZN(n12506) );
  XNOR2_X1 U14317 ( .A(n12505), .B(n12506), .ZN(n13887) );
  INV_X1 U14318 ( .A(n12505), .ZN(n12535) );
  NAND2_X1 U14319 ( .A1(n12535), .A2(n12506), .ZN(n12507) );
  NAND2_X1 U14320 ( .A1(n13881), .A2(n12507), .ZN(n12521) );
  NAND2_X1 U14321 ( .A1(n12508), .A2(n14201), .ZN(n12511) );
  OR2_X1 U14322 ( .A1(n14202), .A2(n12509), .ZN(n12510) );
  XNOR2_X1 U14323 ( .A(n14593), .B(n7463), .ZN(n13772) );
  INV_X1 U14324 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n12531) );
  NAND2_X1 U14325 ( .A1(n12513), .A2(n12531), .ZN(n12514) );
  AND2_X1 U14326 ( .A1(n12524), .A2(n12514), .ZN(n14599) );
  NAND2_X1 U14327 ( .A1(n14599), .A2(n13843), .ZN(n12520) );
  INV_X1 U14328 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n12517) );
  NAND2_X1 U14329 ( .A1(n13902), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n12516) );
  NAND2_X1 U14330 ( .A1(n14181), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n12515) );
  OAI211_X1 U14331 ( .C1(n12517), .C2(n14192), .A(n12516), .B(n12515), .ZN(
        n12518) );
  INV_X1 U14332 ( .A(n12518), .ZN(n12519) );
  NAND2_X1 U14333 ( .A1(n12520), .A2(n12519), .ZN(n14615) );
  NAND2_X1 U14334 ( .A1(n14615), .A2(n7458), .ZN(n13773) );
  XNOR2_X1 U14335 ( .A(n13772), .B(n13773), .ZN(n12534) );
  INV_X1 U14336 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12523) );
  NAND2_X1 U14337 ( .A1(n12524), .A2(n12523), .ZN(n12525) );
  NAND2_X1 U14338 ( .A1(n13803), .A2(n12525), .ZN(n14581) );
  OR2_X1 U14339 ( .A1(n14581), .A2(n10059), .ZN(n12530) );
  INV_X1 U14340 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n14580) );
  NAND2_X1 U14341 ( .A1(n14181), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n12527) );
  NAND2_X1 U14342 ( .A1(n13902), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n12526) );
  OAI211_X1 U14343 ( .C1(n14192), .C2(n14580), .A(n12527), .B(n12526), .ZN(
        n12528) );
  INV_X1 U14344 ( .A(n12528), .ZN(n12529) );
  NAND2_X1 U14345 ( .A1(n12530), .A2(n12529), .ZN(n14431) );
  AOI22_X1 U14346 ( .A1(n14431), .A2(n14614), .B1(n14613), .B2(n14428), .ZN(
        n14590) );
  OAI22_X1 U14347 ( .A1(n14590), .A2(n13975), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12531), .ZN(n12533) );
  INV_X1 U14348 ( .A(n14593), .ZN(n14774) );
  NOR2_X1 U14349 ( .A1(n14774), .A2(n13966), .ZN(n12532) );
  AOI211_X1 U14350 ( .C1(n13972), .C2(n14599), .A(n12533), .B(n12532), .ZN(
        n12539) );
  INV_X1 U14351 ( .A(n12534), .ZN(n12537) );
  INV_X1 U14352 ( .A(n14428), .ZN(n14390) );
  OAI22_X1 U14353 ( .A1(n12535), .A2(n13915), .B1(n14390), .B2(n13967), .ZN(
        n12536) );
  NAND3_X1 U14354 ( .A1(n13881), .A2(n12537), .A3(n12536), .ZN(n12538) );
  OAI211_X1 U14355 ( .C1(n13776), .C2(n13915), .A(n12539), .B(n12538), .ZN(
        P2_U3205) );
  XNOR2_X1 U14356 ( .A(n13027), .B(n7614), .ZN(n13151) );
  MUX2_X1 U14357 ( .A(n13217), .B(n12541), .S(n12540), .Z(n12542) );
  NOR2_X1 U14358 ( .A1(n12542), .A2(n13151), .ZN(n13150) );
  AOI21_X1 U14359 ( .B1(n13151), .B2(n12542), .A(n13150), .ZN(n12550) );
  OAI22_X1 U14360 ( .A1(n13198), .A2(n12920), .B1(n12543), .B2(n13187), .ZN(
        n12544) );
  AOI211_X1 U14361 ( .C1(n12546), .C2(n13168), .A(n12545), .B(n12544), .ZN(
        n12549) );
  NAND2_X1 U14362 ( .A1(n13202), .A2(n12547), .ZN(n12548) );
  OAI211_X1 U14363 ( .C1(n12550), .C2(n13204), .A(n12549), .B(n12548), .ZN(
        P3_U3164) );
  INV_X1 U14364 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12992) );
  OAI222_X1 U14365 ( .A1(n15916), .A2(n12992), .B1(n15919), .B2(n14186), .C1(
        P1_U3086), .C2(n12551), .ZN(P1_U3325) );
  INV_X1 U14366 ( .A(n15395), .ZN(n15173) );
  OR2_X1 U14367 ( .A1(n15456), .A2(n12573), .ZN(n12554) );
  OR2_X1 U14368 ( .A1(n15451), .A2(n12555), .ZN(n12556) );
  AND2_X1 U14369 ( .A1(n15446), .A2(n14950), .ZN(n15285) );
  NOR2_X1 U14370 ( .A1(n15284), .A2(n15285), .ZN(n12557) );
  INV_X1 U14371 ( .A(n15267), .ZN(n15275) );
  NAND2_X1 U14372 ( .A1(n15268), .A2(n15275), .ZN(n12560) );
  OR2_X1 U14373 ( .A1(n15435), .A2(n14891), .ZN(n12559) );
  INV_X1 U14374 ( .A(n15252), .ZN(n15248) );
  INV_X1 U14375 ( .A(n15270), .ZN(n15231) );
  NAND2_X1 U14376 ( .A1(n15257), .A2(n15231), .ZN(n12561) );
  INV_X1 U14377 ( .A(n15237), .ZN(n15228) );
  INV_X1 U14378 ( .A(n15258), .ZN(n15214) );
  OR2_X1 U14379 ( .A1(n15421), .A2(n15214), .ZN(n12562) );
  INV_X1 U14380 ( .A(n15199), .ZN(n15233) );
  OR2_X1 U14381 ( .A1(n12645), .A2(n15233), .ZN(n12563) );
  NAND2_X1 U14382 ( .A1(n15408), .A2(n7885), .ZN(n12564) );
  NAND2_X1 U14383 ( .A1(n12565), .A2(n12564), .ZN(n15181) );
  NAND2_X1 U14384 ( .A1(n15138), .A2(n15143), .ZN(n15137) );
  INV_X1 U14385 ( .A(n15382), .ZN(n15125) );
  NAND2_X1 U14386 ( .A1(n15125), .A2(n15147), .ZN(n12568) );
  INV_X1 U14387 ( .A(n15147), .ZN(n15111) );
  XNOR2_X1 U14388 ( .A(n15091), .B(n12580), .ZN(n12569) );
  AOI22_X1 U14389 ( .A1(n15133), .A2(n15331), .B1(n15329), .B2(n14960), .ZN(
        n12570) );
  INV_X1 U14390 ( .A(n15284), .ZN(n15282) );
  AOI21_X1 U14391 ( .B1(n15258), .B2(n15421), .A(n15426), .ZN(n15218) );
  INV_X1 U14392 ( .A(n15212), .ZN(n15217) );
  NOR2_X1 U14393 ( .A1(n15408), .A2(n14961), .ZN(n12575) );
  NAND2_X1 U14394 ( .A1(n15157), .A2(n12576), .ZN(n15142) );
  NAND2_X1 U14395 ( .A1(n15388), .A2(n15132), .ZN(n12577) );
  NAND2_X1 U14396 ( .A1(n15376), .A2(n14939), .ZN(n12578) );
  NAND2_X1 U14397 ( .A1(n15107), .A2(n12578), .ZN(n12581) );
  INV_X1 U14398 ( .A(n12581), .ZN(n12579) );
  NAND2_X1 U14399 ( .A1(n12579), .A2(n15090), .ZN(n15087) );
  NAND2_X1 U14400 ( .A1(n12581), .A2(n12580), .ZN(n12582) );
  NAND2_X1 U14401 ( .A1(n15370), .A2(n15309), .ZN(n12589) );
  INV_X1 U14402 ( .A(n15440), .ZN(n15298) );
  OR2_X1 U14403 ( .A1(n15435), .A2(n15293), .ZN(n15256) );
  OR2_X1 U14404 ( .A1(n15256), .A2(n15257), .ZN(n15254) );
  NAND2_X1 U14405 ( .A1(n15240), .A2(n8453), .ZN(n15220) );
  OR2_X1 U14406 ( .A1(n12707), .A2(n15114), .ZN(n12583) );
  AND2_X1 U14407 ( .A1(n15093), .A2(n12583), .ZN(n15372) );
  OAI22_X1 U14408 ( .A1(n15338), .A2(n12584), .B1(n12711), .B2(n15312), .ZN(
        n12585) );
  INV_X1 U14409 ( .A(n12585), .ZN(n12586) );
  OAI21_X1 U14410 ( .B1(n12707), .B2(n15310), .A(n12586), .ZN(n12587) );
  AOI21_X1 U14411 ( .B1(n15372), .B2(n15347), .A(n12587), .ZN(n12588) );
  OAI211_X1 U14412 ( .C1(n15374), .C2(n15333), .A(n12589), .B(n12588), .ZN(
        P1_U3265) );
  INV_X1 U14413 ( .A(n12590), .ZN(n12785) );
  OAI222_X1 U14414 ( .A1(n12592), .A2(P1_U3086), .B1(n15919), .B2(n12785), 
        .C1(n12591), .C2(n15916), .ZN(P1_U3336) );
  INV_X1 U14415 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n14187) );
  OAI222_X1 U14416 ( .A1(n14818), .A2(n14187), .B1(P2_U3088), .B2(n12593), 
        .C1(n14816), .C2(n14186), .ZN(P2_U3297) );
  INV_X1 U14417 ( .A(n12594), .ZN(n12597) );
  AOI22_X1 U14418 ( .A1(n15451), .A2(n12687), .B1(n7456), .B2(n15303), .ZN(
        n12598) );
  XOR2_X1 U14419 ( .A(n12705), .B(n12598), .Z(n12599) );
  INV_X1 U14420 ( .A(n12600), .ZN(n12601) );
  AOI22_X1 U14421 ( .A1(n15451), .A2(n7456), .B1(n12698), .B2(n15303), .ZN(
        n14946) );
  NAND2_X1 U14422 ( .A1(n14945), .A2(n14946), .ZN(n14944) );
  INV_X1 U14423 ( .A(n12602), .ZN(n12603) );
  NAND2_X1 U14424 ( .A1(n14944), .A2(n12603), .ZN(n14876) );
  NAND2_X1 U14425 ( .A1(n15446), .A2(n12687), .ZN(n12605) );
  NAND2_X1 U14426 ( .A1(n15330), .A2(n7456), .ZN(n12604) );
  NAND2_X1 U14427 ( .A1(n12605), .A2(n12604), .ZN(n12606) );
  XNOR2_X1 U14428 ( .A(n12606), .B(n12705), .ZN(n12610) );
  NAND2_X1 U14429 ( .A1(n15446), .A2(n7456), .ZN(n12608) );
  NAND2_X1 U14430 ( .A1(n12698), .A2(n15330), .ZN(n12607) );
  NAND2_X1 U14431 ( .A1(n12608), .A2(n12607), .ZN(n12609) );
  NOR2_X1 U14432 ( .A1(n12610), .A2(n12609), .ZN(n12611) );
  AOI21_X1 U14433 ( .B1(n12610), .B2(n12609), .A(n12611), .ZN(n14877) );
  NAND2_X1 U14434 ( .A1(n14876), .A2(n14877), .ZN(n14887) );
  INV_X1 U14435 ( .A(n12611), .ZN(n14886) );
  NAND2_X1 U14436 ( .A1(n15440), .A2(n12687), .ZN(n12613) );
  NAND2_X1 U14437 ( .A1(n15304), .A2(n7456), .ZN(n12612) );
  NAND2_X1 U14438 ( .A1(n12613), .A2(n12612), .ZN(n12614) );
  XNOR2_X1 U14439 ( .A(n12614), .B(n7593), .ZN(n12616) );
  AND2_X1 U14440 ( .A1(n12698), .A2(n15304), .ZN(n12615) );
  AOI21_X1 U14441 ( .B1(n15440), .B2(n7456), .A(n12615), .ZN(n12617) );
  NAND2_X1 U14442 ( .A1(n12616), .A2(n12617), .ZN(n12621) );
  INV_X1 U14443 ( .A(n12616), .ZN(n12619) );
  INV_X1 U14444 ( .A(n12617), .ZN(n12618) );
  NAND2_X1 U14445 ( .A1(n12619), .A2(n12618), .ZN(n12620) );
  NAND2_X1 U14446 ( .A1(n12621), .A2(n12620), .ZN(n14885) );
  AOI21_X2 U14447 ( .B1(n14887), .B2(n14886), .A(n14885), .ZN(n14927) );
  INV_X1 U14448 ( .A(n12621), .ZN(n14926) );
  NAND2_X1 U14449 ( .A1(n15435), .A2(n12687), .ZN(n12623) );
  NAND2_X1 U14450 ( .A1(n15289), .A2(n7456), .ZN(n12622) );
  NAND2_X1 U14451 ( .A1(n12623), .A2(n12622), .ZN(n12624) );
  XNOR2_X1 U14452 ( .A(n12624), .B(n7593), .ZN(n12626) );
  AND2_X1 U14453 ( .A1(n15289), .A2(n12698), .ZN(n12625) );
  AOI21_X1 U14454 ( .B1(n15435), .B2(n7456), .A(n12625), .ZN(n12627) );
  NAND2_X1 U14455 ( .A1(n12626), .A2(n12627), .ZN(n12631) );
  INV_X1 U14456 ( .A(n12626), .ZN(n12629) );
  INV_X1 U14457 ( .A(n12627), .ZN(n12628) );
  NAND2_X1 U14458 ( .A1(n12629), .A2(n12628), .ZN(n12630) );
  AND2_X1 U14459 ( .A1(n12631), .A2(n12630), .ZN(n14925) );
  NAND2_X1 U14460 ( .A1(n15257), .A2(n12687), .ZN(n12633) );
  NAND2_X1 U14461 ( .A1(n15270), .A2(n7456), .ZN(n12632) );
  NAND2_X1 U14462 ( .A1(n12633), .A2(n12632), .ZN(n12634) );
  XNOR2_X1 U14463 ( .A(n12634), .B(n12705), .ZN(n12637) );
  AOI22_X1 U14464 ( .A1(n15257), .A2(n7456), .B1(n12698), .B2(n15270), .ZN(
        n12638) );
  XNOR2_X1 U14465 ( .A(n12637), .B(n12638), .ZN(n14851) );
  AND2_X1 U14466 ( .A1(n15258), .A2(n12698), .ZN(n12635) );
  AOI21_X1 U14467 ( .B1(n15421), .B2(n7456), .A(n12635), .ZN(n12647) );
  AOI22_X1 U14468 ( .A1(n15421), .A2(n12687), .B1(n7456), .B2(n15258), .ZN(
        n12636) );
  XNOR2_X1 U14469 ( .A(n12636), .B(n12705), .ZN(n12646) );
  XOR2_X1 U14470 ( .A(n12647), .B(n12646), .Z(n14908) );
  INV_X1 U14471 ( .A(n12637), .ZN(n12639) );
  NAND2_X1 U14472 ( .A1(n12639), .A2(n12638), .ZN(n14905) );
  NAND2_X1 U14473 ( .A1(n12645), .A2(n12687), .ZN(n12642) );
  NAND2_X1 U14474 ( .A1(n15199), .A2(n7456), .ZN(n12641) );
  NAND2_X1 U14475 ( .A1(n12642), .A2(n12641), .ZN(n12643) );
  XNOR2_X1 U14476 ( .A(n12643), .B(n12705), .ZN(n12651) );
  AND2_X1 U14477 ( .A1(n15199), .A2(n12698), .ZN(n12644) );
  AOI21_X1 U14478 ( .B1(n12645), .B2(n7456), .A(n12644), .ZN(n12652) );
  XNOR2_X1 U14479 ( .A(n12651), .B(n12652), .ZN(n14857) );
  INV_X1 U14480 ( .A(n12646), .ZN(n12649) );
  INV_X1 U14481 ( .A(n12647), .ZN(n12648) );
  NAND2_X1 U14482 ( .A1(n12649), .A2(n12648), .ZN(n14858) );
  INV_X1 U14483 ( .A(n12651), .ZN(n12653) );
  NAND2_X1 U14484 ( .A1(n15408), .A2(n12687), .ZN(n12655) );
  NAND2_X1 U14485 ( .A1(n14961), .A2(n7456), .ZN(n12654) );
  NAND2_X1 U14486 ( .A1(n12655), .A2(n12654), .ZN(n12656) );
  XNOR2_X1 U14487 ( .A(n12656), .B(n12705), .ZN(n12667) );
  AND2_X1 U14488 ( .A1(n14961), .A2(n12698), .ZN(n12657) );
  AOI21_X1 U14489 ( .B1(n15408), .B2(n7456), .A(n12657), .ZN(n12665) );
  XNOR2_X1 U14490 ( .A(n12667), .B(n12665), .ZN(n14917) );
  NAND2_X1 U14491 ( .A1(n15183), .A2(n12687), .ZN(n12659) );
  NAND2_X1 U14492 ( .A1(n15198), .A2(n7456), .ZN(n12658) );
  NAND2_X1 U14493 ( .A1(n12659), .A2(n12658), .ZN(n12660) );
  XNOR2_X1 U14494 ( .A(n12660), .B(n12705), .ZN(n12664) );
  NAND2_X1 U14495 ( .A1(n15183), .A2(n7456), .ZN(n12662) );
  NAND2_X1 U14496 ( .A1(n15198), .A2(n12698), .ZN(n12661) );
  NAND2_X1 U14497 ( .A1(n12662), .A2(n12661), .ZN(n12663) );
  NOR2_X1 U14498 ( .A1(n12664), .A2(n12663), .ZN(n12668) );
  AOI21_X1 U14499 ( .B1(n12664), .B2(n12663), .A(n12668), .ZN(n14830) );
  INV_X1 U14500 ( .A(n12665), .ZN(n12666) );
  NAND2_X1 U14501 ( .A1(n12667), .A2(n12666), .ZN(n14831) );
  INV_X1 U14502 ( .A(n12668), .ZN(n12669) );
  NAND2_X1 U14503 ( .A1(n14829), .A2(n12669), .ZN(n14897) );
  NAND2_X1 U14504 ( .A1(n15395), .A2(n12687), .ZN(n12671) );
  NAND2_X1 U14505 ( .A1(n7456), .A2(n15146), .ZN(n12670) );
  NAND2_X1 U14506 ( .A1(n12671), .A2(n12670), .ZN(n12672) );
  XNOR2_X1 U14507 ( .A(n12672), .B(n12705), .ZN(n12676) );
  NAND2_X1 U14508 ( .A1(n15395), .A2(n7456), .ZN(n12674) );
  NAND2_X1 U14509 ( .A1(n12698), .A2(n15146), .ZN(n12673) );
  NAND2_X1 U14510 ( .A1(n12674), .A2(n12673), .ZN(n12675) );
  NOR2_X1 U14511 ( .A1(n12676), .A2(n12675), .ZN(n12677) );
  AOI21_X1 U14512 ( .B1(n12676), .B2(n12675), .A(n12677), .ZN(n14898) );
  INV_X1 U14513 ( .A(n12677), .ZN(n12678) );
  NAND2_X1 U14514 ( .A1(n15388), .A2(n12687), .ZN(n12680) );
  NAND2_X1 U14515 ( .A1(n7456), .A2(n15132), .ZN(n12679) );
  NAND2_X1 U14516 ( .A1(n12680), .A2(n12679), .ZN(n12681) );
  XNOR2_X1 U14517 ( .A(n12681), .B(n12705), .ZN(n12685) );
  NAND2_X1 U14518 ( .A1(n15388), .A2(n7456), .ZN(n12683) );
  NAND2_X1 U14519 ( .A1(n12698), .A2(n15132), .ZN(n12682) );
  NAND2_X1 U14520 ( .A1(n12683), .A2(n12682), .ZN(n12684) );
  NOR2_X1 U14521 ( .A1(n12685), .A2(n12684), .ZN(n12686) );
  AOI21_X1 U14522 ( .B1(n12685), .B2(n12684), .A(n12686), .ZN(n14869) );
  NAND2_X1 U14523 ( .A1(n15382), .A2(n12687), .ZN(n12689) );
  NAND2_X1 U14524 ( .A1(n7456), .A2(n15147), .ZN(n12688) );
  NAND2_X1 U14525 ( .A1(n12689), .A2(n12688), .ZN(n12690) );
  XNOR2_X1 U14526 ( .A(n12690), .B(n12705), .ZN(n12694) );
  NAND2_X1 U14527 ( .A1(n15382), .A2(n7456), .ZN(n12692) );
  NAND2_X1 U14528 ( .A1(n12698), .A2(n15147), .ZN(n12691) );
  NAND2_X1 U14529 ( .A1(n12692), .A2(n12691), .ZN(n12693) );
  NOR2_X1 U14530 ( .A1(n12694), .A2(n12693), .ZN(n12695) );
  AOI21_X1 U14531 ( .B1(n12694), .B2(n12693), .A(n12695), .ZN(n14936) );
  NAND2_X1 U14532 ( .A1(n14935), .A2(n14936), .ZN(n14934) );
  INV_X1 U14533 ( .A(n12695), .ZN(n12696) );
  NAND2_X1 U14534 ( .A1(n14934), .A2(n12696), .ZN(n14821) );
  OAI22_X1 U14535 ( .A1(n15376), .A2(n10644), .B1(n14939), .B2(n7468), .ZN(
        n12697) );
  XNOR2_X1 U14536 ( .A(n12697), .B(n12705), .ZN(n12702) );
  OR2_X1 U14537 ( .A1(n15376), .A2(n7468), .ZN(n12700) );
  NAND2_X1 U14538 ( .A1(n12698), .A2(n15133), .ZN(n12699) );
  NAND2_X1 U14539 ( .A1(n12700), .A2(n12699), .ZN(n12701) );
  NOR2_X1 U14540 ( .A1(n12702), .A2(n12701), .ZN(n12703) );
  AOI21_X1 U14541 ( .B1(n12702), .B2(n12701), .A(n12703), .ZN(n14822) );
  NAND2_X1 U14542 ( .A1(n14821), .A2(n14822), .ZN(n14820) );
  INV_X1 U14543 ( .A(n12703), .ZN(n12704) );
  AOI22_X1 U14544 ( .A1(n15371), .A2(n7456), .B1(n12698), .B2(n15085), .ZN(
        n12706) );
  XNOR2_X1 U14545 ( .A(n12706), .B(n12705), .ZN(n12709) );
  OAI22_X1 U14546 ( .A1(n12707), .A2(n10644), .B1(n15112), .B2(n7468), .ZN(
        n12708) );
  XNOR2_X1 U14547 ( .A(n12709), .B(n12708), .ZN(n12710) );
  NOR2_X1 U14548 ( .A1(n14952), .A2(n12711), .ZN(n12715) );
  AOI22_X1 U14549 ( .A1(n14955), .A2(n15133), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12712) );
  OAI21_X1 U14550 ( .B1(n12713), .B2(n14951), .A(n12712), .ZN(n12714) );
  AOI211_X1 U14551 ( .C1(n15371), .C2(n14844), .A(n12715), .B(n12714), .ZN(
        n12716) );
  AOI22_X1 U14552 ( .A1(n13950), .A2(n14309), .B1(n13888), .B2(n14311), .ZN(
        n12718) );
  OAI211_X1 U14553 ( .C1(n12719), .C2(n13943), .A(n12718), .B(n12717), .ZN(
        n12726) );
  INV_X1 U14554 ( .A(n12720), .ZN(n12724) );
  AOI22_X1 U14555 ( .A1(n12721), .A2(n13977), .B1(n13957), .B2(n14311), .ZN(
        n12723) );
  NOR3_X1 U14556 ( .A1(n12724), .A2(n12723), .A3(n12722), .ZN(n12725) );
  AOI211_X1 U14557 ( .C1(n14084), .C2(n13952), .A(n12726), .B(n12725), .ZN(
        n12727) );
  OAI21_X1 U14558 ( .B1(n12728), .B2(n13915), .A(n12727), .ZN(P2_U3196) );
  AOI22_X1 U14559 ( .A1(n13888), .A2(n14309), .B1(n13950), .B2(n14307), .ZN(
        n12729) );
  NAND2_X1 U14560 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n16196)
         );
  OAI211_X1 U14561 ( .C1(n12730), .C2(n13943), .A(n12729), .B(n16196), .ZN(
        n12737) );
  INV_X1 U14562 ( .A(n12731), .ZN(n12735) );
  AOI22_X1 U14563 ( .A1(n12732), .A2(n13977), .B1(n13957), .B2(n14309), .ZN(
        n12734) );
  NOR3_X1 U14564 ( .A1(n12735), .A2(n12734), .A3(n12733), .ZN(n12736) );
  AOI211_X1 U14565 ( .C1(n14102), .C2(n13952), .A(n12737), .B(n12736), .ZN(
        n12738) );
  OAI21_X1 U14566 ( .B1(n12739), .B2(n13915), .A(n12738), .ZN(P2_U3187) );
  NOR2_X1 U14567 ( .A1(n13943), .A2(n12740), .ZN(n12744) );
  OAI22_X1 U14568 ( .A1(n13975), .A2(n12742), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12741), .ZN(n12743) );
  AOI211_X1 U14569 ( .C1(n14789), .C2(n13952), .A(n12744), .B(n12743), .ZN(
        n12752) );
  INV_X1 U14570 ( .A(n12745), .ZN(n12749) );
  OAI22_X1 U14571 ( .A1(n12747), .A2(n13915), .B1(n12746), .B2(n13967), .ZN(
        n12748) );
  NAND3_X1 U14572 ( .A1(n12750), .A2(n12749), .A3(n12748), .ZN(n12751) );
  OAI211_X1 U14573 ( .C1(n12753), .C2(n13915), .A(n12752), .B(n12751), .ZN(
        P2_U3198) );
  NAND2_X1 U14574 ( .A1(n13972), .A2(n12754), .ZN(n12755) );
  NAND2_X1 U14575 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n14328) );
  OAI211_X1 U14576 ( .C1(n13975), .C2(n12756), .A(n12755), .B(n14328), .ZN(
        n12765) );
  INV_X1 U14577 ( .A(n12757), .ZN(n12761) );
  NOR3_X1 U14578 ( .A1(n13967), .A2(n12759), .A3(n12758), .ZN(n12760) );
  AOI21_X1 U14579 ( .B1(n12761), .B2(n13977), .A(n12760), .ZN(n12763) );
  NOR2_X1 U14580 ( .A1(n12763), .A2(n12762), .ZN(n12764) );
  AOI211_X1 U14581 ( .C1(n14044), .C2(n13952), .A(n12765), .B(n12764), .ZN(
        n12766) );
  OAI21_X1 U14582 ( .B1(n12767), .B2(n13915), .A(n12766), .ZN(P2_U3185) );
  NAND3_X1 U14583 ( .A1(n13957), .A2(n14319), .A3(n12768), .ZN(n12769) );
  OAI21_X1 U14584 ( .B1(n13915), .B2(n12770), .A(n12769), .ZN(n12778) );
  INV_X1 U14585 ( .A(n12771), .ZN(n12777) );
  AOI22_X1 U14586 ( .A1(n13945), .A2(n12772), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12774) );
  NAND2_X1 U14587 ( .A1(n13952), .A2(n14026), .ZN(n12773) );
  OAI211_X1 U14588 ( .C1(n13943), .C2(n12775), .A(n12774), .B(n12773), .ZN(
        n12776) );
  AOI21_X1 U14589 ( .B1(n12778), .B2(n12777), .A(n12776), .ZN(n12779) );
  OAI21_X1 U14590 ( .B1(n12780), .B2(n13915), .A(n12779), .ZN(P2_U3202) );
  INV_X1 U14591 ( .A(n14802), .ZN(n12782) );
  OAI222_X1 U14592 ( .A1(n9943), .A2(P1_U3086), .B1(n15919), .B2(n12782), .C1(
        n12781), .C2(n15916), .ZN(P1_U3327) );
  OAI222_X1 U14593 ( .A1(n13750), .A2(n12784), .B1(n13745), .B2(n15498), .C1(
        P3_U3151), .C2(n7728), .ZN(P3_U3267) );
  OAI222_X1 U14594 ( .A1(n14818), .A2(n12786), .B1(n14816), .B2(n12785), .C1(
        n14366), .C2(P2_U3088), .ZN(P2_U3308) );
  INV_X1 U14595 ( .A(n12789), .ZN(n12790) );
  XNOR2_X1 U14596 ( .A(n13726), .B(n7614), .ZN(n12791) );
  NAND2_X1 U14597 ( .A1(n12791), .A2(n13568), .ZN(n13191) );
  NAND2_X1 U14598 ( .A1(n13193), .A2(n13191), .ZN(n12793) );
  INV_X1 U14599 ( .A(n12791), .ZN(n12792) );
  NAND2_X1 U14600 ( .A1(n12792), .A2(n13213), .ZN(n13192) );
  XNOR2_X1 U14601 ( .A(n13118), .B(n7614), .ZN(n12794) );
  XNOR2_X1 U14602 ( .A(n12794), .B(n13584), .ZN(n13120) );
  NAND2_X1 U14603 ( .A1(n12794), .A2(n13212), .ZN(n12795) );
  NAND2_X1 U14604 ( .A1(n13119), .A2(n12795), .ZN(n13128) );
  XNOR2_X1 U14605 ( .A(n13644), .B(n7614), .ZN(n12796) );
  XNOR2_X1 U14606 ( .A(n12796), .B(n13211), .ZN(n13127) );
  INV_X1 U14607 ( .A(n12796), .ZN(n12797) );
  NAND2_X1 U14608 ( .A1(n12797), .A2(n13211), .ZN(n12798) );
  XNOR2_X1 U14609 ( .A(n13171), .B(n7614), .ZN(n12799) );
  XNOR2_X1 U14610 ( .A(n12799), .B(n13548), .ZN(n13173) );
  NAND2_X1 U14611 ( .A1(n12799), .A2(n13210), .ZN(n12800) );
  XNOR2_X1 U14612 ( .A(n13085), .B(n7614), .ZN(n12801) );
  XNOR2_X1 U14613 ( .A(n12801), .B(n13540), .ZN(n13087) );
  NAND2_X1 U14614 ( .A1(n12801), .A2(n13209), .ZN(n12802) );
  NAND2_X1 U14615 ( .A1(n13086), .A2(n12802), .ZN(n13145) );
  XNOR2_X1 U14616 ( .A(n13142), .B(n7614), .ZN(n12803) );
  XNOR2_X1 U14617 ( .A(n12803), .B(n13527), .ZN(n13144) );
  NAND2_X1 U14618 ( .A1(n12803), .A2(n13501), .ZN(n12804) );
  NAND2_X1 U14619 ( .A1(n13143), .A2(n12804), .ZN(n13097) );
  INV_X1 U14620 ( .A(n12852), .ZN(n12807) );
  INV_X1 U14621 ( .A(n12805), .ZN(n12806) );
  MUX2_X1 U14622 ( .A(n12807), .B(n12806), .S(n7614), .Z(n13095) );
  MUX2_X1 U14623 ( .A(n12853), .B(n12808), .S(n7614), .Z(n13093) );
  XOR2_X1 U14624 ( .A(n7614), .B(n13486), .Z(n12809) );
  NAND2_X1 U14625 ( .A1(n12810), .A2(n12809), .ZN(n12813) );
  INV_X1 U14626 ( .A(n13164), .ZN(n12812) );
  NAND2_X1 U14627 ( .A1(n13162), .A2(n12813), .ZN(n12817) );
  INV_X1 U14628 ( .A(n12817), .ZN(n12815) );
  XOR2_X1 U14629 ( .A(n7614), .B(n13469), .Z(n12816) );
  NAND2_X1 U14630 ( .A1(n12815), .A2(n12814), .ZN(n12818) );
  NAND2_X1 U14631 ( .A1(n12817), .A2(n12816), .ZN(n13133) );
  XNOR2_X1 U14632 ( .A(n13687), .B(n7614), .ZN(n12819) );
  NAND2_X1 U14633 ( .A1(n12819), .A2(n13439), .ZN(n13107) );
  INV_X1 U14634 ( .A(n12819), .ZN(n12820) );
  NAND2_X1 U14635 ( .A1(n12820), .A2(n13466), .ZN(n12821) );
  NAND2_X1 U14636 ( .A1(n12822), .A2(n13134), .ZN(n13105) );
  NAND2_X1 U14637 ( .A1(n13105), .A2(n13107), .ZN(n12827) );
  XNOR2_X1 U14638 ( .A(n13104), .B(n12823), .ZN(n12824) );
  NAND2_X1 U14639 ( .A1(n12824), .A2(n13453), .ZN(n12828) );
  INV_X1 U14640 ( .A(n12824), .ZN(n12825) );
  NAND2_X1 U14641 ( .A1(n12825), .A2(n13208), .ZN(n12826) );
  NAND2_X1 U14642 ( .A1(n12827), .A2(n13108), .ZN(n13110) );
  NAND2_X1 U14643 ( .A1(n13110), .A2(n12828), .ZN(n13181) );
  XNOR2_X1 U14644 ( .A(n13179), .B(n7614), .ZN(n12829) );
  NOR2_X1 U14645 ( .A1(n12829), .A2(n13207), .ZN(n12830) );
  AOI21_X1 U14646 ( .B1(n13207), .B2(n12829), .A(n12830), .ZN(n13182) );
  INV_X1 U14647 ( .A(n12830), .ZN(n12831) );
  XNOR2_X1 U14648 ( .A(n13412), .B(n7614), .ZN(n12832) );
  NOR2_X1 U14649 ( .A1(n12832), .A2(n13392), .ZN(n12833) );
  XNOR2_X1 U14650 ( .A(n13387), .B(n7614), .ZN(n12835) );
  NAND2_X1 U14651 ( .A1(n13202), .A2(n13396), .ZN(n12837) );
  AOI22_X1 U14652 ( .A1(n13185), .A2(n13392), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12836) );
  OAI211_X1 U14653 ( .C1(n12838), .C2(n13187), .A(n12837), .B(n12836), .ZN(
        n12839) );
  AOI21_X1 U14654 ( .B1(n12978), .B2(n13168), .A(n12839), .ZN(n12840) );
  INV_X1 U14655 ( .A(n13687), .ZN(n12842) );
  NAND2_X1 U14656 ( .A1(n12842), .A2(n13439), .ZN(n12969) );
  INV_X1 U14657 ( .A(n12843), .ZN(n12846) );
  INV_X1 U14658 ( .A(n12844), .ZN(n12845) );
  AOI211_X1 U14659 ( .C1(n13424), .C2(n12847), .A(n12846), .B(n12845), .ZN(
        n12850) );
  INV_X1 U14660 ( .A(n12848), .ZN(n12849) );
  NOR2_X1 U14661 ( .A1(n12850), .A2(n12849), .ZN(n12974) );
  MUX2_X1 U14662 ( .A(n12851), .B(n13462), .S(n12961), .Z(n12959) );
  INV_X1 U14663 ( .A(n13482), .ZN(n13475) );
  MUX2_X1 U14664 ( .A(n12853), .B(n12852), .S(n12975), .Z(n12957) );
  NAND4_X1 U14665 ( .A1(n13017), .A2(n12855), .A3(n12858), .A4(n12854), .ZN(
        n12862) );
  NAND2_X1 U14666 ( .A1(n12857), .A2(n12856), .ZN(n12860) );
  AND2_X1 U14667 ( .A1(n12858), .A2(n12961), .ZN(n12859) );
  NAND2_X1 U14668 ( .A1(n12860), .A2(n12859), .ZN(n12864) );
  INV_X1 U14669 ( .A(n12864), .ZN(n12861) );
  AOI21_X1 U14670 ( .B1(n12863), .B2(n12862), .A(n12861), .ZN(n12874) );
  NAND2_X1 U14671 ( .A1(n12864), .A2(n13017), .ZN(n12866) );
  NAND3_X1 U14672 ( .A1(n12866), .A2(n12865), .A3(n12870), .ZN(n12869) );
  NAND2_X1 U14673 ( .A1(n12871), .A2(n12867), .ZN(n12868) );
  MUX2_X1 U14674 ( .A(n12869), .B(n12868), .S(n12975), .Z(n12873) );
  MUX2_X1 U14675 ( .A(n12871), .B(n12870), .S(n12975), .Z(n12872) );
  OAI21_X1 U14676 ( .B1(n12874), .B2(n12873), .A(n12872), .ZN(n12875) );
  NAND2_X1 U14677 ( .A1(n12875), .A2(n13016), .ZN(n12879) );
  MUX2_X1 U14678 ( .A(n12877), .B(n12876), .S(n12975), .Z(n12878) );
  NAND3_X1 U14679 ( .A1(n12879), .A2(n13015), .A3(n12878), .ZN(n12883) );
  MUX2_X1 U14680 ( .A(n12881), .B(n12880), .S(n12975), .Z(n12882) );
  NAND3_X1 U14681 ( .A1(n12883), .A2(n13023), .A3(n12882), .ZN(n12889) );
  NAND2_X1 U14682 ( .A1(n13222), .A2(n12975), .ZN(n12886) );
  NAND2_X1 U14683 ( .A1(n12884), .A2(n12961), .ZN(n12885) );
  MUX2_X1 U14684 ( .A(n12886), .B(n12885), .S(n16470), .Z(n12887) );
  NAND3_X1 U14685 ( .A1(n12889), .A2(n12888), .A3(n12887), .ZN(n12894) );
  MUX2_X1 U14686 ( .A(n12975), .B(n13221), .S(n12890), .Z(n12891) );
  OAI21_X1 U14687 ( .B1(n12892), .B2(n12961), .A(n12891), .ZN(n12893) );
  NAND3_X1 U14688 ( .A1(n12894), .A2(n13022), .A3(n12893), .ZN(n12898) );
  NAND2_X1 U14689 ( .A1(n13220), .A2(n16485), .ZN(n12896) );
  MUX2_X1 U14690 ( .A(n12896), .B(n12895), .S(n12961), .Z(n12897) );
  NAND3_X1 U14691 ( .A1(n12898), .A2(n13014), .A3(n12897), .ZN(n12902) );
  MUX2_X1 U14692 ( .A(n12900), .B(n12899), .S(n12975), .Z(n12901) );
  NAND3_X1 U14693 ( .A1(n12902), .A2(n9070), .A3(n12901), .ZN(n12908) );
  MUX2_X1 U14694 ( .A(n12904), .B(n12903), .S(n12975), .Z(n12906) );
  AND2_X1 U14695 ( .A1(n12906), .A2(n12905), .ZN(n12907) );
  NAND2_X1 U14696 ( .A1(n12908), .A2(n12907), .ZN(n12918) );
  NAND3_X1 U14697 ( .A1(n12918), .A2(n12921), .A3(n12909), .ZN(n12910) );
  NAND3_X1 U14698 ( .A1(n12910), .A2(n12917), .A3(n12975), .ZN(n12911) );
  NAND2_X1 U14699 ( .A1(n12911), .A2(n13029), .ZN(n12913) );
  NAND3_X1 U14700 ( .A1(n13659), .A2(n13215), .A3(n12975), .ZN(n12912) );
  NAND2_X1 U14701 ( .A1(n12913), .A2(n12912), .ZN(n12914) );
  NAND3_X1 U14702 ( .A1(n12914), .A2(n13034), .A3(n13580), .ZN(n12916) );
  NAND3_X1 U14703 ( .A1(n13726), .A2(n13213), .A3(n12975), .ZN(n12915) );
  NAND2_X1 U14704 ( .A1(n12916), .A2(n12915), .ZN(n12924) );
  OAI211_X1 U14705 ( .C1(n12920), .C2(n12919), .A(n12918), .B(n12917), .ZN(
        n12922) );
  NAND3_X1 U14706 ( .A1(n12922), .A2(n12961), .A3(n12921), .ZN(n12923) );
  NAND2_X1 U14707 ( .A1(n12924), .A2(n12923), .ZN(n12932) );
  AOI21_X1 U14708 ( .B1(n12926), .B2(n12925), .A(n12975), .ZN(n12928) );
  MUX2_X1 U14709 ( .A(n12975), .B(n12928), .S(n12927), .Z(n12930) );
  AOI22_X1 U14710 ( .A1(n13580), .A2(n12930), .B1(n8407), .B2(n12961), .ZN(
        n12931) );
  NAND2_X1 U14711 ( .A1(n12932), .A2(n12931), .ZN(n12940) );
  MUX2_X1 U14712 ( .A(n13212), .B(n13118), .S(n12975), .Z(n12936) );
  NAND2_X1 U14713 ( .A1(n12936), .A2(n12933), .ZN(n12939) );
  INV_X1 U14714 ( .A(n12934), .ZN(n12935) );
  OR2_X1 U14715 ( .A1(n12936), .A2(n12935), .ZN(n12937) );
  NAND4_X1 U14716 ( .A1(n12946), .A2(n12944), .A3(n13557), .A4(n12937), .ZN(
        n12938) );
  AOI21_X1 U14717 ( .B1(n12940), .B2(n12939), .A(n12938), .ZN(n12951) );
  INV_X1 U14718 ( .A(n12946), .ZN(n12943) );
  INV_X1 U14719 ( .A(n12941), .ZN(n13011) );
  OAI211_X1 U14720 ( .C1(n12943), .C2(n12942), .A(n13011), .B(n12944), .ZN(
        n12948) );
  NAND3_X1 U14721 ( .A1(n12944), .A2(n13211), .A3(n13644), .ZN(n12945) );
  NAND3_X1 U14722 ( .A1(n13012), .A2(n12946), .A3(n12945), .ZN(n12947) );
  MUX2_X1 U14723 ( .A(n12948), .B(n12947), .S(n12961), .Z(n12950) );
  MUX2_X1 U14724 ( .A(n13011), .B(n13012), .S(n12975), .Z(n12949) );
  OAI211_X1 U14725 ( .C1(n12951), .C2(n12950), .A(n13512), .B(n12949), .ZN(
        n12955) );
  MUX2_X1 U14726 ( .A(n12953), .B(n12952), .S(n12961), .Z(n12954) );
  NAND3_X1 U14727 ( .A1(n12955), .A2(n13494), .A3(n12954), .ZN(n12956) );
  NAND3_X1 U14728 ( .A1(n13475), .A2(n12957), .A3(n12956), .ZN(n12958) );
  NAND3_X1 U14729 ( .A1(n12960), .A2(n12959), .A3(n12958), .ZN(n12965) );
  NAND2_X1 U14730 ( .A1(n13478), .A2(n12975), .ZN(n12963) );
  NAND2_X1 U14731 ( .A1(n13454), .A2(n12961), .ZN(n12962) );
  MUX2_X1 U14732 ( .A(n12963), .B(n12962), .S(n13469), .Z(n12964) );
  NAND2_X1 U14733 ( .A1(n12965), .A2(n12964), .ZN(n12966) );
  NAND2_X1 U14734 ( .A1(n13447), .A2(n12966), .ZN(n12967) );
  INV_X1 U14735 ( .A(n12972), .ZN(n12968) );
  OAI211_X1 U14736 ( .C1(n12970), .C2(n12969), .A(n12974), .B(n12968), .ZN(
        n12976) );
  INV_X1 U14737 ( .A(n12970), .ZN(n13039) );
  NAND2_X1 U14738 ( .A1(n13039), .A2(n12971), .ZN(n12973) );
  INV_X1 U14739 ( .A(n12977), .ZN(n12980) );
  NAND2_X1 U14740 ( .A1(n13673), .A2(n13404), .ZN(n12979) );
  OAI211_X1 U14741 ( .C1(n12981), .C2(n12980), .A(n13051), .B(n12979), .ZN(
        n12989) );
  NAND2_X1 U14742 ( .A1(n12983), .A2(n12982), .ZN(n12985) );
  INV_X1 U14743 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15907) );
  NAND2_X1 U14744 ( .A1(n15907), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12984) );
  XNOR2_X1 U14745 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n12990) );
  INV_X1 U14746 ( .A(n12990), .ZN(n12986) );
  XNOR2_X1 U14747 ( .A(n12991), .B(n12986), .ZN(n13068) );
  NAND2_X1 U14748 ( .A1(n13068), .A2(n12997), .ZN(n12988) );
  INV_X1 U14749 ( .A(SI_30_), .ZN(n13070) );
  OR2_X1 U14750 ( .A1(n7461), .A2(n13070), .ZN(n12987) );
  NAND2_X1 U14751 ( .A1(n12988), .A2(n12987), .ZN(n13006) );
  NAND2_X1 U14752 ( .A1(n13006), .A2(n13007), .ZN(n13047) );
  NAND3_X1 U14753 ( .A1(n12989), .A2(n13048), .A3(n13047), .ZN(n13010) );
  NAND2_X1 U14754 ( .A1(n12991), .A2(n12990), .ZN(n12994) );
  NAND2_X1 U14755 ( .A1(n12992), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12993) );
  NAND2_X1 U14756 ( .A1(n12994), .A2(n12993), .ZN(n12996) );
  INV_X1 U14757 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n14794) );
  XNOR2_X1 U14758 ( .A(n14794), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n12995) );
  XNOR2_X1 U14759 ( .A(n12996), .B(n12995), .ZN(n13740) );
  NAND2_X1 U14760 ( .A1(n13740), .A2(n12997), .ZN(n12999) );
  INV_X1 U14761 ( .A(SI_31_), .ZN(n13746) );
  OR2_X1 U14762 ( .A1(n7461), .A2(n13746), .ZN(n12998) );
  NAND2_X1 U14763 ( .A1(n9009), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n13003) );
  NAND2_X1 U14764 ( .A1(n9010), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n13002) );
  NAND2_X1 U14765 ( .A1(n13000), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13001) );
  NAND4_X1 U14766 ( .A1(n13004), .A2(n13003), .A3(n13002), .A4(n13001), .ZN(
        n13375) );
  INV_X1 U14767 ( .A(n13375), .ZN(n13005) );
  AND2_X1 U14768 ( .A1(n13054), .A2(n13005), .ZN(n13053) );
  INV_X1 U14769 ( .A(n13053), .ZN(n13009) );
  INV_X1 U14770 ( .A(n13007), .ZN(n13206) );
  AND2_X1 U14771 ( .A1(n13670), .A2(n13206), .ZN(n13055) );
  INV_X1 U14772 ( .A(n13055), .ZN(n13008) );
  AND2_X1 U14773 ( .A1(n13667), .A2(n13375), .ZN(n13050) );
  AOI21_X1 U14774 ( .B1(n13010), .B2(n13042), .A(n13050), .ZN(n13059) );
  INV_X1 U14775 ( .A(n13494), .ZN(n13496) );
  NAND2_X1 U14776 ( .A1(n13012), .A2(n13011), .ZN(n13525) );
  NAND4_X1 U14777 ( .A1(n13016), .A2(n13015), .A3(n13014), .A4(n13013), .ZN(
        n13021) );
  INV_X1 U14778 ( .A(n16370), .ZN(n13019) );
  NAND3_X1 U14779 ( .A1(n13019), .A2(n13018), .A3(n13017), .ZN(n13020) );
  NOR2_X1 U14780 ( .A1(n13021), .A2(n13020), .ZN(n13028) );
  AND2_X1 U14781 ( .A1(n13023), .A2(n13022), .ZN(n13026) );
  NOR2_X1 U14782 ( .A1(n13024), .A2(n8399), .ZN(n13025) );
  NAND4_X1 U14783 ( .A1(n13028), .A2(n13027), .A3(n13026), .A4(n13025), .ZN(
        n13032) );
  INV_X1 U14784 ( .A(n13029), .ZN(n13030) );
  NOR3_X1 U14785 ( .A1(n13032), .A2(n13031), .A3(n13030), .ZN(n13033) );
  NAND4_X1 U14786 ( .A1(n13564), .A2(n13580), .A3(n13034), .A4(n13033), .ZN(
        n13035) );
  OR4_X1 U14787 ( .A1(n13525), .A2(n8859), .A3(n8349), .A4(n13035), .ZN(n13036) );
  OR4_X1 U14788 ( .A1(n13482), .A2(n13037), .A3(n13496), .A4(n13036), .ZN(
        n13038) );
  OAI211_X1 U14789 ( .C1(n13670), .C2(n13375), .A(n13048), .B(n13047), .ZN(
        n13049) );
  NOR2_X1 U14790 ( .A1(n13057), .A2(n13056), .ZN(n13058) );
  NAND3_X1 U14791 ( .A1(n13062), .A2(n13061), .A3(n13357), .ZN(n13063) );
  OAI211_X1 U14792 ( .C1(n13064), .C2(n13066), .A(n13063), .B(P3_B_REG_SCAN_IN), .ZN(n13065) );
  OAI21_X1 U14793 ( .B1(n13067), .B2(n13066), .A(n13065), .ZN(P3_U3296) );
  INV_X1 U14794 ( .A(n13068), .ZN(n13069) );
  OAI222_X1 U14795 ( .A1(n13071), .A2(P3_U3151), .B1(n13745), .B2(n13070), 
        .C1(n13750), .C2(n13069), .ZN(P3_U3265) );
  INV_X1 U14796 ( .A(n13412), .ZN(n13677) );
  AOI22_X1 U14797 ( .A1(n13185), .A2(n13207), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13075) );
  OAI21_X1 U14798 ( .B1(n13076), .B2(n13187), .A(n13075), .ZN(n13077) );
  AOI21_X1 U14799 ( .B1(n13408), .B2(n13202), .A(n13077), .ZN(n13078) );
  AOI21_X1 U14800 ( .B1(n13478), .B2(n13079), .A(n7471), .ZN(n13084) );
  NAND2_X1 U14801 ( .A1(n13202), .A2(n13470), .ZN(n13081) );
  AOI22_X1 U14802 ( .A1(n13185), .A2(n13499), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13080) );
  OAI211_X1 U14803 ( .C1(n13439), .C2(n13187), .A(n13081), .B(n13080), .ZN(
        n13082) );
  AOI21_X1 U14804 ( .B1(n13469), .B2(n13168), .A(n13082), .ZN(n13083) );
  OAI21_X1 U14805 ( .B1(n13084), .B2(n13204), .A(n13083), .ZN(P3_U3156) );
  INV_X1 U14806 ( .A(n13085), .ZN(n13713) );
  OAI211_X1 U14807 ( .C1(n13088), .C2(n13087), .A(n13086), .B(n13183), .ZN(
        n13092) );
  NAND2_X1 U14808 ( .A1(n13185), .A2(n13210), .ZN(n13089) );
  NAND2_X1 U14809 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13367)
         );
  OAI211_X1 U14810 ( .C1(n13527), .C2(n13187), .A(n13089), .B(n13367), .ZN(
        n13090) );
  AOI21_X1 U14811 ( .B1(n13528), .B2(n13202), .A(n13090), .ZN(n13091) );
  OAI211_X1 U14812 ( .C1(n13713), .C2(n13199), .A(n13092), .B(n13091), .ZN(
        P3_U3159) );
  INV_X1 U14813 ( .A(n13093), .ZN(n13094) );
  NOR2_X1 U14814 ( .A1(n13095), .A2(n13094), .ZN(n13096) );
  XNOR2_X1 U14815 ( .A(n13097), .B(n13096), .ZN(n13103) );
  NAND2_X1 U14816 ( .A1(n13202), .A2(n13507), .ZN(n13099) );
  AOI22_X1 U14817 ( .A1(n13185), .A2(n13501), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13098) );
  OAI211_X1 U14818 ( .C1(n13100), .C2(n13187), .A(n13099), .B(n13098), .ZN(
        n13101) );
  AOI21_X1 U14819 ( .B1(n13702), .B2(n13168), .A(n13101), .ZN(n13102) );
  OAI21_X1 U14820 ( .B1(n13103), .B2(n13204), .A(n13102), .ZN(P3_U3163) );
  INV_X1 U14821 ( .A(n13106), .ZN(n13136) );
  INV_X1 U14822 ( .A(n13107), .ZN(n13109) );
  NOR3_X1 U14823 ( .A1(n13136), .A2(n13109), .A3(n13108), .ZN(n13113) );
  INV_X1 U14824 ( .A(n13111), .ZN(n13112) );
  OAI21_X1 U14825 ( .B1(n13113), .B2(n13112), .A(n13183), .ZN(n13117) );
  AOI22_X1 U14826 ( .A1(n13196), .A2(n13207), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13114) );
  OAI21_X1 U14827 ( .B1(n13439), .B2(n13198), .A(n13114), .ZN(n13115) );
  AOI21_X1 U14828 ( .B1(n13442), .B2(n13202), .A(n13115), .ZN(n13116) );
  OAI211_X1 U14829 ( .C1(n13685), .C2(n13199), .A(n13117), .B(n13116), .ZN(
        P3_U3165) );
  INV_X1 U14830 ( .A(n13118), .ZN(n13722) );
  OAI211_X1 U14831 ( .C1(n13121), .C2(n13120), .A(n13119), .B(n13183), .ZN(
        n13125) );
  NAND2_X1 U14832 ( .A1(n13185), .A2(n13213), .ZN(n13122) );
  NAND2_X1 U14833 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n13281)
         );
  OAI211_X1 U14834 ( .C1(n13569), .C2(n13187), .A(n13122), .B(n13281), .ZN(
        n13123) );
  AOI21_X1 U14835 ( .B1(n13570), .B2(n13202), .A(n13123), .ZN(n13124) );
  OAI211_X1 U14836 ( .C1(n13722), .C2(n13199), .A(n13125), .B(n13124), .ZN(
        P3_U3166) );
  OAI211_X1 U14837 ( .C1(n13128), .C2(n13127), .A(n13126), .B(n13183), .ZN(
        n13132) );
  NAND2_X1 U14838 ( .A1(n13185), .A2(n13212), .ZN(n13129) );
  NAND2_X1 U14839 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13313)
         );
  OAI211_X1 U14840 ( .C1(n13548), .C2(n13187), .A(n13129), .B(n13313), .ZN(
        n13130) );
  AOI21_X1 U14841 ( .B1(n13551), .B2(n13202), .A(n13130), .ZN(n13131) );
  OAI211_X1 U14842 ( .C1(n13199), .C2(n13644), .A(n13132), .B(n13131), .ZN(
        P3_U3168) );
  INV_X1 U14843 ( .A(n13133), .ZN(n13135) );
  NOR3_X1 U14844 ( .A1(n7471), .A2(n13135), .A3(n13134), .ZN(n13137) );
  OAI21_X1 U14845 ( .B1(n13137), .B2(n13136), .A(n13183), .ZN(n13141) );
  AOI22_X1 U14846 ( .A1(n13196), .A2(n13208), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13138) );
  OAI21_X1 U14847 ( .B1(n13454), .B2(n13198), .A(n13138), .ZN(n13139) );
  AOI21_X1 U14848 ( .B1(n13449), .B2(n13202), .A(n13139), .ZN(n13140) );
  OAI211_X1 U14849 ( .C1(n13199), .C2(n13687), .A(n13141), .B(n13140), .ZN(
        P3_U3169) );
  INV_X1 U14850 ( .A(n13142), .ZN(n13628) );
  OAI211_X1 U14851 ( .C1(n13145), .C2(n13144), .A(n13143), .B(n13183), .ZN(
        n13149) );
  AOI22_X1 U14852 ( .A1(n13196), .A2(n13479), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13146) );
  OAI21_X1 U14853 ( .B1(n13540), .B2(n13198), .A(n13146), .ZN(n13147) );
  AOI21_X1 U14854 ( .B1(n13518), .B2(n13202), .A(n13147), .ZN(n13148) );
  OAI211_X1 U14855 ( .C1(n13628), .C2(n13199), .A(n13149), .B(n13148), .ZN(
        P3_U3173) );
  AOI21_X1 U14856 ( .B1(n13151), .B2(n13157), .A(n13150), .ZN(n13154) );
  OAI211_X1 U14857 ( .C1(n13154), .C2(n13153), .A(n13183), .B(n13152), .ZN(
        n13161) );
  AOI21_X1 U14858 ( .B1(n13196), .B2(n13214), .A(n13155), .ZN(n13156) );
  OAI21_X1 U14859 ( .B1(n13157), .B2(n13198), .A(n13156), .ZN(n13158) );
  AOI21_X1 U14860 ( .B1(n13159), .B2(n13202), .A(n13158), .ZN(n13160) );
  OAI211_X1 U14861 ( .C1(n13199), .C2(n13659), .A(n13161), .B(n13160), .ZN(
        P3_U3174) );
  INV_X1 U14862 ( .A(n13162), .ZN(n13163) );
  AOI21_X1 U14863 ( .B1(n13499), .B2(n13164), .A(n13163), .ZN(n13170) );
  NAND2_X1 U14864 ( .A1(n13202), .A2(n13487), .ZN(n13166) );
  AOI22_X1 U14865 ( .A1(n13185), .A2(n13479), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13165) );
  OAI211_X1 U14866 ( .C1(n13454), .C2(n13187), .A(n13166), .B(n13165), .ZN(
        n13167) );
  AOI21_X1 U14867 ( .B1(n13486), .B2(n13168), .A(n13167), .ZN(n13169) );
  OAI21_X1 U14868 ( .B1(n13170), .B2(n13204), .A(n13169), .ZN(P3_U3175) );
  INV_X1 U14869 ( .A(n13171), .ZN(n13717) );
  OAI211_X1 U14870 ( .C1(n13174), .C2(n13173), .A(n13172), .B(n13183), .ZN(
        n13178) );
  AND2_X1 U14871 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13340) );
  AOI21_X1 U14872 ( .B1(n13196), .B2(n13209), .A(n13340), .ZN(n13175) );
  OAI21_X1 U14873 ( .B1(n13569), .B2(n13198), .A(n13175), .ZN(n13176) );
  AOI21_X1 U14874 ( .B1(n13541), .B2(n13202), .A(n13176), .ZN(n13177) );
  OAI211_X1 U14875 ( .C1(n13717), .C2(n13199), .A(n13178), .B(n13177), .ZN(
        P3_U3178) );
  NAND2_X1 U14876 ( .A1(n13184), .A2(n13183), .ZN(n13190) );
  AOI22_X1 U14877 ( .A1(n13185), .A2(n13208), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13186) );
  OAI21_X1 U14878 ( .B1(n13421), .B2(n13187), .A(n13186), .ZN(n13188) );
  AOI21_X1 U14879 ( .B1(n13429), .B2(n13202), .A(n13188), .ZN(n13189) );
  OAI211_X1 U14880 ( .C1(n13681), .C2(n13199), .A(n13190), .B(n13189), .ZN(
        P3_U3180) );
  NAND2_X1 U14881 ( .A1(n13192), .A2(n13191), .ZN(n13194) );
  XOR2_X1 U14882 ( .A(n13194), .B(n13193), .Z(n13205) );
  INV_X1 U14883 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n13195) );
  NOR2_X1 U14884 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13195), .ZN(n13259) );
  AOI21_X1 U14885 ( .B1(n13196), .B2(n13212), .A(n13259), .ZN(n13197) );
  OAI21_X1 U14886 ( .B1(n13583), .B2(n13198), .A(n13197), .ZN(n13201) );
  NOR2_X1 U14887 ( .A1(n13726), .A2(n13199), .ZN(n13200) );
  AOI211_X1 U14888 ( .C1(n13585), .C2(n13202), .A(n13201), .B(n13200), .ZN(
        n13203) );
  OAI21_X1 U14889 ( .B1(n13205), .B2(n13204), .A(n13203), .ZN(P3_U3181) );
  MUX2_X1 U14890 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n13375), .S(n16079), .Z(
        P3_U3522) );
  MUX2_X1 U14891 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n13206), .S(n16079), .Z(
        P3_U3521) );
  MUX2_X1 U14892 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n13393), .S(n16079), .Z(
        P3_U3520) );
  MUX2_X1 U14893 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n13404), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14894 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n13392), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14895 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n13207), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14896 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n13208), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14897 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n13466), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14898 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n13478), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14899 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n13499), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14900 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n13479), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14901 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13501), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14902 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n13209), .S(n16079), .Z(
        P3_U3510) );
  MUX2_X1 U14903 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13210), .S(n16079), .Z(
        P3_U3509) );
  MUX2_X1 U14904 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13211), .S(n16079), .Z(
        P3_U3508) );
  MUX2_X1 U14905 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13212), .S(n16079), .Z(
        P3_U3507) );
  MUX2_X1 U14906 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n13213), .S(n16079), .Z(
        P3_U3506) );
  MUX2_X1 U14907 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n13214), .S(n16079), .Z(
        P3_U3505) );
  MUX2_X1 U14908 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n13215), .S(n16079), .Z(
        P3_U3504) );
  MUX2_X1 U14909 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13216), .S(n16079), .Z(
        P3_U3503) );
  MUX2_X1 U14910 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n13217), .S(n16079), .Z(
        P3_U3502) );
  MUX2_X1 U14911 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n13218), .S(n16079), .Z(
        P3_U3501) );
  MUX2_X1 U14912 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n13219), .S(n16079), .Z(
        P3_U3500) );
  MUX2_X1 U14913 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n13220), .S(n16079), .Z(
        P3_U3499) );
  MUX2_X1 U14914 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n13221), .S(n16079), .Z(
        P3_U3498) );
  MUX2_X1 U14915 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13222), .S(n16079), .Z(
        P3_U3497) );
  MUX2_X1 U14916 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n13223), .S(n16079), .Z(
        P3_U3496) );
  MUX2_X1 U14917 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n13224), .S(n16079), .Z(
        P3_U3495) );
  MUX2_X1 U14918 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n13225), .S(n16079), .Z(
        P3_U3494) );
  MUX2_X1 U14919 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13226), .S(n16079), .Z(
        P3_U3493) );
  MUX2_X1 U14920 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n13227), .S(n16079), .Z(
        P3_U3492) );
  MUX2_X1 U14921 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n13228), .S(n16079), .Z(
        P3_U3491) );
  INV_X1 U14922 ( .A(n13268), .ZN(n13254) );
  INV_X1 U14923 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n13655) );
  AOI22_X1 U14924 ( .A1(P3_REG1_REG_14__SCAN_IN), .A2(n13254), .B1(n13268), 
        .B2(n13655), .ZN(n13230) );
  NOR2_X1 U14925 ( .A1(n13231), .A2(n13230), .ZN(n13257) );
  AOI21_X1 U14926 ( .B1(n13231), .B2(n13230), .A(n13257), .ZN(n13256) );
  MUX2_X1 U14927 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n13357), .Z(n13232) );
  AND2_X1 U14928 ( .A1(n13268), .A2(n13232), .ZN(n13261) );
  NOR2_X1 U14929 ( .A1(n13268), .A2(n13232), .ZN(n13233) );
  OR2_X1 U14930 ( .A1(n13261), .A2(n13233), .ZN(n13239) );
  OR2_X1 U14931 ( .A1(n13235), .A2(n13234), .ZN(n13237) );
  NAND2_X1 U14932 ( .A1(n13237), .A2(n13236), .ZN(n13238) );
  NAND2_X1 U14933 ( .A1(n13239), .A2(n13238), .ZN(n13241) );
  INV_X1 U14934 ( .A(n13260), .ZN(n13240) );
  NAND3_X1 U14935 ( .A1(n13342), .A2(n13241), .A3(n13240), .ZN(n13244) );
  AOI21_X1 U14936 ( .B1(n16330), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n13242), 
        .ZN(n13243) );
  NAND2_X1 U14937 ( .A1(n13244), .A2(n13243), .ZN(n13253) );
  NOR2_X1 U14938 ( .A1(n8029), .A2(n13245), .ZN(n13247) );
  INV_X1 U14939 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13248) );
  AOI22_X1 U14940 ( .A1(P3_REG2_REG_14__SCAN_IN), .A2(n13254), .B1(n13268), 
        .B2(n13248), .ZN(n13249) );
  AOI21_X1 U14941 ( .B1(n13250), .B2(n13249), .A(n13267), .ZN(n13251) );
  NOR2_X1 U14942 ( .A1(n13251), .A2(n13368), .ZN(n13252) );
  AOI211_X1 U14943 ( .C1(n13370), .C2(n13254), .A(n13253), .B(n13252), .ZN(
        n13255) );
  OAI21_X1 U14944 ( .B1(n13256), .B2(n16328), .A(n13255), .ZN(P3_U3196) );
  INV_X1 U14945 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n13651) );
  AOI21_X1 U14946 ( .B1(n13651), .B2(n13258), .A(n13277), .ZN(n13275) );
  AOI21_X1 U14947 ( .B1(n16330), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n13259), 
        .ZN(n13266) );
  INV_X1 U14948 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13269) );
  MUX2_X1 U14949 ( .A(n13269), .B(n13651), .S(n13357), .Z(n13262) );
  NAND2_X1 U14950 ( .A1(n13263), .A2(n13262), .ZN(n13283) );
  OAI21_X1 U14951 ( .B1(n13263), .B2(n13262), .A(n13283), .ZN(n13264) );
  NAND2_X1 U14952 ( .A1(n13342), .A2(n13264), .ZN(n13265) );
  NAND2_X1 U14953 ( .A1(n13266), .A2(n13265), .ZN(n13273) );
  AOI21_X1 U14954 ( .B1(n13270), .B2(n13269), .A(n13293), .ZN(n13271) );
  NOR2_X1 U14955 ( .A1(n13271), .A2(n13368), .ZN(n13272) );
  AOI211_X1 U14956 ( .C1(n13370), .C2(n13292), .A(n13273), .B(n13272), .ZN(
        n13274) );
  OAI21_X1 U14957 ( .B1(n13275), .B2(n16328), .A(n13274), .ZN(P3_U3197) );
  NOR2_X1 U14958 ( .A1(n13292), .A2(n13276), .ZN(n13278) );
  INV_X1 U14959 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13647) );
  AOI22_X1 U14960 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n13296), .B1(n13316), 
        .B2(n13647), .ZN(n13279) );
  NOR2_X1 U14961 ( .A1(n13280), .A2(n13279), .ZN(n13302) );
  AOI21_X1 U14962 ( .B1(n13280), .B2(n13279), .A(n13302), .ZN(n13301) );
  INV_X1 U14963 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n16026) );
  OAI21_X1 U14964 ( .B1(n13345), .B2(n16026), .A(n13281), .ZN(n13290) );
  NAND2_X1 U14965 ( .A1(n13292), .A2(n13282), .ZN(n13284) );
  NAND2_X1 U14966 ( .A1(n13284), .A2(n13283), .ZN(n13288) );
  INV_X1 U14967 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13295) );
  MUX2_X1 U14968 ( .A(n13295), .B(n13647), .S(n13357), .Z(n13285) );
  NOR2_X1 U14969 ( .A1(n13296), .A2(n13285), .ZN(n13308) );
  AOI21_X1 U14970 ( .B1(n13296), .B2(n13285), .A(n13308), .ZN(n13286) );
  INV_X1 U14971 ( .A(n13286), .ZN(n13287) );
  NOR2_X1 U14972 ( .A1(n13287), .A2(n13288), .ZN(n13307) );
  AOI211_X1 U14973 ( .C1(n13288), .C2(n13287), .A(n13307), .B(n16327), .ZN(
        n13289) );
  AOI211_X1 U14974 ( .C1(n13370), .C2(n13296), .A(n13290), .B(n13289), .ZN(
        n13300) );
  AOI22_X1 U14975 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n13296), .B1(n13316), 
        .B2(n13295), .ZN(n13297) );
  AOI21_X1 U14976 ( .B1(n7524), .B2(n13297), .A(n13315), .ZN(n13298) );
  OR2_X1 U14977 ( .A1(n13298), .A2(n13368), .ZN(n13299) );
  OAI211_X1 U14978 ( .C1(n13301), .C2(n16328), .A(n13300), .B(n13299), .ZN(
        P3_U3198) );
  INV_X1 U14979 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13304) );
  AOI21_X1 U14980 ( .B1(P3_REG1_REG_16__SCAN_IN), .B2(n13316), .A(n13302), 
        .ZN(n13323) );
  AOI21_X1 U14981 ( .B1(n13304), .B2(n13303), .A(n13324), .ZN(n13322) );
  INV_X1 U14982 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n15967) );
  INV_X1 U14983 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13553) );
  MUX2_X1 U14984 ( .A(n13553), .B(n13304), .S(n13357), .Z(n13305) );
  NOR2_X1 U14985 ( .A1(n13328), .A2(n13305), .ZN(n13336) );
  AND2_X1 U14986 ( .A1(n13328), .A2(n13305), .ZN(n13306) );
  OR2_X1 U14987 ( .A1(n13336), .A2(n13306), .ZN(n13309) );
  NOR2_X1 U14988 ( .A1(n13308), .A2(n13307), .ZN(n13310) );
  NAND2_X1 U14989 ( .A1(n13309), .A2(n13310), .ZN(n13312) );
  NOR2_X1 U14990 ( .A1(n13310), .A2(n13309), .ZN(n13335) );
  NOR2_X1 U14991 ( .A1(n16327), .A2(n13335), .ZN(n13311) );
  NAND2_X1 U14992 ( .A1(n13312), .A2(n13311), .ZN(n13314) );
  OAI211_X1 U14993 ( .C1(n15967), .C2(n13345), .A(n13314), .B(n13313), .ZN(
        n13320) );
  XNOR2_X1 U14994 ( .A(n13327), .B(n13328), .ZN(n13317) );
  AOI21_X1 U14995 ( .B1(n13317), .B2(n13553), .A(n13329), .ZN(n13318) );
  NOR2_X1 U14996 ( .A1(n13318), .A2(n13368), .ZN(n13319) );
  AOI211_X1 U14997 ( .C1(n13370), .C2(n13328), .A(n13320), .B(n13319), .ZN(
        n13321) );
  OAI21_X1 U14998 ( .B1(n13322), .B2(n16328), .A(n13321), .ZN(P3_U3199) );
  NOR2_X1 U14999 ( .A1(n13328), .A2(n13323), .ZN(n13325) );
  INV_X1 U15000 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13639) );
  AOI22_X1 U15001 ( .A1(n13353), .A2(P3_REG1_REG_18__SCAN_IN), .B1(n13639), 
        .B2(n13364), .ZN(n13326) );
  AOI21_X1 U15002 ( .B1(n7510), .B2(n13326), .A(n13350), .ZN(n13349) );
  NOR2_X1 U15003 ( .A1(n13328), .A2(n13327), .ZN(n13330) );
  NAND2_X1 U15004 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n13364), .ZN(n13331) );
  OAI21_X1 U15005 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n13364), .A(n13331), 
        .ZN(n13332) );
  AOI21_X1 U15006 ( .B1(n13333), .B2(n13332), .A(n13363), .ZN(n13334) );
  NOR2_X1 U15007 ( .A1(n13334), .A2(n13368), .ZN(n13347) );
  INV_X1 U15008 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n16038) );
  NAND2_X1 U15009 ( .A1(n13370), .A2(n13353), .ZN(n13344) );
  INV_X1 U15010 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13337) );
  MUX2_X1 U15011 ( .A(n13337), .B(n13639), .S(n13357), .Z(n13338) );
  OAI21_X1 U15012 ( .B1(n13339), .B2(n13338), .A(n13355), .ZN(n13341) );
  AOI21_X1 U15013 ( .B1(n13342), .B2(n13341), .A(n13340), .ZN(n13343) );
  OAI211_X1 U15014 ( .C1(n16038), .C2(n13345), .A(n13344), .B(n13343), .ZN(
        n13346) );
  NOR2_X1 U15015 ( .A1(n13347), .A2(n13346), .ZN(n13348) );
  OAI21_X1 U15016 ( .B1(n13349), .B2(n16328), .A(n13348), .ZN(P3_U3200) );
  XNOR2_X1 U15017 ( .A(n13369), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13356) );
  XNOR2_X1 U15018 ( .A(n13351), .B(n13356), .ZN(n13371) );
  NAND2_X1 U15019 ( .A1(n13353), .A2(n13352), .ZN(n13354) );
  NAND2_X1 U15020 ( .A1(n13355), .A2(n13354), .ZN(n13361) );
  XNOR2_X1 U15021 ( .A(n13369), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n13365) );
  INV_X1 U15022 ( .A(n13365), .ZN(n13359) );
  INV_X1 U15023 ( .A(n13356), .ZN(n13358) );
  MUX2_X1 U15024 ( .A(n13359), .B(n13358), .S(n13357), .Z(n13360) );
  XNOR2_X1 U15025 ( .A(n13361), .B(n13360), .ZN(n13362) );
  NAND2_X1 U15026 ( .A1(n16330), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n13366) );
  NOR2_X1 U15027 ( .A1(n16405), .A2(n13372), .ZN(n13382) );
  INV_X1 U15028 ( .A(n13373), .ZN(n13374) );
  NAND2_X1 U15029 ( .A1(n13375), .A2(n13374), .ZN(n13665) );
  INV_X1 U15030 ( .A(n13665), .ZN(n13376) );
  NOR3_X1 U15031 ( .A1(n16414), .A2(n13382), .A3(n13376), .ZN(n13379) );
  NOR2_X1 U15032 ( .A1(n16411), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n13377) );
  OAI22_X1 U15033 ( .A1(n13667), .A2(n13587), .B1(n13379), .B2(n13377), .ZN(
        P3_U3202) );
  NOR2_X1 U15034 ( .A1(n16411), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n13378) );
  OAI22_X1 U15035 ( .A1(n13670), .A2(n13587), .B1(n13379), .B2(n13378), .ZN(
        P3_U3203) );
  NOR2_X1 U15036 ( .A1(n13380), .A2(n13587), .ZN(n13381) );
  AOI211_X1 U15037 ( .C1(n13492), .C2(P3_REG2_REG_29__SCAN_IN), .A(n13382), 
        .B(n13381), .ZN(n13385) );
  NAND2_X1 U15038 ( .A1(n13383), .A2(n13559), .ZN(n13384) );
  OAI211_X1 U15039 ( .C1(n7530), .C2(n16414), .A(n13385), .B(n13384), .ZN(
        P3_U3204) );
  OAI21_X1 U15040 ( .B1(n13388), .B2(n13387), .A(n13386), .ZN(n13596) );
  INV_X1 U15041 ( .A(n13596), .ZN(n13400) );
  AOI21_X1 U15042 ( .B1(n13403), .B2(n13391), .A(n13390), .ZN(n13395) );
  AOI22_X1 U15043 ( .A1(n13498), .A2(n13393), .B1(n13392), .B2(n13500), .ZN(
        n13394) );
  AOI22_X1 U15044 ( .A1(n13492), .A2(P3_REG2_REG_28__SCAN_IN), .B1(n16388), 
        .B2(n13396), .ZN(n13397) );
  OAI21_X1 U15045 ( .B1(n13673), .B2(n13587), .A(n13397), .ZN(n13398) );
  AOI21_X1 U15046 ( .B1(n13595), .B2(n16411), .A(n13398), .ZN(n13399) );
  OAI21_X1 U15047 ( .B1(n13400), .B2(n13590), .A(n13399), .ZN(P3_U3205) );
  OR2_X1 U15048 ( .A1(n13401), .A2(n13413), .ZN(n13402) );
  NAND2_X1 U15049 ( .A1(n13403), .A2(n13402), .ZN(n13407) );
  NAND2_X1 U15050 ( .A1(n13404), .A2(n13498), .ZN(n13405) );
  OAI21_X1 U15051 ( .B1(n13438), .B2(n16374), .A(n13405), .ZN(n13406) );
  AOI21_X1 U15052 ( .B1(n13407), .B2(n16377), .A(n13406), .ZN(n13600) );
  INV_X1 U15053 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n13410) );
  INV_X1 U15054 ( .A(n13408), .ZN(n13409) );
  OAI22_X1 U15055 ( .A1(n16411), .A2(n13410), .B1(n13409), .B2(n16405), .ZN(
        n13411) );
  AOI21_X1 U15056 ( .B1(n13412), .B2(n13555), .A(n13411), .ZN(n13418) );
  NAND2_X1 U15057 ( .A1(n13414), .A2(n13413), .ZN(n13415) );
  NAND2_X1 U15058 ( .A1(n13416), .A2(n13415), .ZN(n13598) );
  NAND2_X1 U15059 ( .A1(n13598), .A2(n13559), .ZN(n13417) );
  OAI211_X1 U15060 ( .C1(n13600), .C2(n16414), .A(n13418), .B(n13417), .ZN(
        P3_U3206) );
  INV_X1 U15061 ( .A(n13425), .ZN(n13419) );
  XNOR2_X1 U15062 ( .A(n13420), .B(n13419), .ZN(n13423) );
  OAI22_X1 U15063 ( .A1(n13453), .A2(n16374), .B1(n13421), .B2(n16372), .ZN(
        n13422) );
  AOI21_X1 U15064 ( .B1(n13423), .B2(n16377), .A(n13422), .ZN(n13606) );
  NAND2_X1 U15065 ( .A1(n13434), .A2(n13424), .ZN(n13426) );
  NAND2_X1 U15066 ( .A1(n13426), .A2(n13425), .ZN(n13428) );
  NAND2_X1 U15067 ( .A1(n13428), .A2(n13427), .ZN(n13604) );
  INV_X1 U15068 ( .A(n13604), .ZN(n13432) );
  AOI22_X1 U15069 ( .A1(n13492), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n13429), 
        .B2(n16388), .ZN(n13430) );
  OAI21_X1 U15070 ( .B1(n13681), .B2(n13587), .A(n13430), .ZN(n13431) );
  AOI21_X1 U15071 ( .B1(n13432), .B2(n13559), .A(n13431), .ZN(n13433) );
  OAI21_X1 U15072 ( .B1(n13492), .B2(n13606), .A(n13433), .ZN(P3_U3207) );
  OAI21_X1 U15073 ( .B1(n7514), .B2(n9083), .A(n13434), .ZN(n13610) );
  INV_X1 U15074 ( .A(n13610), .ZN(n13446) );
  INV_X1 U15075 ( .A(n13435), .ZN(n13436) );
  AOI211_X1 U15076 ( .C1(n9083), .C2(n13437), .A(n13582), .B(n13436), .ZN(
        n13441) );
  OAI22_X1 U15077 ( .A1(n13439), .A2(n16374), .B1(n13438), .B2(n16372), .ZN(
        n13440) );
  OR2_X1 U15078 ( .A1(n13441), .A2(n13440), .ZN(n13609) );
  AOI22_X1 U15079 ( .A1(n13492), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n16388), 
        .B2(n13442), .ZN(n13443) );
  OAI21_X1 U15080 ( .B1(n13685), .B2(n13587), .A(n13443), .ZN(n13444) );
  AOI21_X1 U15081 ( .B1(n13609), .B2(n16411), .A(n13444), .ZN(n13445) );
  OAI21_X1 U15082 ( .B1(n13446), .B2(n13590), .A(n13445), .ZN(P3_U3208) );
  XNOR2_X1 U15083 ( .A(n13448), .B(n13447), .ZN(n13688) );
  INV_X1 U15084 ( .A(n13688), .ZN(n13460) );
  INV_X1 U15085 ( .A(n13449), .ZN(n13450) );
  OAI22_X1 U15086 ( .A1(n13687), .A2(n13587), .B1(n13450), .B2(n16405), .ZN(
        n13459) );
  OAI21_X1 U15087 ( .B1(n7496), .B2(n13452), .A(n13451), .ZN(n13456) );
  OAI22_X1 U15088 ( .A1(n13454), .A2(n16374), .B1(n13453), .B2(n16372), .ZN(
        n13455) );
  AOI21_X1 U15089 ( .B1(n13456), .B2(n16377), .A(n13455), .ZN(n13457) );
  OAI21_X1 U15090 ( .B1(n13688), .B2(n16380), .A(n13457), .ZN(n13686) );
  MUX2_X1 U15091 ( .A(P3_REG2_REG_24__SCAN_IN), .B(n13686), .S(n16411), .Z(
        n13458) );
  AOI211_X1 U15092 ( .C1(n16390), .C2(n13460), .A(n13459), .B(n13458), .ZN(
        n13461) );
  INV_X1 U15093 ( .A(n13461), .ZN(P3_U3209) );
  OR2_X1 U15094 ( .A1(n13483), .A2(n13482), .ZN(n13485) );
  NAND2_X1 U15095 ( .A1(n13485), .A2(n13462), .ZN(n13463) );
  XNOR2_X1 U15096 ( .A(n13463), .B(n9080), .ZN(n13616) );
  INV_X1 U15097 ( .A(n13616), .ZN(n13474) );
  OAI211_X1 U15098 ( .C1(n13465), .C2(n9080), .A(n13464), .B(n16377), .ZN(
        n13468) );
  AOI22_X1 U15099 ( .A1(n13500), .A2(n13499), .B1(n13466), .B2(n13498), .ZN(
        n13467) );
  NAND2_X1 U15100 ( .A1(n13468), .A2(n13467), .ZN(n13615) );
  INV_X1 U15101 ( .A(n13469), .ZN(n13694) );
  AOI22_X1 U15102 ( .A1(n13492), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n16388), 
        .B2(n13470), .ZN(n13471) );
  OAI21_X1 U15103 ( .B1(n13694), .B2(n13587), .A(n13471), .ZN(n13472) );
  AOI21_X1 U15104 ( .B1(n13615), .B2(n16411), .A(n13472), .ZN(n13473) );
  OAI21_X1 U15105 ( .B1(n13474), .B2(n13590), .A(n13473), .ZN(P3_U3210) );
  XNOR2_X1 U15106 ( .A(n13476), .B(n13475), .ZN(n13477) );
  NAND2_X1 U15107 ( .A1(n13477), .A2(n16377), .ZN(n13481) );
  AOI22_X1 U15108 ( .A1(n13479), .A2(n13500), .B1(n13498), .B2(n13478), .ZN(
        n13480) );
  NAND2_X1 U15109 ( .A1(n13481), .A2(n13480), .ZN(n13619) );
  INV_X1 U15110 ( .A(n13619), .ZN(n13491) );
  NAND2_X1 U15111 ( .A1(n13483), .A2(n13482), .ZN(n13484) );
  AND2_X1 U15112 ( .A1(n13485), .A2(n13484), .ZN(n13620) );
  INV_X1 U15113 ( .A(n13486), .ZN(n13698) );
  AOI22_X1 U15114 ( .A1(n16414), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n16388), 
        .B2(n13487), .ZN(n13488) );
  OAI21_X1 U15115 ( .B1(n13698), .B2(n13587), .A(n13488), .ZN(n13489) );
  AOI21_X1 U15116 ( .B1(n13620), .B2(n13559), .A(n13489), .ZN(n13490) );
  OAI21_X1 U15117 ( .B1(n13492), .B2(n13491), .A(n13490), .ZN(P3_U3211) );
  OAI21_X1 U15118 ( .B1(n13495), .B2(n13494), .A(n13493), .ZN(n13505) );
  INV_X1 U15119 ( .A(n13505), .ZN(n13705) );
  INV_X1 U15120 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n13506) );
  XNOR2_X1 U15121 ( .A(n13497), .B(n13496), .ZN(n13503) );
  AOI22_X1 U15122 ( .A1(n13501), .A2(n13500), .B1(n13499), .B2(n13498), .ZN(
        n13502) );
  OAI21_X1 U15123 ( .B1(n13503), .B2(n13582), .A(n13502), .ZN(n13504) );
  AOI21_X1 U15124 ( .B1(n13505), .B2(n13661), .A(n13504), .ZN(n13699) );
  MUX2_X1 U15125 ( .A(n13506), .B(n13699), .S(n16411), .Z(n13509) );
  AOI22_X1 U15126 ( .A1(n13702), .A2(n13555), .B1(n16388), .B2(n13507), .ZN(
        n13508) );
  OAI211_X1 U15127 ( .C1(n13705), .C2(n13510), .A(n13509), .B(n13508), .ZN(
        P3_U3212) );
  OAI21_X1 U15128 ( .B1(n7597), .B2(n13512), .A(n13511), .ZN(n13630) );
  INV_X1 U15129 ( .A(n13630), .ZN(n13709) );
  AOI21_X1 U15130 ( .B1(n13513), .B2(n13512), .A(n13582), .ZN(n13517) );
  OAI22_X1 U15131 ( .A1(n13540), .A2(n16374), .B1(n13514), .B2(n16372), .ZN(
        n13515) );
  AOI21_X1 U15132 ( .B1(n13517), .B2(n13516), .A(n13515), .ZN(n13627) );
  INV_X1 U15133 ( .A(n13627), .ZN(n13521) );
  AOI22_X1 U15134 ( .A1(n16414), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n16388), 
        .B2(n13518), .ZN(n13519) );
  OAI21_X1 U15135 ( .B1(n13628), .B2(n13587), .A(n13519), .ZN(n13520) );
  AOI21_X1 U15136 ( .B1(n13521), .B2(n16411), .A(n13520), .ZN(n13522) );
  OAI21_X1 U15137 ( .B1(n13709), .B2(n13590), .A(n13522), .ZN(P3_U3213) );
  XOR2_X1 U15138 ( .A(n13525), .B(n13523), .Z(n13634) );
  INV_X1 U15139 ( .A(n13634), .ZN(n13532) );
  XOR2_X1 U15140 ( .A(n13525), .B(n13524), .Z(n13526) );
  OAI222_X1 U15141 ( .A1(n16374), .A2(n13548), .B1(n16372), .B2(n13527), .C1(
        n13582), .C2(n13526), .ZN(n13633) );
  AOI22_X1 U15142 ( .A1(n16414), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n16388), 
        .B2(n13528), .ZN(n13529) );
  OAI21_X1 U15143 ( .B1(n13713), .B2(n13587), .A(n13529), .ZN(n13530) );
  AOI21_X1 U15144 ( .B1(n13633), .B2(n16411), .A(n13530), .ZN(n13531) );
  OAI21_X1 U15145 ( .B1(n13590), .B2(n13532), .A(n13531), .ZN(P3_U3214) );
  XNOR2_X1 U15146 ( .A(n13533), .B(n13535), .ZN(n13638) );
  INV_X1 U15147 ( .A(n13638), .ZN(n13545) );
  INV_X1 U15148 ( .A(n13534), .ZN(n13546) );
  OAI21_X1 U15149 ( .B1(n13546), .B2(n13536), .A(n13535), .ZN(n13538) );
  AND2_X1 U15150 ( .A1(n13538), .A2(n13537), .ZN(n13539) );
  OAI222_X1 U15151 ( .A1(n16372), .A2(n13540), .B1(n16374), .B2(n13569), .C1(
        n13582), .C2(n13539), .ZN(n13637) );
  AOI22_X1 U15152 ( .A1(n16414), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n16388), 
        .B2(n13541), .ZN(n13542) );
  OAI21_X1 U15153 ( .B1(n13717), .B2(n13587), .A(n13542), .ZN(n13543) );
  AOI21_X1 U15154 ( .B1(n13637), .B2(n16411), .A(n13543), .ZN(n13544) );
  OAI21_X1 U15155 ( .B1(n13590), .B2(n13545), .A(n13544), .ZN(P3_U3215) );
  AOI211_X1 U15156 ( .C1(n13557), .C2(n13547), .A(n13582), .B(n13546), .ZN(
        n13550) );
  OAI22_X1 U15157 ( .A1(n13584), .A2(n16374), .B1(n13548), .B2(n16372), .ZN(
        n13549) );
  NOR2_X1 U15158 ( .A1(n13550), .A2(n13549), .ZN(n13643) );
  INV_X1 U15159 ( .A(n13644), .ZN(n13556) );
  INV_X1 U15160 ( .A(n13551), .ZN(n13552) );
  OAI22_X1 U15161 ( .A1(n16411), .A2(n13553), .B1(n13552), .B2(n16405), .ZN(
        n13554) );
  AOI21_X1 U15162 ( .B1(n13556), .B2(n13555), .A(n13554), .ZN(n13561) );
  XNOR2_X1 U15163 ( .A(n13558), .B(n13557), .ZN(n13641) );
  NAND2_X1 U15164 ( .A1(n13641), .A2(n13559), .ZN(n13560) );
  OAI211_X1 U15165 ( .C1(n13643), .C2(n16414), .A(n13561), .B(n13560), .ZN(
        P3_U3216) );
  XNOR2_X1 U15166 ( .A(n13562), .B(n13564), .ZN(n13646) );
  INV_X1 U15167 ( .A(n13646), .ZN(n13574) );
  NAND3_X1 U15168 ( .A1(n13577), .A2(n13564), .A3(n13563), .ZN(n13565) );
  AND2_X1 U15169 ( .A1(n13566), .A2(n13565), .ZN(n13567) );
  OAI222_X1 U15170 ( .A1(n16372), .A2(n13569), .B1(n16374), .B2(n13568), .C1(
        n13582), .C2(n13567), .ZN(n13645) );
  AOI22_X1 U15171 ( .A1(n16414), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n16388), 
        .B2(n13570), .ZN(n13571) );
  OAI21_X1 U15172 ( .B1(n13722), .B2(n13587), .A(n13571), .ZN(n13572) );
  AOI21_X1 U15173 ( .B1(n13645), .B2(n16411), .A(n13572), .ZN(n13573) );
  OAI21_X1 U15174 ( .B1(n13574), .B2(n13590), .A(n13573), .ZN(P3_U3217) );
  XNOR2_X1 U15175 ( .A(n13576), .B(n13575), .ZN(n13650) );
  INV_X1 U15176 ( .A(n13650), .ZN(n13591) );
  INV_X1 U15177 ( .A(n13577), .ZN(n13578) );
  AOI21_X1 U15178 ( .B1(n13580), .B2(n13579), .A(n13578), .ZN(n13581) );
  OAI222_X1 U15179 ( .A1(n16372), .A2(n13584), .B1(n16374), .B2(n13583), .C1(
        n13582), .C2(n13581), .ZN(n13649) );
  AOI22_X1 U15180 ( .A1(n16414), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n16388), 
        .B2(n13585), .ZN(n13586) );
  OAI21_X1 U15181 ( .B1(n13726), .B2(n13587), .A(n13586), .ZN(n13588) );
  AOI21_X1 U15182 ( .B1(n13649), .B2(n16411), .A(n13588), .ZN(n13589) );
  OAI21_X1 U15183 ( .B1(n13591), .B2(n13590), .A(n13589), .ZN(P3_U3218) );
  NOR2_X1 U15184 ( .A1(n16563), .A2(n13665), .ZN(n13593) );
  AOI21_X1 U15185 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n16563), .A(n13593), 
        .ZN(n13592) );
  OAI21_X1 U15186 ( .B1(n13667), .B2(n13657), .A(n13592), .ZN(P3_U3490) );
  AOI21_X1 U15187 ( .B1(P3_REG1_REG_30__SCAN_IN), .B2(n16563), .A(n13593), 
        .ZN(n13594) );
  OAI21_X1 U15188 ( .B1(n13670), .B2(n13657), .A(n13594), .ZN(P3_U3489) );
  INV_X1 U15189 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13597) );
  NAND2_X1 U15190 ( .A1(n13598), .A2(n16561), .ZN(n13599) );
  NAND2_X1 U15191 ( .A1(n13600), .A2(n13599), .ZN(n13674) );
  MUX2_X1 U15192 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n13674), .S(n16565), .Z(
        n13601) );
  INV_X1 U15193 ( .A(n13601), .ZN(n13602) );
  OAI21_X1 U15194 ( .B1(n13677), .B2(n13657), .A(n13602), .ZN(P3_U3486) );
  INV_X1 U15195 ( .A(n16561), .ZN(n13603) );
  NAND2_X1 U15196 ( .A1(n13606), .A2(n13605), .ZN(n13678) );
  MUX2_X1 U15197 ( .A(n13678), .B(P3_REG1_REG_26__SCAN_IN), .S(n16563), .Z(
        n13607) );
  INV_X1 U15198 ( .A(n13607), .ZN(n13608) );
  OAI21_X1 U15199 ( .B1(n13681), .B2(n13657), .A(n13608), .ZN(P3_U3485) );
  INV_X1 U15200 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13611) );
  AOI21_X1 U15201 ( .B1(n16561), .B2(n13610), .A(n13609), .ZN(n13682) );
  MUX2_X1 U15202 ( .A(n13611), .B(n13682), .S(n16565), .Z(n13612) );
  OAI21_X1 U15203 ( .B1(n13685), .B2(n13657), .A(n13612), .ZN(P3_U3484) );
  MUX2_X1 U15204 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13686), .S(n16565), .Z(
        n13614) );
  OAI22_X1 U15205 ( .A1(n13688), .A2(n13664), .B1(n13687), .B2(n13657), .ZN(
        n13613) );
  OR2_X1 U15206 ( .A1(n13614), .A2(n13613), .ZN(P3_U3483) );
  INV_X1 U15207 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13617) );
  AOI21_X1 U15208 ( .B1(n13616), .B2(n16561), .A(n13615), .ZN(n13691) );
  MUX2_X1 U15209 ( .A(n13617), .B(n13691), .S(n16565), .Z(n13618) );
  OAI21_X1 U15210 ( .B1(n13694), .B2(n13657), .A(n13618), .ZN(P3_U3482) );
  INV_X1 U15211 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13621) );
  AOI21_X1 U15212 ( .B1(n13620), .B2(n16561), .A(n13619), .ZN(n13695) );
  MUX2_X1 U15213 ( .A(n13621), .B(n13695), .S(n16565), .Z(n13622) );
  OAI21_X1 U15214 ( .B1(n13698), .B2(n13657), .A(n13622), .ZN(P3_U3481) );
  INV_X1 U15215 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13623) );
  MUX2_X1 U15216 ( .A(n13623), .B(n13699), .S(n16565), .Z(n13626) );
  NAND2_X1 U15217 ( .A1(n13702), .A2(n13624), .ZN(n13625) );
  OAI211_X1 U15218 ( .C1(n13705), .C2(n13664), .A(n13626), .B(n13625), .ZN(
        P3_U3480) );
  INV_X1 U15219 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13631) );
  OAI21_X1 U15220 ( .B1(n13628), .B2(n16558), .A(n13627), .ZN(n13629) );
  AOI21_X1 U15221 ( .B1(n13630), .B2(n13661), .A(n13629), .ZN(n13706) );
  MUX2_X1 U15222 ( .A(n13631), .B(n13706), .S(n16565), .Z(n13632) );
  OAI21_X1 U15223 ( .B1(n13709), .B2(n13664), .A(n13632), .ZN(P3_U3479) );
  INV_X1 U15224 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13635) );
  AOI21_X1 U15225 ( .B1(n13634), .B2(n16561), .A(n13633), .ZN(n13710) );
  MUX2_X1 U15226 ( .A(n13635), .B(n13710), .S(n16565), .Z(n13636) );
  OAI21_X1 U15227 ( .B1(n13713), .B2(n13657), .A(n13636), .ZN(P3_U3478) );
  AOI21_X1 U15228 ( .B1(n13638), .B2(n16561), .A(n13637), .ZN(n13714) );
  MUX2_X1 U15229 ( .A(n13639), .B(n13714), .S(n16565), .Z(n13640) );
  OAI21_X1 U15230 ( .B1(n13717), .B2(n13657), .A(n13640), .ZN(P3_U3477) );
  NAND2_X1 U15231 ( .A1(n13641), .A2(n16561), .ZN(n13642) );
  OAI211_X1 U15232 ( .C1(n16558), .C2(n13644), .A(n13643), .B(n13642), .ZN(
        n13718) );
  MUX2_X1 U15233 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13718), .S(n16565), .Z(
        P3_U3476) );
  AOI21_X1 U15234 ( .B1(n16561), .B2(n13646), .A(n13645), .ZN(n13719) );
  MUX2_X1 U15235 ( .A(n13647), .B(n13719), .S(n16565), .Z(n13648) );
  OAI21_X1 U15236 ( .B1(n13722), .B2(n13657), .A(n13648), .ZN(P3_U3475) );
  AOI21_X1 U15237 ( .B1(n16561), .B2(n13650), .A(n13649), .ZN(n13723) );
  MUX2_X1 U15238 ( .A(n13651), .B(n13723), .S(n16565), .Z(n13652) );
  OAI21_X1 U15239 ( .B1(n13657), .B2(n13726), .A(n13652), .ZN(P3_U3474) );
  AOI21_X1 U15240 ( .B1(n13654), .B2(n16561), .A(n13653), .ZN(n13727) );
  MUX2_X1 U15241 ( .A(n13655), .B(n13727), .S(n16565), .Z(n13656) );
  OAI21_X1 U15242 ( .B1(n13657), .B2(n13730), .A(n13656), .ZN(P3_U3473) );
  OAI21_X1 U15243 ( .B1(n13659), .B2(n16558), .A(n13658), .ZN(n13660) );
  AOI21_X1 U15244 ( .B1(n13662), .B2(n13661), .A(n13660), .ZN(n13732) );
  MUX2_X1 U15245 ( .A(n12296), .B(n13732), .S(n16565), .Z(n13663) );
  OAI21_X1 U15246 ( .B1(n13736), .B2(n13664), .A(n13663), .ZN(P3_U3472) );
  NOR2_X1 U15247 ( .A1(n16566), .A2(n13665), .ZN(n13668) );
  AOI21_X1 U15248 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n16566), .A(n13668), 
        .ZN(n13666) );
  OAI21_X1 U15249 ( .B1(n13667), .B2(n13731), .A(n13666), .ZN(P3_U3458) );
  AOI21_X1 U15250 ( .B1(P3_REG0_REG_30__SCAN_IN), .B2(n16566), .A(n13668), 
        .ZN(n13669) );
  OAI21_X1 U15251 ( .B1(n13670), .B2(n13731), .A(n13669), .ZN(P3_U3457) );
  INV_X1 U15252 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13671) );
  MUX2_X1 U15253 ( .A(n13671), .B(n7568), .S(n16569), .Z(n13672) );
  OAI21_X1 U15254 ( .B1(n13673), .B2(n13731), .A(n13672), .ZN(P3_U3455) );
  MUX2_X1 U15255 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n13674), .S(n16569), .Z(
        n13675) );
  INV_X1 U15256 ( .A(n13675), .ZN(n13676) );
  OAI21_X1 U15257 ( .B1(n13677), .B2(n13731), .A(n13676), .ZN(P3_U3454) );
  MUX2_X1 U15258 ( .A(n13678), .B(P3_REG0_REG_26__SCAN_IN), .S(n16566), .Z(
        n13679) );
  INV_X1 U15259 ( .A(n13679), .ZN(n13680) );
  OAI21_X1 U15260 ( .B1(n13681), .B2(n13731), .A(n13680), .ZN(P3_U3453) );
  INV_X1 U15261 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13683) );
  MUX2_X1 U15262 ( .A(n13683), .B(n13682), .S(n16569), .Z(n13684) );
  OAI21_X1 U15263 ( .B1(n13685), .B2(n13731), .A(n13684), .ZN(P3_U3452) );
  MUX2_X1 U15264 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n13686), .S(n16569), .Z(
        n13690) );
  OAI22_X1 U15265 ( .A1(n13688), .A2(n13735), .B1(n13687), .B2(n13731), .ZN(
        n13689) );
  OR2_X1 U15266 ( .A1(n13690), .A2(n13689), .ZN(P3_U3451) );
  INV_X1 U15267 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13692) );
  MUX2_X1 U15268 ( .A(n13692), .B(n13691), .S(n16569), .Z(n13693) );
  OAI21_X1 U15269 ( .B1(n13694), .B2(n13731), .A(n13693), .ZN(P3_U3450) );
  INV_X1 U15270 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13696) );
  MUX2_X1 U15271 ( .A(n13696), .B(n13695), .S(n16569), .Z(n13697) );
  OAI21_X1 U15272 ( .B1(n13698), .B2(n13731), .A(n13697), .ZN(P3_U3449) );
  INV_X1 U15273 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13700) );
  MUX2_X1 U15274 ( .A(n13700), .B(n13699), .S(n16569), .Z(n13704) );
  NAND2_X1 U15275 ( .A1(n13702), .A2(n13701), .ZN(n13703) );
  OAI211_X1 U15276 ( .C1(n13705), .C2(n13735), .A(n13704), .B(n13703), .ZN(
        P3_U3448) );
  INV_X1 U15277 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13707) );
  MUX2_X1 U15278 ( .A(n13707), .B(n13706), .S(n16569), .Z(n13708) );
  OAI21_X1 U15279 ( .B1(n13709), .B2(n13735), .A(n13708), .ZN(P3_U3447) );
  INV_X1 U15280 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13711) );
  MUX2_X1 U15281 ( .A(n13711), .B(n13710), .S(n16569), .Z(n13712) );
  OAI21_X1 U15282 ( .B1(n13713), .B2(n13731), .A(n13712), .ZN(P3_U3446) );
  INV_X1 U15283 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13715) );
  MUX2_X1 U15284 ( .A(n13715), .B(n13714), .S(n16569), .Z(n13716) );
  OAI21_X1 U15285 ( .B1(n13717), .B2(n13731), .A(n13716), .ZN(P3_U3444) );
  MUX2_X1 U15286 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n13718), .S(n16569), .Z(
        P3_U3441) );
  INV_X1 U15287 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13720) );
  MUX2_X1 U15288 ( .A(n13720), .B(n13719), .S(n16569), .Z(n13721) );
  OAI21_X1 U15289 ( .B1(n13722), .B2(n13731), .A(n13721), .ZN(P3_U3438) );
  INV_X1 U15290 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13724) );
  MUX2_X1 U15291 ( .A(n13724), .B(n13723), .S(n16569), .Z(n13725) );
  OAI21_X1 U15292 ( .B1(n13731), .B2(n13726), .A(n13725), .ZN(P3_U3435) );
  INV_X1 U15293 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n13728) );
  MUX2_X1 U15294 ( .A(n13728), .B(n13727), .S(n16569), .Z(n13729) );
  OAI21_X1 U15295 ( .B1(n13731), .B2(n13730), .A(n13729), .ZN(P3_U3432) );
  INV_X1 U15296 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n13733) );
  MUX2_X1 U15297 ( .A(n13733), .B(n13732), .S(n16569), .Z(n13734) );
  OAI21_X1 U15298 ( .B1(n13736), .B2(n13735), .A(n13734), .ZN(P3_U3429) );
  MUX2_X1 U15299 ( .A(P3_D_REG_1__SCAN_IN), .B(n13738), .S(n13737), .Z(
        P3_U3377) );
  NAND2_X1 U15300 ( .A1(n13740), .A2(n13739), .ZN(n13744) );
  OR4_X1 U15301 ( .A1(n13742), .A2(P3_IR_REG_30__SCAN_IN), .A3(n8638), .A4(
        P3_U3151), .ZN(n13743) );
  OAI211_X1 U15302 ( .C1(n13746), .C2(n13745), .A(n13744), .B(n13743), .ZN(
        P3_U3264) );
  INV_X1 U15303 ( .A(n13747), .ZN(n13749) );
  OAI222_X1 U15304 ( .A1(n13750), .A2(n13749), .B1(P3_U3151), .B2(n13748), 
        .C1(n15696), .C2(n13745), .ZN(P3_U3266) );
  MUX2_X1 U15305 ( .A(n13752), .B(n13751), .S(P3_STATE_REG_SCAN_IN), .Z(
        P3_U3294) );
  NAND2_X1 U15306 ( .A1(n14806), .A2(n14201), .ZN(n13754) );
  OR2_X1 U15307 ( .A1(n14202), .A2(n14808), .ZN(n13753) );
  INV_X1 U15308 ( .A(n14672), .ZN(n13870) );
  NAND2_X1 U15309 ( .A1(n14810), .A2(n14201), .ZN(n13756) );
  OR2_X1 U15310 ( .A1(n14202), .A2(n14811), .ZN(n13755) );
  XNOR2_X1 U15311 ( .A(n14677), .B(n13816), .ZN(n13842) );
  NAND2_X1 U15312 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .ZN(n13757) );
  INV_X1 U15313 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13930) );
  INV_X1 U15314 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13759) );
  NAND2_X1 U15315 ( .A1(n13829), .A2(n13759), .ZN(n13760) );
  NAND2_X1 U15316 ( .A1(n14494), .A2(n13843), .ZN(n13766) );
  INV_X1 U15317 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13763) );
  NAND2_X1 U15318 ( .A1(n13902), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n13762) );
  NAND2_X1 U15319 ( .A1(n14181), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n13761) );
  OAI211_X1 U15320 ( .C1(n13763), .C2(n14192), .A(n13762), .B(n13761), .ZN(
        n13764) );
  INV_X1 U15321 ( .A(n13764), .ZN(n13765) );
  NAND2_X1 U15322 ( .A1(n13766), .A2(n13765), .ZN(n14507) );
  NAND2_X1 U15323 ( .A1(n14507), .A2(n7458), .ZN(n13841) );
  NAND2_X1 U15324 ( .A1(n13767), .A2(n14201), .ZN(n13770) );
  OR2_X1 U15325 ( .A1(n14202), .A2(n13768), .ZN(n13769) );
  XNOR2_X1 U15326 ( .A(n14693), .B(n7463), .ZN(n13801) );
  INV_X1 U15327 ( .A(n13772), .ZN(n13774) );
  NAND2_X1 U15328 ( .A1(n13774), .A2(n13773), .ZN(n13775) );
  NAND2_X1 U15329 ( .A1(n13777), .A2(n14201), .ZN(n13780) );
  OR2_X1 U15330 ( .A1(n14202), .A2(n13778), .ZN(n13779) );
  XNOR2_X1 U15331 ( .A(n14708), .B(n13816), .ZN(n13781) );
  NAND2_X1 U15332 ( .A1(n14431), .A2(n7458), .ZN(n13782) );
  XNOR2_X1 U15333 ( .A(n13781), .B(n13782), .ZN(n13922) );
  INV_X1 U15334 ( .A(n13781), .ZN(n13784) );
  INV_X1 U15335 ( .A(n13782), .ZN(n13783) );
  NAND2_X1 U15336 ( .A1(n13784), .A2(n13783), .ZN(n13785) );
  NAND2_X1 U15337 ( .A1(n13786), .A2(n14201), .ZN(n13789) );
  OR2_X1 U15338 ( .A1(n14202), .A2(n13787), .ZN(n13788) );
  XNOR2_X1 U15339 ( .A(n14564), .B(n13816), .ZN(n13796) );
  XNOR2_X1 U15340 ( .A(n13803), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n14565) );
  NAND2_X1 U15341 ( .A1(n14565), .A2(n13843), .ZN(n13795) );
  INV_X1 U15342 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13792) );
  NAND2_X1 U15343 ( .A1(n14181), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n13791) );
  NAND2_X1 U15344 ( .A1(n13902), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n13790) );
  OAI211_X1 U15345 ( .C1(n13846), .C2(n13792), .A(n13791), .B(n13790), .ZN(
        n13793) );
  INV_X1 U15346 ( .A(n13793), .ZN(n13794) );
  NAND2_X1 U15347 ( .A1(n13795), .A2(n13794), .ZN(n14434) );
  NAND2_X1 U15348 ( .A1(n14434), .A2(n7458), .ZN(n13958) );
  INV_X1 U15349 ( .A(n13796), .ZN(n13797) );
  NOR2_X1 U15350 ( .A1(n13798), .A2(n13797), .ZN(n13799) );
  AOI21_X2 U15351 ( .B1(n13959), .B2(n13958), .A(n13799), .ZN(n13800) );
  INV_X1 U15352 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13962) );
  INV_X1 U15353 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13802) );
  OAI21_X1 U15354 ( .B1(n13803), .B2(n13962), .A(n13802), .ZN(n13804) );
  AND2_X1 U15355 ( .A1(n13804), .A2(n13817), .ZN(n14550) );
  NAND2_X1 U15356 ( .A1(n14550), .A2(n13843), .ZN(n13810) );
  INV_X1 U15357 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13807) );
  NAND2_X1 U15358 ( .A1(n13902), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n13806) );
  NAND2_X1 U15359 ( .A1(n14181), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n13805) );
  OAI211_X1 U15360 ( .C1(n13807), .C2(n14192), .A(n13806), .B(n13805), .ZN(
        n13808) );
  INV_X1 U15361 ( .A(n13808), .ZN(n13809) );
  NAND2_X1 U15362 ( .A1(n13810), .A2(n13809), .ZN(n14437) );
  NAND2_X1 U15363 ( .A1(n13812), .A2(n14201), .ZN(n13815) );
  OR2_X1 U15364 ( .A1(n14202), .A2(n13813), .ZN(n13814) );
  XNOR2_X1 U15365 ( .A(n14688), .B(n13816), .ZN(n13927) );
  INV_X1 U15366 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13942) );
  NAND2_X1 U15367 ( .A1(n13817), .A2(n13942), .ZN(n13818) );
  NAND2_X1 U15368 ( .A1(n13827), .A2(n13818), .ZN(n14535) );
  OR2_X1 U15369 ( .A1(n14535), .A2(n10059), .ZN(n13823) );
  INV_X1 U15370 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n14534) );
  NAND2_X1 U15371 ( .A1(n13902), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n13820) );
  NAND2_X1 U15372 ( .A1(n14181), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n13819) );
  OAI211_X1 U15373 ( .C1(n14534), .C2(n14192), .A(n13820), .B(n13819), .ZN(
        n13821) );
  INV_X1 U15374 ( .A(n13821), .ZN(n13822) );
  NAND2_X1 U15375 ( .A1(n13823), .A2(n13822), .ZN(n14506) );
  NAND2_X1 U15376 ( .A1(n14506), .A2(n7458), .ZN(n13824) );
  NOR2_X1 U15377 ( .A1(n13927), .A2(n13824), .ZN(n13825) );
  AOI21_X1 U15378 ( .B1(n13927), .B2(n13824), .A(n13825), .ZN(n13939) );
  OR2_X1 U15379 ( .A1(n14202), .A2(n14817), .ZN(n13826) );
  XNOR2_X1 U15380 ( .A(n14760), .B(n7463), .ZN(n13835) );
  NAND2_X1 U15381 ( .A1(n13827), .A2(n13930), .ZN(n13828) );
  AND2_X1 U15382 ( .A1(n13829), .A2(n13828), .ZN(n14517) );
  NAND2_X1 U15383 ( .A1(n14517), .A2(n13843), .ZN(n13834) );
  INV_X1 U15384 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n14519) );
  NAND2_X1 U15385 ( .A1(n13902), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n13831) );
  NAND2_X1 U15386 ( .A1(n14181), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n13830) );
  OAI211_X1 U15387 ( .C1(n14519), .C2(n14192), .A(n13831), .B(n13830), .ZN(
        n13832) );
  INV_X1 U15388 ( .A(n13832), .ZN(n13833) );
  NAND2_X1 U15389 ( .A1(n13834), .A2(n13833), .ZN(n14442) );
  AND2_X1 U15390 ( .A1(n14442), .A2(n7458), .ZN(n13836) );
  NAND2_X1 U15391 ( .A1(n13835), .A2(n13836), .ZN(n13839) );
  INV_X1 U15392 ( .A(n13835), .ZN(n13968) );
  INV_X1 U15393 ( .A(n13836), .ZN(n13837) );
  NAND2_X1 U15394 ( .A1(n13968), .A2(n13837), .ZN(n13838) );
  NAND2_X1 U15395 ( .A1(n13839), .A2(n13838), .ZN(n13926) );
  INV_X1 U15396 ( .A(n13839), .ZN(n13840) );
  XNOR2_X1 U15397 ( .A(n13842), .B(n13841), .ZN(n13971) );
  XNOR2_X1 U15398 ( .A(n14672), .B(n13816), .ZN(n13851) );
  XNOR2_X1 U15399 ( .A(n13857), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n14477) );
  NAND2_X1 U15400 ( .A1(n14477), .A2(n13843), .ZN(n13849) );
  INV_X1 U15401 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n14479) );
  NAND2_X1 U15402 ( .A1(n13902), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n13845) );
  NAND2_X1 U15403 ( .A1(n14181), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n13844) );
  OAI211_X1 U15404 ( .C1(n14479), .C2(n14192), .A(n13845), .B(n13844), .ZN(
        n13847) );
  INV_X1 U15405 ( .A(n13847), .ZN(n13848) );
  NAND2_X1 U15406 ( .A1(n14447), .A2(n7458), .ZN(n13850) );
  NOR2_X1 U15407 ( .A1(n13851), .A2(n13850), .ZN(n13893) );
  AOI21_X1 U15408 ( .B1(n13851), .B2(n13850), .A(n13893), .ZN(n13852) );
  NAND2_X1 U15409 ( .A1(n13853), .A2(n13852), .ZN(n13895) );
  OAI211_X1 U15410 ( .C1(n13853), .C2(n13852), .A(n13895), .B(n13977), .ZN(
        n13869) );
  INV_X1 U15411 ( .A(n13857), .ZN(n13855) );
  AND2_X1 U15412 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n13854) );
  NAND2_X1 U15413 ( .A1(n13855), .A2(n13854), .ZN(n14420) );
  INV_X1 U15414 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n13865) );
  INV_X1 U15415 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n13856) );
  OAI21_X1 U15416 ( .B1(n13857), .B2(n13865), .A(n13856), .ZN(n13858) );
  NAND2_X1 U15417 ( .A1(n14420), .A2(n13858), .ZN(n14463) );
  OR2_X1 U15418 ( .A1(n14463), .A2(n10059), .ZN(n13863) );
  INV_X1 U15419 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n14462) );
  NAND2_X1 U15420 ( .A1(n14181), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n13860) );
  NAND2_X1 U15421 ( .A1(n13902), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n13859) );
  OAI211_X1 U15422 ( .C1(n14462), .C2(n14192), .A(n13860), .B(n13859), .ZN(
        n13861) );
  INV_X1 U15423 ( .A(n13861), .ZN(n13862) );
  INV_X1 U15424 ( .A(n14412), .ZN(n13864) );
  INV_X1 U15425 ( .A(n14507), .ZN(n14407) );
  OAI22_X1 U15426 ( .A1(n13864), .A2(n14374), .B1(n14407), .B2(n13941), .ZN(
        n14471) );
  INV_X1 U15427 ( .A(n14477), .ZN(n13866) );
  OAI22_X1 U15428 ( .A1(n13866), .A2(n13943), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13865), .ZN(n13867) );
  AOI21_X1 U15429 ( .B1(n14471), .B2(n13945), .A(n13867), .ZN(n13868) );
  OAI211_X1 U15430 ( .C1(n13870), .C2(n13966), .A(n13869), .B(n13868), .ZN(
        P2_U3186) );
  AOI22_X1 U15431 ( .A1(n13871), .A2(n13977), .B1(n13957), .B2(n14437), .ZN(
        n13880) );
  INV_X1 U15432 ( .A(n13872), .ZN(n13879) );
  NAND2_X1 U15433 ( .A1(n14506), .A2(n14614), .ZN(n13874) );
  NAND2_X1 U15434 ( .A1(n14434), .A2(n14613), .ZN(n13873) );
  NAND2_X1 U15435 ( .A1(n13874), .A2(n13873), .ZN(n14544) );
  INV_X1 U15436 ( .A(n14544), .ZN(n13876) );
  AOI22_X1 U15437 ( .A1(n14550), .A2(n13972), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13875) );
  OAI21_X1 U15438 ( .B1(n13876), .B2(n13975), .A(n13875), .ZN(n13877) );
  AOI21_X1 U15439 ( .B1(n14693), .B2(n13952), .A(n13877), .ZN(n13878) );
  OAI21_X1 U15440 ( .B1(n13880), .B2(n13879), .A(n13878), .ZN(P2_U3188) );
  OAI21_X1 U15441 ( .B1(n13882), .B2(n13887), .A(n13881), .ZN(n13883) );
  NAND2_X1 U15442 ( .A1(n13883), .A2(n13977), .ZN(n13892) );
  INV_X1 U15443 ( .A(n14615), .ZN(n14392) );
  NOR2_X1 U15444 ( .A1(n13933), .A2(n14392), .ZN(n13885) );
  NAND2_X1 U15445 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3088), .ZN(n14365)
         );
  OAI21_X1 U15446 ( .B1(n13943), .B2(n14623), .A(n14365), .ZN(n13884) );
  AOI211_X1 U15447 ( .C1(n14621), .C2(n13952), .A(n13885), .B(n13884), .ZN(
        n13891) );
  NOR3_X1 U15448 ( .A1(n13887), .A2(n13886), .A3(n13967), .ZN(n13889) );
  OAI21_X1 U15449 ( .B1(n13889), .B2(n13888), .A(n14612), .ZN(n13890) );
  NAND3_X1 U15450 ( .A1(n13892), .A2(n13891), .A3(n13890), .ZN(P2_U3191) );
  INV_X1 U15451 ( .A(n13893), .ZN(n13894) );
  NAND2_X1 U15452 ( .A1(n13895), .A2(n13894), .ZN(n13901) );
  NAND2_X1 U15453 ( .A1(n14802), .A2(n14201), .ZN(n13897) );
  OR2_X1 U15454 ( .A1(n14202), .A2(n14805), .ZN(n13896) );
  NAND2_X1 U15455 ( .A1(n14412), .A2(n7458), .ZN(n13898) );
  XNOR2_X1 U15456 ( .A(n13898), .B(n7463), .ZN(n13899) );
  XNOR2_X1 U15457 ( .A(n14465), .B(n13899), .ZN(n13900) );
  XNOR2_X1 U15458 ( .A(n13901), .B(n13900), .ZN(n13916) );
  NAND2_X1 U15459 ( .A1(n14447), .A2(n14613), .ZN(n13910) );
  OR2_X1 U15460 ( .A1(n14420), .A2(n10059), .ZN(n13908) );
  INV_X1 U15461 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n13905) );
  NAND2_X1 U15462 ( .A1(n13902), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n13904) );
  NAND2_X1 U15463 ( .A1(n14181), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n13903) );
  OAI211_X1 U15464 ( .C1(n13905), .C2(n14192), .A(n13904), .B(n13903), .ZN(
        n13906) );
  INV_X1 U15465 ( .A(n13906), .ZN(n13907) );
  NAND2_X1 U15466 ( .A1(n13908), .A2(n13907), .ZN(n14304) );
  NAND2_X1 U15467 ( .A1(n14304), .A2(n14614), .ZN(n13909) );
  AND2_X1 U15468 ( .A1(n13910), .A2(n13909), .ZN(n14455) );
  INV_X1 U15469 ( .A(n14463), .ZN(n13911) );
  AOI22_X1 U15470 ( .A1(n13911), .A2(n13972), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13912) );
  OAI21_X1 U15471 ( .B1(n14455), .B2(n13975), .A(n13912), .ZN(n13913) );
  AOI21_X1 U15472 ( .B1(n14465), .B2(n13952), .A(n13913), .ZN(n13914) );
  OAI21_X1 U15473 ( .B1(n13916), .B2(n13915), .A(n13914), .ZN(P2_U3192) );
  AOI22_X1 U15474 ( .A1(n14434), .A2(n14614), .B1(n14613), .B2(n14615), .ZN(
        n14575) );
  INV_X1 U15475 ( .A(n14581), .ZN(n13917) );
  AOI22_X1 U15476 ( .A1(n13972), .A2(n13917), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13918) );
  OAI21_X1 U15477 ( .B1(n14575), .B2(n13975), .A(n13918), .ZN(n13924) );
  INV_X1 U15478 ( .A(n13919), .ZN(n13920) );
  AOI211_X1 U15479 ( .C1(n13922), .C2(n13921), .A(n13915), .B(n13920), .ZN(
        n13923) );
  AOI211_X1 U15480 ( .C1(n14708), .C2(n13952), .A(n13924), .B(n13923), .ZN(
        n13925) );
  INV_X1 U15481 ( .A(n13925), .ZN(P2_U3195) );
  AOI21_X1 U15482 ( .B1(n13938), .B2(n13926), .A(n13915), .ZN(n13929) );
  INV_X1 U15483 ( .A(n14506), .ZN(n14404) );
  NOR3_X1 U15484 ( .A1(n13927), .A2(n14404), .A3(n13967), .ZN(n13928) );
  NOR2_X1 U15485 ( .A1(n13929), .A2(n13928), .ZN(n13937) );
  INV_X1 U15486 ( .A(n14517), .ZN(n13931) );
  OAI22_X1 U15487 ( .A1(n13931), .A2(n13943), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13930), .ZN(n13935) );
  OAI22_X1 U15488 ( .A1(n14407), .A2(n13933), .B1(n14404), .B2(n13932), .ZN(
        n13934) );
  AOI211_X1 U15489 ( .C1(n14760), .C2(n13952), .A(n13935), .B(n13934), .ZN(
        n13936) );
  OAI21_X1 U15490 ( .B1(n13937), .B2(n13970), .A(n13936), .ZN(P2_U3197) );
  INV_X1 U15491 ( .A(n14688), .ZN(n14533) );
  OAI211_X1 U15492 ( .C1(n13940), .C2(n13939), .A(n13938), .B(n13977), .ZN(
        n13947) );
  INV_X1 U15493 ( .A(n14437), .ZN(n14402) );
  OAI22_X1 U15494 ( .A1(n7855), .A2(n14374), .B1(n14402), .B2(n13941), .ZN(
        n14531) );
  OAI22_X1 U15495 ( .A1(n14535), .A2(n13943), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13942), .ZN(n13944) );
  AOI21_X1 U15496 ( .B1(n14531), .B2(n13945), .A(n13944), .ZN(n13946) );
  OAI211_X1 U15497 ( .C1(n14533), .C2(n13966), .A(n13947), .B(n13946), .ZN(
        P2_U3201) );
  INV_X1 U15498 ( .A(n13948), .ZN(n13949) );
  AOI22_X1 U15499 ( .A1(n13950), .A2(n14321), .B1(n13949), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n13956) );
  AOI21_X1 U15500 ( .B1(n14323), .B2(n7458), .A(n13915), .ZN(n13953) );
  OAI21_X1 U15501 ( .B1(n13953), .B2(n13952), .A(n13951), .ZN(n13955) );
  NAND3_X1 U15502 ( .A1(n13957), .A2(n14323), .A3(n13987), .ZN(n13954) );
  NAND3_X1 U15503 ( .A1(n13956), .A2(n13955), .A3(n13954), .ZN(P2_U3204) );
  NAND2_X1 U15504 ( .A1(n13957), .A2(n14434), .ZN(n13961) );
  NAND2_X1 U15505 ( .A1(n13958), .A2(n13977), .ZN(n13960) );
  MUX2_X1 U15506 ( .A(n13961), .B(n13960), .S(n13959), .Z(n13965) );
  AOI22_X1 U15507 ( .A1(n14437), .A2(n14614), .B1(n14613), .B2(n14431), .ZN(
        n14559) );
  OAI22_X1 U15508 ( .A1(n14559), .A2(n13975), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13962), .ZN(n13963) );
  AOI21_X1 U15509 ( .B1(n14565), .B2(n13972), .A(n13963), .ZN(n13964) );
  OAI211_X1 U15510 ( .C1(n14769), .C2(n13966), .A(n13965), .B(n13964), .ZN(
        P2_U3207) );
  NOR3_X1 U15511 ( .A1(n13968), .A2(n7855), .A3(n13967), .ZN(n13969) );
  AOI21_X1 U15512 ( .B1(n13970), .B2(n13977), .A(n13969), .ZN(n13981) );
  INV_X1 U15513 ( .A(n13971), .ZN(n13980) );
  AOI22_X1 U15514 ( .A1(n14447), .A2(n14614), .B1(n14613), .B2(n14442), .ZN(
        n14488) );
  NAND2_X1 U15515 ( .A1(n14677), .A2(n13952), .ZN(n13974) );
  AOI22_X1 U15516 ( .A1(n14494), .A2(n13972), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13973) );
  OAI211_X1 U15517 ( .C1(n14488), .C2(n13975), .A(n13974), .B(n13973), .ZN(
        n13976) );
  AOI21_X1 U15518 ( .B1(n13978), .B2(n13977), .A(n13976), .ZN(n13979) );
  OAI21_X1 U15519 ( .B1(n13981), .B2(n13980), .A(n13979), .ZN(P2_U3212) );
  NAND2_X1 U15520 ( .A1(n13983), .A2(n10126), .ZN(n13985) );
  NAND2_X1 U15521 ( .A1(n13987), .A2(n13986), .ZN(n13989) );
  NAND3_X1 U15522 ( .A1(n13989), .A2(n13988), .A3(n14217), .ZN(n13990) );
  NAND2_X1 U15523 ( .A1(n13991), .A2(n13990), .ZN(n13997) );
  NAND2_X1 U15524 ( .A1(n14321), .A2(n14004), .ZN(n13998) );
  NAND2_X1 U15525 ( .A1(n14207), .A2(n13992), .ZN(n13999) );
  NAND2_X1 U15526 ( .A1(n13998), .A2(n13999), .ZN(n13993) );
  NAND2_X1 U15527 ( .A1(n14321), .A2(n14212), .ZN(n13994) );
  INV_X1 U15528 ( .A(n13997), .ZN(n14001) );
  AND2_X1 U15529 ( .A1(n13999), .A2(n13998), .ZN(n14000) );
  NAND2_X1 U15530 ( .A1(n14001), .A2(n14000), .ZN(n14002) );
  INV_X1 U15531 ( .A(n14004), .ZN(n14217) );
  NAND2_X1 U15532 ( .A1(n14320), .A2(n14207), .ZN(n14007) );
  NAND2_X1 U15533 ( .A1(n14113), .A2(n14005), .ZN(n14006) );
  NAND2_X1 U15534 ( .A1(n14007), .A2(n14006), .ZN(n14012) );
  NAND2_X1 U15535 ( .A1(n14011), .A2(n14012), .ZN(n14010) );
  NAND2_X1 U15536 ( .A1(n14320), .A2(n14004), .ZN(n14008) );
  OAI21_X1 U15537 ( .B1(n14113), .B2(n16418), .A(n14008), .ZN(n14009) );
  NAND2_X1 U15538 ( .A1(n14010), .A2(n14009), .ZN(n14016) );
  INV_X1 U15539 ( .A(n14011), .ZN(n14014) );
  INV_X1 U15540 ( .A(n14012), .ZN(n14013) );
  NAND2_X1 U15541 ( .A1(n14014), .A2(n14013), .ZN(n14015) );
  NAND2_X1 U15542 ( .A1(n14019), .A2(n14238), .ZN(n14018) );
  NAND2_X1 U15543 ( .A1(n14319), .A2(n14113), .ZN(n14017) );
  NAND2_X1 U15544 ( .A1(n14018), .A2(n14017), .ZN(n14021) );
  INV_X1 U15545 ( .A(n14004), .ZN(n14207) );
  AOI22_X1 U15546 ( .A1(n14113), .A2(n14019), .B1(n14319), .B2(n14238), .ZN(
        n14020) );
  NAND2_X1 U15547 ( .A1(n14026), .A2(n14113), .ZN(n14025) );
  INV_X1 U15548 ( .A(n14004), .ZN(n14212) );
  NAND2_X1 U15549 ( .A1(n14318), .A2(n14238), .ZN(n14024) );
  NAND2_X1 U15550 ( .A1(n14026), .A2(n14238), .ZN(n14027) );
  OAI21_X1 U15551 ( .B1(n14028), .B2(n14238), .A(n14027), .ZN(n14029) );
  NAND2_X1 U15552 ( .A1(n14032), .A2(n14238), .ZN(n14031) );
  NAND2_X1 U15553 ( .A1(n14317), .A2(n14004), .ZN(n14030) );
  NAND2_X1 U15554 ( .A1(n14031), .A2(n14030), .ZN(n14034) );
  AOI22_X1 U15555 ( .A1(n14032), .A2(n14113), .B1(n14238), .B2(n14317), .ZN(
        n14033) );
  NAND2_X1 U15556 ( .A1(n14038), .A2(n14206), .ZN(n14037) );
  NAND2_X1 U15557 ( .A1(n14316), .A2(n7451), .ZN(n14036) );
  NAND2_X1 U15558 ( .A1(n14037), .A2(n14036), .ZN(n14040) );
  AOI22_X1 U15559 ( .A1(n14038), .A2(n14176), .B1(n14206), .B2(n14316), .ZN(
        n14039) );
  NAND2_X1 U15560 ( .A1(n14044), .A2(n7452), .ZN(n14043) );
  NAND2_X1 U15561 ( .A1(n14315), .A2(n14004), .ZN(n14042) );
  NAND2_X1 U15562 ( .A1(n14043), .A2(n14042), .ZN(n14048) );
  NAND2_X1 U15563 ( .A1(n14044), .A2(n14004), .ZN(n14045) );
  OAI21_X1 U15564 ( .B1(n14206), .B2(n14046), .A(n14045), .ZN(n14047) );
  INV_X1 U15565 ( .A(n14048), .ZN(n14049) );
  NAND2_X1 U15566 ( .A1(n14052), .A2(n14206), .ZN(n14051) );
  NAND2_X1 U15567 ( .A1(n14314), .A2(n7452), .ZN(n14050) );
  NAND2_X1 U15568 ( .A1(n14051), .A2(n14050), .ZN(n14054) );
  AOI22_X1 U15569 ( .A1(n14052), .A2(n14176), .B1(n14206), .B2(n14314), .ZN(
        n14053) );
  AOI21_X1 U15570 ( .B1(n14055), .B2(n14054), .A(n14053), .ZN(n14057) );
  NOR2_X1 U15571 ( .A1(n14055), .A2(n14054), .ZN(n14056) );
  NAND2_X1 U15572 ( .A1(n14060), .A2(n14176), .ZN(n14059) );
  NAND2_X1 U15573 ( .A1(n14313), .A2(n14206), .ZN(n14058) );
  NAND2_X1 U15574 ( .A1(n14059), .A2(n14058), .ZN(n14064) );
  NAND2_X1 U15575 ( .A1(n14060), .A2(n14206), .ZN(n14061) );
  OAI21_X1 U15576 ( .B1(n14206), .B2(n14062), .A(n14061), .ZN(n14063) );
  INV_X1 U15577 ( .A(n14064), .ZN(n14065) );
  NAND2_X1 U15578 ( .A1(n14068), .A2(n14206), .ZN(n14067) );
  NAND2_X1 U15579 ( .A1(n14312), .A2(n14176), .ZN(n14066) );
  NAND2_X1 U15580 ( .A1(n14067), .A2(n14066), .ZN(n14070) );
  AOI22_X1 U15581 ( .A1(n14068), .A2(n7452), .B1(n14206), .B2(n14312), .ZN(
        n14069) );
  NAND2_X1 U15582 ( .A1(n14072), .A2(n7522), .ZN(n14079) );
  NAND2_X1 U15583 ( .A1(n14075), .A2(n14176), .ZN(n14074) );
  NAND2_X1 U15584 ( .A1(n14311), .A2(n14206), .ZN(n14073) );
  NAND2_X1 U15585 ( .A1(n14074), .A2(n14073), .ZN(n14080) );
  NAND2_X1 U15586 ( .A1(n14075), .A2(n14206), .ZN(n14076) );
  OAI21_X1 U15587 ( .B1(n14206), .B2(n14077), .A(n14076), .ZN(n14078) );
  NAND2_X1 U15588 ( .A1(n14084), .A2(n14206), .ZN(n14083) );
  NAND2_X1 U15589 ( .A1(n14310), .A2(n7452), .ZN(n14082) );
  NAND2_X1 U15590 ( .A1(n14083), .A2(n14082), .ZN(n14086) );
  AOI22_X1 U15591 ( .A1(n14084), .A2(n14176), .B1(n14206), .B2(n14310), .ZN(
        n14085) );
  NAND2_X1 U15592 ( .A1(n14089), .A2(n14176), .ZN(n14088) );
  NAND2_X1 U15593 ( .A1(n14309), .A2(n14206), .ZN(n14087) );
  NAND2_X1 U15594 ( .A1(n14088), .A2(n14087), .ZN(n14095) );
  NAND2_X1 U15595 ( .A1(n14094), .A2(n14095), .ZN(n14093) );
  NAND2_X1 U15596 ( .A1(n14089), .A2(n14206), .ZN(n14090) );
  OAI21_X1 U15597 ( .B1(n14206), .B2(n14091), .A(n14090), .ZN(n14092) );
  NAND2_X1 U15598 ( .A1(n14093), .A2(n14092), .ZN(n14099) );
  INV_X1 U15599 ( .A(n14094), .ZN(n14097) );
  NAND2_X1 U15600 ( .A1(n14097), .A2(n14096), .ZN(n14098) );
  NAND2_X1 U15601 ( .A1(n14102), .A2(n14206), .ZN(n14101) );
  NAND2_X1 U15602 ( .A1(n14308), .A2(n7452), .ZN(n14100) );
  NAND2_X1 U15603 ( .A1(n14101), .A2(n14100), .ZN(n14104) );
  AOI22_X1 U15604 ( .A1(n14102), .A2(n14176), .B1(n14206), .B2(n14308), .ZN(
        n14103) );
  NAND2_X1 U15605 ( .A1(n14108), .A2(n14176), .ZN(n14107) );
  NAND2_X1 U15606 ( .A1(n14307), .A2(n14206), .ZN(n14106) );
  NAND2_X1 U15607 ( .A1(n14107), .A2(n14106), .ZN(n14110) );
  AOI22_X1 U15608 ( .A1(n14108), .A2(n14206), .B1(n14176), .B2(n14307), .ZN(
        n14109) );
  AOI21_X1 U15609 ( .B1(n14111), .B2(n14110), .A(n14109), .ZN(n14112) );
  NAND2_X1 U15610 ( .A1(n14789), .A2(n14206), .ZN(n14115) );
  NAND2_X1 U15611 ( .A1(n14306), .A2(n14176), .ZN(n14114) );
  NAND2_X1 U15612 ( .A1(n14115), .A2(n14114), .ZN(n14119) );
  NAND2_X1 U15613 ( .A1(n14789), .A2(n7452), .ZN(n14117) );
  NAND2_X1 U15614 ( .A1(n14306), .A2(n14206), .ZN(n14116) );
  NAND2_X1 U15615 ( .A1(n14117), .A2(n14116), .ZN(n14118) );
  NAND2_X1 U15616 ( .A1(n14728), .A2(n14176), .ZN(n14121) );
  NAND2_X1 U15617 ( .A1(n14305), .A2(n14206), .ZN(n14120) );
  NAND2_X1 U15618 ( .A1(n14121), .A2(n14120), .ZN(n14126) );
  NAND2_X1 U15619 ( .A1(n14125), .A2(n14126), .ZN(n14124) );
  AOI22_X1 U15620 ( .A1(n14728), .A2(n14206), .B1(n14176), .B2(n14305), .ZN(
        n14122) );
  NAND2_X1 U15621 ( .A1(n14426), .A2(n14206), .ZN(n14129) );
  NAND2_X1 U15622 ( .A1(n14612), .A2(n7452), .ZN(n14128) );
  NAND2_X1 U15623 ( .A1(n14426), .A2(n14176), .ZN(n14130) );
  OAI21_X1 U15624 ( .B1(n14386), .B2(n7452), .A(n14130), .ZN(n14131) );
  NAND2_X1 U15625 ( .A1(n14621), .A2(n7452), .ZN(n14133) );
  NAND2_X1 U15626 ( .A1(n14428), .A2(n14206), .ZN(n14132) );
  NAND2_X1 U15627 ( .A1(n14133), .A2(n14132), .ZN(n14135) );
  AOI22_X1 U15628 ( .A1(n14621), .A2(n14206), .B1(n7452), .B2(n14428), .ZN(
        n14134) );
  AOI21_X1 U15629 ( .B1(n14136), .B2(n14135), .A(n14134), .ZN(n14137) );
  AND2_X1 U15630 ( .A1(n14615), .A2(n14176), .ZN(n14138) );
  AOI21_X1 U15631 ( .B1(n14593), .B2(n14206), .A(n14138), .ZN(n14139) );
  INV_X1 U15632 ( .A(n14139), .ZN(n14140) );
  NAND2_X1 U15633 ( .A1(n14593), .A2(n14176), .ZN(n14141) );
  OAI21_X1 U15634 ( .B1(n14392), .B2(n14176), .A(n14141), .ZN(n14142) );
  NAND2_X1 U15635 ( .A1(n14708), .A2(n7452), .ZN(n14144) );
  NAND2_X1 U15636 ( .A1(n14431), .A2(n14206), .ZN(n14143) );
  NAND2_X1 U15637 ( .A1(n14144), .A2(n14143), .ZN(n14146) );
  AOI22_X1 U15638 ( .A1(n14708), .A2(n14206), .B1(n7452), .B2(n14431), .ZN(
        n14145) );
  NOR2_X1 U15639 ( .A1(n14147), .A2(n14146), .ZN(n14148) );
  NAND2_X1 U15640 ( .A1(n14564), .A2(n14206), .ZN(n14151) );
  NAND2_X1 U15641 ( .A1(n14434), .A2(n14176), .ZN(n14150) );
  NAND2_X1 U15642 ( .A1(n14151), .A2(n14150), .ZN(n14153) );
  AOI22_X1 U15643 ( .A1(n14564), .A2(n14176), .B1(n14206), .B2(n14434), .ZN(
        n14152) );
  NAND2_X1 U15644 ( .A1(n14693), .A2(n7452), .ZN(n14156) );
  NAND2_X1 U15645 ( .A1(n14437), .A2(n14206), .ZN(n14155) );
  NAND2_X1 U15646 ( .A1(n14156), .A2(n14155), .ZN(n14161) );
  NAND2_X1 U15647 ( .A1(n14693), .A2(n14206), .ZN(n14158) );
  NAND2_X1 U15648 ( .A1(n14437), .A2(n14238), .ZN(n14157) );
  NAND2_X1 U15649 ( .A1(n14158), .A2(n14157), .ZN(n14159) );
  NAND2_X1 U15650 ( .A1(n14688), .A2(n14206), .ZN(n14164) );
  NAND2_X1 U15651 ( .A1(n14506), .A2(n14176), .ZN(n14163) );
  AOI22_X1 U15652 ( .A1(n14688), .A2(n7452), .B1(n14206), .B2(n14506), .ZN(
        n14165) );
  NAND2_X1 U15653 ( .A1(n14760), .A2(n7452), .ZN(n14167) );
  NAND2_X1 U15654 ( .A1(n14442), .A2(n14206), .ZN(n14166) );
  NAND2_X1 U15655 ( .A1(n14167), .A2(n14166), .ZN(n14171) );
  NAND2_X1 U15656 ( .A1(n14172), .A2(n14171), .ZN(n14170) );
  NAND2_X1 U15657 ( .A1(n14760), .A2(n14206), .ZN(n14168) );
  OAI21_X1 U15658 ( .B1(n14206), .B2(n7855), .A(n14168), .ZN(n14169) );
  NAND2_X1 U15659 ( .A1(n14170), .A2(n14169), .ZN(n14173) );
  NAND2_X1 U15660 ( .A1(n14677), .A2(n14206), .ZN(n14175) );
  NAND2_X1 U15661 ( .A1(n14507), .A2(n14217), .ZN(n14174) );
  NAND2_X1 U15662 ( .A1(n14175), .A2(n14174), .ZN(n14178) );
  AOI22_X1 U15663 ( .A1(n14677), .A2(n14207), .B1(n14206), .B2(n14507), .ZN(
        n14177) );
  NAND2_X1 U15664 ( .A1(n14792), .A2(n14201), .ZN(n14180) );
  OR2_X1 U15665 ( .A1(n14202), .A2(n14794), .ZN(n14179) );
  INV_X1 U15666 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n14184) );
  NAND2_X1 U15667 ( .A1(n13902), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n14183) );
  NAND2_X1 U15668 ( .A1(n14181), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n14182) );
  OAI211_X1 U15669 ( .C1(n14192), .C2(n14184), .A(n14183), .B(n14182), .ZN(
        n14375) );
  XNOR2_X1 U15670 ( .A(n14240), .B(n14375), .ZN(n14278) );
  OR2_X1 U15671 ( .A1(n14202), .A2(n14187), .ZN(n14188) );
  AND2_X1 U15672 ( .A1(n14290), .A2(n10125), .ZN(n14190) );
  NAND2_X1 U15673 ( .A1(n14296), .A2(n14295), .ZN(n14281) );
  AND2_X1 U15674 ( .A1(n14190), .A2(n14281), .ZN(n14196) );
  NAND2_X1 U15675 ( .A1(n14375), .A2(n14238), .ZN(n14239) );
  INV_X1 U15676 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n14661) );
  OR2_X1 U15677 ( .A1(n14191), .A2(n14661), .ZN(n14195) );
  INV_X1 U15678 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n14379) );
  OR2_X1 U15679 ( .A1(n14192), .A2(n14379), .ZN(n14194) );
  INV_X1 U15680 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14750) );
  OR2_X1 U15681 ( .A1(n10986), .A2(n14750), .ZN(n14193) );
  AND3_X1 U15682 ( .A1(n14195), .A2(n14194), .A3(n14193), .ZN(n14198) );
  AOI21_X1 U15683 ( .B1(n14196), .B2(n14239), .A(n14198), .ZN(n14197) );
  AOI21_X1 U15684 ( .B1(n14382), .B2(n14206), .A(n14197), .ZN(n14234) );
  NAND2_X1 U15685 ( .A1(n14382), .A2(n14238), .ZN(n14200) );
  INV_X1 U15686 ( .A(n14198), .ZN(n14414) );
  NAND2_X1 U15687 ( .A1(n14414), .A2(n14206), .ZN(n14199) );
  NAND2_X1 U15688 ( .A1(n14200), .A2(n14199), .ZN(n14233) );
  NAND2_X1 U15689 ( .A1(n14798), .A2(n14201), .ZN(n14204) );
  INV_X1 U15690 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14799) );
  OR2_X1 U15691 ( .A1(n14202), .A2(n14799), .ZN(n14203) );
  AND2_X1 U15692 ( .A1(n14304), .A2(n14238), .ZN(n14205) );
  AOI21_X1 U15693 ( .B1(n14664), .B2(n14206), .A(n14205), .ZN(n14231) );
  NAND2_X1 U15694 ( .A1(n14664), .A2(n14217), .ZN(n14209) );
  NAND2_X1 U15695 ( .A1(n14304), .A2(n14206), .ZN(n14208) );
  NAND2_X1 U15696 ( .A1(n14209), .A2(n14208), .ZN(n14230) );
  OAI22_X1 U15697 ( .A1(n14234), .A2(n14233), .B1(n14231), .B2(n14230), .ZN(
        n14210) );
  NAND2_X1 U15698 ( .A1(n14278), .A2(n14210), .ZN(n14236) );
  AND2_X1 U15699 ( .A1(n14412), .A2(n14206), .ZN(n14211) );
  AOI21_X1 U15700 ( .B1(n14465), .B2(n14207), .A(n14211), .ZN(n14227) );
  NAND2_X1 U15701 ( .A1(n14465), .A2(n14206), .ZN(n14214) );
  NAND2_X1 U15702 ( .A1(n14412), .A2(n14238), .ZN(n14213) );
  NAND2_X1 U15703 ( .A1(n14214), .A2(n14213), .ZN(n14226) );
  NAND2_X1 U15704 ( .A1(n14227), .A2(n14226), .ZN(n14215) );
  AND2_X1 U15705 ( .A1(n14236), .A2(n14215), .ZN(n14225) );
  AND2_X1 U15706 ( .A1(n14447), .A2(n14206), .ZN(n14216) );
  AOI21_X1 U15707 ( .B1(n14672), .B2(n14207), .A(n14216), .ZN(n14221) );
  NAND2_X1 U15708 ( .A1(n14672), .A2(n14206), .ZN(n14219) );
  NAND2_X1 U15709 ( .A1(n14447), .A2(n14238), .ZN(n14218) );
  NAND2_X1 U15710 ( .A1(n14219), .A2(n14218), .ZN(n14222) );
  NAND2_X1 U15711 ( .A1(n14221), .A2(n14222), .ZN(n14220) );
  INV_X1 U15712 ( .A(n14221), .ZN(n14224) );
  INV_X1 U15713 ( .A(n14222), .ZN(n14223) );
  INV_X1 U15714 ( .A(n14226), .ZN(n14229) );
  INV_X1 U15715 ( .A(n14227), .ZN(n14228) );
  AOI22_X1 U15716 ( .A1(n14231), .A2(n14230), .B1(n14229), .B2(n14228), .ZN(
        n14232) );
  NAND2_X1 U15717 ( .A1(n14278), .A2(n14232), .ZN(n14235) );
  AOI22_X1 U15718 ( .A1(n14236), .A2(n14235), .B1(n14234), .B2(n14233), .ZN(
        n14237) );
  NAND2_X1 U15719 ( .A1(n14206), .A2(n14375), .ZN(n14242) );
  NAND2_X1 U15720 ( .A1(n14239), .A2(n14238), .ZN(n14241) );
  MUX2_X1 U15721 ( .A(n14242), .B(n14241), .S(n14240), .Z(n14243) );
  XNOR2_X1 U15722 ( .A(n14382), .B(n14414), .ZN(n14276) );
  NAND2_X1 U15723 ( .A1(n14465), .A2(n14412), .ZN(n14448) );
  OR2_X1 U15724 ( .A1(n14465), .A2(n14412), .ZN(n14244) );
  NAND2_X1 U15725 ( .A1(n14448), .A2(n14244), .ZN(n14452) );
  XNOR2_X1 U15726 ( .A(n14688), .B(n14404), .ZN(n14526) );
  XNOR2_X1 U15727 ( .A(n14693), .B(n14402), .ZN(n14540) );
  INV_X1 U15728 ( .A(n14434), .ZN(n14399) );
  XNOR2_X1 U15729 ( .A(n14564), .B(n14399), .ZN(n14562) );
  INV_X1 U15730 ( .A(n14431), .ZN(n14245) );
  OR2_X1 U15731 ( .A1(n14708), .A2(n14245), .ZN(n14395) );
  NAND2_X1 U15732 ( .A1(n14708), .A2(n14245), .ZN(n14396) );
  NAND4_X1 U15733 ( .A1(n14249), .A2(n14248), .A3(n14247), .A4(n14246), .ZN(
        n14251) );
  NOR2_X1 U15734 ( .A1(n14251), .A2(n14250), .ZN(n14254) );
  NAND4_X1 U15735 ( .A1(n14255), .A2(n14254), .A3(n14253), .A4(n14252), .ZN(
        n14256) );
  OR4_X1 U15736 ( .A1(n14259), .A2(n14258), .A3(n14257), .A4(n14256), .ZN(
        n14260) );
  NOR2_X1 U15737 ( .A1(n14261), .A2(n14260), .ZN(n14263) );
  NAND4_X1 U15738 ( .A1(n14265), .A2(n14264), .A3(n14263), .A4(n14262), .ZN(
        n14266) );
  NOR2_X1 U15739 ( .A1(n14267), .A2(n14266), .ZN(n14269) );
  NAND4_X1 U15740 ( .A1(n14638), .A2(n14270), .A3(n14269), .A4(n14268), .ZN(
        n14271) );
  NOR2_X1 U15741 ( .A1(n14272), .A2(n14271), .ZN(n14273) );
  XNOR2_X1 U15742 ( .A(n14621), .B(n14428), .ZN(n14610) );
  XNOR2_X1 U15743 ( .A(n14593), .B(n14615), .ZN(n14589) );
  NAND4_X1 U15744 ( .A1(n14574), .A2(n14273), .A3(n14610), .A4(n14589), .ZN(
        n14274) );
  OR2_X1 U15745 ( .A1(n14677), .A2(n14507), .ZN(n14446) );
  NAND2_X1 U15746 ( .A1(n14677), .A2(n14507), .ZN(n14444) );
  NAND2_X1 U15747 ( .A1(n14446), .A2(n14444), .ZN(n14498) );
  AND4_X1 U15748 ( .A1(n14452), .A2(n7500), .A3(n14510), .A4(n14498), .ZN(
        n14275) );
  XNOR2_X1 U15749 ( .A(n14664), .B(n14304), .ZN(n14449) );
  XNOR2_X1 U15750 ( .A(n14672), .B(n14447), .ZN(n14473) );
  AND4_X1 U15751 ( .A1(n14276), .A2(n14275), .A3(n14449), .A4(n14473), .ZN(
        n14277) );
  AOI21_X1 U15752 ( .B1(n14279), .B2(n10130), .A(n10125), .ZN(n14300) );
  INV_X1 U15753 ( .A(n14279), .ZN(n14280) );
  NAND2_X1 U15754 ( .A1(n14280), .A2(n14366), .ZN(n14297) );
  INV_X1 U15755 ( .A(n14281), .ZN(n14284) );
  NOR3_X1 U15756 ( .A1(n14282), .A2(n14287), .A3(n14366), .ZN(n14283) );
  AOI211_X1 U15757 ( .C1(n14300), .C2(n14297), .A(n14284), .B(n14283), .ZN(
        n14285) );
  INV_X1 U15758 ( .A(n14294), .ZN(n14299) );
  INV_X1 U15759 ( .A(n13982), .ZN(n14286) );
  OAI211_X1 U15760 ( .C1(n10130), .C2(n14287), .A(n14286), .B(n14290), .ZN(
        n14288) );
  INV_X1 U15761 ( .A(n14290), .ZN(n14291) );
  NAND4_X1 U15762 ( .A1(n16076), .A2(n14292), .A3(n14291), .A4(n14613), .ZN(
        n14293) );
  OAI211_X1 U15763 ( .C1(n14295), .C2(n14294), .A(n14293), .B(P2_B_REG_SCAN_IN), .ZN(n14302) );
  INV_X1 U15764 ( .A(n14296), .ZN(n14298) );
  NAND4_X1 U15765 ( .A1(n14300), .A2(n14299), .A3(n14298), .A4(n14297), .ZN(
        n14301) );
  MUX2_X1 U15766 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n14375), .S(n14322), .Z(
        P2_U3562) );
  MUX2_X1 U15767 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n14414), .S(n14322), .Z(
        P2_U3561) );
  MUX2_X1 U15768 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n14304), .S(n14322), .Z(
        P2_U3560) );
  MUX2_X1 U15769 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n14412), .S(n14322), .Z(
        P2_U3559) );
  MUX2_X1 U15770 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n14447), .S(n14322), .Z(
        P2_U3558) );
  MUX2_X1 U15771 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n14507), .S(n14322), .Z(
        P2_U3557) );
  MUX2_X1 U15772 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n14442), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15773 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n14506), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15774 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n14437), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U15775 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n14434), .S(P2_U3947), .Z(
        P2_U3553) );
  MUX2_X1 U15776 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n14431), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15777 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n14615), .S(P2_U3947), .Z(
        P2_U3551) );
  MUX2_X1 U15778 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n14428), .S(P2_U3947), .Z(
        P2_U3550) );
  MUX2_X1 U15779 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n14612), .S(n14322), .Z(
        P2_U3549) );
  MUX2_X1 U15780 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n14305), .S(n14322), .Z(
        P2_U3548) );
  MUX2_X1 U15781 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n14306), .S(n14322), .Z(
        P2_U3547) );
  MUX2_X1 U15782 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n14307), .S(n14322), .Z(
        P2_U3546) );
  MUX2_X1 U15783 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n14308), .S(n14322), .Z(
        P2_U3545) );
  MUX2_X1 U15784 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n14309), .S(n14322), .Z(
        P2_U3544) );
  MUX2_X1 U15785 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n14310), .S(n14322), .Z(
        P2_U3543) );
  MUX2_X1 U15786 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n14311), .S(n14322), .Z(
        P2_U3542) );
  MUX2_X1 U15787 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n14312), .S(n14322), .Z(
        P2_U3541) );
  MUX2_X1 U15788 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n14313), .S(n14322), .Z(
        P2_U3540) );
  MUX2_X1 U15789 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n14314), .S(n14322), .Z(
        P2_U3539) );
  MUX2_X1 U15790 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n14315), .S(n14322), .Z(
        P2_U3538) );
  MUX2_X1 U15791 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n14316), .S(n14322), .Z(
        P2_U3537) );
  MUX2_X1 U15792 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n14317), .S(n14322), .Z(
        P2_U3536) );
  MUX2_X1 U15793 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n14318), .S(n14322), .Z(
        P2_U3535) );
  MUX2_X1 U15794 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n14319), .S(n14322), .Z(
        P2_U3534) );
  MUX2_X1 U15795 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n14320), .S(n14322), .Z(
        P2_U3533) );
  MUX2_X1 U15796 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n14321), .S(n14322), .Z(
        P2_U3532) );
  MUX2_X1 U15797 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n14323), .S(n14322), .Z(
        P2_U3531) );
  AOI211_X1 U15798 ( .C1(n14326), .C2(n14325), .A(n16228), .B(n14324), .ZN(
        n14327) );
  INV_X1 U15799 ( .A(n14327), .ZN(n14337) );
  INV_X1 U15800 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14329) );
  OAI21_X1 U15801 ( .B1(n16254), .B2(n14329), .A(n14328), .ZN(n14330) );
  AOI21_X1 U15802 ( .B1(n14331), .B2(n16234), .A(n14330), .ZN(n14336) );
  OAI211_X1 U15803 ( .C1(n14334), .C2(n14333), .A(n16222), .B(n14332), .ZN(
        n14335) );
  NAND3_X1 U15804 ( .A1(n14337), .A2(n14336), .A3(n14335), .ZN(P2_U3221) );
  XNOR2_X1 U15805 ( .A(n16218), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n16214) );
  NOR2_X1 U15806 ( .A1(n14345), .A2(n14338), .ZN(n14340) );
  NOR2_X1 U15807 ( .A1(n14340), .A2(n14339), .ZN(n16201) );
  NAND2_X1 U15808 ( .A1(n16207), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n14341) );
  OAI21_X1 U15809 ( .B1(n16207), .B2(P2_REG2_REG_16__SCAN_IN), .A(n14341), 
        .ZN(n16200) );
  NOR2_X1 U15810 ( .A1(n16201), .A2(n16200), .ZN(n16199) );
  AOI21_X1 U15811 ( .B1(n16207), .B2(P2_REG2_REG_16__SCAN_IN), .A(n16199), 
        .ZN(n16215) );
  NOR2_X1 U15812 ( .A1(n16214), .A2(n16215), .ZN(n16213) );
  AOI21_X1 U15813 ( .B1(n16218), .B2(P2_REG2_REG_17__SCAN_IN), .A(n16213), 
        .ZN(n14360) );
  XNOR2_X1 U15814 ( .A(n14360), .B(n14359), .ZN(n14358) );
  XNOR2_X1 U15815 ( .A(n14358), .B(n12457), .ZN(n14353) );
  INV_X1 U15816 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n14343) );
  NAND2_X1 U15817 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3088), .ZN(n14342)
         );
  OAI21_X1 U15818 ( .B1(n16254), .B2(n14343), .A(n14342), .ZN(n14344) );
  AOI21_X1 U15819 ( .B1(n14349), .B2(n16234), .A(n14344), .ZN(n14352) );
  XNOR2_X1 U15820 ( .A(n16218), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n16211) );
  NOR2_X1 U15821 ( .A1(n14346), .A2(n14345), .ZN(n14348) );
  XNOR2_X1 U15822 ( .A(n16207), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n16203) );
  NOR2_X1 U15823 ( .A1(n16211), .A2(n16212), .ZN(n16210) );
  XNOR2_X1 U15824 ( .A(n14355), .B(n14349), .ZN(n14350) );
  NAND2_X1 U15825 ( .A1(n14350), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n14354) );
  OAI211_X1 U15826 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n14350), .A(n16250), 
        .B(n14354), .ZN(n14351) );
  OAI211_X1 U15827 ( .C1(n16247), .C2(n14353), .A(n14352), .B(n14351), .ZN(
        P2_U3232) );
  OAI21_X1 U15828 ( .B1(n14355), .B2(n14359), .A(n14354), .ZN(n14357) );
  INV_X1 U15829 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n14721) );
  XNOR2_X1 U15830 ( .A(n10130), .B(n14721), .ZN(n14356) );
  XNOR2_X1 U15831 ( .A(n14357), .B(n14356), .ZN(n14370) );
  MUX2_X1 U15832 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n14624), .S(n10130), .Z(
        n14363) );
  INV_X1 U15833 ( .A(n14358), .ZN(n14361) );
  AOI22_X1 U15834 ( .A1(n14361), .A2(n12457), .B1(n14360), .B2(n14359), .ZN(
        n14362) );
  XOR2_X1 U15835 ( .A(n14363), .B(n14362), .Z(n14368) );
  NAND2_X1 U15836 ( .A1(n16097), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n14364) );
  OAI211_X1 U15837 ( .C1(n16189), .C2(n14366), .A(n14365), .B(n14364), .ZN(
        n14367) );
  AOI21_X1 U15838 ( .B1(n16222), .B2(n14368), .A(n14367), .ZN(n14369) );
  OAI21_X1 U15839 ( .B1(n14370), .B2(n16228), .A(n14369), .ZN(P2_U3233) );
  INV_X1 U15840 ( .A(n14677), .ZN(n14496) );
  OR2_X2 U15841 ( .A1(n14620), .A2(n14621), .ZN(n14618) );
  INV_X1 U15842 ( .A(n14708), .ZN(n14577) );
  NAND2_X1 U15843 ( .A1(n14496), .A2(n14516), .ZN(n14491) );
  XNOR2_X1 U15844 ( .A(n14240), .B(n14378), .ZN(n14371) );
  NAND2_X1 U15845 ( .A1(n14656), .A2(n14650), .ZN(n14377) );
  NOR2_X1 U15846 ( .A1(n14807), .A2(n14372), .ZN(n14373) );
  NOR2_X1 U15847 ( .A1(n14374), .A2(n14373), .ZN(n14413) );
  AND2_X1 U15848 ( .A1(n14375), .A2(n14413), .ZN(n14655) );
  INV_X1 U15849 ( .A(n14655), .ZN(n14659) );
  NOR2_X1 U15850 ( .A1(n14571), .A2(n14659), .ZN(n14380) );
  AOI21_X1 U15851 ( .B1(n14571), .B2(P2_REG2_REG_31__SCAN_IN), .A(n14380), 
        .ZN(n14376) );
  OAI211_X1 U15852 ( .C1(n14749), .C2(n14622), .A(n14377), .B(n14376), .ZN(
        P2_U3234) );
  OAI211_X1 U15853 ( .C1(n14753), .C2(n14419), .A(n14594), .B(n14378), .ZN(
        n14660) );
  NOR2_X1 U15854 ( .A1(n14644), .A2(n14379), .ZN(n14381) );
  AOI211_X1 U15855 ( .C1(n14382), .C2(n14646), .A(n14381), .B(n14380), .ZN(
        n14383) );
  OAI21_X1 U15856 ( .B1(n14660), .B2(n14553), .A(n14383), .ZN(P2_U3235) );
  NAND2_X1 U15857 ( .A1(n14426), .A2(n14386), .ZN(n14384) );
  NAND2_X1 U15858 ( .A1(n14385), .A2(n14384), .ZN(n14388) );
  OR2_X1 U15859 ( .A1(n14426), .A2(n14386), .ZN(n14387) );
  NOR2_X1 U15860 ( .A1(n14621), .A2(n14390), .ZN(n14389) );
  NAND2_X1 U15861 ( .A1(n14621), .A2(n14390), .ZN(n14391) );
  NAND2_X1 U15862 ( .A1(n14593), .A2(n14392), .ZN(n14393) );
  NAND2_X1 U15863 ( .A1(n14394), .A2(n14393), .ZN(n14573) );
  NAND2_X1 U15864 ( .A1(n14573), .A2(n14395), .ZN(n14397) );
  NAND2_X1 U15865 ( .A1(n14397), .A2(n14396), .ZN(n14558) );
  OR2_X1 U15866 ( .A1(n14564), .A2(n14399), .ZN(n14398) );
  NAND2_X1 U15867 ( .A1(n14564), .A2(n14399), .ZN(n14400) );
  AND2_X1 U15868 ( .A1(n14693), .A2(n14402), .ZN(n14401) );
  OR2_X1 U15869 ( .A1(n14402), .A2(n14693), .ZN(n14403) );
  NAND2_X1 U15870 ( .A1(n14688), .A2(n14404), .ZN(n14405) );
  OR2_X1 U15871 ( .A1(n14760), .A2(n7855), .ZN(n14406) );
  NAND2_X1 U15872 ( .A1(n14677), .A2(n14407), .ZN(n14408) );
  INV_X1 U15873 ( .A(n14447), .ZN(n14410) );
  AND2_X1 U15874 ( .A1(n14672), .A2(n14410), .ZN(n14411) );
  NAND2_X1 U15875 ( .A1(n14412), .A2(n14613), .ZN(n14416) );
  NAND2_X1 U15876 ( .A1(n14414), .A2(n14413), .ZN(n14415) );
  AOI211_X1 U15877 ( .C1(n14664), .C2(n14460), .A(n7458), .B(n14419), .ZN(
        n14663) );
  INV_X1 U15878 ( .A(n14664), .ZN(n14423) );
  INV_X1 U15879 ( .A(n14420), .ZN(n14421) );
  AOI22_X1 U15880 ( .A1(n14421), .A2(n14598), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14571), .ZN(n14422) );
  OAI21_X1 U15881 ( .B1(n14423), .B2(n14622), .A(n14422), .ZN(n14450) );
  OR2_X1 U15882 ( .A1(n14426), .A2(n14612), .ZN(n14427) );
  NAND2_X1 U15883 ( .A1(n14621), .A2(n14428), .ZN(n14429) );
  AND2_X1 U15884 ( .A1(n14593), .A2(n14615), .ZN(n14430) );
  NAND2_X1 U15885 ( .A1(n14708), .A2(n14431), .ZN(n14432) );
  NAND2_X1 U15886 ( .A1(n14433), .A2(n14432), .ZN(n14561) );
  NAND2_X1 U15887 ( .A1(n14561), .A2(n14562), .ZN(n14436) );
  NAND2_X1 U15888 ( .A1(n14564), .A2(n14434), .ZN(n14435) );
  NAND2_X1 U15889 ( .A1(n14693), .A2(n14437), .ZN(n14438) );
  INV_X1 U15890 ( .A(n14526), .ZN(n14440) );
  OR2_X1 U15891 ( .A1(n14688), .A2(n14506), .ZN(n14441) );
  NAND2_X1 U15892 ( .A1(n14760), .A2(n14442), .ZN(n14443) );
  INV_X1 U15893 ( .A(n14444), .ZN(n14445) );
  INV_X1 U15894 ( .A(n14452), .ZN(n14458) );
  OAI21_X1 U15895 ( .B1(n14666), .B2(n14571), .A(n14451), .ZN(P2_U3236) );
  OAI21_X1 U15896 ( .B1(n14453), .B2(n14452), .A(n7449), .ZN(n14454) );
  OAI21_X1 U15897 ( .B1(n14459), .B2(n14458), .A(n14457), .ZN(n14670) );
  INV_X1 U15898 ( .A(n14670), .ZN(n14468) );
  AOI21_X1 U15899 ( .B1(n14465), .B2(n14481), .A(n7458), .ZN(n14461) );
  NAND2_X1 U15900 ( .A1(n14461), .A2(n14460), .ZN(n14668) );
  OAI22_X1 U15901 ( .A1(n14463), .A2(n14641), .B1(n14462), .B2(n14644), .ZN(
        n14464) );
  AOI21_X1 U15902 ( .B1(n14465), .B2(n14646), .A(n14464), .ZN(n14466) );
  OAI21_X1 U15903 ( .B1(n14668), .B2(n14553), .A(n14466), .ZN(n14467) );
  AOI21_X1 U15904 ( .B1(n14468), .B2(n14640), .A(n14467), .ZN(n14469) );
  OAI21_X1 U15905 ( .B1(n14669), .B2(n14571), .A(n14469), .ZN(P2_U3237) );
  XNOR2_X1 U15906 ( .A(n14470), .B(n14473), .ZN(n14472) );
  AOI21_X1 U15907 ( .B1(n14472), .B2(n7449), .A(n14471), .ZN(n14674) );
  NAND2_X1 U15908 ( .A1(n14474), .A2(n14473), .ZN(n14475) );
  NAND2_X1 U15909 ( .A1(n14476), .A2(n14475), .ZN(n14675) );
  NAND2_X1 U15910 ( .A1(n14477), .A2(n14598), .ZN(n14478) );
  OAI21_X1 U15911 ( .B1(n14644), .B2(n14479), .A(n14478), .ZN(n14480) );
  AOI21_X1 U15912 ( .B1(n14672), .B2(n14646), .A(n14480), .ZN(n14484) );
  AOI21_X1 U15913 ( .B1(n14491), .B2(n14672), .A(n7458), .ZN(n14482) );
  AND2_X1 U15914 ( .A1(n14482), .A2(n14481), .ZN(n14671) );
  NAND2_X1 U15915 ( .A1(n14671), .A2(n14650), .ZN(n14483) );
  OAI211_X1 U15916 ( .C1(n14675), .C2(n14604), .A(n14484), .B(n14483), .ZN(
        n14485) );
  INV_X1 U15917 ( .A(n14485), .ZN(n14486) );
  OAI21_X1 U15918 ( .B1(n14571), .B2(n14674), .A(n14486), .ZN(P2_U3238) );
  XOR2_X1 U15919 ( .A(n14498), .B(n14487), .Z(n14490) );
  INV_X1 U15920 ( .A(n14488), .ZN(n14489) );
  AOI21_X1 U15921 ( .B1(n14490), .B2(n7449), .A(n14489), .ZN(n14679) );
  INV_X1 U15922 ( .A(n14516), .ZN(n14493) );
  INV_X1 U15923 ( .A(n14491), .ZN(n14492) );
  AOI211_X1 U15924 ( .C1(n14677), .C2(n14493), .A(n7458), .B(n14492), .ZN(
        n14676) );
  AOI22_X1 U15925 ( .A1(n14494), .A2(n14598), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14571), .ZN(n14495) );
  OAI21_X1 U15926 ( .B1(n14496), .B2(n14622), .A(n14495), .ZN(n14500) );
  XOR2_X1 U15927 ( .A(n14498), .B(n14497), .Z(n14680) );
  NOR2_X1 U15928 ( .A1(n14680), .A2(n14604), .ZN(n14499) );
  AOI211_X1 U15929 ( .C1(n14676), .C2(n14650), .A(n14500), .B(n14499), .ZN(
        n14501) );
  OAI21_X1 U15930 ( .B1(n14571), .B2(n14679), .A(n14501), .ZN(P2_U3239) );
  NAND2_X1 U15931 ( .A1(n14503), .A2(n14502), .ZN(n14504) );
  NAND3_X1 U15932 ( .A1(n14505), .A2(n7449), .A3(n14504), .ZN(n14509) );
  AOI22_X1 U15933 ( .A1(n14507), .A2(n14614), .B1(n14613), .B2(n14506), .ZN(
        n14508) );
  AND2_X1 U15934 ( .A1(n14509), .A2(n14508), .ZN(n14682) );
  NAND2_X1 U15935 ( .A1(n14511), .A2(n14510), .ZN(n14512) );
  NAND2_X1 U15936 ( .A1(n14513), .A2(n14512), .ZN(n14683) );
  INV_X1 U15937 ( .A(n14683), .ZN(n14523) );
  NAND2_X1 U15938 ( .A1(n14760), .A2(n14532), .ZN(n14514) );
  NAND2_X1 U15939 ( .A1(n14514), .A2(n14594), .ZN(n14515) );
  OR2_X1 U15940 ( .A1(n14516), .A2(n14515), .ZN(n14681) );
  NAND2_X1 U15941 ( .A1(n14517), .A2(n14598), .ZN(n14518) );
  OAI21_X1 U15942 ( .B1(n14644), .B2(n14519), .A(n14518), .ZN(n14520) );
  AOI21_X1 U15943 ( .B1(n14760), .B2(n14646), .A(n14520), .ZN(n14521) );
  OAI21_X1 U15944 ( .B1(n14681), .B2(n14553), .A(n14521), .ZN(n14522) );
  AOI21_X1 U15945 ( .B1(n14523), .B2(n14640), .A(n14522), .ZN(n14524) );
  OAI21_X1 U15946 ( .B1(n14571), .B2(n14682), .A(n14524), .ZN(P2_U3240) );
  OAI21_X1 U15947 ( .B1(n7519), .B2(n14526), .A(n14525), .ZN(n14686) );
  NAND2_X1 U15948 ( .A1(n14527), .A2(n14526), .ZN(n14528) );
  AOI21_X1 U15949 ( .B1(n14529), .B2(n14528), .A(n14591), .ZN(n14530) );
  AOI211_X1 U15950 ( .C1(n14686), .C2(n10128), .A(n14531), .B(n14530), .ZN(
        n14690) );
  AOI211_X1 U15951 ( .C1(n14688), .C2(n14548), .A(n7458), .B(n7994), .ZN(
        n14687) );
  NOR2_X1 U15952 ( .A1(n14533), .A2(n14622), .ZN(n14537) );
  OAI22_X1 U15953 ( .A1(n14535), .A2(n14641), .B1(n14534), .B2(n14644), .ZN(
        n14536) );
  AOI211_X1 U15954 ( .C1(n14687), .C2(n14650), .A(n14537), .B(n14536), .ZN(
        n14539) );
  INV_X1 U15955 ( .A(n14629), .ZN(n14555) );
  NAND2_X1 U15956 ( .A1(n14686), .A2(n14555), .ZN(n14538) );
  OAI211_X1 U15957 ( .C1(n14690), .C2(n14571), .A(n14539), .B(n14538), .ZN(
        P2_U3241) );
  INV_X1 U15958 ( .A(n14540), .ZN(n14542) );
  XNOR2_X1 U15959 ( .A(n14541), .B(n14542), .ZN(n14694) );
  NAND2_X1 U15960 ( .A1(n14694), .A2(n10128), .ZN(n14547) );
  XNOR2_X1 U15961 ( .A(n14543), .B(n14542), .ZN(n14545) );
  AOI21_X1 U15962 ( .B1(n14545), .B2(n7449), .A(n14544), .ZN(n14546) );
  NAND2_X1 U15963 ( .A1(n14547), .A2(n14546), .ZN(n14698) );
  INV_X1 U15964 ( .A(n14698), .ZN(n14557) );
  AOI21_X1 U15965 ( .B1(n14693), .B2(n14563), .A(n7458), .ZN(n14549) );
  NAND2_X1 U15966 ( .A1(n14549), .A2(n14548), .ZN(n14695) );
  AOI22_X1 U15967 ( .A1(n14550), .A2(n14598), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n14571), .ZN(n14552) );
  NAND2_X1 U15968 ( .A1(n14693), .A2(n14646), .ZN(n14551) );
  OAI211_X1 U15969 ( .C1(n14695), .C2(n14553), .A(n14552), .B(n14551), .ZN(
        n14554) );
  AOI21_X1 U15970 ( .B1(n14694), .B2(n14555), .A(n14554), .ZN(n14556) );
  OAI21_X1 U15971 ( .B1(n14557), .B2(n14571), .A(n14556), .ZN(P2_U3242) );
  XNOR2_X1 U15972 ( .A(n14558), .B(n14562), .ZN(n14560) );
  OAI21_X1 U15973 ( .B1(n14560), .B2(n14591), .A(n14559), .ZN(n14701) );
  INV_X1 U15974 ( .A(n14701), .ZN(n14570) );
  XOR2_X1 U15975 ( .A(n14562), .B(n14561), .Z(n14703) );
  AOI211_X1 U15976 ( .C1(n14564), .C2(n14578), .A(n7458), .B(n7996), .ZN(
        n14702) );
  NAND2_X1 U15977 ( .A1(n14702), .A2(n14650), .ZN(n14567) );
  AOI22_X1 U15978 ( .A1(n14565), .A2(n14598), .B1(n14571), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n14566) );
  OAI211_X1 U15979 ( .C1(n14769), .C2(n14622), .A(n14567), .B(n14566), .ZN(
        n14568) );
  AOI21_X1 U15980 ( .B1(n14703), .B2(n14640), .A(n14568), .ZN(n14569) );
  OAI21_X1 U15981 ( .B1(n14571), .B2(n14570), .A(n14569), .ZN(P2_U3243) );
  XNOR2_X1 U15982 ( .A(n14572), .B(n14574), .ZN(n14711) );
  XOR2_X1 U15983 ( .A(n14573), .B(n14574), .Z(n14576) );
  OAI21_X1 U15984 ( .B1(n14576), .B2(n14591), .A(n14575), .ZN(n14706) );
  OR2_X1 U15985 ( .A1(n14597), .A2(n14577), .ZN(n14579) );
  AND3_X1 U15986 ( .A1(n14579), .A2(n14578), .A3(n14594), .ZN(n14707) );
  NAND2_X1 U15987 ( .A1(n14707), .A2(n14650), .ZN(n14584) );
  OAI22_X1 U15988 ( .A1(n14581), .A2(n14641), .B1(n14644), .B2(n14580), .ZN(
        n14582) );
  AOI21_X1 U15989 ( .B1(n14708), .B2(n14646), .A(n14582), .ZN(n14583) );
  NAND2_X1 U15990 ( .A1(n14584), .A2(n14583), .ZN(n14585) );
  AOI21_X1 U15991 ( .B1(n14706), .B2(n14644), .A(n14585), .ZN(n14586) );
  OAI21_X1 U15992 ( .B1(n14711), .B2(n14604), .A(n14586), .ZN(P2_U3244) );
  XNOR2_X1 U15993 ( .A(n14587), .B(n14589), .ZN(n14714) );
  INV_X1 U15994 ( .A(n14714), .ZN(n14605) );
  XOR2_X1 U15995 ( .A(n14588), .B(n14589), .Z(n14592) );
  OAI21_X1 U15996 ( .B1(n14592), .B2(n14591), .A(n14590), .ZN(n14712) );
  NAND2_X1 U15997 ( .A1(n14618), .A2(n14593), .ZN(n14595) );
  NAND2_X1 U15998 ( .A1(n14595), .A2(n14594), .ZN(n14596) );
  NOR2_X1 U15999 ( .A1(n14597), .A2(n14596), .ZN(n14713) );
  NAND2_X1 U16000 ( .A1(n14713), .A2(n14650), .ZN(n14601) );
  AOI22_X1 U16001 ( .A1(n14571), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14599), 
        .B2(n14598), .ZN(n14600) );
  OAI211_X1 U16002 ( .C1(n14774), .C2(n14622), .A(n14601), .B(n14600), .ZN(
        n14602) );
  AOI21_X1 U16003 ( .B1(n14712), .B2(n14644), .A(n14602), .ZN(n14603) );
  OAI21_X1 U16004 ( .B1(n14605), .B2(n14604), .A(n14603), .ZN(P2_U3245) );
  NAND2_X1 U16005 ( .A1(n14606), .A2(n14610), .ZN(n14607) );
  NAND2_X1 U16006 ( .A1(n14608), .A2(n14607), .ZN(n14717) );
  XOR2_X1 U16007 ( .A(n14609), .B(n14610), .Z(n14611) );
  NAND2_X1 U16008 ( .A1(n14611), .A2(n7449), .ZN(n14617) );
  AOI22_X1 U16009 ( .A1(n14615), .A2(n14614), .B1(n14613), .B2(n14612), .ZN(
        n14616) );
  OAI211_X1 U16010 ( .C1(n14717), .C2(n8139), .A(n14617), .B(n14616), .ZN(
        n14718) );
  NAND2_X1 U16011 ( .A1(n14718), .A2(n14644), .ZN(n14628) );
  INV_X1 U16012 ( .A(n14618), .ZN(n14619) );
  AOI211_X1 U16013 ( .C1(n14621), .C2(n14620), .A(n7458), .B(n14619), .ZN(
        n14719) );
  INV_X1 U16014 ( .A(n14621), .ZN(n14778) );
  NOR2_X1 U16015 ( .A1(n14778), .A2(n14622), .ZN(n14626) );
  OAI22_X1 U16016 ( .A1(n14644), .A2(n14624), .B1(n14623), .B2(n14641), .ZN(
        n14625) );
  AOI211_X1 U16017 ( .C1(n14719), .C2(n14650), .A(n14626), .B(n14625), .ZN(
        n14627) );
  OAI211_X1 U16018 ( .C1(n14717), .C2(n14629), .A(n14628), .B(n14627), .ZN(
        P2_U3246) );
  NAND3_X1 U16019 ( .A1(n14632), .A2(n14631), .A3(n14630), .ZN(n14633) );
  NAND3_X1 U16020 ( .A1(n14635), .A2(n7449), .A3(n14633), .ZN(n14637) );
  NAND2_X1 U16021 ( .A1(n14637), .A2(n14636), .ZN(n14729) );
  NAND2_X1 U16022 ( .A1(n14729), .A2(n14644), .ZN(n14654) );
  XNOR2_X1 U16023 ( .A(n14639), .B(n14638), .ZN(n14731) );
  NAND2_X1 U16024 ( .A1(n14731), .A2(n14640), .ZN(n14653) );
  OAI22_X1 U16025 ( .A1(n14644), .A2(n14643), .B1(n14642), .B2(n14641), .ZN(
        n14645) );
  AOI21_X1 U16026 ( .B1(n14728), .B2(n14646), .A(n14645), .ZN(n14652) );
  AOI21_X1 U16027 ( .B1(n14647), .B2(n14728), .A(n7458), .ZN(n14649) );
  AND2_X1 U16028 ( .A1(n14649), .A2(n14648), .ZN(n14730) );
  NAND2_X1 U16029 ( .A1(n14730), .A2(n14650), .ZN(n14651) );
  NAND4_X1 U16030 ( .A1(n14654), .A2(n14653), .A3(n14652), .A4(n14651), .ZN(
        P2_U3248) );
  INV_X1 U16031 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n14657) );
  NOR2_X1 U16032 ( .A1(n14656), .A2(n14655), .ZN(n14746) );
  OAI21_X1 U16033 ( .B1(n14749), .B2(n14734), .A(n14658), .ZN(P2_U3530) );
  AND2_X1 U16034 ( .A1(n14660), .A2(n14659), .ZN(n14751) );
  MUX2_X1 U16035 ( .A(n14751), .B(n14661), .S(n16584), .Z(n14662) );
  OAI21_X1 U16036 ( .B1(n14753), .B2(n14734), .A(n14662), .ZN(P2_U3529) );
  AOI21_X1 U16037 ( .B1(n14709), .B2(n14664), .A(n14663), .ZN(n14665) );
  MUX2_X1 U16038 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n14754), .S(n14740), .Z(
        P2_U3528) );
  AOI21_X1 U16039 ( .B1(n14709), .B2(n14672), .A(n14671), .ZN(n14673) );
  OAI211_X1 U16040 ( .C1(n14675), .C2(n14735), .A(n14674), .B(n14673), .ZN(
        n14756) );
  MUX2_X1 U16041 ( .A(n14756), .B(P2_REG1_REG_27__SCAN_IN), .S(n16584), .Z(
        P2_U3526) );
  AOI21_X1 U16042 ( .B1(n14709), .B2(n14677), .A(n14676), .ZN(n14678) );
  OAI211_X1 U16043 ( .C1(n14680), .C2(n14735), .A(n14679), .B(n14678), .ZN(
        n14757) );
  MUX2_X1 U16044 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14757), .S(n14740), .Z(
        P2_U3525) );
  OAI211_X1 U16045 ( .C1(n14683), .C2(n14735), .A(n14682), .B(n14681), .ZN(
        n14758) );
  MUX2_X1 U16046 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14758), .S(n14740), .Z(
        n14684) );
  AOI21_X1 U16047 ( .B1(n14742), .B2(n14760), .A(n14684), .ZN(n14685) );
  INV_X1 U16048 ( .A(n14685), .ZN(P2_U3524) );
  INV_X1 U16049 ( .A(n14686), .ZN(n14692) );
  AOI21_X1 U16050 ( .B1(n14709), .B2(n14688), .A(n14687), .ZN(n14689) );
  OAI211_X1 U16051 ( .C1(n14692), .C2(n14691), .A(n14690), .B(n14689), .ZN(
        n14762) );
  MUX2_X1 U16052 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14762), .S(n14740), .Z(
        P2_U3523) );
  INV_X1 U16053 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n14699) );
  NAND2_X1 U16054 ( .A1(n14694), .A2(n16532), .ZN(n14696) );
  NAND2_X1 U16055 ( .A1(n14696), .A2(n14695), .ZN(n14697) );
  NOR2_X1 U16056 ( .A1(n14698), .A2(n14697), .ZN(n14763) );
  MUX2_X1 U16057 ( .A(n14699), .B(n14763), .S(n14740), .Z(n14700) );
  OAI21_X1 U16058 ( .B1(n7995), .B2(n14734), .A(n14700), .ZN(P2_U3522) );
  INV_X1 U16059 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n14704) );
  AOI211_X1 U16060 ( .C1(n16583), .C2(n14703), .A(n14702), .B(n14701), .ZN(
        n14766) );
  MUX2_X1 U16061 ( .A(n14704), .B(n14766), .S(n14740), .Z(n14705) );
  OAI21_X1 U16062 ( .B1(n14769), .B2(n14734), .A(n14705), .ZN(P2_U3521) );
  AOI211_X1 U16063 ( .C1(n14709), .C2(n14708), .A(n14707), .B(n14706), .ZN(
        n14710) );
  OAI21_X1 U16064 ( .B1(n14735), .B2(n14711), .A(n14710), .ZN(n14770) );
  MUX2_X1 U16065 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14770), .S(n14740), .Z(
        P2_U3520) );
  INV_X1 U16066 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n14715) );
  AOI211_X1 U16067 ( .C1(n16583), .C2(n14714), .A(n14713), .B(n14712), .ZN(
        n14771) );
  MUX2_X1 U16068 ( .A(n14715), .B(n14771), .S(n14740), .Z(n14716) );
  OAI21_X1 U16069 ( .B1(n14774), .B2(n14734), .A(n14716), .ZN(P2_U3519) );
  INV_X1 U16070 ( .A(n14717), .ZN(n14720) );
  AOI211_X1 U16071 ( .C1(n14720), .C2(n16532), .A(n14719), .B(n14718), .ZN(
        n14775) );
  MUX2_X1 U16072 ( .A(n14721), .B(n14775), .S(n14740), .Z(n14722) );
  OAI21_X1 U16073 ( .B1(n14778), .B2(n14734), .A(n14722), .ZN(P2_U3518) );
  INV_X1 U16074 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14726) );
  AOI211_X1 U16075 ( .C1(n16583), .C2(n14725), .A(n14724), .B(n14723), .ZN(
        n14779) );
  MUX2_X1 U16076 ( .A(n14726), .B(n14779), .S(n14740), .Z(n14727) );
  OAI21_X1 U16077 ( .B1(n7992), .B2(n14734), .A(n14727), .ZN(P2_U3517) );
  INV_X1 U16078 ( .A(n14728), .ZN(n14786) );
  INV_X1 U16079 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n14732) );
  AOI211_X1 U16080 ( .C1(n16583), .C2(n14731), .A(n14730), .B(n14729), .ZN(
        n14782) );
  MUX2_X1 U16081 ( .A(n14732), .B(n14782), .S(n14740), .Z(n14733) );
  OAI21_X1 U16082 ( .B1(n14786), .B2(n14734), .A(n14733), .ZN(P2_U3516) );
  NOR2_X1 U16083 ( .A1(n14736), .A2(n14735), .ZN(n14739) );
  MUX2_X1 U16084 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14787), .S(n14740), .Z(
        n14741) );
  AOI21_X1 U16085 ( .B1(n14742), .B2(n14789), .A(n14741), .ZN(n14743) );
  INV_X1 U16086 ( .A(n14743), .ZN(P2_U3515) );
  MUX2_X1 U16087 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n14744), .S(n14740), .Z(
        P2_U3505) );
  MUX2_X1 U16088 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n14745), .S(n14740), .Z(
        P2_U3503) );
  INV_X1 U16089 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n14747) );
  MUX2_X1 U16090 ( .A(n14747), .B(n14746), .S(n16534), .Z(n14748) );
  MUX2_X1 U16091 ( .A(n14751), .B(n14750), .S(n16585), .Z(n14752) );
  OAI21_X1 U16092 ( .B1(n14753), .B2(n14785), .A(n14752), .ZN(P2_U3497) );
  MUX2_X1 U16093 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n14754), .S(n16534), .Z(
        P2_U3496) );
  MUX2_X1 U16094 ( .A(n14756), .B(P2_REG0_REG_27__SCAN_IN), .S(n16585), .Z(
        P2_U3494) );
  MUX2_X1 U16095 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14757), .S(n16534), .Z(
        P2_U3493) );
  MUX2_X1 U16096 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14758), .S(n16534), .Z(
        n14759) );
  AOI21_X1 U16097 ( .B1(n14790), .B2(n14760), .A(n14759), .ZN(n14761) );
  INV_X1 U16098 ( .A(n14761), .ZN(P2_U3492) );
  MUX2_X1 U16099 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14762), .S(n16534), .Z(
        P2_U3491) );
  INV_X1 U16100 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n14764) );
  MUX2_X1 U16101 ( .A(n14764), .B(n14763), .S(n16534), .Z(n14765) );
  OAI21_X1 U16102 ( .B1(n7995), .B2(n14785), .A(n14765), .ZN(P2_U3490) );
  INV_X1 U16103 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n14767) );
  MUX2_X1 U16104 ( .A(n14767), .B(n14766), .S(n16534), .Z(n14768) );
  OAI21_X1 U16105 ( .B1(n14769), .B2(n14785), .A(n14768), .ZN(P2_U3489) );
  MUX2_X1 U16106 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14770), .S(n16534), .Z(
        P2_U3488) );
  INV_X1 U16107 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n14772) );
  MUX2_X1 U16108 ( .A(n14772), .B(n14771), .S(n16534), .Z(n14773) );
  OAI21_X1 U16109 ( .B1(n14774), .B2(n14785), .A(n14773), .ZN(P2_U3487) );
  INV_X1 U16110 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n14776) );
  MUX2_X1 U16111 ( .A(n14776), .B(n14775), .S(n16534), .Z(n14777) );
  OAI21_X1 U16112 ( .B1(n14778), .B2(n14785), .A(n14777), .ZN(P2_U3486) );
  INV_X1 U16113 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n14780) );
  MUX2_X1 U16114 ( .A(n14780), .B(n14779), .S(n16534), .Z(n14781) );
  OAI21_X1 U16115 ( .B1(n7992), .B2(n14785), .A(n14781), .ZN(P2_U3484) );
  INV_X1 U16116 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n14783) );
  MUX2_X1 U16117 ( .A(n14783), .B(n14782), .S(n16534), .Z(n14784) );
  OAI21_X1 U16118 ( .B1(n14786), .B2(n14785), .A(n14784), .ZN(P2_U3481) );
  MUX2_X1 U16119 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14787), .S(n16534), .Z(
        n14788) );
  AOI21_X1 U16120 ( .B1(n14790), .B2(n14789), .A(n14788), .ZN(n14791) );
  INV_X1 U16121 ( .A(n14791), .ZN(P2_U3478) );
  INV_X1 U16122 ( .A(n14792), .ZN(n15906) );
  NAND3_X1 U16123 ( .A1(n14793), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n14795) );
  OAI22_X1 U16124 ( .A1(n10016), .A2(n14795), .B1(n14794), .B2(n14818), .ZN(
        n14796) );
  INV_X1 U16125 ( .A(n14796), .ZN(n14797) );
  OAI21_X1 U16126 ( .B1(n15906), .B2(n14816), .A(n14797), .ZN(P2_U3296) );
  INV_X1 U16127 ( .A(n14798), .ZN(n15908) );
  OAI222_X1 U16128 ( .A1(P2_U3088), .A2(n14800), .B1(n14816), .B2(n15908), 
        .C1(n14799), .C2(n14818), .ZN(P2_U3298) );
  NAND2_X1 U16129 ( .A1(n14802), .A2(n14801), .ZN(n14804) );
  OAI211_X1 U16130 ( .C1(n14818), .C2(n14805), .A(n14804), .B(n14803), .ZN(
        P2_U3299) );
  INV_X1 U16131 ( .A(n14806), .ZN(n15911) );
  OAI222_X1 U16132 ( .A1(n14818), .A2(n14808), .B1(n14816), .B2(n15911), .C1(
        n14807), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U16133 ( .A(n14809), .ZN(n14812) );
  INV_X1 U16134 ( .A(n14810), .ZN(n15914) );
  OAI222_X1 U16135 ( .A1(n14812), .A2(P2_U3088), .B1(n14816), .B2(n15914), 
        .C1(n14811), .C2(n14818), .ZN(P2_U3301) );
  INV_X1 U16136 ( .A(n14813), .ZN(n15918) );
  INV_X1 U16137 ( .A(n14814), .ZN(n14815) );
  OAI222_X1 U16138 ( .A1(n14818), .A2(n14817), .B1(n14816), .B2(n15918), .C1(
        n14815), .C2(P2_U3088), .ZN(P2_U3302) );
  MUX2_X1 U16139 ( .A(n14819), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI21_X1 U16140 ( .B1(n14822), .B2(n14821), .A(n14820), .ZN(n14823) );
  NAND2_X1 U16141 ( .A1(n14823), .A2(n14947), .ZN(n14828) );
  OAI22_X1 U16142 ( .A1(n14951), .A2(n15112), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14824), .ZN(n14826) );
  NOR2_X1 U16143 ( .A1(n14952), .A2(n15116), .ZN(n14825) );
  AOI211_X1 U16144 ( .C1(n14955), .C2(n15147), .A(n14826), .B(n14825), .ZN(
        n14827) );
  OAI211_X1 U16145 ( .C1(n15376), .C2(n14958), .A(n14828), .B(n14827), .ZN(
        P1_U3214) );
  INV_X1 U16146 ( .A(n14829), .ZN(n14833) );
  AOI21_X1 U16147 ( .B1(n14916), .B2(n14831), .A(n14830), .ZN(n14832) );
  OAI21_X1 U16148 ( .B1(n14833), .B2(n14832), .A(n14915), .ZN(n14839) );
  AND2_X1 U16149 ( .A1(n15146), .A2(n15329), .ZN(n14834) );
  AOI21_X1 U16150 ( .B1(n14961), .B2(n15331), .A(n14834), .ZN(n15400) );
  INV_X1 U16151 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14835) );
  OAI22_X1 U16152 ( .A1(n15400), .A2(n14836), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14835), .ZN(n14837) );
  AOI21_X1 U16153 ( .B1(n15187), .B2(n14893), .A(n14837), .ZN(n14838) );
  OAI211_X1 U16154 ( .C1(n15402), .C2(n14958), .A(n14839), .B(n14838), .ZN(
        P1_U3216) );
  OAI211_X1 U16155 ( .C1(n14842), .C2(n14841), .A(n14840), .B(n14947), .ZN(
        n14849) );
  AOI22_X1 U16156 ( .A1(n14844), .A2(n14843), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14848) );
  AOI22_X1 U16157 ( .A1(n14845), .A2(n14972), .B1(n14955), .B2(n9332), .ZN(
        n14847) );
  INV_X1 U16158 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14991) );
  NAND2_X1 U16159 ( .A1(n14893), .A2(n14991), .ZN(n14846) );
  NAND4_X1 U16160 ( .A1(n14849), .A2(n14848), .A3(n14847), .A4(n14846), .ZN(
        P1_U3218) );
  OAI21_X1 U16161 ( .B1(n14851), .B2(n14850), .A(n14906), .ZN(n14852) );
  NAND2_X1 U16162 ( .A1(n14852), .A2(n14915), .ZN(n14856) );
  NAND2_X1 U16163 ( .A1(n14955), .A2(n15289), .ZN(n14853) );
  NAND2_X1 U16164 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n15070)
         );
  OAI211_X1 U16165 ( .C1(n15214), .C2(n14951), .A(n14853), .B(n15070), .ZN(
        n14854) );
  AOI21_X1 U16166 ( .B1(n14893), .B2(n15259), .A(n14854), .ZN(n14855) );
  OAI211_X1 U16167 ( .C1(n8482), .C2(n14958), .A(n14856), .B(n14855), .ZN(
        P1_U3219) );
  AOI21_X1 U16168 ( .B1(n14907), .B2(n14858), .A(n14857), .ZN(n14859) );
  OAI21_X1 U16169 ( .B1(n14860), .B2(n14859), .A(n14915), .ZN(n14866) );
  NOR2_X1 U16170 ( .A1(n14861), .A2(n15214), .ZN(n14864) );
  OAI22_X1 U16171 ( .A1(n7885), .A2(n14951), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14862), .ZN(n14863) );
  AOI211_X1 U16172 ( .C1(n15222), .C2(n14893), .A(n14864), .B(n14863), .ZN(
        n14865) );
  OAI211_X1 U16173 ( .C1(n8453), .C2(n14958), .A(n14866), .B(n14865), .ZN(
        P1_U3223) );
  OAI21_X1 U16174 ( .B1(n14869), .B2(n14868), .A(n14867), .ZN(n14870) );
  NAND2_X1 U16175 ( .A1(n14870), .A2(n14947), .ZN(n14875) );
  INV_X1 U16176 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14871) );
  OAI22_X1 U16177 ( .A1(n14951), .A2(n15111), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14871), .ZN(n14873) );
  NOR2_X1 U16178 ( .A1(n14952), .A2(n15150), .ZN(n14872) );
  AOI211_X1 U16179 ( .C1(n14955), .C2(n15146), .A(n14873), .B(n14872), .ZN(
        n14874) );
  OAI211_X1 U16180 ( .C1(n8011), .C2(n14958), .A(n14875), .B(n14874), .ZN(
        P1_U3225) );
  INV_X1 U16181 ( .A(n15446), .ZN(n15311) );
  OAI21_X1 U16182 ( .B1(n14877), .B2(n14876), .A(n14887), .ZN(n14878) );
  NAND2_X1 U16183 ( .A1(n14878), .A2(n14947), .ZN(n14884) );
  OAI21_X1 U16184 ( .B1(n14951), .B2(n14880), .A(n14879), .ZN(n14882) );
  NOR2_X1 U16185 ( .A1(n14952), .A2(n15313), .ZN(n14881) );
  AOI211_X1 U16186 ( .C1(n14955), .C2(n15303), .A(n14882), .B(n14881), .ZN(
        n14883) );
  OAI211_X1 U16187 ( .C1(n15311), .C2(n14958), .A(n14884), .B(n14883), .ZN(
        P1_U3226) );
  AND3_X1 U16188 ( .A1(n14887), .A2(n14886), .A3(n14885), .ZN(n14888) );
  OAI21_X1 U16189 ( .B1(n14927), .B2(n14888), .A(n14915), .ZN(n14895) );
  NAND2_X1 U16190 ( .A1(n14955), .A2(n15330), .ZN(n14890) );
  OAI211_X1 U16191 ( .C1(n14891), .C2(n14951), .A(n14890), .B(n14889), .ZN(
        n14892) );
  AOI21_X1 U16192 ( .B1(n14893), .B2(n15294), .A(n14892), .ZN(n14894) );
  OAI211_X1 U16193 ( .C1(n15298), .C2(n14958), .A(n14895), .B(n14894), .ZN(
        P1_U3228) );
  OAI21_X1 U16194 ( .B1(n14898), .B2(n14897), .A(n14896), .ZN(n14899) );
  NAND2_X1 U16195 ( .A1(n14899), .A2(n14947), .ZN(n14904) );
  INV_X1 U16196 ( .A(n15132), .ZN(n15162) );
  INV_X1 U16197 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n14900) );
  OAI22_X1 U16198 ( .A1(n14951), .A2(n15162), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14900), .ZN(n14902) );
  NOR2_X1 U16199 ( .A1(n14952), .A2(n15168), .ZN(n14901) );
  AOI211_X1 U16200 ( .C1(n14955), .C2(n15198), .A(n14902), .B(n14901), .ZN(
        n14903) );
  OAI211_X1 U16201 ( .C1(n15173), .C2(n14958), .A(n14904), .B(n14903), .ZN(
        P1_U3229) );
  INV_X1 U16202 ( .A(n15421), .ZN(n15244) );
  AND2_X1 U16203 ( .A1(n14906), .A2(n14905), .ZN(n14909) );
  OAI211_X1 U16204 ( .C1(n14909), .C2(n14908), .A(n14915), .B(n14907), .ZN(
        n14914) );
  OAI22_X1 U16205 ( .A1(n14951), .A2(n15233), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14910), .ZN(n14912) );
  NOR2_X1 U16206 ( .A1(n14952), .A2(n15241), .ZN(n14911) );
  AOI211_X1 U16207 ( .C1(n14955), .C2(n15270), .A(n14912), .B(n14911), .ZN(
        n14913) );
  OAI211_X1 U16208 ( .C1(n15244), .C2(n14958), .A(n14914), .B(n14913), .ZN(
        P1_U3233) );
  OAI211_X1 U16209 ( .C1(n14918), .C2(n14917), .A(n14916), .B(n14915), .ZN(
        n14923) );
  OAI22_X1 U16210 ( .A1(n15163), .A2(n14951), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14919), .ZN(n14921) );
  NOR2_X1 U16211 ( .A1(n14952), .A2(n15202), .ZN(n14920) );
  AOI211_X1 U16212 ( .C1(n14955), .C2(n15199), .A(n14921), .B(n14920), .ZN(
        n14922) );
  OAI211_X1 U16213 ( .C1(n14958), .C2(n15206), .A(n14923), .B(n14922), .ZN(
        P1_U3235) );
  INV_X1 U16214 ( .A(n14924), .ZN(n14929) );
  NOR3_X1 U16215 ( .A1(n14927), .A2(n14926), .A3(n14925), .ZN(n14928) );
  OAI21_X1 U16216 ( .B1(n14929), .B2(n14928), .A(n14947), .ZN(n14933) );
  NAND2_X1 U16217 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n16269)
         );
  OAI21_X1 U16218 ( .B1(n14951), .B2(n15231), .A(n16269), .ZN(n14931) );
  NOR2_X1 U16219 ( .A1(n14952), .A2(n15271), .ZN(n14930) );
  AOI211_X1 U16220 ( .C1(n14955), .C2(n15304), .A(n14931), .B(n14930), .ZN(
        n14932) );
  OAI211_X1 U16221 ( .C1(n15274), .C2(n14958), .A(n14933), .B(n14932), .ZN(
        P1_U3238) );
  OAI21_X1 U16222 ( .B1(n14936), .B2(n14935), .A(n14934), .ZN(n14937) );
  NAND2_X1 U16223 ( .A1(n14937), .A2(n14947), .ZN(n14943) );
  OAI22_X1 U16224 ( .A1(n14951), .A2(n14939), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14938), .ZN(n14941) );
  NOR2_X1 U16225 ( .A1(n14952), .A2(n15126), .ZN(n14940) );
  AOI211_X1 U16226 ( .C1(n14955), .C2(n15132), .A(n14941), .B(n14940), .ZN(
        n14942) );
  OAI211_X1 U16227 ( .C1(n15125), .C2(n14958), .A(n14943), .B(n14942), .ZN(
        P1_U3240) );
  INV_X1 U16228 ( .A(n15451), .ZN(n15325) );
  OAI21_X1 U16229 ( .B1(n14946), .B2(n14945), .A(n14944), .ZN(n14948) );
  NAND2_X1 U16230 ( .A1(n14948), .A2(n14947), .ZN(n14957) );
  OAI21_X1 U16231 ( .B1(n14951), .B2(n14950), .A(n14949), .ZN(n14954) );
  NOR2_X1 U16232 ( .A1(n14952), .A2(n15322), .ZN(n14953) );
  AOI211_X1 U16233 ( .C1(n14955), .C2(n15332), .A(n14954), .B(n14953), .ZN(
        n14956) );
  OAI211_X1 U16234 ( .C1(n15325), .C2(n14958), .A(n14957), .B(n14956), .ZN(
        P1_U3241) );
  MUX2_X1 U16235 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14959), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16236 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n15095), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16237 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14960), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16238 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n15085), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16239 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n15133), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16240 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n15147), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16241 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n15132), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16242 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n15146), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16243 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n15198), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16244 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14961), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16245 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n15199), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16246 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n15258), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16247 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n15270), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16248 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n15289), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16249 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n15304), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16250 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n15330), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16251 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n15303), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16252 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n15332), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16253 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14962), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16254 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14963), .S(n14964), .Z(
        P1_U3572) );
  MUX2_X1 U16255 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14965), .S(n14964), .Z(
        P1_U3571) );
  MUX2_X1 U16256 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14966), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16257 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14967), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16258 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14968), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16259 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14969), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16260 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14970), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16261 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14971), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16262 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14972), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16263 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14973), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16264 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9332), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16265 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n10517), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16266 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14974), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U16267 ( .C1(n10316), .C2(n14977), .A(n16347), .B(n14976), .ZN(
        n14986) );
  AOI22_X1 U16268 ( .A1(n14978), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14985) );
  OAI211_X1 U16269 ( .C1(n14981), .C2(n14980), .A(n16354), .B(n14979), .ZN(
        n14984) );
  NAND2_X1 U16270 ( .A1(n15065), .A2(n14982), .ZN(n14983) );
  NAND4_X1 U16271 ( .A1(n14986), .A2(n14985), .A3(n14984), .A4(n14983), .ZN(
        P1_U3244) );
  MUX2_X1 U16272 ( .A(n11119), .B(P1_REG2_REG_3__SCAN_IN), .S(n14993), .Z(
        n14988) );
  NAND3_X1 U16273 ( .A1(n14989), .A2(n14988), .A3(n14987), .ZN(n14990) );
  NAND3_X1 U16274 ( .A1(n16347), .A2(n16344), .A3(n14990), .ZN(n15000) );
  OAI22_X1 U16275 ( .A1(n16364), .A2(n15992), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14991), .ZN(n14992) );
  AOI21_X1 U16276 ( .B1(n14993), .B2(n15065), .A(n14992), .ZN(n14999) );
  MUX2_X1 U16277 ( .A(n10307), .B(P1_REG1_REG_3__SCAN_IN), .S(n14993), .Z(
        n14995) );
  NAND3_X1 U16278 ( .A1(n14996), .A2(n14995), .A3(n14994), .ZN(n14997) );
  NAND3_X1 U16279 ( .A1(n16354), .A2(n16351), .A3(n14997), .ZN(n14998) );
  NAND3_X1 U16280 ( .A1(n15000), .A2(n14999), .A3(n14998), .ZN(P1_U3246) );
  NOR2_X1 U16281 ( .A1(n15002), .A2(n15001), .ZN(n15003) );
  OAI21_X1 U16282 ( .B1(n15003), .B2(n15018), .A(n16354), .ZN(n15014) );
  INV_X1 U16283 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n15005) );
  OAI21_X1 U16284 ( .B1(n16364), .B2(n15005), .A(n15004), .ZN(n15006) );
  AOI21_X1 U16285 ( .B1(n15007), .B2(n15065), .A(n15006), .ZN(n15013) );
  MUX2_X1 U16286 ( .A(n10385), .B(P1_REG2_REG_8__SCAN_IN), .S(n15007), .Z(
        n15008) );
  NAND3_X1 U16287 ( .A1(n15010), .A2(n15009), .A3(n15008), .ZN(n15011) );
  NAND3_X1 U16288 ( .A1(n16347), .A2(n15027), .A3(n15011), .ZN(n15012) );
  NAND3_X1 U16289 ( .A1(n15014), .A2(n15013), .A3(n15012), .ZN(P1_U3251) );
  INV_X1 U16290 ( .A(n15015), .ZN(n15020) );
  NOR3_X1 U16291 ( .A1(n15018), .A2(n15017), .A3(n15016), .ZN(n15019) );
  OAI21_X1 U16292 ( .B1(n15020), .B2(n15019), .A(n16354), .ZN(n15032) );
  INV_X1 U16293 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n15022) );
  OAI21_X1 U16294 ( .B1(n16364), .B2(n15022), .A(n15021), .ZN(n15023) );
  AOI21_X1 U16295 ( .B1(n15024), .B2(n15065), .A(n15023), .ZN(n15031) );
  MUX2_X1 U16296 ( .A(n10388), .B(P1_REG2_REG_9__SCAN_IN), .S(n15024), .Z(
        n15025) );
  NAND3_X1 U16297 ( .A1(n15027), .A2(n15026), .A3(n15025), .ZN(n15028) );
  NAND3_X1 U16298 ( .A1(n16347), .A2(n15029), .A3(n15028), .ZN(n15030) );
  NAND3_X1 U16299 ( .A1(n15032), .A2(n15031), .A3(n15030), .ZN(P1_U3252) );
  NOR2_X1 U16300 ( .A1(n15034), .A2(n15033), .ZN(n15036) );
  OAI21_X1 U16301 ( .B1(n15036), .B2(n15035), .A(n16354), .ZN(n15047) );
  INV_X1 U16302 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n15923) );
  OAI21_X1 U16303 ( .B1(n16364), .B2(n15923), .A(n15037), .ZN(n15038) );
  AOI21_X1 U16304 ( .B1(n15039), .B2(n15065), .A(n15038), .ZN(n15046) );
  MUX2_X1 U16305 ( .A(n11867), .B(P1_REG2_REG_11__SCAN_IN), .S(n15039), .Z(
        n15040) );
  NAND3_X1 U16306 ( .A1(n15042), .A2(n15041), .A3(n15040), .ZN(n15043) );
  NAND3_X1 U16307 ( .A1(n16347), .A2(n15044), .A3(n15043), .ZN(n15045) );
  NAND3_X1 U16308 ( .A1(n15047), .A2(n15046), .A3(n15045), .ZN(P1_U3254) );
  NAND2_X1 U16309 ( .A1(n15059), .A2(n15051), .ZN(n15052) );
  XNOR2_X1 U16310 ( .A(n16267), .B(n15051), .ZN(n16260) );
  NAND2_X1 U16311 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n16260), .ZN(n16259) );
  INV_X1 U16312 ( .A(n15053), .ZN(n15057) );
  INV_X1 U16313 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n15054) );
  OAI22_X1 U16314 ( .A1(n15057), .A2(n15056), .B1(n15055), .B2(n15054), .ZN(
        n15058) );
  NAND2_X1 U16315 ( .A1(n15059), .A2(n15058), .ZN(n15060) );
  XOR2_X1 U16316 ( .A(n15059), .B(n15058), .Z(n16262) );
  NAND2_X1 U16317 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n16262), .ZN(n16261) );
  NAND2_X1 U16318 ( .A1(n15060), .A2(n16261), .ZN(n15061) );
  XOR2_X1 U16319 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n15061), .Z(n15062) );
  AOI22_X1 U16320 ( .A1(n15063), .A2(n16354), .B1(n16347), .B2(n15062), .ZN(
        n15069) );
  INV_X1 U16321 ( .A(n15062), .ZN(n15066) );
  NOR2_X1 U16322 ( .A1(n15063), .A2(n16266), .ZN(n15064) );
  AOI211_X1 U16323 ( .C1(n15067), .C2(n15066), .A(n15065), .B(n15064), .ZN(
        n15068) );
  MUX2_X1 U16324 ( .A(n15069), .B(n15068), .S(n15185), .Z(n15071) );
  OAI211_X1 U16325 ( .C1(n15072), .C2(n16364), .A(n15071), .B(n15070), .ZN(
        P1_U3262) );
  INV_X1 U16326 ( .A(n15351), .ZN(n15078) );
  NOR2_X1 U16327 ( .A1(n15080), .A2(n15081), .ZN(n15079) );
  XNOR2_X1 U16328 ( .A(n15079), .B(n15351), .ZN(n15354) );
  NAND2_X1 U16329 ( .A1(n15354), .A2(n15347), .ZN(n15077) );
  NAND2_X1 U16330 ( .A1(n15073), .A2(P1_B_REG_SCAN_IN), .ZN(n15074) );
  NAND2_X1 U16331 ( .A1(n15329), .A2(n15074), .ZN(n15096) );
  OR2_X1 U16332 ( .A1(n15075), .A2(n15096), .ZN(n15358) );
  NOR2_X1 U16333 ( .A1(n15333), .A2(n15358), .ZN(n15082) );
  AOI21_X1 U16334 ( .B1(n15295), .B2(P1_REG2_REG_31__SCAN_IN), .A(n15082), 
        .ZN(n15076) );
  OAI211_X1 U16335 ( .C1(n15078), .C2(n15310), .A(n15077), .B(n15076), .ZN(
        P1_U3263) );
  INV_X1 U16336 ( .A(n15081), .ZN(n15360) );
  AOI21_X1 U16337 ( .B1(n15081), .B2(n15080), .A(n15079), .ZN(n15357) );
  NAND2_X1 U16338 ( .A1(n15357), .A2(n15347), .ZN(n15084) );
  AOI21_X1 U16339 ( .B1(n15333), .B2(P1_REG2_REG_30__SCAN_IN), .A(n15082), 
        .ZN(n15083) );
  OAI211_X1 U16340 ( .C1(n15360), .C2(n15310), .A(n15084), .B(n15083), .ZN(
        P1_U3264) );
  NAND2_X1 U16341 ( .A1(n15371), .A2(n15085), .ZN(n15086) );
  NAND2_X1 U16342 ( .A1(n15087), .A2(n15086), .ZN(n15088) );
  XNOR2_X1 U16343 ( .A(n15088), .B(n15092), .ZN(n15362) );
  INV_X1 U16344 ( .A(n15362), .ZN(n15106) );
  XNOR2_X1 U16345 ( .A(n15094), .B(n15093), .ZN(n15363) );
  NOR2_X1 U16346 ( .A1(n15363), .A2(n15221), .ZN(n15104) );
  INV_X1 U16347 ( .A(n15095), .ZN(n15097) );
  OR2_X1 U16348 ( .A1(n15097), .A2(n15096), .ZN(n15365) );
  OAI22_X1 U16349 ( .A1(n15099), .A2(n15365), .B1(n15098), .B2(n15312), .ZN(
        n15101) );
  OR2_X1 U16350 ( .A1(n15112), .A2(n15230), .ZN(n15364) );
  NOR2_X1 U16351 ( .A1(n15333), .A2(n15364), .ZN(n15100) );
  AOI211_X1 U16352 ( .C1(n15295), .C2(P1_REG2_REG_29__SCAN_IN), .A(n15101), 
        .B(n15100), .ZN(n15102) );
  OAI21_X1 U16353 ( .B1(n15366), .B2(n15310), .A(n15102), .ZN(n15103) );
  AOI211_X1 U16354 ( .C1(n15368), .C2(n15265), .A(n15104), .B(n15103), .ZN(
        n15105) );
  OAI21_X1 U16355 ( .B1(n15106), .B2(n15337), .A(n15105), .ZN(P1_U3356) );
  OAI21_X1 U16356 ( .B1(n15108), .B2(n15110), .A(n15107), .ZN(n15379) );
  OAI22_X1 U16357 ( .A1(n15112), .A2(n15232), .B1(n15111), .B2(n15230), .ZN(
        n15113) );
  INV_X1 U16358 ( .A(n15114), .ZN(n15115) );
  OAI21_X1 U16359 ( .B1(n15376), .B2(n15124), .A(n15115), .ZN(n15377) );
  NOR2_X1 U16360 ( .A1(n15377), .A2(n15221), .ZN(n15120) );
  INV_X1 U16361 ( .A(n15116), .ZN(n15117) );
  AOI22_X1 U16362 ( .A1(n15295), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n15117), 
        .B2(n15341), .ZN(n15118) );
  OAI21_X1 U16363 ( .B1(n15376), .B2(n15310), .A(n15118), .ZN(n15119) );
  AOI211_X1 U16364 ( .C1(n15379), .C2(n15345), .A(n15120), .B(n15119), .ZN(
        n15121) );
  OAI21_X1 U16365 ( .B1(n15381), .B2(n15333), .A(n15121), .ZN(P1_U3266) );
  XNOR2_X1 U16366 ( .A(n15123), .B(n15122), .ZN(n15386) );
  AOI21_X1 U16367 ( .B1(n15382), .B2(n15145), .A(n15124), .ZN(n15383) );
  NOR2_X1 U16368 ( .A1(n15125), .A2(n15310), .ZN(n15129) );
  OAI22_X1 U16369 ( .A1(n15338), .A2(n15127), .B1(n15126), .B2(n15312), .ZN(
        n15128) );
  AOI211_X1 U16370 ( .C1(n15383), .C2(n15347), .A(n15129), .B(n15128), .ZN(
        n15136) );
  XNOR2_X1 U16371 ( .A(n15131), .B(n15130), .ZN(n15134) );
  AOI222_X1 U16372 ( .A1(n15431), .A2(n15134), .B1(n15133), .B2(n15329), .C1(
        n15132), .C2(n15331), .ZN(n15385) );
  OR2_X1 U16373 ( .A1(n15385), .A2(n15295), .ZN(n15135) );
  OAI211_X1 U16374 ( .C1(n15386), .C2(n15337), .A(n15136), .B(n15135), .ZN(
        P1_U3267) );
  OAI21_X1 U16375 ( .B1(n15138), .B2(n15143), .A(n15137), .ZN(n15139) );
  INV_X1 U16376 ( .A(n15139), .ZN(n15394) );
  INV_X1 U16377 ( .A(n15140), .ZN(n15141) );
  AOI21_X1 U16378 ( .B1(n15143), .B2(n15142), .A(n15141), .ZN(n15392) );
  NAND2_X1 U16379 ( .A1(n15388), .A2(n15170), .ZN(n15144) );
  NAND2_X1 U16380 ( .A1(n15145), .A2(n15144), .ZN(n15390) );
  NOR2_X1 U16381 ( .A1(n15390), .A2(n15221), .ZN(n15155) );
  NAND2_X1 U16382 ( .A1(n15146), .A2(n15331), .ZN(n15149) );
  NAND2_X1 U16383 ( .A1(n15147), .A2(n15329), .ZN(n15148) );
  NAND2_X1 U16384 ( .A1(n15149), .A2(n15148), .ZN(n15387) );
  INV_X1 U16385 ( .A(n15150), .ZN(n15151) );
  AOI22_X1 U16386 ( .A1(n15338), .A2(n15387), .B1(n15151), .B2(n15341), .ZN(
        n15153) );
  NAND2_X1 U16387 ( .A1(n15295), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n15152) );
  OAI211_X1 U16388 ( .C1(n8011), .C2(n15310), .A(n15153), .B(n15152), .ZN(
        n15154) );
  AOI211_X1 U16389 ( .C1(n15392), .C2(n15309), .A(n15155), .B(n15154), .ZN(
        n15156) );
  OAI21_X1 U16390 ( .B1(n15394), .B2(n15211), .A(n15156), .ZN(P1_U3268) );
  OAI21_X1 U16391 ( .B1(n15158), .B2(n15161), .A(n15157), .ZN(n15167) );
  INV_X1 U16392 ( .A(n15167), .ZN(n15399) );
  AOI211_X1 U16393 ( .C1(n15161), .C2(n15160), .A(n16449), .B(n15159), .ZN(
        n15165) );
  OAI22_X1 U16394 ( .A1(n15163), .A2(n15230), .B1(n15162), .B2(n15232), .ZN(
        n15164) );
  AOI211_X1 U16395 ( .C1(n15167), .C2(n15166), .A(n15165), .B(n15164), .ZN(
        n15398) );
  OAI21_X1 U16396 ( .B1(n15168), .B2(n15312), .A(n15398), .ZN(n15169) );
  NAND2_X1 U16397 ( .A1(n15169), .A2(n15338), .ZN(n15176) );
  AOI21_X1 U16398 ( .B1(n15395), .B2(n15171), .A(n8012), .ZN(n15396) );
  OAI22_X1 U16399 ( .A1(n15173), .A2(n15310), .B1(n15172), .B2(n15338), .ZN(
        n15174) );
  AOI21_X1 U16400 ( .B1(n15396), .B2(n15347), .A(n15174), .ZN(n15175) );
  OAI211_X1 U16401 ( .C1(n15399), .C2(n15177), .A(n15176), .B(n15175), .ZN(
        P1_U3269) );
  XNOR2_X1 U16402 ( .A(n15178), .B(n15180), .ZN(n15405) );
  OAI21_X1 U16403 ( .B1(n15181), .B2(n15180), .A(n15179), .ZN(n15182) );
  AND2_X1 U16404 ( .A1(n15182), .A2(n15431), .ZN(n15404) );
  XNOR2_X1 U16405 ( .A(n15197), .B(n15183), .ZN(n15184) );
  NAND2_X1 U16406 ( .A1(n15184), .A2(n15471), .ZN(n15401) );
  OAI21_X1 U16407 ( .B1(n15401), .B2(n15185), .A(n15400), .ZN(n15186) );
  OAI21_X1 U16408 ( .B1(n15404), .B2(n15186), .A(n15338), .ZN(n15189) );
  AOI22_X1 U16409 ( .A1(n15295), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n15187), 
        .B2(n15341), .ZN(n15188) );
  OAI211_X1 U16410 ( .C1(n15402), .C2(n15310), .A(n15189), .B(n15188), .ZN(
        n15190) );
  AOI21_X1 U16411 ( .B1(n15405), .B2(n15309), .A(n15190), .ZN(n15191) );
  INV_X1 U16412 ( .A(n15191), .ZN(P1_U3270) );
  INV_X1 U16413 ( .A(n15194), .ZN(n15192) );
  XNOR2_X1 U16414 ( .A(n15193), .B(n15192), .ZN(n15414) );
  XNOR2_X1 U16415 ( .A(n15195), .B(n15194), .ZN(n15412) );
  NAND2_X1 U16416 ( .A1(n15412), .A2(n15309), .ZN(n15210) );
  AND2_X1 U16417 ( .A1(n15408), .A2(n15220), .ZN(n15196) );
  OR2_X1 U16418 ( .A1(n15197), .A2(n15196), .ZN(n15410) );
  INV_X1 U16419 ( .A(n15410), .ZN(n15208) );
  NAND2_X1 U16420 ( .A1(n15198), .A2(n15329), .ZN(n15201) );
  NAND2_X1 U16421 ( .A1(n15199), .A2(n15331), .ZN(n15200) );
  NAND2_X1 U16422 ( .A1(n15201), .A2(n15200), .ZN(n15407) );
  INV_X1 U16423 ( .A(n15202), .ZN(n15203) );
  AOI22_X1 U16424 ( .A1(n15407), .A2(n15338), .B1(n15203), .B2(n15341), .ZN(
        n15205) );
  NAND2_X1 U16425 ( .A1(n15295), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n15204) );
  OAI211_X1 U16426 ( .C1(n15206), .C2(n15310), .A(n15205), .B(n15204), .ZN(
        n15207) );
  AOI21_X1 U16427 ( .B1(n15208), .B2(n15347), .A(n15207), .ZN(n15209) );
  OAI211_X1 U16428 ( .C1(n15414), .C2(n15211), .A(n15210), .B(n15209), .ZN(
        P1_U3271) );
  XNOR2_X1 U16429 ( .A(n15213), .B(n15212), .ZN(n15215) );
  OAI222_X1 U16430 ( .A1(n15232), .A2(n7885), .B1(n15215), .B2(n16449), .C1(
        n15230), .C2(n15214), .ZN(n15417) );
  INV_X1 U16431 ( .A(n15417), .ZN(n15227) );
  OAI21_X1 U16432 ( .B1(n15218), .B2(n15217), .A(n15216), .ZN(n15418) );
  OR2_X1 U16433 ( .A1(n15240), .A2(n8453), .ZN(n15219) );
  NAND2_X1 U16434 ( .A1(n15220), .A2(n15219), .ZN(n15415) );
  NOR2_X1 U16435 ( .A1(n15415), .A2(n15221), .ZN(n15225) );
  AOI22_X1 U16436 ( .A1(n15295), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n15222), 
        .B2(n15341), .ZN(n15223) );
  OAI21_X1 U16437 ( .B1(n8453), .B2(n15310), .A(n15223), .ZN(n15224) );
  AOI211_X1 U16438 ( .C1(n15418), .C2(n15309), .A(n15225), .B(n15224), .ZN(
        n15226) );
  OAI21_X1 U16439 ( .B1(n15295), .B2(n15227), .A(n15226), .ZN(P1_U3272) );
  AOI21_X1 U16440 ( .B1(n15229), .B2(n15228), .A(n16449), .ZN(n15236) );
  OAI22_X1 U16441 ( .A1(n15233), .A2(n15232), .B1(n15231), .B2(n15230), .ZN(
        n15234) );
  AOI21_X1 U16442 ( .B1(n15236), .B2(n15235), .A(n15234), .ZN(n15424) );
  INV_X1 U16443 ( .A(n15426), .ZN(n15239) );
  NAND2_X1 U16444 ( .A1(n15238), .A2(n15237), .ZN(n15420) );
  NAND3_X1 U16445 ( .A1(n15239), .A2(n15309), .A3(n15420), .ZN(n15247) );
  AOI21_X1 U16446 ( .B1(n15421), .B2(n15254), .A(n15240), .ZN(n15422) );
  INV_X1 U16447 ( .A(n15241), .ZN(n15242) );
  AOI22_X1 U16448 ( .A1(n15295), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n15242), 
        .B2(n15341), .ZN(n15243) );
  OAI21_X1 U16449 ( .B1(n15244), .B2(n15310), .A(n15243), .ZN(n15245) );
  AOI21_X1 U16450 ( .B1(n15422), .B2(n15347), .A(n15245), .ZN(n15246) );
  OAI211_X1 U16451 ( .C1(n15333), .C2(n15424), .A(n15247), .B(n15246), .ZN(
        P1_U3273) );
  XNOR2_X1 U16452 ( .A(n15249), .B(n15248), .ZN(n15434) );
  INV_X1 U16453 ( .A(n15250), .ZN(n15253) );
  OAI21_X1 U16454 ( .B1(n15253), .B2(n15252), .A(n15251), .ZN(n15432) );
  INV_X1 U16455 ( .A(n15254), .ZN(n15255) );
  AOI21_X1 U16456 ( .B1(n15257), .B2(n15256), .A(n15255), .ZN(n15427) );
  NAND2_X1 U16457 ( .A1(n15427), .A2(n15347), .ZN(n15263) );
  AOI22_X1 U16458 ( .A1(n15258), .A2(n15329), .B1(n15331), .B2(n15289), .ZN(
        n15428) );
  INV_X1 U16459 ( .A(n15259), .ZN(n15260) );
  OAI22_X1 U16460 ( .A1(n15295), .A2(n15428), .B1(n15260), .B2(n15312), .ZN(
        n15261) );
  AOI21_X1 U16461 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(n15333), .A(n15261), 
        .ZN(n15262) );
  OAI211_X1 U16462 ( .C1(n8482), .C2(n15310), .A(n15263), .B(n15262), .ZN(
        n15264) );
  AOI21_X1 U16463 ( .B1(n15432), .B2(n15265), .A(n15264), .ZN(n15266) );
  OAI21_X1 U16464 ( .B1(n15434), .B2(n15337), .A(n15266), .ZN(P1_U3274) );
  XNOR2_X1 U16465 ( .A(n15268), .B(n15267), .ZN(n15269) );
  AOI222_X1 U16466 ( .A1(n15304), .A2(n15331), .B1(n15270), .B2(n15329), .C1(
        n15431), .C2(n15269), .ZN(n15438) );
  XNOR2_X1 U16467 ( .A(n15274), .B(n15293), .ZN(n15436) );
  INV_X1 U16468 ( .A(n15271), .ZN(n15272) );
  AOI22_X1 U16469 ( .A1(n15295), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n15272), 
        .B2(n15341), .ZN(n15273) );
  OAI21_X1 U16470 ( .B1(n15274), .B2(n15310), .A(n15273), .ZN(n15278) );
  XNOR2_X1 U16471 ( .A(n15276), .B(n15275), .ZN(n15439) );
  NOR2_X1 U16472 ( .A1(n15439), .A2(n15337), .ZN(n15277) );
  AOI211_X1 U16473 ( .C1(n15436), .C2(n15347), .A(n15278), .B(n15277), .ZN(
        n15279) );
  OAI21_X1 U16474 ( .B1(n15295), .B2(n15438), .A(n15279), .ZN(P1_U3275) );
  AOI21_X1 U16475 ( .B1(n15282), .B2(n15281), .A(n15280), .ZN(n15283) );
  INV_X1 U16476 ( .A(n15283), .ZN(n15444) );
  INV_X1 U16477 ( .A(n15302), .ZN(n15286) );
  OAI21_X1 U16478 ( .B1(n15286), .B2(n15285), .A(n15284), .ZN(n15288) );
  NAND3_X1 U16479 ( .A1(n15288), .A2(n15431), .A3(n15287), .ZN(n15291) );
  AOI22_X1 U16480 ( .A1(n15289), .A2(n15329), .B1(n15331), .B2(n15330), .ZN(
        n15290) );
  AND2_X1 U16481 ( .A1(n15291), .A2(n15290), .ZN(n15443) );
  INV_X1 U16482 ( .A(n15443), .ZN(n15300) );
  OR2_X1 U16483 ( .A1(n15298), .A2(n7595), .ZN(n15292) );
  AND2_X1 U16484 ( .A1(n15293), .A2(n15292), .ZN(n15441) );
  NAND2_X1 U16485 ( .A1(n15441), .A2(n15347), .ZN(n15297) );
  AOI22_X1 U16486 ( .A1(n15295), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n15294), 
        .B2(n15341), .ZN(n15296) );
  OAI211_X1 U16487 ( .C1(n15298), .C2(n15310), .A(n15297), .B(n15296), .ZN(
        n15299) );
  AOI21_X1 U16488 ( .B1(n15300), .B2(n15338), .A(n15299), .ZN(n15301) );
  OAI21_X1 U16489 ( .B1(n15444), .B2(n15337), .A(n15301), .ZN(P1_U3276) );
  OAI21_X1 U16490 ( .B1(n7598), .B2(n8430), .A(n15302), .ZN(n15305) );
  AOI222_X1 U16491 ( .A1(n15431), .A2(n15305), .B1(n15304), .B2(n15329), .C1(
        n15303), .C2(n15331), .ZN(n15449) );
  OAI21_X1 U16492 ( .B1(n15308), .B2(n15307), .A(n15306), .ZN(n15445) );
  NAND2_X1 U16493 ( .A1(n15445), .A2(n15309), .ZN(n15317) );
  AOI21_X1 U16494 ( .B1(n15446), .B2(n15319), .A(n7595), .ZN(n15447) );
  NOR2_X1 U16495 ( .A1(n15311), .A2(n15310), .ZN(n15315) );
  OAI22_X1 U16496 ( .A1(n15338), .A2(n11578), .B1(n15313), .B2(n15312), .ZN(
        n15314) );
  AOI211_X1 U16497 ( .C1(n15447), .C2(n15347), .A(n15315), .B(n15314), .ZN(
        n15316) );
  OAI211_X1 U16498 ( .C1(n15333), .C2(n15449), .A(n15317), .B(n15316), .ZN(
        P1_U3277) );
  XOR2_X1 U16499 ( .A(n15318), .B(n15327), .Z(n15455) );
  INV_X1 U16500 ( .A(n15319), .ZN(n15320) );
  AOI21_X1 U16501 ( .B1(n15451), .B2(n15321), .A(n15320), .ZN(n15452) );
  INV_X1 U16502 ( .A(n15322), .ZN(n15323) );
  AOI22_X1 U16503 ( .A1(n15333), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n15323), 
        .B2(n15341), .ZN(n15324) );
  OAI21_X1 U16504 ( .B1(n15325), .B2(n15310), .A(n15324), .ZN(n15335) );
  XOR2_X1 U16505 ( .A(n15327), .B(n15326), .Z(n15328) );
  AOI222_X1 U16506 ( .A1(n15332), .A2(n15331), .B1(n15330), .B2(n15329), .C1(
        n15431), .C2(n15328), .ZN(n15454) );
  NOR2_X1 U16507 ( .A1(n15454), .A2(n15333), .ZN(n15334) );
  AOI211_X1 U16508 ( .C1(n15452), .C2(n15347), .A(n15335), .B(n15334), .ZN(
        n15336) );
  OAI21_X1 U16509 ( .B1(n15455), .B2(n15337), .A(n15336), .ZN(P1_U3278) );
  MUX2_X1 U16510 ( .A(n15340), .B(n15339), .S(n15338), .Z(n15350) );
  AOI22_X1 U16511 ( .A1(n15343), .A2(n15342), .B1(n15341), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n15349) );
  AOI22_X1 U16512 ( .A1(n15347), .A2(n15346), .B1(n15345), .B2(n15344), .ZN(
        n15348) );
  NAND3_X1 U16513 ( .A1(n15350), .A2(n15349), .A3(n15348), .ZN(P1_U3291) );
  NAND2_X1 U16514 ( .A1(n15351), .A2(n16445), .ZN(n15352) );
  NAND2_X1 U16515 ( .A1(n15352), .A2(n15358), .ZN(n15353) );
  AOI21_X1 U16516 ( .B1(n15354), .B2(n15471), .A(n15353), .ZN(n15477) );
  MUX2_X1 U16517 ( .A(n15355), .B(n15477), .S(n16553), .Z(n15356) );
  INV_X1 U16518 ( .A(n15356), .ZN(P1_U3559) );
  NAND2_X1 U16519 ( .A1(n15357), .A2(n15471), .ZN(n15359) );
  OAI211_X1 U16520 ( .C1(n15360), .C2(n16542), .A(n15359), .B(n15358), .ZN(
        n15480) );
  MUX2_X1 U16521 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15480), .S(n16553), .Z(
        P1_U3558) );
  NAND2_X1 U16522 ( .A1(n15362), .A2(n16547), .ZN(n15369) );
  OAI211_X1 U16523 ( .C1(n15366), .C2(n16542), .A(n15365), .B(n15364), .ZN(
        n15367) );
  MUX2_X1 U16524 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n15481), .S(n16553), .Z(
        P1_U3557) );
  NAND2_X1 U16525 ( .A1(n15370), .A2(n16547), .ZN(n15375) );
  AOI22_X1 U16526 ( .A1(n15372), .A2(n15471), .B1(n15371), .B2(n16445), .ZN(
        n15373) );
  MUX2_X1 U16527 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15482), .S(n16553), .Z(
        P1_U3556) );
  INV_X1 U16528 ( .A(n15475), .ZN(n16495) );
  OAI22_X1 U16529 ( .A1(n15377), .A2(n16544), .B1(n15376), .B2(n16542), .ZN(
        n15378) );
  AOI21_X1 U16530 ( .B1(n15379), .B2(n16495), .A(n15378), .ZN(n15380) );
  MUX2_X1 U16531 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n15483), .S(n16553), .Z(
        P1_U3555) );
  AOI22_X1 U16532 ( .A1(n15383), .A2(n15471), .B1(n15382), .B2(n16445), .ZN(
        n15384) );
  OAI211_X1 U16533 ( .C1(n15386), .C2(n15463), .A(n15385), .B(n15384), .ZN(
        n15484) );
  MUX2_X1 U16534 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15484), .S(n16553), .Z(
        P1_U3554) );
  AOI21_X1 U16535 ( .B1(n15388), .B2(n16445), .A(n15387), .ZN(n15389) );
  OAI21_X1 U16536 ( .B1(n15390), .B2(n16544), .A(n15389), .ZN(n15391) );
  AOI21_X1 U16537 ( .B1(n15392), .B2(n16547), .A(n15391), .ZN(n15393) );
  OAI21_X1 U16538 ( .B1(n16449), .B2(n15394), .A(n15393), .ZN(n15485) );
  MUX2_X1 U16539 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n15485), .S(n16553), .Z(
        P1_U3553) );
  AOI22_X1 U16540 ( .A1(n15396), .A2(n15471), .B1(n15395), .B2(n16445), .ZN(
        n15397) );
  OAI211_X1 U16541 ( .C1(n15399), .C2(n15475), .A(n15398), .B(n15397), .ZN(
        n15486) );
  MUX2_X1 U16542 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n15486), .S(n16553), .Z(
        P1_U3552) );
  OAI211_X1 U16543 ( .C1(n15402), .C2(n16542), .A(n15401), .B(n15400), .ZN(
        n15403) );
  AOI211_X1 U16544 ( .C1(n15405), .C2(n16547), .A(n15404), .B(n15403), .ZN(
        n15406) );
  INV_X1 U16545 ( .A(n15406), .ZN(n15487) );
  MUX2_X1 U16546 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15487), .S(n16553), .Z(
        P1_U3551) );
  AOI21_X1 U16547 ( .B1(n15408), .B2(n16445), .A(n15407), .ZN(n15409) );
  OAI21_X1 U16548 ( .B1(n15410), .B2(n16544), .A(n15409), .ZN(n15411) );
  AOI21_X1 U16549 ( .B1(n15412), .B2(n16547), .A(n15411), .ZN(n15413) );
  OAI21_X1 U16550 ( .B1(n16449), .B2(n15414), .A(n15413), .ZN(n15488) );
  MUX2_X1 U16551 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15488), .S(n16553), .Z(
        P1_U3550) );
  OAI22_X1 U16552 ( .A1(n15415), .A2(n16544), .B1(n8453), .B2(n16542), .ZN(
        n15416) );
  AOI211_X1 U16553 ( .C1(n15418), .C2(n16547), .A(n15417), .B(n15416), .ZN(
        n15419) );
  INV_X1 U16554 ( .A(n15419), .ZN(n15489) );
  MUX2_X1 U16555 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15489), .S(n16553), .Z(
        P1_U3549) );
  NAND2_X1 U16556 ( .A1(n15420), .A2(n16547), .ZN(n15425) );
  AOI22_X1 U16557 ( .A1(n15422), .A2(n15471), .B1(n15421), .B2(n16445), .ZN(
        n15423) );
  OAI211_X1 U16558 ( .C1(n15426), .C2(n15425), .A(n15424), .B(n15423), .ZN(
        n15490) );
  MUX2_X1 U16559 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15490), .S(n16553), .Z(
        P1_U3548) );
  NAND2_X1 U16560 ( .A1(n15427), .A2(n15471), .ZN(n15429) );
  OAI211_X1 U16561 ( .C1(n8482), .C2(n16542), .A(n15429), .B(n15428), .ZN(
        n15430) );
  AOI21_X1 U16562 ( .B1(n15432), .B2(n15431), .A(n15430), .ZN(n15433) );
  OAI21_X1 U16563 ( .B1(n15434), .B2(n15463), .A(n15433), .ZN(n15491) );
  MUX2_X1 U16564 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15491), .S(n16553), .Z(
        P1_U3547) );
  AOI22_X1 U16565 ( .A1(n15436), .A2(n15471), .B1(n15435), .B2(n16445), .ZN(
        n15437) );
  OAI211_X1 U16566 ( .C1(n15439), .C2(n15463), .A(n15438), .B(n15437), .ZN(
        n15492) );
  MUX2_X1 U16567 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15492), .S(n16553), .Z(
        P1_U3546) );
  AOI22_X1 U16568 ( .A1(n15441), .A2(n15471), .B1(n15440), .B2(n16445), .ZN(
        n15442) );
  OAI211_X1 U16569 ( .C1(n15444), .C2(n15463), .A(n15443), .B(n15442), .ZN(
        n15493) );
  MUX2_X1 U16570 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15493), .S(n16553), .Z(
        P1_U3545) );
  INV_X1 U16571 ( .A(n15445), .ZN(n15450) );
  AOI22_X1 U16572 ( .A1(n15447), .A2(n15471), .B1(n15446), .B2(n16445), .ZN(
        n15448) );
  OAI211_X1 U16573 ( .C1(n15450), .C2(n15463), .A(n15449), .B(n15448), .ZN(
        n15494) );
  MUX2_X1 U16574 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n15494), .S(n16553), .Z(
        P1_U3544) );
  AOI22_X1 U16575 ( .A1(n15452), .A2(n15471), .B1(n15451), .B2(n16445), .ZN(
        n15453) );
  OAI211_X1 U16576 ( .C1(n15455), .C2(n15463), .A(n15454), .B(n15453), .ZN(
        n15896) );
  MUX2_X1 U16577 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15896), .S(n16553), .Z(
        P1_U3543) );
  AOI22_X1 U16578 ( .A1(n15457), .A2(n15471), .B1(n15456), .B2(n16445), .ZN(
        n15458) );
  OAI211_X1 U16579 ( .C1(n15460), .C2(n15463), .A(n15459), .B(n15458), .ZN(
        n15899) );
  MUX2_X1 U16580 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15899), .S(n16553), .Z(
        P1_U3542) );
  OAI21_X1 U16581 ( .B1(n15462), .B2(n16542), .A(n15461), .ZN(n15466) );
  NOR2_X1 U16582 ( .A1(n15464), .A2(n15463), .ZN(n15465) );
  AOI211_X1 U16583 ( .C1(n15471), .C2(n15467), .A(n15466), .B(n15465), .ZN(
        n15468) );
  OAI21_X1 U16584 ( .B1(n16449), .B2(n15469), .A(n15468), .ZN(n15900) );
  MUX2_X1 U16585 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15900), .S(n16553), .Z(
        P1_U3541) );
  AOI22_X1 U16586 ( .A1(n15472), .A2(n15471), .B1(n15470), .B2(n16445), .ZN(
        n15473) );
  OAI211_X1 U16587 ( .C1(n15476), .C2(n15475), .A(n15474), .B(n15473), .ZN(
        n15901) );
  MUX2_X1 U16588 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n15901), .S(n16553), .Z(
        P1_U3540) );
  MUX2_X1 U16589 ( .A(n15478), .B(n15477), .S(n16556), .Z(n15479) );
  INV_X1 U16590 ( .A(n15479), .ZN(P1_U3527) );
  MUX2_X1 U16591 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15480), .S(n16556), .Z(
        P1_U3526) );
  MUX2_X1 U16592 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n15481), .S(n16556), .Z(
        P1_U3525) );
  MUX2_X1 U16593 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15482), .S(n16556), .Z(
        P1_U3524) );
  MUX2_X1 U16594 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n15483), .S(n16556), .Z(
        P1_U3523) );
  MUX2_X1 U16595 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15484), .S(n16556), .Z(
        P1_U3522) );
  MUX2_X1 U16596 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n15485), .S(n16556), .Z(
        P1_U3521) );
  MUX2_X1 U16597 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n15486), .S(n16556), .Z(
        P1_U3520) );
  MUX2_X1 U16598 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15487), .S(n16556), .Z(
        P1_U3519) );
  MUX2_X1 U16599 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15488), .S(n16556), .Z(
        P1_U3518) );
  MUX2_X1 U16600 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15489), .S(n16556), .Z(
        P1_U3517) );
  MUX2_X1 U16601 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15490), .S(n16556), .Z(
        P1_U3516) );
  MUX2_X1 U16602 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15491), .S(n16556), .Z(
        P1_U3515) );
  MUX2_X1 U16603 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15492), .S(n16556), .Z(
        P1_U3513) );
  MUX2_X1 U16604 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15493), .S(n16556), .Z(
        P1_U3510) );
  MUX2_X1 U16605 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n15494), .S(n16556), .Z(
        P1_U3507) );
  XNOR2_X1 U16606 ( .A(keyinput_128), .B(P3_WR_REG_SCAN_IN), .ZN(n15497) );
  XNOR2_X1 U16607 ( .A(SI_31_), .B(keyinput_129), .ZN(n15496) );
  XOR2_X1 U16608 ( .A(SI_30_), .B(keyinput_130), .Z(n15495) );
  OAI21_X1 U16609 ( .B1(n15497), .B2(n15496), .A(n15495), .ZN(n15501) );
  XNOR2_X1 U16610 ( .A(SI_29_), .B(keyinput_131), .ZN(n15500) );
  XNOR2_X1 U16611 ( .A(n15498), .B(keyinput_132), .ZN(n15499) );
  AOI21_X1 U16612 ( .B1(n15501), .B2(n15500), .A(n15499), .ZN(n15505) );
  XNOR2_X1 U16613 ( .A(n15502), .B(keyinput_134), .ZN(n15504) );
  XNOR2_X1 U16614 ( .A(SI_27_), .B(keyinput_133), .ZN(n15503) );
  NOR3_X1 U16615 ( .A1(n15505), .A2(n15504), .A3(n15503), .ZN(n15508) );
  XNOR2_X1 U16616 ( .A(n15704), .B(keyinput_135), .ZN(n15507) );
  XNOR2_X1 U16617 ( .A(SI_24_), .B(keyinput_136), .ZN(n15506) );
  NOR3_X1 U16618 ( .A1(n15508), .A2(n15507), .A3(n15506), .ZN(n15511) );
  XOR2_X1 U16619 ( .A(SI_23_), .B(keyinput_137), .Z(n15510) );
  XOR2_X1 U16620 ( .A(SI_22_), .B(keyinput_138), .Z(n15509) );
  NOR3_X1 U16621 ( .A1(n15511), .A2(n15510), .A3(n15509), .ZN(n15516) );
  XNOR2_X1 U16622 ( .A(n15512), .B(keyinput_141), .ZN(n15515) );
  XNOR2_X1 U16623 ( .A(SI_20_), .B(keyinput_140), .ZN(n15514) );
  XNOR2_X1 U16624 ( .A(SI_21_), .B(keyinput_139), .ZN(n15513) );
  NOR4_X1 U16625 ( .A1(n15516), .A2(n15515), .A3(n15514), .A4(n15513), .ZN(
        n15519) );
  XNOR2_X1 U16626 ( .A(n15716), .B(keyinput_142), .ZN(n15518) );
  XNOR2_X1 U16627 ( .A(n15717), .B(keyinput_143), .ZN(n15517) );
  OAI21_X1 U16628 ( .B1(n15519), .B2(n15518), .A(n15517), .ZN(n15524) );
  XNOR2_X1 U16629 ( .A(n15520), .B(keyinput_144), .ZN(n15523) );
  XNOR2_X1 U16630 ( .A(n15521), .B(keyinput_145), .ZN(n15522) );
  AOI21_X1 U16631 ( .B1(n15524), .B2(n15523), .A(n15522), .ZN(n15528) );
  XNOR2_X1 U16632 ( .A(n15525), .B(keyinput_146), .ZN(n15527) );
  XNOR2_X1 U16633 ( .A(SI_13_), .B(keyinput_147), .ZN(n15526) );
  OAI21_X1 U16634 ( .B1(n15528), .B2(n15527), .A(n15526), .ZN(n15531) );
  XNOR2_X1 U16635 ( .A(SI_12_), .B(keyinput_148), .ZN(n15530) );
  XNOR2_X1 U16636 ( .A(SI_11_), .B(keyinput_149), .ZN(n15529) );
  AOI21_X1 U16637 ( .B1(n15531), .B2(n15530), .A(n15529), .ZN(n15534) );
  XOR2_X1 U16638 ( .A(SI_9_), .B(keyinput_151), .Z(n15533) );
  XNOR2_X1 U16639 ( .A(SI_10_), .B(keyinput_150), .ZN(n15532) );
  NOR3_X1 U16640 ( .A1(n15534), .A2(n15533), .A3(n15532), .ZN(n15537) );
  XOR2_X1 U16641 ( .A(SI_8_), .B(keyinput_152), .Z(n15536) );
  XNOR2_X1 U16642 ( .A(SI_7_), .B(keyinput_153), .ZN(n15535) );
  OAI21_X1 U16643 ( .B1(n15537), .B2(n15536), .A(n15535), .ZN(n15540) );
  XOR2_X1 U16644 ( .A(SI_6_), .B(keyinput_154), .Z(n15539) );
  XOR2_X1 U16645 ( .A(SI_5_), .B(keyinput_155), .Z(n15538) );
  AOI21_X1 U16646 ( .B1(n15540), .B2(n15539), .A(n15538), .ZN(n15543) );
  XOR2_X1 U16647 ( .A(SI_3_), .B(keyinput_157), .Z(n15542) );
  XNOR2_X1 U16648 ( .A(SI_4_), .B(keyinput_156), .ZN(n15541) );
  NOR3_X1 U16649 ( .A1(n15543), .A2(n15542), .A3(n15541), .ZN(n15551) );
  XNOR2_X1 U16650 ( .A(n15544), .B(keyinput_158), .ZN(n15550) );
  XOR2_X1 U16651 ( .A(keyinput_161), .B(P3_RD_REG_SCAN_IN), .Z(n15548) );
  XNOR2_X1 U16652 ( .A(n15545), .B(keyinput_159), .ZN(n15547) );
  XNOR2_X1 U16653 ( .A(SI_0_), .B(keyinput_160), .ZN(n15546) );
  NOR3_X1 U16654 ( .A1(n15548), .A2(n15547), .A3(n15546), .ZN(n15549) );
  OAI21_X1 U16655 ( .B1(n15551), .B2(n15550), .A(n15549), .ZN(n15554) );
  XNOR2_X1 U16656 ( .A(P3_U3151), .B(keyinput_162), .ZN(n15553) );
  XNOR2_X1 U16657 ( .A(P3_REG3_REG_7__SCAN_IN), .B(keyinput_163), .ZN(n15552)
         );
  NAND3_X1 U16658 ( .A1(n15554), .A2(n15553), .A3(n15552), .ZN(n15557) );
  XOR2_X1 U16659 ( .A(P3_REG3_REG_14__SCAN_IN), .B(keyinput_165), .Z(n15556)
         );
  XNOR2_X1 U16660 ( .A(P3_REG3_REG_27__SCAN_IN), .B(keyinput_164), .ZN(n15555)
         );
  NAND3_X1 U16661 ( .A1(n15557), .A2(n15556), .A3(n15555), .ZN(n15561) );
  XOR2_X1 U16662 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput_166), .Z(n15560)
         );
  XNOR2_X1 U16663 ( .A(P3_REG3_REG_3__SCAN_IN), .B(keyinput_168), .ZN(n15559)
         );
  XNOR2_X1 U16664 ( .A(P3_REG3_REG_10__SCAN_IN), .B(keyinput_167), .ZN(n15558)
         );
  AOI211_X1 U16665 ( .C1(n15561), .C2(n15560), .A(n15559), .B(n15558), .ZN(
        n15568) );
  XOR2_X1 U16666 ( .A(P3_REG3_REG_19__SCAN_IN), .B(keyinput_169), .Z(n15567)
         );
  XOR2_X1 U16667 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_172), .Z(n15565) );
  XNOR2_X1 U16668 ( .A(n15761), .B(keyinput_173), .ZN(n15564) );
  XNOR2_X1 U16669 ( .A(P3_REG3_REG_28__SCAN_IN), .B(keyinput_170), .ZN(n15563)
         );
  XNOR2_X1 U16670 ( .A(P3_REG3_REG_8__SCAN_IN), .B(keyinput_171), .ZN(n15562)
         );
  NOR4_X1 U16671 ( .A1(n15565), .A2(n15564), .A3(n15563), .A4(n15562), .ZN(
        n15566) );
  OAI21_X1 U16672 ( .B1(n15568), .B2(n15567), .A(n15566), .ZN(n15571) );
  XOR2_X1 U16673 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput_174), .Z(n15570)
         );
  XNOR2_X1 U16674 ( .A(P3_REG3_REG_25__SCAN_IN), .B(keyinput_175), .ZN(n15569)
         );
  AOI21_X1 U16675 ( .B1(n15571), .B2(n15570), .A(n15569), .ZN(n15574) );
  XNOR2_X1 U16676 ( .A(P3_REG3_REG_16__SCAN_IN), .B(keyinput_176), .ZN(n15573)
         );
  XNOR2_X1 U16677 ( .A(P3_REG3_REG_5__SCAN_IN), .B(keyinput_177), .ZN(n15572)
         );
  OAI21_X1 U16678 ( .B1(n15574), .B2(n15573), .A(n15572), .ZN(n15580) );
  XNOR2_X1 U16679 ( .A(n15575), .B(keyinput_178), .ZN(n15579) );
  XOR2_X1 U16680 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput_180), .Z(n15578) );
  XNOR2_X1 U16681 ( .A(n15576), .B(keyinput_179), .ZN(n15577) );
  AOI211_X1 U16682 ( .C1(n15580), .C2(n15579), .A(n15578), .B(n15577), .ZN(
        n15583) );
  XNOR2_X1 U16683 ( .A(n15782), .B(keyinput_181), .ZN(n15582) );
  XNOR2_X1 U16684 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_182), .ZN(n15581)
         );
  NOR3_X1 U16685 ( .A1(n15583), .A2(n15582), .A3(n15581), .ZN(n15590) );
  AOI22_X1 U16686 ( .A1(n8771), .A2(keyinput_184), .B1(n15585), .B2(
        keyinput_185), .ZN(n15584) );
  OAI221_X1 U16687 ( .B1(n8771), .B2(keyinput_184), .C1(n15585), .C2(
        keyinput_185), .A(n15584), .ZN(n15589) );
  INV_X1 U16688 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n16404) );
  AOI22_X1 U16689 ( .A1(n16404), .A2(keyinput_187), .B1(n15788), .B2(
        keyinput_183), .ZN(n15586) );
  OAI221_X1 U16690 ( .B1(n16404), .B2(keyinput_187), .C1(n15788), .C2(
        keyinput_183), .A(n15586), .ZN(n15588) );
  XNOR2_X1 U16691 ( .A(P3_REG3_REG_11__SCAN_IN), .B(keyinput_186), .ZN(n15587)
         );
  NOR4_X1 U16692 ( .A1(n15590), .A2(n15589), .A3(n15588), .A4(n15587), .ZN(
        n15593) );
  XOR2_X1 U16693 ( .A(P3_REG3_REG_18__SCAN_IN), .B(keyinput_188), .Z(n15592)
         );
  XNOR2_X1 U16694 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput_189), .ZN(n15591)
         );
  NOR3_X1 U16695 ( .A1(n15593), .A2(n15592), .A3(n15591), .ZN(n15596) );
  XOR2_X1 U16696 ( .A(P3_REG3_REG_15__SCAN_IN), .B(keyinput_191), .Z(n15595)
         );
  XNOR2_X1 U16697 ( .A(n15795), .B(keyinput_190), .ZN(n15594) );
  NOR3_X1 U16698 ( .A1(n15596), .A2(n15595), .A3(n15594), .ZN(n15599) );
  XOR2_X1 U16699 ( .A(P3_B_REG_SCAN_IN), .B(keyinput_192), .Z(n15598) );
  XOR2_X1 U16700 ( .A(keyinput_193), .B(P3_DATAO_REG_31__SCAN_IN), .Z(n15597)
         );
  OAI21_X1 U16701 ( .B1(n15599), .B2(n15598), .A(n15597), .ZN(n15605) );
  XOR2_X1 U16702 ( .A(keyinput_194), .B(P3_DATAO_REG_30__SCAN_IN), .Z(n15604)
         );
  XOR2_X1 U16703 ( .A(keyinput_197), .B(P3_DATAO_REG_27__SCAN_IN), .Z(n15602)
         );
  XOR2_X1 U16704 ( .A(keyinput_196), .B(P3_DATAO_REG_28__SCAN_IN), .Z(n15601)
         );
  XNOR2_X1 U16705 ( .A(keyinput_195), .B(P3_DATAO_REG_29__SCAN_IN), .ZN(n15600) );
  NAND3_X1 U16706 ( .A1(n15602), .A2(n15601), .A3(n15600), .ZN(n15603) );
  AOI21_X1 U16707 ( .B1(n15605), .B2(n15604), .A(n15603), .ZN(n15608) );
  XOR2_X1 U16708 ( .A(keyinput_198), .B(P3_DATAO_REG_26__SCAN_IN), .Z(n15607)
         );
  XNOR2_X1 U16709 ( .A(keyinput_199), .B(P3_DATAO_REG_25__SCAN_IN), .ZN(n15606) );
  OAI21_X1 U16710 ( .B1(n15608), .B2(n15607), .A(n15606), .ZN(n15612) );
  XOR2_X1 U16711 ( .A(keyinput_200), .B(P3_DATAO_REG_24__SCAN_IN), .Z(n15611)
         );
  XOR2_X1 U16712 ( .A(keyinput_201), .B(P3_DATAO_REG_23__SCAN_IN), .Z(n15610)
         );
  XOR2_X1 U16713 ( .A(keyinput_202), .B(P3_DATAO_REG_22__SCAN_IN), .Z(n15609)
         );
  AOI211_X1 U16714 ( .C1(n15612), .C2(n15611), .A(n15610), .B(n15609), .ZN(
        n15615) );
  XOR2_X1 U16715 ( .A(keyinput_203), .B(P3_DATAO_REG_21__SCAN_IN), .Z(n15614)
         );
  XOR2_X1 U16716 ( .A(keyinput_204), .B(P3_DATAO_REG_20__SCAN_IN), .Z(n15613)
         );
  OAI21_X1 U16717 ( .B1(n15615), .B2(n15614), .A(n15613), .ZN(n15618) );
  XNOR2_X1 U16718 ( .A(keyinput_205), .B(P3_DATAO_REG_19__SCAN_IN), .ZN(n15617) );
  XNOR2_X1 U16719 ( .A(keyinput_206), .B(P3_DATAO_REG_18__SCAN_IN), .ZN(n15616) );
  NAND3_X1 U16720 ( .A1(n15618), .A2(n15617), .A3(n15616), .ZN(n15622) );
  XOR2_X1 U16721 ( .A(keyinput_209), .B(P3_DATAO_REG_15__SCAN_IN), .Z(n15621)
         );
  XOR2_X1 U16722 ( .A(keyinput_207), .B(P3_DATAO_REG_17__SCAN_IN), .Z(n15620)
         );
  XNOR2_X1 U16723 ( .A(keyinput_208), .B(P3_DATAO_REG_16__SCAN_IN), .ZN(n15619) );
  NAND4_X1 U16724 ( .A1(n15622), .A2(n15621), .A3(n15620), .A4(n15619), .ZN(
        n15625) );
  XOR2_X1 U16725 ( .A(keyinput_211), .B(P3_DATAO_REG_13__SCAN_IN), .Z(n15624)
         );
  XNOR2_X1 U16726 ( .A(keyinput_210), .B(P3_DATAO_REG_14__SCAN_IN), .ZN(n15623) );
  NAND3_X1 U16727 ( .A1(n15625), .A2(n15624), .A3(n15623), .ZN(n15628) );
  XOR2_X1 U16728 ( .A(keyinput_213), .B(P3_DATAO_REG_11__SCAN_IN), .Z(n15627)
         );
  XNOR2_X1 U16729 ( .A(keyinput_212), .B(P3_DATAO_REG_12__SCAN_IN), .ZN(n15626) );
  NAND3_X1 U16730 ( .A1(n15628), .A2(n15627), .A3(n15626), .ZN(n15631) );
  XOR2_X1 U16731 ( .A(keyinput_214), .B(P3_DATAO_REG_10__SCAN_IN), .Z(n15630)
         );
  XOR2_X1 U16732 ( .A(keyinput_215), .B(P3_DATAO_REG_9__SCAN_IN), .Z(n15629)
         );
  NAND3_X1 U16733 ( .A1(n15631), .A2(n15630), .A3(n15629), .ZN(n15635) );
  XNOR2_X1 U16734 ( .A(keyinput_216), .B(P3_DATAO_REG_8__SCAN_IN), .ZN(n15634)
         );
  XNOR2_X1 U16735 ( .A(keyinput_217), .B(P3_DATAO_REG_7__SCAN_IN), .ZN(n15633)
         );
  XNOR2_X1 U16736 ( .A(keyinput_218), .B(P3_DATAO_REG_6__SCAN_IN), .ZN(n15632)
         );
  AOI211_X1 U16737 ( .C1(n15635), .C2(n15634), .A(n15633), .B(n15632), .ZN(
        n15638) );
  XOR2_X1 U16738 ( .A(keyinput_219), .B(P3_DATAO_REG_5__SCAN_IN), .Z(n15637)
         );
  XNOR2_X1 U16739 ( .A(keyinput_220), .B(P3_DATAO_REG_4__SCAN_IN), .ZN(n15636)
         );
  OAI21_X1 U16740 ( .B1(n15638), .B2(n15637), .A(n15636), .ZN(n15642) );
  XNOR2_X1 U16741 ( .A(keyinput_221), .B(P3_DATAO_REG_3__SCAN_IN), .ZN(n15641)
         );
  XOR2_X1 U16742 ( .A(keyinput_223), .B(P3_DATAO_REG_1__SCAN_IN), .Z(n15640)
         );
  XOR2_X1 U16743 ( .A(keyinput_222), .B(P3_DATAO_REG_2__SCAN_IN), .Z(n15639)
         );
  AOI211_X1 U16744 ( .C1(n15642), .C2(n15641), .A(n15640), .B(n15639), .ZN(
        n15646) );
  XNOR2_X1 U16745 ( .A(keyinput_225), .B(P3_ADDR_REG_0__SCAN_IN), .ZN(n15645)
         );
  XNOR2_X1 U16746 ( .A(keyinput_226), .B(P3_ADDR_REG_1__SCAN_IN), .ZN(n15644)
         );
  XNOR2_X1 U16747 ( .A(keyinput_224), .B(P3_DATAO_REG_0__SCAN_IN), .ZN(n15643)
         );
  NOR4_X1 U16748 ( .A1(n15646), .A2(n15645), .A3(n15644), .A4(n15643), .ZN(
        n15650) );
  XOR2_X1 U16749 ( .A(keyinput_227), .B(P3_ADDR_REG_2__SCAN_IN), .Z(n15649) );
  XOR2_X1 U16750 ( .A(keyinput_229), .B(P3_ADDR_REG_4__SCAN_IN), .Z(n15648) );
  XOR2_X1 U16751 ( .A(keyinput_228), .B(P3_ADDR_REG_3__SCAN_IN), .Z(n15647) );
  OAI211_X1 U16752 ( .C1(n15650), .C2(n15649), .A(n15648), .B(n15647), .ZN(
        n15658) );
  XOR2_X1 U16753 ( .A(keyinput_233), .B(P3_ADDR_REG_8__SCAN_IN), .Z(n15654) );
  XOR2_X1 U16754 ( .A(keyinput_232), .B(P3_ADDR_REG_7__SCAN_IN), .Z(n15653) );
  XOR2_X1 U16755 ( .A(keyinput_231), .B(P3_ADDR_REG_6__SCAN_IN), .Z(n15652) );
  XNOR2_X1 U16756 ( .A(keyinput_230), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n15651)
         );
  NOR4_X1 U16757 ( .A1(n15654), .A2(n15653), .A3(n15652), .A4(n15651), .ZN(
        n15657) );
  XOR2_X1 U16758 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_235), .Z(n15656) );
  XOR2_X1 U16759 ( .A(keyinput_234), .B(P3_ADDR_REG_9__SCAN_IN), .Z(n15655) );
  AOI211_X1 U16760 ( .C1(n15658), .C2(n15657), .A(n15656), .B(n15655), .ZN(
        n15662) );
  XNOR2_X1 U16761 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_236), .ZN(n15661) );
  XNOR2_X1 U16762 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_238), .ZN(n15660) );
  XNOR2_X1 U16763 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_237), .ZN(n15659) );
  OAI211_X1 U16764 ( .C1(n15662), .C2(n15661), .A(n15660), .B(n15659), .ZN(
        n15666) );
  XNOR2_X1 U16765 ( .A(n15867), .B(keyinput_240), .ZN(n15665) );
  XOR2_X1 U16766 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_239), .Z(n15664) );
  XNOR2_X1 U16767 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_241), .ZN(n15663) );
  NAND4_X1 U16768 ( .A1(n15666), .A2(n15665), .A3(n15664), .A4(n15663), .ZN(
        n15668) );
  XNOR2_X1 U16769 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_242), .ZN(n15667) );
  NAND2_X1 U16770 ( .A1(n15668), .A2(n15667), .ZN(n15683) );
  INV_X1 U16771 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n15674) );
  INV_X1 U16772 ( .A(keyinput_249), .ZN(n15673) );
  AOI22_X1 U16773 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(keyinput_243), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput_245), .ZN(n15672) );
  OAI22_X1 U16774 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput_244), .B1(
        P1_IR_REG_14__SCAN_IN), .B2(keyinput_249), .ZN(n15670) );
  OAI22_X1 U16775 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput_245), .B1(
        P1_IR_REG_8__SCAN_IN), .B2(keyinput_243), .ZN(n15669) );
  AOI211_X1 U16776 ( .C1(keyinput_244), .C2(P1_IR_REG_9__SCAN_IN), .A(n15670), 
        .B(n15669), .ZN(n15671) );
  OAI211_X1 U16777 ( .C1(n15674), .C2(n15673), .A(n15672), .B(n15671), .ZN(
        n15679) );
  XOR2_X1 U16778 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_246), .Z(n15678) );
  XNOR2_X1 U16779 ( .A(n15675), .B(keyinput_248), .ZN(n15677) );
  XNOR2_X1 U16780 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_247), .ZN(n15676)
         );
  NOR4_X1 U16781 ( .A1(n15679), .A2(n15678), .A3(n15677), .A4(n15676), .ZN(
        n15682) );
  XOR2_X1 U16782 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_251), .Z(n15681) );
  XNOR2_X1 U16783 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_250), .ZN(n15680)
         );
  AOI211_X1 U16784 ( .C1(n15683), .C2(n15682), .A(n15681), .B(n15680), .ZN(
        n15687) );
  XNOR2_X1 U16785 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_252), .ZN(n15686)
         );
  XNOR2_X1 U16786 ( .A(n15684), .B(keyinput_253), .ZN(n15685) );
  OAI21_X1 U16787 ( .B1(n15687), .B2(n15686), .A(n15685), .ZN(n15691) );
  XNOR2_X1 U16788 ( .A(n15688), .B(keyinput_255), .ZN(n15690) );
  XNOR2_X1 U16789 ( .A(n15692), .B(keyinput_254), .ZN(n15689) );
  NAND3_X1 U16790 ( .A1(n15691), .A2(n15690), .A3(n15689), .ZN(n15895) );
  XNOR2_X1 U16791 ( .A(n15692), .B(keyinput_126), .ZN(n15894) );
  XOR2_X1 U16792 ( .A(P3_WR_REG_SCAN_IN), .B(keyinput_0), .Z(n15695) );
  XOR2_X1 U16793 ( .A(SI_31_), .B(keyinput_1), .Z(n15694) );
  XOR2_X1 U16794 ( .A(SI_30_), .B(keyinput_2), .Z(n15693) );
  AOI21_X1 U16795 ( .B1(n15695), .B2(n15694), .A(n15693), .ZN(n15699) );
  XNOR2_X1 U16796 ( .A(n15696), .B(keyinput_3), .ZN(n15698) );
  XNOR2_X1 U16797 ( .A(SI_28_), .B(keyinput_4), .ZN(n15697) );
  OAI21_X1 U16798 ( .B1(n15699), .B2(n15698), .A(n15697), .ZN(n15703) );
  XNOR2_X1 U16799 ( .A(n15700), .B(keyinput_5), .ZN(n15702) );
  XNOR2_X1 U16800 ( .A(SI_26_), .B(keyinput_6), .ZN(n15701) );
  NAND3_X1 U16801 ( .A1(n15703), .A2(n15702), .A3(n15701), .ZN(n15708) );
  XNOR2_X1 U16802 ( .A(n15704), .B(keyinput_7), .ZN(n15707) );
  XNOR2_X1 U16803 ( .A(n15705), .B(keyinput_8), .ZN(n15706) );
  NAND3_X1 U16804 ( .A1(n15708), .A2(n15707), .A3(n15706), .ZN(n15711) );
  XOR2_X1 U16805 ( .A(SI_22_), .B(keyinput_10), .Z(n15710) );
  XOR2_X1 U16806 ( .A(SI_23_), .B(keyinput_9), .Z(n15709) );
  NAND3_X1 U16807 ( .A1(n15711), .A2(n15710), .A3(n15709), .ZN(n15715) );
  XNOR2_X1 U16808 ( .A(SI_19_), .B(keyinput_13), .ZN(n15714) );
  XNOR2_X1 U16809 ( .A(SI_20_), .B(keyinput_12), .ZN(n15713) );
  XNOR2_X1 U16810 ( .A(SI_21_), .B(keyinput_11), .ZN(n15712) );
  NAND4_X1 U16811 ( .A1(n15715), .A2(n15714), .A3(n15713), .A4(n15712), .ZN(
        n15720) );
  XNOR2_X1 U16812 ( .A(n15716), .B(keyinput_14), .ZN(n15719) );
  XNOR2_X1 U16813 ( .A(n15717), .B(keyinput_15), .ZN(n15718) );
  AOI21_X1 U16814 ( .B1(n15720), .B2(n15719), .A(n15718), .ZN(n15723) );
  XNOR2_X1 U16815 ( .A(SI_16_), .B(keyinput_16), .ZN(n15722) );
  XNOR2_X1 U16816 ( .A(SI_15_), .B(keyinput_17), .ZN(n15721) );
  OAI21_X1 U16817 ( .B1(n15723), .B2(n15722), .A(n15721), .ZN(n15727) );
  XNOR2_X1 U16818 ( .A(SI_14_), .B(keyinput_18), .ZN(n15726) );
  XNOR2_X1 U16819 ( .A(n15724), .B(keyinput_19), .ZN(n15725) );
  AOI21_X1 U16820 ( .B1(n15727), .B2(n15726), .A(n15725), .ZN(n15731) );
  XNOR2_X1 U16821 ( .A(n15728), .B(keyinput_20), .ZN(n15730) );
  XNOR2_X1 U16822 ( .A(SI_11_), .B(keyinput_21), .ZN(n15729) );
  OAI21_X1 U16823 ( .B1(n15731), .B2(n15730), .A(n15729), .ZN(n15734) );
  XOR2_X1 U16824 ( .A(SI_10_), .B(keyinput_22), .Z(n15733) );
  XOR2_X1 U16825 ( .A(SI_9_), .B(keyinput_23), .Z(n15732) );
  NAND3_X1 U16826 ( .A1(n15734), .A2(n15733), .A3(n15732), .ZN(n15737) );
  XOR2_X1 U16827 ( .A(SI_8_), .B(keyinput_24), .Z(n15736) );
  XNOR2_X1 U16828 ( .A(SI_7_), .B(keyinput_25), .ZN(n15735) );
  AOI21_X1 U16829 ( .B1(n15737), .B2(n15736), .A(n15735), .ZN(n15740) );
  XOR2_X1 U16830 ( .A(SI_6_), .B(keyinput_26), .Z(n15739) );
  XNOR2_X1 U16831 ( .A(SI_5_), .B(keyinput_27), .ZN(n15738) );
  OAI21_X1 U16832 ( .B1(n15740), .B2(n15739), .A(n15738), .ZN(n15743) );
  XOR2_X1 U16833 ( .A(SI_3_), .B(keyinput_29), .Z(n15742) );
  XNOR2_X1 U16834 ( .A(SI_4_), .B(keyinput_28), .ZN(n15741) );
  NAND3_X1 U16835 ( .A1(n15743), .A2(n15742), .A3(n15741), .ZN(n15749) );
  XNOR2_X1 U16836 ( .A(SI_2_), .B(keyinput_30), .ZN(n15748) );
  XOR2_X1 U16837 ( .A(P3_RD_REG_SCAN_IN), .B(keyinput_33), .Z(n15746) );
  XNOR2_X1 U16838 ( .A(SI_0_), .B(keyinput_32), .ZN(n15745) );
  XNOR2_X1 U16839 ( .A(SI_1_), .B(keyinput_31), .ZN(n15744) );
  NAND3_X1 U16840 ( .A1(n15746), .A2(n15745), .A3(n15744), .ZN(n15747) );
  AOI21_X1 U16841 ( .B1(n15749), .B2(n15748), .A(n15747), .ZN(n15752) );
  XNOR2_X1 U16842 ( .A(P3_U3151), .B(keyinput_34), .ZN(n15751) );
  XNOR2_X1 U16843 ( .A(P3_REG3_REG_7__SCAN_IN), .B(keyinput_35), .ZN(n15750)
         );
  NOR3_X1 U16844 ( .A1(n15752), .A2(n15751), .A3(n15750), .ZN(n15755) );
  XOR2_X1 U16845 ( .A(P3_REG3_REG_27__SCAN_IN), .B(keyinput_36), .Z(n15754) );
  XNOR2_X1 U16846 ( .A(P3_REG3_REG_14__SCAN_IN), .B(keyinput_37), .ZN(n15753)
         );
  NOR3_X1 U16847 ( .A1(n15755), .A2(n15754), .A3(n15753), .ZN(n15760) );
  XNOR2_X1 U16848 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput_38), .ZN(n15759)
         );
  XNOR2_X1 U16849 ( .A(n15756), .B(keyinput_40), .ZN(n15758) );
  XNOR2_X1 U16850 ( .A(P3_REG3_REG_10__SCAN_IN), .B(keyinput_39), .ZN(n15757)
         );
  OAI211_X1 U16851 ( .C1(n15760), .C2(n15759), .A(n15758), .B(n15757), .ZN(
        n15769) );
  XNOR2_X1 U16852 ( .A(P3_REG3_REG_19__SCAN_IN), .B(keyinput_41), .ZN(n15768)
         );
  XOR2_X1 U16853 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_44), .Z(n15766) );
  XNOR2_X1 U16854 ( .A(n15761), .B(keyinput_45), .ZN(n15765) );
  XNOR2_X1 U16855 ( .A(n15762), .B(keyinput_42), .ZN(n15764) );
  XNOR2_X1 U16856 ( .A(P3_REG3_REG_8__SCAN_IN), .B(keyinput_43), .ZN(n15763)
         );
  NAND4_X1 U16857 ( .A1(n15766), .A2(n15765), .A3(n15764), .A4(n15763), .ZN(
        n15767) );
  AOI21_X1 U16858 ( .B1(n15769), .B2(n15768), .A(n15767), .ZN(n15772) );
  XNOR2_X1 U16859 ( .A(P3_REG3_REG_12__SCAN_IN), .B(keyinput_46), .ZN(n15771)
         );
  XNOR2_X1 U16860 ( .A(P3_REG3_REG_25__SCAN_IN), .B(keyinput_47), .ZN(n15770)
         );
  OAI21_X1 U16861 ( .B1(n15772), .B2(n15771), .A(n15770), .ZN(n15777) );
  XNOR2_X1 U16862 ( .A(n15773), .B(keyinput_48), .ZN(n15776) );
  XNOR2_X1 U16863 ( .A(n15774), .B(keyinput_49), .ZN(n15775) );
  AOI21_X1 U16864 ( .B1(n15777), .B2(n15776), .A(n15775), .ZN(n15781) );
  XNOR2_X1 U16865 ( .A(P3_REG3_REG_17__SCAN_IN), .B(keyinput_50), .ZN(n15780)
         );
  XNOR2_X1 U16866 ( .A(P3_REG3_REG_24__SCAN_IN), .B(keyinput_51), .ZN(n15779)
         );
  XNOR2_X1 U16867 ( .A(P3_REG3_REG_4__SCAN_IN), .B(keyinput_52), .ZN(n15778)
         );
  OAI211_X1 U16868 ( .C1(n15781), .C2(n15780), .A(n15779), .B(n15778), .ZN(
        n15785) );
  XNOR2_X1 U16869 ( .A(n15782), .B(keyinput_53), .ZN(n15784) );
  XOR2_X1 U16870 ( .A(P3_REG3_REG_0__SCAN_IN), .B(keyinput_54), .Z(n15783) );
  NAND3_X1 U16871 ( .A1(n15785), .A2(n15784), .A3(n15783), .ZN(n15792) );
  OAI22_X1 U16872 ( .A1(n8771), .A2(keyinput_56), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(keyinput_57), .ZN(n15786) );
  AOI221_X1 U16873 ( .B1(n8771), .B2(keyinput_56), .C1(keyinput_57), .C2(
        P3_REG3_REG_22__SCAN_IN), .A(n15786), .ZN(n15791) );
  XOR2_X1 U16874 ( .A(P3_REG3_REG_11__SCAN_IN), .B(keyinput_58), .Z(n15790) );
  OAI22_X1 U16875 ( .A1(n15788), .A2(keyinput_55), .B1(keyinput_59), .B2(
        P3_REG3_REG_2__SCAN_IN), .ZN(n15787) );
  AOI221_X1 U16876 ( .B1(n15788), .B2(keyinput_55), .C1(P3_REG3_REG_2__SCAN_IN), .C2(keyinput_59), .A(n15787), .ZN(n15789) );
  NAND4_X1 U16877 ( .A1(n15792), .A2(n15791), .A3(n15790), .A4(n15789), .ZN(
        n15799) );
  XOR2_X1 U16878 ( .A(P3_REG3_REG_18__SCAN_IN), .B(keyinput_60), .Z(n15794) );
  XNOR2_X1 U16879 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput_61), .ZN(n15793)
         );
  NOR2_X1 U16880 ( .A1(n15794), .A2(n15793), .ZN(n15798) );
  XOR2_X1 U16881 ( .A(P3_REG3_REG_15__SCAN_IN), .B(keyinput_63), .Z(n15797) );
  XNOR2_X1 U16882 ( .A(n15795), .B(keyinput_62), .ZN(n15796) );
  AOI211_X1 U16883 ( .C1(n15799), .C2(n15798), .A(n15797), .B(n15796), .ZN(
        n15802) );
  XOR2_X1 U16884 ( .A(P3_B_REG_SCAN_IN), .B(keyinput_64), .Z(n15801) );
  XOR2_X1 U16885 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .Z(n15800)
         );
  OAI21_X1 U16886 ( .B1(n15802), .B2(n15801), .A(n15800), .ZN(n15808) );
  XNOR2_X1 U16887 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(keyinput_66), .ZN(n15807)
         );
  XOR2_X1 U16888 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .Z(n15805)
         );
  XNOR2_X1 U16889 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(keyinput_69), .ZN(n15804)
         );
  XNOR2_X1 U16890 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .ZN(n15803)
         );
  NAND3_X1 U16891 ( .A1(n15805), .A2(n15804), .A3(n15803), .ZN(n15806) );
  AOI21_X1 U16892 ( .B1(n15808), .B2(n15807), .A(n15806), .ZN(n15811) );
  XNOR2_X1 U16893 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(keyinput_70), .ZN(n15810)
         );
  XOR2_X1 U16894 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .Z(n15809)
         );
  OAI21_X1 U16895 ( .B1(n15811), .B2(n15810), .A(n15809), .ZN(n15815) );
  XOR2_X1 U16896 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .Z(n15814)
         );
  XOR2_X1 U16897 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .Z(n15813)
         );
  XOR2_X1 U16898 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .Z(n15812)
         );
  AOI211_X1 U16899 ( .C1(n15815), .C2(n15814), .A(n15813), .B(n15812), .ZN(
        n15818) );
  XOR2_X1 U16900 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .Z(n15817)
         );
  XNOR2_X1 U16901 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(keyinput_76), .ZN(n15816)
         );
  OAI21_X1 U16902 ( .B1(n15818), .B2(n15817), .A(n15816), .ZN(n15821) );
  XNOR2_X1 U16903 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .ZN(n15820)
         );
  XNOR2_X1 U16904 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .ZN(n15819)
         );
  NAND3_X1 U16905 ( .A1(n15821), .A2(n15820), .A3(n15819), .ZN(n15825) );
  XNOR2_X1 U16906 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .ZN(n15824)
         );
  XNOR2_X1 U16907 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .ZN(n15823)
         );
  XNOR2_X1 U16908 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(keyinput_80), .ZN(n15822)
         );
  NAND4_X1 U16909 ( .A1(n15825), .A2(n15824), .A3(n15823), .A4(n15822), .ZN(
        n15828) );
  XOR2_X1 U16910 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(keyinput_82), .Z(n15827)
         );
  XOR2_X1 U16911 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(keyinput_83), .Z(n15826)
         );
  NAND3_X1 U16912 ( .A1(n15828), .A2(n15827), .A3(n15826), .ZN(n15831) );
  XOR2_X1 U16913 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(keyinput_84), .Z(n15830)
         );
  XNOR2_X1 U16914 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .ZN(n15829)
         );
  NAND3_X1 U16915 ( .A1(n15831), .A2(n15830), .A3(n15829), .ZN(n15834) );
  XNOR2_X1 U16916 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(keyinput_87), .ZN(n15833)
         );
  XNOR2_X1 U16917 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(keyinput_86), .ZN(n15832)
         );
  NAND3_X1 U16918 ( .A1(n15834), .A2(n15833), .A3(n15832), .ZN(n15838) );
  XNOR2_X1 U16919 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .ZN(n15837)
         );
  XNOR2_X1 U16920 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(keyinput_90), .ZN(n15836)
         );
  XNOR2_X1 U16921 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .ZN(n15835)
         );
  AOI211_X1 U16922 ( .C1(n15838), .C2(n15837), .A(n15836), .B(n15835), .ZN(
        n15841) );
  XNOR2_X1 U16923 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(keyinput_91), .ZN(n15840)
         );
  XNOR2_X1 U16924 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(keyinput_92), .ZN(n15839)
         );
  OAI21_X1 U16925 ( .B1(n15841), .B2(n15840), .A(n15839), .ZN(n15845) );
  XNOR2_X1 U16926 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(keyinput_93), .ZN(n15844)
         );
  XOR2_X1 U16927 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(keyinput_94), .Z(n15843) );
  XNOR2_X1 U16928 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(keyinput_95), .ZN(n15842)
         );
  AOI211_X1 U16929 ( .C1(n15845), .C2(n15844), .A(n15843), .B(n15842), .ZN(
        n15849) );
  XOR2_X1 U16930 ( .A(P3_ADDR_REG_0__SCAN_IN), .B(keyinput_97), .Z(n15848) );
  XNOR2_X1 U16931 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(keyinput_98), .ZN(n15847)
         );
  XNOR2_X1 U16932 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(keyinput_96), .ZN(n15846)
         );
  NOR4_X1 U16933 ( .A1(n15849), .A2(n15848), .A3(n15847), .A4(n15846), .ZN(
        n15853) );
  XNOR2_X1 U16934 ( .A(P3_ADDR_REG_2__SCAN_IN), .B(keyinput_99), .ZN(n15852)
         );
  XOR2_X1 U16935 ( .A(P3_ADDR_REG_3__SCAN_IN), .B(keyinput_100), .Z(n15851) );
  XNOR2_X1 U16936 ( .A(P3_ADDR_REG_4__SCAN_IN), .B(keyinput_101), .ZN(n15850)
         );
  OAI211_X1 U16937 ( .C1(n15853), .C2(n15852), .A(n15851), .B(n15850), .ZN(
        n15861) );
  XOR2_X1 U16938 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(keyinput_104), .Z(n15857) );
  XOR2_X1 U16939 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(keyinput_102), .Z(n15856) );
  XOR2_X1 U16940 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(keyinput_105), .Z(n15855) );
  XNOR2_X1 U16941 ( .A(P3_ADDR_REG_6__SCAN_IN), .B(keyinput_103), .ZN(n15854)
         );
  NOR4_X1 U16942 ( .A1(n15857), .A2(n15856), .A3(n15855), .A4(n15854), .ZN(
        n15860) );
  XOR2_X1 U16943 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(keyinput_106), .Z(n15859) );
  XOR2_X1 U16944 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_107), .Z(n15858) );
  AOI211_X1 U16945 ( .C1(n15861), .C2(n15860), .A(n15859), .B(n15858), .ZN(
        n15866) );
  XNOR2_X1 U16946 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_108), .ZN(n15865) );
  XOR2_X1 U16947 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_110), .Z(n15864) );
  XNOR2_X1 U16948 ( .A(n15862), .B(keyinput_109), .ZN(n15863) );
  OAI211_X1 U16949 ( .C1(n15866), .C2(n15865), .A(n15864), .B(n15863), .ZN(
        n15872) );
  XNOR2_X1 U16950 ( .A(n15867), .B(keyinput_112), .ZN(n15871) );
  XNOR2_X1 U16951 ( .A(n15868), .B(keyinput_113), .ZN(n15870) );
  XOR2_X1 U16952 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_111), .Z(n15869) );
  NAND4_X1 U16953 ( .A1(n15872), .A2(n15871), .A3(n15870), .A4(n15869), .ZN(
        n15884) );
  XOR2_X1 U16954 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_114), .Z(n15883) );
  OAI22_X1 U16955 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput_116), .B1(
        keyinput_121), .B2(P1_IR_REG_14__SCAN_IN), .ZN(n15873) );
  AOI221_X1 U16956 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput_116), .C1(
        P1_IR_REG_14__SCAN_IN), .C2(keyinput_121), .A(n15873), .ZN(n15881) );
  XOR2_X1 U16957 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_118), .Z(n15877) );
  XNOR2_X1 U16958 ( .A(n15874), .B(keyinput_115), .ZN(n15876) );
  XNOR2_X1 U16959 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_119), .ZN(n15875)
         );
  NOR3_X1 U16960 ( .A1(n15877), .A2(n15876), .A3(n15875), .ZN(n15880) );
  XNOR2_X1 U16961 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_120), .ZN(n15879)
         );
  XNOR2_X1 U16962 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_117), .ZN(n15878)
         );
  NAND4_X1 U16963 ( .A1(n15881), .A2(n15880), .A3(n15879), .A4(n15878), .ZN(
        n15882) );
  AOI21_X1 U16964 ( .B1(n15884), .B2(n15883), .A(n15882), .ZN(n15888) );
  XNOR2_X1 U16965 ( .A(n15885), .B(keyinput_122), .ZN(n15887) );
  XNOR2_X1 U16966 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_123), .ZN(n15886)
         );
  NOR3_X1 U16967 ( .A1(n15888), .A2(n15887), .A3(n15886), .ZN(n15891) );
  XNOR2_X1 U16968 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_124), .ZN(n15890)
         );
  XNOR2_X1 U16969 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_125), .ZN(n15889)
         );
  OAI21_X1 U16970 ( .B1(n15891), .B2(n15890), .A(n15889), .ZN(n15893) );
  XNOR2_X1 U16971 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_127), .ZN(n15892)
         );
  NAND4_X1 U16972 ( .A1(n15895), .A2(n15894), .A3(n15893), .A4(n15892), .ZN(
        n15898) );
  MUX2_X1 U16973 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15896), .S(n16556), .Z(
        n15897) );
  XNOR2_X1 U16974 ( .A(n15898), .B(n15897), .ZN(P1_U3504) );
  MUX2_X1 U16975 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15899), .S(n16556), .Z(
        P1_U3501) );
  MUX2_X1 U16976 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n15900), .S(n16556), .Z(
        P1_U3498) );
  MUX2_X1 U16977 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n15901), .S(n16556), .Z(
        P1_U3495) );
  NOR4_X1 U16978 ( .A1(n15902), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n9361), .ZN(n15903) );
  AOI21_X1 U16979 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n15904), .A(n15903), 
        .ZN(n15905) );
  OAI21_X1 U16980 ( .B1(n15906), .B2(n15919), .A(n15905), .ZN(P1_U3324) );
  OAI222_X1 U16981 ( .A1(P1_U3086), .A2(n15909), .B1(n15919), .B2(n15908), 
        .C1(n15907), .C2(n15916), .ZN(P1_U3326) );
  OAI222_X1 U16982 ( .A1(n15912), .A2(P1_U3086), .B1(n15919), .B2(n15911), 
        .C1(n15910), .C2(n15916), .ZN(P1_U3328) );
  OAI222_X1 U16983 ( .A1(n15915), .A2(P1_U3086), .B1(n15919), .B2(n15914), 
        .C1(n15913), .C2(n15916), .ZN(P1_U3329) );
  OAI222_X1 U16984 ( .A1(P1_U3086), .A2(n15920), .B1(n15919), .B2(n15918), 
        .C1(n15917), .C2(n15916), .ZN(P1_U3330) );
  MUX2_X1 U16985 ( .A(n15921), .B(n9838), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U16986 ( .A(n15922), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16987 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n15954) );
  INV_X1 U16988 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n15952) );
  INV_X1 U16989 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n15950) );
  XNOR2_X1 U16990 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(n15923), .ZN(n15972) );
  INV_X1 U16991 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n15948) );
  NOR2_X1 U16992 ( .A1(n16001), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n16000) );
  NOR2_X1 U16993 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n15977), .ZN(n15934) );
  NAND2_X1 U16994 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n15925), .ZN(n15927) );
  NAND2_X1 U16995 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n15928), .ZN(n15929) );
  NAND2_X1 U16996 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n15930), .ZN(n15933) );
  INV_X1 U16997 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n15931) );
  NAND2_X1 U16998 ( .A1(n15980), .A2(n16363), .ZN(n15932) );
  NAND2_X1 U16999 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n15977), .ZN(n15976) );
  INV_X1 U17000 ( .A(n16003), .ZN(n15935) );
  NAND2_X1 U17001 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n15946), .ZN(n15944) );
  OAI21_X1 U17002 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n15946), .A(n15944), .ZN(
        n15973) );
  XOR2_X1 U17003 ( .A(n15948), .B(P1_ADDR_REG_10__SCAN_IN), .Z(n16011) );
  NAND2_X1 U17004 ( .A1(n16012), .A2(n16011), .ZN(n15947) );
  AOI21_X2 U17005 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n15950), .A(n15949), 
        .ZN(n16015) );
  XOR2_X1 U17006 ( .A(n15952), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n16014) );
  NAND2_X1 U17007 ( .A1(n16015), .A2(n16014), .ZN(n15951) );
  INV_X1 U17008 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15968) );
  NAND2_X1 U17009 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n15968), .ZN(n15953) );
  XNOR2_X1 U17010 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n15956), .ZN(n16018) );
  NOR2_X1 U17011 ( .A1(n16019), .A2(n16018), .ZN(n15955) );
  AOI21_X1 U17012 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n15956), .A(n15955), 
        .ZN(n16022) );
  XOR2_X1 U17013 ( .A(P3_ADDR_REG_15__SCAN_IN), .B(n15958), .Z(n16021) );
  NAND2_X1 U17014 ( .A1(n16022), .A2(n16021), .ZN(n15957) );
  NOR2_X1 U17015 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n15959), .ZN(n15961) );
  XOR2_X1 U17016 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n15959), .Z(n16025) );
  NOR2_X1 U17017 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n15962), .ZN(n15964) );
  XOR2_X1 U17018 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n15962), .Z(n15966) );
  AND2_X1 U17019 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n15966), .ZN(n15963) );
  NAND2_X1 U17020 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n16038), .ZN(n15965) );
  OAI21_X1 U17021 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n16038), .A(n15965), 
        .ZN(n16036) );
  XOR2_X1 U17022 ( .A(n16035), .B(n16036), .Z(n16031) );
  XOR2_X1 U17023 ( .A(n15967), .B(n15966), .Z(n16029) );
  NAND2_X1 U17024 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n16029), .ZN(n16030) );
  INV_X1 U17025 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n16024) );
  INV_X1 U17026 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n16198) );
  XOR2_X1 U17027 ( .A(n15968), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n15970) );
  XNOR2_X1 U17028 ( .A(n15970), .B(n15969), .ZN(n16303) );
  INV_X1 U17029 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n16184) );
  XOR2_X1 U17030 ( .A(n15972), .B(n15971), .Z(n16299) );
  INV_X1 U17031 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n16255) );
  XOR2_X1 U17032 ( .A(n15974), .B(n15973), .Z(n16289) );
  XOR2_X1 U17033 ( .A(n15005), .B(n15975), .Z(n16008) );
  INV_X1 U17034 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n16159) );
  OAI21_X1 U17035 ( .B1(n15977), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n15976), .ZN(
        n15979) );
  XOR2_X1 U17036 ( .A(n15979), .B(n15978), .Z(n15998) );
  NAND2_X1 U17037 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n15981), .ZN(n15997) );
  INV_X1 U17038 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n15990) );
  NAND2_X1 U17039 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n15983), .ZN(n15987) );
  AOI21_X1 U17040 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n15985), .A(n15984), .ZN(
        n16272) );
  NOR2_X1 U17041 ( .A1(n16272), .A2(n10284), .ZN(n16325) );
  NAND2_X1 U17042 ( .A1(n16326), .A2(n16325), .ZN(n15986) );
  NAND2_X1 U17043 ( .A1(n15987), .A2(n15986), .ZN(n16274) );
  XNOR2_X1 U17044 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n15988), .ZN(n16275) );
  NAND2_X1 U17045 ( .A1(n16274), .A2(n16275), .ZN(n15989) );
  NOR2_X1 U17046 ( .A1(n16274), .A2(n16275), .ZN(n16273) );
  XNOR2_X1 U17047 ( .A(n15992), .B(n15991), .ZN(n15994) );
  NOR2_X1 U17048 ( .A1(n15993), .A2(n15994), .ZN(n15996) );
  XNOR2_X1 U17049 ( .A(n15994), .B(n15993), .ZN(n16277) );
  NOR2_X1 U17050 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(n16277), .ZN(n15995) );
  NOR2_X1 U17051 ( .A1(n15996), .A2(n15995), .ZN(n16279) );
  NOR2_X1 U17052 ( .A1(n15998), .A2(n15999), .ZN(n16281) );
  AOI21_X1 U17053 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n16001), .A(n16000), .ZN(
        n16002) );
  XOR2_X1 U17054 ( .A(n16003), .B(n16002), .Z(n16322) );
  NAND2_X1 U17055 ( .A1(n16323), .A2(n16322), .ZN(n16004) );
  XNOR2_X1 U17056 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n16006), .ZN(n16284) );
  NOR2_X1 U17057 ( .A1(n16008), .A2(n16007), .ZN(n16010) );
  XNOR2_X1 U17058 ( .A(n16012), .B(n16011), .ZN(n16294) );
  INV_X1 U17059 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n16295) );
  NAND2_X1 U17060 ( .A1(n16299), .A2(n16298), .ZN(n16013) );
  XNOR2_X1 U17061 ( .A(n16015), .B(n16014), .ZN(n16017) );
  XNOR2_X1 U17062 ( .A(n16019), .B(n16018), .ZN(n16307) );
  NAND2_X1 U17063 ( .A1(n16308), .A2(n16307), .ZN(n16020) );
  NOR2_X1 U17064 ( .A1(n16308), .A2(n16307), .ZN(n16306) );
  XOR2_X1 U17065 ( .A(n16022), .B(n16021), .Z(n16312) );
  NAND2_X1 U17066 ( .A1(n16311), .A2(n16312), .ZN(n16023) );
  XOR2_X1 U17067 ( .A(n16026), .B(n16025), .Z(n16028) );
  XOR2_X1 U17068 ( .A(n16029), .B(P2_ADDR_REG_17__SCAN_IN), .Z(n16318) );
  NAND2_X1 U17069 ( .A1(n16031), .A2(n16032), .ZN(n16034) );
  NAND2_X1 U17070 ( .A1(n16320), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n16033) );
  NOR2_X1 U17071 ( .A1(n16036), .A2(n16035), .ZN(n16037) );
  AOI21_X1 U17072 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n16038), .A(n16037), 
        .ZN(n16041) );
  XNOR2_X1 U17073 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n16039) );
  XNOR2_X1 U17074 ( .A(n16039), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n16040) );
  XNOR2_X1 U17075 ( .A(n16041), .B(n16040), .ZN(n16042) );
  INV_X1 U17076 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n16043) );
  NOR2_X1 U17077 ( .A1(n16073), .A2(n16043), .ZN(P1_U3323) );
  INV_X1 U17078 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n16044) );
  NOR2_X1 U17079 ( .A1(n16073), .A2(n16044), .ZN(P1_U3322) );
  INV_X1 U17080 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n16045) );
  NOR2_X1 U17081 ( .A1(n16073), .A2(n16045), .ZN(P1_U3321) );
  INV_X1 U17082 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n16046) );
  NOR2_X1 U17083 ( .A1(n16073), .A2(n16046), .ZN(P1_U3320) );
  INV_X1 U17084 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n16047) );
  NOR2_X1 U17085 ( .A1(n16073), .A2(n16047), .ZN(P1_U3319) );
  INV_X1 U17086 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n16048) );
  NOR2_X1 U17087 ( .A1(n16073), .A2(n16048), .ZN(P1_U3318) );
  INV_X1 U17088 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n16049) );
  NOR2_X1 U17089 ( .A1(n16073), .A2(n16049), .ZN(P1_U3317) );
  INV_X1 U17090 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n16050) );
  NOR2_X1 U17091 ( .A1(n16073), .A2(n16050), .ZN(P1_U3316) );
  INV_X1 U17092 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n16051) );
  NOR2_X1 U17093 ( .A1(n16073), .A2(n16051), .ZN(P1_U3315) );
  INV_X1 U17094 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n16052) );
  NOR2_X1 U17095 ( .A1(n16073), .A2(n16052), .ZN(P1_U3314) );
  INV_X1 U17096 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n16053) );
  NOR2_X1 U17097 ( .A1(n16073), .A2(n16053), .ZN(P1_U3313) );
  INV_X1 U17098 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n16054) );
  NOR2_X1 U17099 ( .A1(n16073), .A2(n16054), .ZN(P1_U3312) );
  INV_X1 U17100 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n16055) );
  NOR2_X1 U17101 ( .A1(n16073), .A2(n16055), .ZN(P1_U3311) );
  INV_X1 U17102 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n16056) );
  NOR2_X1 U17103 ( .A1(n16073), .A2(n16056), .ZN(P1_U3310) );
  INV_X1 U17104 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n16057) );
  NOR2_X1 U17105 ( .A1(n16073), .A2(n16057), .ZN(P1_U3309) );
  INV_X1 U17106 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n16058) );
  NOR2_X1 U17107 ( .A1(n16073), .A2(n16058), .ZN(P1_U3308) );
  INV_X1 U17108 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n16059) );
  NOR2_X1 U17109 ( .A1(n16073), .A2(n16059), .ZN(P1_U3307) );
  INV_X1 U17110 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n16060) );
  NOR2_X1 U17111 ( .A1(n16073), .A2(n16060), .ZN(P1_U3306) );
  INV_X1 U17112 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n16061) );
  NOR2_X1 U17113 ( .A1(n16073), .A2(n16061), .ZN(P1_U3305) );
  INV_X1 U17114 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n16062) );
  NOR2_X1 U17115 ( .A1(n16073), .A2(n16062), .ZN(P1_U3304) );
  INV_X1 U17116 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n16063) );
  NOR2_X1 U17117 ( .A1(n16073), .A2(n16063), .ZN(P1_U3303) );
  INV_X1 U17118 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n16064) );
  NOR2_X1 U17119 ( .A1(n16073), .A2(n16064), .ZN(P1_U3302) );
  INV_X1 U17120 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n16065) );
  NOR2_X1 U17121 ( .A1(n16073), .A2(n16065), .ZN(P1_U3301) );
  INV_X1 U17122 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n16066) );
  NOR2_X1 U17123 ( .A1(n16073), .A2(n16066), .ZN(P1_U3300) );
  INV_X1 U17124 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n16067) );
  NOR2_X1 U17125 ( .A1(n16073), .A2(n16067), .ZN(P1_U3299) );
  INV_X1 U17126 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n16068) );
  NOR2_X1 U17127 ( .A1(n16073), .A2(n16068), .ZN(P1_U3298) );
  INV_X1 U17128 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n16069) );
  NOR2_X1 U17129 ( .A1(n16073), .A2(n16069), .ZN(P1_U3297) );
  INV_X1 U17130 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n16070) );
  NOR2_X1 U17131 ( .A1(n16073), .A2(n16070), .ZN(P1_U3296) );
  INV_X1 U17132 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n16071) );
  NOR2_X1 U17133 ( .A1(n16073), .A2(n16071), .ZN(P1_U3295) );
  INV_X1 U17134 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n16072) );
  NOR2_X1 U17135 ( .A1(n16073), .A2(n16072), .ZN(P1_U3294) );
  INV_X1 U17136 ( .A(n16074), .ZN(n16075) );
  AOI22_X1 U17137 ( .A1(n16078), .A2(n16082), .B1(n16077), .B2(n16080), .ZN(
        P2_U3417) );
  AND2_X1 U17138 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n16080), .ZN(P2_U3295) );
  AND2_X1 U17139 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n16080), .ZN(P2_U3294) );
  AND2_X1 U17140 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n16080), .ZN(P2_U3293) );
  AND2_X1 U17141 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n16080), .ZN(P2_U3292) );
  AND2_X1 U17142 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n16080), .ZN(P2_U3291) );
  AND2_X1 U17143 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n16080), .ZN(P2_U3290) );
  AND2_X1 U17144 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n16080), .ZN(P2_U3289) );
  AND2_X1 U17145 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n16080), .ZN(P2_U3288) );
  AND2_X1 U17146 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n16080), .ZN(P2_U3287) );
  AND2_X1 U17147 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n16080), .ZN(P2_U3286) );
  AND2_X1 U17148 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n16080), .ZN(P2_U3285) );
  AND2_X1 U17149 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n16080), .ZN(P2_U3284) );
  AND2_X1 U17150 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n16080), .ZN(P2_U3283) );
  AND2_X1 U17151 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n16080), .ZN(P2_U3282) );
  AND2_X1 U17152 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n16080), .ZN(P2_U3281) );
  AND2_X1 U17153 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n16080), .ZN(P2_U3280) );
  AND2_X1 U17154 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n16080), .ZN(P2_U3279) );
  AND2_X1 U17155 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n16080), .ZN(P2_U3278) );
  AND2_X1 U17156 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n16080), .ZN(P2_U3277) );
  AND2_X1 U17157 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n16080), .ZN(P2_U3276) );
  AND2_X1 U17158 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n16080), .ZN(P2_U3275) );
  AND2_X1 U17159 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n16080), .ZN(P2_U3274) );
  AND2_X1 U17160 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n16080), .ZN(P2_U3273) );
  AND2_X1 U17161 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n16080), .ZN(P2_U3272) );
  AND2_X1 U17162 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n16080), .ZN(P2_U3271) );
  AND2_X1 U17163 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n16080), .ZN(P2_U3270) );
  AND2_X1 U17164 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n16080), .ZN(P2_U3269) );
  AND2_X1 U17165 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n16080), .ZN(P2_U3268) );
  AND2_X1 U17166 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n16080), .ZN(P2_U3267) );
  AND2_X1 U17167 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n16080), .ZN(P2_U3266) );
  NOR2_X1 U17168 ( .A1(n16097), .A2(P2_U3947), .ZN(P2_U3087) );
  NOR2_X1 U17169 ( .A1(n16079), .A2(n16330), .ZN(P3_U3150) );
  AOI22_X1 U17170 ( .A1(n16083), .A2(n16082), .B1(n16081), .B2(n16080), .ZN(
        P2_U3416) );
  AOI22_X1 U17171 ( .A1(n16097), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n16096) );
  NAND2_X1 U17172 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n16088) );
  INV_X1 U17173 ( .A(n16084), .ZN(n16087) );
  INV_X1 U17174 ( .A(n16085), .ZN(n16086) );
  AOI211_X1 U17175 ( .C1(n16088), .C2(n16087), .A(n16086), .B(n16247), .ZN(
        n16093) );
  NAND2_X1 U17176 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n16091) );
  AOI211_X1 U17177 ( .C1(n16091), .C2(n16090), .A(n16089), .B(n16228), .ZN(
        n16092) );
  AOI211_X1 U17178 ( .C1(n16234), .C2(n16094), .A(n16093), .B(n16092), .ZN(
        n16095) );
  NAND2_X1 U17179 ( .A1(n16096), .A2(n16095), .ZN(P2_U3215) );
  AOI22_X1 U17180 ( .A1(n16097), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n16109) );
  OAI211_X1 U17181 ( .C1(n16100), .C2(n16099), .A(n16222), .B(n16098), .ZN(
        n16101) );
  INV_X1 U17182 ( .A(n16101), .ZN(n16106) );
  AOI211_X1 U17183 ( .C1(n16104), .C2(n16103), .A(n16102), .B(n16228), .ZN(
        n16105) );
  AOI211_X1 U17184 ( .C1(n16234), .C2(n16107), .A(n16106), .B(n16105), .ZN(
        n16108) );
  NAND2_X1 U17185 ( .A1(n16109), .A2(n16108), .ZN(P2_U3216) );
  INV_X1 U17186 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n16278) );
  AOI211_X1 U17187 ( .C1(n16112), .C2(n16111), .A(n16110), .B(n16228), .ZN(
        n16119) );
  OAI211_X1 U17188 ( .C1(n16115), .C2(n16114), .A(n16222), .B(n16113), .ZN(
        n16116) );
  OAI21_X1 U17189 ( .B1(n16189), .B2(n16117), .A(n16116), .ZN(n16118) );
  NOR2_X1 U17190 ( .A1(n16119), .A2(n16118), .ZN(n16121) );
  NAND2_X1 U17191 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n16120) );
  OAI211_X1 U17192 ( .C1(n16254), .C2(n16278), .A(n16121), .B(n16120), .ZN(
        P2_U3217) );
  AOI211_X1 U17193 ( .C1(n16124), .C2(n16123), .A(n16228), .B(n16122), .ZN(
        n16131) );
  OAI211_X1 U17194 ( .C1(n16127), .C2(n16126), .A(n16222), .B(n16125), .ZN(
        n16128) );
  OAI21_X1 U17195 ( .B1(n16189), .B2(n16129), .A(n16128), .ZN(n16130) );
  NOR2_X1 U17196 ( .A1(n16131), .A2(n16130), .ZN(n16133) );
  NAND2_X1 U17197 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n16132) );
  OAI211_X1 U17198 ( .C1(n16254), .C2(n7979), .A(n16133), .B(n16132), .ZN(
        P2_U3218) );
  INV_X1 U17199 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n16146) );
  AOI211_X1 U17200 ( .C1(n16136), .C2(n16135), .A(n16228), .B(n16134), .ZN(
        n16143) );
  OAI211_X1 U17201 ( .C1(n16139), .C2(n16138), .A(n16222), .B(n16137), .ZN(
        n16140) );
  OAI21_X1 U17202 ( .B1(n16189), .B2(n16141), .A(n16140), .ZN(n16142) );
  NOR2_X1 U17203 ( .A1(n16143), .A2(n16142), .ZN(n16145) );
  OAI211_X1 U17204 ( .C1(n16254), .C2(n16146), .A(n16145), .B(n16144), .ZN(
        P2_U3219) );
  OAI211_X1 U17205 ( .C1(n16149), .C2(n16148), .A(n16222), .B(n16147), .ZN(
        n16150) );
  INV_X1 U17206 ( .A(n16150), .ZN(n16155) );
  AOI211_X1 U17207 ( .C1(n16153), .C2(n16152), .A(n16228), .B(n16151), .ZN(
        n16154) );
  AOI211_X1 U17208 ( .C1(n16234), .C2(n16156), .A(n16155), .B(n16154), .ZN(
        n16158) );
  NAND2_X1 U17209 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n16157) );
  OAI211_X1 U17210 ( .C1(n16254), .C2(n16159), .A(n16158), .B(n16157), .ZN(
        P2_U3220) );
  INV_X1 U17211 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n16287) );
  OAI211_X1 U17212 ( .C1(n16162), .C2(n16161), .A(n16222), .B(n16160), .ZN(
        n16163) );
  INV_X1 U17213 ( .A(n16163), .ZN(n16168) );
  AOI211_X1 U17214 ( .C1(n16166), .C2(n16165), .A(n16228), .B(n16164), .ZN(
        n16167) );
  AOI211_X1 U17215 ( .C1(n16234), .C2(n16169), .A(n16168), .B(n16167), .ZN(
        n16171) );
  NAND2_X1 U17216 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n16170) );
  OAI211_X1 U17217 ( .C1(n16287), .C2(n16254), .A(n16171), .B(n16170), .ZN(
        P2_U3222) );
  AOI21_X1 U17218 ( .B1(n16174), .B2(n16173), .A(n16172), .ZN(n16175) );
  NOR2_X1 U17219 ( .A1(n16175), .A2(n16247), .ZN(n16180) );
  AOI211_X1 U17220 ( .C1(n16178), .C2(n16177), .A(n16228), .B(n16176), .ZN(
        n16179) );
  AOI211_X1 U17221 ( .C1(n16234), .C2(n16181), .A(n16180), .B(n16179), .ZN(
        n16183) );
  OAI211_X1 U17222 ( .C1(n16184), .C2(n16254), .A(n16183), .B(n16182), .ZN(
        P2_U3225) );
  OAI21_X1 U17223 ( .B1(n16187), .B2(n16186), .A(n16185), .ZN(n16195) );
  NOR2_X1 U17224 ( .A1(n16189), .A2(n16188), .ZN(n16194) );
  AOI211_X1 U17225 ( .C1(n16192), .C2(n16191), .A(n16190), .B(n16228), .ZN(
        n16193) );
  AOI211_X1 U17226 ( .C1(n16222), .C2(n16195), .A(n16194), .B(n16193), .ZN(
        n16197) );
  OAI211_X1 U17227 ( .C1(n16198), .C2(n16254), .A(n16197), .B(n16196), .ZN(
        P2_U3228) );
  INV_X1 U17228 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n16317) );
  AOI211_X1 U17229 ( .C1(n16201), .C2(n16200), .A(n16199), .B(n16247), .ZN(
        n16206) );
  AOI211_X1 U17230 ( .C1(n16204), .C2(n16203), .A(n16202), .B(n16228), .ZN(
        n16205) );
  AOI211_X1 U17231 ( .C1(n16207), .C2(n16234), .A(n16206), .B(n16205), .ZN(
        n16209) );
  NAND2_X1 U17232 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n16208)
         );
  OAI211_X1 U17233 ( .C1(n16317), .C2(n16254), .A(n16209), .B(n16208), .ZN(
        P2_U3230) );
  INV_X1 U17234 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n16221) );
  AOI211_X1 U17235 ( .C1(n16212), .C2(n16211), .A(n16210), .B(n16228), .ZN(
        n16217) );
  AOI211_X1 U17236 ( .C1(n16215), .C2(n16214), .A(n16213), .B(n16247), .ZN(
        n16216) );
  AOI211_X1 U17237 ( .C1(n16234), .C2(n16218), .A(n16217), .B(n16216), .ZN(
        n16220) );
  NAND2_X1 U17238 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3088), .ZN(n16219)
         );
  OAI211_X1 U17239 ( .C1(n16221), .C2(n16254), .A(n16220), .B(n16219), .ZN(
        P2_U3231) );
  OAI211_X1 U17240 ( .C1(n16225), .C2(n16224), .A(n16223), .B(n16222), .ZN(
        n16226) );
  INV_X1 U17241 ( .A(n16226), .ZN(n16232) );
  AOI211_X1 U17242 ( .C1(n16230), .C2(n16229), .A(n16228), .B(n16227), .ZN(
        n16231) );
  AOI211_X1 U17243 ( .C1(n16234), .C2(n16233), .A(n16232), .B(n16231), .ZN(
        n16236) );
  OAI211_X1 U17244 ( .C1(n16295), .C2(n16254), .A(n16236), .B(n16235), .ZN(
        P2_U3224) );
  INV_X1 U17245 ( .A(n16237), .ZN(n16239) );
  OAI21_X1 U17246 ( .B1(n16239), .B2(n16238), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n16240) );
  OAI21_X1 U17247 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n16240), .ZN(n16253) );
  OAI21_X1 U17248 ( .B1(n16243), .B2(n16242), .A(n16241), .ZN(n16251) );
  AOI21_X1 U17249 ( .B1(n16246), .B2(n16245), .A(n16244), .ZN(n16248) );
  NOR2_X1 U17250 ( .A1(n16248), .A2(n16247), .ZN(n16249) );
  AOI21_X1 U17251 ( .B1(n16251), .B2(n16250), .A(n16249), .ZN(n16252) );
  OAI211_X1 U17252 ( .C1(n16255), .C2(n16254), .A(n16253), .B(n16252), .ZN(
        P2_U3223) );
  INV_X1 U17253 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n16257) );
  AOI21_X1 U17254 ( .B1(n16258), .B2(n16257), .A(n16256), .ZN(P1_U3445) );
  INV_X1 U17255 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n16271) );
  OAI21_X1 U17256 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n16260), .A(n16259), 
        .ZN(n16265) );
  OAI21_X1 U17257 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n16262), .A(n16261), 
        .ZN(n16263) );
  OAI222_X1 U17258 ( .A1(n16358), .A2(n16267), .B1(n16266), .B2(n16265), .C1(
        n16264), .C2(n16263), .ZN(n16268) );
  INV_X1 U17259 ( .A(n16268), .ZN(n16270) );
  OAI211_X1 U17260 ( .C1(n16271), .C2(n16364), .A(n16270), .B(n16269), .ZN(
        P1_U3261) );
  AOI21_X1 U17261 ( .B1(n16272), .B2(n10284), .A(n16325), .ZN(SUB_1596_U53) );
  AOI21_X1 U17262 ( .B1(n16275), .B2(n16274), .A(n16273), .ZN(n16276) );
  XOR2_X1 U17263 ( .A(n16276), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  XOR2_X1 U17264 ( .A(n16278), .B(n16277), .Z(SUB_1596_U60) );
  XOR2_X1 U17265 ( .A(n16280), .B(n16279), .Z(SUB_1596_U59) );
  NOR2_X1 U17266 ( .A1(n16282), .A2(n16281), .ZN(n16283) );
  XOR2_X1 U17267 ( .A(n16283), .B(P2_ADDR_REG_5__SCAN_IN), .Z(SUB_1596_U58) );
  XNOR2_X1 U17268 ( .A(n16285), .B(n16284), .ZN(SUB_1596_U56) );
  XOR2_X1 U17269 ( .A(n16287), .B(n16286), .Z(SUB_1596_U55) );
  AOI21_X1 U17270 ( .B1(n16290), .B2(n16289), .A(n16288), .ZN(n16291) );
  XOR2_X1 U17271 ( .A(n16291), .B(P2_ADDR_REG_9__SCAN_IN), .Z(SUB_1596_U54) );
  OAI21_X1 U17272 ( .B1(n16294), .B2(n16293), .A(n16292), .ZN(n16296) );
  XOR2_X1 U17273 ( .A(n16296), .B(n16295), .Z(SUB_1596_U70) );
  AOI21_X1 U17274 ( .B1(n16299), .B2(n16298), .A(n16297), .ZN(n16300) );
  XOR2_X1 U17275 ( .A(n16300), .B(P2_ADDR_REG_11__SCAN_IN), .Z(SUB_1596_U69)
         );
  XNOR2_X1 U17276 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n16301), .ZN(SUB_1596_U68)
         );
  AOI21_X1 U17277 ( .B1(n16304), .B2(n16303), .A(n16302), .ZN(n16305) );
  XOR2_X1 U17278 ( .A(n16305), .B(P2_ADDR_REG_13__SCAN_IN), .Z(SUB_1596_U67)
         );
  AOI21_X1 U17279 ( .B1(n16308), .B2(n16307), .A(n16306), .ZN(n16309) );
  XOR2_X1 U17280 ( .A(n16309), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  AOI21_X1 U17281 ( .B1(n16312), .B2(n16311), .A(n16310), .ZN(n16313) );
  XOR2_X1 U17282 ( .A(n16313), .B(P2_ADDR_REG_15__SCAN_IN), .Z(SUB_1596_U65)
         );
  NOR2_X1 U17283 ( .A1(n16315), .A2(n16314), .ZN(n16316) );
  XNOR2_X1 U17284 ( .A(n16317), .B(n16316), .ZN(SUB_1596_U64) );
  XOR2_X1 U17285 ( .A(n16319), .B(n16318), .Z(SUB_1596_U63) );
  XOR2_X1 U17286 ( .A(n16320), .B(P2_ADDR_REG_18__SCAN_IN), .Z(SUB_1596_U62)
         );
  AOI21_X1 U17287 ( .B1(n16323), .B2(n16322), .A(n16321), .ZN(n16324) );
  XOR2_X1 U17288 ( .A(n16324), .B(P2_ADDR_REG_6__SCAN_IN), .Z(SUB_1596_U57) );
  XOR2_X1 U17289 ( .A(n16326), .B(n16325), .Z(SUB_1596_U5) );
  NAND2_X1 U17290 ( .A1(n16328), .A2(n16327), .ZN(n16332) );
  INV_X1 U17291 ( .A(n16331), .ZN(n16329) );
  NAND2_X1 U17292 ( .A1(n16332), .A2(n16329), .ZN(n16340) );
  AOI22_X1 U17293 ( .A1(n16330), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n16339) );
  OAI21_X1 U17294 ( .B1(n16336), .B2(n16332), .A(n16331), .ZN(n16334) );
  NAND2_X1 U17295 ( .A1(n16334), .A2(n16333), .ZN(n16337) );
  AOI22_X1 U17296 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n16337), .B1(n16336), .B2(
        n16335), .ZN(n16338) );
  OAI211_X1 U17297 ( .C1(P3_IR_REG_0__SCAN_IN), .C2(n16340), .A(n16339), .B(
        n16338), .ZN(P3_U3182) );
  MUX2_X1 U17298 ( .A(n10321), .B(P1_REG2_REG_4__SCAN_IN), .S(n16341), .Z(
        n16342) );
  NAND3_X1 U17299 ( .A1(n16344), .A2(n16343), .A3(n16342), .ZN(n16345) );
  NAND3_X1 U17300 ( .A1(n16347), .A2(n16346), .A3(n16345), .ZN(n16356) );
  INV_X1 U17301 ( .A(n16348), .ZN(n16353) );
  NAND3_X1 U17302 ( .A1(n16351), .A2(n16350), .A3(n16349), .ZN(n16352) );
  NAND3_X1 U17303 ( .A1(n16354), .A2(n16353), .A3(n16352), .ZN(n16355) );
  OAI211_X1 U17304 ( .C1(n16358), .C2(n16357), .A(n16356), .B(n16355), .ZN(
        n16359) );
  NOR2_X1 U17305 ( .A1(n16360), .A2(n16359), .ZN(n16362) );
  OAI211_X1 U17306 ( .C1(n16364), .C2(n16363), .A(n16362), .B(n16361), .ZN(
        P1_U3247) );
  INV_X1 U17307 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n16365) );
  AOI22_X1 U17308 ( .A1(n16556), .A2(n16366), .B1(n16365), .B2(n16554), .ZN(
        P1_U3459) );
  XNOR2_X1 U17309 ( .A(n16367), .B(n16370), .ZN(n16389) );
  NOR2_X1 U17310 ( .A1(n16368), .A2(n16558), .ZN(n16387) );
  INV_X1 U17311 ( .A(n16389), .ZN(n16381) );
  OAI21_X1 U17312 ( .B1(n16371), .B2(n16370), .A(n16369), .ZN(n16378) );
  OAI22_X1 U17313 ( .A1(n16375), .A2(n16374), .B1(n16373), .B2(n16372), .ZN(
        n16376) );
  AOI21_X1 U17314 ( .B1(n16378), .B2(n16377), .A(n16376), .ZN(n16379) );
  OAI21_X1 U17315 ( .B1(n16381), .B2(n16380), .A(n16379), .ZN(n16385) );
  AOI211_X1 U17316 ( .C1(n8515), .C2(n16389), .A(n16387), .B(n16385), .ZN(
        n16384) );
  AOI22_X1 U17317 ( .A1(n16565), .A2(n16384), .B1(n16382), .B2(n16563), .ZN(
        P3_U3460) );
  INV_X1 U17318 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n16383) );
  AOI22_X1 U17319 ( .A1(n16569), .A2(n16384), .B1(n16383), .B2(n16566), .ZN(
        P3_U3393) );
  INV_X1 U17320 ( .A(n16411), .ZN(n16414) );
  AOI21_X1 U17321 ( .B1(n16387), .B2(n16386), .A(n16385), .ZN(n16393) );
  AOI22_X1 U17322 ( .A1(n16390), .A2(n16389), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n16388), .ZN(n16391) );
  OAI221_X1 U17323 ( .B1(n16414), .B2(n16393), .C1(n16411), .C2(n16392), .A(
        n16391), .ZN(P3_U3232) );
  OAI22_X1 U17324 ( .A1(n16395), .A2(n16544), .B1(n16394), .B2(n16542), .ZN(
        n16397) );
  AOI211_X1 U17325 ( .C1(n16495), .C2(n16398), .A(n16397), .B(n16396), .ZN(
        n16399) );
  AOI22_X1 U17326 ( .A1(n16553), .A2(n16399), .B1(n10304), .B2(n16551), .ZN(
        P1_U3529) );
  AOI22_X1 U17327 ( .A1(n16556), .A2(n16399), .B1(n9276), .B2(n16554), .ZN(
        P1_U3462) );
  INV_X1 U17328 ( .A(n16400), .ZN(n16401) );
  NAND2_X1 U17329 ( .A1(n16402), .A2(n16401), .ZN(n16403) );
  OAI21_X1 U17330 ( .B1(n16405), .B2(n16404), .A(n16403), .ZN(n16408) );
  INV_X1 U17331 ( .A(n16406), .ZN(n16407) );
  AOI211_X1 U17332 ( .C1(n16410), .C2(n16409), .A(n16408), .B(n16407), .ZN(
        n16412) );
  AOI22_X1 U17333 ( .A1(n16414), .A2(n16413), .B1(n16412), .B2(n16411), .ZN(
        P3_U3231) );
  INV_X1 U17334 ( .A(n16415), .ZN(n16420) );
  OAI211_X1 U17335 ( .C1(n16418), .C2(n16579), .A(n16417), .B(n16416), .ZN(
        n16419) );
  AOI21_X1 U17336 ( .B1(n16420), .B2(n16583), .A(n16419), .ZN(n16421) );
  AOI22_X1 U17337 ( .A1(n14740), .A2(n16421), .B1(n11182), .B2(n16584), .ZN(
        P2_U3501) );
  AOI22_X1 U17338 ( .A1(n16534), .A2(n16421), .B1(n10044), .B2(n16585), .ZN(
        P2_U3436) );
  AOI22_X1 U17339 ( .A1(n16423), .A2(n8515), .B1(n16422), .B2(n16471), .ZN(
        n16424) );
  AND2_X1 U17340 ( .A1(n16425), .A2(n16424), .ZN(n16428) );
  AOI22_X1 U17341 ( .A1(n16565), .A2(n16428), .B1(n16426), .B2(n16563), .ZN(
        P3_U3462) );
  INV_X1 U17342 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n16427) );
  AOI22_X1 U17343 ( .A1(n16569), .A2(n16428), .B1(n16427), .B2(n16566), .ZN(
        P3_U3399) );
  OAI22_X1 U17344 ( .A1(n16430), .A2(n16544), .B1(n16429), .B2(n16542), .ZN(
        n16433) );
  INV_X1 U17345 ( .A(n16431), .ZN(n16432) );
  AOI211_X1 U17346 ( .C1(n16495), .C2(n16434), .A(n16433), .B(n16432), .ZN(
        n16436) );
  AOI22_X1 U17347 ( .A1(n16553), .A2(n16436), .B1(n10307), .B2(n16551), .ZN(
        P1_U3531) );
  INV_X1 U17348 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n16435) );
  AOI22_X1 U17349 ( .A1(n16556), .A2(n16436), .B1(n16435), .B2(n16554), .ZN(
        P1_U3468) );
  AOI22_X1 U17350 ( .A1(n16438), .A2(n16561), .B1(n16437), .B2(n16471), .ZN(
        n16440) );
  AND2_X1 U17351 ( .A1(n16440), .A2(n16439), .ZN(n16443) );
  AOI22_X1 U17352 ( .A1(n16565), .A2(n16443), .B1(n16441), .B2(n16563), .ZN(
        P3_U3463) );
  INV_X1 U17353 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n16442) );
  AOI22_X1 U17354 ( .A1(n16569), .A2(n16443), .B1(n16442), .B2(n16566), .ZN(
        P3_U3402) );
  AOI21_X1 U17355 ( .B1(n16446), .B2(n16445), .A(n16444), .ZN(n16447) );
  OAI21_X1 U17356 ( .B1(n16448), .B2(n16544), .A(n16447), .ZN(n16452) );
  NOR2_X1 U17357 ( .A1(n16450), .A2(n16449), .ZN(n16451) );
  AOI211_X1 U17358 ( .C1(n16547), .C2(n16453), .A(n16452), .B(n16451), .ZN(
        n16455) );
  AOI22_X1 U17359 ( .A1(n16553), .A2(n16455), .B1(n9343), .B2(n16551), .ZN(
        P1_U3532) );
  INV_X1 U17360 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n16454) );
  AOI22_X1 U17361 ( .A1(n16556), .A2(n16455), .B1(n16454), .B2(n16554), .ZN(
        P1_U3471) );
  AOI22_X1 U17362 ( .A1(n16457), .A2(n8515), .B1(n16456), .B2(n16471), .ZN(
        n16458) );
  AND2_X1 U17363 ( .A1(n16459), .A2(n16458), .ZN(n16462) );
  AOI22_X1 U17364 ( .A1(n16565), .A2(n16462), .B1(n16460), .B2(n16563), .ZN(
        P3_U3464) );
  INV_X1 U17365 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n16461) );
  AOI22_X1 U17366 ( .A1(n16569), .A2(n16462), .B1(n16461), .B2(n16566), .ZN(
        P3_U3405) );
  OAI22_X1 U17367 ( .A1(n16464), .A2(n16544), .B1(n16463), .B2(n16542), .ZN(
        n16467) );
  INV_X1 U17368 ( .A(n16465), .ZN(n16466) );
  AOI211_X1 U17369 ( .C1(n16495), .C2(n16468), .A(n16467), .B(n16466), .ZN(
        n16469) );
  AOI22_X1 U17370 ( .A1(n16553), .A2(n16469), .B1(n9367), .B2(n16551), .ZN(
        P1_U3533) );
  AOI22_X1 U17371 ( .A1(n16556), .A2(n16469), .B1(n9366), .B2(n16554), .ZN(
        P1_U3474) );
  AOI22_X1 U17372 ( .A1(n16472), .A2(n8515), .B1(n16471), .B2(n16470), .ZN(
        n16473) );
  AND2_X1 U17373 ( .A1(n16474), .A2(n16473), .ZN(n16477) );
  AOI22_X1 U17374 ( .A1(n16565), .A2(n16477), .B1(n16475), .B2(n16563), .ZN(
        P3_U3465) );
  INV_X1 U17375 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n16476) );
  AOI22_X1 U17376 ( .A1(n16569), .A2(n16477), .B1(n16476), .B2(n16566), .ZN(
        P3_U3408) );
  INV_X1 U17377 ( .A(n16478), .ZN(n16479) );
  OAI22_X1 U17378 ( .A1(n16480), .A2(n16544), .B1(n16479), .B2(n16542), .ZN(
        n16482) );
  AOI211_X1 U17379 ( .C1(n16495), .C2(n16483), .A(n16482), .B(n16481), .ZN(
        n16484) );
  AOI22_X1 U17380 ( .A1(n16553), .A2(n16484), .B1(n9399), .B2(n16551), .ZN(
        P1_U3535) );
  AOI22_X1 U17381 ( .A1(n16556), .A2(n16484), .B1(n9403), .B2(n16554), .ZN(
        P1_U3480) );
  NOR2_X1 U17382 ( .A1(n16485), .A2(n16558), .ZN(n16487) );
  AOI211_X1 U17383 ( .C1(n16561), .C2(n16488), .A(n16487), .B(n16486), .ZN(
        n16490) );
  AOI22_X1 U17384 ( .A1(n16565), .A2(n16490), .B1(n11269), .B2(n16563), .ZN(
        P3_U3467) );
  INV_X1 U17385 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n16489) );
  AOI22_X1 U17386 ( .A1(n16569), .A2(n16490), .B1(n16489), .B2(n16566), .ZN(
        P3_U3414) );
  OAI22_X1 U17387 ( .A1(n16491), .A2(n16544), .B1(n8004), .B2(n16542), .ZN(
        n16493) );
  AOI211_X1 U17388 ( .C1(n16495), .C2(n16494), .A(n16493), .B(n16492), .ZN(
        n16497) );
  AOI22_X1 U17389 ( .A1(n16553), .A2(n16497), .B1(n16496), .B2(n16551), .ZN(
        P1_U3536) );
  AOI22_X1 U17390 ( .A1(n16556), .A2(n16497), .B1(n9419), .B2(n16554), .ZN(
        P1_U3483) );
  NOR2_X1 U17391 ( .A1(n16498), .A2(n16558), .ZN(n16499) );
  AOI21_X1 U17392 ( .B1(n16500), .B2(n8515), .A(n16499), .ZN(n16501) );
  AND2_X1 U17393 ( .A1(n16502), .A2(n16501), .ZN(n16505) );
  AOI22_X1 U17394 ( .A1(n16565), .A2(n16505), .B1(n16503), .B2(n16563), .ZN(
        P3_U3468) );
  INV_X1 U17395 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n16504) );
  AOI22_X1 U17396 ( .A1(n16569), .A2(n16505), .B1(n16504), .B2(n16566), .ZN(
        P3_U3417) );
  INV_X1 U17397 ( .A(n16506), .ZN(n16507) );
  OAI21_X1 U17398 ( .B1(n16508), .B2(n16542), .A(n16507), .ZN(n16510) );
  AOI211_X1 U17399 ( .C1(n16547), .C2(n16511), .A(n16510), .B(n16509), .ZN(
        n16512) );
  AOI22_X1 U17400 ( .A1(n16553), .A2(n16512), .B1(n9435), .B2(n16551), .ZN(
        P1_U3537) );
  AOI22_X1 U17401 ( .A1(n16556), .A2(n16512), .B1(n9439), .B2(n16554), .ZN(
        P1_U3486) );
  NOR2_X1 U17402 ( .A1(n16513), .A2(n16558), .ZN(n16515) );
  AOI211_X1 U17403 ( .C1(n16516), .C2(n16561), .A(n16515), .B(n16514), .ZN(
        n16519) );
  INV_X1 U17404 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n16517) );
  AOI22_X1 U17405 ( .A1(n16565), .A2(n16519), .B1(n16517), .B2(n16563), .ZN(
        P3_U3469) );
  INV_X1 U17406 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n16518) );
  AOI22_X1 U17407 ( .A1(n16569), .A2(n16519), .B1(n16518), .B2(n16566), .ZN(
        P3_U3420) );
  OAI21_X1 U17408 ( .B1(n16521), .B2(n16542), .A(n16520), .ZN(n16523) );
  AOI211_X1 U17409 ( .C1(n16547), .C2(n16524), .A(n16523), .B(n16522), .ZN(
        n16526) );
  AOI22_X1 U17410 ( .A1(n16553), .A2(n16526), .B1(n16525), .B2(n16551), .ZN(
        P1_U3538) );
  AOI22_X1 U17411 ( .A1(n16556), .A2(n16526), .B1(n9456), .B2(n16554), .ZN(
        P1_U3489) );
  INV_X1 U17412 ( .A(n16527), .ZN(n16531) );
  OAI21_X1 U17413 ( .B1(n7988), .B2(n16579), .A(n16528), .ZN(n16530) );
  AOI211_X1 U17414 ( .C1(n16532), .C2(n16531), .A(n16530), .B(n16529), .ZN(
        n16533) );
  AOI22_X1 U17415 ( .A1(n14740), .A2(n16533), .B1(n11193), .B2(n16584), .ZN(
        P2_U3509) );
  AOI22_X1 U17416 ( .A1(n16534), .A2(n16533), .B1(n10985), .B2(n16585), .ZN(
        P2_U3460) );
  OAI21_X1 U17417 ( .B1(n16536), .B2(n16558), .A(n16535), .ZN(n16537) );
  AOI21_X1 U17418 ( .B1(n16538), .B2(n16561), .A(n16537), .ZN(n16541) );
  AOI22_X1 U17419 ( .A1(n16565), .A2(n16541), .B1(n16539), .B2(n16563), .ZN(
        P3_U3470) );
  INV_X1 U17420 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n16540) );
  AOI22_X1 U17421 ( .A1(n16569), .A2(n16541), .B1(n16540), .B2(n16566), .ZN(
        P3_U3423) );
  OAI22_X1 U17422 ( .A1(n16545), .A2(n16544), .B1(n16543), .B2(n16542), .ZN(
        n16546) );
  AOI21_X1 U17423 ( .B1(n16548), .B2(n16547), .A(n16546), .ZN(n16549) );
  AOI22_X1 U17424 ( .A1(n16553), .A2(n16555), .B1(n16552), .B2(n16551), .ZN(
        P1_U3539) );
  AOI22_X1 U17425 ( .A1(n16556), .A2(n16555), .B1(n9481), .B2(n16554), .ZN(
        P1_U3492) );
  OAI21_X1 U17426 ( .B1(n16559), .B2(n16558), .A(n16557), .ZN(n16560) );
  AOI21_X1 U17427 ( .B1(n16562), .B2(n16561), .A(n16560), .ZN(n16568) );
  AOI22_X1 U17428 ( .A1(n16565), .A2(n16568), .B1(n16564), .B2(n16563), .ZN(
        P3_U3471) );
  INV_X1 U17429 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n16567) );
  AOI22_X1 U17430 ( .A1(n16569), .A2(n16568), .B1(n16567), .B2(n16566), .ZN(
        P3_U3426) );
  AND2_X1 U17431 ( .A1(n16570), .A2(n16583), .ZN(n16574) );
  OAI21_X1 U17432 ( .B1(n16572), .B2(n16579), .A(n16571), .ZN(n16573) );
  NOR3_X1 U17433 ( .A1(n16575), .A2(n16574), .A3(n16573), .ZN(n16577) );
  AOI22_X1 U17434 ( .A1(n14740), .A2(n16577), .B1(n11610), .B2(n16584), .ZN(
        P2_U3511) );
  INV_X1 U17435 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n16576) );
  AOI22_X1 U17436 ( .A1(n16534), .A2(n16577), .B1(n16576), .B2(n16585), .ZN(
        P2_U3466) );
  OAI21_X1 U17437 ( .B1(n7739), .B2(n16579), .A(n16578), .ZN(n16581) );
  AOI211_X1 U17438 ( .C1(n16583), .C2(n16582), .A(n16581), .B(n16580), .ZN(
        n16586) );
  AOI22_X1 U17439 ( .A1(n14740), .A2(n16586), .B1(n12271), .B2(n16584), .ZN(
        P2_U3513) );
  AOI22_X1 U17440 ( .A1(n16534), .A2(n16586), .B1(n11907), .B2(n16585), .ZN(
        P2_U3472) );
  AOI21_X1 U17441 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n16587) );
  OAI21_X1 U17442 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n16587), 
        .ZN(U28) );
  AND3_X1 U7595 ( .A1(n7897), .A2(n7896), .A3(n9950), .ZN(n9951) );
  NAND2_X2 U7601 ( .A1(n10927), .A2(n10196), .ZN(n9027) );
  INV_X2 U7552 ( .A(n14238), .ZN(n14113) );
  CLKBUF_X1 U7554 ( .A(n13800), .Z(n13811) );
  CLKBUF_X2 U7574 ( .A(n12834), .Z(n7614) );
  CLKBUF_X1 U7575 ( .A(n8951), .Z(n9010) );
  CLKBUF_X1 U7588 ( .A(n8631), .Z(n13000) );
  AND3_X1 U7596 ( .A1(n8607), .A2(n8606), .A3(n8605), .ZN(n16437) );
  NAND2_X1 U7600 ( .A1(n14529), .A2(n8189), .ZN(n14505) );
  CLKBUF_X1 U7642 ( .A(n9326), .Z(n9803) );
  CLKBUF_X1 U7658 ( .A(n13983), .Z(n13951) );
  NAND2_X1 U7659 ( .A1(n10439), .A2(n11126), .ZN(n10522) );
endmodule

