

module b21_C_SARLock_k_128_1 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227;

  NAND2_X1 U4907 ( .A1(n8029), .A2(n8028), .ZN(n8489) );
  INV_X1 U4908 ( .A(n6769), .ZN(n7787) );
  CLKBUF_X2 U4909 ( .A(n7032), .Z(n7771) );
  NAND2_X1 U4910 ( .A1(n5890), .A2(n8683), .ZN(n7032) );
  INV_X1 U4911 ( .A(n8393), .ZN(n8385) );
  XNOR2_X1 U4912 ( .A(n5157), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5163) );
  AND4_X1 U4913 ( .A1(n5831), .A2(n5828), .A3(n5830), .A4(n5829), .ZN(n5835)
         );
  INV_X1 U4914 ( .A(n5405), .ZN(n5378) );
  INV_X1 U4915 ( .A(n7994), .ZN(n7833) );
  INV_X1 U4916 ( .A(n5796), .ZN(n5261) );
  INV_X1 U4917 ( .A(n5318), .ZN(n7415) );
  AND2_X2 U4918 ( .A1(n5868), .A2(n6486), .ZN(n5934) );
  INV_X1 U4919 ( .A(n7802), .ZN(n4407) );
  NAND2_X2 U4920 ( .A1(n8037), .A2(n7402), .ZN(n6143) );
  INV_X1 U4921 ( .A(n5801), .ZN(n5732) );
  AND4_X1 U4923 ( .A1(n5730), .A2(n5729), .A3(n5728), .A4(n5727), .ZN(n9053)
         );
  INV_X2 U4924 ( .A(n5799), .ZN(n4581) );
  INV_X1 U4925 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U4926 ( .A1(n8105), .A2(n8104), .ZN(n8238) );
  OAI21_X1 U4928 ( .B1(n8775), .B2(n4465), .A(n5438), .ZN(n7260) );
  BUF_X2 U4929 ( .A(n5222), .Z(n4404) );
  INV_X1 U4930 ( .A(n6636), .ZN(n7622) );
  XNOR2_X1 U4931 ( .A(n5856), .B(n5855), .ZN(n7819) );
  INV_X1 U4932 ( .A(n6832), .ZN(n9681) );
  INV_X1 U4933 ( .A(n9087), .ZN(n8929) );
  NAND2_X1 U4934 ( .A1(n5191), .A2(n7411), .ZN(n5318) );
  OAI21_X2 U4935 ( .B1(n9457), .B2(n4865), .A(n4863), .ZN(n8947) );
  NAND2_X2 U4936 ( .A1(n7269), .A2(n7268), .ZN(n9457) );
  NAND2_X1 U4937 ( .A1(n5890), .A2(n5889), .ZN(n7746) );
  INV_X1 U4938 ( .A(n5889), .ZN(n8683) );
  AOI21_X2 U4939 ( .B1(n9762), .B2(n6504), .A(n4999), .ZN(n6511) );
  OR2_X2 U4940 ( .A1(n9763), .A2(n5905), .ZN(n6248) );
  AND2_X4 U4941 ( .A1(n9780), .A2(n8003), .ZN(n5905) );
  BUF_X4 U4942 ( .A(n7799), .Z(n4401) );
  AND2_X2 U4943 ( .A1(n5888), .A2(n8683), .ZN(n7799) );
  NOR2_X2 U4944 ( .A1(n5124), .A2(n5123), .ZN(n5125) );
  XNOR2_X2 U4945 ( .A(n5192), .B(P1_IR_REG_1__SCAN_IN), .ZN(n8855) );
  AND2_X1 U4946 ( .A1(n5868), .A2(n6486), .ZN(n4402) );
  NAND2_X2 U4947 ( .A1(n8675), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5884) );
  OAI22_X2 U4948 ( .A1(n8489), .A2(n8030), .B1(n8492), .B2(n8481), .ZN(n8470)
         );
  NOR2_X2 U4949 ( .A1(n5357), .A2(n4896), .ZN(n4895) );
  NAND2_X1 U4951 ( .A1(n9064), .A2(n9072), .ZN(n9063) );
  NAND2_X1 U4952 ( .A1(n4493), .A2(n4480), .ZN(n9124) );
  NAND2_X1 U4953 ( .A1(n9251), .A2(n8973), .ZN(n9228) );
  INV_X1 U4954 ( .A(n9710), .ZN(n7053) );
  NAND2_X1 U4955 ( .A1(n6613), .A2(n6562), .ZN(n6614) );
  NAND3_X1 U4956 ( .A1(n5195), .A2(n5197), .A3(n5196), .ZN(n4495) );
  CLKBUF_X2 U4957 ( .A(n7746), .Z(n7768) );
  CLKBUF_X2 U4958 ( .A(n5249), .Z(n7421) );
  INV_X2 U4959 ( .A(n5191), .ZN(n5359) );
  NAND2_X2 U4960 ( .A1(n5773), .A2(n6274), .ZN(n5191) );
  INV_X2 U4961 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U4962 ( .A1(n9281), .A2(n4710), .ZN(n4709) );
  INV_X1 U4963 ( .A(n8237), .ZN(n8105) );
  AND2_X1 U4964 ( .A1(n9021), .A2(n9020), .ZN(n9284) );
  INV_X1 U4965 ( .A(n9280), .ZN(n4712) );
  NAND2_X1 U4966 ( .A1(n9063), .A2(n4847), .ZN(n4846) );
  NOR2_X1 U4967 ( .A1(n8366), .A2(n7942), .ZN(n8353) );
  NAND2_X1 U4968 ( .A1(n8399), .A2(n4993), .ZN(n8376) );
  NAND2_X1 U4969 ( .A1(n7812), .A2(n7811), .ZN(n8570) );
  NAND2_X1 U4970 ( .A1(n8400), .A2(n4947), .ZN(n8399) );
  INV_X1 U4971 ( .A(n4937), .ZN(n4936) );
  AND2_X1 U4972 ( .A1(n7945), .A2(n7806), .ZN(n4828) );
  NAND2_X1 U4973 ( .A1(n4942), .A2(n8033), .ZN(n4939) );
  AND2_X1 U4974 ( .A1(n7392), .A2(n5521), .ZN(n4808) );
  NAND2_X1 U4975 ( .A1(n4735), .A2(n4733), .ZN(n8221) );
  NAND2_X1 U4976 ( .A1(n7794), .A2(n7793), .ZN(n8582) );
  OAI21_X1 U4977 ( .B1(n5461), .B2(n4587), .A(n4417), .ZN(n7393) );
  NAND2_X1 U4978 ( .A1(n5724), .A2(n5723), .ZN(n9291) );
  OR2_X1 U4979 ( .A1(n9249), .A2(n9248), .ZN(n9251) );
  NAND2_X1 U4980 ( .A1(n7027), .A2(n7026), .ZN(n7092) );
  OAI21_X1 U4981 ( .B1(n7290), .B2(n4816), .A(n4814), .ZN(n7686) );
  AOI21_X1 U4982 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9624), .A(n9619), .ZN(
        n6402) );
  NOR2_X1 U4983 ( .A1(n7980), .A2(n4986), .ZN(n4985) );
  OR2_X1 U4984 ( .A1(n6937), .A2(n7493), .ZN(n7044) );
  NAND2_X1 U4985 ( .A1(n5940), .A2(n5939), .ZN(n8206) );
  INV_X2 U4986 ( .A(n9839), .ZN(n4405) );
  OAI21_X1 U4987 ( .B1(n6746), .B2(n6703), .A(n7448), .ZN(n7082) );
  AND2_X2 U4988 ( .A1(n6568), .A2(n6553), .ZN(n9853) );
  AND2_X1 U4989 ( .A1(n9571), .A2(n6289), .ZN(n8882) );
  NAND3_X1 U4990 ( .A1(n5949), .A2(n5948), .A3(n5947), .ZN(n8283) );
  AND2_X1 U4991 ( .A1(n5973), .A2(n5972), .ZN(n9808) );
  OR2_X1 U4992 ( .A1(n6505), .A2(n9758), .ZN(n7843) );
  NOR2_X2 U4993 ( .A1(n4991), .A2(n5253), .ZN(n6749) );
  INV_X1 U4994 ( .A(n6748), .ZN(n8845) );
  NAND2_X1 U4995 ( .A1(n4456), .A2(n5925), .ZN(n8284) );
  NAND2_X2 U4996 ( .A1(n6623), .A2(n5171), .ZN(n5799) );
  INV_X1 U4997 ( .A(n4495), .ZN(n6636) );
  AND2_X2 U4998 ( .A1(n5776), .A2(n5171), .ZN(n5796) );
  NAND4_X1 U4999 ( .A1(n5226), .A2(n5225), .A3(n5224), .A4(n5223), .ZN(n6679)
         );
  AND4_X1 U5000 ( .A1(n5274), .A2(n5273), .A3(n5272), .A4(n5271), .ZN(n7676)
         );
  AND3_X1 U5001 ( .A1(n5913), .A2(n5912), .A3(n5911), .ZN(n9789) );
  NAND4_X1 U5002 ( .A1(n5918), .A2(n5917), .A3(n5916), .A4(n5915), .ZN(n6506)
         );
  NAND4_X1 U5003 ( .A1(n5205), .A2(n5204), .A3(n5203), .A4(n5202), .ZN(n6634)
         );
  NAND2_X1 U5004 ( .A1(n4585), .A2(n7013), .ZN(n5171) );
  AND3_X1 U5005 ( .A1(n5188), .A2(n5187), .A3(n5189), .ZN(n4494) );
  INV_X1 U5006 ( .A(n9779), .ZN(n9759) );
  INV_X1 U5007 ( .A(n5864), .ZN(n9780) );
  INV_X2 U5008 ( .A(n5221), .ZN(n5812) );
  INV_X2 U5009 ( .A(n5178), .ZN(n7418) );
  AND2_X1 U5010 ( .A1(n7992), .A2(n8385), .ZN(n8003) );
  INV_X1 U5011 ( .A(n7819), .ZN(n8007) );
  AND2_X2 U5012 ( .A1(n9373), .A2(n8087), .ZN(n5221) );
  NAND2_X1 U5013 ( .A1(n8087), .A2(n5161), .ZN(n5249) );
  INV_X1 U5014 ( .A(n5163), .ZN(n8087) );
  NAND2_X1 U5015 ( .A1(n5139), .A2(n5141), .ZN(n7391) );
  INV_X1 U5016 ( .A(n5161), .ZN(n9373) );
  NAND2_X1 U5017 ( .A1(n5874), .A2(n5873), .ZN(n7402) );
  XNOR2_X1 U5018 ( .A(n5160), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5161) );
  MUX2_X1 U5019 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5140), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n5141) );
  XNOR2_X1 U5020 ( .A(n5148), .B(n5147), .ZN(n7232) );
  NAND2_X1 U5021 ( .A1(n9365), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U5022 ( .A1(n4502), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5160) );
  MUX2_X1 U5023 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5875), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5877) );
  MUX2_X1 U5024 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5871), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n5874) );
  OAI21_X1 U5025 ( .B1(n5869), .B2(P2_IR_REG_26__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5875) );
  INV_X2 U5026 ( .A(n8679), .ZN(n8131) );
  OR2_X1 U5027 ( .A1(n5159), .A2(n5464), .ZN(n4635) );
  AND2_X1 U5028 ( .A1(n4885), .A2(n5158), .ZN(n4503) );
  AND2_X1 U5029 ( .A1(n4879), .A2(n4719), .ZN(n4633) );
  AND2_X1 U5030 ( .A1(n4992), .A2(n4880), .ZN(n4879) );
  NAND2_X1 U5031 ( .A1(n4672), .A2(n4671), .ZN(n5016) );
  AND2_X2 U5032 ( .A1(n4918), .A2(n4919), .ZN(n5880) );
  AND3_X1 U5033 ( .A1(n4801), .A2(n4800), .A3(n4799), .ZN(n4992) );
  NOR2_X1 U5034 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5829) );
  NOR2_X1 U5035 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P1_RD_REG_SCAN_IN), .ZN(
        n5009) );
  NOR2_X1 U5036 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5830) );
  NOR2_X1 U5037 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5828) );
  INV_X1 U5038 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5147) );
  NOR2_X1 U5039 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5120) );
  INV_X1 U5040 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6436) );
  INV_X1 U5041 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6226) );
  NOR2_X2 U5042 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5878) );
  INV_X1 U5043 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5505) );
  INV_X1 U5044 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5130) );
  INV_X1 U5045 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6134) );
  INV_X1 U5046 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5567) );
  NOR2_X1 U5047 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4801) );
  NOR2_X1 U5048 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n4800) );
  INV_X1 U5049 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5118) );
  NOR2_X1 U5050 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n4799) );
  NOR2_X1 U5051 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5832) );
  INV_X4 U5052 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U5053 ( .A(n7802), .ZN(n4406) );
  NAND2_X2 U5054 ( .A1(n6484), .A2(n9779), .ZN(n9763) );
  NAND4_X4 U5055 ( .A1(n5901), .A2(n5900), .A3(n5899), .A4(n5898), .ZN(n6484)
         );
  NOR2_X4 U5056 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5229) );
  AND2_X1 U5057 ( .A1(n9373), .A2(n8087), .ZN(n4408) );
  AND2_X1 U5058 ( .A1(n9373), .A2(n8087), .ZN(n4409) );
  AND2_X2 U5059 ( .A1(n5878), .A2(n5832), .ZN(n5941) );
  OAI21_X2 U5060 ( .B1(n7218), .B2(n4747), .A(n4744), .ZN(n8174) );
  NAND2_X2 U5061 ( .A1(n7094), .A2(n7093), .ZN(n7218) );
  AOI21_X2 U5062 ( .B1(n9242), .B2(n9255), .A(n9226), .ZN(n9213) );
  XNOR2_X2 U5063 ( .A(n6625), .B(n4495), .ZN(n7491) );
  NAND2_X1 U5064 ( .A1(n5163), .A2(n5161), .ZN(n5222) );
  INV_X1 U5065 ( .A(n7954), .ZN(n4829) );
  OR2_X1 U5066 ( .A1(n9302), .A2(n9083), .ZN(n7593) );
  AOI21_X1 U5067 ( .B1(n4964), .B2(n4963), .A(n4452), .ZN(n4962) );
  INV_X1 U5068 ( .A(n5171), .ZN(n4584) );
  NAND2_X1 U5069 ( .A1(n4874), .A2(n9168), .ZN(n4871) );
  AOI21_X1 U5070 ( .B1(n4870), .B2(n9168), .A(n4876), .ZN(n4869) );
  AOI21_X1 U5071 ( .B1(n7871), .B2(n7870), .A(n7869), .ZN(n7878) );
  NAND2_X1 U5072 ( .A1(n7915), .A2(n7921), .ZN(n4547) );
  NAND2_X1 U5073 ( .A1(n4544), .A2(n4443), .ZN(n4543) );
  NAND2_X1 U5074 ( .A1(n7924), .A2(n7923), .ZN(n4544) );
  AOI21_X1 U5075 ( .B1(n4541), .B2(n7929), .A(n4454), .ZN(n7934) );
  INV_X1 U5076 ( .A(n8722), .ZN(n4789) );
  OAI21_X1 U5077 ( .B1(n4673), .B2(n4448), .A(n7947), .ZN(n7949) );
  AOI21_X1 U5078 ( .B1(n4901), .B2(n4900), .A(n4425), .ZN(n4673) );
  XNOR2_X1 U5079 ( .A(n9796), .B(n5934), .ZN(n5935) );
  AND2_X1 U5080 ( .A1(n6552), .A2(n6489), .ZN(n6035) );
  INV_X1 U5081 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5836) );
  OR2_X1 U5082 ( .A1(n8593), .A2(n8367), .ZN(n7931) );
  NOR2_X1 U5083 ( .A1(n4631), .A2(n8608), .ZN(n4630) );
  INV_X1 U5084 ( .A(n4632), .ZN(n4631) );
  NOR2_X1 U5085 ( .A1(n8613), .A2(n8619), .ZN(n4632) );
  OR2_X1 U5086 ( .A1(n8624), .A2(n8461), .ZN(n7917) );
  OR2_X1 U5087 ( .A1(n8565), .A2(n8260), .ZN(n4621) );
  NOR2_X1 U5088 ( .A1(n7884), .A2(n4818), .ZN(n4817) );
  NAND2_X1 U5089 ( .A1(n4819), .A2(n7324), .ZN(n4818) );
  NAND2_X1 U5090 ( .A1(n7979), .A2(n4820), .ZN(n4819) );
  INV_X1 U5091 ( .A(n7875), .ZN(n4820) );
  NAND2_X1 U5092 ( .A1(n7289), .A2(n7872), .ZN(n7290) );
  OR2_X1 U5093 ( .A1(n7162), .A2(n7161), .ZN(n7864) );
  AOI21_X1 U5094 ( .B1(n4410), .B2(n4837), .A(n4836), .ZN(n4835) );
  INV_X1 U5095 ( .A(n7858), .ZN(n4836) );
  INV_X1 U5096 ( .A(n4839), .ZN(n4837) );
  OR2_X1 U5097 ( .A1(n6506), .A2(n9789), .ZN(n7842) );
  NAND2_X1 U5098 ( .A1(n4767), .A2(n5564), .ZN(n5585) );
  INV_X1 U5099 ( .A(n8744), .ZN(n4768) );
  OR2_X1 U5100 ( .A1(n9282), .A2(n9013), .ZN(n7518) );
  OR2_X1 U5101 ( .A1(n9307), .A2(n9074), .ZN(n7588) );
  OR2_X1 U5102 ( .A1(n9322), .A2(n9119), .ZN(n7586) );
  OR2_X1 U5103 ( .A1(n4691), .A2(n8977), .ZN(n4688) );
  OR2_X1 U5104 ( .A1(n9466), .A2(n8700), .ZN(n7457) );
  INV_X1 U5105 ( .A(n5736), .ZN(n4585) );
  OR2_X1 U5106 ( .A1(n7478), .A2(n9971), .ZN(n5195) );
  NAND2_X1 U5107 ( .A1(n7410), .A2(n7409), .ZN(n7477) );
  OAI21_X1 U5108 ( .B1(n5663), .B2(n5662), .A(n5661), .ZN(n5687) );
  AND2_X1 U5109 ( .A1(n5100), .A2(n5099), .ZN(n5173) );
  INV_X1 U5110 ( .A(n5565), .ZN(n5088) );
  NOR2_X1 U5111 ( .A1(n5068), .A2(n4915), .ZN(n4914) );
  INV_X1 U5112 ( .A(n5066), .ZN(n4915) );
  INV_X1 U5113 ( .A(n5484), .ZN(n5068) );
  XNOR2_X1 U5114 ( .A(n5069), .B(SI_14_), .ZN(n5484) );
  INV_X1 U5115 ( .A(n4930), .ZN(n4929) );
  OAI21_X1 U5116 ( .B1(n4933), .B2(n4931), .A(n5061), .ZN(n4930) );
  NAND2_X1 U5117 ( .A1(n4932), .A2(n5055), .ZN(n4931) );
  AND2_X1 U5118 ( .A1(n5066), .A2(n5065), .ZN(n5001) );
  INV_X1 U5119 ( .A(n4555), .ZN(n4557) );
  INV_X1 U5120 ( .A(n4559), .ZN(n4558) );
  OAI21_X1 U5121 ( .B1(n4891), .B2(n4560), .A(n5045), .ZN(n4555) );
  INV_X1 U5122 ( .A(n5019), .ZN(n4659) );
  AND2_X1 U5123 ( .A1(n4523), .A2(n4522), .ZN(n5021) );
  NAND2_X1 U5124 ( .A1(n5016), .A2(n6061), .ZN(n4522) );
  NAND2_X1 U5125 ( .A1(n4524), .A2(n6073), .ZN(n4523) );
  INV_X1 U5126 ( .A(n5016), .ZN(n4524) );
  NAND2_X1 U5127 ( .A1(n5206), .A2(n5011), .ZN(n5013) );
  AND2_X1 U5128 ( .A1(n4730), .A2(n8121), .ZN(n4729) );
  NAND2_X1 U5129 ( .A1(n4728), .A2(n8113), .ZN(n4730) );
  OR3_X1 U5130 ( .A1(n7230), .A2(n7387), .A3(n7342), .ZN(n6038) );
  AND2_X1 U5131 ( .A1(n6035), .A2(n9771), .ZN(n6050) );
  NAND2_X1 U5132 ( .A1(n4826), .A2(n4828), .ZN(n4825) );
  NAND2_X1 U5133 ( .A1(n4829), .A2(n4489), .ZN(n4826) );
  NAND2_X1 U5134 ( .A1(n7819), .A2(n7994), .ZN(n5864) );
  INV_X1 U5135 ( .A(n7998), .ZN(n7999) );
  AND2_X1 U5136 ( .A1(n7774), .A2(n7773), .ZN(n8200) );
  OR2_X1 U5137 ( .A1(n8396), .A2(n7768), .ZN(n7774) );
  AOI21_X1 U5138 ( .B1(n4942), .B2(n4941), .A(n4468), .ZN(n4940) );
  INV_X1 U5139 ( .A(n4948), .ZN(n4941) );
  AOI21_X1 U5140 ( .B1(n4969), .B2(n4414), .A(n4460), .ZN(n4968) );
  OAI21_X1 U5141 ( .B1(n7686), .B2(n7982), .A(n7891), .ZN(n8547) );
  NAND2_X1 U5142 ( .A1(n9814), .A2(n6963), .ZN(n7858) );
  INV_X2 U5143 ( .A(n6143), .ZN(n7714) );
  NAND2_X1 U5144 ( .A1(n4785), .A2(n8685), .ZN(n4784) );
  INV_X1 U5145 ( .A(n5654), .ZN(n4785) );
  INV_X1 U5146 ( .A(n8685), .ZN(n4783) );
  NAND2_X1 U5147 ( .A1(n5585), .A2(n5584), .ZN(n8788) );
  NAND2_X1 U5148 ( .A1(n4577), .A2(n5290), .ZN(n8798) );
  NOR2_X1 U5149 ( .A1(n8964), .A2(n4848), .ZN(n4847) );
  INV_X1 U5150 ( .A(n8963), .ZN(n4848) );
  AOI21_X1 U5151 ( .B1(n9073), .B2(n8990), .A(n8989), .ZN(n9051) );
  OR2_X1 U5152 ( .A1(n9302), .A2(n8962), .ZN(n8963) );
  AOI21_X1 U5153 ( .B1(n4411), .B2(n4860), .A(n4469), .ZN(n4852) );
  INV_X1 U5154 ( .A(n4859), .ZN(n4858) );
  OAI21_X1 U5155 ( .B1(n9127), .B2(n4860), .A(n4862), .ZN(n4859) );
  NAND2_X1 U5156 ( .A1(n9112), .A2(n9130), .ZN(n4862) );
  INV_X1 U5157 ( .A(n9124), .ZN(n4856) );
  AOI21_X1 U5158 ( .B1(n4874), .B2(n4877), .A(n4458), .ZN(n4872) );
  AOI21_X1 U5159 ( .B1(n4866), .B2(n4864), .A(n4447), .ZN(n4863) );
  INV_X1 U5160 ( .A(n4866), .ZN(n4865) );
  INV_X1 U5161 ( .A(n9234), .ZN(n9470) );
  INV_X1 U5162 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5137) );
  NAND2_X1 U5163 ( .A1(n4904), .A2(n4540), .ZN(n5317) );
  AOI21_X1 U5164 ( .B1(n4905), .B2(n5298), .A(n4463), .ZN(n4904) );
  AND2_X1 U5165 ( .A1(n4725), .A2(n4723), .ZN(n4722) );
  INV_X1 U5166 ( .A(n4729), .ZN(n4723) );
  NAND2_X1 U5167 ( .A1(n6217), .A2(n6218), .ZN(n6216) );
  AOI21_X1 U5168 ( .B1(n8042), .B2(n9748), .A(n8041), .ZN(n8581) );
  NAND2_X1 U5169 ( .A1(n8813), .A2(n4994), .ZN(n5791) );
  OR2_X1 U5170 ( .A1(n5712), .A2(n5711), .ZN(n4994) );
  XNOR2_X1 U5171 ( .A(n4500), .B(n4499), .ZN(n7541) );
  NAND2_X1 U5172 ( .A1(n4501), .A2(n7635), .ZN(n4500) );
  OAI21_X1 U5173 ( .B1(n7528), .B2(n7527), .A(n4446), .ZN(n4501) );
  NOR2_X1 U5174 ( .A1(n7879), .A2(n7841), .ZN(n4669) );
  OAI21_X1 U5175 ( .B1(n7880), .B2(n7821), .A(n7979), .ZN(n4670) );
  NOR2_X1 U5176 ( .A1(n7884), .A2(n7885), .ZN(n4668) );
  NAND2_X1 U5177 ( .A1(n7903), .A2(n4455), .ZN(n4549) );
  INV_X1 U5178 ( .A(n7902), .ZN(n4550) );
  NOR2_X1 U5179 ( .A1(n7908), .A2(n7907), .ZN(n7910) );
  OAI21_X1 U5180 ( .B1(n4516), .B2(n4515), .A(n4513), .ZN(n4512) );
  NOR2_X1 U5181 ( .A1(n4514), .A2(n4692), .ZN(n4513) );
  NOR2_X1 U5182 ( .A1(n7562), .A2(n4499), .ZN(n4516) );
  OAI21_X1 U5183 ( .B1(n7563), .B2(n7602), .A(n9227), .ZN(n4515) );
  AND2_X1 U5184 ( .A1(n9196), .A2(n7567), .ZN(n4511) );
  NAND2_X1 U5185 ( .A1(n4547), .A2(n4546), .ZN(n4545) );
  OAI21_X1 U5186 ( .B1(n7937), .B2(n4424), .A(n4462), .ZN(n4902) );
  NAND2_X1 U5187 ( .A1(n4902), .A2(n8368), .ZN(n4901) );
  NOR2_X1 U5188 ( .A1(n6959), .A2(n7831), .ZN(n4839) );
  AOI21_X1 U5189 ( .B1(n4788), .B2(n4794), .A(n4459), .ZN(n4787) );
  NAND2_X1 U5190 ( .A1(n4428), .A2(n4413), .ZN(n4593) );
  AOI21_X1 U5191 ( .B1(n4519), .B2(n4517), .A(n7592), .ZN(n7598) );
  AOI21_X1 U5192 ( .B1(n4520), .B2(n4481), .A(n4427), .ZN(n4519) );
  OAI21_X1 U5193 ( .B1(n4518), .B2(n7587), .A(n4482), .ZN(n4517) );
  NOR2_X1 U5194 ( .A1(n9330), .A2(n9325), .ZN(n4638) );
  INV_X1 U5195 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5133) );
  AND2_X1 U5196 ( .A1(n4927), .A2(n5173), .ZN(n4926) );
  NAND2_X1 U5197 ( .A1(n5586), .A2(n5095), .ZN(n4927) );
  INV_X1 U5198 ( .A(n5095), .ZN(n4924) );
  NOR2_X1 U5199 ( .A1(n8227), .A2(n4742), .ZN(n4741) );
  INV_X1 U5200 ( .A(n8187), .ZN(n4742) );
  INV_X1 U5201 ( .A(n7217), .ZN(n4746) );
  NAND2_X1 U5202 ( .A1(n7957), .A2(n7956), .ZN(n4890) );
  INV_X1 U5203 ( .A(n7988), .ZN(n7950) );
  NOR2_X1 U5204 ( .A1(n4554), .A2(n7953), .ZN(n4552) );
  INV_X1 U5205 ( .A(n4890), .ZN(n4554) );
  NAND2_X1 U5206 ( .A1(n8582), .A2(n8368), .ZN(n7940) );
  OR2_X1 U5207 ( .A1(n8587), .A2(n8240), .ZN(n7791) );
  NOR2_X1 U5208 ( .A1(n8582), .A2(n4614), .ZN(n4613) );
  INV_X1 U5209 ( .A(n4615), .ZN(n4614) );
  OAI21_X1 U5210 ( .B1(n4940), .B2(n4938), .A(n4464), .ZN(n4937) );
  NOR2_X1 U5211 ( .A1(n8587), .A2(n8593), .ZN(n4615) );
  OR2_X1 U5212 ( .A1(n8602), .A2(n8426), .ZN(n7929) );
  NOR2_X1 U5213 ( .A1(n8447), .A2(n4970), .ZN(n4969) );
  NOR2_X1 U5214 ( .A1(n4414), .A2(n8031), .ZN(n4970) );
  OR2_X1 U5215 ( .A1(n8641), .A2(n8551), .ZN(n7899) );
  OR2_X1 U5216 ( .A1(n8260), .A2(n8549), .ZN(n7891) );
  NAND2_X1 U5217 ( .A1(n9832), .A2(n4627), .ZN(n4626) );
  NOR2_X1 U5218 ( .A1(n7196), .A2(n7162), .ZN(n4627) );
  INV_X1 U5219 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6797) );
  NAND2_X1 U5220 ( .A1(n6729), .A2(n4839), .ZN(n4838) );
  NAND2_X1 U5221 ( .A1(n4536), .A2(n4535), .ZN(n7853) );
  NAND2_X1 U5222 ( .A1(n8283), .A2(n9803), .ZN(n7823) );
  NOR2_X1 U5223 ( .A1(n8423), .A2(n7925), .ZN(n8415) );
  NAND2_X1 U5224 ( .A1(n8415), .A2(n8414), .ZN(n8413) );
  OR2_X1 U5225 ( .A1(n6222), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6223) );
  INV_X1 U5226 ( .A(n5501), .ZN(n4591) );
  NOR2_X1 U5227 ( .A1(n7248), .A2(n4590), .ZN(n4589) );
  INV_X1 U5228 ( .A(n5462), .ZN(n4590) );
  NAND2_X1 U5229 ( .A1(n7393), .A2(n7395), .ZN(n4809) );
  AND2_X1 U5230 ( .A1(n7013), .A2(n8929), .ZN(n7668) );
  OR2_X1 U5231 ( .A1(n9285), .A2(n9037), .ZN(n8993) );
  NAND2_X1 U5232 ( .A1(n9228), .A2(n8976), .ZN(n4693) );
  NOR2_X1 U5233 ( .A1(n8700), .A2(n7233), .ZN(n4644) );
  AND2_X1 U5234 ( .A1(n7150), .A2(n4473), .ZN(n4884) );
  NAND2_X1 U5235 ( .A1(n7044), .A2(n7043), .ZN(n7143) );
  NOR2_X1 U5236 ( .A1(n5306), .A2(n5305), .ZN(n5334) );
  NAND2_X1 U5237 ( .A1(n8847), .A2(n6758), .ZN(n7448) );
  NOR2_X1 U5238 ( .A1(n7153), .A2(n7233), .ZN(n7243) );
  INV_X1 U5239 ( .A(n7391), .ZN(n5745) );
  NAND2_X1 U5240 ( .A1(n5793), .A2(n5792), .ZN(n7406) );
  NAND2_X1 U5241 ( .A1(n5720), .A2(n5719), .ZN(n5793) );
  NOR2_X1 U5242 ( .A1(n4888), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n4887) );
  NAND2_X1 U5243 ( .A1(n5147), .A2(n4889), .ZN(n4888) );
  INV_X1 U5244 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4889) );
  NAND2_X1 U5245 ( .A1(n5643), .A2(n5116), .ZN(n5663) );
  NAND2_X1 U5246 ( .A1(n4803), .A2(n4802), .ZN(n5134) );
  AOI21_X1 U5247 ( .B1(n4805), .B2(n5464), .A(n5464), .ZN(n4802) );
  AND2_X1 U5248 ( .A1(n4806), .A2(n5137), .ZN(n4805) );
  NAND2_X1 U5249 ( .A1(n5134), .A2(n5133), .ZN(n5150) );
  AND2_X1 U5250 ( .A1(n5132), .A2(n5122), .ZN(n4807) );
  OAI21_X1 U5251 ( .B1(n5546), .B2(n5087), .A(n5086), .ZN(n5566) );
  NOR2_X2 U5252 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5275) );
  OR2_X1 U5253 ( .A1(n7778), .A2(n10185), .ZN(n7795) );
  AND2_X1 U5254 ( .A1(n4749), .A2(n7222), .ZN(n4748) );
  INV_X1 U5255 ( .A(n7224), .ZN(n4749) );
  OAI21_X1 U5256 ( .B1(n8227), .B2(n4740), .A(n4743), .ZN(n4739) );
  INV_X1 U5257 ( .A(n8061), .ZN(n4740) );
  NAND3_X1 U5258 ( .A1(n5864), .A2(n7991), .A3(n7994), .ZN(n5868) );
  NAND2_X1 U5259 ( .A1(n6372), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n7766) );
  INV_X1 U5260 ( .A(n6344), .ZN(n5939) );
  NOR2_X1 U5261 ( .A1(n8151), .A2(n4739), .ZN(n4737) );
  OR2_X1 U5262 ( .A1(n6923), .A2(n6922), .ZN(n7030) );
  NAND2_X1 U5263 ( .A1(n8074), .A2(n8073), .ZN(n8075) );
  OR2_X1 U5264 ( .A1(n6798), .A2(n6797), .ZN(n6898) );
  INV_X1 U5265 ( .A(n6794), .ZN(n4753) );
  INV_X1 U5266 ( .A(n6916), .ZN(n4752) );
  AND2_X1 U5267 ( .A1(n6895), .A2(n6892), .ZN(n4755) );
  OR2_X1 U5268 ( .A1(n8165), .A2(n8166), .ZN(n4756) );
  AND2_X1 U5269 ( .A1(n8165), .A2(n8166), .ZN(n4757) );
  INV_X1 U5270 ( .A(n7771), .ZN(n7798) );
  OR2_X1 U5271 ( .A1(n8294), .A2(n8293), .ZN(n4573) );
  XNOR2_X1 U5272 ( .A(n4571), .B(n8323), .ZN(n8309) );
  NAND2_X1 U5273 ( .A1(n4573), .A2(n4572), .ZN(n4571) );
  NAND2_X1 U5274 ( .A1(n8308), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4572) );
  NAND2_X1 U5275 ( .A1(n8309), .A2(n7708), .ZN(n8320) );
  INV_X1 U5276 ( .A(n8377), .ZN(n4944) );
  NOR2_X1 U5277 ( .A1(n4951), .A2(n4949), .ZN(n4948) );
  INV_X1 U5278 ( .A(n4953), .ZN(n4949) );
  AND2_X1 U5279 ( .A1(n7931), .A2(n8364), .ZN(n8377) );
  NAND2_X1 U5280 ( .A1(n4952), .A2(n4947), .ZN(n4946) );
  NAND2_X1 U5281 ( .A1(n8413), .A2(n7929), .ZN(n8400) );
  OR2_X1 U5282 ( .A1(n8602), .A2(n8268), .ZN(n4953) );
  NAND2_X1 U5283 ( .A1(n8456), .A2(n4969), .ZN(n4967) );
  AND2_X1 U5284 ( .A1(n8447), .A2(n7919), .ZN(n4833) );
  AND2_X1 U5285 ( .A1(n7923), .A2(n7921), .ZN(n8447) );
  AND2_X1 U5286 ( .A1(n4834), .A2(n7919), .ZN(n8448) );
  NAND2_X1 U5287 ( .A1(n8471), .A2(n4632), .ZN(n8440) );
  INV_X1 U5288 ( .A(n7724), .ZN(n6122) );
  OR2_X1 U5289 ( .A1(n8459), .A2(n8458), .ZN(n4834) );
  AND2_X1 U5290 ( .A1(n8491), .A2(n8476), .ZN(n8471) );
  NOR2_X1 U5291 ( .A1(n8631), .A2(n8515), .ZN(n8030) );
  NAND2_X1 U5292 ( .A1(n6121), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7717) );
  OR2_X1 U5293 ( .A1(n8634), .A2(n8027), .ZN(n8498) );
  NOR2_X1 U5294 ( .A1(n8506), .A2(n8631), .ZN(n8491) );
  NAND2_X1 U5295 ( .A1(n8025), .A2(n4620), .ZN(n4619) );
  NOR2_X1 U5296 ( .A1(n4621), .A2(n8634), .ZN(n4620) );
  NAND2_X1 U5297 ( .A1(n8565), .A2(n8273), .ZN(n4982) );
  NAND2_X1 U5298 ( .A1(n8024), .A2(n8023), .ZN(n8543) );
  AND2_X1 U5299 ( .A1(n7890), .A2(n7894), .ZN(n8542) );
  OR2_X1 U5300 ( .A1(n8543), .A2(n8542), .ZN(n4983) );
  NOR2_X1 U5301 ( .A1(n7378), .A2(n8260), .ZN(n8559) );
  NAND2_X1 U5302 ( .A1(n7887), .A2(n7979), .ZN(n4816) );
  NAND2_X1 U5303 ( .A1(n4815), .A2(n7887), .ZN(n4814) );
  INV_X1 U5304 ( .A(n4817), .ZN(n4815) );
  OR2_X1 U5305 ( .A1(n7196), .A2(n7186), .ZN(n7863) );
  NAND2_X1 U5306 ( .A1(n4526), .A2(n4528), .ZN(n7183) );
  AOI21_X1 U5307 ( .B1(n7973), .B2(n4530), .A(n4529), .ZN(n4528) );
  INV_X1 U5308 ( .A(n7864), .ZN(n4529) );
  AND2_X1 U5309 ( .A1(n7974), .A2(n7113), .ZN(n4987) );
  NAND2_X1 U5310 ( .A1(n7116), .A2(n7861), .ZN(n7165) );
  NAND2_X1 U5311 ( .A1(n6977), .A2(n4988), .ZN(n7114) );
  AND2_X1 U5312 ( .A1(n7973), .A2(n6957), .ZN(n4988) );
  NAND2_X1 U5313 ( .A1(n4838), .A2(n4410), .ZN(n6982) );
  INV_X1 U5314 ( .A(n6959), .ZN(n7971) );
  NAND2_X1 U5315 ( .A1(n7852), .A2(n7853), .ZN(n6959) );
  NAND2_X1 U5316 ( .A1(n6559), .A2(n6558), .ZN(n6646) );
  INV_X1 U5317 ( .A(n7828), .ZN(n6561) );
  NAND2_X1 U5318 ( .A1(n6511), .A2(n6560), .ZN(n6555) );
  NAND2_X1 U5319 ( .A1(n7991), .A2(n7817), .ZN(n9748) );
  NAND2_X1 U5320 ( .A1(n9747), .A2(n9763), .ZN(n9762) );
  OR2_X1 U5321 ( .A1(n6484), .A2(n9759), .ZN(n9749) );
  NAND2_X1 U5322 ( .A1(n7742), .A2(n7741), .ZN(n8608) );
  OR2_X1 U5323 ( .A1(n6071), .A2(n6769), .ZN(n4677) );
  NOR2_X1 U5324 ( .A1(n4440), .A2(n4676), .ZN(n4675) );
  NOR2_X1 U5325 ( .A1(n4492), .A2(n6205), .ZN(n4676) );
  AND2_X1 U5326 ( .A1(n6488), .A2(n9771), .ZN(n6567) );
  AND2_X1 U5327 ( .A1(n6012), .A2(n6015), .ZN(n9769) );
  NOR2_X1 U5328 ( .A1(n4978), .A2(n4844), .ZN(n4843) );
  INV_X1 U5329 ( .A(n5848), .ZN(n4840) );
  NAND2_X1 U5330 ( .A1(n5850), .A2(n5872), .ZN(n4844) );
  NAND2_X1 U5331 ( .A1(n5852), .A2(n4842), .ZN(n5876) );
  NOR2_X1 U5332 ( .A1(n4978), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4842) );
  NAND2_X1 U5333 ( .A1(n5839), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5854) );
  XNOR2_X1 U5334 ( .A(n5854), .B(P2_IR_REG_23__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U5335 ( .A1(n5838), .A2(n4995), .ZN(n5857) );
  INV_X1 U5336 ( .A(n5860), .ZN(n5838) );
  NAND2_X1 U5337 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4576) );
  NAND2_X1 U5338 ( .A1(n4763), .A2(n5369), .ZN(n8712) );
  NAND2_X1 U5339 ( .A1(n5348), .A2(n6873), .ZN(n4763) );
  NOR2_X1 U5340 ( .A1(n8766), .A2(n4774), .ZN(n4786) );
  NOR2_X1 U5341 ( .A1(n4775), .A2(n4778), .ZN(n4774) );
  AOI21_X1 U5342 ( .B1(n8765), .B2(n4777), .A(n4780), .ZN(n4776) );
  NOR2_X1 U5343 ( .A1(n4781), .A2(n4778), .ZN(n4777) );
  XNOR2_X1 U5344 ( .A(n5262), .B(n4581), .ZN(n5263) );
  NAND2_X1 U5345 ( .A1(n4765), .A2(n4762), .ZN(n4761) );
  INV_X1 U5346 ( .A(n4434), .ZN(n4762) );
  NOR2_X1 U5347 ( .A1(n4796), .A2(n8758), .ZN(n4795) );
  NOR2_X1 U5348 ( .A1(n4797), .A2(n8705), .ZN(n4796) );
  NAND2_X1 U5349 ( .A1(n5392), .A2(n5391), .ZN(n8775) );
  XNOR2_X1 U5350 ( .A(n5240), .B(n4581), .ZN(n5245) );
  OAI21_X1 U5351 ( .B1(n4497), .B2(n4496), .A(n4453), .ZN(n7605) );
  AND4_X1 U5352 ( .A1(n5296), .A2(n5295), .A3(n5294), .A4(n5293), .ZN(n6748)
         );
  NOR2_X1 U5353 ( .A1(n9546), .A2(n9545), .ZN(n9544) );
  AOI21_X1 U5354 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n6323), .A(n6318), .ZN(
        n6396) );
  NAND2_X1 U5355 ( .A1(n7480), .A2(n7479), .ZN(n9282) );
  AND2_X1 U5356 ( .A1(n7518), .A2(n7658), .ZN(n8995) );
  OR2_X1 U5357 ( .A1(n9051), .A2(n4698), .ZN(n4695) );
  NAND2_X1 U5358 ( .A1(n8992), .A2(n4699), .ZN(n4698) );
  NAND2_X1 U5359 ( .A1(n4697), .A2(n8992), .ZN(n4696) );
  INV_X1 U5360 ( .A(n4700), .ZN(n4697) );
  AND2_X1 U5361 ( .A1(n4695), .A2(n4694), .ZN(n9010) );
  AND2_X1 U5362 ( .A1(n4696), .A2(n9018), .ZN(n4694) );
  INV_X1 U5363 ( .A(n9044), .ZN(n9076) );
  OR2_X1 U5364 ( .A1(n9094), .A2(n9307), .ZN(n9084) );
  INV_X1 U5365 ( .A(n4704), .ZN(n4703) );
  OAI22_X1 U5366 ( .A1(n4707), .A2(n7510), .B1(n8986), .B2(n8985), .ZN(n4704)
         );
  OR2_X1 U5367 ( .A1(n9317), .A2(n9130), .ZN(n9101) );
  INV_X1 U5368 ( .A(n9125), .ZN(n4706) );
  INV_X1 U5369 ( .A(n8959), .ZN(n4861) );
  NAND2_X1 U5370 ( .A1(n9322), .A2(n9142), .ZN(n8959) );
  NOR2_X1 U5371 ( .A1(n9126), .A2(n9127), .ZN(n9125) );
  NAND2_X1 U5372 ( .A1(n9138), .A2(n8957), .ZN(n4493) );
  OR2_X1 U5373 ( .A1(n9325), .A2(n9163), .ZN(n8957) );
  AOI21_X1 U5374 ( .B1(n4685), .B2(n4683), .A(n4682), .ZN(n4681) );
  INV_X1 U5375 ( .A(n4685), .ZN(n4684) );
  INV_X1 U5376 ( .A(n8978), .ZN(n4682) );
  NOR2_X1 U5377 ( .A1(n9187), .A2(n9335), .ZN(n9170) );
  INV_X1 U5378 ( .A(n4877), .ZN(n4875) );
  AND2_X1 U5379 ( .A1(n9220), .A2(n9230), .ZN(n4877) );
  INV_X1 U5380 ( .A(n7565), .ZN(n9196) );
  NOR2_X1 U5381 ( .A1(n9213), .A2(n9212), .ZN(n9211) );
  NOR2_X1 U5382 ( .A1(n7355), .A2(n9499), .ZN(n9260) );
  INV_X1 U5383 ( .A(n4715), .ZN(n4714) );
  OAI21_X1 U5384 ( .B1(n7043), .B2(n4717), .A(n7543), .ZN(n4715) );
  AND2_X1 U5385 ( .A1(n5398), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U5386 ( .A1(n4883), .A2(n4881), .ZN(n7267) );
  AOI21_X1 U5387 ( .B1(n7149), .B2(n4884), .A(n4882), .ZN(n4881) );
  NAND2_X1 U5388 ( .A1(n7148), .A2(n4884), .ZN(n4883) );
  NOR2_X1 U5389 ( .A1(n7233), .A2(n8841), .ZN(n4882) );
  INV_X1 U5390 ( .A(n7478), .ZN(n5588) );
  OR2_X1 U5391 ( .A1(n5350), .A2(n5349), .ZN(n5371) );
  OAI21_X1 U5392 ( .B1(n7076), .B2(n7085), .A(n6944), .ZN(n6945) );
  AND2_X1 U5393 ( .A1(n6629), .A2(n6628), .ZN(n9253) );
  AND2_X1 U5394 ( .A1(n7633), .A2(n7447), .ZN(n6718) );
  NAND2_X1 U5395 ( .A1(n6822), .A2(n7630), .ZN(n6746) );
  OR2_X1 U5396 ( .A1(n7610), .A2(n6628), .ZN(n9467) );
  INV_X1 U5397 ( .A(n9253), .ZN(n9465) );
  AND2_X1 U5398 ( .A1(n6631), .A2(n6630), .ZN(n9234) );
  NAND2_X1 U5399 ( .A1(n5738), .A2(n8929), .ZN(n6623) );
  INV_X1 U5400 ( .A(n9467), .ZN(n9254) );
  AND2_X1 U5401 ( .A1(n4879), .A2(n5125), .ZN(n4720) );
  NAND2_X1 U5402 ( .A1(n4917), .A2(n5642), .ZN(n5643) );
  NAND2_X1 U5403 ( .A1(n4461), .A2(n5130), .ZN(n4604) );
  INV_X1 U5404 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4605) );
  INV_X1 U5405 ( .A(n4807), .ZN(n4606) );
  AND2_X1 U5406 ( .A1(n4879), .A2(n4878), .ZN(n5465) );
  AND2_X1 U5407 ( .A1(n5465), .A2(n5130), .ZN(n5486) );
  NOR2_X1 U5408 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5131) );
  NAND2_X1 U5409 ( .A1(n4913), .A2(n5071), .ZN(n5504) );
  NAND2_X1 U5410 ( .A1(n5067), .A2(n4914), .ZN(n4913) );
  NAND2_X1 U5411 ( .A1(n5067), .A2(n5066), .ZN(n5485) );
  NAND2_X1 U5412 ( .A1(n4928), .A2(n5055), .ZN(n5440) );
  NAND2_X1 U5413 ( .A1(n5051), .A2(n4933), .ZN(n4928) );
  INV_X1 U5414 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U5415 ( .A1(n4897), .A2(n5034), .ZN(n5358) );
  NAND2_X1 U5416 ( .A1(n5342), .A2(n5341), .ZN(n4897) );
  NOR2_X1 U5417 ( .A1(n4659), .A2(n4658), .ZN(n4655) );
  INV_X1 U5418 ( .A(SI_3_), .ZN(n4521) );
  NAND2_X1 U5419 ( .A1(n5015), .A2(n5014), .ZN(n5228) );
  NAND2_X1 U5420 ( .A1(n8034), .A2(n7942), .ZN(n4539) );
  AOI21_X1 U5421 ( .B1(n4729), .B2(n4731), .A(n4726), .ZN(n4725) );
  OAI21_X1 U5422 ( .B1(n8123), .B2(n4727), .A(n8122), .ZN(n4726) );
  NAND2_X1 U5423 ( .A1(n4728), .A2(n8113), .ZN(n4727) );
  AND4_X1 U5424 ( .A1(n6049), .A2(n6048), .A3(n6047), .A4(n6046), .ZN(n6963)
         );
  INV_X1 U5425 ( .A(n8449), .ZN(n8482) );
  NAND2_X1 U5426 ( .A1(n7723), .A2(n7722), .ZN(n8624) );
  NAND2_X1 U5427 ( .A1(n7735), .A2(n7734), .ZN(n8613) );
  OR2_X1 U5428 ( .A1(n6070), .A2(n6769), .ZN(n5973) );
  INV_X1 U5429 ( .A(n8259), .ZN(n8248) );
  NOR2_X1 U5430 ( .A1(n6052), .A2(n6051), .ZN(n8245) );
  AND2_X1 U5431 ( .A1(n4824), .A2(n4822), .ZN(n7815) );
  INV_X1 U5432 ( .A(n4823), .ZN(n4822) );
  NAND2_X1 U5433 ( .A1(n8001), .A2(n8000), .ZN(n4811) );
  OR2_X1 U5434 ( .A1(n7032), .A2(n10101), .ZN(n5917) );
  OR2_X1 U5435 ( .A1(n7746), .A2(n5914), .ZN(n5916) );
  NAND2_X1 U5436 ( .A1(n6200), .A2(n4477), .ZN(n6217) );
  NAND2_X1 U5437 ( .A1(n4841), .A2(n5837), .ZN(n6738) );
  NAND2_X1 U5438 ( .A1(n9768), .A2(n6495), .ZN(n8538) );
  AND2_X1 U5439 ( .A1(n8579), .A2(n9815), .ZN(n4610) );
  NOR2_X1 U5440 ( .A1(n8578), .A2(n8644), .ZN(n4611) );
  NOR2_X1 U5441 ( .A1(n6083), .A2(P2_U3152), .ZN(n9777) );
  NAND2_X1 U5442 ( .A1(n8798), .A2(n5324), .ZN(n5332) );
  NAND2_X1 U5443 ( .A1(n4601), .A2(n4600), .ZN(n4596) );
  NAND2_X1 U5444 ( .A1(n5791), .A2(n5790), .ZN(n5823) );
  INV_X1 U5445 ( .A(n5823), .ZN(n4580) );
  NAND2_X1 U5446 ( .A1(n5198), .A2(n4583), .ZN(n4582) );
  OR2_X1 U5447 ( .A1(n5261), .A2(n6636), .ZN(n5198) );
  NAND2_X1 U5448 ( .A1(n5378), .A2(n6625), .ZN(n4583) );
  AND4_X1 U5449 ( .A1(n5169), .A2(n5168), .A3(n5167), .A4(n5166), .ZN(n9074)
         );
  NAND2_X1 U5450 ( .A1(n5669), .A2(n5668), .ZN(n9302) );
  INV_X1 U5451 ( .A(n8837), .ZN(n9121) );
  AND4_X1 U5452 ( .A1(n5621), .A2(n5620), .A3(n5619), .A4(n5618), .ZN(n9119)
         );
  INV_X1 U5453 ( .A(n9181), .ZN(n8955) );
  AND2_X1 U5454 ( .A1(n7063), .A2(n9709), .ZN(n8819) );
  OR2_X1 U5455 ( .A1(n7609), .A2(n8929), .ZN(n4509) );
  INV_X1 U5456 ( .A(n7670), .ZN(n4508) );
  NOR2_X1 U5457 ( .A1(n4419), .A2(n7671), .ZN(n4510) );
  AND4_X1 U5458 ( .A1(n5816), .A2(n5815), .A3(n5814), .A4(n5813), .ZN(n9013)
         );
  INV_X1 U5459 ( .A(n9074), .ZN(n9106) );
  INV_X1 U5460 ( .A(n9119), .ZN(n9142) );
  INV_X1 U5461 ( .A(n9208), .ZN(n9255) );
  AOI21_X1 U5462 ( .B1(n9363), .B2(n7415), .A(n7432), .ZN(n8939) );
  NAND2_X1 U5463 ( .A1(n9686), .A2(n6663), .ZN(n9476) );
  INV_X1 U5464 ( .A(n7840), .ZN(n4662) );
  INV_X1 U5465 ( .A(n7839), .ZN(n4663) );
  OAI21_X1 U5466 ( .B1(n7839), .B2(n4450), .A(n4666), .ZN(n4665) );
  NOR2_X1 U5467 ( .A1(n7832), .A2(n7831), .ZN(n4666) );
  AOI21_X1 U5468 ( .B1(n4664), .B2(n4661), .A(n4660), .ZN(n7849) );
  NAND2_X1 U5469 ( .A1(n7847), .A2(n7848), .ZN(n4660) );
  NAND2_X1 U5470 ( .A1(n4665), .A2(n7821), .ZN(n4664) );
  NAND2_X1 U5471 ( .A1(n4663), .A2(n4662), .ZN(n4661) );
  NAND2_X1 U5472 ( .A1(n4562), .A2(n7841), .ZN(n4561) );
  NAND2_X1 U5473 ( .A1(n7865), .A2(n7864), .ZN(n4562) );
  AOI21_X1 U5474 ( .B1(n4667), .B2(n4420), .A(n4548), .ZN(n7908) );
  NAND2_X1 U5475 ( .A1(n4550), .A2(n4549), .ZN(n4548) );
  INV_X1 U5476 ( .A(n7564), .ZN(n4514) );
  NOR2_X1 U5477 ( .A1(n4831), .A2(n7821), .ZN(n4546) );
  NAND2_X1 U5478 ( .A1(n4512), .A2(n4511), .ZN(n7572) );
  INV_X1 U5479 ( .A(n7943), .ZN(n4903) );
  NOR2_X1 U5480 ( .A1(n7944), .A2(n4899), .ZN(n4898) );
  NOR2_X1 U5481 ( .A1(n7841), .A2(n8582), .ZN(n4899) );
  AOI21_X1 U5482 ( .B1(n7585), .B2(n8981), .A(n8983), .ZN(n4518) );
  OAI21_X1 U5483 ( .B1(n7585), .B2(n7583), .A(n7582), .ZN(n4520) );
  NOR2_X1 U5484 ( .A1(n9242), .A2(n9265), .ZN(n4647) );
  OR2_X1 U5485 ( .A1(n4807), .A2(n5464), .ZN(n4806) );
  INV_X1 U5486 ( .A(n5071), .ZN(n4912) );
  INV_X1 U5487 ( .A(n4914), .ZN(n4909) );
  INV_X1 U5488 ( .A(n5076), .ZN(n4908) );
  NAND2_X1 U5489 ( .A1(n5079), .A2(n5078), .ZN(n5082) );
  INV_X1 U5490 ( .A(n5439), .ZN(n4932) );
  NAND2_X1 U5491 ( .A1(n5058), .A2(n5057), .ZN(n5061) );
  INV_X1 U5492 ( .A(n5002), .ZN(n4560) );
  AOI21_X1 U5493 ( .B1(n4891), .B2(n4894), .A(n4560), .ZN(n4559) );
  INV_X1 U5494 ( .A(n5034), .ZN(n4896) );
  OR2_X1 U5495 ( .A1(n8570), .A2(n7814), .ZN(n7818) );
  INV_X1 U5496 ( .A(n4969), .ZN(n4963) );
  NAND2_X1 U5497 ( .A1(n4968), .A2(n4966), .ZN(n4965) );
  INV_X1 U5498 ( .A(n7338), .ZN(n4986) );
  INV_X1 U5499 ( .A(n7861), .ZN(n4531) );
  NOR2_X1 U5500 ( .A1(n6645), .A2(n4956), .ZN(n4955) );
  INV_X1 U5501 ( .A(n6558), .ZN(n4956) );
  AND2_X1 U5502 ( .A1(n6726), .A2(n6643), .ZN(n4954) );
  NOR2_X1 U5503 ( .A1(n6652), .A2(n6728), .ZN(n6731) );
  NAND2_X1 U5504 ( .A1(n4617), .A2(n6587), .ZN(n6652) );
  INV_X1 U5505 ( .A(n6564), .ZN(n4617) );
  NAND2_X1 U5506 ( .A1(n4678), .A2(n6643), .ZN(n7830) );
  INV_X1 U5507 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U5508 ( .A1(n5870), .A2(n4979), .ZN(n4978) );
  INV_X1 U5509 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5870) );
  NOR2_X1 U5510 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n4732) );
  INV_X1 U5511 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5861) );
  INV_X1 U5512 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5833) );
  OR2_X1 U5513 ( .A1(n6137), .A2(n6136), .ZN(n6222) );
  OR2_X1 U5514 ( .A1(n6090), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U5515 ( .A1(n5607), .A2(n5608), .ZN(n4798) );
  INV_X1 U5516 ( .A(n8767), .ZN(n4778) );
  INV_X1 U5517 ( .A(n4595), .ZN(n4594) );
  OAI21_X1 U5518 ( .B1(n4597), .B2(n4485), .A(n4787), .ZN(n4595) );
  INV_X1 U5519 ( .A(n5584), .ZN(n4598) );
  INV_X1 U5520 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5305) );
  AOI21_X1 U5521 ( .B1(n7600), .B2(n4498), .A(n7601), .ZN(n4497) );
  AND2_X1 U5522 ( .A1(n9018), .A2(n7599), .ZN(n4498) );
  NOR2_X1 U5523 ( .A1(n7658), .A2(n7602), .ZN(n4496) );
  NOR2_X1 U5524 ( .A1(n9297), .A2(n9302), .ZN(n4652) );
  NAND2_X1 U5525 ( .A1(n4652), .A2(n9036), .ZN(n4651) );
  NAND2_X1 U5526 ( .A1(n4708), .A2(n4416), .ZN(n4707) );
  INV_X1 U5527 ( .A(n8985), .ZN(n4708) );
  INV_X1 U5528 ( .A(n4707), .ZN(n4705) );
  INV_X1 U5529 ( .A(n8961), .ZN(n4853) );
  AND2_X1 U5530 ( .A1(n4688), .A2(n4686), .ZN(n4685) );
  INV_X1 U5531 ( .A(n8979), .ZN(n4686) );
  INV_X1 U5532 ( .A(n4689), .ZN(n4683) );
  INV_X1 U5533 ( .A(n4872), .ZN(n4870) );
  NOR2_X1 U5534 ( .A1(n8977), .A2(n4690), .ZN(n4689) );
  AND2_X1 U5535 ( .A1(n5573), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5591) );
  NOR2_X1 U5536 ( .A1(n4692), .A2(n8975), .ZN(n4691) );
  OR2_X1 U5537 ( .A1(n9265), .A2(n7454), .ZN(n8973) );
  OR2_X1 U5538 ( .A1(n5470), .A2(n5469), .ZN(n5490) );
  AND2_X1 U5539 ( .A1(n7347), .A2(n4867), .ZN(n4866) );
  INV_X1 U5540 ( .A(n7270), .ZN(n4864) );
  NAND2_X1 U5541 ( .A1(n9513), .A2(n4644), .ZN(n4643) );
  NAND2_X1 U5542 ( .A1(n5419), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5446) );
  NAND2_X1 U5543 ( .A1(n9170), .A2(n4638), .ZN(n9145) );
  NAND2_X1 U5544 ( .A1(n9260), .A2(n4647), .ZN(n9238) );
  AND2_X1 U5545 ( .A1(n4887), .A2(n5126), .ZN(n4885) );
  AND2_X1 U5546 ( .A1(n5792), .A2(n5718), .ZN(n5719) );
  OAI21_X1 U5547 ( .B1(n5687), .B2(n5686), .A(n5685), .ZN(n5693) );
  AND2_X1 U5548 ( .A1(n5713), .A2(n5691), .ZN(n5692) );
  NAND2_X1 U5549 ( .A1(n5105), .A2(n5104), .ZN(n5629) );
  AOI21_X1 U5550 ( .B1(n4926), .B2(n4924), .A(n4923), .ZN(n4922) );
  INV_X1 U5551 ( .A(n4926), .ZN(n4925) );
  INV_X1 U5552 ( .A(n5100), .ZN(n4923) );
  OAI21_X1 U5553 ( .B1(n5067), .B2(n4910), .A(n4907), .ZN(n5527) );
  INV_X1 U5554 ( .A(n4911), .ZN(n4910) );
  AOI21_X1 U5555 ( .B1(n4909), .B2(n4911), .A(n4908), .ZN(n4907) );
  NOR2_X1 U5556 ( .A1(n5503), .A2(n4912), .ZN(n4911) );
  NAND2_X1 U5557 ( .A1(n5063), .A2(n5062), .ZN(n5066) );
  NOR2_X1 U5558 ( .A1(n5056), .A2(n4934), .ZN(n4933) );
  INV_X1 U5559 ( .A(n5050), .ZN(n4934) );
  INV_X1 U5560 ( .A(n4895), .ZN(n4894) );
  AOI21_X1 U5561 ( .B1(n4895), .B2(n4893), .A(n4892), .ZN(n4891) );
  INV_X1 U5562 ( .A(n5039), .ZN(n4892) );
  INV_X1 U5563 ( .A(n5341), .ZN(n4893) );
  INV_X1 U5564 ( .A(n5025), .ZN(n4905) );
  INV_X1 U5565 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4921) );
  NAND2_X1 U5566 ( .A1(n7218), .A2(n7217), .ZN(n4750) );
  NAND2_X1 U5567 ( .A1(n8188), .A2(n4741), .ZN(n4738) );
  INV_X1 U5568 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U5569 ( .A1(n6371), .A2(n6370), .ZN(n7756) );
  INV_X1 U5570 ( .A(n7744), .ZN(n6371) );
  INV_X1 U5571 ( .A(n8093), .ZN(n8096) );
  NAND2_X1 U5572 ( .A1(n6795), .A2(n6794), .ZN(n6893) );
  INV_X1 U5573 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7029) );
  OR2_X1 U5574 ( .A1(n7030), .A2(n7029), .ZN(n7100) );
  NAND2_X1 U5575 ( .A1(n6102), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6923) );
  AND2_X1 U5576 ( .A1(n8060), .A2(n8059), .ZN(n8061) );
  AOI21_X1 U5577 ( .B1(n4748), .B2(n4746), .A(n4745), .ZN(n4744) );
  INV_X1 U5578 ( .A(n4748), .ZN(n4747) );
  INV_X1 U5579 ( .A(n8048), .ZN(n4745) );
  NAND2_X1 U5580 ( .A1(n6103), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7102) );
  INV_X1 U5581 ( .A(n7100), .ZN(n6103) );
  AND2_X1 U5582 ( .A1(n7818), .A2(n7948), .ZN(n7988) );
  OAI22_X1 U5583 ( .A1(n4829), .A2(n7946), .B1(n4827), .B2(n4489), .ZN(n4823)
         );
  NOR2_X1 U5584 ( .A1(n8340), .A2(n7809), .ZN(n4827) );
  AOI21_X1 U5585 ( .B1(n4422), .B2(n4890), .A(n7964), .ZN(n4553) );
  OR2_X1 U5586 ( .A1(n6038), .A2(P2_U3152), .ZN(n6141) );
  AND2_X1 U5587 ( .A1(n6357), .A2(n4570), .ZN(n6360) );
  NAND2_X1 U5588 ( .A1(n6771), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4570) );
  NOR2_X1 U5589 ( .A1(n6360), .A2(n6359), .ZN(n6409) );
  NAND2_X1 U5590 ( .A1(n7003), .A2(n4564), .ZN(n7004) );
  OR2_X1 U5591 ( .A1(n7096), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4564) );
  NAND2_X1 U5592 ( .A1(n7004), .A2(n7005), .ZN(n7132) );
  NAND2_X1 U5593 ( .A1(n7132), .A2(n4563), .ZN(n7313) );
  OR2_X1 U5594 ( .A1(n7209), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4563) );
  CLKBUF_X1 U5595 ( .A(n5849), .Z(n6499) );
  CLKBUF_X1 U5596 ( .A(n6143), .Z(n4492) );
  AND2_X1 U5597 ( .A1(n8391), .A2(n4429), .ZN(n8338) );
  AND2_X1 U5598 ( .A1(n4539), .A2(n7806), .ZN(n4537) );
  NAND2_X1 U5599 ( .A1(n8391), .A2(n4613), .ZN(n8345) );
  AND2_X1 U5600 ( .A1(n7795), .A2(n7779), .ZN(n8384) );
  NOR2_X1 U5601 ( .A1(n8602), .A2(n4629), .ZN(n4628) );
  INV_X1 U5602 ( .A(n4630), .ZN(n4629) );
  INV_X1 U5603 ( .A(n4965), .ZN(n4964) );
  AND2_X1 U5604 ( .A1(n7762), .A2(n7761), .ZN(n8426) );
  NAND2_X1 U5605 ( .A1(n4832), .A2(n4830), .ZN(n8424) );
  AOI21_X1 U5606 ( .B1(n4833), .B2(n8458), .A(n4831), .ZN(n4830) );
  OR2_X1 U5607 ( .A1(n7717), .A2(n10040), .ZN(n7724) );
  AND2_X1 U5608 ( .A1(n7904), .A2(n8479), .ZN(n8497) );
  AOI21_X1 U5609 ( .B1(n4415), .B2(n8542), .A(n4451), .ZN(n4981) );
  AND2_X1 U5610 ( .A1(n8498), .A2(n7906), .ZN(n8512) );
  OR2_X1 U5611 ( .A1(n7695), .A2(n6120), .ZN(n7706) );
  NAND2_X1 U5612 ( .A1(n6104), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7695) );
  INV_X1 U5613 ( .A(n7102), .ZN(n6104) );
  NOR2_X1 U5614 ( .A1(n7378), .A2(n4621), .ZN(n8561) );
  AND4_X1 U5615 ( .A1(n7375), .A2(n7374), .A3(n7373), .A4(n7372), .ZN(n8047)
         );
  OR2_X1 U5616 ( .A1(n7290), .A2(n4821), .ZN(n4813) );
  AND2_X1 U5617 ( .A1(n7291), .A2(n7979), .ZN(n7325) );
  NOR2_X1 U5618 ( .A1(n4626), .A2(n7337), .ZN(n4624) );
  AND4_X1 U5619 ( .A1(n7106), .A2(n7105), .A3(n7104), .A4(n7103), .ZN(n7377)
         );
  AND4_X1 U5620 ( .A1(n6928), .A2(n6927), .A3(n6926), .A4(n6925), .ZN(n7293)
         );
  NOR2_X1 U5621 ( .A1(n7123), .A2(n4626), .ZN(n7299) );
  AND2_X1 U5622 ( .A1(n7876), .A2(n7875), .ZN(n7978) );
  NOR2_X1 U5623 ( .A1(n7123), .A2(n4625), .ZN(n7188) );
  INV_X1 U5624 ( .A(n4627), .ZN(n4625) );
  AND4_X1 U5625 ( .A1(n6904), .A2(n6903), .A3(n6902), .A4(n6901), .ZN(n7186)
         );
  NAND2_X1 U5626 ( .A1(n6101), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6798) );
  INV_X1 U5627 ( .A(n6787), .ZN(n6101) );
  OR2_X1 U5628 ( .A1(n6043), .A2(n6042), .ZN(n6787) );
  AND4_X1 U5629 ( .A1(n6803), .A2(n6802), .A3(n6801), .A4(n6800), .ZN(n7161)
         );
  NAND2_X1 U5630 ( .A1(n4527), .A2(n4835), .ZN(n4532) );
  NAND2_X1 U5631 ( .A1(n4838), .A2(n7853), .ZN(n6980) );
  AND4_X1 U5632 ( .A1(n6792), .A2(n6791), .A3(n6790), .A4(n6789), .ZN(n7117)
         );
  AND2_X1 U5633 ( .A1(n6989), .A2(n6993), .ZN(n6991) );
  AND2_X1 U5634 ( .A1(n6731), .A2(n4536), .ZN(n6989) );
  INV_X1 U5635 ( .A(n4976), .ZN(n4975) );
  OAI21_X1 U5636 ( .B1(n7836), .B2(n6554), .A(n6556), .ZN(n4976) );
  NOR2_X1 U5637 ( .A1(n9757), .A2(n8020), .ZN(n6573) );
  INV_X1 U5638 ( .A(n9748), .ZN(n8529) );
  INV_X1 U5639 ( .A(n9758), .ZN(n6504) );
  AND2_X1 U5640 ( .A1(n6485), .A2(n8385), .ZN(n6978) );
  AND2_X1 U5641 ( .A1(n9773), .A2(n6014), .ZN(n6552) );
  OR2_X1 U5642 ( .A1(n6140), .A2(n8003), .ZN(n6551) );
  NAND2_X1 U5643 ( .A1(n7790), .A2(n7789), .ZN(n8587) );
  NAND2_X1 U5644 ( .A1(n7765), .A2(n7764), .ZN(n8599) );
  AND2_X1 U5645 ( .A1(n8418), .A2(n8417), .ZN(n8605) );
  AND2_X1 U5646 ( .A1(n9780), .A2(n7992), .ZN(n9816) );
  AND2_X1 U5647 ( .A1(n9780), .A2(n6051), .ZN(n9815) );
  AND3_X1 U5648 ( .A1(n5945), .A2(n5944), .A3(n5943), .ZN(n9803) );
  INV_X1 U5649 ( .A(n9815), .ZN(n9831) );
  NOR2_X1 U5650 ( .A1(n6550), .A2(n6549), .ZN(n6568) );
  OAI21_X2 U5651 ( .B1(n5857), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5856) );
  INV_X1 U5652 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5855) );
  INV_X1 U5653 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5866) );
  INV_X1 U5654 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5989) );
  INV_X1 U5655 ( .A(n4589), .ZN(n4587) );
  NAND2_X1 U5656 ( .A1(n7261), .A2(n4589), .ZN(n4586) );
  NAND2_X1 U5657 ( .A1(n4588), .A2(n7249), .ZN(n5502) );
  NAND2_X1 U5658 ( .A1(n7258), .A2(n4589), .ZN(n4588) );
  INV_X1 U5659 ( .A(n5633), .ZN(n5615) );
  NAND2_X1 U5660 ( .A1(n4793), .A2(n4798), .ZN(n4792) );
  INV_X1 U5661 ( .A(n4795), .ZN(n4793) );
  NAND2_X1 U5662 ( .A1(n4486), .A2(n4798), .ZN(n4794) );
  AND2_X1 U5663 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5292) );
  NAND2_X1 U5664 ( .A1(n4770), .A2(n8737), .ZN(n4769) );
  AND2_X1 U5665 ( .A1(n8824), .A2(n4772), .ZN(n4771) );
  INV_X1 U5666 ( .A(n6477), .ZN(n5217) );
  NAND2_X1 U5667 ( .A1(n4599), .A2(n4598), .ZN(n4601) );
  INV_X1 U5668 ( .A(n5585), .ZN(n4599) );
  INV_X1 U5669 ( .A(n9206), .ZN(n8953) );
  NOR2_X1 U5670 ( .A1(n5490), .A2(n5489), .ZN(n5511) );
  AND2_X1 U5671 ( .A1(n7514), .A2(n7612), .ZN(n7608) );
  OR4_X1 U5672 ( .A1(n7617), .A2(n7662), .A3(n7657), .A4(n7513), .ZN(n7514) );
  INV_X1 U5673 ( .A(n7421), .ZN(n5697) );
  OR2_X1 U5674 ( .A1(n9544), .A2(n6287), .ZN(n9562) );
  OR2_X1 U5675 ( .A1(n5394), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5395) );
  AOI21_X1 U5676 ( .B1(n6397), .B2(n6396), .A(n6395), .ZN(n9622) );
  AND2_X1 U5677 ( .A1(n9622), .A2(n9621), .ZN(n9619) );
  NOR2_X1 U5678 ( .A1(n8906), .A2(n9634), .ZN(n9648) );
  AOI21_X1 U5679 ( .B1(n8910), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9659), .ZN(
        n8911) );
  NOR2_X1 U5680 ( .A1(n9022), .A2(n9282), .ZN(n9001) );
  NOR2_X1 U5681 ( .A1(n9038), .A2(n4850), .ZN(n4845) );
  NOR2_X1 U5682 ( .A1(n9084), .A2(n4650), .ZN(n9054) );
  INV_X1 U5683 ( .A(n4652), .ZN(n4650) );
  NOR2_X1 U5684 ( .A1(n9084), .A2(n9302), .ZN(n9066) );
  INV_X1 U5685 ( .A(n4604), .ZN(n4602) );
  INV_X1 U5686 ( .A(n5646), .ZN(n5164) );
  NAND2_X1 U5687 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n5164), .ZN(n5672) );
  NAND2_X1 U5688 ( .A1(n7588), .A2(n8987), .ZN(n9081) );
  NOR2_X1 U5689 ( .A1(n5615), .A2(n8769), .ZN(n5647) );
  AND2_X1 U5690 ( .A1(n9170), .A2(n4636), .ZN(n9111) );
  AND2_X1 U5691 ( .A1(n9112), .A2(n4412), .ZN(n4636) );
  NAND2_X1 U5692 ( .A1(n5593), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U5693 ( .A1(n9170), .A2(n9158), .ZN(n9152) );
  AND2_X1 U5694 ( .A1(n7573), .A2(n8980), .ZN(n9161) );
  NAND2_X1 U5695 ( .A1(n4687), .A2(n4688), .ZN(n9178) );
  NAND2_X1 U5696 ( .A1(n9228), .A2(n4689), .ZN(n4687) );
  AND4_X1 U5697 ( .A1(n5578), .A2(n5577), .A3(n5576), .A4(n5575), .ZN(n9200)
         );
  NAND2_X1 U5698 ( .A1(n9260), .A2(n4645), .ZN(n9187) );
  AND2_X1 U5699 ( .A1(n4418), .A2(n9189), .ZN(n4645) );
  NAND2_X1 U5700 ( .A1(n9260), .A2(n4418), .ZN(n9216) );
  OR2_X1 U5701 ( .A1(n5533), .A2(n5532), .ZN(n5551) );
  AND2_X1 U5702 ( .A1(n4693), .A2(n4691), .ZN(n9205) );
  AND2_X1 U5703 ( .A1(n4693), .A2(n8974), .ZN(n9203) );
  AND2_X1 U5704 ( .A1(n9260), .A2(n9494), .ZN(n9258) );
  NOR2_X1 U5705 ( .A1(n7153), .A2(n4642), .ZN(n9458) );
  INV_X1 U5706 ( .A(n4644), .ZN(n4642) );
  AND4_X1 U5707 ( .A1(n5452), .A2(n5451), .A3(n5450), .A4(n5449), .ZN(n9468)
         );
  NAND2_X1 U5708 ( .A1(n7143), .A2(n4716), .ZN(n7278) );
  NOR2_X1 U5709 ( .A1(n5371), .A2(n5370), .ZN(n5398) );
  AND4_X1 U5710 ( .A1(n5404), .A2(n5403), .A3(n5402), .A4(n5401), .ZN(n9466)
         );
  AND2_X1 U5711 ( .A1(n7143), .A2(n7539), .ZN(n7235) );
  INV_X1 U5712 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5349) );
  AND2_X1 U5713 ( .A1(n7537), .A2(n7539), .ZN(n7149) );
  AND4_X1 U5714 ( .A1(n5339), .A2(n5338), .A3(n5337), .A4(n5336), .ZN(n7049)
         );
  NAND2_X1 U5715 ( .A1(n7083), .A2(n7447), .ZN(n7528) );
  NAND2_X1 U5716 ( .A1(n4640), .A2(n7681), .ZN(n7078) );
  INV_X1 U5717 ( .A(n6756), .ZN(n4640) );
  AND4_X1 U5718 ( .A1(n5312), .A2(n5311), .A3(n5310), .A4(n5309), .ZN(n6943)
         );
  NAND2_X1 U5719 ( .A1(n6829), .A2(n9681), .ZN(n6828) );
  OR2_X1 U5720 ( .A1(n6828), .A2(n6812), .ZN(n6756) );
  NAND2_X1 U5721 ( .A1(n7446), .A2(n6823), .ZN(n6822) );
  NOR2_X1 U5722 ( .A1(n6687), .A2(n5237), .ZN(n6829) );
  NOR2_X1 U5723 ( .A1(n4404), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n4991) );
  NOR2_X1 U5724 ( .A1(n5171), .A2(n8929), .ZN(n6696) );
  OR2_X1 U5725 ( .A1(n6623), .A2(n5171), .ZN(n6721) );
  NAND2_X1 U5726 ( .A1(n7417), .A2(n7416), .ZN(n9275) );
  AOI211_X1 U5727 ( .C1(n9022), .C2(n9282), .A(n9723), .B(n9001), .ZN(n9281)
         );
  NAND2_X1 U5728 ( .A1(n9282), .A2(n9709), .ZN(n4711) );
  NAND2_X1 U5729 ( .A1(n5795), .A2(n5794), .ZN(n9285) );
  INV_X1 U5730 ( .A(n6952), .ZN(n9706) );
  NAND2_X2 U5731 ( .A1(n6673), .A2(n5737), .ZN(n9709) );
  AND2_X1 U5732 ( .A1(n5774), .A2(n6671), .ZN(n6336) );
  OAI21_X1 U5733 ( .B1(n9677), .B2(P1_D_REG_0__SCAN_IN), .A(n5759), .ZN(n6948)
         );
  XNOR2_X1 U5734 ( .A(n7477), .B(n7476), .ZN(n8681) );
  AND2_X1 U5735 ( .A1(n4887), .A2(n4719), .ZN(n4718) );
  INV_X1 U5736 ( .A(n4888), .ZN(n4886) );
  XNOR2_X1 U5737 ( .A(n5687), .B(n5686), .ZN(n7763) );
  OAI21_X1 U5738 ( .B1(n5629), .B2(n5628), .A(n5110), .ZN(n4917) );
  AND2_X1 U5739 ( .A1(n5116), .A2(n5115), .ZN(n5642) );
  NAND2_X1 U5740 ( .A1(n5150), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U5741 ( .A1(n5135), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n5136) );
  NAND2_X1 U5742 ( .A1(n5031), .A2(n5030), .ZN(n5342) );
  OAI21_X1 U5743 ( .B1(n5020), .B2(n4657), .A(n4656), .ZN(n5282) );
  AND3_X1 U5744 ( .A1(n5229), .A2(n5275), .A3(n5118), .ZN(n5279) );
  NAND2_X1 U5745 ( .A1(n5016), .A2(n5010), .ZN(n5206) );
  AND2_X1 U5746 ( .A1(n7805), .A2(n7804), .ZN(n8368) );
  AND4_X1 U5747 ( .A1(n7036), .A2(n7035), .A3(n7034), .A4(n7033), .ZN(n7326)
         );
  NAND2_X1 U5748 ( .A1(n4750), .A2(n7222), .ZN(n7223) );
  AND2_X1 U5749 ( .A1(n6893), .A2(n6892), .ZN(n6894) );
  NAND2_X1 U5750 ( .A1(n4738), .A2(n4736), .ZN(n8152) );
  INV_X1 U5751 ( .A(n4739), .ZN(n4736) );
  NAND2_X1 U5752 ( .A1(n7716), .A2(n7715), .ZN(n8631) );
  AND3_X1 U5753 ( .A1(n7729), .A2(n7728), .A3(n7727), .ZN(n8461) );
  NAND2_X1 U5754 ( .A1(n7018), .A2(n7017), .ZN(n7285) );
  NAND2_X1 U5755 ( .A1(n8206), .A2(n5951), .ZN(n8205) );
  XNOR2_X1 U5756 ( .A(n8100), .B(n8098), .ZN(n8196) );
  NAND2_X1 U5757 ( .A1(n4734), .A2(n8066), .ZN(n4733) );
  INV_X1 U5758 ( .A(n4737), .ZN(n4734) );
  AOI21_X1 U5759 ( .B1(n8443), .B2(n7780), .A(n7739), .ZN(n8462) );
  INV_X1 U5760 ( .A(n4755), .ZN(n4754) );
  AOI21_X1 U5761 ( .B1(n4755), .B2(n4753), .A(n4752), .ZN(n4751) );
  NAND2_X1 U5762 ( .A1(n6913), .A2(n6912), .ZN(n7196) );
  AOI21_X1 U5763 ( .B1(n8188), .B2(n8187), .A(n8061), .ZN(n8228) );
  NAND2_X1 U5764 ( .A1(n7705), .A2(n7704), .ZN(n8634) );
  CLKBUF_X1 U5765 ( .A(n6348), .Z(n6425) );
  OR2_X1 U5766 ( .A1(n8263), .A2(n5905), .ZN(n8255) );
  NAND2_X1 U5767 ( .A1(n6034), .A2(n8556), .ZN(n8259) );
  NAND2_X1 U5768 ( .A1(n7370), .A2(n7369), .ZN(n8260) );
  INV_X1 U5769 ( .A(n8368), .ZN(n8266) );
  AOI21_X1 U5770 ( .B1(n8361), .B2(n7780), .A(n6449), .ZN(n8240) );
  NOR2_X1 U5771 ( .A1(n6141), .A2(n6083), .ZN(n8264) );
  INV_X1 U5772 ( .A(n8264), .ZN(n8271) );
  OR2_X1 U5773 ( .A1(n7802), .A2(n5897), .ZN(n5898) );
  OR2_X1 U5774 ( .A1(n6302), .A2(n4569), .ZN(n6241) );
  NAND2_X1 U5775 ( .A1(n6241), .A2(n6242), .ZN(n6240) );
  AOI21_X1 U5776 ( .B1(n4569), .B2(n6242), .A(n4467), .ZN(n4568) );
  NAND2_X1 U5777 ( .A1(n6216), .A2(n4483), .ZN(n6190) );
  NAND2_X1 U5778 ( .A1(n6190), .A2(n6191), .ZN(n6189) );
  NAND2_X1 U5779 ( .A1(n6177), .A2(n6178), .ZN(n6357) );
  NOR2_X1 U5780 ( .A1(n9892), .A2(n4566), .ZN(n6412) );
  AND2_X1 U5781 ( .A1(n6882), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4566) );
  NAND2_X1 U5782 ( .A1(n6412), .A2(n6413), .ZN(n6528) );
  AND2_X1 U5783 ( .A1(n6528), .A2(n4565), .ZN(n6530) );
  NAND2_X1 U5784 ( .A1(n6529), .A2(n6900), .ZN(n4565) );
  XNOR2_X1 U5785 ( .A(n7313), .B(n7368), .ZN(n7133) );
  INV_X1 U5786 ( .A(n4573), .ZN(n8307) );
  INV_X1 U5787 ( .A(n4571), .ZN(n8318) );
  OAI21_X1 U5788 ( .B1(n8406), .B2(n4943), .A(n4940), .ZN(n8359) );
  NAND2_X1 U5789 ( .A1(n4945), .A2(n4946), .ZN(n8374) );
  NAND2_X1 U5790 ( .A1(n8406), .A2(n4948), .ZN(n4945) );
  INV_X1 U5791 ( .A(n8599), .ZN(n8394) );
  NAND2_X1 U5792 ( .A1(n8406), .A2(n4953), .ZN(n8390) );
  NAND2_X1 U5793 ( .A1(n4967), .A2(n4968), .ZN(n8435) );
  AND2_X1 U5794 ( .A1(n8452), .A2(n8451), .ZN(n8616) );
  NAND2_X1 U5795 ( .A1(n4834), .A2(n4833), .ZN(n8446) );
  NAND2_X1 U5796 ( .A1(n8471), .A2(n8466), .ZN(n8442) );
  AOI21_X1 U5797 ( .B1(n8456), .B2(n8031), .A(n4414), .ZN(n8439) );
  NAND2_X1 U5798 ( .A1(n4983), .A2(n4415), .ZN(n8523) );
  AND2_X1 U5799 ( .A1(n4983), .A2(n4982), .ZN(n8524) );
  NAND2_X1 U5800 ( .A1(n7211), .A2(n7210), .ZN(n7365) );
  NAND2_X1 U5801 ( .A1(n7339), .A2(n7338), .ZN(n7364) );
  AND2_X1 U5802 ( .A1(n7114), .A2(n7113), .ZN(n7115) );
  NAND2_X1 U5803 ( .A1(n6884), .A2(n6883), .ZN(n7162) );
  AND2_X1 U5804 ( .A1(n6977), .A2(n6957), .ZN(n6958) );
  NAND2_X1 U5805 ( .A1(n6729), .A2(n7851), .ZN(n6960) );
  AND2_X1 U5806 ( .A1(n7204), .A2(n9816), .ZN(n8521) );
  OR2_X1 U5807 ( .A1(n6646), .A2(n6645), .ZN(n4957) );
  NAND2_X1 U5808 ( .A1(n6555), .A2(n6554), .ZN(n6572) );
  INV_X1 U5809 ( .A(n8538), .ZN(n8566) );
  CLKBUF_X1 U5810 ( .A(n8518), .Z(n8535) );
  NAND2_X1 U5811 ( .A1(n9771), .A2(n9770), .ZN(n9775) );
  INV_X1 U5812 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8676) );
  NAND2_X1 U5813 ( .A1(n5876), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5871) );
  INV_X1 U5814 ( .A(n6015), .ZN(n7387) );
  INV_X1 U5815 ( .A(n6016), .ZN(n7342) );
  XNOR2_X1 U5816 ( .A(n5843), .B(n5842), .ZN(n7230) );
  INV_X1 U5817 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7067) );
  INV_X1 U5818 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5858) );
  INV_X1 U5819 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10070) );
  INV_X1 U5820 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6857) );
  INV_X1 U5821 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6501) );
  INV_X1 U5822 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6445) );
  INV_X1 U5823 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6440) );
  INV_X1 U5824 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6229) );
  INV_X1 U5825 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9970) );
  INV_X1 U5826 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10117) );
  INV_X1 U5827 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6078) );
  INV_X1 U5828 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10158) );
  INV_X1 U5829 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9981) );
  INV_X1 U5830 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10104) );
  INV_X1 U5831 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U5832 ( .A1(n4574), .A2(n5879), .ZN(n6164) );
  INV_X1 U5833 ( .A(n4575), .ZN(n4574) );
  OAI22_X1 U5834 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .B1(
        n5992), .B2(n4576), .ZN(n4575) );
  AND4_X1 U5835 ( .A1(n5356), .A2(n5355), .A3(n5354), .A4(n5353), .ZN(n7145)
         );
  NAND2_X1 U5836 ( .A1(n5645), .A2(n5644), .ZN(n9310) );
  NAND2_X1 U5837 ( .A1(n5247), .A2(n5246), .ZN(n6597) );
  NAND2_X1 U5838 ( .A1(n5348), .A2(n4434), .ZN(n5008) );
  NAND2_X1 U5839 ( .A1(n4790), .A2(n4792), .ZN(n8723) );
  OR2_X1 U5840 ( .A1(n8707), .A2(n4794), .ZN(n4790) );
  NAND2_X1 U5841 ( .A1(n5444), .A2(n5443), .ZN(n9508) );
  AND4_X1 U5842 ( .A1(n5517), .A2(n5516), .A3(n5515), .A4(n5514), .ZN(n9208)
         );
  NAND2_X1 U5843 ( .A1(n8828), .A2(n8824), .ZN(n8739) );
  NAND2_X1 U5844 ( .A1(n5544), .A2(n4769), .ZN(n8745) );
  NAND2_X1 U5845 ( .A1(n4779), .A2(n4782), .ZN(n8751) );
  NAND2_X1 U5846 ( .A1(n4786), .A2(n4784), .ZN(n4779) );
  INV_X1 U5847 ( .A(n6604), .ZN(n5287) );
  NAND2_X1 U5848 ( .A1(n4760), .A2(n4759), .ZN(n7059) );
  NAND2_X1 U5849 ( .A1(n4764), .A2(n4766), .ZN(n4759) );
  OR2_X1 U5850 ( .A1(n8707), .A2(n4797), .ZN(n4791) );
  AOI21_X1 U5851 ( .B1(n8707), .B2(n8705), .A(n4797), .ZN(n8759) );
  NAND2_X1 U5852 ( .A1(n5176), .A2(n5175), .ZN(n9325) );
  NAND2_X1 U5853 ( .A1(n7258), .A2(n5462), .ZN(n7252) );
  NAND2_X1 U5854 ( .A1(n5468), .A2(n5467), .ZN(n9499) );
  NAND2_X1 U5855 ( .A1(n5418), .A2(n5417), .ZN(n8783) );
  NAND2_X1 U5856 ( .A1(n5572), .A2(n5571), .ZN(n9335) );
  INV_X1 U5857 ( .A(n8825), .ZN(n8812) );
  INV_X1 U5858 ( .A(n8806), .ZN(n8831) );
  OR2_X1 U5859 ( .A1(n5597), .A2(n5596), .ZN(n9181) );
  INV_X1 U5860 ( .A(n9200), .ZN(n9162) );
  INV_X1 U5861 ( .A(n9468), .ZN(n8838) );
  NAND2_X1 U5862 ( .A1(n7418), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5190) );
  OR2_X1 U5863 ( .A1(n5178), .A2(n5201), .ZN(n5204) );
  NAND2_X1 U5864 ( .A1(n6460), .A2(n6461), .ZN(n6459) );
  INV_X1 U5865 ( .A(n9275), .ZN(n8942) );
  OAI21_X1 U5866 ( .B1(n4713), .B2(n9234), .A(n9000), .ZN(n9280) );
  XNOR2_X1 U5867 ( .A(n8997), .B(n8996), .ZN(n4713) );
  NAND2_X1 U5868 ( .A1(n4695), .A2(n4696), .ZN(n9012) );
  AND2_X1 U5869 ( .A1(n4701), .A2(n4700), .ZN(n9041) );
  INV_X1 U5870 ( .A(n9291), .ZN(n9036) );
  NAND2_X1 U5871 ( .A1(n4846), .A2(n4849), .ZN(n9031) );
  NAND2_X1 U5872 ( .A1(n9063), .A2(n8963), .ZN(n9048) );
  NAND2_X1 U5873 ( .A1(n5129), .A2(n5128), .ZN(n9307) );
  NAND2_X1 U5874 ( .A1(n4706), .A2(n4416), .ZN(n9102) );
  INV_X1 U5875 ( .A(n9310), .ZN(n9100) );
  NAND2_X1 U5876 ( .A1(n4854), .A2(n4858), .ZN(n9093) );
  NAND2_X1 U5877 ( .A1(n4856), .A2(n4855), .ZN(n4854) );
  NOR2_X1 U5878 ( .A1(n9125), .A2(n8983), .ZN(n9118) );
  NAND2_X1 U5879 ( .A1(n9124), .A2(n9127), .ZN(n4857) );
  OAI21_X1 U5880 ( .B1(n9213), .B2(n4873), .A(n4872), .ZN(n9169) );
  NOR2_X1 U5881 ( .A1(n9211), .A2(n4877), .ZN(n9186) );
  NAND2_X1 U5882 ( .A1(n5382), .A2(n5381), .ZN(n7233) );
  OAI21_X1 U5883 ( .B1(n7148), .B2(n7149), .A(n7150), .ZN(n7234) );
  INV_X1 U5884 ( .A(n9271), .ZN(n9214) );
  NAND2_X1 U5885 ( .A1(n6744), .A2(n6717), .ZN(n6719) );
  AND2_X1 U5886 ( .A1(n9193), .A2(n9711), .ZN(n9461) );
  INV_X1 U5887 ( .A(n9475), .ZN(n9264) );
  NAND2_X1 U5888 ( .A1(n9269), .A2(n6674), .ZN(n9475) );
  INV_X1 U5889 ( .A(n9737), .ZN(n9735) );
  INV_X1 U5890 ( .A(n9729), .ZN(n9727) );
  AND2_X1 U5891 ( .A1(n5776), .A2(n5741), .ZN(n9678) );
  XNOR2_X1 U5892 ( .A(n7431), .B(n7430), .ZN(n9363) );
  NAND2_X1 U5893 ( .A1(n7427), .A2(n7426), .ZN(n7431) );
  INV_X1 U5894 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7179) );
  NAND2_X1 U5895 ( .A1(n5643), .A2(n4916), .ZN(n7740) );
  OR2_X1 U5896 ( .A1(n4917), .A2(n5642), .ZN(n4916) );
  NOR2_X1 U5897 ( .A1(n5880), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7176) );
  INV_X1 U5898 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7129) );
  CLKBUF_X1 U5899 ( .A(n5736), .Z(n7612) );
  NAND2_X1 U5900 ( .A1(n4804), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5138) );
  NOR2_X1 U5901 ( .A1(n4604), .A2(n4606), .ZN(n4603) );
  INV_X1 U5902 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10058) );
  INV_X1 U5903 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U5904 ( .A1(n5486), .A2(n5131), .ZN(n5528) );
  INV_X1 U5905 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10060) );
  INV_X1 U5906 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10026) );
  INV_X1 U5907 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6132) );
  INV_X1 U5908 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6114) );
  INV_X1 U5909 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6099) );
  INV_X1 U5910 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6080) );
  OR2_X1 U5911 ( .A1(n5365), .A2(n5364), .ZN(n9587) );
  INV_X1 U5912 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6074) );
  INV_X1 U5913 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6064) );
  XNOR2_X1 U5914 ( .A(n5317), .B(n5316), .ZN(n6070) );
  INV_X1 U5915 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5314) );
  INV_X1 U5916 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9979) );
  NAND2_X1 U5917 ( .A1(n4906), .A2(n5025), .ZN(n5299) );
  INV_X1 U5918 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U5919 ( .A1(n5020), .A2(n5019), .ZN(n5257) );
  NOR2_X1 U5920 ( .A1(n9434), .A2(n10209), .ZN(n9881) );
  AOI21_X1 U5921 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9879), .ZN(n9878) );
  NOR2_X1 U5922 ( .A1(n9878), .A2(n9877), .ZN(n9876) );
  NAND2_X1 U5923 ( .A1(n4725), .A2(n4478), .ZN(n4724) );
  OAI21_X1 U5924 ( .B1(n4680), .B2(n4679), .A(n8008), .ZN(P2_U3244) );
  NOR2_X1 U5925 ( .A1(n4811), .A2(n4490), .ZN(n4679) );
  OAI21_X1 U5926 ( .B1(n4811), .B2(n4810), .A(n8002), .ZN(n4680) );
  INV_X1 U5927 ( .A(n8046), .ZN(n4533) );
  OR2_X1 U5928 ( .A1(n9853), .A2(n4973), .ZN(n4972) );
  NAND2_X1 U5929 ( .A1(n8659), .A2(n9853), .ZN(n4974) );
  INV_X1 U5930 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n4973) );
  NAND2_X1 U5931 ( .A1(n9839), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4607) );
  NAND2_X1 U5932 ( .A1(n8659), .A2(n4405), .ZN(n4608) );
  NOR2_X1 U5933 ( .A1(n4989), .A2(n5007), .ZN(n5787) );
  NAND2_X1 U5934 ( .A1(n5824), .A2(n4578), .ZN(P1_U3218) );
  NAND2_X1 U5935 ( .A1(n4580), .A2(n4579), .ZN(n4578) );
  NOR2_X1 U5936 ( .A1(n5806), .A2(n8825), .ZN(n4579) );
  NAND2_X1 U5937 ( .A1(n7667), .A2(n4436), .ZN(n4507) );
  INV_X1 U5938 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8934) );
  AND2_X1 U5939 ( .A1(n7970), .A2(n7853), .ZN(n4410) );
  AND2_X1 U5940 ( .A1(n4858), .A2(n4853), .ZN(n4411) );
  AND2_X1 U5941 ( .A1(n4638), .A2(n4637), .ZN(n4412) );
  INV_X1 U5942 ( .A(n8582), .ZN(n8350) );
  OR2_X1 U5943 ( .A1(n4597), .A2(n8791), .ZN(n4413) );
  OR2_X1 U5944 ( .A1(n9242), .A2(n9208), .ZN(n8974) );
  INV_X1 U5945 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5992) );
  AND2_X1 U5946 ( .A1(n8466), .A2(n8482), .ZN(n4414) );
  INV_X1 U5947 ( .A(n4486), .ZN(n4797) );
  AND2_X1 U5948 ( .A1(n8526), .A2(n4982), .ZN(n4415) );
  INV_X1 U5949 ( .A(n8032), .ZN(n4947) );
  AND2_X1 U5950 ( .A1(n8984), .A2(n7584), .ZN(n4416) );
  OR2_X1 U5951 ( .A1(n9291), .A2(n9053), .ZN(n8992) );
  OR2_X1 U5952 ( .A1(n7365), .A2(n7377), .ZN(n7887) );
  AND2_X1 U5953 ( .A1(n4466), .A2(n4586), .ZN(n4417) );
  AND2_X1 U5954 ( .A1(n4647), .A2(n4646), .ZN(n4418) );
  INV_X1 U5955 ( .A(n8033), .ZN(n4938) );
  AND2_X1 U5956 ( .A1(n7666), .A2(n7013), .ZN(n4419) );
  XNOR2_X1 U5957 ( .A(n5021), .B(n4521), .ZN(n5258) );
  AND2_X1 U5958 ( .A1(n7806), .A2(n7940), .ZN(n8034) );
  AND2_X1 U5959 ( .A1(n7903), .A2(n4445), .ZN(n4420) );
  AND2_X1 U5960 ( .A1(n4786), .A2(n5654), .ZN(n4421) );
  AND2_X1 U5961 ( .A1(n7958), .A2(n7956), .ZN(n4422) );
  NAND2_X1 U5962 ( .A1(n5510), .A2(n5509), .ZN(n9242) );
  AND4_X1 U5963 ( .A1(n6006), .A2(n6005), .A3(n6004), .A4(n6003), .ZN(n6983)
         );
  INV_X1 U5964 ( .A(n6983), .ZN(n4535) );
  AND2_X1 U5965 ( .A1(n7683), .A2(n7682), .ZN(n8577) );
  NAND2_X1 U5966 ( .A1(n9265), .A2(n9229), .ZN(n4423) );
  AND2_X1 U5967 ( .A1(n8992), .A2(n7488), .ZN(n9038) );
  INV_X1 U5968 ( .A(n4860), .ZN(n4855) );
  OR2_X1 U5969 ( .A1(n8960), .A2(n4861), .ZN(n4860) );
  OR2_X1 U5970 ( .A1(n8033), .A2(n4439), .ZN(n4424) );
  AND2_X1 U5971 ( .A1(n7945), .A2(n7841), .ZN(n4425) );
  AND2_X1 U5972 ( .A1(n8057), .A2(n8056), .ZN(n4426) );
  INV_X1 U5973 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5837) );
  OR2_X1 U5974 ( .A1(n9081), .A2(n9103), .ZN(n4427) );
  NAND2_X1 U5975 ( .A1(n5745), .A2(n5149), .ZN(n5776) );
  NAND2_X1 U5976 ( .A1(n4788), .A2(n5584), .ZN(n4428) );
  AND2_X1 U5977 ( .A1(n4613), .A2(n4612), .ZN(n4429) );
  AND2_X1 U5978 ( .A1(n6704), .A2(n6717), .ZN(n4430) );
  AND2_X1 U5979 ( .A1(n4534), .A2(n4533), .ZN(n4431) );
  AND2_X1 U5980 ( .A1(n5631), .A2(n5630), .ZN(n9112) );
  INV_X1 U5981 ( .A(n9112), .ZN(n9317) );
  NAND2_X1 U5982 ( .A1(n7611), .A2(n8929), .ZN(n4432) );
  AND2_X1 U5983 ( .A1(n7786), .A2(n7785), .ZN(n8367) );
  NAND2_X1 U5984 ( .A1(n4677), .A2(n4675), .ZN(n6643) );
  INV_X1 U5985 ( .A(n6643), .ZN(n6587) );
  OR2_X1 U5986 ( .A1(n7153), .A2(n4643), .ZN(n4433) );
  INV_X1 U5987 ( .A(n5369), .ZN(n4766) );
  NAND2_X1 U5988 ( .A1(n9373), .A2(n5163), .ZN(n5178) );
  AND2_X1 U5989 ( .A1(n4766), .A2(n6873), .ZN(n4434) );
  AND2_X1 U5990 ( .A1(n7887), .A2(n7886), .ZN(n7980) );
  NAND2_X1 U5991 ( .A1(n4944), .A2(n4946), .ZN(n4943) );
  INV_X1 U5992 ( .A(n8434), .ZN(n4966) );
  AND2_X1 U5993 ( .A1(n4538), .A2(n4537), .ZN(n4435) );
  OR2_X1 U5994 ( .A1(n4510), .A2(n4508), .ZN(n4436) );
  INV_X1 U5995 ( .A(n4717), .ZN(n4716) );
  NAND2_X1 U5996 ( .A1(n7539), .A2(n7538), .ZN(n4717) );
  AND2_X1 U5997 ( .A1(n4857), .A2(n8959), .ZN(n4437) );
  AND2_X1 U5998 ( .A1(n4938), .A2(n8364), .ZN(n4438) );
  AND3_X1 U5999 ( .A1(n5933), .A2(n5932), .A3(n5931), .ZN(n9796) );
  INV_X1 U6000 ( .A(n9796), .ZN(n4812) );
  INV_X1 U6001 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n10008) );
  INV_X1 U6002 ( .A(n8765), .ZN(n4775) );
  AND2_X1 U6003 ( .A1(n7938), .A2(n7956), .ZN(n4439) );
  INV_X1 U6004 ( .A(n7836), .ZN(n7967) );
  NAND2_X1 U6005 ( .A1(n5590), .A2(n5589), .ZN(n9330) );
  NAND2_X1 U6006 ( .A1(n7754), .A2(n7753), .ZN(n8602) );
  NAND2_X1 U6007 ( .A1(n7595), .A2(n9039), .ZN(n9050) );
  INV_X1 U6008 ( .A(n9050), .ZN(n4699) );
  NAND2_X1 U6009 ( .A1(n5696), .A2(n5695), .ZN(n9297) );
  NOR2_X1 U6010 ( .A1(n7810), .A2(n10104), .ZN(n4440) );
  NOR2_X1 U6011 ( .A1(n7032), .A2(n6171), .ZN(n4441) );
  NOR3_X1 U6012 ( .A1(n9084), .A2(n9285), .A3(n4651), .ZN(n4648) );
  NAND2_X1 U6013 ( .A1(n5145), .A2(n4886), .ZN(n4442) );
  INV_X1 U6014 ( .A(n9130), .ZN(n9107) );
  AND4_X1 U6015 ( .A1(n5638), .A2(n5637), .A3(n5636), .A4(n5635), .ZN(n9130)
         );
  NOR2_X1 U6016 ( .A1(n7922), .A2(n7841), .ZN(n4443) );
  INV_X1 U6017 ( .A(n7979), .ZN(n4821) );
  AND2_X1 U6018 ( .A1(n7881), .A2(n7324), .ZN(n7979) );
  AND2_X1 U6019 ( .A1(n4955), .A2(n6726), .ZN(n4444) );
  OR2_X1 U6020 ( .A1(n9808), .A2(n8281), .ZN(n7851) );
  INV_X1 U6021 ( .A(n8619), .ZN(n8466) );
  NAND2_X1 U6022 ( .A1(n7732), .A2(n7731), .ZN(n8619) );
  NAND2_X1 U6023 ( .A1(n8391), .A2(n4615), .ZN(n4616) );
  INV_X1 U6024 ( .A(n5022), .ZN(n4658) );
  AND2_X1 U6025 ( .A1(n7889), .A2(n7888), .ZN(n4445) );
  AND2_X1 U6026 ( .A1(n7526), .A2(n7634), .ZN(n4446) );
  INV_X1 U6027 ( .A(n4649), .ZN(n9032) );
  NOR2_X1 U6028 ( .A1(n9084), .A2(n4651), .ZN(n4649) );
  AND2_X1 U6029 ( .A1(n9508), .A2(n8838), .ZN(n4447) );
  AND3_X1 U6030 ( .A1(n5236), .A2(n5235), .A3(n5234), .ZN(n6712) );
  INV_X1 U6031 ( .A(n4850), .ZN(n4849) );
  AND2_X1 U6032 ( .A1(n4902), .A2(n4898), .ZN(n4448) );
  NAND2_X1 U6033 ( .A1(n7777), .A2(n7776), .ZN(n8593) );
  INV_X1 U6034 ( .A(n8593), .ZN(n4950) );
  OR2_X1 U6035 ( .A1(n8613), .A2(n8462), .ZN(n7923) );
  INV_X1 U6036 ( .A(n7923), .ZN(n4831) );
  AND2_X1 U6037 ( .A1(n4791), .A2(n4795), .ZN(n4449) );
  AND2_X1 U6038 ( .A1(n7829), .A2(n7828), .ZN(n4450) );
  AND2_X1 U6039 ( .A1(n8025), .A2(n8551), .ZN(n4451) );
  AND2_X1 U6040 ( .A1(n8608), .A2(n8450), .ZN(n4452) );
  AND2_X1 U6041 ( .A1(n7604), .A2(n7603), .ZN(n4453) );
  AND2_X1 U6042 ( .A1(n7928), .A2(n7841), .ZN(n4454) );
  NAND2_X1 U6043 ( .A1(n7893), .A2(n8542), .ZN(n4455) );
  AND3_X1 U6044 ( .A1(n5928), .A2(n5926), .A3(n5927), .ZN(n4456) );
  AND2_X1 U6045 ( .A1(n8281), .A2(n6728), .ZN(n4457) );
  NOR2_X1 U6046 ( .A1(n9189), .A2(n8953), .ZN(n4458) );
  NOR2_X1 U6047 ( .A1(n5627), .A2(n5626), .ZN(n4459) );
  NOR2_X1 U6048 ( .A1(n8613), .A2(n8269), .ZN(n4460) );
  AND2_X1 U6049 ( .A1(n4634), .A2(n4633), .ZN(n5145) );
  INV_X1 U6050 ( .A(n4874), .ZN(n4873) );
  AOI21_X1 U6051 ( .B1(n9212), .B2(n4875), .A(n8954), .ZN(n4874) );
  AND2_X1 U6052 ( .A1(n5131), .A2(n4605), .ZN(n4461) );
  AND2_X1 U6053 ( .A1(n7865), .A2(n7861), .ZN(n6961) );
  AND2_X1 U6054 ( .A1(n4903), .A2(n7806), .ZN(n4462) );
  AND2_X1 U6055 ( .A1(n5027), .A2(SI_5_), .ZN(n4463) );
  NAND2_X1 U6056 ( .A1(n8363), .A2(n8240), .ZN(n4464) );
  OR2_X1 U6057 ( .A1(n8774), .A2(n5437), .ZN(n4465) );
  OAI21_X1 U6058 ( .B1(n4784), .B2(n4781), .A(n8752), .ZN(n4780) );
  AND2_X1 U6059 ( .A1(n4591), .A2(n7249), .ZN(n4466) );
  NOR2_X1 U6060 ( .A1(n6170), .A2(n6171), .ZN(n4467) );
  INV_X1 U6061 ( .A(n4765), .ZN(n4764) );
  OAI21_X1 U6062 ( .B1(n6873), .B2(n4766), .A(n8714), .ZN(n4765) );
  AND2_X1 U6063 ( .A1(n4950), .A2(n8367), .ZN(n4468) );
  AND2_X1 U6064 ( .A1(n7857), .A2(n7858), .ZN(n7970) );
  OR2_X1 U6065 ( .A1(n8579), .A2(n8124), .ZN(n7945) );
  INV_X1 U6066 ( .A(n4943), .ZN(n4942) );
  NAND2_X1 U6067 ( .A1(n7945), .A2(n7946), .ZN(n8036) );
  INV_X1 U6068 ( .A(n8036), .ZN(n4900) );
  INV_X1 U6069 ( .A(n4952), .ZN(n4951) );
  NAND2_X1 U6070 ( .A1(n8394), .A2(n8200), .ZN(n4952) );
  AND2_X1 U6071 ( .A1(n9310), .A2(n8837), .ZN(n4469) );
  AND2_X1 U6072 ( .A1(n4792), .A2(n4789), .ZN(n4788) );
  OR2_X1 U6073 ( .A1(n8582), .A2(n8368), .ZN(n7806) );
  XNOR2_X1 U6074 ( .A(n8608), .B(n8450), .ZN(n8434) );
  AND2_X1 U6075 ( .A1(n4509), .A2(n7670), .ZN(n4470) );
  OR2_X1 U6076 ( .A1(n7861), .A2(n7841), .ZN(n4471) );
  NOR2_X1 U6077 ( .A1(n4786), .A2(n5654), .ZN(n4472) );
  NAND2_X1 U6078 ( .A1(n8841), .A2(n7233), .ZN(n4473) );
  AND2_X1 U6079 ( .A1(n8066), .A2(n4741), .ZN(n4474) );
  NOR2_X1 U6080 ( .A1(n7974), .A2(n4531), .ZN(n4530) );
  INV_X1 U6081 ( .A(n9018), .ZN(n9011) );
  AND2_X1 U6082 ( .A1(n8993), .A2(n7516), .ZN(n9018) );
  INV_X1 U6083 ( .A(n4782), .ZN(n4781) );
  NAND2_X1 U6084 ( .A1(n5654), .A2(n4783), .ZN(n4782) );
  AND2_X1 U6085 ( .A1(n8034), .A2(n4438), .ZN(n4475) );
  INV_X1 U6086 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5126) );
  INV_X1 U6087 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4920) );
  INV_X2 U6088 ( .A(n7810), .ZN(n7703) );
  NAND2_X1 U6089 ( .A1(n5998), .A2(n5997), .ZN(n6955) );
  INV_X1 U6090 ( .A(n6955), .ZN(n4536) );
  AND2_X1 U6091 ( .A1(n8471), .A2(n4630), .ZN(n4476) );
  NAND2_X1 U6092 ( .A1(n7692), .A2(n7691), .ZN(n8641) );
  INV_X1 U6093 ( .A(n8791), .ZN(n4600) );
  NAND4_X1 U6094 ( .A1(n5835), .A2(n5834), .A3(n5941), .A4(n5836), .ZN(n5849)
         );
  INV_X1 U6095 ( .A(n8113), .ZN(n4731) );
  OR2_X1 U6096 ( .A1(n6205), .A2(n6586), .ZN(n4477) );
  NAND4_X1 U6097 ( .A1(n5229), .A2(n5275), .A3(n5118), .A4(n5119), .ZN(n5313)
         );
  INV_X1 U6098 ( .A(n5313), .ZN(n4878) );
  INV_X1 U6099 ( .A(n8976), .ZN(n4690) );
  NAND2_X1 U6100 ( .A1(n7290), .A2(n7875), .ZN(n7291) );
  NAND2_X1 U6101 ( .A1(n7689), .A2(n7688), .ZN(n8565) );
  OR2_X1 U6102 ( .A1(n8123), .A2(n4731), .ZN(n4478) );
  AND2_X1 U6103 ( .A1(n4813), .A2(n4817), .ZN(n4479) );
  AND2_X1 U6104 ( .A1(n8113), .A2(n8111), .ZN(n8132) );
  INV_X1 U6105 ( .A(n8132), .ZN(n4728) );
  NAND2_X1 U6106 ( .A1(n4878), .A2(n4992), .ZN(n5441) );
  OR2_X1 U6107 ( .A1(n8958), .A2(n9129), .ZN(n4480) );
  INV_X1 U6108 ( .A(n4618), .ZN(n8531) );
  NOR3_X1 U6109 ( .A1(n7378), .A2(n8641), .A3(n4621), .ZN(n4618) );
  NAND2_X1 U6110 ( .A1(n7808), .A2(n7807), .ZN(n8579) );
  INV_X1 U6111 ( .A(n8579), .ZN(n4612) );
  NOR2_X1 U6112 ( .A1(n7378), .A2(n4619), .ZN(n4622) );
  NAND2_X1 U6113 ( .A1(n5397), .A2(n5396), .ZN(n8700) );
  AND2_X1 U6114 ( .A1(n9101), .A2(n4499), .ZN(n4481) );
  NAND2_X1 U6115 ( .A1(n5488), .A2(n5487), .ZN(n9265) );
  AND2_X1 U6116 ( .A1(n8984), .A2(n7602), .ZN(n4482) );
  OR2_X1 U6117 ( .A1(n6221), .A2(n6172), .ZN(n4483) );
  NAND2_X1 U6118 ( .A1(n5550), .A2(n5549), .ZN(n9342) );
  AND2_X1 U6119 ( .A1(n7566), .A2(n9194), .ZN(n9212) );
  INV_X1 U6120 ( .A(n9212), .ZN(n4692) );
  NAND2_X1 U6121 ( .A1(n9170), .A2(n4412), .ZN(n4639) );
  NAND2_X1 U6122 ( .A1(n7098), .A2(n7097), .ZN(n7337) );
  AND2_X1 U6123 ( .A1(n4738), .A2(n4737), .ZN(n4484) );
  OR2_X1 U6124 ( .A1(n4598), .A2(n8791), .ZN(n4485) );
  NAND2_X1 U6125 ( .A1(n4967), .A2(n4964), .ZN(n4971) );
  INV_X1 U6126 ( .A(n8641), .ZN(n8025) );
  NAND2_X1 U6127 ( .A1(n6568), .A2(n6567), .ZN(n9839) );
  AND2_X1 U6128 ( .A1(n5170), .A2(n9087), .ZN(n7602) );
  INV_X1 U6129 ( .A(n7602), .ZN(n4499) );
  NAND2_X1 U6130 ( .A1(n6893), .A2(n4755), .ZN(n6917) );
  NAND2_X1 U6131 ( .A1(n5531), .A2(n5530), .ZN(n9220) );
  INV_X1 U6132 ( .A(n9220), .ZN(n4646) );
  INV_X1 U6133 ( .A(n5170), .ZN(n5738) );
  INV_X1 U6134 ( .A(n8518), .ZN(n9768) );
  AND2_X1 U6135 ( .A1(n6490), .A2(n8556), .ZN(n8518) );
  INV_X1 U6136 ( .A(n7013), .ZN(n7615) );
  XNOR2_X1 U6137 ( .A(n5138), .B(n5137), .ZN(n7013) );
  OR2_X1 U6138 ( .A1(n5604), .A2(n5603), .ZN(n4486) );
  NAND2_X1 U6139 ( .A1(n5613), .A2(n5612), .ZN(n9322) );
  INV_X1 U6140 ( .A(n9322), .ZN(n4637) );
  AOI21_X1 U6141 ( .B1(n6576), .B2(n7836), .A(n6561), .ZN(n6613) );
  OR2_X1 U6142 ( .A1(n7123), .A2(n7162), .ZN(n4487) );
  NAND2_X1 U6143 ( .A1(n4532), .A2(n6961), .ZN(n7116) );
  NOR3_X1 U6144 ( .A1(n7153), .A2(n9508), .A3(n4643), .ZN(n4641) );
  NAND2_X1 U6145 ( .A1(n4720), .A2(n4878), .ZN(n5739) );
  AND2_X1 U6146 ( .A1(n4750), .A2(n4748), .ZN(n4488) );
  INV_X1 U6147 ( .A(n6729), .ZN(n4525) );
  INV_X1 U6148 ( .A(n8282), .ZN(n4678) );
  NAND2_X1 U6149 ( .A1(n7843), .A2(n7959), .ZN(n9747) );
  OR2_X1 U6150 ( .A1(n8335), .A2(n7994), .ZN(n4489) );
  INV_X1 U6151 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4719) );
  NAND2_X1 U6152 ( .A1(n7829), .A2(n7823), .ZN(n7966) );
  NAND2_X1 U6153 ( .A1(n8092), .A2(n7817), .ZN(n4490) );
  XNOR2_X1 U6154 ( .A(n5867), .B(n5866), .ZN(n7992) );
  AND2_X1 U6155 ( .A1(n8205), .A2(n5955), .ZN(n4491) );
  XNOR2_X1 U6156 ( .A(n5154), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9087) );
  INV_X1 U6157 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5151) );
  INV_X1 U6158 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4979) );
  INV_X1 U6159 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4880) );
  NAND2_X1 U6160 ( .A1(n5885), .A2(n5886), .ZN(n8675) );
  NAND2_X1 U6161 ( .A1(n8007), .A2(n8393), .ZN(n7991) );
  AND2_X1 U6162 ( .A1(n5865), .A2(n5863), .ZN(n8393) );
  OR2_X1 U6163 ( .A1(n8578), .A2(n8541), .ZN(n4534) );
  NAND2_X1 U6164 ( .A1(n6540), .A2(n9262), .ZN(n8902) );
  XNOR2_X1 U6165 ( .A(n8901), .B(n6541), .ZN(n6540) );
  NAND2_X1 U6166 ( .A1(n8856), .A2(n6282), .ZN(n6460) );
  OAI21_X1 U6167 ( .B1(n6795), .B2(n4754), .A(n4751), .ZN(n6919) );
  NAND2_X2 U6168 ( .A1(n8238), .A2(n8106), .ZN(n8112) );
  NOR2_X2 U6169 ( .A1(n8181), .A2(n4426), .ZN(n8188) );
  AOI21_X2 U6170 ( .B1(n8055), .B2(n8054), .A(n8053), .ZN(n8181) );
  NAND2_X1 U6171 ( .A1(n8022), .A2(n5924), .ZN(n6343) );
  NAND2_X1 U6172 ( .A1(n6742), .A2(n6745), .ZN(n6744) );
  NAND2_X2 U6173 ( .A1(n7051), .A2(n7050), .ZN(n7148) );
  AOI22_X2 U6174 ( .A1(n9079), .A2(n9081), .B1(n9106), .B2(n9307), .ZN(n9064)
         );
  NAND2_X1 U6175 ( .A1(n8947), .A2(n8946), .ZN(n8949) );
  INV_X1 U6176 ( .A(n7491), .ZN(n6632) );
  NAND2_X1 U6177 ( .A1(n9283), .A2(n4711), .ZN(n4710) );
  OAI21_X1 U6178 ( .B1(n9213), .B2(n4871), .A(n4869), .ZN(n4868) );
  NAND2_X1 U6179 ( .A1(n4712), .A2(n4709), .ZN(n9348) );
  OAI22_X2 U6180 ( .A1(n7286), .A2(n7978), .B1(n7285), .B2(n8276), .ZN(n7287)
         );
  NAND2_X2 U6181 ( .A1(n8408), .A2(n8407), .ZN(n8406) );
  NAND2_X1 U6182 ( .A1(n4608), .A2(n4607), .ZN(P2_U3517) );
  NAND2_X1 U6183 ( .A1(n4974), .A2(n4972), .ZN(P2_U3549) );
  NAND2_X1 U6184 ( .A1(n5009), .A2(n4920), .ZN(n4672) );
  NAND2_X1 U6185 ( .A1(n8581), .A2(n4609), .ZN(n8659) );
  NAND2_X1 U6186 ( .A1(n4959), .A2(n4958), .ZN(n6956) );
  XNOR2_X1 U6187 ( .A(n8035), .B(n4900), .ZN(n8578) );
  NAND2_X1 U6188 ( .A1(n6681), .A2(n7491), .ZN(n6683) );
  NAND2_X4 U6189 ( .A1(n4494), .A2(n5190), .ZN(n6625) );
  AND3_X2 U6190 ( .A1(n4634), .A2(n4633), .A3(n4885), .ZN(n5159) );
  NAND3_X1 U6191 ( .A1(n4634), .A2(n4633), .A3(n4503), .ZN(n4502) );
  AND2_X2 U6192 ( .A1(n4878), .A2(n5125), .ZN(n4634) );
  NAND2_X1 U6193 ( .A1(n4507), .A2(n4504), .ZN(P1_U3240) );
  NAND2_X1 U6194 ( .A1(n4436), .A2(n4505), .ZN(n4504) );
  NAND3_X1 U6195 ( .A1(n4506), .A2(n4470), .A3(n4432), .ZN(n4505) );
  OR3_X1 U6196 ( .A1(n7614), .A2(n7610), .A3(n8929), .ZN(n4506) );
  NAND2_X1 U6197 ( .A1(n4410), .A2(n4525), .ZN(n4527) );
  NAND3_X1 U6198 ( .A1(n4527), .A2(n4835), .A3(n4530), .ZN(n4526) );
  OAI21_X1 U6199 ( .B1(n8581), .B2(n8518), .A(n4431), .ZN(P2_U3267) );
  NAND2_X1 U6200 ( .A1(n8376), .A2(n4475), .ZN(n4538) );
  NAND2_X1 U6201 ( .A1(n4538), .A2(n4539), .ZN(n8351) );
  AND2_X1 U6202 ( .A1(n8376), .A2(n4438), .ZN(n8366) );
  NAND3_X1 U6203 ( .A1(n5282), .A2(n5298), .A3(n5283), .ZN(n4540) );
  NAND3_X1 U6204 ( .A1(n4542), .A2(n7927), .A3(n7926), .ZN(n4541) );
  NAND3_X1 U6205 ( .A1(n4545), .A2(n4543), .A3(n8434), .ZN(n4542) );
  NAND2_X1 U6206 ( .A1(n4674), .A2(n4552), .ZN(n4551) );
  NAND2_X1 U6207 ( .A1(n4551), .A2(n4553), .ZN(n7998) );
  OR2_X1 U6208 ( .A1(n5342), .A2(n4894), .ZN(n4556) );
  NAND2_X1 U6209 ( .A1(n4556), .A2(n4891), .ZN(n5379) );
  OAI21_X2 U6210 ( .B1(n5342), .B2(n4558), .A(n4557), .ZN(n5393) );
  NAND3_X1 U6211 ( .A1(n4561), .A2(n7862), .A3(n4471), .ZN(n7866) );
  NAND2_X2 U6212 ( .A1(P2_U3152), .A2(n7428), .ZN(n7404) );
  INV_X2 U6213 ( .A(n5880), .ZN(n7428) );
  MUX2_X1 U6214 ( .A(n9979), .B(n10104), .S(n5880), .Z(n5026) );
  MUX2_X1 U6215 ( .A(n6062), .B(n6069), .S(n5880), .Z(n5023) );
  MUX2_X1 U6216 ( .A(n7129), .B(n7131), .S(n5880), .Z(n5107) );
  MUX2_X1 U6217 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n5880), .Z(n5660) );
  MUX2_X1 U6218 ( .A(n5722), .B(n5715), .S(n5880), .Z(n5716) );
  MUX2_X1 U6219 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n5880), .Z(n7424) );
  NAND2_X1 U6220 ( .A1(n6302), .A2(n6242), .ZN(n4567) );
  NAND2_X1 U6221 ( .A1(n4567), .A2(n4568), .ZN(n6201) );
  NOR2_X1 U6222 ( .A1(n6311), .A2(n6169), .ZN(n4569) );
  NAND2_X1 U6223 ( .A1(n6605), .A2(n4577), .ZN(n6609) );
  NAND2_X1 U6224 ( .A1(n4758), .A2(n5287), .ZN(n4577) );
  XNOR2_X1 U6225 ( .A(n4582), .B(n4581), .ZN(n6477) );
  NAND2_X2 U6226 ( .A1(n5776), .A2(n4584), .ZN(n5405) );
  NAND2_X1 U6227 ( .A1(n5461), .A2(n5460), .ZN(n7258) );
  NAND2_X1 U6228 ( .A1(n5585), .A2(n4593), .ZN(n4592) );
  NAND2_X1 U6229 ( .A1(n4592), .A2(n4594), .ZN(n5641) );
  NAND2_X1 U6230 ( .A1(n4596), .A2(n8788), .ZN(n8707) );
  INV_X1 U6231 ( .A(n4788), .ZN(n4597) );
  INV_X1 U6232 ( .A(n4601), .ZN(n8790) );
  AND2_X1 U6233 ( .A1(n5465), .A2(n4602), .ZN(n5547) );
  NAND2_X1 U6234 ( .A1(n5465), .A2(n4603), .ZN(n4804) );
  NOR2_X2 U6235 ( .A1(n5849), .A2(n5848), .ZN(n5852) );
  AOI211_X2 U6236 ( .C1(n8580), .C2(n9816), .A(n4611), .B(n4610), .ZN(n4609)
         );
  NAND2_X1 U6237 ( .A1(n8391), .A2(n4950), .ZN(n8381) );
  INV_X1 U6238 ( .A(n4616), .ZN(n8360) );
  INV_X1 U6239 ( .A(n4622), .ZN(n8506) );
  INV_X1 U6240 ( .A(n7123), .ZN(n4623) );
  NAND2_X1 U6241 ( .A1(n4623), .A2(n4624), .ZN(n7332) );
  NAND2_X1 U6242 ( .A1(n8471), .A2(n4628), .ZN(n8392) );
  XNOR2_X2 U6243 ( .A(n4635), .B(n5158), .ZN(n5773) );
  INV_X1 U6244 ( .A(n4639), .ZN(n9131) );
  INV_X1 U6245 ( .A(n4641), .ZN(n7355) );
  INV_X1 U6246 ( .A(n4648), .ZN(n9022) );
  NAND2_X1 U6247 ( .A1(n5020), .A2(n4655), .ZN(n4654) );
  NAND3_X1 U6248 ( .A1(n4654), .A2(n5283), .A3(n4653), .ZN(n4906) );
  NAND2_X1 U6249 ( .A1(n4657), .A2(n5022), .ZN(n4653) );
  AOI21_X1 U6250 ( .B1(n5258), .B2(n4659), .A(n4658), .ZN(n4656) );
  INV_X1 U6251 ( .A(n5258), .ZN(n4657) );
  OAI21_X1 U6252 ( .B1(n4670), .B2(n4669), .A(n4668), .ZN(n4667) );
  NAND3_X1 U6253 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .A3(n4921), .ZN(n4671) );
  NAND2_X1 U6254 ( .A1(n7952), .A2(n7951), .ZN(n4674) );
  OAI21_X1 U6255 ( .B1(n9228), .B2(n4684), .A(n4681), .ZN(n9160) );
  OR2_X1 U6256 ( .A1(n9051), .A2(n9050), .ZN(n4701) );
  INV_X1 U6257 ( .A(n4701), .ZN(n9049) );
  NOR2_X1 U6258 ( .A1(n9030), .A2(n8991), .ZN(n4700) );
  NAND2_X1 U6259 ( .A1(n9126), .A2(n4705), .ZN(n4702) );
  NAND2_X1 U6260 ( .A1(n4702), .A2(n4703), .ZN(n9080) );
  OAI21_X1 U6261 ( .B1(n7044), .B2(n4717), .A(n4714), .ZN(n7279) );
  NAND4_X1 U6262 ( .A1(n4878), .A2(n4879), .A3(n4718), .A4(n5125), .ZN(n5139)
         );
  OR2_X1 U6263 ( .A1(n7810), .A2(n10182), .ZN(n5881) );
  NAND2_X2 U6264 ( .A1(n6143), .A2(n7428), .ZN(n7810) );
  NAND2_X2 U6265 ( .A1(n5877), .A2(n5876), .ZN(n8037) );
  NAND2_X1 U6266 ( .A1(n8112), .A2(n4722), .ZN(n4721) );
  OAI211_X1 U6267 ( .C1(n8112), .C2(n4724), .A(n4721), .B(n8129), .ZN(P2_U3222) );
  NAND2_X1 U6268 ( .A1(n8112), .A2(n8132), .ZN(n8135) );
  NAND2_X1 U6269 ( .A1(n4841), .A2(n4732), .ZN(n5860) );
  NAND2_X1 U6270 ( .A1(n8188), .A2(n4474), .ZN(n4735) );
  OR2_X1 U6271 ( .A1(n8063), .A2(n8062), .ZN(n4743) );
  NAND2_X1 U6272 ( .A1(n6348), .A2(n5983), .ZN(n6424) );
  NAND3_X1 U6273 ( .A1(n8205), .A2(n6349), .A3(n5955), .ZN(n6348) );
  OAI21_X2 U6274 ( .B1(n8168), .B2(n4757), .A(n4756), .ZN(n8237) );
  OR2_X1 U6275 ( .A1(n6769), .A2(n6076), .ZN(n5882) );
  NAND2_X1 U6276 ( .A1(n7279), .A2(n7457), .ZN(n9463) );
  OAI21_X2 U6277 ( .B1(n9139), .B2(n8982), .A(n8981), .ZN(n9126) );
  INV_X1 U6278 ( .A(n8174), .ZN(n8055) );
  XNOR2_X2 U6279 ( .A(n4402), .B(n9758), .ZN(n8014) );
  INV_X1 U6280 ( .A(n6603), .ZN(n4758) );
  NAND2_X1 U6281 ( .A1(n5348), .A2(n4761), .ZN(n4760) );
  NAND3_X1 U6282 ( .A1(n5544), .A2(n4768), .A3(n4769), .ZN(n4767) );
  NAND2_X1 U6283 ( .A1(n4771), .A2(n8828), .ZN(n4770) );
  INV_X1 U6284 ( .A(n8736), .ZN(n4772) );
  NAND2_X1 U6285 ( .A1(n8766), .A2(n4782), .ZN(n4773) );
  NAND2_X1 U6286 ( .A1(n4776), .A2(n4773), .ZN(n8750) );
  MUX2_X1 U6287 ( .A(n6624), .B(n6623), .S(n5171), .Z(n9473) );
  NAND2_X1 U6288 ( .A1(n5547), .A2(n4805), .ZN(n4803) );
  NAND2_X1 U6289 ( .A1(n5547), .A2(n5132), .ZN(n5153) );
  NAND2_X1 U6290 ( .A1(n4809), .A2(n7392), .ZN(n5525) );
  NAND2_X1 U6291 ( .A1(n4809), .A2(n4808), .ZN(n8822) );
  XNOR2_X1 U6292 ( .A(n7816), .B(n8385), .ZN(n4810) );
  XNOR2_X2 U6293 ( .A(n8284), .B(n4812), .ZN(n7836) );
  OR2_X1 U6294 ( .A1(n8351), .A2(n4825), .ZN(n4824) );
  NAND2_X1 U6295 ( .A1(n8459), .A2(n4833), .ZN(n4832) );
  INV_X1 U6296 ( .A(n4834), .ZN(n8457) );
  INV_X1 U6297 ( .A(n5849), .ZN(n4841) );
  AND3_X2 U6298 ( .A1(n4841), .A2(n4843), .A3(n4840), .ZN(n5885) );
  NAND2_X1 U6299 ( .A1(n5852), .A2(n5850), .ZN(n5869) );
  NAND2_X1 U6300 ( .A1(n4846), .A2(n4845), .ZN(n9017) );
  NOR2_X1 U6301 ( .A1(n9060), .A2(n9076), .ZN(n4850) );
  NAND2_X1 U6302 ( .A1(n9124), .A2(n4411), .ZN(n4851) );
  NAND2_X1 U6303 ( .A1(n4851), .A2(n4852), .ZN(n9079) );
  OAI21_X1 U6304 ( .B1(n9457), .B2(n7271), .A(n7270), .ZN(n7348) );
  NAND2_X1 U6305 ( .A1(n7271), .A2(n7270), .ZN(n4867) );
  INV_X1 U6306 ( .A(n4868), .ZN(n9151) );
  AND2_X1 U6307 ( .A1(n9335), .A2(n9162), .ZN(n4876) );
  NAND2_X1 U6308 ( .A1(n6744), .A2(n4430), .ZN(n6942) );
  NAND2_X1 U6309 ( .A1(n5145), .A2(n5147), .ZN(n5142) );
  NAND2_X1 U6310 ( .A1(n5009), .A2(n4920), .ZN(n4918) );
  NAND3_X1 U6311 ( .A1(n4921), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4919) );
  OAI21_X1 U6312 ( .B1(n5587), .B2(n4925), .A(n4922), .ZN(n5610) );
  OAI21_X1 U6313 ( .B1(n5587), .B2(n5586), .A(n5095), .ZN(n5174) );
  NAND2_X1 U6314 ( .A1(n5051), .A2(n5050), .ZN(n5412) );
  OAI21_X2 U6315 ( .B1(n5051), .B2(n4931), .A(n4929), .ZN(n5463) );
  INV_X1 U6316 ( .A(n4935), .ZN(n8344) );
  OAI21_X2 U6317 ( .B1(n8406), .B2(n4939), .A(n4936), .ZN(n4935) );
  NAND2_X1 U6318 ( .A1(n6505), .A2(n9758), .ZN(n7959) );
  NAND2_X1 U6319 ( .A1(n6559), .A2(n4444), .ZN(n4959) );
  NAND2_X1 U6320 ( .A1(n6644), .A2(n6643), .ZN(n4960) );
  AOI21_X1 U6321 ( .B1(n4954), .B2(n6644), .A(n4457), .ZN(n4958) );
  NAND2_X1 U6322 ( .A1(n4957), .A2(n4960), .ZN(n6727) );
  OR2_X1 U6323 ( .A1(n8456), .A2(n4965), .ZN(n4961) );
  AND2_X2 U6324 ( .A1(n4961), .A2(n4962), .ZN(n8408) );
  INV_X1 U6325 ( .A(n4971), .ZN(n8433) );
  NAND2_X1 U6326 ( .A1(n4977), .A2(n4975), .ZN(n6612) );
  NAND3_X1 U6327 ( .A1(n6511), .A2(n6560), .A3(n7967), .ZN(n4977) );
  NAND2_X1 U6328 ( .A1(n8543), .A2(n4415), .ZN(n4980) );
  NAND2_X1 U6329 ( .A1(n4980), .A2(n4981), .ZN(n8505) );
  INV_X1 U6330 ( .A(n4983), .ZN(n8545) );
  NAND3_X1 U6331 ( .A1(n5835), .A2(n5834), .A3(n5941), .ZN(n6442) );
  NAND2_X1 U6332 ( .A1(n7339), .A2(n4985), .ZN(n4984) );
  NAND2_X1 U6333 ( .A1(n4984), .A2(n7366), .ZN(n7371) );
  NAND2_X1 U6334 ( .A1(n7114), .A2(n4987), .ZN(n7164) );
  NAND2_X1 U6335 ( .A1(n6380), .A2(n6381), .ZN(n6379) );
  XNOR2_X1 U6336 ( .A(n7423), .B(SI_30_), .ZN(n8086) );
  NAND2_X1 U6337 ( .A1(n6778), .A2(n6862), .ZN(n6795) );
  XNOR2_X1 U6338 ( .A(n8089), .B(n8076), .ZN(n8081) );
  NAND2_X1 U6339 ( .A1(n7791), .A2(n7939), .ZN(n8033) );
  NAND2_X1 U6340 ( .A1(n5714), .A2(n5713), .ZN(n5720) );
  NAND2_X1 U6341 ( .A1(n5693), .A2(n5692), .ZN(n5714) );
  NAND2_X1 U6342 ( .A1(n5463), .A2(n5001), .ZN(n5067) );
  NAND2_X1 U6343 ( .A1(n5083), .A2(n5082), .ZN(n5546) );
  NAND2_X1 U6344 ( .A1(n5527), .A2(n5526), .ZN(n5083) );
  XNOR2_X1 U6345 ( .A(n5393), .B(n5000), .ZN(n6881) );
  BUF_X4 U6346 ( .A(n5016), .Z(n7411) );
  AOI21_X1 U6347 ( .B1(n5823), .B2(n4990), .A(n5822), .ZN(n5824) );
  NAND2_X1 U6348 ( .A1(n5880), .A2(n5005), .ZN(n5011) );
  NAND2_X1 U6349 ( .A1(n8950), .A2(n4423), .ZN(n8952) );
  NAND2_X1 U6350 ( .A1(n8822), .A2(n8823), .ZN(n8828) );
  OR2_X1 U6351 ( .A1(n5885), .A2(n5992), .ZN(n5887) );
  OR2_X1 U6352 ( .A1(n7802), .A2(n6146), .ZN(n5915) );
  NAND2_X1 U6353 ( .A1(n4401), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5918) );
  AOI21_X1 U6354 ( .B1(n8547), .B2(n7894), .A(n7896), .ZN(n8527) );
  INV_X1 U6355 ( .A(n6625), .ZN(n6592) );
  INV_X1 U6356 ( .A(n5773), .ZN(n6628) );
  OR2_X1 U6357 ( .A1(n5785), .A2(n5784), .ZN(n4989) );
  AND3_X1 U6358 ( .A1(n5807), .A2(n5806), .A3(n8812), .ZN(n4990) );
  AND2_X1 U6359 ( .A1(n8377), .A2(n8375), .ZN(n4993) );
  AND2_X1 U6360 ( .A1(n5861), .A2(n5866), .ZN(n4995) );
  AND2_X1 U6361 ( .A1(n8052), .A2(n8051), .ZN(n4996) );
  AND2_X1 U6362 ( .A1(n8478), .A2(n8479), .ZN(n4997) );
  AND2_X1 U6363 ( .A1(n4407), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4998) );
  AND2_X1 U6364 ( .A1(n6510), .A2(n6505), .ZN(n4999) );
  INV_X1 U6365 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5850) );
  INV_X1 U6366 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5886) );
  AND2_X1 U6367 ( .A1(n5050), .A2(n5049), .ZN(n5000) );
  AND4_X1 U6368 ( .A1(n5769), .A2(n5768), .A3(n5767), .A4(n5766), .ZN(n9037)
         );
  AND2_X1 U6369 ( .A1(n5045), .A2(n5044), .ZN(n5002) );
  OR2_X1 U6370 ( .A1(n8462), .A2(n5905), .ZN(n5003) );
  AND4_X1 U6371 ( .A1(n7701), .A2(n7700), .A3(n7699), .A4(n7698), .ZN(n8551)
         );
  AND2_X1 U6372 ( .A1(n5209), .A2(n5208), .ZN(n5004) );
  XNOR2_X1 U6373 ( .A(n7406), .B(n7405), .ZN(n7792) );
  AND2_X1 U6374 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n5005) );
  INV_X1 U6375 ( .A(n8939), .ZN(n7485) );
  AND2_X1 U6376 ( .A1(n8497), .A2(n8498), .ZN(n5006) );
  AND2_X1 U6377 ( .A1(n9291), .A2(n8819), .ZN(n5007) );
  INV_X1 U6378 ( .A(n9038), .ZN(n9030) );
  INV_X1 U6379 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5122) );
  NAND2_X1 U6380 ( .A1(n7950), .A2(n7841), .ZN(n7951) );
  OAI22_X1 U6381 ( .A1(n6749), .A2(n5405), .B1(n9681), .B2(n5261), .ZN(n5262)
         );
  INV_X1 U6382 ( .A(n9037), .ZN(n8966) );
  INV_X1 U6383 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5119) );
  INV_X1 U6384 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6922) );
  INV_X1 U6385 ( .A(n8094), .ZN(n8095) );
  AOI21_X1 U6386 ( .B1(n7815), .B2(n7988), .A(n7953), .ZN(n7816) );
  INV_X1 U6387 ( .A(n7706), .ZN(n6121) );
  NAND2_X1 U6388 ( .A1(n8334), .A2(n8265), .ZN(n8039) );
  INV_X1 U6389 ( .A(n7756), .ZN(n6372) );
  NAND2_X1 U6390 ( .A1(n5239), .A2(n5238), .ZN(n5240) );
  INV_X1 U6391 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5370) );
  INV_X1 U6392 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5158) );
  INV_X1 U6393 ( .A(n5610), .ZN(n5101) );
  INV_X1 U6394 ( .A(n6030), .ZN(n6028) );
  NAND2_X1 U6395 ( .A1(n8096), .A2(n8095), .ZN(n8097) );
  NAND2_X1 U6396 ( .A1(n6122), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7726) );
  OR2_X1 U6397 ( .A1(n7726), .A2(n8159), .ZN(n7744) );
  INV_X1 U6398 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10040) );
  NAND2_X1 U6399 ( .A1(n8040), .A2(n8039), .ZN(n8041) );
  OR2_X1 U6400 ( .A1(n7766), .A2(n8169), .ZN(n7778) );
  NAND2_X1 U6401 ( .A1(n7851), .A2(n7848), .ZN(n6726) );
  INV_X1 U6402 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n5611) );
  INV_X1 U6403 ( .A(n7261), .ZN(n5460) );
  INV_X1 U6404 ( .A(n5524), .ZN(n5521) );
  NAND2_X1 U6405 ( .A1(n5698), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5761) );
  AND2_X1 U6406 ( .A1(n5591), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U6407 ( .A1(n4408), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5189) );
  NOR2_X1 U6408 ( .A1(n5614), .A2(n8724), .ZN(n5633) );
  NOR2_X1 U6409 ( .A1(n5551), .A2(n10190), .ZN(n5573) );
  OR2_X1 U6410 ( .A1(n5446), .A2(n5445), .ZN(n5470) );
  AND2_X1 U6411 ( .A1(n8974), .A2(n8976), .ZN(n9227) );
  NAND2_X1 U6412 ( .A1(n7406), .A2(n7405), .ZN(n7410) );
  NAND2_X1 U6413 ( .A1(n6000), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6043) );
  OR2_X1 U6414 ( .A1(n8120), .A2(n8119), .ZN(n8121) );
  AND2_X1 U6415 ( .A1(n8069), .A2(n8068), .ZN(n8070) );
  OR2_X1 U6416 ( .A1(n8179), .A2(n4996), .ZN(n8053) );
  INV_X1 U6417 ( .A(n8088), .ZN(n8076) );
  INV_X1 U6418 ( .A(n8236), .ZN(n8104) );
  OR2_X1 U6419 ( .A1(n8347), .A2(n7746), .ZN(n7805) );
  INV_X1 U6420 ( .A(n4401), .ZN(n7783) );
  INV_X1 U6421 ( .A(n6493), .ZN(n6489) );
  AND2_X1 U6422 ( .A1(n6081), .A2(n6053), .ZN(n9751) );
  NAND2_X1 U6423 ( .A1(n8477), .A2(n4997), .ZN(n8484) );
  INV_X1 U6424 ( .A(n9751), .ZN(n8548) );
  NAND2_X1 U6425 ( .A1(n5738), .A2(n4585), .ZN(n7610) );
  OR2_X1 U6426 ( .A1(n5805), .A2(n5804), .ZN(n5790) );
  XNOR2_X1 U6427 ( .A(n5245), .B(n5243), .ZN(n6469) );
  OR2_X1 U6428 ( .A1(n5782), .A2(n6628), .ZN(n8830) );
  OR2_X1 U6429 ( .A1(n5782), .A2(n5773), .ZN(n8816) );
  INV_X1 U6430 ( .A(n5776), .ZN(n5825) );
  INV_X1 U6431 ( .A(n9663), .ZN(n9645) );
  INV_X1 U6432 ( .A(n9297), .ZN(n9060) );
  NAND2_X1 U6433 ( .A1(n7593), .A2(n8988), .ZN(n9072) );
  NOR2_X1 U6434 ( .A1(n9112), .A2(n9130), .ZN(n8960) );
  INV_X1 U6435 ( .A(n9223), .ZN(n9479) );
  AND2_X1 U6436 ( .A1(n6671), .A2(n6670), .ZN(n6949) );
  INV_X1 U6437 ( .A(n9723), .ZN(n9711) );
  INV_X1 U6438 ( .A(n9709), .ZN(n9705) );
  AND2_X1 U6439 ( .A1(n5777), .A2(n9678), .ZN(n6671) );
  NAND2_X1 U6440 ( .A1(n5139), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5127) );
  NAND2_X1 U6441 ( .A1(n5091), .A2(n5090), .ZN(n5587) );
  AND2_X1 U6442 ( .A1(n5082), .A2(n5081), .ZN(n5526) );
  NAND2_X1 U6443 ( .A1(n8011), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8253) );
  NAND2_X1 U6444 ( .A1(n6424), .A2(n5987), .ZN(n6031) );
  INV_X1 U6445 ( .A(n8550), .ZN(n9752) );
  INV_X1 U6446 ( .A(n7768), .ZN(n7780) );
  INV_X1 U6447 ( .A(n9896), .ZN(n9740) );
  INV_X1 U6448 ( .A(n9741), .ZN(n9891) );
  AND2_X1 U6449 ( .A1(n6176), .A2(n6175), .ZN(n9896) );
  INV_X1 U6450 ( .A(n8034), .ZN(n8352) );
  INV_X1 U6451 ( .A(n8489), .ZN(n8490) );
  NAND2_X1 U6452 ( .A1(n7863), .A2(n7874), .ZN(n7976) );
  INV_X1 U6453 ( .A(n9756), .ZN(n8556) );
  INV_X1 U6454 ( .A(n8535), .ZN(n8555) );
  AND2_X1 U6455 ( .A1(n9771), .A2(n6033), .ZN(n9756) );
  AND3_X1 U6456 ( .A1(n9771), .A2(n6552), .A3(n6551), .ZN(n6553) );
  INV_X1 U6457 ( .A(n9816), .ZN(n9833) );
  AND2_X1 U6458 ( .A1(n6032), .A2(n7819), .ZN(n9829) );
  INV_X1 U6459 ( .A(n8644), .ZN(n9837) );
  AND2_X1 U6460 ( .A1(n6038), .A2(n9777), .ZN(n9771) );
  XNOR2_X1 U6461 ( .A(n5851), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6015) );
  AND2_X1 U6462 ( .A1(n5786), .A2(n6671), .ZN(n7063) );
  INV_X1 U6463 ( .A(n8830), .ZN(n8807) );
  INV_X1 U6464 ( .A(n8816), .ZN(n8833) );
  AND4_X1 U6465 ( .A1(n5678), .A2(n5677), .A3(n5676), .A4(n5675), .ZN(n9083)
         );
  AND4_X1 U6466 ( .A1(n5538), .A2(n5537), .A3(n5536), .A4(n5535), .ZN(n9198)
         );
  AND2_X1 U6467 ( .A1(n9614), .A2(n9613), .ZN(n9616) );
  INV_X1 U6468 ( .A(n9675), .ZN(n9581) );
  AND2_X1 U6469 ( .A1(n9529), .A2(n6628), .ZN(n9663) );
  INV_X1 U6470 ( .A(n9630), .ZN(n9670) );
  AND2_X1 U6471 ( .A1(n9101), .A2(n8984), .ZN(n9117) );
  AND2_X1 U6472 ( .A1(n9479), .A2(n8929), .ZN(n9193) );
  AND2_X1 U6473 ( .A1(n7634), .A2(n7525), .ZN(n7085) );
  INV_X1 U6474 ( .A(n9223), .ZN(n9269) );
  INV_X1 U6475 ( .A(n9686), .ZN(n9715) );
  OR2_X1 U6476 ( .A1(n6635), .A2(n7615), .ZN(n9723) );
  INV_X1 U6477 ( .A(n9725), .ZN(n9687) );
  NAND2_X1 U6478 ( .A1(n9473), .A2(n9715), .ZN(n9725) );
  AND2_X1 U6479 ( .A1(n7602), .A2(n7013), .ZN(n9686) );
  NAND2_X1 U6480 ( .A1(n5746), .A2(n5745), .ZN(n9677) );
  XNOR2_X1 U6481 ( .A(n5127), .B(n5126), .ZN(n6274) );
  XNOR2_X1 U6482 ( .A(n5152), .B(n5151), .ZN(n5170) );
  INV_X1 U6483 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9994) );
  INV_X1 U6484 ( .A(n9888), .ZN(n9739) );
  NAND2_X1 U6485 ( .A1(n6050), .A2(n6027), .ZN(n8263) );
  INV_X1 U6486 ( .A(n8200), .ZN(n8416) );
  AND4_X1 U6487 ( .A1(n6111), .A2(n6110), .A3(n6109), .A4(n6108), .ZN(n8549)
         );
  OR2_X1 U6488 ( .A1(n8545), .A2(n8544), .ZN(n9441) );
  INV_X1 U6489 ( .A(n9775), .ZN(n9772) );
  INV_X1 U6490 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U6491 ( .A1(n5760), .A2(n5772), .ZN(n8825) );
  INV_X1 U6492 ( .A(n9083), .ZN(n8962) );
  INV_X1 U6493 ( .A(n9198), .ZN(n9230) );
  INV_X1 U6494 ( .A(n7049), .ZN(n8843) );
  OR2_X1 U6495 ( .A1(n9528), .A2(n8936), .ZN(n9630) );
  INV_X1 U6496 ( .A(n9461), .ZN(n9239) );
  NAND2_X1 U6497 ( .A1(n9479), .A2(n6723), .ZN(n9271) );
  AND2_X2 U6498 ( .A1(n6672), .A2(n9476), .ZN(n9223) );
  AND2_X2 U6499 ( .A1(n6336), .A2(n6335), .ZN(n9737) );
  AND3_X1 U6500 ( .A1(n9694), .A2(n9693), .A3(n9692), .ZN(n9731) );
  AND2_X2 U6501 ( .A1(n6336), .A2(n6332), .ZN(n9729) );
  AND2_X1 U6502 ( .A1(n9678), .A2(n9677), .ZN(n9679) );
  INV_X1 U6503 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7344) );
  INV_X1 U6504 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7012) );
  INV_X1 U6505 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6230) );
  INV_X1 U6506 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10161) );
  NOR2_X1 U6507 ( .A1(n10211), .A2(n10210), .ZN(n10209) );
  NOR2_X1 U6508 ( .A1(n9881), .A2(n9880), .ZN(n9879) );
  INV_X1 U6509 ( .A(n8271), .ZN(P2_U3966) );
  INV_X1 U6510 ( .A(n8846), .ZN(P1_U4006) );
  AND2_X1 U6511 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n5010) );
  INV_X1 U6512 ( .A(SI_1_), .ZN(n5012) );
  XNOR2_X1 U6513 ( .A(n5013), .B(n5012), .ZN(n5194) );
  MUX2_X1 U6514 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5016), .Z(n5193) );
  NAND2_X1 U6515 ( .A1(n5194), .A2(n5193), .ZN(n5015) );
  NAND2_X1 U6516 ( .A1(n5013), .A2(SI_1_), .ZN(n5014) );
  INV_X1 U6517 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6067) );
  INV_X1 U6518 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6059) );
  MUX2_X1 U6519 ( .A(n6067), .B(n6059), .S(n5016), .Z(n5017) );
  XNOR2_X1 U6520 ( .A(n5017), .B(SI_2_), .ZN(n5227) );
  NAND2_X1 U6521 ( .A1(n5228), .A2(n5227), .ZN(n5020) );
  INV_X1 U6522 ( .A(n5017), .ZN(n5018) );
  NAND2_X1 U6523 ( .A1(n5018), .A2(SI_2_), .ZN(n5019) );
  INV_X1 U6524 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6073) );
  INV_X1 U6525 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U6526 ( .A1(n5021), .A2(SI_3_), .ZN(n5022) );
  XNOR2_X1 U6527 ( .A(n5023), .B(SI_4_), .ZN(n5283) );
  INV_X1 U6528 ( .A(n5023), .ZN(n5024) );
  NAND2_X1 U6529 ( .A1(n5024), .A2(SI_4_), .ZN(n5025) );
  XNOR2_X1 U6530 ( .A(n5026), .B(SI_5_), .ZN(n5298) );
  INV_X1 U6531 ( .A(n5026), .ZN(n5027) );
  MUX2_X1 U6532 ( .A(n9981), .B(n6064), .S(n7411), .Z(n5028) );
  XNOR2_X1 U6533 ( .A(n5028), .B(SI_6_), .ZN(n5316) );
  NAND2_X1 U6534 ( .A1(n5317), .A2(n5316), .ZN(n5031) );
  INV_X1 U6535 ( .A(n5028), .ZN(n5029) );
  NAND2_X1 U6536 ( .A1(n5029), .A2(SI_6_), .ZN(n5030) );
  MUX2_X1 U6537 ( .A(n10158), .B(n6074), .S(n7411), .Z(n5032) );
  XNOR2_X1 U6538 ( .A(n5032), .B(SI_7_), .ZN(n5341) );
  INV_X1 U6539 ( .A(n5032), .ZN(n5033) );
  NAND2_X1 U6540 ( .A1(n5033), .A2(SI_7_), .ZN(n5034) );
  MUX2_X1 U6541 ( .A(n6078), .B(n6080), .S(n7411), .Z(n5036) );
  INV_X1 U6542 ( .A(SI_8_), .ZN(n5035) );
  NAND2_X1 U6543 ( .A1(n5036), .A2(n5035), .ZN(n5039) );
  INV_X1 U6544 ( .A(n5036), .ZN(n5037) );
  NAND2_X1 U6545 ( .A1(n5037), .A2(SI_8_), .ZN(n5038) );
  NAND2_X1 U6546 ( .A1(n5039), .A2(n5038), .ZN(n5357) );
  INV_X1 U6547 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5040) );
  MUX2_X1 U6548 ( .A(n5040), .B(n10161), .S(n7411), .Z(n5042) );
  INV_X1 U6549 ( .A(SI_9_), .ZN(n5041) );
  NAND2_X1 U6550 ( .A1(n5042), .A2(n5041), .ZN(n5045) );
  INV_X1 U6551 ( .A(n5042), .ZN(n5043) );
  NAND2_X1 U6552 ( .A1(n5043), .A2(SI_9_), .ZN(n5044) );
  MUX2_X1 U6553 ( .A(n10117), .B(n6099), .S(n7411), .Z(n5047) );
  INV_X1 U6554 ( .A(SI_10_), .ZN(n5046) );
  NAND2_X1 U6555 ( .A1(n5047), .A2(n5046), .ZN(n5050) );
  INV_X1 U6556 ( .A(n5047), .ZN(n5048) );
  NAND2_X1 U6557 ( .A1(n5048), .A2(SI_10_), .ZN(n5049) );
  NAND2_X1 U6558 ( .A1(n5393), .A2(n5000), .ZN(n5051) );
  INV_X1 U6559 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5052) );
  MUX2_X1 U6560 ( .A(n5052), .B(n6114), .S(n7411), .Z(n5053) );
  XNOR2_X1 U6561 ( .A(n5053), .B(SI_11_), .ZN(n5411) );
  INV_X1 U6562 ( .A(n5411), .ZN(n5056) );
  INV_X1 U6563 ( .A(n5053), .ZN(n5054) );
  NAND2_X1 U6564 ( .A1(n5054), .A2(SI_11_), .ZN(n5055) );
  MUX2_X1 U6565 ( .A(n9970), .B(n6132), .S(n7411), .Z(n5058) );
  INV_X1 U6566 ( .A(SI_12_), .ZN(n5057) );
  INV_X1 U6567 ( .A(n5058), .ZN(n5059) );
  NAND2_X1 U6568 ( .A1(n5059), .A2(SI_12_), .ZN(n5060) );
  NAND2_X1 U6569 ( .A1(n5061), .A2(n5060), .ZN(n5439) );
  MUX2_X1 U6570 ( .A(n6224), .B(n10026), .S(n7428), .Z(n5063) );
  INV_X1 U6571 ( .A(SI_13_), .ZN(n5062) );
  INV_X1 U6572 ( .A(n5063), .ZN(n5064) );
  NAND2_X1 U6573 ( .A1(n5064), .A2(SI_13_), .ZN(n5065) );
  MUX2_X1 U6574 ( .A(n6229), .B(n6230), .S(n7428), .Z(n5069) );
  INV_X1 U6575 ( .A(n5069), .ZN(n5070) );
  NAND2_X1 U6576 ( .A1(n5070), .A2(SI_14_), .ZN(n5071) );
  MUX2_X1 U6577 ( .A(n6440), .B(n10060), .S(n7428), .Z(n5073) );
  INV_X1 U6578 ( .A(SI_15_), .ZN(n5072) );
  NAND2_X1 U6579 ( .A1(n5073), .A2(n5072), .ZN(n5076) );
  INV_X1 U6580 ( .A(n5073), .ZN(n5074) );
  NAND2_X1 U6581 ( .A1(n5074), .A2(SI_15_), .ZN(n5075) );
  NAND2_X1 U6582 ( .A1(n5076), .A2(n5075), .ZN(n5503) );
  INV_X1 U6583 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5077) );
  MUX2_X1 U6584 ( .A(n6445), .B(n5077), .S(n7428), .Z(n5079) );
  INV_X1 U6585 ( .A(SI_16_), .ZN(n5078) );
  INV_X1 U6586 ( .A(n5079), .ZN(n5080) );
  NAND2_X1 U6587 ( .A1(n5080), .A2(SI_16_), .ZN(n5081) );
  MUX2_X1 U6588 ( .A(n6501), .B(n6503), .S(n7428), .Z(n5084) );
  XNOR2_X1 U6589 ( .A(n5084), .B(SI_17_), .ZN(n5545) );
  INV_X1 U6590 ( .A(n5545), .ZN(n5087) );
  INV_X1 U6591 ( .A(n5084), .ZN(n5085) );
  NAND2_X1 U6592 ( .A1(n5085), .A2(SI_17_), .ZN(n5086) );
  MUX2_X1 U6593 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7428), .Z(n5089) );
  XNOR2_X1 U6594 ( .A(n5089), .B(SI_18_), .ZN(n5565) );
  NAND2_X1 U6595 ( .A1(n5566), .A2(n5088), .ZN(n5091) );
  NAND2_X1 U6596 ( .A1(n5089), .A2(SI_18_), .ZN(n5090) );
  MUX2_X1 U6597 ( .A(n6857), .B(n10058), .S(n7428), .Z(n5092) );
  INV_X1 U6598 ( .A(SI_19_), .ZN(n10163) );
  NAND2_X1 U6599 ( .A1(n5092), .A2(n10163), .ZN(n5095) );
  INV_X1 U6600 ( .A(n5092), .ZN(n5093) );
  NAND2_X1 U6601 ( .A1(n5093), .A2(SI_19_), .ZN(n5094) );
  NAND2_X1 U6602 ( .A1(n5095), .A2(n5094), .ZN(n5586) );
  MUX2_X1 U6603 ( .A(n10070), .B(n7012), .S(n7428), .Z(n5097) );
  INV_X1 U6604 ( .A(SI_20_), .ZN(n5096) );
  NAND2_X1 U6605 ( .A1(n5097), .A2(n5096), .ZN(n5100) );
  INV_X1 U6606 ( .A(n5097), .ZN(n5098) );
  NAND2_X1 U6607 ( .A1(n5098), .A2(SI_20_), .ZN(n5099) );
  MUX2_X1 U6608 ( .A(n7067), .B(n5611), .S(n7428), .Z(n5102) );
  XNOR2_X1 U6609 ( .A(n5102), .B(SI_21_), .ZN(n5609) );
  NAND2_X1 U6610 ( .A1(n5101), .A2(n5609), .ZN(n5105) );
  INV_X1 U6611 ( .A(n5102), .ZN(n5103) );
  NAND2_X1 U6612 ( .A1(n5103), .A2(SI_21_), .ZN(n5104) );
  INV_X1 U6613 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7131) );
  INV_X1 U6614 ( .A(SI_22_), .ZN(n5106) );
  NAND2_X1 U6615 ( .A1(n5107), .A2(n5106), .ZN(n5110) );
  INV_X1 U6616 ( .A(n5107), .ZN(n5108) );
  NAND2_X1 U6617 ( .A1(n5108), .A2(SI_22_), .ZN(n5109) );
  NAND2_X1 U6618 ( .A1(n5110), .A2(n5109), .ZN(n5628) );
  INV_X1 U6619 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5111) );
  MUX2_X1 U6620 ( .A(n5111), .B(n7179), .S(n7428), .Z(n5113) );
  INV_X1 U6621 ( .A(SI_23_), .ZN(n5112) );
  NAND2_X1 U6622 ( .A1(n5113), .A2(n5112), .ZN(n5116) );
  INV_X1 U6623 ( .A(n5113), .ZN(n5114) );
  NAND2_X1 U6624 ( .A1(n5114), .A2(SI_23_), .ZN(n5115) );
  INV_X1 U6625 ( .A(SI_24_), .ZN(n5117) );
  XNOR2_X1 U6626 ( .A(n5660), .B(n5117), .ZN(n5659) );
  XNOR2_X1 U6627 ( .A(n5663), .B(n5659), .ZN(n7752) );
  NOR2_X1 U6628 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5121) );
  NAND4_X1 U6629 ( .A1(n5121), .A2(n5120), .A3(n5133), .A4(n5567), .ZN(n5124)
         );
  NAND4_X1 U6630 ( .A1(n5151), .A2(n5122), .A3(n5505), .A4(n5130), .ZN(n5123)
         );
  NAND2_X1 U6631 ( .A1(n7752), .A2(n7415), .ZN(n5129) );
  NAND2_X4 U6632 ( .A1(n5191), .A2(n5880), .ZN(n7478) );
  INV_X1 U6633 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10071) );
  OR2_X1 U6634 ( .A1(n7478), .A2(n10071), .ZN(n5128) );
  NOR2_X1 U6635 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5132) );
  INV_X1 U6636 ( .A(n5134), .ZN(n5135) );
  NAND2_X1 U6637 ( .A1(n5150), .A2(n5136), .ZN(n5736) );
  NAND2_X1 U6638 ( .A1(n4442), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5140) );
  NAND2_X1 U6639 ( .A1(n5142), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5143) );
  MUX2_X1 U6640 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5143), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5144) );
  NAND2_X1 U6641 ( .A1(n5144), .A2(n4442), .ZN(n7346) );
  INV_X1 U6642 ( .A(n5145), .ZN(n5146) );
  NAND2_X1 U6643 ( .A1(n5146), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5148) );
  NOR2_X1 U6644 ( .A1(n7346), .A2(n7232), .ZN(n5149) );
  NAND2_X1 U6645 ( .A1(n5153), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U6646 ( .A1(n5170), .A2(n7668), .ZN(n5155) );
  NOR2_X1 U6647 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n5156) );
  NAND2_X1 U6648 ( .A1(n5159), .A2(n5156), .ZN(n9365) );
  NAND2_X1 U6649 ( .A1(n5697), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5169) );
  INV_X1 U6650 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n5162) );
  OR2_X1 U6651 ( .A1(n5670), .A2(n5162), .ZN(n5168) );
  NAND2_X1 U6652 ( .A1(n5292), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6653 ( .A1(n5334), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5350) );
  INV_X1 U6654 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5445) );
  INV_X1 U6655 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5469) );
  INV_X1 U6656 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5489) );
  NAND2_X1 U6657 ( .A1(n5511), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5533) );
  INV_X1 U6658 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5532) );
  INV_X1 U6659 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n10190) );
  INV_X1 U6660 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8724) );
  INV_X1 U6661 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8769) );
  NAND2_X1 U6662 ( .A1(n5647), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5646) );
  OAI21_X1 U6663 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n5164), .A(n5672), .ZN(
        n9086) );
  OR2_X1 U6664 ( .A1(n4404), .A2(n9086), .ZN(n5167) );
  INV_X1 U6665 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n5165) );
  OR2_X1 U6666 ( .A1(n5812), .A2(n5165), .ZN(n5166) );
  AOI22_X1 U6667 ( .A1(n9307), .A2(n5734), .B1(n5801), .B2(n9106), .ZN(n5656)
         );
  INV_X1 U6668 ( .A(n5656), .ZN(n5658) );
  INV_X2 U6669 ( .A(n5405), .ZN(n5734) );
  AOI22_X1 U6670 ( .A1(n9307), .A2(n5796), .B1(n5734), .B2(n9106), .ZN(n5172)
         );
  XNOR2_X1 U6671 ( .A(n5172), .B(n5799), .ZN(n5655) );
  INV_X1 U6672 ( .A(n5655), .ZN(n5657) );
  XNOR2_X1 U6673 ( .A(n5174), .B(n5173), .ZN(n7721) );
  NAND2_X1 U6674 ( .A1(n7721), .A2(n7415), .ZN(n5176) );
  OR2_X1 U6675 ( .A1(n7478), .A2(n7012), .ZN(n5175) );
  INV_X1 U6676 ( .A(n9325), .ZN(n8958) );
  OR2_X1 U6677 ( .A1(n5593), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6678 ( .A1(n5177), .A2(n5614), .ZN(n9143) );
  NAND2_X1 U6679 ( .A1(n5697), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5180) );
  NAND2_X1 U6680 ( .A1(n7418), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5179) );
  AND2_X1 U6681 ( .A1(n5180), .A2(n5179), .ZN(n5182) );
  NAND2_X1 U6682 ( .A1(n5221), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5181) );
  OAI211_X1 U6683 ( .C1(n9143), .C2(n4404), .A(n5182), .B(n5181), .ZN(n9163)
         );
  INV_X1 U6684 ( .A(n9163), .ZN(n9129) );
  OAI22_X1 U6685 ( .A1(n8958), .A2(n5405), .B1(n9129), .B2(n5732), .ZN(n5605)
         );
  INV_X1 U6686 ( .A(n5605), .ZN(n5608) );
  NAND2_X1 U6687 ( .A1(n9325), .A2(n5796), .ZN(n5184) );
  NAND2_X1 U6688 ( .A1(n9163), .A2(n5734), .ZN(n5183) );
  NAND2_X1 U6689 ( .A1(n5184), .A2(n5183), .ZN(n5185) );
  XNOR2_X1 U6690 ( .A(n5185), .B(n5799), .ZN(n5606) );
  INV_X1 U6691 ( .A(n5606), .ZN(n5607) );
  INV_X1 U6692 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6664) );
  OR2_X1 U6693 ( .A1(n5222), .A2(n6664), .ZN(n5188) );
  INV_X1 U6694 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5186) );
  OR2_X1 U6695 ( .A1(n5249), .A2(n5186), .ZN(n5187) );
  NAND2_X1 U6696 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5192) );
  NAND2_X1 U6697 ( .A1(n5359), .A2(n8855), .ZN(n5197) );
  XNOR2_X1 U6698 ( .A(n5194), .B(n5193), .ZN(n6076) );
  OR2_X1 U6699 ( .A1(n5318), .A2(n6076), .ZN(n5196) );
  INV_X1 U6700 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9971) );
  NAND2_X1 U6701 ( .A1(n6625), .A2(n5801), .ZN(n5200) );
  NAND2_X1 U6702 ( .A1(n7622), .A2(n5378), .ZN(n5199) );
  NAND2_X1 U6703 ( .A1(n5200), .A2(n5199), .ZN(n5218) );
  NAND2_X1 U6704 ( .A1(n5217), .A2(n5218), .ZN(n5216) );
  INV_X1 U6705 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5210) );
  OR2_X1 U6706 ( .A1(n5249), .A2(n5210), .ZN(n5205) );
  INV_X1 U6707 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U6708 ( .A1(n5221), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5203) );
  OR2_X1 U6709 ( .A1(n4404), .A2(n9538), .ZN(n5202) );
  NAND2_X1 U6710 ( .A1(n6634), .A2(n5801), .ZN(n5209) );
  INV_X1 U6711 ( .A(SI_0_), .ZN(n5902) );
  INV_X1 U6712 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n10127) );
  OAI21_X1 U6713 ( .B1(n5880), .B2(n5902), .A(n10127), .ZN(n5207) );
  AND2_X1 U6714 ( .A1(n5207), .A2(n5206), .ZN(n9375) );
  MUX2_X1 U6715 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9375), .S(n5191), .Z(n6626) );
  AOI22_X1 U6716 ( .A1(n6626), .A2(n5378), .B1(n5825), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5208) );
  NAND2_X1 U6717 ( .A1(n6634), .A2(n5378), .ZN(n5213) );
  NOR2_X1 U6718 ( .A1(n5776), .A2(n5210), .ZN(n5211) );
  AOI21_X1 U6719 ( .B1(n6626), .B2(n5796), .A(n5211), .ZN(n5212) );
  NAND2_X1 U6720 ( .A1(n5213), .A2(n5212), .ZN(n6453) );
  NAND2_X1 U6721 ( .A1(n5004), .A2(n6453), .ZN(n6452) );
  INV_X1 U6722 ( .A(n6453), .ZN(n5214) );
  NAND2_X1 U6723 ( .A1(n5214), .A2(n5799), .ZN(n5215) );
  NAND2_X1 U6724 ( .A1(n6452), .A2(n5215), .ZN(n6476) );
  NAND2_X1 U6725 ( .A1(n5216), .A2(n6476), .ZN(n5220) );
  INV_X1 U6726 ( .A(n5218), .ZN(n6475) );
  NAND2_X1 U6727 ( .A1(n6477), .A2(n6475), .ZN(n5219) );
  NAND2_X1 U6728 ( .A1(n5220), .A2(n5219), .ZN(n6470) );
  NAND2_X1 U6729 ( .A1(n7418), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U6730 ( .A1(n4409), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5225) );
  INV_X1 U6731 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6691) );
  OR2_X1 U6732 ( .A1(n4404), .A2(n6691), .ZN(n5224) );
  INV_X1 U6733 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6253) );
  OR2_X1 U6734 ( .A1(n5249), .A2(n6253), .ZN(n5223) );
  NAND2_X1 U6735 ( .A1(n6679), .A2(n5378), .ZN(n5239) );
  XNOR2_X1 U6736 ( .A(n5228), .B(n5227), .ZN(n6066) );
  OR2_X1 U6737 ( .A1(n5318), .A2(n6066), .ZN(n5236) );
  OR2_X1 U6738 ( .A1(n7478), .A2(n6059), .ZN(n5235) );
  NOR2_X1 U6739 ( .A1(n5229), .A2(n5464), .ZN(n5230) );
  NAND2_X1 U6740 ( .A1(n5230), .A2(P1_IR_REG_2__SCAN_IN), .ZN(n5233) );
  INV_X1 U6741 ( .A(n5230), .ZN(n5232) );
  INV_X1 U6742 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5231) );
  NAND2_X1 U6743 ( .A1(n5232), .A2(n5231), .ZN(n5254) );
  AND2_X1 U6744 ( .A1(n5233), .A2(n5254), .ZN(n6462) );
  NAND2_X1 U6745 ( .A1(n5359), .A2(n6462), .ZN(n5234) );
  INV_X1 U6746 ( .A(n6712), .ZN(n5237) );
  NAND2_X1 U6747 ( .A1(n5237), .A2(n5796), .ZN(n5238) );
  NAND2_X1 U6748 ( .A1(n6679), .A2(n5801), .ZN(n5242) );
  NAND2_X1 U6749 ( .A1(n5237), .A2(n5378), .ZN(n5241) );
  NAND2_X1 U6750 ( .A1(n5242), .A2(n5241), .ZN(n5243) );
  NAND2_X1 U6751 ( .A1(n6470), .A2(n6469), .ZN(n5247) );
  INV_X1 U6752 ( .A(n5243), .ZN(n5244) );
  NAND2_X1 U6753 ( .A1(n5245), .A2(n5244), .ZN(n5246) );
  INV_X1 U6754 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5248) );
  OR2_X1 U6755 ( .A1(n5812), .A2(n5248), .ZN(n5252) );
  INV_X1 U6756 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6257) );
  OR2_X1 U6757 ( .A1(n5249), .A2(n6257), .ZN(n5251) );
  NAND2_X1 U6758 ( .A1(n7418), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5250) );
  NAND3_X1 U6759 ( .A1(n5252), .A2(n5251), .A3(n5250), .ZN(n5253) );
  NAND2_X1 U6760 ( .A1(n5254), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5256) );
  INV_X1 U6761 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5255) );
  XNOR2_X1 U6762 ( .A(n5256), .B(n5255), .ZN(n6284) );
  OR2_X1 U6763 ( .A1(n7478), .A2(n6061), .ZN(n5260) );
  XNOR2_X1 U6764 ( .A(n5257), .B(n5258), .ZN(n6072) );
  OR2_X1 U6765 ( .A1(n5318), .A2(n6072), .ZN(n5259) );
  OAI211_X1 U6766 ( .C1(n5191), .C2(n6284), .A(n5260), .B(n5259), .ZN(n6832)
         );
  OAI22_X1 U6767 ( .A1(n6749), .A2(n5732), .B1(n9681), .B2(n5405), .ZN(n5264)
         );
  XNOR2_X1 U6768 ( .A(n5263), .B(n5264), .ZN(n6596) );
  NAND2_X1 U6769 ( .A1(n6597), .A2(n6596), .ZN(n5267) );
  INV_X1 U6770 ( .A(n5263), .ZN(n5265) );
  OR2_X1 U6771 ( .A1(n5265), .A2(n5264), .ZN(n5266) );
  NAND2_X1 U6772 ( .A1(n5267), .A2(n5266), .ZN(n6603) );
  NAND2_X1 U6773 ( .A1(n7418), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5274) );
  INV_X1 U6774 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6259) );
  OR2_X1 U6775 ( .A1(n7421), .A2(n6259), .ZN(n5273) );
  INV_X1 U6776 ( .A(n5292), .ZN(n5269) );
  INV_X1 U6777 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10006) );
  INV_X1 U6778 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U6779 ( .A1(n10006), .A2(n6599), .ZN(n5268) );
  NAND2_X1 U6780 ( .A1(n5269), .A2(n5268), .ZN(n6757) );
  OR2_X1 U6781 ( .A1(n4404), .A2(n6757), .ZN(n5272) );
  INV_X1 U6782 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5270) );
  OR2_X1 U6783 ( .A1(n5812), .A2(n5270), .ZN(n5271) );
  AND2_X1 U6784 ( .A1(n5275), .A2(n5229), .ZN(n5276) );
  NOR2_X1 U6785 ( .A1(n5276), .A2(n5464), .ZN(n5277) );
  MUX2_X1 U6786 ( .A(n5464), .B(n5277), .S(P1_IR_REG_4__SCAN_IN), .Z(n5278) );
  INV_X1 U6787 ( .A(n5278), .ZN(n5281) );
  INV_X1 U6788 ( .A(n5279), .ZN(n5280) );
  NAND2_X1 U6789 ( .A1(n5281), .A2(n5280), .ZN(n9547) );
  OR2_X1 U6790 ( .A1(n7478), .A2(n6062), .ZN(n5285) );
  XNOR2_X1 U6791 ( .A(n5282), .B(n5283), .ZN(n6068) );
  OR2_X1 U6792 ( .A1(n5318), .A2(n6068), .ZN(n5284) );
  OAI211_X1 U6793 ( .C1(n5191), .C2(n9547), .A(n5285), .B(n5284), .ZN(n6812)
         );
  INV_X1 U6794 ( .A(n6812), .ZN(n6758) );
  OAI22_X1 U6795 ( .A1(n7676), .A2(n5405), .B1(n6758), .B2(n5261), .ZN(n5286)
         );
  XNOR2_X1 U6796 ( .A(n5286), .B(n5799), .ZN(n5289) );
  OAI22_X1 U6797 ( .A1(n7676), .A2(n5732), .B1(n6758), .B2(n5405), .ZN(n5288)
         );
  XNOR2_X1 U6798 ( .A(n5289), .B(n5288), .ZN(n6604) );
  NAND2_X1 U6799 ( .A1(n5289), .A2(n5288), .ZN(n5290) );
  NAND2_X1 U6800 ( .A1(n5221), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5296) );
  INV_X1 U6801 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5291) );
  OR2_X1 U6802 ( .A1(n7421), .A2(n5291), .ZN(n5295) );
  INV_X1 U6803 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6707) );
  OR2_X1 U6804 ( .A1(n5670), .A2(n6707), .ZN(n5294) );
  OAI21_X1 U6805 ( .B1(n5292), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5306), .ZN(
        n7677) );
  OR2_X1 U6806 ( .A1(n4404), .A2(n7677), .ZN(n5293) );
  OR2_X1 U6807 ( .A1(n6748), .A2(n5732), .ZN(n5303) );
  OR2_X1 U6808 ( .A1(n5279), .A2(n5464), .ZN(n5297) );
  XNOR2_X1 U6809 ( .A(n5297), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9566) );
  INV_X1 U6810 ( .A(n9566), .ZN(n6063) );
  XNOR2_X1 U6811 ( .A(n5299), .B(n5298), .ZN(n6071) );
  OR2_X1 U6812 ( .A1(n5318), .A2(n6071), .ZN(n5301) );
  OR2_X1 U6813 ( .A1(n7478), .A2(n9979), .ZN(n5300) );
  OAI211_X1 U6814 ( .C1(n5191), .C2(n6063), .A(n5301), .B(n5300), .ZN(n9689)
         );
  NAND2_X1 U6815 ( .A1(n9689), .A2(n5378), .ZN(n5302) );
  NAND2_X1 U6816 ( .A1(n5303), .A2(n5302), .ZN(n5325) );
  INV_X1 U6817 ( .A(n5325), .ZN(n7674) );
  INV_X1 U6818 ( .A(n9689), .ZN(n7681) );
  OAI22_X1 U6819 ( .A1(n6748), .A2(n5405), .B1(n7681), .B2(n5261), .ZN(n5304)
         );
  XNOR2_X1 U6820 ( .A(n5304), .B(n4581), .ZN(n7672) );
  NAND2_X1 U6821 ( .A1(n7418), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5312) );
  INV_X1 U6822 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6262) );
  OR2_X1 U6823 ( .A1(n7421), .A2(n6262), .ZN(n5311) );
  AND2_X1 U6824 ( .A1(n5306), .A2(n5305), .ZN(n5307) );
  OR2_X1 U6825 ( .A1(n5307), .A2(n5334), .ZN(n7079) );
  OR2_X1 U6826 ( .A1(n4404), .A2(n7079), .ZN(n5310) );
  INV_X1 U6827 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5308) );
  OR2_X1 U6828 ( .A1(n5812), .A2(n5308), .ZN(n5309) );
  NAND2_X1 U6829 ( .A1(n5313), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5315) );
  XNOR2_X1 U6830 ( .A(n5315), .B(n5314), .ZN(n9580) );
  OR2_X1 U6831 ( .A1(n7478), .A2(n6064), .ZN(n5320) );
  OR2_X1 U6832 ( .A1(n5318), .A2(n6070), .ZN(n5319) );
  OAI211_X1 U6833 ( .C1(n5191), .C2(n9580), .A(n5320), .B(n5319), .ZN(n9696)
         );
  INV_X1 U6834 ( .A(n9696), .ZN(n7081) );
  OAI22_X1 U6835 ( .A1(n6943), .A2(n5405), .B1(n7081), .B2(n5261), .ZN(n5321)
         );
  XNOR2_X1 U6836 ( .A(n5321), .B(n4581), .ZN(n8801) );
  OR2_X1 U6837 ( .A1(n6943), .A2(n5732), .ZN(n5323) );
  NAND2_X1 U6838 ( .A1(n9696), .A2(n5378), .ZN(n5322) );
  NAND2_X1 U6839 ( .A1(n5323), .A2(n5322), .ZN(n8800) );
  INV_X1 U6840 ( .A(n8800), .ZN(n5326) );
  AOI22_X1 U6841 ( .A1(n7674), .A2(n7672), .B1(n8801), .B2(n5326), .ZN(n5324)
         );
  INV_X1 U6842 ( .A(n8801), .ZN(n5330) );
  INV_X1 U6843 ( .A(n7672), .ZN(n8799) );
  NAND2_X1 U6844 ( .A1(n8799), .A2(n5325), .ZN(n5327) );
  NAND2_X1 U6845 ( .A1(n5327), .A2(n5326), .ZN(n5329) );
  INV_X1 U6846 ( .A(n5327), .ZN(n5328) );
  AOI22_X1 U6847 ( .A1(n5330), .A2(n5329), .B1(n5328), .B2(n8800), .ZN(n5331)
         );
  NAND2_X1 U6848 ( .A1(n5332), .A2(n5331), .ZN(n6875) );
  NAND2_X1 U6849 ( .A1(n4409), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5339) );
  INV_X1 U6850 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5333) );
  OR2_X1 U6851 ( .A1(n7421), .A2(n5333), .ZN(n5338) );
  INV_X1 U6852 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6947) );
  OR2_X1 U6853 ( .A1(n5670), .A2(n6947), .ZN(n5337) );
  OR2_X1 U6854 ( .A1(n5334), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U6855 ( .A1(n5350), .A2(n5335), .ZN(n6946) );
  OR2_X1 U6856 ( .A1(n4404), .A2(n6946), .ZN(n5336) );
  OR2_X1 U6857 ( .A1(n5313), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U6858 ( .A1(n5360), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5340) );
  XNOR2_X1 U6859 ( .A(n5340), .B(P1_IR_REG_7__SCAN_IN), .ZN(n8878) );
  INV_X1 U6860 ( .A(n8878), .ZN(n6279) );
  XNOR2_X1 U6861 ( .A(n5342), .B(n5341), .ZN(n6075) );
  OR2_X1 U6862 ( .A1(n5318), .A2(n6075), .ZN(n5344) );
  OR2_X1 U6863 ( .A1(n7478), .A2(n6074), .ZN(n5343) );
  OAI211_X1 U6864 ( .C1(n5191), .C2(n6279), .A(n5344), .B(n5343), .ZN(n6952)
         );
  OAI22_X1 U6865 ( .A1(n7049), .A2(n5405), .B1(n9706), .B2(n5261), .ZN(n5345)
         );
  XNOR2_X1 U6866 ( .A(n5345), .B(n5799), .ZN(n5347) );
  OAI22_X1 U6867 ( .A1(n7049), .A2(n5732), .B1(n9706), .B2(n5405), .ZN(n5346)
         );
  OR2_X1 U6868 ( .A1(n5347), .A2(n5346), .ZN(n6874) );
  NAND2_X1 U6869 ( .A1(n6875), .A2(n6874), .ZN(n5348) );
  NAND2_X1 U6870 ( .A1(n5347), .A2(n5346), .ZN(n6873) );
  NAND2_X1 U6871 ( .A1(n7418), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5356) );
  INV_X1 U6872 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6266) );
  OR2_X1 U6873 ( .A1(n7421), .A2(n6266), .ZN(n5355) );
  NAND2_X1 U6874 ( .A1(n5350), .A2(n5349), .ZN(n5351) );
  NAND2_X1 U6875 ( .A1(n5371), .A2(n5351), .ZN(n8716) );
  OR2_X1 U6876 ( .A1(n4404), .A2(n8716), .ZN(n5354) );
  INV_X1 U6877 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5352) );
  OR2_X1 U6878 ( .A1(n5812), .A2(n5352), .ZN(n5353) );
  XNOR2_X1 U6879 ( .A(n5358), .B(n5357), .ZN(n6770) );
  NAND2_X1 U6880 ( .A1(n6770), .A2(n7415), .ZN(n5367) );
  NOR2_X1 U6881 ( .A1(n5360), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5363) );
  NOR2_X1 U6882 ( .A1(n5363), .A2(n5464), .ZN(n5361) );
  MUX2_X1 U6883 ( .A(n5464), .B(n5361), .S(P1_IR_REG_8__SCAN_IN), .Z(n5365) );
  INV_X1 U6884 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6885 ( .A1(n5363), .A2(n5362), .ZN(n5394) );
  INV_X1 U6886 ( .A(n5394), .ZN(n5364) );
  INV_X1 U6887 ( .A(n9587), .ZN(n9600) );
  NAND2_X1 U6888 ( .A1(n5359), .A2(n9600), .ZN(n5366) );
  OAI211_X1 U6889 ( .C1(n7478), .C2(n6080), .A(n5367), .B(n5366), .ZN(n9710)
         );
  OAI22_X1 U6890 ( .A1(n7145), .A2(n5732), .B1(n7053), .B2(n5405), .ZN(n5369)
         );
  OAI22_X1 U6891 ( .A1(n7145), .A2(n5405), .B1(n7053), .B2(n5261), .ZN(n5368)
         );
  XNOR2_X1 U6892 ( .A(n5368), .B(n4581), .ZN(n8714) );
  NAND2_X1 U6893 ( .A1(n7418), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U6894 ( .A1(n5221), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5376) );
  AND2_X1 U6895 ( .A1(n5371), .A2(n5370), .ZN(n5372) );
  OR2_X1 U6896 ( .A1(n5372), .A2(n5398), .ZN(n7151) );
  OR2_X1 U6897 ( .A1(n4404), .A2(n7151), .ZN(n5375) );
  INV_X1 U6898 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5373) );
  OR2_X1 U6899 ( .A1(n7421), .A2(n5373), .ZN(n5374) );
  NAND4_X1 U6900 ( .A1(n5377), .A2(n5376), .A3(n5375), .A4(n5374), .ZN(n8841)
         );
  NAND2_X1 U6901 ( .A1(n8841), .A2(n5378), .ZN(n5384) );
  XNOR2_X1 U6902 ( .A(n5379), .B(n5002), .ZN(n6781) );
  NAND2_X1 U6903 ( .A1(n6781), .A2(n7415), .ZN(n5382) );
  NAND2_X1 U6904 ( .A1(n5394), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5380) );
  XNOR2_X1 U6905 ( .A(n5380), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6295) );
  AOI22_X1 U6906 ( .A1(n5588), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5359), .B2(
        n6295), .ZN(n5381) );
  NAND2_X1 U6907 ( .A1(n7233), .A2(n5796), .ZN(n5383) );
  NAND2_X1 U6908 ( .A1(n5384), .A2(n5383), .ZN(n5385) );
  XNOR2_X1 U6909 ( .A(n5385), .B(n4581), .ZN(n5390) );
  NAND2_X1 U6910 ( .A1(n8841), .A2(n5801), .ZN(n5387) );
  NAND2_X1 U6911 ( .A1(n7233), .A2(n5734), .ZN(n5386) );
  NAND2_X1 U6912 ( .A1(n5387), .A2(n5386), .ZN(n5388) );
  XNOR2_X1 U6913 ( .A(n5390), .B(n5388), .ZN(n7058) );
  NAND2_X1 U6914 ( .A1(n7059), .A2(n7058), .ZN(n5392) );
  INV_X1 U6915 ( .A(n5388), .ZN(n5389) );
  NAND2_X1 U6916 ( .A1(n5390), .A2(n5389), .ZN(n5391) );
  NAND2_X1 U6917 ( .A1(n6881), .A2(n7415), .ZN(n5397) );
  NAND2_X1 U6918 ( .A1(n5395), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5414) );
  XNOR2_X1 U6919 ( .A(n5414), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6323) );
  AOI22_X1 U6920 ( .A1(n5588), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5359), .B2(
        n6323), .ZN(n5396) );
  NAND2_X1 U6921 ( .A1(n8700), .A2(n5796), .ZN(n5407) );
  NAND2_X1 U6922 ( .A1(n4409), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5404) );
  INV_X1 U6923 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7241) );
  OR2_X1 U6924 ( .A1(n5670), .A2(n7241), .ZN(n5403) );
  NOR2_X1 U6925 ( .A1(n5398), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5399) );
  OR2_X1 U6926 ( .A1(n5419), .A2(n5399), .ZN(n8698) );
  OR2_X1 U6927 ( .A1(n4404), .A2(n8698), .ZN(n5402) );
  INV_X1 U6928 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5400) );
  OR2_X1 U6929 ( .A1(n7421), .A2(n5400), .ZN(n5401) );
  OR2_X1 U6930 ( .A1(n9466), .A2(n5405), .ZN(n5406) );
  NAND2_X1 U6931 ( .A1(n5407), .A2(n5406), .ZN(n5408) );
  XNOR2_X1 U6932 ( .A(n5408), .B(n4581), .ZN(n8693) );
  OR2_X1 U6933 ( .A1(n9466), .A2(n5732), .ZN(n5410) );
  NAND2_X1 U6934 ( .A1(n8700), .A2(n5734), .ZN(n5409) );
  AND2_X1 U6935 ( .A1(n5410), .A2(n5409), .ZN(n5433) );
  AND2_X1 U6936 ( .A1(n8693), .A2(n5433), .ZN(n8774) );
  XNOR2_X1 U6937 ( .A(n5412), .B(n5411), .ZN(n6910) );
  NAND2_X1 U6938 ( .A1(n6910), .A2(n7415), .ZN(n5418) );
  NAND2_X1 U6939 ( .A1(n5414), .A2(n5413), .ZN(n5415) );
  NAND2_X1 U6940 ( .A1(n5415), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5416) );
  XNOR2_X1 U6941 ( .A(n5416), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6394) );
  AOI22_X1 U6942 ( .A1(n5588), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5359), .B2(
        n6394), .ZN(n5417) );
  NAND2_X1 U6943 ( .A1(n8783), .A2(n5796), .ZN(n5426) );
  NAND2_X1 U6944 ( .A1(n5221), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U6945 ( .A1(n5697), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5423) );
  INV_X1 U6946 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9478) );
  OR2_X1 U6947 ( .A1(n5670), .A2(n9478), .ZN(n5422) );
  OR2_X1 U6948 ( .A1(n5419), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6949 ( .A1(n5446), .A2(n5420), .ZN(n9477) );
  OR2_X1 U6950 ( .A1(n4404), .A2(n9477), .ZN(n5421) );
  NAND4_X1 U6951 ( .A1(n5424), .A2(n5423), .A3(n5422), .A4(n5421), .ZN(n8839)
         );
  NAND2_X1 U6952 ( .A1(n8839), .A2(n5734), .ZN(n5425) );
  NAND2_X1 U6953 ( .A1(n5426), .A2(n5425), .ZN(n5427) );
  XNOR2_X1 U6954 ( .A(n5427), .B(n5799), .ZN(n5431) );
  AND2_X1 U6955 ( .A1(n8839), .A2(n5801), .ZN(n5428) );
  AOI21_X1 U6956 ( .B1(n8783), .B2(n5734), .A(n5428), .ZN(n5430) );
  INV_X1 U6957 ( .A(n5430), .ZN(n5429) );
  NAND2_X1 U6958 ( .A1(n5431), .A2(n5429), .ZN(n5435) );
  INV_X1 U6959 ( .A(n5435), .ZN(n5432) );
  XNOR2_X1 U6960 ( .A(n5431), .B(n5430), .ZN(n8779) );
  NOR2_X1 U6961 ( .A1(n5432), .A2(n8779), .ZN(n5437) );
  INV_X1 U6962 ( .A(n8693), .ZN(n5434) );
  INV_X1 U6963 ( .A(n5433), .ZN(n8692) );
  NAND2_X1 U6964 ( .A1(n5434), .A2(n8692), .ZN(n8776) );
  AND2_X1 U6965 ( .A1(n8776), .A2(n5435), .ZN(n5436) );
  OR2_X1 U6966 ( .A1(n5437), .A2(n5436), .ZN(n5438) );
  INV_X1 U6967 ( .A(n7260), .ZN(n5461) );
  XNOR2_X1 U6968 ( .A(n5440), .B(n5439), .ZN(n7015) );
  NAND2_X1 U6969 ( .A1(n7015), .A2(n7415), .ZN(n5444) );
  NAND2_X1 U6970 ( .A1(n5441), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5442) );
  XNOR2_X1 U6971 ( .A(n5442), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9624) );
  AOI22_X1 U6972 ( .A1(n5588), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5359), .B2(
        n9624), .ZN(n5443) );
  NAND2_X1 U6973 ( .A1(n9508), .A2(n5796), .ZN(n5454) );
  NAND2_X1 U6974 ( .A1(n7418), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5452) );
  INV_X1 U6975 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6389) );
  OR2_X1 U6976 ( .A1(n7421), .A2(n6389), .ZN(n5451) );
  NAND2_X1 U6977 ( .A1(n5446), .A2(n5445), .ZN(n5447) );
  NAND2_X1 U6978 ( .A1(n5470), .A2(n5447), .ZN(n7273) );
  OR2_X1 U6979 ( .A1(n4404), .A2(n7273), .ZN(n5450) );
  INV_X1 U6980 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5448) );
  OR2_X1 U6981 ( .A1(n5812), .A2(n5448), .ZN(n5449) );
  NAND2_X1 U6982 ( .A1(n8838), .A2(n5734), .ZN(n5453) );
  NAND2_X1 U6983 ( .A1(n5454), .A2(n5453), .ZN(n5455) );
  XNOR2_X1 U6984 ( .A(n5455), .B(n4581), .ZN(n5458) );
  NOR2_X1 U6985 ( .A1(n9468), .A2(n5732), .ZN(n5456) );
  AOI21_X1 U6986 ( .B1(n9508), .B2(n5734), .A(n5456), .ZN(n5457) );
  NAND2_X1 U6987 ( .A1(n5458), .A2(n5457), .ZN(n5462) );
  OR2_X1 U6988 ( .A1(n5458), .A2(n5457), .ZN(n5459) );
  NAND2_X1 U6989 ( .A1(n5462), .A2(n5459), .ZN(n7261) );
  XNOR2_X1 U6990 ( .A(n5463), .B(n5001), .ZN(n7095) );
  NAND2_X1 U6991 ( .A1(n7095), .A2(n7415), .ZN(n5468) );
  OR2_X1 U6992 ( .A1(n5465), .A2(n5464), .ZN(n5466) );
  XNOR2_X1 U6993 ( .A(n5466), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6539) );
  AOI22_X1 U6994 ( .A1(n5588), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5359), .B2(
        n6539), .ZN(n5467) );
  NAND2_X1 U6995 ( .A1(n9499), .A2(n5796), .ZN(n5477) );
  NAND2_X1 U6996 ( .A1(n5697), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5475) );
  NAND2_X1 U6997 ( .A1(n4409), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5474) );
  INV_X1 U6998 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7358) );
  OR2_X1 U6999 ( .A1(n5670), .A2(n7358), .ZN(n5473) );
  NAND2_X1 U7000 ( .A1(n5470), .A2(n5469), .ZN(n5471) );
  NAND2_X1 U7001 ( .A1(n5490), .A2(n5471), .ZN(n7357) );
  OR2_X1 U7002 ( .A1(n4404), .A2(n7357), .ZN(n5472) );
  NAND4_X1 U7003 ( .A1(n5475), .A2(n5474), .A3(n5473), .A4(n5472), .ZN(n9252)
         );
  NAND2_X1 U7004 ( .A1(n9252), .A2(n5734), .ZN(n5476) );
  NAND2_X1 U7005 ( .A1(n5477), .A2(n5476), .ZN(n5478) );
  XNOR2_X1 U7006 ( .A(n5478), .B(n4581), .ZN(n5480) );
  AND2_X1 U7007 ( .A1(n9252), .A2(n5801), .ZN(n5479) );
  AOI21_X1 U7008 ( .B1(n9499), .B2(n5734), .A(n5479), .ZN(n5481) );
  AND2_X1 U7009 ( .A1(n5480), .A2(n5481), .ZN(n7248) );
  INV_X1 U7010 ( .A(n5480), .ZN(n5483) );
  INV_X1 U7011 ( .A(n5481), .ZN(n5482) );
  NAND2_X1 U7012 ( .A1(n5483), .A2(n5482), .ZN(n7249) );
  XNOR2_X1 U7013 ( .A(n5485), .B(n5484), .ZN(n7208) );
  NAND2_X1 U7014 ( .A1(n7208), .A2(n7415), .ZN(n5488) );
  OR2_X1 U7015 ( .A1(n5486), .A2(n5464), .ZN(n5506) );
  XNOR2_X1 U7016 ( .A(n5506), .B(P1_IR_REG_14__SCAN_IN), .ZN(n6541) );
  AOI22_X1 U7017 ( .A1(n5588), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5359), .B2(
        n6541), .ZN(n5487) );
  NAND2_X1 U7018 ( .A1(n9265), .A2(n5796), .ZN(n5497) );
  NAND2_X1 U7019 ( .A1(n5697), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U7020 ( .A1(n5221), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5494) );
  AND2_X1 U7021 ( .A1(n5490), .A2(n5489), .ZN(n5491) );
  OR2_X1 U7022 ( .A1(n5491), .A2(n5511), .ZN(n9261) );
  OR2_X1 U7023 ( .A1(n4404), .A2(n9261), .ZN(n5493) );
  INV_X1 U7024 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9262) );
  OR2_X1 U7025 ( .A1(n5670), .A2(n9262), .ZN(n5492) );
  NAND4_X1 U7026 ( .A1(n5495), .A2(n5494), .A3(n5493), .A4(n5492), .ZN(n9229)
         );
  NAND2_X1 U7027 ( .A1(n9229), .A2(n5734), .ZN(n5496) );
  NAND2_X1 U7028 ( .A1(n5497), .A2(n5496), .ZN(n5498) );
  XNOR2_X1 U7029 ( .A(n5498), .B(n5799), .ZN(n5501) );
  NAND2_X1 U7030 ( .A1(n9265), .A2(n5734), .ZN(n5500) );
  NAND2_X1 U7031 ( .A1(n9229), .A2(n5801), .ZN(n5499) );
  NAND2_X1 U7032 ( .A1(n5500), .A2(n5499), .ZN(n7395) );
  NAND2_X1 U7033 ( .A1(n5502), .A2(n5501), .ZN(n7392) );
  XNOR2_X1 U7034 ( .A(n5504), .B(n5503), .ZN(n7367) );
  NAND2_X1 U7035 ( .A1(n7367), .A2(n7415), .ZN(n5510) );
  NAND2_X1 U7036 ( .A1(n5506), .A2(n5505), .ZN(n5507) );
  NAND2_X1 U7037 ( .A1(n5507), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5508) );
  XNOR2_X1 U7038 ( .A(n5508), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9638) );
  AOI22_X1 U7039 ( .A1(n5588), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5359), .B2(
        n9638), .ZN(n5509) );
  NAND2_X1 U7040 ( .A1(n9242), .A2(n5796), .ZN(n5519) );
  NAND2_X1 U7041 ( .A1(n4409), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5517) );
  INV_X1 U7042 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9236) );
  OR2_X1 U7043 ( .A1(n5670), .A2(n9236), .ZN(n5516) );
  OR2_X1 U7044 ( .A1(n5511), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U7045 ( .A1(n5533), .A2(n5512), .ZN(n9235) );
  OR2_X1 U7046 ( .A1(n4404), .A2(n9235), .ZN(n5515) );
  INV_X1 U7047 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5513) );
  OR2_X1 U7048 ( .A1(n7421), .A2(n5513), .ZN(n5514) );
  NAND2_X1 U7049 ( .A1(n9255), .A2(n5734), .ZN(n5518) );
  NAND2_X1 U7050 ( .A1(n5519), .A2(n5518), .ZN(n5520) );
  XNOR2_X1 U7051 ( .A(n5520), .B(n5799), .ZN(n5524) );
  NAND2_X1 U7052 ( .A1(n9242), .A2(n5734), .ZN(n5523) );
  NAND2_X1 U7053 ( .A1(n9255), .A2(n5801), .ZN(n5522) );
  NAND2_X1 U7054 ( .A1(n5523), .A2(n5522), .ZN(n8823) );
  NAND2_X1 U7055 ( .A1(n5525), .A2(n5524), .ZN(n8824) );
  XNOR2_X1 U7056 ( .A(n5527), .B(n5526), .ZN(n7687) );
  NAND2_X1 U7057 ( .A1(n7687), .A2(n7415), .ZN(n5531) );
  NAND2_X1 U7058 ( .A1(n5528), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5529) );
  XNOR2_X1 U7059 ( .A(n5529), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9652) );
  AOI22_X1 U7060 ( .A1(n5588), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5359), .B2(
        n9652), .ZN(n5530) );
  NAND2_X1 U7061 ( .A1(n9220), .A2(n5796), .ZN(n5540) );
  NAND2_X1 U7062 ( .A1(n7418), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5538) );
  OR2_X1 U7063 ( .A1(n5812), .A2(n9518), .ZN(n5537) );
  NAND2_X1 U7064 ( .A1(n5533), .A2(n5532), .ZN(n5534) );
  NAND2_X1 U7065 ( .A1(n5551), .A2(n5534), .ZN(n9215) );
  OR2_X1 U7066 ( .A1(n4404), .A2(n9215), .ZN(n5536) );
  INV_X1 U7067 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8888) );
  OR2_X1 U7068 ( .A1(n7421), .A2(n8888), .ZN(n5535) );
  NAND2_X1 U7069 ( .A1(n9230), .A2(n5734), .ZN(n5539) );
  NAND2_X1 U7070 ( .A1(n5540), .A2(n5539), .ZN(n5541) );
  XNOR2_X1 U7071 ( .A(n5541), .B(n5799), .ZN(n8736) );
  NAND2_X1 U7072 ( .A1(n9220), .A2(n5734), .ZN(n5543) );
  NAND2_X1 U7073 ( .A1(n9230), .A2(n5801), .ZN(n5542) );
  NAND2_X1 U7074 ( .A1(n5543), .A2(n5542), .ZN(n8737) );
  NAND2_X1 U7075 ( .A1(n8739), .A2(n8736), .ZN(n5544) );
  XNOR2_X1 U7076 ( .A(n5546), .B(n5545), .ZN(n7690) );
  NAND2_X1 U7077 ( .A1(n7690), .A2(n7415), .ZN(n5550) );
  INV_X1 U7078 ( .A(n5547), .ZN(n5548) );
  NAND2_X1 U7079 ( .A1(n5548), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5568) );
  XNOR2_X1 U7080 ( .A(n5568), .B(n5567), .ZN(n9667) );
  INV_X1 U7081 ( .A(n9667), .ZN(n8910) );
  AOI22_X1 U7082 ( .A1(n5588), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5359), .B2(
        n8910), .ZN(n5549) );
  NAND2_X1 U7083 ( .A1(n9342), .A2(n5796), .ZN(n5559) );
  AND2_X1 U7084 ( .A1(n5551), .A2(n10190), .ZN(n5552) );
  OR2_X1 U7085 ( .A1(n5552), .A2(n5573), .ZN(n9190) );
  OR2_X1 U7086 ( .A1(n4404), .A2(n9190), .ZN(n5557) );
  NAND2_X1 U7087 ( .A1(n7418), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5556) );
  INV_X1 U7088 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n5553) );
  OR2_X1 U7089 ( .A1(n5812), .A2(n5553), .ZN(n5555) );
  INV_X1 U7090 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8893) );
  OR2_X1 U7091 ( .A1(n7421), .A2(n8893), .ZN(n5554) );
  NAND4_X1 U7092 ( .A1(n5557), .A2(n5556), .A3(n5555), .A4(n5554), .ZN(n9206)
         );
  NAND2_X1 U7093 ( .A1(n9206), .A2(n5734), .ZN(n5558) );
  NAND2_X1 U7094 ( .A1(n5559), .A2(n5558), .ZN(n5560) );
  XNOR2_X1 U7095 ( .A(n5560), .B(n4581), .ZN(n5563) );
  AND2_X1 U7096 ( .A1(n9206), .A2(n5801), .ZN(n5561) );
  AOI21_X1 U7097 ( .B1(n9342), .B2(n5734), .A(n5561), .ZN(n5562) );
  XNOR2_X1 U7098 ( .A(n5563), .B(n5562), .ZN(n8744) );
  NAND2_X1 U7099 ( .A1(n5563), .A2(n5562), .ZN(n5564) );
  XNOR2_X1 U7100 ( .A(n5566), .B(n5565), .ZN(n7702) );
  NAND2_X1 U7101 ( .A1(n7702), .A2(n7415), .ZN(n5572) );
  NAND2_X1 U7102 ( .A1(n5568), .A2(n5567), .ZN(n5569) );
  NAND2_X1 U7103 ( .A1(n5569), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5570) );
  XNOR2_X1 U7104 ( .A(n5570), .B(P1_IR_REG_18__SCAN_IN), .ZN(n8918) );
  AOI22_X1 U7105 ( .A1(n5588), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5359), .B2(
        n8918), .ZN(n5571) );
  NAND2_X1 U7106 ( .A1(n9335), .A2(n5796), .ZN(n5580) );
  NAND2_X1 U7107 ( .A1(n5221), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5578) );
  INV_X1 U7108 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8922) );
  OR2_X1 U7109 ( .A1(n7421), .A2(n8922), .ZN(n5577) );
  NOR2_X1 U7110 ( .A1(n5573), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5574) );
  OR2_X1 U7111 ( .A1(n5591), .A2(n5574), .ZN(n9171) );
  OR2_X1 U7112 ( .A1(n9171), .A2(n4404), .ZN(n5576) );
  INV_X1 U7113 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8898) );
  OR2_X1 U7114 ( .A1(n5670), .A2(n8898), .ZN(n5575) );
  NAND2_X1 U7115 ( .A1(n9162), .A2(n5734), .ZN(n5579) );
  NAND2_X1 U7116 ( .A1(n5580), .A2(n5579), .ZN(n5581) );
  XNOR2_X1 U7117 ( .A(n5581), .B(n4581), .ZN(n5584) );
  NAND2_X1 U7118 ( .A1(n9335), .A2(n5734), .ZN(n5583) );
  NAND2_X1 U7119 ( .A1(n9162), .A2(n5801), .ZN(n5582) );
  NAND2_X1 U7120 ( .A1(n5583), .A2(n5582), .ZN(n8791) );
  XNOR2_X1 U7121 ( .A(n5587), .B(n5586), .ZN(n7713) );
  NAND2_X1 U7122 ( .A1(n7713), .A2(n7415), .ZN(n5590) );
  AOI22_X1 U7123 ( .A1(n5588), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9087), .B2(
        n5359), .ZN(n5589) );
  NAND2_X1 U7124 ( .A1(n9330), .A2(n5796), .ZN(n5599) );
  NOR2_X1 U7125 ( .A1(n5591), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5592) );
  OR2_X1 U7126 ( .A1(n5593), .A2(n5592), .ZN(n9155) );
  INV_X1 U7127 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8924) );
  OAI22_X1 U7128 ( .A1(n9155), .A2(n4404), .B1(n7421), .B2(n8924), .ZN(n5597)
         );
  INV_X1 U7129 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7130 ( .A1(n4409), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5594) );
  OAI21_X1 U7131 ( .B1(n5595), .B2(n5670), .A(n5594), .ZN(n5596) );
  NAND2_X1 U7132 ( .A1(n9181), .A2(n5734), .ZN(n5598) );
  NAND2_X1 U7133 ( .A1(n5599), .A2(n5598), .ZN(n5600) );
  XNOR2_X1 U7134 ( .A(n5600), .B(n5799), .ZN(n5604) );
  NAND2_X1 U7135 ( .A1(n9330), .A2(n5734), .ZN(n5602) );
  NAND2_X1 U7136 ( .A1(n9181), .A2(n5801), .ZN(n5601) );
  NAND2_X1 U7137 ( .A1(n5602), .A2(n5601), .ZN(n5603) );
  NAND2_X1 U7138 ( .A1(n5604), .A2(n5603), .ZN(n8705) );
  XNOR2_X1 U7139 ( .A(n5606), .B(n5605), .ZN(n8758) );
  XNOR2_X1 U7140 ( .A(n5610), .B(n5609), .ZN(n7730) );
  NAND2_X1 U7141 ( .A1(n7730), .A2(n7415), .ZN(n5613) );
  OR2_X1 U7142 ( .A1(n7478), .A2(n5611), .ZN(n5612) );
  NAND2_X1 U7143 ( .A1(n7418), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5621) );
  INV_X1 U7144 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9973) );
  OR2_X1 U7145 ( .A1(n5812), .A2(n9973), .ZN(n5620) );
  INV_X1 U7146 ( .A(n5614), .ZN(n5616) );
  OAI21_X1 U7147 ( .B1(P1_REG3_REG_21__SCAN_IN), .B2(n5616), .A(n5615), .ZN(
        n9132) );
  OR2_X1 U7148 ( .A1(n4404), .A2(n9132), .ZN(n5619) );
  INV_X1 U7149 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5617) );
  OR2_X1 U7150 ( .A1(n7421), .A2(n5617), .ZN(n5618) );
  AOI22_X1 U7151 ( .A1(n9322), .A2(n5734), .B1(n5801), .B2(n9142), .ZN(n5625)
         );
  NAND2_X1 U7152 ( .A1(n9322), .A2(n5796), .ZN(n5623) );
  NAND2_X1 U7153 ( .A1(n9142), .A2(n5734), .ZN(n5622) );
  NAND2_X1 U7154 ( .A1(n5623), .A2(n5622), .ZN(n5624) );
  XNOR2_X1 U7155 ( .A(n5624), .B(n5799), .ZN(n5627) );
  XOR2_X1 U7156 ( .A(n5625), .B(n5627), .Z(n8722) );
  INV_X1 U7157 ( .A(n5625), .ZN(n5626) );
  XNOR2_X1 U7158 ( .A(n5629), .B(n5628), .ZN(n7733) );
  NAND2_X1 U7159 ( .A1(n7733), .A2(n7415), .ZN(n5631) );
  OR2_X1 U7160 ( .A1(n7478), .A2(n7129), .ZN(n5630) );
  NAND2_X1 U7161 ( .A1(n5697), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5638) );
  INV_X1 U7162 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9114) );
  OR2_X1 U7163 ( .A1(n5670), .A2(n9114), .ZN(n5637) );
  INV_X1 U7164 ( .A(n5647), .ZN(n5632) );
  OAI21_X1 U7165 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n5633), .A(n5632), .ZN(
        n9113) );
  OR2_X1 U7166 ( .A1(n4404), .A2(n9113), .ZN(n5636) );
  INV_X1 U7167 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n5634) );
  OR2_X1 U7168 ( .A1(n5812), .A2(n5634), .ZN(n5635) );
  AOI22_X1 U7169 ( .A1(n9317), .A2(n5734), .B1(n5801), .B2(n9107), .ZN(n5640)
         );
  NAND2_X1 U7170 ( .A1(n5641), .A2(n5640), .ZN(n8765) );
  OAI22_X1 U7171 ( .A1(n9112), .A2(n5261), .B1(n9130), .B2(n5405), .ZN(n5639)
         );
  XNOR2_X1 U7172 ( .A(n5639), .B(n5799), .ZN(n8767) );
  NOR2_X1 U7173 ( .A1(n5641), .A2(n5640), .ZN(n8766) );
  NAND2_X1 U7174 ( .A1(n7740), .A2(n7415), .ZN(n5645) );
  OR2_X1 U7175 ( .A1(n7478), .A2(n7179), .ZN(n5644) );
  NAND2_X1 U7176 ( .A1(n5221), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5652) );
  NAND2_X1 U7177 ( .A1(n5697), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5651) );
  OAI21_X1 U7178 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n5647), .A(n5646), .ZN(
        n9097) );
  OR2_X1 U7179 ( .A1(n4404), .A2(n9097), .ZN(n5650) );
  INV_X1 U7180 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5648) );
  OR2_X1 U7181 ( .A1(n5670), .A2(n5648), .ZN(n5649) );
  NAND4_X1 U7182 ( .A1(n5652), .A2(n5651), .A3(n5650), .A4(n5649), .ZN(n8837)
         );
  OAI22_X1 U7183 ( .A1(n9100), .A2(n5261), .B1(n9121), .B2(n5405), .ZN(n5653)
         );
  XOR2_X1 U7184 ( .A(n5799), .B(n5653), .Z(n5654) );
  OAI22_X1 U7185 ( .A1(n9100), .A2(n5405), .B1(n9121), .B2(n5732), .ZN(n8685)
         );
  XOR2_X1 U7186 ( .A(n5656), .B(n5655), .Z(n8752) );
  OAI21_X1 U7187 ( .B1(n5658), .B2(n5657), .A(n8750), .ZN(n8729) );
  INV_X1 U7188 ( .A(n5659), .ZN(n5662) );
  NAND2_X1 U7189 ( .A1(n5660), .A2(SI_24_), .ZN(n5661) );
  INV_X1 U7190 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7343) );
  MUX2_X1 U7191 ( .A(n7343), .B(n7344), .S(n7428), .Z(n5665) );
  INV_X1 U7192 ( .A(SI_25_), .ZN(n5664) );
  NAND2_X1 U7193 ( .A1(n5665), .A2(n5664), .ZN(n5685) );
  INV_X1 U7194 ( .A(n5665), .ZN(n5666) );
  NAND2_X1 U7195 ( .A1(n5666), .A2(SI_25_), .ZN(n5667) );
  NAND2_X1 U7196 ( .A1(n5685), .A2(n5667), .ZN(n5686) );
  NAND2_X1 U7197 ( .A1(n7763), .A2(n7415), .ZN(n5669) );
  OR2_X1 U7198 ( .A1(n7478), .A2(n7344), .ZN(n5668) );
  NAND2_X1 U7199 ( .A1(n9302), .A2(n5796), .ZN(n5680) );
  NAND2_X1 U7200 ( .A1(n5697), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5678) );
  INV_X1 U7201 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9069) );
  OR2_X1 U7202 ( .A1(n5670), .A2(n9069), .ZN(n5677) );
  INV_X1 U7203 ( .A(n5672), .ZN(n5671) );
  NAND2_X1 U7204 ( .A1(n5671), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5699) );
  INV_X1 U7205 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U7206 ( .A1(n5672), .A2(n8731), .ZN(n5673) );
  NAND2_X1 U7207 ( .A1(n5699), .A2(n5673), .ZN(n9068) );
  OR2_X1 U7208 ( .A1(n4404), .A2(n9068), .ZN(n5676) );
  INV_X1 U7209 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n5674) );
  OR2_X1 U7210 ( .A1(n5812), .A2(n5674), .ZN(n5675) );
  NAND2_X1 U7211 ( .A1(n8962), .A2(n5734), .ZN(n5679) );
  NAND2_X1 U7212 ( .A1(n5680), .A2(n5679), .ZN(n5681) );
  XNOR2_X1 U7213 ( .A(n5681), .B(n5799), .ZN(n5682) );
  AOI22_X1 U7214 ( .A1(n9302), .A2(n5734), .B1(n5801), .B2(n8962), .ZN(n5683)
         );
  XNOR2_X1 U7215 ( .A(n5682), .B(n5683), .ZN(n8730) );
  INV_X1 U7216 ( .A(n5682), .ZN(n5684) );
  AOI22_X1 U7217 ( .A1(n8729), .A2(n8730), .B1(n5684), .B2(n5683), .ZN(n8815)
         );
  INV_X1 U7218 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7388) );
  INV_X1 U7219 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7389) );
  MUX2_X1 U7220 ( .A(n7388), .B(n7389), .S(n7411), .Z(n5689) );
  INV_X1 U7221 ( .A(SI_26_), .ZN(n5688) );
  NAND2_X1 U7222 ( .A1(n5689), .A2(n5688), .ZN(n5713) );
  INV_X1 U7223 ( .A(n5689), .ZN(n5690) );
  NAND2_X1 U7224 ( .A1(n5690), .A2(SI_26_), .ZN(n5691) );
  OR2_X1 U7225 ( .A1(n5693), .A2(n5692), .ZN(n5694) );
  NAND2_X1 U7226 ( .A1(n5714), .A2(n5694), .ZN(n7775) );
  NAND2_X1 U7227 ( .A1(n7775), .A2(n7415), .ZN(n5696) );
  OR2_X1 U7228 ( .A1(n7478), .A2(n7389), .ZN(n5695) );
  NAND2_X1 U7229 ( .A1(n5697), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U7230 ( .A1(n7418), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5704) );
  INV_X1 U7231 ( .A(n5699), .ZN(n5698) );
  INV_X1 U7232 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9965) );
  NAND2_X1 U7233 ( .A1(n5699), .A2(n9965), .ZN(n5700) );
  NAND2_X1 U7234 ( .A1(n5761), .A2(n5700), .ZN(n9056) );
  OR2_X1 U7235 ( .A1(n4404), .A2(n9056), .ZN(n5703) );
  INV_X1 U7236 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n5701) );
  OR2_X1 U7237 ( .A1(n5812), .A2(n5701), .ZN(n5702) );
  NAND4_X1 U7238 ( .A1(n5705), .A2(n5704), .A3(n5703), .A4(n5702), .ZN(n9044)
         );
  OAI22_X1 U7239 ( .A1(n9060), .A2(n5405), .B1(n9076), .B2(n5732), .ZN(n5710)
         );
  NAND2_X1 U7240 ( .A1(n9297), .A2(n5796), .ZN(n5707) );
  NAND2_X1 U7241 ( .A1(n9044), .A2(n5734), .ZN(n5706) );
  NAND2_X1 U7242 ( .A1(n5707), .A2(n5706), .ZN(n5708) );
  XNOR2_X1 U7243 ( .A(n5708), .B(n5799), .ZN(n5709) );
  XOR2_X1 U7244 ( .A(n5710), .B(n5709), .Z(n8814) );
  NAND2_X1 U7245 ( .A1(n8815), .A2(n8814), .ZN(n8813) );
  INV_X1 U7246 ( .A(n5709), .ZN(n5712) );
  INV_X1 U7247 ( .A(n5710), .ZN(n5711) );
  INV_X1 U7248 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5715) );
  INV_X1 U7249 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5722) );
  INV_X1 U7250 ( .A(SI_27_), .ZN(n9999) );
  NAND2_X1 U7251 ( .A1(n5716), .A2(n9999), .ZN(n5792) );
  INV_X1 U7252 ( .A(n5716), .ZN(n5717) );
  NAND2_X1 U7253 ( .A1(n5717), .A2(SI_27_), .ZN(n5718) );
  OR2_X1 U7254 ( .A1(n5720), .A2(n5719), .ZN(n5721) );
  NAND2_X1 U7255 ( .A1(n5793), .A2(n5721), .ZN(n7788) );
  NAND2_X1 U7256 ( .A1(n7788), .A2(n7415), .ZN(n5724) );
  OR2_X1 U7257 ( .A1(n7478), .A2(n5722), .ZN(n5723) );
  NAND2_X1 U7258 ( .A1(n7418), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5730) );
  INV_X1 U7259 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5725) );
  OR2_X1 U7260 ( .A1(n7421), .A2(n5725), .ZN(n5729) );
  INV_X1 U7261 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5783) );
  XNOR2_X1 U7262 ( .A(n5761), .B(n5783), .ZN(n5780) );
  OR2_X1 U7263 ( .A1(n4404), .A2(n5780), .ZN(n5728) );
  INV_X1 U7264 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n5726) );
  OR2_X1 U7265 ( .A1(n5812), .A2(n5726), .ZN(n5727) );
  OAI22_X1 U7266 ( .A1(n9036), .A2(n5261), .B1(n9053), .B2(n5405), .ZN(n5731)
         );
  XNOR2_X1 U7267 ( .A(n5731), .B(n5799), .ZN(n5805) );
  NOR2_X1 U7268 ( .A1(n9053), .A2(n5732), .ZN(n5733) );
  AOI21_X1 U7269 ( .B1(n9291), .B2(n5734), .A(n5733), .ZN(n5789) );
  XNOR2_X1 U7270 ( .A(n5805), .B(n5789), .ZN(n5735) );
  XNOR2_X1 U7271 ( .A(n5791), .B(n5735), .ZN(n5788) );
  NAND2_X1 U7272 ( .A1(n5170), .A2(n7612), .ZN(n6635) );
  OR2_X1 U7273 ( .A1(n6635), .A2(n7013), .ZN(n6673) );
  OR2_X1 U7274 ( .A1(n6635), .A2(n8929), .ZN(n5737) );
  NAND2_X1 U7275 ( .A1(n5739), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5740) );
  XNOR2_X1 U7276 ( .A(n5740), .B(n4719), .ZN(n5826) );
  AND2_X1 U7277 ( .A1(n5826), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5741) );
  NAND2_X1 U7278 ( .A1(n7610), .A2(n9678), .ZN(n5742) );
  NOR2_X1 U7279 ( .A1(n9709), .A2(n5742), .ZN(n5760) );
  NAND2_X1 U7280 ( .A1(n7346), .A2(P1_B_REG_SCAN_IN), .ZN(n5744) );
  INV_X1 U7281 ( .A(n7232), .ZN(n5743) );
  MUX2_X1 U7282 ( .A(n5744), .B(P1_B_REG_SCAN_IN), .S(n5743), .Z(n5746) );
  NAND2_X1 U7283 ( .A1(n7391), .A2(n7346), .ZN(n5747) );
  OAI21_X1 U7284 ( .B1(n9677), .B2(P1_D_REG_1__SCAN_IN), .A(n5747), .ZN(n6331)
         );
  INV_X1 U7285 ( .A(n6331), .ZN(n9361) );
  INV_X1 U7286 ( .A(n9677), .ZN(n5758) );
  NOR4_X1 U7287 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n5756) );
  NOR4_X1 U7288 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5755) );
  INV_X1 U7289 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n9967) );
  INV_X1 U7290 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9983) );
  INV_X1 U7291 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10007) );
  INV_X1 U7292 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10054) );
  NAND4_X1 U7293 ( .A1(n9967), .A2(n9983), .A3(n10007), .A4(n10054), .ZN(n5753) );
  NOR4_X1 U7294 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5751) );
  NOR4_X1 U7295 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n5750) );
  NOR4_X1 U7296 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5749) );
  NOR4_X1 U7297 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5748) );
  NAND4_X1 U7298 ( .A1(n5751), .A2(n5750), .A3(n5749), .A4(n5748), .ZN(n5752)
         );
  NOR4_X1 U7299 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5753), .A4(n5752), .ZN(n5754) );
  NAND3_X1 U7300 ( .A1(n5756), .A2(n5755), .A3(n5754), .ZN(n5757) );
  NAND2_X1 U7301 ( .A1(n5758), .A2(n5757), .ZN(n6330) );
  NAND2_X1 U7302 ( .A1(n9361), .A2(n6330), .ZN(n6669) );
  NAND2_X1 U7303 ( .A1(n7391), .A2(n7232), .ZN(n5759) );
  OR2_X1 U7304 ( .A1(n6669), .A2(n6948), .ZN(n5775) );
  INV_X1 U7305 ( .A(n5775), .ZN(n5772) );
  NAND2_X1 U7306 ( .A1(n7418), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5769) );
  INV_X1 U7307 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10103) );
  OR2_X1 U7308 ( .A1(n7421), .A2(n10103), .ZN(n5768) );
  INV_X1 U7309 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5817) );
  OAI21_X1 U7310 ( .B1(n5761), .B2(n5783), .A(n5817), .ZN(n5764) );
  INV_X1 U7311 ( .A(n5761), .ZN(n5763) );
  AND2_X1 U7312 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5762) );
  NAND2_X1 U7313 ( .A1(n5763), .A2(n5762), .ZN(n9002) );
  NAND2_X1 U7314 ( .A1(n5764), .A2(n9002), .ZN(n9023) );
  OR2_X1 U7315 ( .A1(n4404), .A2(n9023), .ZN(n5767) );
  INV_X1 U7316 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5765) );
  OR2_X1 U7317 ( .A1(n5812), .A2(n5765), .ZN(n5766) );
  INV_X1 U7318 ( .A(n9678), .ZN(n5770) );
  NOR2_X1 U7319 ( .A1(n6721), .A2(n5770), .ZN(n5771) );
  NAND2_X1 U7320 ( .A1(n5772), .A2(n5771), .ZN(n5782) );
  NAND2_X1 U7321 ( .A1(n9686), .A2(n7612), .ZN(n5774) );
  OR2_X1 U7322 ( .A1(n7610), .A2(n7668), .ZN(n5777) );
  NAND2_X1 U7323 ( .A1(n6336), .A2(n5775), .ZN(n5786) );
  NAND3_X1 U7324 ( .A1(n5777), .A2(n5776), .A3(n5826), .ZN(n5778) );
  NAND2_X1 U7325 ( .A1(n5778), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5779) );
  NAND2_X1 U7326 ( .A1(n5786), .A2(n5779), .ZN(n8806) );
  INV_X1 U7327 ( .A(n5780), .ZN(n9034) );
  NAND2_X1 U7328 ( .A1(n8806), .A2(n9034), .ZN(n5781) );
  OAI21_X1 U7329 ( .B1(n9037), .B2(n8830), .A(n5781), .ZN(n5785) );
  OAI22_X1 U7330 ( .A1(n8816), .A2(n9076), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5783), .ZN(n5784) );
  OAI21_X1 U7331 ( .B1(n5788), .B2(n8825), .A(n5787), .ZN(P1_U3212) );
  INV_X1 U7332 ( .A(n5789), .ZN(n5804) );
  INV_X1 U7333 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7403) );
  INV_X1 U7334 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8084) );
  MUX2_X1 U7335 ( .A(n7403), .B(n8084), .S(n7411), .Z(n7408) );
  XNOR2_X1 U7336 ( .A(n7408), .B(SI_28_), .ZN(n7405) );
  NAND2_X1 U7337 ( .A1(n7792), .A2(n7415), .ZN(n5795) );
  OR2_X1 U7338 ( .A1(n7478), .A2(n8084), .ZN(n5794) );
  NAND2_X1 U7339 ( .A1(n9285), .A2(n5796), .ZN(n5798) );
  NAND2_X1 U7340 ( .A1(n8966), .A2(n5734), .ZN(n5797) );
  NAND2_X1 U7341 ( .A1(n5798), .A2(n5797), .ZN(n5800) );
  XNOR2_X1 U7342 ( .A(n5800), .B(n5799), .ZN(n5803) );
  AOI22_X1 U7343 ( .A1(n9285), .A2(n5734), .B1(n5801), .B2(n8966), .ZN(n5802)
         );
  XNOR2_X1 U7344 ( .A(n5803), .B(n5802), .ZN(n5806) );
  NAND2_X1 U7345 ( .A1(n5805), .A2(n5804), .ZN(n5807) );
  INV_X1 U7346 ( .A(n5806), .ZN(n5809) );
  INV_X1 U7347 ( .A(n5807), .ZN(n5808) );
  NAND3_X1 U7348 ( .A1(n5809), .A2(n5808), .A3(n8812), .ZN(n5821) );
  NAND2_X1 U7349 ( .A1(n7418), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5816) );
  INV_X1 U7350 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5810) );
  OR2_X1 U7351 ( .A1(n7421), .A2(n5810), .ZN(n5815) );
  OR2_X1 U7352 ( .A1(n4404), .A2(n9002), .ZN(n5814) );
  INV_X1 U7353 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5811) );
  OR2_X1 U7354 ( .A1(n5812), .A2(n5811), .ZN(n5813) );
  OAI22_X1 U7355 ( .A1(n8830), .A2(n9013), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5817), .ZN(n5819) );
  OAI22_X1 U7356 ( .A1(n8831), .A2(n9023), .B1(n9053), .B2(n8816), .ZN(n5818)
         );
  AOI211_X1 U7357 ( .C1(n9285), .C2(n8819), .A(n5819), .B(n5818), .ZN(n5820)
         );
  NAND2_X1 U7358 ( .A1(n5821), .A2(n5820), .ZN(n5822) );
  NAND2_X1 U7359 ( .A1(n5825), .A2(n5826), .ZN(n6275) );
  OR2_X2 U7360 ( .A1(n6275), .A2(P1_U3084), .ZN(n8846) );
  INV_X1 U7361 ( .A(n5826), .ZN(n7177) );
  OR2_X1 U7362 ( .A1(n7610), .A2(n7177), .ZN(n5827) );
  NAND2_X1 U7363 ( .A1(n5827), .A2(n6275), .ZN(n6273) );
  OAI21_X1 U7364 ( .B1(n6273), .B2(n5359), .A(P1_STATE_REG_SCAN_IN), .ZN(
        P1_U3083) );
  NOR2_X1 U7365 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5831) );
  AND4_X2 U7366 ( .A1(n6226), .A2(n6436), .A3(n6134), .A4(n5833), .ZN(n5834)
         );
  NAND2_X1 U7367 ( .A1(n5856), .A2(n5855), .ZN(n5839) );
  INV_X1 U7368 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U7369 ( .A1(n5854), .A2(n5840), .ZN(n5841) );
  NAND2_X1 U7370 ( .A1(n5841), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5843) );
  INV_X1 U7371 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5842) );
  NOR2_X1 U7372 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5847) );
  NOR2_X1 U7373 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n5846) );
  NOR2_X1 U7374 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5845) );
  NOR2_X1 U7375 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5844) );
  NAND4_X1 U7376 ( .A1(n5847), .A2(n5846), .A3(n5845), .A4(n5844), .ZN(n5848)
         );
  NAND2_X1 U7377 ( .A1(n5869), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5851) );
  OR2_X1 U7378 ( .A1(n5852), .A2(n5992), .ZN(n5853) );
  XNOR2_X1 U7379 ( .A(n5853), .B(P2_IR_REG_25__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7380 ( .A1(n5857), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5859) );
  XNOR2_X2 U7381 ( .A(n5859), .B(n5858), .ZN(n7994) );
  NAND2_X1 U7382 ( .A1(n5860), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U7383 ( .A1(n5862), .A2(n5861), .ZN(n5865) );
  OR2_X1 U7384 ( .A1(n5862), .A2(n5861), .ZN(n5863) );
  NAND2_X1 U7385 ( .A1(n5865), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U7386 ( .A1(n7992), .A2(n7833), .ZN(n6486) );
  INV_X1 U7387 ( .A(n5885), .ZN(n5873) );
  INV_X1 U7388 ( .A(n5878), .ZN(n5879) );
  INV_X1 U7389 ( .A(n6164), .ZN(n9381) );
  NAND2_X1 U7390 ( .A1(n7714), .A2(n9381), .ZN(n5883) );
  INV_X1 U7392 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10182) );
  AND3_X2 U7393 ( .A1(n5883), .A2(n5882), .A3(n5881), .ZN(n9758) );
  XNOR2_X2 U7394 ( .A(n5884), .B(n8676), .ZN(n5888) );
  XNOR2_X2 U7395 ( .A(n5887), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5889) );
  NAND2_X1 U7396 ( .A1(n4401), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5895) );
  NAND2_X4 U7397 ( .A1(n5888), .A2(n5889), .ZN(n7802) );
  INV_X1 U7398 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7399 ( .A1(n4406), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5894) );
  INV_X1 U7400 ( .A(n5888), .ZN(n5890) );
  INV_X1 U7401 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6165) );
  OR2_X1 U7402 ( .A1(n7032), .A2(n6165), .ZN(n5893) );
  INV_X1 U7403 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n5891) );
  OR2_X1 U7404 ( .A1(n7746), .A2(n5891), .ZN(n5892) );
  NAND4_X2 U7405 ( .A1(n5895), .A2(n5894), .A3(n5893), .A4(n5892), .ZN(n6505)
         );
  INV_X1 U7406 ( .A(n5905), .ZN(n5919) );
  NAND2_X1 U7407 ( .A1(n6505), .A2(n5919), .ZN(n5907) );
  XNOR2_X1 U7408 ( .A(n8014), .B(n5907), .ZN(n6380) );
  INV_X1 U7409 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5896) );
  OR2_X1 U7410 ( .A1(n7032), .A2(n5896), .ZN(n5901) );
  INV_X1 U7411 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6245) );
  OR2_X1 U7412 ( .A1(n7746), .A2(n6245), .ZN(n5900) );
  NAND2_X1 U7413 ( .A1(n7799), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5899) );
  INV_X1 U7414 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5897) );
  NOR2_X1 U7415 ( .A1(n7428), .A2(n5902), .ZN(n5904) );
  INV_X1 U7416 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5903) );
  XNOR2_X1 U7417 ( .A(n5904), .B(n5903), .ZN(n8684) );
  MUX2_X1 U7418 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8684), .S(n6143), .Z(n9779) );
  NAND2_X1 U7419 ( .A1(n9759), .A2(n5934), .ZN(n5906) );
  AND2_X2 U7420 ( .A1(n6248), .A2(n5906), .ZN(n6381) );
  INV_X1 U7421 ( .A(n8014), .ZN(n5908) );
  NAND2_X1 U7422 ( .A1(n5908), .A2(n5907), .ZN(n5909) );
  NAND2_X1 U7423 ( .A1(n6379), .A2(n5909), .ZN(n5920) );
  OR2_X1 U7424 ( .A1(n6769), .A2(n6066), .ZN(n5913) );
  OR2_X1 U7425 ( .A1(n7810), .A2(n6067), .ZN(n5912) );
  OR2_X1 U7426 ( .A1(n5878), .A2(n5992), .ZN(n5910) );
  XNOR2_X1 U7427 ( .A(n5910), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9394) );
  NAND2_X1 U7428 ( .A1(n7714), .A2(n9394), .ZN(n5911) );
  XNOR2_X1 U7429 ( .A(n9789), .B(n5934), .ZN(n5921) );
  INV_X1 U7430 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5914) );
  INV_X1 U7431 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6146) );
  BUF_X2 U7432 ( .A(n5919), .Z(n8092) );
  NAND2_X1 U7433 ( .A1(n6506), .A2(n8092), .ZN(n5922) );
  XNOR2_X1 U7434 ( .A(n5921), .B(n5922), .ZN(n8015) );
  NAND2_X1 U7435 ( .A1(n5920), .A2(n8015), .ZN(n8022) );
  INV_X1 U7436 ( .A(n5921), .ZN(n5923) );
  NAND2_X1 U7437 ( .A1(n5923), .A2(n5922), .ZN(n5924) );
  INV_X1 U7438 ( .A(n6343), .ZN(n5940) );
  NAND2_X1 U7439 ( .A1(n4401), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5928) );
  OR2_X1 U7440 ( .A1(n7746), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5927) );
  INV_X1 U7441 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6169) );
  OR2_X1 U7442 ( .A1(n7032), .A2(n6169), .ZN(n5926) );
  INV_X1 U7443 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6145) );
  OR2_X1 U7444 ( .A1(n7802), .A2(n6145), .ZN(n5925) );
  AND2_X1 U7445 ( .A1(n8284), .A2(n8092), .ZN(n5936) );
  OR2_X1 U7446 ( .A1(n6769), .A2(n6072), .ZN(n5933) );
  OR2_X1 U7447 ( .A1(n7810), .A2(n6073), .ZN(n5932) );
  OR3_X1 U7448 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U7449 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5929), .ZN(n5930) );
  XNOR2_X1 U7450 ( .A(n5930), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7451 ( .A1(n7714), .A2(n6168), .ZN(n5931) );
  NAND2_X1 U7452 ( .A1(n5936), .A2(n5935), .ZN(n5950) );
  INV_X1 U7453 ( .A(n5935), .ZN(n8213) );
  INV_X1 U7454 ( .A(n5936), .ZN(n5937) );
  NAND2_X1 U7455 ( .A1(n8213), .A2(n5937), .ZN(n5938) );
  NAND2_X1 U7456 ( .A1(n5950), .A2(n5938), .ZN(n6344) );
  OR2_X1 U7457 ( .A1(n6769), .A2(n6068), .ZN(n5945) );
  OR2_X1 U7458 ( .A1(n7810), .A2(n6069), .ZN(n5944) );
  OR2_X1 U7459 ( .A1(n5941), .A2(n5992), .ZN(n5942) );
  XNOR2_X1 U7460 ( .A(n5942), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7461 ( .A1(n7714), .A2(n6239), .ZN(n5943) );
  XNOR2_X1 U7462 ( .A(n9803), .B(n5934), .ZN(n5952) );
  INV_X1 U7463 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5946) );
  OR2_X1 U7464 ( .A1(n7783), .A2(n5946), .ZN(n5949) );
  NAND2_X1 U7465 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5958) );
  OAI21_X1 U7466 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5958), .ZN(n8210) );
  OR2_X1 U7467 ( .A1(n7768), .A2(n8210), .ZN(n5948) );
  INV_X1 U7468 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6171) );
  NOR2_X1 U7469 ( .A1(n4998), .A2(n4441), .ZN(n5947) );
  NAND2_X1 U7470 ( .A1(n8283), .A2(n8092), .ZN(n5953) );
  XNOR2_X1 U7471 ( .A(n5952), .B(n5953), .ZN(n8214) );
  AND2_X1 U7472 ( .A1(n8214), .A2(n5950), .ZN(n5951) );
  INV_X1 U7473 ( .A(n5952), .ZN(n5954) );
  NAND2_X1 U7474 ( .A1(n5954), .A2(n5953), .ZN(n5955) );
  NAND2_X1 U7475 ( .A1(n4401), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5963) );
  INV_X1 U7476 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5956) );
  OR2_X1 U7477 ( .A1(n7802), .A2(n5956), .ZN(n5962) );
  INV_X1 U7478 ( .A(n5958), .ZN(n5957) );
  NAND2_X1 U7479 ( .A1(n5957), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5976) );
  INV_X1 U7480 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10132) );
  NAND2_X1 U7481 ( .A1(n5958), .A2(n10132), .ZN(n5959) );
  NAND2_X1 U7482 ( .A1(n5976), .A2(n5959), .ZN(n6585) );
  OR2_X1 U7483 ( .A1(n7768), .A2(n6585), .ZN(n5961) );
  INV_X1 U7484 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6586) );
  OR2_X1 U7485 ( .A1(n7771), .A2(n6586), .ZN(n5960) );
  NAND4_X1 U7486 ( .A1(n5963), .A2(n5962), .A3(n5961), .A4(n5960), .ZN(n8282)
         );
  AND2_X1 U7487 ( .A1(n8282), .A2(n8092), .ZN(n5965) );
  INV_X1 U7488 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U7489 ( .A1(n5941), .A2(n5964), .ZN(n5991) );
  NAND2_X1 U7490 ( .A1(n5991), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5969) );
  XNOR2_X1 U7491 ( .A(n5969), .B(n5989), .ZN(n6205) );
  INV_X2 U7492 ( .A(n5934), .ZN(n8114) );
  XNOR2_X1 U7493 ( .A(n6643), .B(n8114), .ZN(n5966) );
  NAND2_X1 U7494 ( .A1(n5965), .A2(n5966), .ZN(n5982) );
  INV_X1 U7495 ( .A(n5965), .ZN(n5967) );
  INV_X1 U7496 ( .A(n5966), .ZN(n6426) );
  NAND2_X1 U7497 ( .A1(n5967), .A2(n6426), .ZN(n5968) );
  AND2_X1 U7498 ( .A1(n5982), .A2(n5968), .ZN(n6349) );
  NAND2_X1 U7499 ( .A1(n5969), .A2(n5989), .ZN(n5970) );
  NAND2_X1 U7500 ( .A1(n5970), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5971) );
  XNOR2_X1 U7501 ( .A(n5971), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6207) );
  AOI22_X1 U7502 ( .A1(n7703), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7714), .B2(
        n6207), .ZN(n5972) );
  XNOR2_X1 U7503 ( .A(n9808), .B(n5934), .ZN(n5984) );
  NAND2_X1 U7504 ( .A1(n4401), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5981) );
  INV_X1 U7505 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6208) );
  OR2_X1 U7506 ( .A1(n7802), .A2(n6208), .ZN(n5980) );
  INV_X1 U7507 ( .A(n5976), .ZN(n5974) );
  NAND2_X1 U7508 ( .A1(n5974), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6001) );
  INV_X1 U7509 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U7510 ( .A1(n5976), .A2(n5975), .ZN(n5977) );
  NAND2_X1 U7511 ( .A1(n6001), .A2(n5977), .ZN(n6654) );
  OR2_X1 U7512 ( .A1(n7768), .A2(n6654), .ZN(n5979) );
  INV_X1 U7513 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6172) );
  OR2_X1 U7514 ( .A1(n7771), .A2(n6172), .ZN(n5978) );
  NAND4_X1 U7515 ( .A1(n5981), .A2(n5980), .A3(n5979), .A4(n5978), .ZN(n8281)
         );
  NAND2_X1 U7516 ( .A1(n8281), .A2(n8092), .ZN(n5985) );
  XNOR2_X1 U7517 ( .A(n5984), .B(n5985), .ZN(n6427) );
  AND2_X1 U7518 ( .A1(n6427), .A2(n5982), .ZN(n5983) );
  INV_X1 U7519 ( .A(n5984), .ZN(n5986) );
  NAND2_X1 U7520 ( .A1(n5986), .A2(n5985), .ZN(n5987) );
  OR2_X1 U7521 ( .A1(n6075), .A2(n6769), .ZN(n5998) );
  INV_X1 U7522 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U7523 ( .A1(n5989), .A2(n5988), .ZN(n5990) );
  NOR2_X1 U7524 ( .A1(n5991), .A2(n5990), .ZN(n5995) );
  OR2_X1 U7525 ( .A1(n5995), .A2(n5992), .ZN(n5993) );
  MUX2_X1 U7526 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5993), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5996) );
  INV_X1 U7527 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U7528 ( .A1(n5995), .A2(n5994), .ZN(n6090) );
  AND2_X1 U7529 ( .A1(n5996), .A2(n6090), .ZN(n6173) );
  AOI22_X1 U7530 ( .A1(n7703), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7714), .B2(
        n6173), .ZN(n5997) );
  XNOR2_X1 U7531 ( .A(n6955), .B(n8114), .ZN(n6861) );
  NAND2_X1 U7532 ( .A1(n4407), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6006) );
  INV_X1 U7533 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5999) );
  OR2_X1 U7534 ( .A1(n7783), .A2(n5999), .ZN(n6005) );
  INV_X1 U7535 ( .A(n6001), .ZN(n6000) );
  INV_X1 U7536 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7537 ( .A1(n6001), .A2(n6181), .ZN(n6002) );
  NAND2_X1 U7538 ( .A1(n6043), .A2(n6002), .ZN(n6733) );
  OR2_X1 U7539 ( .A1(n7768), .A2(n6733), .ZN(n6004) );
  INV_X1 U7540 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6174) );
  OR2_X1 U7541 ( .A1(n7771), .A2(n6174), .ZN(n6003) );
  NOR2_X1 U7542 ( .A1(n6983), .A2(n5905), .ZN(n6007) );
  NAND2_X1 U7543 ( .A1(n6861), .A2(n6007), .ZN(n6767) );
  INV_X1 U7544 ( .A(n6861), .ZN(n6009) );
  INV_X1 U7545 ( .A(n6007), .ZN(n6008) );
  NAND2_X1 U7546 ( .A1(n6009), .A2(n6008), .ZN(n6010) );
  NAND2_X1 U7547 ( .A1(n6767), .A2(n6010), .ZN(n6030) );
  NAND2_X1 U7548 ( .A1(n7230), .A2(n7387), .ZN(n9773) );
  XNOR2_X1 U7549 ( .A(n7230), .B(P2_B_REG_SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7550 ( .A1(n7342), .A2(n6011), .ZN(n6012) );
  INV_X1 U7551 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U7552 ( .A1(n9769), .A2(n6013), .ZN(n6014) );
  INV_X1 U7553 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9776) );
  NOR2_X1 U7554 ( .A1(n6016), .A2(n6015), .ZN(n9778) );
  AOI21_X1 U7555 ( .B1(n9769), .B2(n9776), .A(n9778), .ZN(n6549) );
  NOR4_X1 U7556 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6020) );
  NOR4_X1 U7557 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6019) );
  NOR4_X1 U7558 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6018) );
  NOR4_X1 U7559 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6017) );
  NAND4_X1 U7560 ( .A1(n6020), .A2(n6019), .A3(n6018), .A4(n6017), .ZN(n6026)
         );
  NOR2_X1 U7561 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .ZN(
        n6024) );
  NOR4_X1 U7562 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n6023) );
  NOR4_X1 U7563 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n6022) );
  NOR4_X1 U7564 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6021) );
  NAND4_X1 U7565 ( .A1(n6024), .A2(n6023), .A3(n6022), .A4(n6021), .ZN(n6025)
         );
  OAI21_X1 U7566 ( .B1(n6026), .B2(n6025), .A(n9769), .ZN(n6548) );
  NAND2_X1 U7567 ( .A1(n6549), .A2(n6548), .ZN(n6493) );
  INV_X1 U7568 ( .A(n8003), .ZN(n6051) );
  NAND2_X1 U7569 ( .A1(n8007), .A2(n7833), .ZN(n6140) );
  INV_X1 U7570 ( .A(n6140), .ZN(n6081) );
  NOR2_X1 U7571 ( .A1(n9815), .A2(n6081), .ZN(n6027) );
  INV_X1 U7572 ( .A(n6031), .ZN(n6029) );
  NAND2_X1 U7573 ( .A1(n6029), .A2(n6028), .ZN(n6768) );
  INV_X1 U7574 ( .A(n6768), .ZN(n6863) );
  AOI211_X1 U7575 ( .C1(n6031), .C2(n6030), .A(n8263), .B(n6863), .ZN(n6057)
         );
  INV_X1 U7576 ( .A(n7992), .ZN(n7964) );
  AND2_X1 U7577 ( .A1(n9780), .A2(n7964), .ZN(n6495) );
  NAND2_X1 U7578 ( .A1(n6050), .A2(n6495), .ZN(n6034) );
  AND2_X1 U7579 ( .A1(n7992), .A2(n8393), .ZN(n6032) );
  NAND2_X1 U7580 ( .A1(n9829), .A2(n7994), .ZN(n6547) );
  INV_X1 U7581 ( .A(n6547), .ZN(n6033) );
  NOR2_X1 U7582 ( .A1(n8248), .A2(n4536), .ZN(n6056) );
  INV_X1 U7583 ( .A(n6035), .ZN(n6036) );
  NAND2_X1 U7584 ( .A1(n6036), .A2(n6547), .ZN(n6040) );
  INV_X1 U7585 ( .A(n6083), .ZN(n6037) );
  AND3_X1 U7586 ( .A1(n6038), .A2(n6037), .A3(n6551), .ZN(n6039) );
  NAND2_X1 U7587 ( .A1(n6040), .A2(n6039), .ZN(n8011) );
  OAI22_X1 U7588 ( .A1(n8253), .A2(n6733), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6181), .ZN(n6055) );
  NAND2_X1 U7589 ( .A1(n4407), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6049) );
  INV_X1 U7590 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6041) );
  OR2_X1 U7591 ( .A1(n7783), .A2(n6041), .ZN(n6048) );
  NAND2_X1 U7592 ( .A1(n6043), .A2(n6042), .ZN(n6044) );
  NAND2_X1 U7593 ( .A1(n6787), .A2(n6044), .ZN(n6992) );
  OR2_X1 U7594 ( .A1(n7768), .A2(n6992), .ZN(n6047) );
  INV_X1 U7595 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6045) );
  OR2_X1 U7596 ( .A1(n7771), .A2(n6045), .ZN(n6046) );
  INV_X1 U7597 ( .A(n6050), .ZN(n6052) );
  NAND2_X1 U7598 ( .A1(n6081), .A2(n7402), .ZN(n8550) );
  NAND2_X1 U7599 ( .A1(n8245), .A2(n9752), .ZN(n8230) );
  INV_X1 U7600 ( .A(n7402), .ZN(n6053) );
  NAND2_X1 U7601 ( .A1(n8245), .A2(n9751), .ZN(n8231) );
  INV_X1 U7602 ( .A(n8281), .ZN(n6350) );
  OAI22_X1 U7603 ( .A1(n6963), .A2(n8230), .B1(n8231), .B2(n6350), .ZN(n6054)
         );
  OR4_X1 U7604 ( .A1(n6057), .A2(n6056), .A3(n6055), .A4(n6054), .ZN(P2_U3215)
         );
  NOR2_X1 U7605 ( .A1(n7428), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9367) );
  INV_X2 U7606 ( .A(n9367), .ZN(n9371) );
  INV_X2 U7607 ( .A(n7176), .ZN(n9369) );
  INV_X1 U7608 ( .A(n6462), .ZN(n6058) );
  OAI222_X1 U7609 ( .A1(n9371), .A2(n6059), .B1(n9369), .B2(n6066), .C1(n6058), 
        .C2(P1_U3084), .ZN(P1_U3351) );
  INV_X1 U7610 ( .A(n8855), .ZN(n6060) );
  OAI222_X1 U7611 ( .A1(n9371), .A2(n9971), .B1(n9369), .B2(n6076), .C1(n6060), 
        .C2(P1_U3084), .ZN(P1_U3352) );
  OAI222_X1 U7612 ( .A1(n9371), .A2(n6061), .B1(n9369), .B2(n6072), .C1(n6284), 
        .C2(P1_U3084), .ZN(P1_U3350) );
  OAI222_X1 U7613 ( .A1(n9371), .A2(n6062), .B1(n9369), .B2(n6068), .C1(n9547), 
        .C2(P1_U3084), .ZN(P1_U3349) );
  OAI222_X1 U7614 ( .A1(n6063), .A2(P1_U3084), .B1(n9369), .B2(n6071), .C1(
        n9979), .C2(n9371), .ZN(P1_U3348) );
  OAI222_X1 U7615 ( .A1(n9371), .A2(n6064), .B1(n9369), .B2(n6070), .C1(n9580), 
        .C2(P1_U3084), .ZN(P1_U3347) );
  INV_X1 U7616 ( .A(n7404), .ZN(n7173) );
  NOR2_X1 U7617 ( .A1(n7428), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8679) );
  INV_X1 U7618 ( .A(n9394), .ZN(n6065) );
  OAI222_X1 U7619 ( .A1(n7404), .A2(n6067), .B1(n8131), .B2(n6066), .C1(
        P2_U3152), .C2(n6065), .ZN(P2_U3356) );
  INV_X1 U7620 ( .A(n6239), .ZN(n6170) );
  OAI222_X1 U7621 ( .A1(n7404), .A2(n6069), .B1(n8131), .B2(n6068), .C1(
        P2_U3152), .C2(n6170), .ZN(P2_U3354) );
  INV_X1 U7622 ( .A(n6207), .ZN(n6221) );
  OAI222_X1 U7623 ( .A1(n7404), .A2(n9981), .B1(n8131), .B2(n6070), .C1(
        P2_U3152), .C2(n6221), .ZN(P2_U3352) );
  OAI222_X1 U7624 ( .A1(n7404), .A2(n10104), .B1(n8131), .B2(n6071), .C1(
        P2_U3152), .C2(n6205), .ZN(P2_U3353) );
  INV_X1 U7625 ( .A(n6168), .ZN(n6311) );
  OAI222_X1 U7626 ( .A1(n7404), .A2(n6073), .B1(n8131), .B2(n6072), .C1(
        P2_U3152), .C2(n6311), .ZN(P2_U3355) );
  OAI222_X1 U7627 ( .A1(n6279), .A2(P1_U3084), .B1(n9369), .B2(n6075), .C1(
        n6074), .C2(n9371), .ZN(P1_U3346) );
  INV_X1 U7628 ( .A(n6173), .ZN(n6194) );
  OAI222_X1 U7629 ( .A1(n7404), .A2(n10158), .B1(n8131), .B2(n6075), .C1(
        P2_U3152), .C2(n6194), .ZN(P2_U3351) );
  OAI222_X1 U7630 ( .A1(n7404), .A2(n10182), .B1(n8131), .B2(n6076), .C1(
        P2_U3152), .C2(n6164), .ZN(P2_U3357) );
  INV_X1 U7631 ( .A(n6770), .ZN(n6079) );
  NAND2_X1 U7632 ( .A1(n6090), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6077) );
  XNOR2_X1 U7633 ( .A(n6077), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6771) );
  INV_X1 U7634 ( .A(n6771), .ZN(n6365) );
  OAI222_X1 U7635 ( .A1(n7404), .A2(n6078), .B1(n8131), .B2(n6079), .C1(
        P2_U3152), .C2(n6365), .ZN(P2_U3350) );
  OAI222_X1 U7636 ( .A1(n9371), .A2(n6080), .B1(n9369), .B2(n6079), .C1(n9587), 
        .C2(P1_U3084), .ZN(P1_U3345) );
  NAND2_X1 U7637 ( .A1(n9771), .A2(n6081), .ZN(n6082) );
  NAND2_X1 U7638 ( .A1(n6082), .A2(n4492), .ZN(n6085) );
  AND2_X1 U7639 ( .A1(n6083), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8002) );
  OR2_X1 U7640 ( .A1(n9771), .A2(n8002), .ZN(n6084) );
  NAND2_X1 U7641 ( .A1(n6085), .A2(n6084), .ZN(n9888) );
  NOR2_X1 U7642 ( .A1(n9739), .A2(n8264), .ZN(P2_U3151) );
  INV_X1 U7643 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10000) );
  INV_X1 U7644 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8333) );
  NAND2_X1 U7645 ( .A1(n4401), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6088) );
  INV_X1 U7646 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6086) );
  OR2_X1 U7647 ( .A1(n7802), .A2(n6086), .ZN(n6087) );
  OAI211_X1 U7648 ( .C1(n7771), .C2(n8333), .A(n6088), .B(n6087), .ZN(n8335)
         );
  NAND2_X1 U7649 ( .A1(n8264), .A2(n8335), .ZN(n6089) );
  OAI21_X1 U7650 ( .B1(n8264), .B2(n10000), .A(n6089), .ZN(P2_U3583) );
  INV_X1 U7651 ( .A(n6781), .ZN(n6092) );
  NAND2_X1 U7652 ( .A1(n6137), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6093) );
  XNOR2_X1 U7653 ( .A(n6093), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6782) );
  AOI22_X1 U7654 ( .A1(n6782), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n7173), .ZN(n6091) );
  OAI21_X1 U7655 ( .B1(n6092), .B2(n8131), .A(n6091), .ZN(P2_U3349) );
  INV_X1 U7656 ( .A(n6295), .ZN(n9611) );
  OAI222_X1 U7657 ( .A1(P1_U3084), .A2(n9611), .B1(n9369), .B2(n6092), .C1(
        n10161), .C2(n9371), .ZN(P1_U3344) );
  INV_X1 U7658 ( .A(n6910), .ZN(n6113) );
  NAND2_X1 U7659 ( .A1(n6093), .A2(n6134), .ZN(n6094) );
  NAND2_X1 U7660 ( .A1(n6094), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6098) );
  INV_X1 U7661 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7662 ( .A1(n6098), .A2(n6135), .ZN(n6095) );
  NAND2_X1 U7663 ( .A1(n6095), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6096) );
  XNOR2_X1 U7664 ( .A(n6096), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6911) );
  AOI22_X1 U7665 ( .A1(n6911), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n7173), .ZN(n6097) );
  OAI21_X1 U7666 ( .B1(n6113), .B2(n8131), .A(n6097), .ZN(P2_U3347) );
  INV_X1 U7667 ( .A(n6881), .ZN(n6100) );
  XNOR2_X1 U7668 ( .A(n6098), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6882) );
  INV_X1 U7669 ( .A(n6882), .ZN(n9899) );
  OAI222_X1 U7670 ( .A1(n7404), .A2(n10117), .B1(n8131), .B2(n6100), .C1(n9899), .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7671 ( .A(n6323), .ZN(n6269) );
  OAI222_X1 U7672 ( .A1(P1_U3084), .A2(n6269), .B1(n9369), .B2(n6100), .C1(
        n6099), .C2(n9371), .ZN(P1_U3343) );
  NAND2_X1 U7673 ( .A1(n4401), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6111) );
  INV_X1 U7674 ( .A(n6898), .ZN(n6102) );
  INV_X1 U7675 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7676 ( .A1(n7102), .A2(n6105), .ZN(n6106) );
  NAND2_X1 U7677 ( .A1(n7695), .A2(n6106), .ZN(n8254) );
  OR2_X1 U7678 ( .A1(n7768), .A2(n8254), .ZN(n6110) );
  INV_X1 U7679 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7381) );
  OR2_X1 U7680 ( .A1(n7771), .A2(n7381), .ZN(n6109) );
  INV_X1 U7681 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6107) );
  OR2_X1 U7682 ( .A1(n7802), .A2(n6107), .ZN(n6108) );
  NAND2_X1 U7683 ( .A1(n8271), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n6112) );
  OAI21_X1 U7684 ( .B1(n8271), .B2(n8549), .A(n6112), .ZN(P2_U3567) );
  INV_X1 U7685 ( .A(n6394), .ZN(n6388) );
  OAI222_X1 U7686 ( .A1(n9371), .A2(n6114), .B1(n9369), .B2(n6113), .C1(
        P1_U3084), .C2(n6388), .ZN(P1_U3342) );
  INV_X1 U7687 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6119) );
  INV_X1 U7688 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U7689 ( .A1(n7418), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U7690 ( .A1(n4409), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6115) );
  OAI211_X1 U7691 ( .C1(n7421), .C2(n6117), .A(n6116), .B(n6115), .ZN(n8938)
         );
  NAND2_X1 U7692 ( .A1(n8938), .A2(P1_U4006), .ZN(n6118) );
  OAI21_X1 U7693 ( .B1(P1_U4006), .B2(n6119), .A(n6118), .ZN(P1_U3586) );
  NAND2_X1 U7694 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_17__SCAN_IN), 
        .ZN(n6120) );
  INV_X1 U7695 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8159) );
  NAND2_X1 U7696 ( .A1(n7726), .A2(n8159), .ZN(n6123) );
  AND2_X1 U7697 ( .A1(n7744), .A2(n6123), .ZN(n8463) );
  NAND2_X1 U7698 ( .A1(n8463), .A2(n7780), .ZN(n6129) );
  INV_X1 U7699 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n6126) );
  NAND2_X1 U7700 ( .A1(n4407), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6125) );
  NAND2_X1 U7701 ( .A1(n4401), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6124) );
  OAI211_X1 U7702 ( .C1(n6126), .C2(n7771), .A(n6125), .B(n6124), .ZN(n6127)
         );
  INV_X1 U7703 ( .A(n6127), .ZN(n6128) );
  NAND2_X1 U7704 ( .A1(n6129), .A2(n6128), .ZN(n8449) );
  NAND2_X1 U7705 ( .A1(n8449), .A2(n8264), .ZN(n6130) );
  OAI21_X1 U7706 ( .B1(n8264), .B2(n5611), .A(n6130), .ZN(P2_U3573) );
  NAND2_X1 U7707 ( .A1(n6634), .A2(P1_U4006), .ZN(n6131) );
  OAI21_X1 U7708 ( .B1(P1_U4006), .B2(n5903), .A(n6131), .ZN(P1_U3555) );
  INV_X1 U7709 ( .A(n9624), .ZN(n6390) );
  INV_X1 U7710 ( .A(n7015), .ZN(n6139) );
  OAI222_X1 U7711 ( .A1(n6390), .A2(P1_U3084), .B1(n9369), .B2(n6139), .C1(
        n6132), .C2(n9371), .ZN(P1_U3341) );
  INV_X1 U7712 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6133) );
  NAND3_X1 U7713 ( .A1(n6135), .A2(n6134), .A3(n6133), .ZN(n6136) );
  NAND2_X1 U7714 ( .A1(n6222), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6138) );
  XNOR2_X1 U7715 ( .A(n6138), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7016) );
  INV_X1 U7716 ( .A(n7016), .ZN(n6838) );
  OAI222_X1 U7717 ( .A1(n7404), .A2(n9970), .B1(n8131), .B2(n6139), .C1(
        P2_U3152), .C2(n6838), .ZN(P2_U3346) );
  NAND2_X1 U7718 ( .A1(n9771), .A2(n6140), .ZN(n6142) );
  INV_X1 U7719 ( .A(n8002), .ZN(n8006) );
  NAND3_X1 U7720 ( .A1(n6142), .A2(n8006), .A3(n6141), .ZN(n6144) );
  NAND2_X1 U7721 ( .A1(n6144), .A2(n4492), .ZN(n6159) );
  NAND2_X1 U7722 ( .A1(n6159), .A2(n8271), .ZN(n6176) );
  NAND2_X1 U7723 ( .A1(n6176), .A2(n7402), .ZN(n9900) );
  NAND2_X1 U7724 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n6859) );
  INV_X1 U7725 ( .A(n6859), .ZN(n6163) );
  NAND2_X1 U7726 ( .A1(n6168), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6149) );
  MUX2_X1 U7727 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6145), .S(n6168), .Z(n6306)
         );
  NAND2_X1 U7728 ( .A1(n9394), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6148) );
  MUX2_X1 U7729 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6146), .S(n9394), .Z(n9397)
         );
  MUX2_X1 U7730 ( .A(n6147), .B(P2_REG1_REG_1__SCAN_IN), .S(n6164), .Z(n9384)
         );
  NAND3_X1 U7731 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n9384), .ZN(n9383) );
  OAI21_X1 U7732 ( .B1(n6164), .B2(n6147), .A(n9383), .ZN(n9398) );
  NAND2_X1 U7733 ( .A1(n9397), .A2(n9398), .ZN(n9396) );
  NAND2_X1 U7734 ( .A1(n6148), .A2(n9396), .ZN(n6307) );
  NAND2_X1 U7735 ( .A1(n6306), .A2(n6307), .ZN(n6305) );
  NAND2_X1 U7736 ( .A1(n6149), .A2(n6305), .ZN(n6234) );
  INV_X1 U7737 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6150) );
  MUX2_X1 U7738 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6150), .S(n6239), .Z(n6233)
         );
  NAND2_X1 U7739 ( .A1(n6234), .A2(n6233), .ZN(n6232) );
  NAND2_X1 U7740 ( .A1(n6239), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6196) );
  MUX2_X1 U7741 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n5956), .S(n6205), .Z(n6195)
         );
  AOI21_X1 U7742 ( .B1(n6232), .B2(n6196), .A(n6195), .ZN(n6211) );
  INV_X1 U7743 ( .A(n6211), .ZN(n6153) );
  INV_X1 U7744 ( .A(n6205), .ZN(n6151) );
  NAND2_X1 U7745 ( .A1(n6151), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6206) );
  MUX2_X1 U7746 ( .A(n6208), .B(P2_REG1_REG_6__SCAN_IN), .S(n6207), .Z(n6152)
         );
  AOI21_X1 U7747 ( .B1(n6153), .B2(n6206), .A(n6152), .ZN(n6213) );
  INV_X1 U7748 ( .A(n6213), .ZN(n6184) );
  NAND2_X1 U7749 ( .A1(n6207), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6183) );
  INV_X1 U7750 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6872) );
  MUX2_X1 U7751 ( .A(n6872), .B(P2_REG1_REG_7__SCAN_IN), .S(n6173), .Z(n6182)
         );
  AOI21_X1 U7752 ( .B1(n6184), .B2(n6183), .A(n6182), .ZN(n6186) );
  INV_X1 U7753 ( .A(n6186), .ZN(n6155) );
  NAND2_X1 U7754 ( .A1(n6173), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6156) );
  INV_X1 U7755 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9847) );
  MUX2_X1 U7756 ( .A(n9847), .B(P2_REG1_REG_8__SCAN_IN), .S(n6771), .Z(n6154)
         );
  AOI21_X1 U7757 ( .B1(n6155), .B2(n6156), .A(n6154), .ZN(n6363) );
  INV_X1 U7758 ( .A(n6156), .ZN(n6158) );
  MUX2_X1 U7759 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9847), .S(n6771), .Z(n6157)
         );
  NOR3_X1 U7760 ( .A1(n6186), .A2(n6158), .A3(n6157), .ZN(n6161) );
  INV_X1 U7761 ( .A(n6159), .ZN(n6160) );
  NAND2_X1 U7762 ( .A1(n6160), .A2(n8037), .ZN(n9741) );
  NOR3_X1 U7763 ( .A1(n6363), .A2(n6161), .A3(n9741), .ZN(n6162) );
  AOI211_X1 U7764 ( .C1(n9739), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n6163), .B(
        n6162), .ZN(n6180) );
  MUX2_X1 U7765 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6045), .S(n6771), .Z(n6178)
         );
  MUX2_X1 U7766 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6171), .S(n6239), .Z(n6242)
         );
  MUX2_X1 U7767 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6165), .S(n6164), .Z(n9378)
         );
  NAND2_X1 U7768 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9379) );
  NOR2_X1 U7769 ( .A1(n9378), .A2(n9379), .ZN(n9377) );
  AOI21_X1 U7770 ( .B1(n9381), .B2(P2_REG2_REG_1__SCAN_IN), .A(n9377), .ZN(
        n9392) );
  NAND2_X1 U7771 ( .A1(n9394), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6166) );
  OAI21_X1 U7772 ( .B1(n9394), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6166), .ZN(
        n9391) );
  NOR2_X1 U7773 ( .A1(n9392), .A2(n9391), .ZN(n9390) );
  AOI21_X1 U7774 ( .B1(n9394), .B2(P2_REG2_REG_2__SCAN_IN), .A(n9390), .ZN(
        n6304) );
  NAND2_X1 U7775 ( .A1(n6168), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6167) );
  OAI21_X1 U7776 ( .B1(n6168), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6167), .ZN(
        n6303) );
  NOR2_X1 U7777 ( .A1(n6304), .A2(n6303), .ZN(n6302) );
  XNOR2_X1 U7778 ( .A(n6205), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n6202) );
  NAND2_X1 U7779 ( .A1(n6201), .A2(n6202), .ZN(n6200) );
  XOR2_X1 U7780 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6207), .Z(n6218) );
  MUX2_X1 U7781 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6174), .S(n6173), .Z(n6191)
         );
  OAI21_X1 U7782 ( .B1(n6174), .B2(n6194), .A(n6189), .ZN(n6177) );
  NOR2_X1 U7783 ( .A1(n7402), .A2(n8037), .ZN(n6175) );
  OAI211_X1 U7784 ( .C1(n6178), .C2(n6177), .A(n9896), .B(n6357), .ZN(n6179)
         );
  OAI211_X1 U7785 ( .C1(n9900), .C2(n6365), .A(n6180), .B(n6179), .ZN(P2_U3253) );
  NOR2_X1 U7786 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6181), .ZN(n6188) );
  AND3_X1 U7787 ( .A1(n6184), .A2(n6183), .A3(n6182), .ZN(n6185) );
  NOR3_X1 U7788 ( .A1(n6186), .A2(n6185), .A3(n9741), .ZN(n6187) );
  AOI211_X1 U7789 ( .C1(n9739), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n6188), .B(
        n6187), .ZN(n6193) );
  OAI211_X1 U7790 ( .C1(n6191), .C2(n6190), .A(n9896), .B(n6189), .ZN(n6192)
         );
  OAI211_X1 U7791 ( .C1(n9900), .C2(n6194), .A(n6193), .B(n6192), .ZN(P2_U3252) );
  NOR2_X1 U7792 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10132), .ZN(n6199) );
  AND3_X1 U7793 ( .A1(n6232), .A2(n6196), .A3(n6195), .ZN(n6197) );
  NOR3_X1 U7794 ( .A1(n9741), .A2(n6211), .A3(n6197), .ZN(n6198) );
  AOI211_X1 U7795 ( .C1(n9739), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n6199), .B(
        n6198), .ZN(n6204) );
  OAI211_X1 U7796 ( .C1(n6202), .C2(n6201), .A(n9896), .B(n6200), .ZN(n6203)
         );
  OAI211_X1 U7797 ( .C1(n9900), .C2(n6205), .A(n6204), .B(n6203), .ZN(P2_U3250) );
  NAND2_X1 U7798 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n6429) );
  INV_X1 U7799 ( .A(n6429), .ZN(n6215) );
  INV_X1 U7800 ( .A(n6206), .ZN(n6210) );
  MUX2_X1 U7801 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6208), .S(n6207), .Z(n6209)
         );
  NOR3_X1 U7802 ( .A1(n6211), .A2(n6210), .A3(n6209), .ZN(n6212) );
  NOR3_X1 U7803 ( .A1(n9741), .A2(n6213), .A3(n6212), .ZN(n6214) );
  AOI211_X1 U7804 ( .C1(n9739), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n6215), .B(
        n6214), .ZN(n6220) );
  OAI211_X1 U7805 ( .C1(n6218), .C2(n6217), .A(n9896), .B(n6216), .ZN(n6219)
         );
  OAI211_X1 U7806 ( .C1(n9900), .C2(n6221), .A(n6220), .B(n6219), .ZN(P2_U3251) );
  INV_X1 U7807 ( .A(n7095), .ZN(n6225) );
  NAND2_X1 U7808 ( .A1(n6223), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6227) );
  XNOR2_X1 U7809 ( .A(n6227), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7096) );
  INV_X1 U7810 ( .A(n7096), .ZN(n6999) );
  OAI222_X1 U7811 ( .A1(n7404), .A2(n6224), .B1(n8131), .B2(n6225), .C1(n6999), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U7812 ( .A(n6539), .ZN(n6535) );
  OAI222_X1 U7813 ( .A1(P1_U3084), .A2(n6535), .B1(n9369), .B2(n6225), .C1(
        n10026), .C2(n9371), .ZN(P1_U3340) );
  INV_X1 U7814 ( .A(n7208), .ZN(n6231) );
  NAND2_X1 U7815 ( .A1(n6227), .A2(n6226), .ZN(n6228) );
  NAND2_X1 U7816 ( .A1(n6228), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6437) );
  XNOR2_X1 U7817 ( .A(n6437), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7209) );
  INV_X1 U7818 ( .A(n7209), .ZN(n7135) );
  OAI222_X1 U7819 ( .A1(n7404), .A2(n6229), .B1(n8131), .B2(n6231), .C1(n7135), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U7820 ( .A(n6541), .ZN(n8900) );
  OAI222_X1 U7821 ( .A1(P1_U3084), .A2(n8900), .B1(n9369), .B2(n6231), .C1(
        n6230), .C2(n9371), .ZN(P1_U3339) );
  INV_X1 U7822 ( .A(n9900), .ZN(n9395) );
  OAI21_X1 U7823 ( .B1(n6234), .B2(n6233), .A(n6232), .ZN(n6237) );
  AND2_X1 U7824 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6235) );
  AOI21_X1 U7825 ( .B1(n9739), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6235), .ZN(
        n6236) );
  OAI21_X1 U7826 ( .B1(n9741), .B2(n6237), .A(n6236), .ZN(n6238) );
  AOI21_X1 U7827 ( .B1(n6239), .B2(n9395), .A(n6238), .ZN(n6244) );
  OAI211_X1 U7828 ( .C1(n6242), .C2(n6241), .A(n9896), .B(n6240), .ZN(n6243)
         );
  NAND2_X1 U7829 ( .A1(n6244), .A2(n6243), .ZN(P2_U3249) );
  INV_X1 U7830 ( .A(n6505), .ZN(n6252) );
  NOR2_X1 U7831 ( .A1(n6245), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9738) );
  NOR2_X1 U7832 ( .A1(n8248), .A2(n9759), .ZN(n6246) );
  AOI211_X1 U7833 ( .C1(P2_REG3_REG_0__SCAN_IN), .C2(n8011), .A(n9738), .B(
        n6246), .ZN(n6251) );
  INV_X1 U7834 ( .A(n6484), .ZN(n6247) );
  OAI22_X1 U7835 ( .A1(n8255), .A2(n6247), .B1(n9759), .B2(n8263), .ZN(n6249)
         );
  NAND2_X1 U7836 ( .A1(n6249), .A2(n6248), .ZN(n6250) );
  OAI211_X1 U7837 ( .C1(n6252), .C2(n8230), .A(n6251), .B(n6250), .ZN(P2_U3234) );
  NOR2_X1 U7838 ( .A1(n6295), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6268) );
  MUX2_X1 U7839 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n5373), .S(n6295), .Z(n9614)
         );
  OR2_X1 U7840 ( .A1(n8878), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6265) );
  AOI22_X1 U7841 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n8878), .B1(n6279), .B2(
        n5333), .ZN(n8876) );
  XNOR2_X1 U7842 ( .A(n9580), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9575) );
  XNOR2_X1 U7843 ( .A(n6462), .B(n6253), .ZN(n6458) );
  MUX2_X1 U7844 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n5186), .S(n8855), .Z(n8849)
         );
  AND2_X1 U7845 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6254) );
  NAND2_X1 U7846 ( .A1(n8849), .A2(n6254), .ZN(n8850) );
  NAND2_X1 U7847 ( .A1(n8855), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7848 ( .A1(n8850), .A2(n6255), .ZN(n6457) );
  NAND2_X1 U7849 ( .A1(n6458), .A2(n6457), .ZN(n6456) );
  NAND2_X1 U7850 ( .A1(n6462), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U7851 ( .A1(n6456), .A2(n6256), .ZN(n8863) );
  XNOR2_X1 U7852 ( .A(n6284), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n8864) );
  NAND2_X1 U7853 ( .A1(n8863), .A2(n8864), .ZN(n8862) );
  OR2_X1 U7854 ( .A1(n6284), .A2(n6257), .ZN(n6258) );
  NAND2_X1 U7855 ( .A1(n8862), .A2(n6258), .ZN(n9540) );
  MUX2_X1 U7856 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6259), .S(n9547), .Z(n9541)
         );
  NOR2_X1 U7857 ( .A1(n9540), .A2(n9541), .ZN(n9539) );
  AND2_X1 U7858 ( .A1(n9547), .A2(n6259), .ZN(n6260) );
  OR2_X1 U7859 ( .A1(n9539), .A2(n6260), .ZN(n9555) );
  NAND2_X1 U7860 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9566), .ZN(n6261) );
  OAI21_X1 U7861 ( .B1(n9566), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6261), .ZN(
        n9554) );
  NOR2_X1 U7862 ( .A1(n9555), .A2(n9554), .ZN(n9557) );
  AOI21_X1 U7863 ( .B1(n9566), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9557), .ZN(
        n9574) );
  NAND2_X1 U7864 ( .A1(n9575), .A2(n9574), .ZN(n6264) );
  NAND2_X1 U7865 ( .A1(n9580), .A2(n6262), .ZN(n6263) );
  NAND2_X1 U7866 ( .A1(n6264), .A2(n6263), .ZN(n8875) );
  NAND2_X1 U7867 ( .A1(n8876), .A2(n8875), .ZN(n8874) );
  NAND2_X1 U7868 ( .A1(n6265), .A2(n8874), .ZN(n9599) );
  OAI21_X1 U7869 ( .B1(n9587), .B2(n6266), .A(n9599), .ZN(n6267) );
  NAND2_X1 U7870 ( .A1(n9587), .A2(n6266), .ZN(n9585) );
  NAND2_X1 U7871 ( .A1(n6267), .A2(n9585), .ZN(n9613) );
  NOR2_X1 U7872 ( .A1(n6268), .A2(n9616), .ZN(n6316) );
  AOI22_X1 U7873 ( .A1(n6323), .A2(n5400), .B1(P1_REG1_REG_10__SCAN_IN), .B2(
        n6269), .ZN(n6315) );
  NOR2_X1 U7874 ( .A1(n6316), .A2(n6315), .ZN(n6314) );
  AOI21_X1 U7875 ( .B1(n6269), .B2(n5400), .A(n6314), .ZN(n6272) );
  INV_X1 U7876 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6270) );
  MUX2_X1 U7877 ( .A(n6270), .B(P1_REG1_REG_11__SCAN_IN), .S(n6394), .Z(n6271)
         );
  NOR2_X1 U7878 ( .A1(n6272), .A2(n6271), .ZN(n6387) );
  AOI21_X1 U7879 ( .B1(n6272), .B2(n6271), .A(n6387), .ZN(n6301) );
  NOR2_X1 U7880 ( .A1(n6273), .A2(P1_U3084), .ZN(n6278) );
  NAND2_X1 U7881 ( .A1(n6278), .A2(n6628), .ZN(n9528) );
  INV_X1 U7882 ( .A(n6274), .ZN(n8936) );
  INV_X1 U7883 ( .A(n6275), .ZN(n6276) );
  OR2_X1 U7884 ( .A1(P1_U3083), .A2(n6276), .ZN(n9675) );
  INV_X1 U7885 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6277) );
  NOR2_X1 U7886 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6277), .ZN(n8781) );
  NAND2_X1 U7887 ( .A1(n6278), .A2(n8936), .ZN(n6297) );
  INV_X1 U7888 ( .A(n6297), .ZN(n9529) );
  INV_X1 U7889 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6291) );
  MUX2_X1 U7890 ( .A(n6291), .B(P1_REG2_REG_8__SCAN_IN), .S(n9587), .Z(n6290)
         );
  AOI22_X1 U7891 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n8878), .B1(n6279), .B2(
        n6947), .ZN(n8883) );
  INV_X1 U7892 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6288) );
  XNOR2_X1 U7893 ( .A(n9580), .B(n6288), .ZN(n9569) );
  NOR2_X1 U7894 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9566), .ZN(n6280) );
  AOI21_X1 U7895 ( .B1(n9566), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6280), .ZN(
        n9561) );
  INV_X1 U7896 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6692) );
  XNOR2_X1 U7897 ( .A(n6462), .B(n6692), .ZN(n6461) );
  INV_X1 U7898 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6281) );
  MUX2_X1 U7899 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6281), .S(n8855), .Z(n8858)
         );
  AND2_X1 U7900 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n8857) );
  NAND2_X1 U7901 ( .A1(n8858), .A2(n8857), .ZN(n8856) );
  NAND2_X1 U7902 ( .A1(n8855), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6282) );
  NAND2_X1 U7903 ( .A1(n6462), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U7904 ( .A1(n6459), .A2(n6283), .ZN(n8868) );
  XNOR2_X1 U7905 ( .A(n6284), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n8869) );
  NAND2_X1 U7906 ( .A1(n8868), .A2(n8869), .ZN(n8867) );
  INV_X1 U7907 ( .A(n6284), .ZN(n8866) );
  NAND2_X1 U7908 ( .A1(n8866), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7909 ( .A1(n8867), .A2(n6285), .ZN(n9546) );
  INV_X1 U7910 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6286) );
  MUX2_X1 U7911 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6286), .S(n9547), .Z(n9545)
         );
  AND2_X1 U7912 ( .A1(n9547), .A2(n6286), .ZN(n6287) );
  NAND2_X1 U7913 ( .A1(n9561), .A2(n9562), .ZN(n9560) );
  OAI21_X1 U7914 ( .B1(n9566), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9560), .ZN(
        n9570) );
  OR2_X1 U7915 ( .A1(n9569), .A2(n9570), .ZN(n9571) );
  OR2_X1 U7916 ( .A1(n9580), .A2(n6288), .ZN(n6289) );
  NAND2_X1 U7917 ( .A1(n8883), .A2(n8882), .ZN(n8881) );
  OAI21_X1 U7918 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n8878), .A(n8881), .ZN(
        n9588) );
  NAND2_X1 U7919 ( .A1(n6290), .A2(n9588), .ZN(n9592) );
  NAND2_X1 U7920 ( .A1(n9587), .A2(n6291), .ZN(n6292) );
  NAND2_X1 U7921 ( .A1(n9592), .A2(n6292), .ZN(n9606) );
  OR2_X1 U7922 ( .A1(n6295), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6294) );
  NAND2_X1 U7923 ( .A1(n6295), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U7924 ( .A1(n6294), .A2(n6293), .ZN(n9605) );
  NOR2_X1 U7925 ( .A1(n9606), .A2(n9605), .ZN(n9604) );
  AOI21_X1 U7926 ( .B1(n6295), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9604), .ZN(
        n6320) );
  NAND2_X1 U7927 ( .A1(n6323), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6296) );
  OAI21_X1 U7928 ( .B1(n6323), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6296), .ZN(
        n6319) );
  NOR2_X1 U7929 ( .A1(n6320), .A2(n6319), .ZN(n6318) );
  XNOR2_X1 U7930 ( .A(n6394), .B(n9478), .ZN(n6397) );
  XOR2_X1 U7931 ( .A(n6396), .B(n6397), .Z(n6298) );
  OR2_X1 U7932 ( .A1(n6297), .A2(n6628), .ZN(n9666) );
  OAI22_X1 U7933 ( .A1(n9645), .A2(n6298), .B1(n6388), .B2(n9666), .ZN(n6299)
         );
  AOI211_X1 U7934 ( .C1(n9581), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n8781), .B(
        n6299), .ZN(n6300) );
  OAI21_X1 U7935 ( .B1(n6301), .B2(n9630), .A(n6300), .ZN(P1_U3252) );
  AOI211_X1 U7936 ( .C1(n6304), .C2(n6303), .A(n6302), .B(n9740), .ZN(n6313)
         );
  OAI211_X1 U7937 ( .C1(n6307), .C2(n6306), .A(n9891), .B(n6305), .ZN(n6310)
         );
  INV_X1 U7938 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6574) );
  NOR2_X1 U7939 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6574), .ZN(n6308) );
  AOI21_X1 U7940 ( .B1(n9739), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6308), .ZN(
        n6309) );
  OAI211_X1 U7941 ( .C1(n9900), .C2(n6311), .A(n6310), .B(n6309), .ZN(n6312)
         );
  OR2_X1 U7942 ( .A1(n6313), .A2(n6312), .ZN(P2_U3248) );
  AOI21_X1 U7943 ( .B1(n6316), .B2(n6315), .A(n6314), .ZN(n6325) );
  INV_X1 U7944 ( .A(n9666), .ZN(n9651) );
  INV_X1 U7945 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6317) );
  NAND2_X1 U7946 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8696) );
  OAI21_X1 U7947 ( .B1(n9675), .B2(n6317), .A(n8696), .ZN(n6322) );
  AOI211_X1 U7948 ( .C1(n6320), .C2(n6319), .A(n6318), .B(n9645), .ZN(n6321)
         );
  AOI211_X1 U7949 ( .C1(n9651), .C2(n6323), .A(n6322), .B(n6321), .ZN(n6324)
         );
  OAI21_X1 U7950 ( .B1(n6325), .B2(n9630), .A(n6324), .ZN(P1_U3251) );
  INV_X1 U7951 ( .A(n6635), .ZN(n6329) );
  INV_X1 U7952 ( .A(n6626), .ZN(n6762) );
  NOR2_X1 U7953 ( .A1(n6634), .A2(n6762), .ZN(n6681) );
  AND2_X1 U7954 ( .A1(n6634), .A2(n6762), .ZN(n7620) );
  NOR2_X1 U7955 ( .A1(n6681), .A2(n7620), .ZN(n7492) );
  NAND2_X1 U7956 ( .A1(n6721), .A2(n6635), .ZN(n6326) );
  OR2_X1 U7957 ( .A1(n7492), .A2(n6326), .ZN(n6328) );
  NAND2_X1 U7958 ( .A1(n6625), .A2(n9254), .ZN(n6327) );
  NAND2_X1 U7959 ( .A1(n6328), .A2(n6327), .ZN(n6765) );
  AOI21_X1 U7960 ( .B1(n6626), .B2(n6329), .A(n6765), .ZN(n6338) );
  INV_X1 U7961 ( .A(n6948), .ZN(n9362) );
  NAND2_X1 U7962 ( .A1(n6331), .A2(n6330), .ZN(n6334) );
  NOR2_X1 U7963 ( .A1(n9362), .A2(n6334), .ZN(n6332) );
  INV_X1 U7964 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10052) );
  NAND2_X1 U7965 ( .A1(n9727), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6333) );
  OAI21_X1 U7966 ( .B1(n6338), .B2(n9727), .A(n6333), .ZN(P1_U3454) );
  NOR2_X1 U7967 ( .A1(n6334), .A2(n6948), .ZN(n6335) );
  NAND2_X1 U7968 ( .A1(n9735), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6337) );
  OAI21_X1 U7969 ( .B1(n6338), .B2(n9735), .A(n6337), .ZN(P1_U3523) );
  INV_X1 U7970 ( .A(n8253), .ZN(n8211) );
  NAND2_X1 U7971 ( .A1(n6506), .A2(n9751), .ZN(n6340) );
  NAND2_X1 U7972 ( .A1(n8283), .A2(n9752), .ZN(n6339) );
  NAND2_X1 U7973 ( .A1(n6340), .A2(n6339), .ZN(n6577) );
  AOI22_X1 U7974 ( .A1(n8245), .A2(n6577), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3152), .ZN(n6341) );
  OAI21_X1 U7975 ( .B1(n8248), .B2(n9796), .A(n6341), .ZN(n6346) );
  INV_X1 U7976 ( .A(n8206), .ZN(n6342) );
  AOI211_X1 U7977 ( .C1(n6344), .C2(n6343), .A(n8263), .B(n6342), .ZN(n6345)
         );
  AOI211_X1 U7978 ( .C1(n8211), .C2(n6574), .A(n6346), .B(n6345), .ZN(n6347)
         );
  INV_X1 U7979 ( .A(n6347), .ZN(P2_U3220) );
  INV_X1 U7980 ( .A(n8263), .ZN(n8207) );
  OAI211_X1 U7981 ( .C1(n4491), .C2(n6349), .A(n6425), .B(n8207), .ZN(n6354)
         );
  INV_X1 U7982 ( .A(n8231), .ZN(n8249) );
  OAI22_X1 U7983 ( .A1(n8253), .A2(n6585), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10132), .ZN(n6352) );
  OAI22_X1 U7984 ( .A1(n6587), .A2(n8248), .B1(n8230), .B2(n6350), .ZN(n6351)
         );
  AOI211_X1 U7985 ( .C1(n8249), .C2(n8283), .A(n6352), .B(n6351), .ZN(n6353)
         );
  NAND2_X1 U7986 ( .A1(n6354), .A2(n6353), .ZN(P2_U3229) );
  NAND2_X1 U7987 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n6796) );
  INV_X1 U7988 ( .A(n6796), .ZN(n6355) );
  AOI21_X1 U7989 ( .B1(n9739), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n6355), .ZN(
        n6356) );
  INV_X1 U7990 ( .A(n6356), .ZN(n6362) );
  NAND2_X1 U7991 ( .A1(n6782), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6358) );
  OAI21_X1 U7992 ( .B1(n6782), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6358), .ZN(
        n6359) );
  AOI211_X1 U7993 ( .C1(n6360), .C2(n6359), .A(n6409), .B(n9740), .ZN(n6361)
         );
  AOI211_X1 U7994 ( .C1(n9395), .C2(n6782), .A(n6362), .B(n6361), .ZN(n6369)
         );
  INV_X1 U7995 ( .A(n6363), .ZN(n6364) );
  OAI21_X1 U7996 ( .B1(n9847), .B2(n6365), .A(n6364), .ZN(n6367) );
  INV_X1 U7997 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6785) );
  MUX2_X1 U7998 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6785), .S(n6782), .Z(n6366)
         );
  NAND2_X1 U7999 ( .A1(n6366), .A2(n6367), .ZN(n6414) );
  OAI211_X1 U8000 ( .C1(n6367), .C2(n6366), .A(n9891), .B(n6414), .ZN(n6368)
         );
  NAND2_X1 U8001 ( .A1(n6369), .A2(n6368), .ZN(P2_U3254) );
  AND2_X1 U8002 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n6370) );
  INV_X1 U8003 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8169) );
  INV_X1 U8004 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10185) );
  INV_X1 U8005 ( .A(n7795), .ZN(n6374) );
  AND2_X1 U8006 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6373) );
  NAND2_X1 U8007 ( .A1(n6374), .A2(n6373), .ZN(n7797) );
  INV_X1 U8008 ( .A(n7797), .ZN(n8043) );
  INV_X1 U8009 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n10125) );
  NAND2_X1 U8010 ( .A1(n4407), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U8011 ( .A1(n7798), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6375) );
  OAI211_X1 U8012 ( .C1(n7783), .C2(n10125), .A(n6376), .B(n6375), .ZN(n6377)
         );
  AOI21_X1 U8013 ( .B1(n8043), .B2(n7780), .A(n6377), .ZN(n8124) );
  NAND2_X1 U8014 ( .A1(n8271), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6378) );
  OAI21_X1 U8015 ( .B1(n8124), .B2(n8271), .A(n6378), .ZN(P2_U3581) );
  OAI21_X1 U8016 ( .B1(n6381), .B2(n6380), .A(n6379), .ZN(n6385) );
  INV_X1 U8017 ( .A(n8230), .ZN(n8250) );
  AOI22_X1 U8018 ( .A1(n8249), .A2(n6484), .B1(n8250), .B2(n6506), .ZN(n6383)
         );
  AND2_X1 U8019 ( .A1(P2_U3152), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9376) );
  AOI21_X1 U8020 ( .B1(n8011), .B2(P2_REG3_REG_1__SCAN_IN), .A(n9376), .ZN(
        n6382) );
  OAI211_X1 U8021 ( .C1(n9758), .C2(n8248), .A(n6383), .B(n6382), .ZN(n6384)
         );
  AOI21_X1 U8022 ( .B1(n8207), .B2(n6385), .A(n6384), .ZN(n6386) );
  INV_X1 U8023 ( .A(n6386), .ZN(P2_U3224) );
  AOI21_X1 U8024 ( .B1(n6270), .B2(n6388), .A(n6387), .ZN(n9629) );
  MUX2_X1 U8025 ( .A(n6389), .B(P1_REG1_REG_12__SCAN_IN), .S(n9624), .Z(n9628)
         );
  NOR2_X1 U8026 ( .A1(n9629), .A2(n9628), .ZN(n9627) );
  AOI21_X1 U8027 ( .B1(n6389), .B2(n6390), .A(n9627), .ZN(n6392) );
  INV_X1 U8028 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9505) );
  AOI22_X1 U8029 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(n6535), .B1(n6539), .B2(
        n9505), .ZN(n6391) );
  NOR2_X1 U8030 ( .A1(n6392), .A2(n6391), .ZN(n6534) );
  AOI21_X1 U8031 ( .B1(n6392), .B2(n6391), .A(n6534), .ZN(n6406) );
  INV_X1 U8032 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U8033 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3084), .ZN(n7253) );
  OAI21_X1 U8034 ( .B1(n9675), .B2(n6393), .A(n7253), .ZN(n6404) );
  NOR2_X1 U8035 ( .A1(n6394), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6395) );
  OR2_X1 U8036 ( .A1(n9624), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U8037 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9624), .ZN(n6398) );
  AND2_X1 U8038 ( .A1(n6399), .A2(n6398), .ZN(n9621) );
  NOR2_X1 U8039 ( .A1(n6539), .A2(n7358), .ZN(n6400) );
  AOI21_X1 U8040 ( .B1(n6539), .B2(n7358), .A(n6400), .ZN(n6401) );
  NOR2_X1 U8041 ( .A1(n6402), .A2(n6401), .ZN(n6538) );
  AOI211_X1 U8042 ( .C1(n6402), .C2(n6401), .A(n6538), .B(n9645), .ZN(n6403)
         );
  AOI211_X1 U8043 ( .C1(n9651), .C2(n6539), .A(n6404), .B(n6403), .ZN(n6405)
         );
  OAI21_X1 U8044 ( .B1(n6406), .B2(n9630), .A(n6405), .ZN(P1_U3254) );
  INV_X1 U8045 ( .A(n7687), .ZN(n6446) );
  AOI22_X1 U8046 ( .A1(n9652), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9367), .ZN(n6407) );
  OAI21_X1 U8047 ( .B1(n6446), .B2(n9369), .A(n6407), .ZN(P1_U3337) );
  NOR2_X1 U8048 ( .A1(n6911), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6408) );
  AOI21_X1 U8049 ( .B1(n6911), .B2(P2_REG2_REG_11__SCAN_IN), .A(n6408), .ZN(
        n6413) );
  AOI21_X1 U8050 ( .B1(n6782), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6409), .ZN(
        n9893) );
  OR2_X1 U8051 ( .A1(n6882), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6411) );
  NAND2_X1 U8052 ( .A1(n6882), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6410) );
  NAND2_X1 U8053 ( .A1(n6411), .A2(n6410), .ZN(n9894) );
  NOR2_X1 U8054 ( .A1(n9893), .A2(n9894), .ZN(n9892) );
  OAI21_X1 U8055 ( .B1(n6413), .B2(n6412), .A(n6528), .ZN(n6422) );
  INV_X1 U8056 ( .A(n6911), .ZN(n6529) );
  INV_X1 U8057 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10098) );
  MUX2_X1 U8058 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n10098), .S(n6882), .Z(n9884) );
  NAND2_X1 U8059 ( .A1(n6782), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6415) );
  NAND2_X1 U8060 ( .A1(n6415), .A2(n6414), .ZN(n9883) );
  NAND2_X1 U8061 ( .A1(n9884), .A2(n9883), .ZN(n9882) );
  OAI21_X1 U8062 ( .B1(n9899), .B2(n10098), .A(n9882), .ZN(n6417) );
  INV_X1 U8063 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6896) );
  MUX2_X1 U8064 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n6896), .S(n6911), .Z(n6416)
         );
  NAND2_X1 U8065 ( .A1(n6416), .A2(n6417), .ZN(n6520) );
  OAI211_X1 U8066 ( .C1(n6417), .C2(n6416), .A(n9891), .B(n6520), .ZN(n6420)
         );
  AND2_X1 U8067 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6418) );
  AOI21_X1 U8068 ( .B1(n9739), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6418), .ZN(
        n6419) );
  OAI211_X1 U8069 ( .C1(n9900), .C2(n6529), .A(n6420), .B(n6419), .ZN(n6421)
         );
  AOI21_X1 U8070 ( .B1(n9896), .B2(n6422), .A(n6421), .ZN(n6423) );
  INV_X1 U8071 ( .A(n6423), .ZN(P2_U3256) );
  OAI21_X1 U8072 ( .B1(n6427), .B2(n6425), .A(n6424), .ZN(n6434) );
  NOR3_X1 U8073 ( .A1(n6427), .A2(n8255), .A3(n6426), .ZN(n6428) );
  OAI21_X1 U8074 ( .B1(n6428), .B2(n8249), .A(n8282), .ZN(n6432) );
  OAI21_X1 U8075 ( .B1(n8253), .B2(n6654), .A(n6429), .ZN(n6430) );
  AOI21_X1 U8076 ( .B1(n8250), .B2(n4535), .A(n6430), .ZN(n6431) );
  OAI211_X1 U8077 ( .C1(n9808), .C2(n8248), .A(n6432), .B(n6431), .ZN(n6433)
         );
  AOI21_X1 U8078 ( .B1(n6434), .B2(n8207), .A(n6433), .ZN(n6435) );
  INV_X1 U8079 ( .A(n6435), .ZN(P2_U3241) );
  INV_X1 U8080 ( .A(n7367), .ZN(n6441) );
  NAND2_X1 U8081 ( .A1(n6437), .A2(n6436), .ZN(n6438) );
  NAND2_X1 U8082 ( .A1(n6438), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6439) );
  XNOR2_X1 U8083 ( .A(n6439), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7368) );
  INV_X1 U8084 ( .A(n7368), .ZN(n7314) );
  OAI222_X1 U8085 ( .A1(n7404), .A2(n6440), .B1(n8131), .B2(n6441), .C1(
        P2_U3152), .C2(n7314), .ZN(P2_U3343) );
  INV_X1 U8086 ( .A(n9638), .ZN(n8904) );
  OAI222_X1 U8087 ( .A1(n8904), .A2(P1_U3084), .B1(n9369), .B2(n6441), .C1(
        n10060), .C2(n9371), .ZN(P1_U3338) );
  NAND2_X1 U8088 ( .A1(n6442), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6443) );
  MUX2_X1 U8089 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6443), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6444) );
  AND2_X1 U8090 ( .A1(n6444), .A2(n6499), .ZN(n8291) );
  INV_X1 U8091 ( .A(n8291), .ZN(n8286) );
  OAI222_X1 U8092 ( .A1(P2_U3152), .A2(n8286), .B1(n8131), .B2(n6446), .C1(
        n6445), .C2(n7404), .ZN(P2_U3342) );
  XNOR2_X1 U8093 ( .A(n7795), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8361) );
  INV_X1 U8094 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10043) );
  NAND2_X1 U8095 ( .A1(n7798), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6448) );
  INV_X1 U8096 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n10086) );
  OR2_X1 U8097 ( .A1(n7783), .A2(n10086), .ZN(n6447) );
  OAI211_X1 U8098 ( .C1(n7802), .C2(n10043), .A(n6448), .B(n6447), .ZN(n6449)
         );
  INV_X1 U8099 ( .A(n8240), .ZN(n6450) );
  NAND2_X1 U8100 ( .A1(n6450), .A2(n8264), .ZN(n6451) );
  OAI21_X1 U8101 ( .B1(n5722), .B2(n8264), .A(n6451), .ZN(P2_U3579) );
  OAI21_X1 U8102 ( .B1(n5004), .B2(n6453), .A(n6452), .ZN(n6594) );
  INV_X1 U8103 ( .A(n6594), .ZN(n6454) );
  MUX2_X1 U8104 ( .A(n8857), .B(n6454), .S(n6274), .Z(n6455) );
  AOI21_X1 U8105 ( .B1(n8936), .B2(n5201), .A(n5773), .ZN(n9533) );
  NOR2_X1 U8106 ( .A1(n9533), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n9532) );
  AOI211_X1 U8107 ( .C1(n6455), .C2(n6628), .A(n9532), .B(n8846), .ZN(n9551)
         );
  AOI22_X1 U8108 ( .A1(n9581), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3084), .ZN(n6466) );
  OAI211_X1 U8109 ( .C1(n6458), .C2(n6457), .A(n9670), .B(n6456), .ZN(n6465)
         );
  OAI211_X1 U8110 ( .C1(n6461), .C2(n6460), .A(n9663), .B(n6459), .ZN(n6464)
         );
  NAND2_X1 U8111 ( .A1(n9651), .A2(n6462), .ZN(n6463) );
  NAND4_X1 U8112 ( .A1(n6466), .A2(n6465), .A3(n6464), .A4(n6463), .ZN(n6467)
         );
  OR2_X1 U8113 ( .A1(n9551), .A2(n6467), .ZN(P1_U3243) );
  NAND2_X1 U8114 ( .A1(n8846), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6468) );
  OAI21_X1 U8115 ( .B1(n9013), .B2(n8846), .A(n6468), .ZN(P1_U3584) );
  XOR2_X1 U8116 ( .A(n6469), .B(n6470), .Z(n6474) );
  INV_X1 U8117 ( .A(n6749), .ZN(n8848) );
  AOI22_X1 U8118 ( .A1(n8833), .A2(n6625), .B1(n8807), .B2(n8848), .ZN(n6471)
         );
  OAI21_X1 U8119 ( .B1(n7063), .B2(n6691), .A(n6471), .ZN(n6472) );
  AOI21_X1 U8120 ( .B1(n8819), .B2(n5237), .A(n6472), .ZN(n6473) );
  OAI21_X1 U8121 ( .B1(n6474), .B2(n8825), .A(n6473), .ZN(P1_U3235) );
  XNOR2_X1 U8122 ( .A(n6476), .B(n6475), .ZN(n6478) );
  XNOR2_X1 U8123 ( .A(n6478), .B(n6477), .ZN(n6483) );
  NAND2_X1 U8124 ( .A1(n8833), .A2(n6634), .ZN(n6480) );
  NAND2_X1 U8125 ( .A1(n8807), .A2(n6679), .ZN(n6479) );
  OAI211_X1 U8126 ( .C1(n7063), .C2(n6664), .A(n6480), .B(n6479), .ZN(n6481)
         );
  AOI21_X1 U8127 ( .B1(n8819), .B2(n7622), .A(n6481), .ZN(n6482) );
  OAI21_X1 U8128 ( .B1(n6483), .B2(n8825), .A(n6482), .ZN(P1_U3220) );
  NAND2_X1 U8129 ( .A1(n6484), .A2(n9759), .ZN(n7962) );
  NAND2_X1 U8130 ( .A1(n9749), .A2(n7962), .ZN(n9781) );
  INV_X1 U8131 ( .A(n9781), .ZN(n6498) );
  XNOR2_X1 U8132 ( .A(n8007), .B(n6486), .ZN(n6485) );
  NOR2_X1 U8133 ( .A1(n6486), .A2(n8385), .ZN(n6972) );
  INV_X1 U8134 ( .A(n6551), .ZN(n6487) );
  NOR2_X1 U8135 ( .A1(n6552), .A2(n6487), .ZN(n6488) );
  NAND2_X1 U8136 ( .A1(n6567), .A2(n6489), .ZN(n6490) );
  OAI21_X2 U8137 ( .B1(n6978), .B2(n6972), .A(n9768), .ZN(n8541) );
  NAND2_X1 U8138 ( .A1(n7964), .A2(n7833), .ZN(n7817) );
  AOI22_X1 U8139 ( .A1(n9781), .A2(n9748), .B1(n9752), .B2(n6505), .ZN(n9783)
         );
  NAND2_X1 U8140 ( .A1(n9756), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6491) );
  AOI21_X1 U8141 ( .B1(n9783), .B2(n6491), .A(n8535), .ZN(n6492) );
  AOI21_X1 U8142 ( .B1(n8518), .B2(P2_REG2_REG_0__SCAN_IN), .A(n6492), .ZN(
        n6497) );
  NOR2_X1 U8143 ( .A1(n8393), .A2(n6493), .ZN(n6494) );
  AND2_X1 U8144 ( .A1(n6567), .A2(n6494), .ZN(n7204) );
  INV_X1 U8145 ( .A(n8521), .ZN(n8562) );
  NAND2_X1 U8146 ( .A1(n8562), .A2(n8538), .ZN(n9765) );
  NAND2_X1 U8147 ( .A1(n9765), .A2(n9779), .ZN(n6496) );
  OAI211_X1 U8148 ( .C1(n6498), .C2(n8541), .A(n6497), .B(n6496), .ZN(P2_U3296) );
  INV_X1 U8149 ( .A(n7690), .ZN(n6502) );
  NAND2_X1 U8150 ( .A1(n6499), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6500) );
  XNOR2_X1 U8151 ( .A(n6500), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8308) );
  INV_X1 U8152 ( .A(n8308), .ZN(n8303) );
  OAI222_X1 U8153 ( .A1(n7404), .A2(n6501), .B1(n8131), .B2(n6502), .C1(n8303), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  OAI222_X1 U8154 ( .A1(n9371), .A2(n6503), .B1(n9369), .B2(n6502), .C1(
        P1_U3084), .C2(n9667), .ZN(P1_U3336) );
  NAND2_X1 U8155 ( .A1(n7843), .A2(n9749), .ZN(n7961) );
  NAND2_X1 U8156 ( .A1(n7961), .A2(n7959), .ZN(n7835) );
  NAND2_X1 U8157 ( .A1(n6506), .A2(n9789), .ZN(n7845) );
  NAND2_X1 U8158 ( .A1(n7842), .A2(n7845), .ZN(n6560) );
  INV_X1 U8159 ( .A(n6560), .ZN(n7963) );
  XNOR2_X1 U8160 ( .A(n7835), .B(n7963), .ZN(n6509) );
  NAND2_X1 U8161 ( .A1(n8284), .A2(n9752), .ZN(n6508) );
  NAND2_X1 U8162 ( .A1(n6505), .A2(n9751), .ZN(n6507) );
  AND2_X1 U8163 ( .A1(n6508), .A2(n6507), .ZN(n8009) );
  OAI21_X1 U8164 ( .B1(n6509), .B2(n8529), .A(n8009), .ZN(n9790) );
  INV_X1 U8165 ( .A(n9790), .ZN(n6519) );
  INV_X1 U8166 ( .A(n9763), .ZN(n6510) );
  OAI21_X1 U8167 ( .B1(n6511), .B2(n6560), .A(n6555), .ZN(n9792) );
  INV_X1 U8168 ( .A(n8541), .ZN(n9764) );
  NAND2_X1 U8169 ( .A1(n9758), .A2(n9759), .ZN(n9757) );
  INV_X1 U8170 ( .A(n9789), .ZN(n8020) );
  NAND2_X1 U8171 ( .A1(n9757), .A2(n8020), .ZN(n6512) );
  NAND2_X1 U8172 ( .A1(n6512), .A2(n9816), .ZN(n6513) );
  OR2_X1 U8173 ( .A1(n6513), .A2(n6573), .ZN(n9788) );
  INV_X1 U8174 ( .A(n9788), .ZN(n6514) );
  AOI22_X1 U8175 ( .A1(n6514), .A2(n7204), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n9756), .ZN(n6516) );
  OR2_X1 U8176 ( .A1(n9768), .A2(n10101), .ZN(n6515) );
  OAI211_X1 U8177 ( .C1(n8538), .C2(n9789), .A(n6516), .B(n6515), .ZN(n6517)
         );
  AOI21_X1 U8178 ( .B1(n9792), .B2(n9764), .A(n6517), .ZN(n6518) );
  OAI21_X1 U8179 ( .B1(n6519), .B2(n8535), .A(n6518), .ZN(P2_U3294) );
  INV_X1 U8180 ( .A(n6520), .ZN(n6521) );
  AOI21_X1 U8181 ( .B1(n6911), .B2(P2_REG1_REG_11__SCAN_IN), .A(n6521), .ZN(
        n6523) );
  INV_X1 U8182 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9851) );
  MUX2_X1 U8183 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n9851), .S(n7016), .Z(n6522)
         );
  NAND2_X1 U8184 ( .A1(n6523), .A2(n6522), .ZN(n6836) );
  OAI21_X1 U8185 ( .B1(n6523), .B2(n6522), .A(n6836), .ZN(n6527) );
  NAND2_X1 U8186 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7037) );
  INV_X1 U8187 ( .A(n7037), .ZN(n6526) );
  INV_X1 U8188 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n6524) );
  NOR2_X1 U8189 ( .A1(n9888), .A2(n6524), .ZN(n6525) );
  AOI211_X1 U8190 ( .C1(n9891), .C2(n6527), .A(n6526), .B(n6525), .ZN(n6533)
         );
  INV_X1 U8191 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7190) );
  XNOR2_X1 U8192 ( .A(n7016), .B(n7190), .ZN(n6531) );
  INV_X1 U8193 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6900) );
  NAND2_X1 U8194 ( .A1(n6530), .A2(n6531), .ZN(n6844) );
  OAI211_X1 U8195 ( .C1(n6531), .C2(n6530), .A(n9896), .B(n6844), .ZN(n6532)
         );
  OAI211_X1 U8196 ( .C1(n9900), .C2(n6838), .A(n6533), .B(n6532), .ZN(P2_U3257) );
  AOI21_X1 U8197 ( .B1(n9505), .B2(n6535), .A(n6534), .ZN(n6537) );
  INV_X1 U8198 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9498) );
  AOI22_X1 U8199 ( .A1(n6541), .A2(n9498), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n8900), .ZN(n6536) );
  NOR2_X1 U8200 ( .A1(n6537), .A2(n6536), .ZN(n8889) );
  AOI21_X1 U8201 ( .B1(n6537), .B2(n6536), .A(n8889), .ZN(n6546) );
  AOI21_X1 U8202 ( .B1(n6539), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6538), .ZN(
        n8901) );
  OAI21_X1 U8203 ( .B1(n6540), .B2(n9262), .A(n8902), .ZN(n6544) );
  INV_X1 U8204 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10172) );
  NAND2_X1 U8205 ( .A1(n9651), .A2(n6541), .ZN(n6542) );
  NAND2_X1 U8206 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n7396) );
  OAI211_X1 U8207 ( .C1(n10172), .C2(n9675), .A(n6542), .B(n7396), .ZN(n6543)
         );
  AOI21_X1 U8208 ( .B1(n6544), .B2(n9663), .A(n6543), .ZN(n6545) );
  OAI21_X1 U8209 ( .B1(n6546), .B2(n9630), .A(n6545), .ZN(P1_U3255) );
  NAND2_X1 U8210 ( .A1(n6548), .A2(n6547), .ZN(n6550) );
  NOR2_X2 U8211 ( .A1(n6978), .A2(n9829), .ZN(n8644) );
  OR2_X1 U8212 ( .A1(n6506), .A2(n8020), .ZN(n6554) );
  OR2_X1 U8213 ( .A1(n8284), .A2(n4812), .ZN(n6556) );
  INV_X1 U8214 ( .A(n8283), .ZN(n6557) );
  NAND2_X1 U8215 ( .A1(n6557), .A2(n8209), .ZN(n7829) );
  NAND2_X1 U8216 ( .A1(n6612), .A2(n7966), .ZN(n6559) );
  INV_X1 U8217 ( .A(n9803), .ZN(n8209) );
  OR2_X1 U8218 ( .A1(n8283), .A2(n8209), .ZN(n6558) );
  NAND2_X1 U8219 ( .A1(n8282), .A2(n6587), .ZN(n7826) );
  NAND2_X1 U8220 ( .A1(n7830), .A2(n7826), .ZN(n7965) );
  INV_X1 U8221 ( .A(n7965), .ZN(n6644) );
  XNOR2_X1 U8222 ( .A(n6646), .B(n6644), .ZN(n6591) );
  OAI21_X1 U8223 ( .B1(n7835), .B2(n6560), .A(n7842), .ZN(n6576) );
  OR2_X1 U8224 ( .A1(n8284), .A2(n9796), .ZN(n7828) );
  INV_X1 U8225 ( .A(n7966), .ZN(n6562) );
  NAND2_X1 U8226 ( .A1(n6614), .A2(n7823), .ZN(n6647) );
  XNOR2_X1 U8227 ( .A(n6647), .B(n7965), .ZN(n6563) );
  AOI222_X1 U8228 ( .A1(n9748), .A2(n6563), .B1(n8281), .B2(n9752), .C1(n8283), 
        .C2(n9751), .ZN(n6584) );
  NAND2_X1 U8229 ( .A1(n6573), .A2(n9796), .ZN(n6617) );
  OR2_X1 U8230 ( .A1(n6617), .A2(n8209), .ZN(n6564) );
  INV_X1 U8231 ( .A(n6652), .ZN(n6653) );
  AOI211_X1 U8232 ( .C1(n6643), .C2(n6564), .A(n9833), .B(n6653), .ZN(n6582)
         );
  AOI21_X1 U8233 ( .B1(n9815), .B2(n6643), .A(n6582), .ZN(n6565) );
  OAI211_X1 U8234 ( .C1(n8644), .C2(n6591), .A(n6584), .B(n6565), .ZN(n6569)
         );
  NAND2_X1 U8235 ( .A1(n6569), .A2(n9853), .ZN(n6566) );
  OAI21_X1 U8236 ( .B1(n9853), .B2(n5956), .A(n6566), .ZN(P2_U3525) );
  INV_X1 U8237 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6571) );
  NAND2_X1 U8238 ( .A1(n6569), .A2(n4405), .ZN(n6570) );
  OAI21_X1 U8239 ( .B1(n4405), .B2(n6571), .A(n6570), .ZN(P2_U3466) );
  XNOR2_X1 U8240 ( .A(n6572), .B(n7836), .ZN(n9798) );
  INV_X1 U8241 ( .A(n7204), .ZN(n7334) );
  OAI211_X1 U8242 ( .C1(n6573), .C2(n9796), .A(n6617), .B(n9816), .ZN(n9794)
         );
  AOI22_X1 U8243 ( .A1(n8535), .A2(P2_REG2_REG_3__SCAN_IN), .B1(n9756), .B2(
        n6574), .ZN(n6575) );
  OAI21_X1 U8244 ( .B1(n7334), .B2(n9794), .A(n6575), .ZN(n6580) );
  XNOR2_X1 U8245 ( .A(n6576), .B(n7836), .ZN(n6578) );
  AOI21_X1 U8246 ( .B1(n6578), .B2(n9748), .A(n6577), .ZN(n9795) );
  NOR2_X1 U8247 ( .A1(n9795), .A2(n8535), .ZN(n6579) );
  AOI211_X1 U8248 ( .C1(n8566), .C2(n4812), .A(n6580), .B(n6579), .ZN(n6581)
         );
  OAI21_X1 U8249 ( .B1(n8541), .B2(n9798), .A(n6581), .ZN(P2_U3293) );
  NAND2_X1 U8250 ( .A1(n6582), .A2(n8385), .ZN(n6583) );
  OAI211_X1 U8251 ( .C1(n8556), .C2(n6585), .A(n6584), .B(n6583), .ZN(n6589)
         );
  OAI22_X1 U8252 ( .A1(n8538), .A2(n6587), .B1(n9768), .B2(n6586), .ZN(n6588)
         );
  AOI21_X1 U8253 ( .B1(n6589), .B2(n9768), .A(n6588), .ZN(n6590) );
  OAI21_X1 U8254 ( .B1(n6591), .B2(n8541), .A(n6590), .ZN(P2_U3291) );
  INV_X1 U8255 ( .A(n8819), .ZN(n8836) );
  OAI22_X1 U8256 ( .A1(n7063), .A2(n9538), .B1(n6592), .B2(n8830), .ZN(n6593)
         );
  AOI21_X1 U8257 ( .B1(n8812), .B2(n6594), .A(n6593), .ZN(n6595) );
  OAI21_X1 U8258 ( .B1(n6762), .B2(n8836), .A(n6595), .ZN(P1_U3230) );
  XNOR2_X1 U8259 ( .A(n6597), .B(n6596), .ZN(n6598) );
  NAND2_X1 U8260 ( .A1(n6598), .A2(n8812), .ZN(n6602) );
  INV_X1 U8261 ( .A(n7676), .ZN(n8847) );
  NOR2_X1 U8262 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6599), .ZN(n8865) );
  INV_X1 U8263 ( .A(n6679), .ZN(n7625) );
  OAI22_X1 U8264 ( .A1(n8831), .A2(P1_REG3_REG_3__SCAN_IN), .B1(n7625), .B2(
        n8816), .ZN(n6600) );
  AOI211_X1 U8265 ( .C1(n8807), .C2(n8847), .A(n8865), .B(n6600), .ZN(n6601)
         );
  OAI211_X1 U8266 ( .C1(n9681), .C2(n8836), .A(n6602), .B(n6601), .ZN(P1_U3216) );
  AOI21_X1 U8267 ( .B1(n6603), .B2(n6604), .A(n8825), .ZN(n6605) );
  NAND2_X1 U8268 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n9542) );
  INV_X1 U8269 ( .A(n9542), .ZN(n6607) );
  OAI22_X1 U8270 ( .A1(n8831), .A2(n6757), .B1(n6749), .B2(n8816), .ZN(n6606)
         );
  AOI211_X1 U8271 ( .C1(n8807), .C2(n8845), .A(n6607), .B(n6606), .ZN(n6608)
         );
  OAI211_X1 U8272 ( .C1(n6758), .C2(n8836), .A(n6609), .B(n6608), .ZN(P1_U3228) );
  INV_X1 U8273 ( .A(n9053), .ZN(n6610) );
  NAND2_X1 U8274 ( .A1(n6610), .A2(P1_U4006), .ZN(n6611) );
  OAI21_X1 U8275 ( .B1(n5715), .B2(P1_U4006), .A(n6611), .ZN(P1_U3582) );
  XNOR2_X1 U8276 ( .A(n7966), .B(n6612), .ZN(n9807) );
  INV_X1 U8277 ( .A(n9807), .ZN(n6622) );
  OAI211_X1 U8278 ( .C1(n6613), .C2(n6562), .A(n9748), .B(n6614), .ZN(n6616)
         );
  AOI22_X1 U8279 ( .A1(n9752), .A2(n8282), .B1(n8284), .B2(n9751), .ZN(n6615)
         );
  NAND2_X1 U8280 ( .A1(n6616), .A2(n6615), .ZN(n9805) );
  XNOR2_X1 U8281 ( .A(n6617), .B(n8209), .ZN(n9804) );
  OAI22_X1 U8282 ( .A1(n9768), .A2(n6171), .B1(n8210), .B2(n8556), .ZN(n6618)
         );
  AOI21_X1 U8283 ( .B1(n8566), .B2(n8209), .A(n6618), .ZN(n6619) );
  OAI21_X1 U8284 ( .B1(n8562), .B2(n9804), .A(n6619), .ZN(n6620) );
  AOI21_X1 U8285 ( .B1(n9805), .B2(n8555), .A(n6620), .ZN(n6621) );
  OAI21_X1 U8286 ( .B1(n6622), .B2(n8541), .A(n6621), .ZN(P2_U3292) );
  NAND2_X1 U8287 ( .A1(n5170), .A2(n8929), .ZN(n6624) );
  AND2_X1 U8288 ( .A1(n6634), .A2(n6626), .ZN(n6627) );
  NAND2_X1 U8289 ( .A1(n6627), .A2(n6632), .ZN(n6678) );
  OAI21_X1 U8290 ( .B1(n6632), .B2(n6627), .A(n6678), .ZN(n6661) );
  INV_X1 U8291 ( .A(n7610), .ZN(n6629) );
  NAND2_X1 U8292 ( .A1(n5738), .A2(n9087), .ZN(n6631) );
  OR2_X1 U8293 ( .A1(n7612), .A2(n7013), .ZN(n6630) );
  XNOR2_X1 U8294 ( .A(n7491), .B(n6681), .ZN(n6633) );
  AOI222_X1 U8295 ( .A1(n6634), .A2(n9253), .B1(n6679), .B2(n9254), .C1(n9470), 
        .C2(n6633), .ZN(n6660) );
  NAND2_X1 U8296 ( .A1(n6636), .A2(n6762), .ZN(n6687) );
  OAI211_X1 U8297 ( .C1(n6762), .C2(n6636), .A(n9711), .B(n6687), .ZN(n6665)
         );
  INV_X1 U8298 ( .A(n6665), .ZN(n6637) );
  AOI21_X1 U8299 ( .B1(n7622), .B2(n9709), .A(n6637), .ZN(n6638) );
  OAI211_X1 U8300 ( .C1(n9687), .C2(n6661), .A(n6660), .B(n6638), .ZN(n6640)
         );
  NAND2_X1 U8301 ( .A1(n6640), .A2(n9737), .ZN(n6639) );
  OAI21_X1 U8302 ( .B1(n9737), .B2(n5186), .A(n6639), .ZN(P1_U3524) );
  INV_X1 U8303 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6642) );
  NAND2_X1 U8304 ( .A1(n6640), .A2(n9729), .ZN(n6641) );
  OAI21_X1 U8305 ( .B1(n9729), .B2(n6642), .A(n6641), .ZN(P1_U3457) );
  NOR2_X1 U8306 ( .A1(n8282), .A2(n6643), .ZN(n6645) );
  NAND2_X1 U8307 ( .A1(n8281), .A2(n9808), .ZN(n7848) );
  INV_X1 U8308 ( .A(n6726), .ZN(n7969) );
  XNOR2_X1 U8309 ( .A(n6727), .B(n7969), .ZN(n9812) );
  INV_X1 U8310 ( .A(n9812), .ZN(n6659) );
  NAND2_X1 U8311 ( .A1(n6647), .A2(n7830), .ZN(n6648) );
  NAND2_X1 U8312 ( .A1(n6648), .A2(n7826), .ZN(n6650) );
  INV_X1 U8313 ( .A(n6650), .ZN(n6649) );
  NAND2_X1 U8314 ( .A1(n6649), .A2(n7969), .ZN(n6729) );
  AOI21_X1 U8315 ( .B1(n6726), .B2(n6650), .A(n4525), .ZN(n6651) );
  OAI222_X1 U8316 ( .A1(n8550), .A2(n6983), .B1(n8548), .B2(n4678), .C1(n8529), 
        .C2(n6651), .ZN(n9810) );
  INV_X1 U8317 ( .A(n9808), .ZN(n6728) );
  INV_X1 U8318 ( .A(n6731), .ZN(n6732) );
  OAI21_X1 U8319 ( .B1(n9808), .B2(n6653), .A(n6732), .ZN(n9809) );
  OAI22_X1 U8320 ( .A1(n9768), .A2(n6172), .B1(n6654), .B2(n8556), .ZN(n6655)
         );
  AOI21_X1 U8321 ( .B1(n8566), .B2(n6728), .A(n6655), .ZN(n6656) );
  OAI21_X1 U8322 ( .B1(n9809), .B2(n8562), .A(n6656), .ZN(n6657) );
  AOI21_X1 U8323 ( .B1(n9810), .B2(n8555), .A(n6657), .ZN(n6658) );
  OAI21_X1 U8324 ( .B1(n8541), .B2(n6659), .A(n6658), .ZN(P2_U3290) );
  INV_X1 U8325 ( .A(n6660), .ZN(n6668) );
  INV_X1 U8326 ( .A(n6696), .ZN(n6662) );
  AOI21_X1 U8327 ( .B1(n9473), .B2(n6662), .A(n6661), .ZN(n6667) );
  AND2_X1 U8328 ( .A1(n9678), .A2(n7612), .ZN(n6663) );
  OAI22_X1 U8329 ( .A1(n6665), .A2(n9087), .B1(n9476), .B2(n6664), .ZN(n6666)
         );
  NOR3_X1 U8330 ( .A1(n6668), .A2(n6667), .A3(n6666), .ZN(n6676) );
  INV_X1 U8331 ( .A(n6669), .ZN(n6670) );
  NAND2_X1 U8332 ( .A1(n6949), .A2(n6948), .ZN(n6672) );
  INV_X1 U8333 ( .A(n6673), .ZN(n6674) );
  AOI22_X1 U8334 ( .A1(n9264), .A2(n7622), .B1(n9223), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6675) );
  OAI21_X1 U8335 ( .B1(n6676), .B2(n9223), .A(n6675), .ZN(P1_U3290) );
  INV_X1 U8336 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9996) );
  NAND2_X1 U8337 ( .A1(n6625), .A2(n7622), .ZN(n6677) );
  AND2_X1 U8338 ( .A1(n6678), .A2(n6677), .ZN(n6680) );
  XNOR2_X1 U8339 ( .A(n6679), .B(n6712), .ZN(n6701) );
  NAND2_X1 U8340 ( .A1(n6680), .A2(n6701), .ZN(n6714) );
  OAI21_X1 U8341 ( .B1(n6680), .B2(n6701), .A(n6714), .ZN(n6697) );
  INV_X1 U8342 ( .A(n6697), .ZN(n6689) );
  INV_X1 U8343 ( .A(n9473), .ZN(n9719) );
  OAI22_X1 U8344 ( .A1(n6592), .A2(n9465), .B1(n6749), .B2(n9467), .ZN(n6686)
         );
  NAND2_X1 U8345 ( .A1(n6592), .A2(n7622), .ZN(n6682) );
  NAND2_X1 U8346 ( .A1(n6683), .A2(n6682), .ZN(n7627) );
  XNOR2_X1 U8347 ( .A(n7627), .B(n6701), .ZN(n6684) );
  NOR2_X1 U8348 ( .A1(n6684), .A2(n9234), .ZN(n6685) );
  AOI211_X1 U8349 ( .C1(n9719), .C2(n6697), .A(n6686), .B(n6685), .ZN(n6700)
         );
  AOI21_X1 U8350 ( .B1(n5237), .B2(n6687), .A(n6829), .ZN(n6695) );
  AOI22_X1 U8351 ( .A1(n6695), .A2(n9711), .B1(n5237), .B2(n9709), .ZN(n6688)
         );
  OAI211_X1 U8352 ( .C1(n6689), .C2(n9715), .A(n6700), .B(n6688), .ZN(n9345)
         );
  NAND2_X1 U8353 ( .A1(n9345), .A2(n9729), .ZN(n6690) );
  OAI21_X1 U8354 ( .B1(n9729), .B2(n9996), .A(n6690), .ZN(P1_U3460) );
  OAI22_X1 U8355 ( .A1(n9269), .A2(n6692), .B1(n6691), .B2(n9476), .ZN(n6694)
         );
  NOR2_X1 U8356 ( .A1(n9475), .A2(n6712), .ZN(n6693) );
  AOI211_X1 U8357 ( .C1(n6695), .C2(n9461), .A(n6694), .B(n6693), .ZN(n6699)
         );
  NAND2_X1 U8358 ( .A1(n9269), .A2(n6696), .ZN(n9245) );
  INV_X1 U8359 ( .A(n9245), .ZN(n9462) );
  NAND2_X1 U8360 ( .A1(n6697), .A2(n9462), .ZN(n6698) );
  OAI211_X1 U8361 ( .C1(n6700), .C2(n9223), .A(n6699), .B(n6698), .ZN(P1_U3289) );
  INV_X1 U8362 ( .A(n6701), .ZN(n7490) );
  NAND2_X1 U8363 ( .A1(n7627), .A2(n7490), .ZN(n6702) );
  NAND2_X1 U8364 ( .A1(n7625), .A2(n5237), .ZN(n7623) );
  NAND2_X1 U8365 ( .A1(n6702), .A2(n7623), .ZN(n7446) );
  NAND2_X1 U8366 ( .A1(n6749), .A2(n6832), .ZN(n7630) );
  NAND2_X1 U8367 ( .A1(n8848), .A2(n9681), .ZN(n7445) );
  NAND2_X1 U8368 ( .A1(n7630), .A2(n7445), .ZN(n6715) );
  INV_X1 U8369 ( .A(n6715), .ZN(n6823) );
  NAND2_X1 U8370 ( .A1(n7676), .A2(n6812), .ZN(n7632) );
  INV_X1 U8371 ( .A(n7632), .ZN(n6703) );
  NAND2_X1 U8372 ( .A1(n6748), .A2(n9689), .ZN(n7633) );
  NAND2_X1 U8373 ( .A1(n8845), .A2(n7681), .ZN(n7447) );
  INV_X1 U8374 ( .A(n6718), .ZN(n6704) );
  XNOR2_X1 U8375 ( .A(n7082), .B(n6704), .ZN(n6706) );
  OAI22_X1 U8376 ( .A1(n7676), .A2(n9465), .B1(n6943), .B2(n9467), .ZN(n6705)
         );
  AOI21_X1 U8377 ( .B1(n6706), .B2(n9470), .A(n6705), .ZN(n9693) );
  OAI22_X1 U8378 ( .A1(n9269), .A2(n6707), .B1(n7677), .B2(n9476), .ZN(n6711)
         );
  AOI21_X1 U8379 ( .B1(n6756), .B2(n9689), .A(n9723), .ZN(n6708) );
  NAND2_X1 U8380 ( .A1(n6708), .A2(n7078), .ZN(n9691) );
  INV_X1 U8381 ( .A(n9193), .ZN(n6709) );
  NOR2_X1 U8382 ( .A1(n9691), .A2(n6709), .ZN(n6710) );
  AOI211_X1 U8383 ( .C1(n9264), .C2(n9689), .A(n6711), .B(n6710), .ZN(n6725)
         );
  NAND2_X1 U8384 ( .A1(n7625), .A2(n6712), .ZN(n6713) );
  NAND2_X1 U8385 ( .A1(n6714), .A2(n6713), .ZN(n6821) );
  NAND2_X1 U8386 ( .A1(n6821), .A2(n6715), .ZN(n6820) );
  NAND2_X1 U8387 ( .A1(n6749), .A2(n9681), .ZN(n6716) );
  NAND2_X1 U8388 ( .A1(n6820), .A2(n6716), .ZN(n6742) );
  NAND2_X1 U8389 ( .A1(n7632), .A2(n7448), .ZN(n6745) );
  NAND2_X1 U8390 ( .A1(n7676), .A2(n6758), .ZN(n6717) );
  NAND2_X1 U8391 ( .A1(n6719), .A2(n6718), .ZN(n6720) );
  NAND2_X1 U8392 ( .A1(n6942), .A2(n6720), .ZN(n9688) );
  INV_X1 U8393 ( .A(n6721), .ZN(n6722) );
  NOR2_X1 U8394 ( .A1(n6722), .A2(n4581), .ZN(n6723) );
  OR2_X1 U8395 ( .A1(n9688), .A2(n9271), .ZN(n6724) );
  OAI211_X1 U8396 ( .C1(n9693), .C2(n9223), .A(n6725), .B(n6724), .ZN(P1_U3286) );
  NAND2_X1 U8397 ( .A1(n6955), .A2(n6983), .ZN(n7852) );
  XNOR2_X1 U8398 ( .A(n6956), .B(n6959), .ZN(n6855) );
  XNOR2_X1 U8399 ( .A(n6960), .B(n7971), .ZN(n6730) );
  INV_X1 U8400 ( .A(n6963), .ZN(n8280) );
  AOI222_X1 U8401 ( .A1(n9748), .A2(n6730), .B1(n8281), .B2(n9751), .C1(n8280), 
        .C2(n9752), .ZN(n6854) );
  OR2_X1 U8402 ( .A1(n6854), .A2(n8518), .ZN(n6737) );
  AOI21_X1 U8403 ( .B1(n6955), .B2(n6732), .A(n6989), .ZN(n6852) );
  NOR2_X1 U8404 ( .A1(n8538), .A2(n4536), .ZN(n6735) );
  OAI22_X1 U8405 ( .A1(n9768), .A2(n6174), .B1(n6733), .B2(n8556), .ZN(n6734)
         );
  AOI211_X1 U8406 ( .C1(n6852), .C2(n8521), .A(n6735), .B(n6734), .ZN(n6736)
         );
  OAI211_X1 U8407 ( .C1(n6855), .C2(n8541), .A(n6737), .B(n6736), .ZN(P2_U3289) );
  INV_X1 U8408 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6740) );
  INV_X1 U8409 ( .A(n7702), .ZN(n6741) );
  NAND2_X1 U8410 ( .A1(n6738), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6739) );
  XNOR2_X1 U8411 ( .A(n6739), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8314) );
  INV_X1 U8412 ( .A(n8314), .ZN(n8323) );
  OAI222_X1 U8413 ( .A1(n7404), .A2(n6740), .B1(n8131), .B2(n6741), .C1(
        P2_U3152), .C2(n8323), .ZN(P2_U3340) );
  INV_X1 U8414 ( .A(n8918), .ZN(n8921) );
  INV_X1 U8415 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10092) );
  OAI222_X1 U8416 ( .A1(n8921), .A2(P1_U3084), .B1(n9369), .B2(n6741), .C1(
        n10092), .C2(n9371), .ZN(P1_U3335) );
  OR2_X1 U8417 ( .A1(n6742), .A2(n6745), .ZN(n6743) );
  NAND2_X1 U8418 ( .A1(n6744), .A2(n6743), .ZN(n6747) );
  INV_X1 U8419 ( .A(n6747), .ZN(n6816) );
  XNOR2_X1 U8420 ( .A(n6746), .B(n6745), .ZN(n6753) );
  NAND2_X1 U8421 ( .A1(n6747), .A2(n9719), .ZN(n6752) );
  OAI22_X1 U8422 ( .A1(n6749), .A2(n9465), .B1(n6748), .B2(n9467), .ZN(n6750)
         );
  INV_X1 U8423 ( .A(n6750), .ZN(n6751) );
  OAI211_X1 U8424 ( .C1(n9234), .C2(n6753), .A(n6752), .B(n6751), .ZN(n6811)
         );
  MUX2_X1 U8425 ( .A(n6811), .B(P1_REG2_REG_4__SCAN_IN), .S(n9223), .Z(n6754)
         );
  INV_X1 U8426 ( .A(n6754), .ZN(n6761) );
  NAND2_X1 U8427 ( .A1(n6828), .A2(n6812), .ZN(n6755) );
  AND2_X1 U8428 ( .A1(n6756), .A2(n6755), .ZN(n6813) );
  OAI22_X1 U8429 ( .A1(n9475), .A2(n6758), .B1(n6757), .B2(n9476), .ZN(n6759)
         );
  AOI21_X1 U8430 ( .B1(n6813), .B2(n9461), .A(n6759), .ZN(n6760) );
  OAI211_X1 U8431 ( .C1(n6816), .C2(n9245), .A(n6761), .B(n6760), .ZN(P1_U3287) );
  OAI22_X1 U8432 ( .A1(n9269), .A2(n5201), .B1(n9538), .B2(n9476), .ZN(n6764)
         );
  AOI21_X1 U8433 ( .B1(n9239), .B2(n9475), .A(n6762), .ZN(n6763) );
  AOI211_X1 U8434 ( .C1(n9269), .C2(n6765), .A(n6764), .B(n6763), .ZN(n6766)
         );
  INV_X1 U8435 ( .A(n6766), .ZN(P1_U3291) );
  NAND2_X1 U8436 ( .A1(n6768), .A2(n6767), .ZN(n6778) );
  NAND2_X1 U8437 ( .A1(n6770), .A2(n7787), .ZN(n6773) );
  AOI22_X1 U8438 ( .A1(n7703), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7714), .B2(
        n6771), .ZN(n6772) );
  NAND2_X1 U8439 ( .A1(n6773), .A2(n6772), .ZN(n9814) );
  XNOR2_X1 U8440 ( .A(n9814), .B(n8114), .ZN(n6774) );
  NOR2_X1 U8441 ( .A1(n6963), .A2(n5905), .ZN(n6775) );
  NAND2_X1 U8442 ( .A1(n6774), .A2(n6775), .ZN(n6793) );
  INV_X1 U8443 ( .A(n6774), .ZN(n6779) );
  INV_X1 U8444 ( .A(n6775), .ZN(n6776) );
  NAND2_X1 U8445 ( .A1(n6779), .A2(n6776), .ZN(n6777) );
  AND2_X1 U8446 ( .A1(n6793), .A2(n6777), .ZN(n6862) );
  INV_X1 U8447 ( .A(n6795), .ZN(n6864) );
  NOR3_X1 U8448 ( .A1(n6779), .A2(n6963), .A3(n8255), .ZN(n6780) );
  AOI21_X1 U8449 ( .B1(n6864), .B2(n8207), .A(n6780), .ZN(n6810) );
  NAND2_X1 U8450 ( .A1(n6781), .A2(n7787), .ZN(n6784) );
  AOI22_X1 U8451 ( .A1(n7703), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7714), .B2(
        n6782), .ZN(n6783) );
  NAND2_X1 U8452 ( .A1(n6784), .A2(n6783), .ZN(n7112) );
  XNOR2_X1 U8453 ( .A(n7112), .B(n5934), .ZN(n6891) );
  NAND2_X1 U8454 ( .A1(n4401), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6792) );
  OR2_X1 U8455 ( .A1(n7802), .A2(n6785), .ZN(n6791) );
  INV_X1 U8456 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U8457 ( .A1(n6787), .A2(n6786), .ZN(n6788) );
  NAND2_X1 U8458 ( .A1(n6798), .A2(n6788), .ZN(n6968) );
  OR2_X1 U8459 ( .A1(n7768), .A2(n6968), .ZN(n6790) );
  INV_X1 U8460 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6969) );
  OR2_X1 U8461 ( .A1(n7771), .A2(n6969), .ZN(n6789) );
  NOR2_X1 U8462 ( .A1(n7117), .A2(n5905), .ZN(n6889) );
  XNOR2_X1 U8463 ( .A(n6891), .B(n6889), .ZN(n6809) );
  AND2_X1 U8464 ( .A1(n6809), .A2(n6793), .ZN(n6794) );
  NOR2_X1 U8465 ( .A1(n6893), .A2(n8263), .ZN(n6807) );
  AND2_X1 U8466 ( .A1(n7112), .A2(n8259), .ZN(n6806) );
  OAI21_X1 U8467 ( .B1(n8253), .B2(n6968), .A(n6796), .ZN(n6805) );
  NAND2_X1 U8468 ( .A1(n4401), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6803) );
  OR2_X1 U8469 ( .A1(n7802), .A2(n10098), .ZN(n6802) );
  NAND2_X1 U8470 ( .A1(n6798), .A2(n6797), .ZN(n6799) );
  NAND2_X1 U8471 ( .A1(n6898), .A2(n6799), .ZN(n7121) );
  OR2_X1 U8472 ( .A1(n7768), .A2(n7121), .ZN(n6801) );
  INV_X1 U8473 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7122) );
  OR2_X1 U8474 ( .A1(n7771), .A2(n7122), .ZN(n6800) );
  OAI22_X1 U8475 ( .A1(n6963), .A2(n8231), .B1(n8230), .B2(n7161), .ZN(n6804)
         );
  NOR4_X1 U8476 ( .A1(n6807), .A2(n6806), .A3(n6805), .A4(n6804), .ZN(n6808)
         );
  OAI21_X1 U8477 ( .B1(n6810), .B2(n6809), .A(n6808), .ZN(P2_U3233) );
  INV_X1 U8478 ( .A(n6811), .ZN(n6815) );
  AOI22_X1 U8479 ( .A1(n6813), .A2(n9711), .B1(n6812), .B2(n9709), .ZN(n6814)
         );
  OAI211_X1 U8480 ( .C1(n6816), .C2(n9715), .A(n6815), .B(n6814), .ZN(n6818)
         );
  NAND2_X1 U8481 ( .A1(n6818), .A2(n9737), .ZN(n6817) );
  OAI21_X1 U8482 ( .B1(n9737), .B2(n6259), .A(n6817), .ZN(P1_U3527) );
  NAND2_X1 U8483 ( .A1(n6818), .A2(n9729), .ZN(n6819) );
  OAI21_X1 U8484 ( .B1(n9729), .B2(n5270), .A(n6819), .ZN(P1_U3466) );
  OAI21_X1 U8485 ( .B1(n6821), .B2(n6715), .A(n6820), .ZN(n9685) );
  INV_X1 U8486 ( .A(n9685), .ZN(n6835) );
  OAI21_X1 U8487 ( .B1(n6823), .B2(n7446), .A(n6822), .ZN(n6825) );
  OAI22_X1 U8488 ( .A1(n7625), .A2(n9465), .B1(n7676), .B2(n9467), .ZN(n6824)
         );
  AOI21_X1 U8489 ( .B1(n6825), .B2(n9470), .A(n6824), .ZN(n6826) );
  OAI21_X1 U8490 ( .B1(n6835), .B2(n9473), .A(n6826), .ZN(n9683) );
  NAND2_X1 U8491 ( .A1(n9683), .A2(n9269), .ZN(n6834) );
  INV_X1 U8492 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6827) );
  OAI22_X1 U8493 ( .A1(n9269), .A2(n6827), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9476), .ZN(n6831) );
  OAI21_X1 U8494 ( .B1(n6829), .B2(n9681), .A(n6828), .ZN(n9682) );
  NOR2_X1 U8495 ( .A1(n9239), .A2(n9682), .ZN(n6830) );
  AOI211_X1 U8496 ( .C1(n9264), .C2(n6832), .A(n6831), .B(n6830), .ZN(n6833)
         );
  OAI211_X1 U8497 ( .C1(n6835), .C2(n9245), .A(n6834), .B(n6833), .ZN(P1_U3288) );
  NAND2_X1 U8498 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7107) );
  INV_X1 U8499 ( .A(n7107), .ZN(n6843) );
  INV_X1 U8500 ( .A(n6836), .ZN(n6837) );
  AOI21_X1 U8501 ( .B1(n9851), .B2(n6838), .A(n6837), .ZN(n6840) );
  INV_X1 U8502 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6998) );
  AOI22_X1 U8503 ( .A1(n7096), .A2(n6998), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n6999), .ZN(n6839) );
  NOR2_X1 U8504 ( .A1(n6840), .A2(n6839), .ZN(n6997) );
  AOI21_X1 U8505 ( .B1(n6840), .B2(n6839), .A(n6997), .ZN(n6841) );
  NOR2_X1 U8506 ( .A1(n9741), .A2(n6841), .ZN(n6842) );
  AOI211_X1 U8507 ( .C1(n9739), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n6843), .B(
        n6842), .ZN(n6851) );
  INV_X1 U8508 ( .A(n6844), .ZN(n6845) );
  AOI21_X1 U8509 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7016), .A(n6845), .ZN(
        n6848) );
  INV_X1 U8510 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6846) );
  AOI22_X1 U8511 ( .A1(n7096), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n6846), .B2(
        n6999), .ZN(n6847) );
  NAND2_X1 U8512 ( .A1(n6848), .A2(n6847), .ZN(n7003) );
  OAI21_X1 U8513 ( .B1(n6848), .B2(n6847), .A(n7003), .ZN(n6849) );
  NAND2_X1 U8514 ( .A1(n9896), .A2(n6849), .ZN(n6850) );
  OAI211_X1 U8515 ( .C1(n9900), .C2(n6999), .A(n6851), .B(n6850), .ZN(P2_U3258) );
  AOI22_X1 U8516 ( .A1(n6852), .A2(n9816), .B1(n9815), .B2(n6955), .ZN(n6853)
         );
  OAI211_X1 U8517 ( .C1(n8644), .C2(n6855), .A(n6854), .B(n6853), .ZN(n6870)
         );
  NAND2_X1 U8518 ( .A1(n6870), .A2(n4405), .ZN(n6856) );
  OAI21_X1 U8519 ( .B1(n4405), .B2(n5999), .A(n6856), .ZN(P2_U3472) );
  INV_X1 U8520 ( .A(n7713), .ZN(n6858) );
  OAI222_X1 U8521 ( .A1(n7404), .A2(n6857), .B1(n8131), .B2(n6858), .C1(n8385), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U8522 ( .A1(n8929), .A2(P1_U3084), .B1(n9369), .B2(n6858), .C1(
        n10058), .C2(n9371), .ZN(P1_U3334) );
  INV_X1 U8523 ( .A(n7117), .ZN(n8279) );
  AOI22_X1 U8524 ( .A1(n8249), .A2(n4535), .B1(n8250), .B2(n8279), .ZN(n6860)
         );
  OAI211_X1 U8525 ( .C1(n6992), .C2(n8253), .A(n6860), .B(n6859), .ZN(n6868)
         );
  INV_X1 U8526 ( .A(n8255), .ZN(n8194) );
  NAND3_X1 U8527 ( .A1(n8194), .A2(n6861), .A3(n4535), .ZN(n6866) );
  OAI21_X1 U8528 ( .B1(n6863), .B2(n6862), .A(n8207), .ZN(n6865) );
  AOI21_X1 U8529 ( .B1(n6866), .B2(n6865), .A(n6864), .ZN(n6867) );
  AOI211_X1 U8530 ( .C1(n9814), .C2(n8259), .A(n6868), .B(n6867), .ZN(n6869)
         );
  INV_X1 U8531 ( .A(n6869), .ZN(P2_U3223) );
  NAND2_X1 U8532 ( .A1(n6870), .A2(n9853), .ZN(n6871) );
  OAI21_X1 U8533 ( .B1(n9853), .B2(n6872), .A(n6871), .ZN(P2_U3527) );
  NAND2_X1 U8534 ( .A1(n6874), .A2(n6873), .ZN(n6876) );
  XOR2_X1 U8535 ( .A(n6876), .B(n6875), .Z(n6880) );
  NAND2_X1 U8536 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3084), .ZN(n8879) );
  OAI21_X1 U8537 ( .B1(n8830), .B2(n7145), .A(n8879), .ZN(n6878) );
  OAI22_X1 U8538 ( .A1(n8831), .A2(n6946), .B1(n6943), .B2(n8816), .ZN(n6877)
         );
  AOI211_X1 U8539 ( .C1(n8819), .C2(n6952), .A(n6878), .B(n6877), .ZN(n6879)
         );
  OAI21_X1 U8540 ( .B1(n6880), .B2(n8825), .A(n6879), .ZN(P1_U3211) );
  NAND2_X1 U8541 ( .A1(n6881), .A2(n7787), .ZN(n6884) );
  AOI22_X1 U8542 ( .A1(n7703), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7714), .B2(
        n6882), .ZN(n6883) );
  INV_X1 U8543 ( .A(n7162), .ZN(n9824) );
  XNOR2_X1 U8544 ( .A(n7162), .B(n8114), .ZN(n6885) );
  NOR2_X1 U8545 ( .A1(n7161), .A2(n5905), .ZN(n6886) );
  NAND2_X1 U8546 ( .A1(n6885), .A2(n6886), .ZN(n6916) );
  INV_X1 U8547 ( .A(n6885), .ZN(n6915) );
  INV_X1 U8548 ( .A(n6886), .ZN(n6887) );
  NAND2_X1 U8549 ( .A1(n6915), .A2(n6887), .ZN(n6888) );
  AND2_X1 U8550 ( .A1(n6916), .A2(n6888), .ZN(n6895) );
  INV_X1 U8551 ( .A(n6889), .ZN(n6890) );
  NAND2_X1 U8552 ( .A1(n6891), .A2(n6890), .ZN(n6892) );
  OAI211_X1 U8553 ( .C1(n6895), .C2(n6894), .A(n6917), .B(n8207), .ZN(n6909)
         );
  INV_X1 U8554 ( .A(n7121), .ZN(n6907) );
  NAND2_X1 U8555 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n9886) );
  INV_X1 U8556 ( .A(n9886), .ZN(n6906) );
  NAND2_X1 U8557 ( .A1(n4401), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6904) );
  OR2_X1 U8558 ( .A1(n7802), .A2(n6896), .ZN(n6903) );
  INV_X1 U8559 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6897) );
  NAND2_X1 U8560 ( .A1(n6898), .A2(n6897), .ZN(n6899) );
  NAND2_X1 U8561 ( .A1(n6923), .A2(n6899), .ZN(n7197) );
  OR2_X1 U8562 ( .A1(n7768), .A2(n7197), .ZN(n6902) );
  OR2_X1 U8563 ( .A1(n7771), .A2(n6900), .ZN(n6901) );
  OAI22_X1 U8564 ( .A1(n7186), .A2(n8230), .B1(n8231), .B2(n7117), .ZN(n6905)
         );
  AOI211_X1 U8565 ( .C1(n6907), .C2(n8211), .A(n6906), .B(n6905), .ZN(n6908)
         );
  OAI211_X1 U8566 ( .C1(n9824), .C2(n8248), .A(n6909), .B(n6908), .ZN(P2_U3219) );
  NAND2_X1 U8567 ( .A1(n6910), .A2(n7787), .ZN(n6913) );
  AOI22_X1 U8568 ( .A1(n7703), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7714), .B2(
        n6911), .ZN(n6912) );
  XNOR2_X1 U8569 ( .A(n7196), .B(n5934), .ZN(n7023) );
  NOR2_X1 U8570 ( .A1(n7186), .A2(n5905), .ZN(n7024) );
  XNOR2_X1 U8571 ( .A(n7023), .B(n7024), .ZN(n6918) );
  INV_X1 U8572 ( .A(n6918), .ZN(n6914) );
  AOI21_X1 U8573 ( .B1(n6917), .B2(n6914), .A(n8263), .ZN(n6921) );
  NOR3_X1 U8574 ( .A1(n6915), .A2(n7161), .A3(n8255), .ZN(n6920) );
  NAND2_X1 U8575 ( .A1(n6919), .A2(n6918), .ZN(n7027) );
  OAI21_X1 U8576 ( .B1(n6921), .B2(n6920), .A(n7027), .ZN(n6934) );
  NAND2_X1 U8577 ( .A1(n4401), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6928) );
  OR2_X1 U8578 ( .A1(n7802), .A2(n9851), .ZN(n6927) );
  NAND2_X1 U8579 ( .A1(n6923), .A2(n6922), .ZN(n6924) );
  NAND2_X1 U8580 ( .A1(n7030), .A2(n6924), .ZN(n7189) );
  OR2_X1 U8581 ( .A1(n7768), .A2(n7189), .ZN(n6926) );
  OR2_X1 U8582 ( .A1(n7771), .A2(n7190), .ZN(n6925) );
  OR2_X1 U8583 ( .A1(n7293), .A2(n8550), .ZN(n6930) );
  OR2_X1 U8584 ( .A1(n7161), .A2(n8548), .ZN(n6929) );
  NAND2_X1 U8585 ( .A1(n6930), .A2(n6929), .ZN(n7166) );
  AOI22_X1 U8586 ( .A1(n8245), .A2(n7166), .B1(P2_REG3_REG_11__SCAN_IN), .B2(
        P2_U3152), .ZN(n6931) );
  OAI21_X1 U8587 ( .B1(n7197), .B2(n8253), .A(n6931), .ZN(n6932) );
  AOI21_X1 U8588 ( .B1(n7196), .B2(n8259), .A(n6932), .ZN(n6933) );
  NAND2_X1 U8589 ( .A1(n6934), .A2(n6933), .ZN(P2_U3238) );
  NAND2_X1 U8590 ( .A1(n6943), .A2(n9696), .ZN(n7634) );
  NAND3_X1 U8591 ( .A1(n7082), .A2(n7634), .A3(n7633), .ZN(n6936) );
  INV_X1 U8592 ( .A(n6943), .ZN(n8844) );
  NAND2_X1 U8593 ( .A1(n8844), .A2(n7081), .ZN(n7525) );
  NAND2_X1 U8594 ( .A1(n7525), .A2(n7447), .ZN(n6935) );
  NAND2_X1 U8595 ( .A1(n7634), .A2(n6935), .ZN(n7636) );
  NAND2_X1 U8596 ( .A1(n6936), .A2(n7636), .ZN(n6937) );
  NAND2_X1 U8597 ( .A1(n7049), .A2(n6952), .ZN(n7526) );
  NAND2_X1 U8598 ( .A1(n8843), .A2(n9706), .ZN(n7635) );
  NAND2_X1 U8599 ( .A1(n7526), .A2(n7635), .ZN(n7493) );
  NAND2_X1 U8600 ( .A1(n6937), .A2(n7493), .ZN(n6938) );
  NAND2_X1 U8601 ( .A1(n7044), .A2(n6938), .ZN(n6940) );
  OAI22_X1 U8602 ( .A1(n7145), .A2(n9467), .B1(n6943), .B2(n9465), .ZN(n6939)
         );
  AOI21_X1 U8603 ( .B1(n6940), .B2(n9470), .A(n6939), .ZN(n9704) );
  NAND2_X1 U8604 ( .A1(n8845), .A2(n9689), .ZN(n6941) );
  NAND2_X1 U8605 ( .A1(n6942), .A2(n6941), .ZN(n7076) );
  NAND2_X1 U8606 ( .A1(n6943), .A2(n7081), .ZN(n6944) );
  NAND2_X1 U8607 ( .A1(n6945), .A2(n7493), .ZN(n7051) );
  OAI21_X1 U8608 ( .B1(n6945), .B2(n7493), .A(n7051), .ZN(n9708) );
  NAND2_X1 U8609 ( .A1(n9708), .A2(n9214), .ZN(n6954) );
  OAI22_X1 U8610 ( .A1(n9269), .A2(n6947), .B1(n6946), .B2(n9476), .ZN(n6951)
         );
  NOR2_X1 U8611 ( .A1(n7078), .A2(n9696), .ZN(n7077) );
  NAND2_X1 U8612 ( .A1(n7077), .A2(n9706), .ZN(n7052) );
  OAI211_X1 U8613 ( .C1(n7077), .C2(n9706), .A(n7052), .B(n9711), .ZN(n9703)
         );
  NAND3_X1 U8614 ( .A1(n6949), .A2(n8929), .A3(n6948), .ZN(n9267) );
  NOR2_X1 U8615 ( .A1(n9703), .A2(n9267), .ZN(n6950) );
  AOI211_X1 U8616 ( .C1(n9264), .C2(n6952), .A(n6951), .B(n6950), .ZN(n6953)
         );
  OAI211_X1 U8617 ( .C1(n9223), .C2(n9704), .A(n6954), .B(n6953), .ZN(P1_U3284) );
  OAI22_X1 U8618 ( .A1(n6956), .A2(n7971), .B1(n6955), .B2(n4535), .ZN(n6975)
         );
  OR2_X1 U8619 ( .A1(n9814), .A2(n6963), .ZN(n7857) );
  OR2_X2 U8620 ( .A1(n6975), .A2(n7970), .ZN(n6977) );
  NAND2_X1 U8621 ( .A1(n9814), .A2(n8280), .ZN(n6957) );
  OR2_X1 U8622 ( .A1(n7112), .A2(n7117), .ZN(n7865) );
  NAND2_X1 U8623 ( .A1(n7112), .A2(n7117), .ZN(n7861) );
  INV_X1 U8624 ( .A(n6961), .ZN(n7973) );
  OAI21_X1 U8625 ( .B1(n6958), .B2(n7973), .A(n7114), .ZN(n7068) );
  INV_X1 U8626 ( .A(n7970), .ZN(n6979) );
  NAND3_X1 U8627 ( .A1(n6982), .A2(n7858), .A3(n7973), .ZN(n6962) );
  AOI21_X1 U8628 ( .B1(n7116), .B2(n6962), .A(n8529), .ZN(n6965) );
  OAI22_X1 U8629 ( .A1(n6963), .A2(n8548), .B1(n7161), .B2(n8550), .ZN(n6964)
         );
  AOI211_X1 U8630 ( .C1(n7068), .C2(n6978), .A(n6965), .B(n6964), .ZN(n7071)
         );
  INV_X1 U8631 ( .A(n9814), .ZN(n6993) );
  INV_X1 U8632 ( .A(n6991), .ZN(n6966) );
  INV_X1 U8633 ( .A(n7112), .ZN(n6967) );
  NAND2_X1 U8634 ( .A1(n6991), .A2(n6967), .ZN(n7123) );
  AOI21_X1 U8635 ( .B1(n7112), .B2(n6966), .A(n4623), .ZN(n7069) );
  NOR2_X1 U8636 ( .A1(n6967), .A2(n8538), .ZN(n6971) );
  OAI22_X1 U8637 ( .A1(n9768), .A2(n6969), .B1(n6968), .B2(n8556), .ZN(n6970)
         );
  AOI211_X1 U8638 ( .C1(n7069), .C2(n8521), .A(n6971), .B(n6970), .ZN(n6974)
         );
  NAND2_X1 U8639 ( .A1(n9768), .A2(n6972), .ZN(n8569) );
  INV_X1 U8640 ( .A(n8569), .ZN(n7305) );
  NAND2_X1 U8641 ( .A1(n7068), .A2(n7305), .ZN(n6973) );
  OAI211_X1 U8642 ( .C1(n7071), .C2(n8518), .A(n6974), .B(n6973), .ZN(P2_U3287) );
  NAND2_X1 U8643 ( .A1(n6975), .A2(n7970), .ZN(n6976) );
  NAND2_X1 U8644 ( .A1(n6977), .A2(n6976), .ZN(n9820) );
  INV_X1 U8645 ( .A(n6978), .ZN(n9797) );
  OR2_X1 U8646 ( .A1(n9820), .A2(n9797), .ZN(n6987) );
  NAND2_X1 U8647 ( .A1(n6980), .A2(n6979), .ZN(n6981) );
  NAND2_X1 U8648 ( .A1(n6982), .A2(n6981), .ZN(n6985) );
  OAI22_X1 U8649 ( .A1(n6983), .A2(n8548), .B1(n7117), .B2(n8550), .ZN(n6984)
         );
  AOI21_X1 U8650 ( .B1(n6985), .B2(n9748), .A(n6984), .ZN(n6986) );
  NAND2_X1 U8651 ( .A1(n6987), .A2(n6986), .ZN(n9822) );
  MUX2_X1 U8652 ( .A(n9822), .B(P2_REG2_REG_8__SCAN_IN), .S(n8535), .Z(n6988)
         );
  INV_X1 U8653 ( .A(n6988), .ZN(n6996) );
  NOR2_X1 U8654 ( .A1(n6989), .A2(n6993), .ZN(n6990) );
  NOR2_X1 U8655 ( .A1(n6991), .A2(n6990), .ZN(n9817) );
  OAI22_X1 U8656 ( .A1(n8538), .A2(n6993), .B1(n8556), .B2(n6992), .ZN(n6994)
         );
  AOI21_X1 U8657 ( .B1(n9817), .B2(n8521), .A(n6994), .ZN(n6995) );
  OAI211_X1 U8658 ( .C1(n9820), .C2(n8569), .A(n6996), .B(n6995), .ZN(P2_U3288) );
  AOI21_X1 U8659 ( .B1(n6999), .B2(n6998), .A(n6997), .ZN(n7001) );
  INV_X1 U8660 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9452) );
  AOI22_X1 U8661 ( .A1(n7209), .A2(n9452), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7135), .ZN(n7000) );
  NOR2_X1 U8662 ( .A1(n7001), .A2(n7000), .ZN(n7134) );
  AOI21_X1 U8663 ( .B1(n7001), .B2(n7000), .A(n7134), .ZN(n7011) );
  NOR2_X1 U8664 ( .A1(n7209), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7002) );
  AOI21_X1 U8665 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n7209), .A(n7002), .ZN(
        n7005) );
  OAI21_X1 U8666 ( .B1(n7005), .B2(n7004), .A(n7132), .ZN(n7009) );
  INV_X1 U8667 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7007) );
  NAND2_X1 U8668 ( .A1(n9395), .A2(n7209), .ZN(n7006) );
  NAND2_X1 U8669 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7225) );
  OAI211_X1 U8670 ( .C1(n7007), .C2(n9888), .A(n7006), .B(n7225), .ZN(n7008)
         );
  AOI21_X1 U8671 ( .B1(n7009), .B2(n9896), .A(n7008), .ZN(n7010) );
  OAI21_X1 U8672 ( .B1(n7011), .B2(n9741), .A(n7010), .ZN(P2_U3259) );
  INV_X1 U8673 ( .A(n7721), .ZN(n7014) );
  OAI222_X1 U8674 ( .A1(P1_U3084), .A2(n7013), .B1(n9369), .B2(n7014), .C1(
        n7012), .C2(n9371), .ZN(P1_U3333) );
  OAI222_X1 U8675 ( .A1(n7404), .A2(n10070), .B1(P2_U3152), .B2(n7992), .C1(
        n8131), .C2(n7014), .ZN(P2_U3338) );
  NAND2_X1 U8676 ( .A1(n7015), .A2(n7787), .ZN(n7018) );
  AOI22_X1 U8677 ( .A1(n7703), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7714), .B2(
        n7016), .ZN(n7017) );
  XNOR2_X1 U8678 ( .A(n7285), .B(n5934), .ZN(n7019) );
  OR2_X1 U8679 ( .A1(n7293), .A2(n5905), .ZN(n7020) );
  NAND2_X1 U8680 ( .A1(n7019), .A2(n7020), .ZN(n7091) );
  INV_X1 U8681 ( .A(n7019), .ZN(n7022) );
  INV_X1 U8682 ( .A(n7020), .ZN(n7021) );
  NAND2_X1 U8683 ( .A1(n7022), .A2(n7021), .ZN(n7093) );
  NAND2_X1 U8684 ( .A1(n7091), .A2(n7093), .ZN(n7028) );
  INV_X1 U8685 ( .A(n7023), .ZN(n7025) );
  NAND2_X1 U8686 ( .A1(n7025), .A2(n7024), .ZN(n7026) );
  XOR2_X1 U8687 ( .A(n7028), .B(n7092), .Z(n7041) );
  INV_X1 U8688 ( .A(n7186), .ZN(n8277) );
  NAND2_X1 U8689 ( .A1(n4401), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7036) );
  OR2_X1 U8690 ( .A1(n7802), .A2(n6998), .ZN(n7035) );
  NAND2_X1 U8691 ( .A1(n7030), .A2(n7029), .ZN(n7031) );
  NAND2_X1 U8692 ( .A1(n7100), .A2(n7031), .ZN(n7301) );
  OR2_X1 U8693 ( .A1(n7768), .A2(n7301), .ZN(n7034) );
  OR2_X1 U8694 ( .A1(n7032), .A2(n6846), .ZN(n7033) );
  INV_X1 U8695 ( .A(n7326), .ZN(n8275) );
  AOI22_X1 U8696 ( .A1(n8249), .A2(n8277), .B1(n8250), .B2(n8275), .ZN(n7038)
         );
  OAI211_X1 U8697 ( .C1(n7189), .C2(n8253), .A(n7038), .B(n7037), .ZN(n7039)
         );
  AOI21_X1 U8698 ( .B1(n7285), .B2(n8259), .A(n7039), .ZN(n7040) );
  OAI21_X1 U8699 ( .B1(n7041), .B2(n8263), .A(n7040), .ZN(P2_U3226) );
  INV_X1 U8700 ( .A(n7730), .ZN(n7066) );
  OAI222_X1 U8701 ( .A1(P1_U3084), .A2(n7612), .B1(n9371), .B2(n5611), .C1(
        n7066), .C2(n9369), .ZN(P1_U3332) );
  NAND2_X1 U8702 ( .A1(n7145), .A2(n4403), .ZN(n7537) );
  INV_X1 U8703 ( .A(n7145), .ZN(n8842) );
  NAND2_X1 U8704 ( .A1(n8842), .A2(n7053), .ZN(n7539) );
  INV_X1 U8705 ( .A(n7149), .ZN(n7497) );
  INV_X1 U8706 ( .A(n7526), .ZN(n7042) );
  NOR2_X1 U8707 ( .A1(n7497), .A2(n7042), .ZN(n7043) );
  INV_X1 U8708 ( .A(n7143), .ZN(n7046) );
  AOI21_X1 U8709 ( .B1(n7044), .B2(n7526), .A(n7149), .ZN(n7045) );
  NOR3_X1 U8710 ( .A1(n7046), .A2(n7045), .A3(n9234), .ZN(n7048) );
  INV_X1 U8711 ( .A(n8841), .ZN(n7237) );
  OAI22_X1 U8712 ( .A1(n7237), .A2(n9467), .B1(n7049), .B2(n9465), .ZN(n7047)
         );
  NOR2_X1 U8713 ( .A1(n7048), .A2(n7047), .ZN(n9714) );
  NAND2_X1 U8714 ( .A1(n7049), .A2(n9706), .ZN(n7050) );
  XNOR2_X1 U8715 ( .A(n7148), .B(n7149), .ZN(n9716) );
  INV_X1 U8716 ( .A(n9716), .ZN(n9718) );
  NAND2_X1 U8717 ( .A1(n9718), .A2(n9214), .ZN(n7057) );
  OR2_X1 U8718 ( .A1(n7052), .A2(n4403), .ZN(n7153) );
  INV_X1 U8719 ( .A(n7153), .ZN(n7155) );
  AOI21_X1 U8720 ( .B1(n4403), .B2(n7052), .A(n7155), .ZN(n9712) );
  NOR2_X1 U8721 ( .A1(n9475), .A2(n7053), .ZN(n7055) );
  OAI22_X1 U8722 ( .A1(n9269), .A2(n6291), .B1(n8716), .B2(n9476), .ZN(n7054)
         );
  AOI211_X1 U8723 ( .C1(n9712), .C2(n9461), .A(n7055), .B(n7054), .ZN(n7056)
         );
  OAI211_X1 U8724 ( .C1(n9223), .C2(n9714), .A(n7057), .B(n7056), .ZN(P1_U3283) );
  XOR2_X1 U8725 ( .A(n7059), .B(n7058), .Z(n7065) );
  NAND2_X1 U8726 ( .A1(n7233), .A2(n9709), .ZN(n9720) );
  INV_X1 U8727 ( .A(n9720), .ZN(n7062) );
  NAND2_X1 U8728 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3084), .ZN(n9609) );
  OAI21_X1 U8729 ( .B1(n8830), .B2(n9466), .A(n9609), .ZN(n7061) );
  OAI22_X1 U8730 ( .A1(n8831), .A2(n7151), .B1(n7145), .B2(n8816), .ZN(n7060)
         );
  AOI211_X1 U8731 ( .C1(n7063), .C2(n7062), .A(n7061), .B(n7060), .ZN(n7064)
         );
  OAI21_X1 U8732 ( .B1(n7065), .B2(n8825), .A(n7064), .ZN(P1_U3229) );
  OAI222_X1 U8733 ( .A1(n7404), .A2(n7067), .B1(P2_U3152), .B2(n7994), .C1(
        n8131), .C2(n7066), .ZN(P2_U3337) );
  INV_X1 U8734 ( .A(n7068), .ZN(n7072) );
  INV_X1 U8735 ( .A(n9829), .ZN(n9819) );
  AOI22_X1 U8736 ( .A1(n7069), .A2(n9816), .B1(n9815), .B2(n7112), .ZN(n7070)
         );
  OAI211_X1 U8737 ( .C1(n7072), .C2(n9819), .A(n7071), .B(n7070), .ZN(n7074)
         );
  NAND2_X1 U8738 ( .A1(n7074), .A2(n9853), .ZN(n7073) );
  OAI21_X1 U8739 ( .B1(n9853), .B2(n6785), .A(n7073), .ZN(P2_U3529) );
  INV_X1 U8740 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10055) );
  NAND2_X1 U8741 ( .A1(n7074), .A2(n4405), .ZN(n7075) );
  OAI21_X1 U8742 ( .B1(n4405), .B2(n10055), .A(n7075), .ZN(P2_U3478) );
  XOR2_X1 U8743 ( .A(n7076), .B(n7085), .Z(n9700) );
  AOI21_X1 U8744 ( .B1(n9696), .B2(n7078), .A(n7077), .ZN(n9697) );
  INV_X1 U8745 ( .A(n7079), .ZN(n8805) );
  INV_X1 U8746 ( .A(n9476), .ZN(n9172) );
  AOI22_X1 U8747 ( .A1(n9223), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n8805), .B2(
        n9172), .ZN(n7080) );
  OAI21_X1 U8748 ( .B1(n7081), .B2(n9475), .A(n7080), .ZN(n7089) );
  NAND2_X1 U8749 ( .A1(n7082), .A2(n7633), .ZN(n7083) );
  NAND2_X1 U8750 ( .A1(n7528), .A2(n7085), .ZN(n7084) );
  OAI211_X1 U8751 ( .C1(n7528), .C2(n7085), .A(n7084), .B(n9470), .ZN(n7087)
         );
  AOI22_X1 U8752 ( .A1(n9253), .A2(n8845), .B1(n8843), .B2(n9254), .ZN(n7086)
         );
  AND2_X1 U8753 ( .A1(n7087), .A2(n7086), .ZN(n9699) );
  NOR2_X1 U8754 ( .A1(n9699), .A2(n9223), .ZN(n7088) );
  AOI211_X1 U8755 ( .C1(n9697), .C2(n9461), .A(n7089), .B(n7088), .ZN(n7090)
         );
  OAI21_X1 U8756 ( .B1(n9271), .B2(n9700), .A(n7090), .ZN(P1_U3285) );
  NAND2_X1 U8757 ( .A1(n7092), .A2(n7091), .ZN(n7094) );
  NAND2_X1 U8758 ( .A1(n7095), .A2(n7787), .ZN(n7098) );
  AOI22_X1 U8759 ( .A1(n7703), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7714), .B2(
        n7096), .ZN(n7097) );
  XNOR2_X1 U8760 ( .A(n7337), .B(n5934), .ZN(n7219) );
  NOR2_X1 U8761 ( .A1(n7326), .A2(n5905), .ZN(n7220) );
  XNOR2_X1 U8762 ( .A(n7219), .B(n7220), .ZN(n7217) );
  XNOR2_X1 U8763 ( .A(n7218), .B(n7217), .ZN(n7111) );
  INV_X1 U8764 ( .A(n7293), .ZN(n8276) );
  NAND2_X1 U8765 ( .A1(n4401), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7106) );
  OR2_X1 U8766 ( .A1(n7802), .A2(n9452), .ZN(n7105) );
  INV_X1 U8767 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7099) );
  NAND2_X1 U8768 ( .A1(n7100), .A2(n7099), .ZN(n7101) );
  NAND2_X1 U8769 ( .A1(n7102), .A2(n7101), .ZN(n7330) );
  OR2_X1 U8770 ( .A1(n7746), .A2(n7330), .ZN(n7104) );
  INV_X1 U8771 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7331) );
  OR2_X1 U8772 ( .A1(n7771), .A2(n7331), .ZN(n7103) );
  INV_X1 U8773 ( .A(n7377), .ZN(n8274) );
  AOI22_X1 U8774 ( .A1(n8249), .A2(n8276), .B1(n8250), .B2(n8274), .ZN(n7108)
         );
  OAI211_X1 U8775 ( .C1(n8253), .C2(n7301), .A(n7108), .B(n7107), .ZN(n7109)
         );
  AOI21_X1 U8776 ( .B1(n7337), .B2(n8259), .A(n7109), .ZN(n7110) );
  OAI21_X1 U8777 ( .B1(n7111), .B2(n8263), .A(n7110), .ZN(P2_U3236) );
  OR2_X1 U8778 ( .A1(n7112), .A2(n8279), .ZN(n7113) );
  NAND2_X1 U8779 ( .A1(n7162), .A2(n7161), .ZN(n7862) );
  NAND2_X1 U8780 ( .A1(n7864), .A2(n7862), .ZN(n7974) );
  OAI21_X1 U8781 ( .B1(n7115), .B2(n7974), .A(n7164), .ZN(n9823) );
  XOR2_X1 U8782 ( .A(n7974), .B(n7165), .Z(n7119) );
  OAI22_X1 U8783 ( .A1(n7186), .A2(n8550), .B1(n7117), .B2(n8548), .ZN(n7118)
         );
  AOI21_X1 U8784 ( .B1(n7119), .B2(n9748), .A(n7118), .ZN(n7120) );
  OAI21_X1 U8785 ( .B1(n9823), .B2(n9797), .A(n7120), .ZN(n9826) );
  NAND2_X1 U8786 ( .A1(n9826), .A2(n8555), .ZN(n7128) );
  OAI22_X1 U8787 ( .A1(n8555), .A2(n7122), .B1(n7121), .B2(n8556), .ZN(n7126)
         );
  NAND2_X1 U8788 ( .A1(n7123), .A2(n7162), .ZN(n7124) );
  NAND2_X1 U8789 ( .A1(n4487), .A2(n7124), .ZN(n9825) );
  NOR2_X1 U8790 ( .A1(n9825), .A2(n8562), .ZN(n7125) );
  AOI211_X1 U8791 ( .C1(n8566), .C2(n7162), .A(n7126), .B(n7125), .ZN(n7127)
         );
  OAI211_X1 U8792 ( .C1(n9823), .C2(n8569), .A(n7128), .B(n7127), .ZN(P2_U3286) );
  INV_X1 U8793 ( .A(n7733), .ZN(n7130) );
  OAI222_X1 U8794 ( .A1(P1_U3084), .A2(n5170), .B1(n9369), .B2(n7130), .C1(
        n7129), .C2(n9371), .ZN(P1_U3331) );
  OAI222_X1 U8795 ( .A1(n7404), .A2(n7131), .B1(n8131), .B2(n7130), .C1(n7819), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  NAND2_X1 U8796 ( .A1(n7133), .A2(n7381), .ZN(n7315) );
  OAI21_X1 U8797 ( .B1(n7133), .B2(n7381), .A(n7315), .ZN(n7141) );
  AOI21_X1 U8798 ( .B1(n7135), .B2(n9452), .A(n7134), .ZN(n7308) );
  XNOR2_X1 U8799 ( .A(n7308), .B(n7314), .ZN(n7136) );
  NAND2_X1 U8800 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7136), .ZN(n7309) );
  OAI211_X1 U8801 ( .C1(n7136), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9891), .B(
        n7309), .ZN(n7139) );
  NAND2_X1 U8802 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n8251) );
  INV_X1 U8803 ( .A(n8251), .ZN(n7137) );
  AOI21_X1 U8804 ( .B1(n9739), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7137), .ZN(
        n7138) );
  OAI211_X1 U8805 ( .C1(n9900), .C2(n7314), .A(n7139), .B(n7138), .ZN(n7140)
         );
  AOI21_X1 U8806 ( .B1(n9896), .B2(n7141), .A(n7140), .ZN(n7142) );
  INV_X1 U8807 ( .A(n7142), .ZN(P2_U3260) );
  NAND2_X1 U8808 ( .A1(n7237), .A2(n7233), .ZN(n7529) );
  INV_X1 U8809 ( .A(n7233), .ZN(n7156) );
  NAND2_X1 U8810 ( .A1(n7156), .A2(n8841), .ZN(n7538) );
  NAND2_X1 U8811 ( .A1(n7529), .A2(n7538), .ZN(n7498) );
  INV_X1 U8812 ( .A(n7498), .ZN(n7144) );
  XNOR2_X1 U8813 ( .A(n7235), .B(n7144), .ZN(n7147) );
  OAI22_X1 U8814 ( .A1(n7145), .A2(n9465), .B1(n9466), .B2(n9467), .ZN(n7146)
         );
  AOI21_X1 U8815 ( .B1(n7147), .B2(n9470), .A(n7146), .ZN(n9721) );
  NAND2_X1 U8816 ( .A1(n8842), .A2(n4403), .ZN(n7150) );
  XOR2_X1 U8817 ( .A(n7498), .B(n7234), .Z(n9726) );
  NAND2_X1 U8818 ( .A1(n9726), .A2(n9214), .ZN(n7160) );
  INV_X1 U8819 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7152) );
  OAI22_X1 U8820 ( .A1(n9269), .A2(n7152), .B1(n7151), .B2(n9476), .ZN(n7158)
         );
  INV_X1 U8821 ( .A(n7243), .ZN(n7154) );
  OAI21_X1 U8822 ( .B1(n7156), .B2(n7155), .A(n7154), .ZN(n9722) );
  NOR2_X1 U8823 ( .A1(n9722), .A2(n9239), .ZN(n7157) );
  AOI211_X1 U8824 ( .C1(n9264), .C2(n7233), .A(n7158), .B(n7157), .ZN(n7159)
         );
  OAI211_X1 U8825 ( .C1(n9223), .C2(n9721), .A(n7160), .B(n7159), .ZN(P1_U3282) );
  INV_X1 U8826 ( .A(n7161), .ZN(n8278) );
  NAND2_X1 U8827 ( .A1(n7162), .A2(n8278), .ZN(n7163) );
  NAND2_X1 U8828 ( .A1(n7164), .A2(n7163), .ZN(n7180) );
  NAND2_X1 U8829 ( .A1(n7196), .A2(n7186), .ZN(n7874) );
  XNOR2_X1 U8830 ( .A(n7180), .B(n7976), .ZN(n7207) );
  XNOR2_X1 U8831 ( .A(n7183), .B(n7976), .ZN(n7167) );
  AOI21_X1 U8832 ( .B1(n7167), .B2(n9748), .A(n7166), .ZN(n7201) );
  AOI211_X1 U8833 ( .C1(n7196), .C2(n4487), .A(n9833), .B(n7188), .ZN(n7205)
         );
  AOI21_X1 U8834 ( .B1(n9815), .B2(n7196), .A(n7205), .ZN(n7168) );
  OAI211_X1 U8835 ( .C1(n7207), .C2(n8644), .A(n7201), .B(n7168), .ZN(n7170)
         );
  NAND2_X1 U8836 ( .A1(n7170), .A2(n9853), .ZN(n7169) );
  OAI21_X1 U8837 ( .B1(n9853), .B2(n6896), .A(n7169), .ZN(P2_U3531) );
  INV_X1 U8838 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7172) );
  NAND2_X1 U8839 ( .A1(n7170), .A2(n4405), .ZN(n7171) );
  OAI21_X1 U8840 ( .B1(n4405), .B2(n7172), .A(n7171), .ZN(P2_U3484) );
  INV_X1 U8841 ( .A(n7740), .ZN(n7175) );
  AOI21_X1 U8842 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n7173), .A(n8002), .ZN(
        n7174) );
  OAI21_X1 U8843 ( .B1(n7175), .B2(n8131), .A(n7174), .ZN(P2_U3335) );
  NAND2_X1 U8844 ( .A1(n7740), .A2(n7176), .ZN(n7178) );
  NAND2_X1 U8845 ( .A1(n7177), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7671) );
  OAI211_X1 U8846 ( .C1(n7179), .C2(n9371), .A(n7178), .B(n7671), .ZN(P1_U3330) );
  NAND2_X1 U8847 ( .A1(n7180), .A2(n7976), .ZN(n7182) );
  NAND2_X1 U8848 ( .A1(n7196), .A2(n8277), .ZN(n7181) );
  NAND2_X1 U8849 ( .A1(n7182), .A2(n7181), .ZN(n7286) );
  OR2_X1 U8850 ( .A1(n7285), .A2(n7293), .ZN(n7876) );
  NAND2_X1 U8851 ( .A1(n7285), .A2(n7293), .ZN(n7875) );
  XNOR2_X1 U8852 ( .A(n7286), .B(n7978), .ZN(n9838) );
  INV_X1 U8853 ( .A(n9838), .ZN(n7195) );
  NAND2_X1 U8854 ( .A1(n7183), .A2(n7874), .ZN(n7289) );
  NAND2_X1 U8855 ( .A1(n7289), .A2(n7863), .ZN(n7184) );
  XNOR2_X1 U8856 ( .A(n7184), .B(n7978), .ZN(n7185) );
  OAI222_X1 U8857 ( .A1(n8550), .A2(n7326), .B1(n8548), .B2(n7186), .C1(n8529), 
        .C2(n7185), .ZN(n9835) );
  INV_X1 U8858 ( .A(n7285), .ZN(n9832) );
  INV_X1 U8859 ( .A(n7299), .ZN(n7187) );
  OAI21_X1 U8860 ( .B1(n9832), .B2(n7188), .A(n7187), .ZN(n9834) );
  OAI22_X1 U8861 ( .A1(n9768), .A2(n7190), .B1(n7189), .B2(n8556), .ZN(n7191)
         );
  AOI21_X1 U8862 ( .B1(n7285), .B2(n8566), .A(n7191), .ZN(n7192) );
  OAI21_X1 U8863 ( .B1(n9834), .B2(n8562), .A(n7192), .ZN(n7193) );
  AOI21_X1 U8864 ( .B1(n9835), .B2(n9768), .A(n7193), .ZN(n7194) );
  OAI21_X1 U8865 ( .B1(n8541), .B2(n7195), .A(n7194), .ZN(P2_U3284) );
  INV_X1 U8866 ( .A(n7196), .ZN(n7200) );
  INV_X1 U8867 ( .A(n7197), .ZN(n7198) );
  AOI22_X1 U8868 ( .A1(n8535), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7198), .B2(
        n9756), .ZN(n7199) );
  OAI21_X1 U8869 ( .B1(n7200), .B2(n8538), .A(n7199), .ZN(n7203) );
  NOR2_X1 U8870 ( .A1(n7201), .A2(n8535), .ZN(n7202) );
  AOI211_X1 U8871 ( .C1(n7205), .C2(n7204), .A(n7203), .B(n7202), .ZN(n7206)
         );
  OAI21_X1 U8872 ( .B1(n8541), .B2(n7207), .A(n7206), .ZN(P2_U3285) );
  NAND2_X1 U8873 ( .A1(n7208), .A2(n7787), .ZN(n7211) );
  AOI22_X1 U8874 ( .A1(n7703), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7714), .B2(
        n7209), .ZN(n7210) );
  XNOR2_X1 U8875 ( .A(n7365), .B(n5934), .ZN(n7212) );
  OR2_X1 U8876 ( .A1(n7377), .A2(n5905), .ZN(n7213) );
  NAND2_X1 U8877 ( .A1(n7212), .A2(n7213), .ZN(n8048) );
  INV_X1 U8878 ( .A(n7212), .ZN(n7215) );
  INV_X1 U8879 ( .A(n7213), .ZN(n7214) );
  NAND2_X1 U8880 ( .A1(n7215), .A2(n7214), .ZN(n7216) );
  NAND2_X1 U8881 ( .A1(n8048), .A2(n7216), .ZN(n7224) );
  INV_X1 U8882 ( .A(n7219), .ZN(n7221) );
  NAND2_X1 U8883 ( .A1(n7221), .A2(n7220), .ZN(n7222) );
  AOI21_X1 U8884 ( .B1(n7224), .B2(n7223), .A(n4488), .ZN(n7229) );
  OAI21_X1 U8885 ( .B1(n8253), .B2(n7330), .A(n7225), .ZN(n7227) );
  OAI22_X1 U8886 ( .A1(n7326), .A2(n8231), .B1(n8230), .B2(n8549), .ZN(n7226)
         );
  AOI211_X1 U8887 ( .C1(n7365), .C2(n8259), .A(n7227), .B(n7226), .ZN(n7228)
         );
  OAI21_X1 U8888 ( .B1(n7229), .B2(n8263), .A(n7228), .ZN(P2_U3217) );
  INV_X1 U8889 ( .A(n7752), .ZN(n7231) );
  INV_X1 U8890 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n10057) );
  OAI222_X1 U8891 ( .A1(P2_U3152), .A2(n7230), .B1(n8131), .B2(n7231), .C1(
        n10057), .C2(n7404), .ZN(P2_U3334) );
  OAI222_X1 U8892 ( .A1(n7232), .A2(P1_U3084), .B1(n9369), .B2(n7231), .C1(
        n10071), .C2(n9371), .ZN(P1_U3329) );
  NAND2_X1 U8893 ( .A1(n8700), .A2(n9466), .ZN(n7532) );
  NAND2_X1 U8894 ( .A1(n7457), .A2(n7532), .ZN(n7266) );
  INV_X1 U8895 ( .A(n7266), .ZN(n7500) );
  XNOR2_X1 U8896 ( .A(n7267), .B(n7500), .ZN(n9402) );
  NAND2_X1 U8897 ( .A1(n7278), .A2(n7529), .ZN(n7236) );
  XNOR2_X1 U8898 ( .A(n7236), .B(n7500), .ZN(n7239) );
  INV_X1 U8899 ( .A(n8839), .ZN(n7282) );
  OAI22_X1 U8900 ( .A1(n7282), .A2(n9467), .B1(n7237), .B2(n9465), .ZN(n7238)
         );
  AOI21_X1 U8901 ( .B1(n7239), .B2(n9470), .A(n7238), .ZN(n7240) );
  OAI21_X1 U8902 ( .B1(n9402), .B2(n9473), .A(n7240), .ZN(n9405) );
  NAND2_X1 U8903 ( .A1(n9405), .A2(n9269), .ZN(n7247) );
  OAI22_X1 U8904 ( .A1(n9479), .A2(n7241), .B1(n8698), .B2(n9476), .ZN(n7245)
         );
  INV_X1 U8905 ( .A(n8700), .ZN(n9404) );
  INV_X1 U8906 ( .A(n9458), .ZN(n7242) );
  OAI211_X1 U8907 ( .C1(n9404), .C2(n7243), .A(n7242), .B(n9711), .ZN(n9403)
         );
  NOR2_X1 U8908 ( .A1(n9403), .A2(n9267), .ZN(n7244) );
  AOI211_X1 U8909 ( .C1(n9264), .C2(n8700), .A(n7245), .B(n7244), .ZN(n7246)
         );
  OAI211_X1 U8910 ( .C1(n9402), .C2(n9245), .A(n7247), .B(n7246), .ZN(P1_U3281) );
  INV_X1 U8911 ( .A(n7248), .ZN(n7250) );
  NAND2_X1 U8912 ( .A1(n7250), .A2(n7249), .ZN(n7251) );
  XNOR2_X1 U8913 ( .A(n7252), .B(n7251), .ZN(n7257) );
  INV_X1 U8914 ( .A(n9229), .ZN(n7454) );
  OAI21_X1 U8915 ( .B1(n8830), .B2(n7454), .A(n7253), .ZN(n7255) );
  OAI22_X1 U8916 ( .A1(n8831), .A2(n7357), .B1(n9468), .B2(n8816), .ZN(n7254)
         );
  AOI211_X1 U8917 ( .C1(n9499), .C2(n8819), .A(n7255), .B(n7254), .ZN(n7256)
         );
  OAI21_X1 U8918 ( .B1(n7257), .B2(n8825), .A(n7256), .ZN(P1_U3232) );
  INV_X1 U8919 ( .A(n7258), .ZN(n7259) );
  AOI21_X1 U8920 ( .B1(n7261), .B2(n7260), .A(n7259), .ZN(n7265) );
  AND2_X1 U8921 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9623) );
  INV_X1 U8922 ( .A(n9252), .ZN(n7455) );
  OAI22_X1 U8923 ( .A1(n8831), .A2(n7273), .B1(n7455), .B2(n8830), .ZN(n7262)
         );
  AOI211_X1 U8924 ( .C1(n8833), .C2(n8839), .A(n9623), .B(n7262), .ZN(n7264)
         );
  NAND2_X1 U8925 ( .A1(n9508), .A2(n8819), .ZN(n7263) );
  OAI211_X1 U8926 ( .C1(n7265), .C2(n8825), .A(n7264), .B(n7263), .ZN(P1_U3222) );
  NAND2_X1 U8927 ( .A1(n7267), .A2(n7266), .ZN(n7269) );
  INV_X1 U8928 ( .A(n9466), .ZN(n8840) );
  OR2_X1 U8929 ( .A1(n8840), .A2(n8700), .ZN(n7268) );
  NOR2_X1 U8930 ( .A1(n8783), .A2(n8839), .ZN(n7271) );
  NAND2_X1 U8931 ( .A1(n8783), .A2(n8839), .ZN(n7270) );
  OR2_X1 U8932 ( .A1(n9508), .A2(n9468), .ZN(n7554) );
  NAND2_X1 U8933 ( .A1(n9508), .A2(n9468), .ZN(n7533) );
  NAND2_X1 U8934 ( .A1(n7554), .A2(n7533), .ZN(n7347) );
  XNOR2_X1 U8935 ( .A(n7348), .B(n7347), .ZN(n9510) );
  INV_X1 U8936 ( .A(n8783), .ZN(n9513) );
  AOI211_X1 U8937 ( .C1(n9508), .C2(n4433), .A(n9723), .B(n4641), .ZN(n9507)
         );
  INV_X1 U8938 ( .A(n9267), .ZN(n7277) );
  INV_X1 U8939 ( .A(n9508), .ZN(n7272) );
  NOR2_X1 U8940 ( .A1(n7272), .A2(n9475), .ZN(n7276) );
  INV_X1 U8941 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7274) );
  OAI22_X1 U8942 ( .A1(n9479), .A2(n7274), .B1(n7273), .B2(n9476), .ZN(n7275)
         );
  AOI211_X1 U8943 ( .C1(n9507), .C2(n7277), .A(n7276), .B(n7275), .ZN(n7284)
         );
  AND2_X1 U8944 ( .A1(n7532), .A2(n7529), .ZN(n7543) );
  NAND2_X1 U8945 ( .A1(n8783), .A2(n7282), .ZN(n7441) );
  NAND2_X1 U8946 ( .A1(n9463), .A2(n7441), .ZN(n7350) );
  OR2_X1 U8947 ( .A1(n8783), .A2(n7282), .ZN(n7349) );
  NAND2_X1 U8948 ( .A1(n7350), .A2(n7349), .ZN(n7280) );
  INV_X1 U8949 ( .A(n7347), .ZN(n7501) );
  XNOR2_X1 U8950 ( .A(n7280), .B(n7501), .ZN(n7281) );
  OAI222_X1 U8951 ( .A1(n9467), .A2(n7455), .B1(n9465), .B2(n7282), .C1(n9234), 
        .C2(n7281), .ZN(n9506) );
  NAND2_X1 U8952 ( .A1(n9506), .A2(n9269), .ZN(n7283) );
  OAI211_X1 U8953 ( .C1(n9510), .C2(n9271), .A(n7284), .B(n7283), .ZN(P1_U3279) );
  OR2_X1 U8954 ( .A1(n7337), .A2(n7326), .ZN(n7881) );
  NAND2_X1 U8955 ( .A1(n7337), .A2(n7326), .ZN(n7324) );
  OR2_X2 U8956 ( .A1(n7287), .A2(n7979), .ZN(n7339) );
  NAND2_X1 U8957 ( .A1(n7287), .A2(n7979), .ZN(n7288) );
  NAND2_X1 U8958 ( .A1(n7339), .A2(n7288), .ZN(n7298) );
  OR2_X1 U8959 ( .A1(n7298), .A2(n9797), .ZN(n7297) );
  AND2_X1 U8960 ( .A1(n7876), .A2(n7863), .ZN(n7872) );
  NOR2_X1 U8961 ( .A1(n7291), .A2(n7979), .ZN(n7292) );
  OR2_X1 U8962 ( .A1(n7325), .A2(n7292), .ZN(n7295) );
  OAI22_X1 U8963 ( .A1(n7293), .A2(n8548), .B1(n7377), .B2(n8550), .ZN(n7294)
         );
  AOI21_X1 U8964 ( .B1(n7295), .B2(n9748), .A(n7294), .ZN(n7296) );
  AND2_X1 U8965 ( .A1(n7297), .A2(n7296), .ZN(n8656) );
  INV_X1 U8966 ( .A(n7298), .ZN(n8654) );
  INV_X1 U8967 ( .A(n7337), .ZN(n8651) );
  OR2_X1 U8968 ( .A1(n7299), .A2(n8651), .ZN(n7300) );
  NAND2_X1 U8969 ( .A1(n7332), .A2(n7300), .ZN(n8652) );
  OAI22_X1 U8970 ( .A1(n9768), .A2(n6846), .B1(n7301), .B2(n8556), .ZN(n7302)
         );
  AOI21_X1 U8971 ( .B1(n7337), .B2(n8566), .A(n7302), .ZN(n7303) );
  OAI21_X1 U8972 ( .B1(n8652), .B2(n8562), .A(n7303), .ZN(n7304) );
  AOI21_X1 U8973 ( .B1(n8654), .B2(n7305), .A(n7304), .ZN(n7306) );
  OAI21_X1 U8974 ( .B1(n8656), .B2(n8518), .A(n7306), .ZN(P2_U3283) );
  INV_X1 U8975 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n10074) );
  NOR2_X1 U8976 ( .A1(n8291), .A2(n10074), .ZN(n7307) );
  AOI21_X1 U8977 ( .B1(n8291), .B2(n10074), .A(n7307), .ZN(n7312) );
  NAND2_X1 U8978 ( .A1(n7368), .A2(n7308), .ZN(n7310) );
  NAND2_X1 U8979 ( .A1(n7310), .A2(n7309), .ZN(n7311) );
  NOR2_X1 U8980 ( .A1(n7311), .A2(n7312), .ZN(n8285) );
  AOI21_X1 U8981 ( .B1(n7312), .B2(n7311), .A(n8285), .ZN(n7323) );
  NAND2_X1 U8982 ( .A1(n7314), .A2(n7313), .ZN(n7316) );
  NAND2_X1 U8983 ( .A1(n7316), .A2(n7315), .ZN(n7318) );
  XNOR2_X1 U8984 ( .A(n8291), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n7317) );
  NOR2_X1 U8985 ( .A1(n7318), .A2(n7317), .ZN(n8290) );
  AOI211_X1 U8986 ( .C1(n7318), .C2(n7317), .A(n9740), .B(n8290), .ZN(n7321)
         );
  AND2_X1 U8987 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8183) );
  AOI21_X1 U8988 ( .B1(n9739), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8183), .ZN(
        n7319) );
  OAI21_X1 U8989 ( .B1(n9900), .B2(n8286), .A(n7319), .ZN(n7320) );
  NOR2_X1 U8990 ( .A1(n7321), .A2(n7320), .ZN(n7322) );
  OAI21_X1 U8991 ( .B1(n7323), .B2(n9741), .A(n7322), .ZN(P2_U3261) );
  INV_X1 U8992 ( .A(n7324), .ZN(n7883) );
  NAND2_X1 U8993 ( .A1(n7365), .A2(n7377), .ZN(n7886) );
  INV_X1 U8994 ( .A(n7980), .ZN(n7884) );
  NOR2_X1 U8995 ( .A1(n4479), .A2(n8529), .ZN(n7329) );
  OAI21_X1 U8996 ( .B1(n7325), .B2(n7883), .A(n7884), .ZN(n7328) );
  OAI22_X1 U8997 ( .A1(n7326), .A2(n8548), .B1(n8549), .B2(n8550), .ZN(n7327)
         );
  AOI21_X1 U8998 ( .B1(n7329), .B2(n7328), .A(n7327), .ZN(n9448) );
  OAI22_X1 U8999 ( .A1(n8555), .A2(n7331), .B1(n7330), .B2(n8556), .ZN(n7336)
         );
  INV_X1 U9000 ( .A(n7332), .ZN(n7333) );
  INV_X1 U9001 ( .A(n7365), .ZN(n9449) );
  OR2_X1 U9002 ( .A1(n7332), .A2(n7365), .ZN(n7378) );
  OAI211_X1 U9003 ( .C1(n7333), .C2(n9449), .A(n7378), .B(n9816), .ZN(n9447)
         );
  NOR2_X1 U9004 ( .A1(n9447), .A2(n7334), .ZN(n7335) );
  AOI211_X1 U9005 ( .C1(n8566), .C2(n7365), .A(n7336), .B(n7335), .ZN(n7341)
         );
  NAND2_X1 U9006 ( .A1(n7337), .A2(n8275), .ZN(n7338) );
  XNOR2_X1 U9007 ( .A(n7364), .B(n7980), .ZN(n9451) );
  NAND2_X1 U9008 ( .A1(n9451), .A2(n9764), .ZN(n7340) );
  OAI211_X1 U9009 ( .C1(n9448), .C2(n8518), .A(n7341), .B(n7340), .ZN(P2_U3282) );
  INV_X1 U9010 ( .A(n7763), .ZN(n7345) );
  OAI222_X1 U9011 ( .A1(n7404), .A2(n7343), .B1(n8131), .B2(n7345), .C1(
        P2_U3152), .C2(n7342), .ZN(P2_U3333) );
  OAI222_X1 U9012 ( .A1(P1_U3084), .A2(n7346), .B1(n9369), .B2(n7345), .C1(
        n7344), .C2(n9371), .ZN(P1_U3328) );
  XNOR2_X1 U9013 ( .A(n9499), .B(n9252), .ZN(n8969) );
  XNOR2_X1 U9014 ( .A(n8947), .B(n8969), .ZN(n9504) );
  INV_X1 U9015 ( .A(n9504), .ZN(n7363) );
  AND2_X1 U9016 ( .A1(n7554), .A2(n7349), .ZN(n7459) );
  NAND2_X1 U9017 ( .A1(n7350), .A2(n7459), .ZN(n7351) );
  NAND2_X1 U9018 ( .A1(n7351), .A2(n7533), .ZN(n8970) );
  XNOR2_X1 U9019 ( .A(n8970), .B(n8969), .ZN(n7352) );
  NAND2_X1 U9020 ( .A1(n7352), .A2(n9470), .ZN(n7354) );
  AOI22_X1 U9021 ( .A1(n8838), .A2(n9253), .B1(n9254), .B2(n9229), .ZN(n7353)
         );
  NAND2_X1 U9022 ( .A1(n7354), .A2(n7353), .ZN(n9503) );
  AND2_X1 U9023 ( .A1(n7355), .A2(n9499), .ZN(n7356) );
  OR2_X1 U9024 ( .A1(n7356), .A2(n9260), .ZN(n9501) );
  OAI22_X1 U9025 ( .A1(n9479), .A2(n7358), .B1(n7357), .B2(n9476), .ZN(n7359)
         );
  AOI21_X1 U9026 ( .B1(n9499), .B2(n9264), .A(n7359), .ZN(n7360) );
  OAI21_X1 U9027 ( .B1(n9501), .B2(n9239), .A(n7360), .ZN(n7361) );
  AOI21_X1 U9028 ( .B1(n9503), .B2(n9269), .A(n7361), .ZN(n7362) );
  OAI21_X1 U9029 ( .B1(n7363), .B2(n9271), .A(n7362), .ZN(P1_U3278) );
  OR2_X1 U9030 ( .A1(n7365), .A2(n8274), .ZN(n7366) );
  NAND2_X1 U9031 ( .A1(n7367), .A2(n7787), .ZN(n7370) );
  AOI22_X1 U9032 ( .A1(n7703), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7368), .B2(
        n7714), .ZN(n7369) );
  NAND2_X1 U9033 ( .A1(n8260), .A2(n8549), .ZN(n7892) );
  NAND2_X1 U9034 ( .A1(n7891), .A2(n7892), .ZN(n7982) );
  NAND2_X1 U9035 ( .A1(n7371), .A2(n7982), .ZN(n8024) );
  OAI21_X1 U9036 ( .B1(n7371), .B2(n7982), .A(n8024), .ZN(n8649) );
  INV_X1 U9037 ( .A(n8649), .ZN(n7386) );
  NAND2_X1 U9038 ( .A1(n4401), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7375) );
  INV_X1 U9039 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7694) );
  XNOR2_X1 U9040 ( .A(n7695), .B(n7694), .ZN(n8557) );
  OR2_X1 U9041 ( .A1(n8557), .A2(n7768), .ZN(n7374) );
  INV_X1 U9042 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8558) );
  OR2_X1 U9043 ( .A1(n7771), .A2(n8558), .ZN(n7373) );
  OR2_X1 U9044 ( .A1(n7802), .A2(n10074), .ZN(n7372) );
  XNOR2_X1 U9045 ( .A(n7686), .B(n7982), .ZN(n7376) );
  OAI222_X1 U9046 ( .A1(n8548), .A2(n7377), .B1(n8550), .B2(n8047), .C1(n8529), 
        .C2(n7376), .ZN(n8647) );
  INV_X1 U9047 ( .A(n8260), .ZN(n8645) );
  INV_X1 U9048 ( .A(n7378), .ZN(n7380) );
  INV_X1 U9049 ( .A(n8559), .ZN(n7379) );
  OAI21_X1 U9050 ( .B1(n8645), .B2(n7380), .A(n7379), .ZN(n8646) );
  OAI22_X1 U9051 ( .A1(n9768), .A2(n7381), .B1(n8254), .B2(n8556), .ZN(n7382)
         );
  AOI21_X1 U9052 ( .B1(n8260), .B2(n8566), .A(n7382), .ZN(n7383) );
  OAI21_X1 U9053 ( .B1(n8646), .B2(n8562), .A(n7383), .ZN(n7384) );
  AOI21_X1 U9054 ( .B1(n8647), .B2(n9768), .A(n7384), .ZN(n7385) );
  OAI21_X1 U9055 ( .B1(n7386), .B2(n8541), .A(n7385), .ZN(P2_U3281) );
  INV_X1 U9056 ( .A(n7775), .ZN(n7390) );
  OAI222_X1 U9057 ( .A1(n7404), .A2(n7388), .B1(n8131), .B2(n7390), .C1(
        P2_U3152), .C2(n7387), .ZN(P2_U3332) );
  OAI222_X1 U9058 ( .A1(P1_U3084), .A2(n7391), .B1(n9369), .B2(n7390), .C1(
        n7389), .C2(n9371), .ZN(P1_U3327) );
  NAND2_X1 U9059 ( .A1(n7393), .A2(n7392), .ZN(n7394) );
  XOR2_X1 U9060 ( .A(n7395), .B(n7394), .Z(n7400) );
  OAI21_X1 U9061 ( .B1(n8830), .B2(n9208), .A(n7396), .ZN(n7398) );
  OAI22_X1 U9062 ( .A1(n8831), .A2(n9261), .B1(n7455), .B2(n8816), .ZN(n7397)
         );
  AOI211_X1 U9063 ( .C1(n9265), .C2(n8819), .A(n7398), .B(n7397), .ZN(n7399)
         );
  OAI21_X1 U9064 ( .B1(n7400), .B2(n8825), .A(n7399), .ZN(P1_U3213) );
  INV_X1 U9065 ( .A(n7788), .ZN(n7401) );
  OAI222_X1 U9066 ( .A1(P2_U3152), .A2(n8037), .B1(n8131), .B2(n7401), .C1(
        n7404), .C2(n5715), .ZN(P2_U3331) );
  OAI222_X1 U9067 ( .A1(n6274), .A2(P1_U3084), .B1(n9369), .B2(n7401), .C1(
        n9371), .C2(n5722), .ZN(P1_U3326) );
  INV_X1 U9068 ( .A(n7792), .ZN(n8085) );
  OAI222_X1 U9069 ( .A1(n7404), .A2(n7403), .B1(P2_U3152), .B2(n7402), .C1(
        n8131), .C2(n8085), .ZN(P2_U3330) );
  INV_X1 U9070 ( .A(SI_28_), .ZN(n7407) );
  NAND2_X1 U9071 ( .A1(n7408), .A2(n7407), .ZN(n7409) );
  INV_X1 U9072 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8682) );
  INV_X1 U9073 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9372) );
  MUX2_X1 U9074 ( .A(n8682), .B(n9372), .S(n7411), .Z(n7475) );
  INV_X1 U9075 ( .A(SI_29_), .ZN(n10016) );
  AND2_X1 U9076 ( .A1(n7475), .A2(n10016), .ZN(n7414) );
  INV_X1 U9077 ( .A(n7475), .ZN(n7412) );
  NAND2_X1 U9078 ( .A1(n7412), .A2(SI_29_), .ZN(n7413) );
  OAI21_X2 U9079 ( .B1(n7477), .B2(n7414), .A(n7413), .ZN(n7425) );
  XNOR2_X2 U9080 ( .A(n7425), .B(n7424), .ZN(n7423) );
  NAND2_X1 U9081 ( .A1(n8086), .A2(n7415), .ZN(n7417) );
  INV_X1 U9082 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10143) );
  OR2_X1 U9083 ( .A1(n7478), .A2(n10143), .ZN(n7416) );
  INV_X1 U9084 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10183) );
  NAND2_X1 U9085 ( .A1(n7418), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7420) );
  NAND2_X1 U9086 ( .A1(n5221), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7419) );
  OAI211_X1 U9087 ( .C1(n7421), .C2(n10183), .A(n7420), .B(n7419), .ZN(n8999)
         );
  INV_X1 U9088 ( .A(n8999), .ZN(n7487) );
  OR2_X1 U9089 ( .A1(n9275), .A2(n7487), .ZN(n7486) );
  NAND2_X1 U9090 ( .A1(n7486), .A2(n8938), .ZN(n7433) );
  INV_X1 U9091 ( .A(SI_30_), .ZN(n7422) );
  OR2_X2 U9092 ( .A1(n7423), .A2(n7422), .ZN(n7427) );
  NAND2_X1 U9093 ( .A1(n7425), .A2(n7424), .ZN(n7426) );
  MUX2_X1 U9094 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7428), .Z(n7429) );
  XNOR2_X1 U9095 ( .A(n7429), .B(SI_31_), .ZN(n7430) );
  NOR2_X1 U9096 ( .A1(n7478), .A2(n10000), .ZN(n7432) );
  NAND2_X1 U9097 ( .A1(n7433), .A2(n7485), .ZN(n7604) );
  NAND2_X1 U9098 ( .A1(n9297), .A2(n9076), .ZN(n9039) );
  INV_X1 U9099 ( .A(n9039), .ZN(n8991) );
  NAND2_X1 U9100 ( .A1(n9291), .A2(n9053), .ZN(n7488) );
  INV_X1 U9101 ( .A(n7488), .ZN(n7435) );
  NAND2_X1 U9102 ( .A1(n9285), .A2(n9037), .ZN(n7516) );
  INV_X1 U9103 ( .A(n7516), .ZN(n7434) );
  AOI211_X1 U9104 ( .C1(n8991), .C2(n8992), .A(n7435), .B(n7434), .ZN(n7654)
         );
  NAND2_X1 U9105 ( .A1(n9100), .A2(n8837), .ZN(n7589) );
  AND2_X1 U9106 ( .A1(n7589), .A2(n9101), .ZN(n8986) );
  NAND2_X1 U9107 ( .A1(n7588), .A2(n8986), .ZN(n7646) );
  NAND2_X1 U9108 ( .A1(n9317), .A2(n9130), .ZN(n8984) );
  AND2_X1 U9109 ( .A1(n9325), .A2(n9129), .ZN(n8982) );
  NAND2_X1 U9110 ( .A1(n7586), .A2(n8982), .ZN(n7436) );
  NAND2_X1 U9111 ( .A1(n9322), .A2(n9119), .ZN(n7584) );
  AND2_X1 U9112 ( .A1(n7436), .A2(n7584), .ZN(n7437) );
  NAND2_X1 U9113 ( .A1(n8984), .A2(n7437), .ZN(n7648) );
  NAND2_X1 U9114 ( .A1(n9330), .A2(n8955), .ZN(n8980) );
  INV_X1 U9115 ( .A(n8980), .ZN(n7439) );
  OR2_X1 U9116 ( .A1(n9335), .A2(n9200), .ZN(n7574) );
  OR2_X1 U9117 ( .A1(n9342), .A2(n8953), .ZN(n9176) );
  NAND2_X1 U9118 ( .A1(n7574), .A2(n9176), .ZN(n8979) );
  NAND2_X1 U9119 ( .A1(n9335), .A2(n9200), .ZN(n8978) );
  NAND2_X1 U9120 ( .A1(n8979), .A2(n8978), .ZN(n7438) );
  OR2_X1 U9121 ( .A1(n9325), .A2(n9129), .ZN(n8981) );
  OR2_X1 U9122 ( .A1(n9330), .A2(n8955), .ZN(n7573) );
  AND2_X1 U9123 ( .A1(n8981), .A2(n7573), .ZN(n7578) );
  OAI211_X1 U9124 ( .C1(n7439), .C2(n7438), .A(n7586), .B(n7578), .ZN(n7644)
         );
  NAND2_X1 U9125 ( .A1(n9342), .A2(n8953), .ZN(n7568) );
  NAND2_X1 U9126 ( .A1(n9220), .A2(n9198), .ZN(n9194) );
  NAND2_X1 U9127 ( .A1(n7568), .A2(n9194), .ZN(n8977) );
  INV_X1 U9128 ( .A(n8977), .ZN(n7440) );
  NAND2_X1 U9129 ( .A1(n8978), .A2(n7440), .ZN(n7465) );
  NAND2_X1 U9130 ( .A1(n9242), .A2(n9208), .ZN(n8976) );
  NAND2_X1 U9131 ( .A1(n9265), .A2(n7454), .ZN(n7559) );
  NAND2_X1 U9132 ( .A1(n9499), .A2(n7455), .ZN(n8971) );
  NAND2_X1 U9133 ( .A1(n7559), .A2(n8971), .ZN(n7557) );
  NAND2_X1 U9134 ( .A1(n7533), .A2(n7441), .ZN(n7555) );
  INV_X1 U9135 ( .A(n7457), .ZN(n7542) );
  NOR2_X1 U9136 ( .A1(n7543), .A2(n7542), .ZN(n7442) );
  OR2_X1 U9137 ( .A1(n7555), .A2(n7442), .ZN(n7461) );
  NAND2_X1 U9138 ( .A1(n7537), .A2(n7526), .ZN(n7443) );
  OR3_X1 U9139 ( .A1(n7557), .A2(n7461), .A3(n7443), .ZN(n7444) );
  OR3_X1 U9140 ( .A1(n7465), .A2(n4690), .A3(n7444), .ZN(n7619) );
  AND2_X1 U9141 ( .A1(n7448), .A2(n7445), .ZN(n7628) );
  NAND3_X1 U9142 ( .A1(n7446), .A2(n7628), .A3(n7636), .ZN(n7453) );
  NAND2_X1 U9143 ( .A1(n7630), .A2(n7632), .ZN(n7449) );
  NAND3_X1 U9144 ( .A1(n7449), .A2(n7448), .A3(n7447), .ZN(n7450) );
  NAND3_X1 U9145 ( .A1(n7450), .A2(n7634), .A3(n7633), .ZN(n7489) );
  NAND2_X1 U9146 ( .A1(n7489), .A2(n7525), .ZN(n7452) );
  INV_X1 U9147 ( .A(n7635), .ZN(n7451) );
  AOI21_X1 U9148 ( .B1(n7453), .B2(n7452), .A(n7451), .ZN(n7466) );
  OR2_X1 U9149 ( .A1(n9220), .A2(n9198), .ZN(n7566) );
  OR2_X1 U9150 ( .A1(n9499), .A2(n7455), .ZN(n7456) );
  NAND2_X1 U9151 ( .A1(n8973), .A2(n7456), .ZN(n7558) );
  NAND2_X1 U9152 ( .A1(n7457), .A2(n7538), .ZN(n7531) );
  INV_X1 U9153 ( .A(n7539), .ZN(n7530) );
  NOR2_X1 U9154 ( .A1(n7531), .A2(n7530), .ZN(n7460) );
  INV_X1 U9155 ( .A(n7533), .ZN(n7458) );
  OR2_X1 U9156 ( .A1(n7459), .A2(n7458), .ZN(n7549) );
  OAI21_X1 U9157 ( .B1(n7461), .B2(n7460), .A(n7549), .ZN(n7462) );
  NAND2_X1 U9158 ( .A1(n7557), .A2(n8973), .ZN(n7551) );
  OAI211_X1 U9159 ( .C1(n7558), .C2(n7462), .A(n7551), .B(n8976), .ZN(n7463)
         );
  AND3_X1 U9160 ( .A1(n7566), .A2(n8974), .A3(n7463), .ZN(n7464) );
  OR2_X1 U9161 ( .A1(n7465), .A2(n7464), .ZN(n7639) );
  OAI21_X1 U9162 ( .B1(n7619), .B2(n7466), .A(n7639), .ZN(n7467) );
  AND2_X1 U9163 ( .A1(n7467), .A2(n8980), .ZN(n7468) );
  NOR2_X1 U9164 ( .A1(n7644), .A2(n7468), .ZN(n7469) );
  NOR2_X1 U9165 ( .A1(n7648), .A2(n7469), .ZN(n7470) );
  NOR2_X1 U9166 ( .A1(n7646), .A2(n7470), .ZN(n7473) );
  AND2_X1 U9167 ( .A1(n9310), .A2(n9121), .ZN(n8985) );
  NAND2_X1 U9168 ( .A1(n7588), .A2(n8985), .ZN(n7471) );
  NAND2_X1 U9169 ( .A1(n9307), .A2(n9074), .ZN(n8987) );
  AND2_X1 U9170 ( .A1(n7471), .A2(n8987), .ZN(n7472) );
  NAND2_X1 U9171 ( .A1(n9302), .A2(n9083), .ZN(n8988) );
  NAND2_X1 U9172 ( .A1(n7472), .A2(n8988), .ZN(n7618) );
  OR2_X1 U9173 ( .A1(n9297), .A2(n9076), .ZN(n7595) );
  AND2_X1 U9174 ( .A1(n7595), .A2(n7593), .ZN(n7650) );
  OAI211_X1 U9175 ( .C1(n7473), .C2(n7618), .A(n8992), .B(n7650), .ZN(n7474)
         );
  AND2_X1 U9176 ( .A1(n7654), .A2(n7474), .ZN(n7482) );
  XNOR2_X1 U9177 ( .A(n7475), .B(SI_29_), .ZN(n7476) );
  NAND2_X1 U9178 ( .A1(n8681), .A2(n7415), .ZN(n7480) );
  OR2_X1 U9179 ( .A1(n7478), .A2(n9372), .ZN(n7479) );
  NAND2_X1 U9180 ( .A1(n7518), .A2(n8993), .ZN(n7660) );
  NAND2_X1 U9181 ( .A1(n9282), .A2(n9013), .ZN(n7658) );
  NAND2_X1 U9182 ( .A1(n8938), .A2(n8999), .ZN(n7481) );
  NAND2_X1 U9183 ( .A1(n9275), .A2(n7481), .ZN(n7603) );
  OAI211_X1 U9184 ( .C1(n7482), .C2(n7660), .A(n7658), .B(n7603), .ZN(n7483)
         );
  AND2_X1 U9185 ( .A1(n8939), .A2(n8938), .ZN(n7662) );
  AOI211_X1 U9186 ( .C1(n7604), .C2(n7483), .A(n7612), .B(n7662), .ZN(n7515)
         );
  INV_X1 U9187 ( .A(n8938), .ZN(n7484) );
  NAND2_X1 U9188 ( .A1(n7485), .A2(n7484), .ZN(n7523) );
  NAND2_X1 U9189 ( .A1(n7523), .A2(n7486), .ZN(n7617) );
  AND2_X1 U9190 ( .A1(n9275), .A2(n7487), .ZN(n7657) );
  NOR2_X1 U9191 ( .A1(n9310), .A2(n8837), .ZN(n8961) );
  OR2_X1 U9192 ( .A1(n8961), .A2(n4469), .ZN(n9092) );
  NAND2_X1 U9193 ( .A1(n7586), .A2(n7584), .ZN(n9127) );
  INV_X1 U9194 ( .A(n9127), .ZN(n7510) );
  INV_X1 U9195 ( .A(n8982), .ZN(n7575) );
  NAND2_X1 U9196 ( .A1(n7575), .A2(n8981), .ZN(n9140) );
  NAND2_X1 U9197 ( .A1(n7574), .A2(n8978), .ZN(n9168) );
  INV_X1 U9198 ( .A(n9168), .ZN(n9179) );
  NAND2_X1 U9199 ( .A1(n9176), .A2(n7568), .ZN(n7565) );
  NAND2_X1 U9200 ( .A1(n8973), .A2(n7559), .ZN(n9248) );
  INV_X1 U9201 ( .A(n8969), .ZN(n7504) );
  INV_X1 U9202 ( .A(n7489), .ZN(n7496) );
  AND4_X1 U9203 ( .A1(n7492), .A2(n7628), .A3(n7491), .A4(n7490), .ZN(n7495)
         );
  INV_X1 U9204 ( .A(n7493), .ZN(n7494) );
  NAND4_X1 U9205 ( .A1(n7496), .A2(n7495), .A3(n7494), .A4(n7636), .ZN(n7499)
         );
  NOR3_X1 U9206 ( .A1(n7499), .A2(n7498), .A3(n7497), .ZN(n7502) );
  XNOR2_X1 U9207 ( .A(n8783), .B(n8839), .ZN(n9464) );
  NAND4_X1 U9208 ( .A1(n7502), .A2(n7501), .A3(n7500), .A4(n9464), .ZN(n7503)
         );
  NOR3_X1 U9209 ( .A1(n9248), .A2(n7504), .A3(n7503), .ZN(n7505) );
  NAND3_X1 U9210 ( .A1(n9212), .A2(n9227), .A3(n7505), .ZN(n7506) );
  NOR2_X1 U9211 ( .A1(n7565), .A2(n7506), .ZN(n7507) );
  NAND3_X1 U9212 ( .A1(n9161), .A2(n9179), .A3(n7507), .ZN(n7508) );
  NOR2_X1 U9213 ( .A1(n9140), .A2(n7508), .ZN(n7509) );
  NAND4_X1 U9214 ( .A1(n9092), .A2(n9117), .A3(n7510), .A4(n7509), .ZN(n7511)
         );
  NOR4_X1 U9215 ( .A1(n9050), .A2(n9072), .A3(n9081), .A4(n7511), .ZN(n7512)
         );
  NAND4_X1 U9216 ( .A1(n8995), .A2(n9038), .A3(n9018), .A4(n7512), .ZN(n7513)
         );
  NOR2_X1 U9217 ( .A1(n7515), .A2(n7608), .ZN(n7611) );
  MUX2_X1 U9218 ( .A(n7516), .B(n8993), .S(n4499), .Z(n7517) );
  NAND2_X1 U9219 ( .A1(n8995), .A2(n7517), .ZN(n7601) );
  OAI21_X1 U9220 ( .B1(n7601), .B2(n8992), .A(n7518), .ZN(n7519) );
  NAND2_X1 U9221 ( .A1(n7519), .A2(n7603), .ZN(n7520) );
  NAND2_X1 U9222 ( .A1(n7604), .A2(n7520), .ZN(n7521) );
  NAND2_X1 U9223 ( .A1(n7521), .A2(n7602), .ZN(n7607) );
  INV_X1 U9224 ( .A(n7662), .ZN(n7522) );
  OAI21_X1 U9225 ( .B1(n7602), .B2(n7603), .A(n7522), .ZN(n7524) );
  NAND2_X1 U9226 ( .A1(n7524), .A2(n7523), .ZN(n7606) );
  INV_X1 U9227 ( .A(n7525), .ZN(n7527) );
  OAI211_X1 U9228 ( .C1(n7541), .C2(n7530), .A(n7537), .B(n7529), .ZN(n7536)
         );
  INV_X1 U9229 ( .A(n7531), .ZN(n7535) );
  NAND2_X1 U9230 ( .A1(n7533), .A2(n7532), .ZN(n7534) );
  AOI21_X1 U9231 ( .B1(n7536), .B2(n7535), .A(n7534), .ZN(n7546) );
  INV_X1 U9232 ( .A(n7537), .ZN(n7540) );
  OAI211_X1 U9233 ( .C1(n7541), .C2(n7540), .A(n7539), .B(n7538), .ZN(n7544)
         );
  AOI21_X1 U9234 ( .B1(n7544), .B2(n7543), .A(n7542), .ZN(n7545) );
  MUX2_X1 U9235 ( .A(n7546), .B(n7545), .S(n7602), .Z(n7548) );
  AND2_X1 U9236 ( .A1(n7554), .A2(n9464), .ZN(n7547) );
  NAND2_X1 U9237 ( .A1(n7548), .A2(n7547), .ZN(n7561) );
  INV_X1 U9238 ( .A(n7549), .ZN(n7550) );
  NOR2_X1 U9239 ( .A1(n7558), .A2(n7550), .ZN(n7553) );
  INV_X1 U9240 ( .A(n7551), .ZN(n7552) );
  AOI21_X1 U9241 ( .B1(n7561), .B2(n7553), .A(n7552), .ZN(n7563) );
  AND2_X1 U9242 ( .A1(n7555), .A2(n7554), .ZN(n7556) );
  NOR2_X1 U9243 ( .A1(n7557), .A2(n7556), .ZN(n7560) );
  AOI22_X1 U9244 ( .A1(n7561), .A2(n7560), .B1(n7559), .B2(n7558), .ZN(n7562)
         );
  MUX2_X1 U9245 ( .A(n8974), .B(n8976), .S(n7602), .Z(n7564) );
  MUX2_X1 U9246 ( .A(n9194), .B(n7566), .S(n7602), .Z(n7567) );
  NAND2_X1 U9247 ( .A1(n8978), .A2(n7568), .ZN(n7569) );
  MUX2_X1 U9248 ( .A(n8979), .B(n7569), .S(n7602), .Z(n7570) );
  INV_X1 U9249 ( .A(n7570), .ZN(n7571) );
  NAND2_X1 U9250 ( .A1(n7572), .A2(n7571), .ZN(n7577) );
  NAND3_X1 U9251 ( .A1(n7577), .A2(n7574), .A3(n7573), .ZN(n7576) );
  NAND3_X1 U9252 ( .A1(n7576), .A2(n8980), .A3(n7575), .ZN(n7581) );
  NAND3_X1 U9253 ( .A1(n7577), .A2(n8980), .A3(n8978), .ZN(n7579) );
  NAND2_X1 U9254 ( .A1(n7579), .A2(n7578), .ZN(n7580) );
  MUX2_X1 U9255 ( .A(n7581), .B(n7580), .S(n4499), .Z(n7585) );
  INV_X1 U9256 ( .A(n7586), .ZN(n7583) );
  INV_X1 U9257 ( .A(n7648), .ZN(n7582) );
  INV_X1 U9258 ( .A(n7584), .ZN(n8983) );
  NAND2_X1 U9259 ( .A1(n9101), .A2(n7586), .ZN(n7587) );
  INV_X1 U9260 ( .A(n9092), .ZN(n9103) );
  INV_X1 U9261 ( .A(n8987), .ZN(n7590) );
  OAI211_X1 U9262 ( .C1(n7590), .C2(n7589), .A(n7593), .B(n7588), .ZN(n7591)
         );
  MUX2_X1 U9263 ( .A(n7591), .B(n7618), .S(n7602), .Z(n7592) );
  MUX2_X1 U9264 ( .A(n8988), .B(n7593), .S(n7602), .Z(n7594) );
  NAND2_X1 U9265 ( .A1(n4699), .A2(n7594), .ZN(n7597) );
  MUX2_X1 U9266 ( .A(n7595), .B(n9039), .S(n7602), .Z(n7596) );
  OAI211_X1 U9267 ( .C1(n7598), .C2(n7597), .A(n9038), .B(n7596), .ZN(n7600)
         );
  NAND3_X1 U9268 ( .A1(n9291), .A2(n9053), .A3(n4499), .ZN(n7599) );
  NAND3_X1 U9269 ( .A1(n7607), .A2(n7606), .A3(n7605), .ZN(n7614) );
  INV_X1 U9270 ( .A(n7608), .ZN(n7609) );
  NOR3_X1 U9271 ( .A1(n7662), .A2(n5738), .A3(n7612), .ZN(n7613) );
  NAND2_X1 U9272 ( .A1(n7614), .A2(n7613), .ZN(n7616) );
  NAND2_X1 U9273 ( .A1(n7616), .A2(n7615), .ZN(n7667) );
  INV_X1 U9274 ( .A(n7617), .ZN(n7664) );
  INV_X1 U9275 ( .A(n7618), .ZN(n7653) );
  INV_X1 U9276 ( .A(n7619), .ZN(n7642) );
  INV_X1 U9277 ( .A(n7620), .ZN(n7621) );
  OAI211_X1 U9278 ( .C1(n6592), .C2(n7622), .A(n4585), .B(n7621), .ZN(n7624)
         );
  NAND2_X1 U9279 ( .A1(n7624), .A2(n7623), .ZN(n7626) );
  OAI22_X1 U9280 ( .A1(n7627), .A2(n7626), .B1(n7625), .B2(n5237), .ZN(n7631)
         );
  INV_X1 U9281 ( .A(n7628), .ZN(n7629) );
  AOI21_X1 U9282 ( .B1(n7631), .B2(n7630), .A(n7629), .ZN(n7638) );
  NAND3_X1 U9283 ( .A1(n7634), .A2(n7633), .A3(n7632), .ZN(n7637) );
  OAI211_X1 U9284 ( .C1(n7638), .C2(n7637), .A(n7636), .B(n7635), .ZN(n7641)
         );
  INV_X1 U9285 ( .A(n7639), .ZN(n7640) );
  AOI21_X1 U9286 ( .B1(n7642), .B2(n7641), .A(n7640), .ZN(n7643) );
  INV_X1 U9287 ( .A(n7643), .ZN(n7645) );
  AOI21_X1 U9288 ( .B1(n8980), .B2(n7645), .A(n7644), .ZN(n7649) );
  INV_X1 U9289 ( .A(n7646), .ZN(n7647) );
  OAI21_X1 U9290 ( .B1(n7649), .B2(n7648), .A(n7647), .ZN(n7652) );
  INV_X1 U9291 ( .A(n7650), .ZN(n7651) );
  AOI211_X1 U9292 ( .C1(n7653), .C2(n7652), .A(n7651), .B(n9030), .ZN(n7656)
         );
  INV_X1 U9293 ( .A(n7654), .ZN(n7655) );
  NOR2_X1 U9294 ( .A1(n7656), .A2(n7655), .ZN(n7661) );
  INV_X1 U9295 ( .A(n7657), .ZN(n7659) );
  OAI211_X1 U9296 ( .C1(n7661), .C2(n7660), .A(n7659), .B(n7658), .ZN(n7663)
         );
  AOI21_X1 U9297 ( .B1(n7664), .B2(n7663), .A(n7662), .ZN(n7665) );
  XNOR2_X1 U9298 ( .A(n7665), .B(n8929), .ZN(n7666) );
  NAND4_X1 U9299 ( .A1(n9253), .A2(n9678), .A3(n7668), .A4(n8936), .ZN(n7669)
         );
  OAI211_X1 U9300 ( .C1(n5738), .C2(n7671), .A(n7669), .B(P1_B_REG_SCAN_IN), 
        .ZN(n7670) );
  XNOR2_X1 U9301 ( .A(n8798), .B(n7672), .ZN(n7673) );
  NAND2_X1 U9302 ( .A1(n7673), .A2(n7674), .ZN(n8797) );
  OAI21_X1 U9303 ( .B1(n7674), .B2(n7673), .A(n8797), .ZN(n7675) );
  NAND2_X1 U9304 ( .A1(n7675), .A2(n8812), .ZN(n7680) );
  AND2_X1 U9305 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3084), .ZN(n9558) );
  OAI22_X1 U9306 ( .A1(n8831), .A2(n7677), .B1(n7676), .B2(n8816), .ZN(n7678)
         );
  AOI211_X1 U9307 ( .C1(n8807), .C2(n8844), .A(n9558), .B(n7678), .ZN(n7679)
         );
  OAI211_X1 U9308 ( .C1(n7681), .C2(n8836), .A(n7680), .B(n7679), .ZN(P1_U3225) );
  NAND2_X1 U9309 ( .A1(n8086), .A2(n7787), .ZN(n7683) );
  INV_X1 U9310 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9992) );
  OR2_X1 U9311 ( .A1(n7810), .A2(n9992), .ZN(n7682) );
  INV_X1 U9312 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n10068) );
  NAND2_X1 U9313 ( .A1(n4401), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7685) );
  NAND2_X1 U9314 ( .A1(n7798), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7684) );
  OAI211_X1 U9315 ( .C1(n7802), .C2(n10068), .A(n7685), .B(n7684), .ZN(n8265)
         );
  NAND2_X1 U9316 ( .A1(n8577), .A2(n8265), .ZN(n7954) );
  NAND2_X1 U9317 ( .A1(n7687), .A2(n7787), .ZN(n7689) );
  AOI22_X1 U9318 ( .A1(n7703), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7714), .B2(
        n8291), .ZN(n7688) );
  NAND2_X1 U9319 ( .A1(n8565), .A2(n8047), .ZN(n7894) );
  OR2_X1 U9320 ( .A1(n8565), .A2(n8047), .ZN(n7890) );
  INV_X1 U9321 ( .A(n7890), .ZN(n7896) );
  NAND2_X1 U9322 ( .A1(n7690), .A2(n7787), .ZN(n7692) );
  AOI22_X1 U9323 ( .A1(n7703), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7714), .B2(
        n8308), .ZN(n7691) );
  INV_X1 U9324 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7693) );
  OAI21_X1 U9325 ( .B1(n7695), .B2(n7694), .A(n7693), .ZN(n7696) );
  AND2_X1 U9326 ( .A1(n7696), .A2(n7706), .ZN(n8534) );
  NAND2_X1 U9327 ( .A1(n8534), .A2(n7780), .ZN(n7701) );
  NAND2_X1 U9328 ( .A1(n4407), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7700) );
  NAND2_X1 U9329 ( .A1(n4401), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7699) );
  INV_X1 U9330 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7697) );
  OR2_X1 U9331 ( .A1(n7771), .A2(n7697), .ZN(n7698) );
  NAND2_X1 U9332 ( .A1(n8641), .A2(n8551), .ZN(n7898) );
  NAND2_X1 U9333 ( .A1(n7899), .A2(n7898), .ZN(n8526) );
  OAI21_X1 U9334 ( .B1(n8527), .B2(n8526), .A(n7899), .ZN(n8513) );
  NAND2_X1 U9335 ( .A1(n7702), .A2(n7787), .ZN(n7705) );
  AOI22_X1 U9336 ( .A1(n7703), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7714), .B2(
        n8314), .ZN(n7704) );
  INV_X1 U9337 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n10036) );
  INV_X1 U9338 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10150) );
  NAND2_X1 U9339 ( .A1(n7706), .A2(n10150), .ZN(n7707) );
  NAND2_X1 U9340 ( .A1(n7717), .A2(n7707), .ZN(n8507) );
  OR2_X1 U9341 ( .A1(n8507), .A2(n7768), .ZN(n7712) );
  INV_X1 U9342 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n10142) );
  OR2_X1 U9343 ( .A1(n7783), .A2(n10142), .ZN(n7710) );
  INV_X1 U9344 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n7708) );
  OR2_X1 U9345 ( .A1(n7771), .A2(n7708), .ZN(n7709) );
  AND2_X1 U9346 ( .A1(n7710), .A2(n7709), .ZN(n7711) );
  OAI211_X1 U9347 ( .C1(n7802), .C2(n10036), .A(n7712), .B(n7711), .ZN(n8272)
         );
  INV_X1 U9348 ( .A(n8272), .ZN(n8027) );
  NAND2_X1 U9349 ( .A1(n8634), .A2(n8027), .ZN(n7906) );
  NAND2_X1 U9350 ( .A1(n8513), .A2(n8512), .ZN(n8511) );
  NAND2_X1 U9351 ( .A1(n7713), .A2(n7787), .ZN(n7716) );
  AOI22_X1 U9352 ( .A1(n7703), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8393), .B2(
        n7714), .ZN(n7715) );
  NAND2_X1 U9353 ( .A1(n7717), .A2(n10040), .ZN(n7718) );
  NAND2_X1 U9354 ( .A1(n7724), .A2(n7718), .ZN(n8493) );
  AOI22_X1 U9355 ( .A1(n4407), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n4401), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n7720) );
  INV_X1 U9356 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8494) );
  OR2_X1 U9357 ( .A1(n7771), .A2(n8494), .ZN(n7719) );
  OAI211_X1 U9358 ( .C1(n8493), .C2(n7768), .A(n7720), .B(n7719), .ZN(n8515)
         );
  INV_X1 U9359 ( .A(n8515), .ZN(n8481) );
  OR2_X1 U9360 ( .A1(n8631), .A2(n8481), .ZN(n7904) );
  NAND2_X1 U9361 ( .A1(n8631), .A2(n8481), .ZN(n8479) );
  NAND2_X1 U9362 ( .A1(n8511), .A2(n5006), .ZN(n8477) );
  NAND2_X1 U9363 ( .A1(n7721), .A2(n7787), .ZN(n7723) );
  NAND2_X1 U9364 ( .A1(n7703), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7722) );
  INV_X1 U9365 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8222) );
  NAND2_X1 U9366 ( .A1(n7724), .A2(n8222), .ZN(n7725) );
  NAND2_X1 U9367 ( .A1(n7726), .A2(n7725), .ZN(n8473) );
  OR2_X1 U9368 ( .A1(n8473), .A2(n7768), .ZN(n7729) );
  AOI22_X1 U9369 ( .A1(n4407), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n4401), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n7728) );
  NAND2_X1 U9370 ( .A1(n7798), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n7727) );
  NAND2_X1 U9371 ( .A1(n8624), .A2(n8461), .ZN(n7913) );
  NAND2_X1 U9372 ( .A1(n7917), .A2(n7913), .ZN(n8469) );
  INV_X1 U9373 ( .A(n8469), .ZN(n8478) );
  NAND2_X1 U9374 ( .A1(n8484), .A2(n7917), .ZN(n8459) );
  NAND2_X1 U9375 ( .A1(n7730), .A2(n7787), .ZN(n7732) );
  NAND2_X1 U9376 ( .A1(n7703), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7731) );
  OR2_X1 U9377 ( .A1(n8619), .A2(n8482), .ZN(n7916) );
  NAND2_X1 U9378 ( .A1(n8619), .A2(n8482), .ZN(n7919) );
  NAND2_X1 U9379 ( .A1(n7916), .A2(n7919), .ZN(n8458) );
  NAND2_X1 U9380 ( .A1(n7733), .A2(n7787), .ZN(n7735) );
  NAND2_X1 U9381 ( .A1(n7703), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n7734) );
  XNOR2_X1 U9382 ( .A(n7744), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n8443) );
  INV_X1 U9383 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U9384 ( .A1(n4401), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n7737) );
  NAND2_X1 U9385 ( .A1(n4407), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n7736) );
  OAI211_X1 U9386 ( .C1(n7771), .C2(n7738), .A(n7737), .B(n7736), .ZN(n7739)
         );
  NAND2_X1 U9387 ( .A1(n8613), .A2(n8462), .ZN(n7921) );
  NAND2_X1 U9388 ( .A1(n7740), .A2(n7787), .ZN(n7742) );
  NAND2_X1 U9389 ( .A1(n7703), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7741) );
  INV_X1 U9390 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8077) );
  INV_X1 U9391 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7743) );
  OAI21_X1 U9392 ( .B1(n7744), .B2(n8077), .A(n7743), .ZN(n7745) );
  NAND2_X1 U9393 ( .A1(n7756), .A2(n7745), .ZN(n8430) );
  OR2_X1 U9394 ( .A1(n8430), .A2(n7746), .ZN(n7751) );
  INV_X1 U9395 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8429) );
  NAND2_X1 U9396 ( .A1(n4407), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n7748) );
  NAND2_X1 U9397 ( .A1(n4401), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n7747) );
  OAI211_X1 U9398 ( .C1(n8429), .C2(n7771), .A(n7748), .B(n7747), .ZN(n7749)
         );
  INV_X1 U9399 ( .A(n7749), .ZN(n7750) );
  NAND2_X1 U9400 ( .A1(n7751), .A2(n7750), .ZN(n8450) );
  NOR2_X1 U9401 ( .A1(n8424), .A2(n4966), .ZN(n8423) );
  INV_X1 U9402 ( .A(n8450), .ZN(n8199) );
  AND2_X1 U9403 ( .A1(n8608), .A2(n8199), .ZN(n7925) );
  NAND2_X1 U9404 ( .A1(n7752), .A2(n7787), .ZN(n7754) );
  NAND2_X1 U9405 ( .A1(n7703), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7753) );
  INV_X1 U9406 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n7755) );
  NAND2_X1 U9407 ( .A1(n7756), .A2(n7755), .ZN(n7757) );
  NAND2_X1 U9408 ( .A1(n7766), .A2(n7757), .ZN(n8419) );
  OR2_X1 U9409 ( .A1(n8419), .A2(n7746), .ZN(n7762) );
  INV_X1 U9410 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n10160) );
  NAND2_X1 U9411 ( .A1(n7798), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n7759) );
  INV_X1 U9412 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n10091) );
  OR2_X1 U9413 ( .A1(n7783), .A2(n10091), .ZN(n7758) );
  OAI211_X1 U9414 ( .C1(n10160), .C2(n7802), .A(n7759), .B(n7758), .ZN(n7760)
         );
  INV_X1 U9415 ( .A(n7760), .ZN(n7761) );
  NAND2_X1 U9416 ( .A1(n8602), .A2(n8426), .ZN(n7926) );
  NAND2_X1 U9417 ( .A1(n7929), .A2(n7926), .ZN(n8407) );
  INV_X1 U9418 ( .A(n8407), .ZN(n8414) );
  NAND2_X1 U9419 ( .A1(n7763), .A2(n7787), .ZN(n7765) );
  NAND2_X1 U9420 ( .A1(n7703), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7764) );
  NAND2_X1 U9421 ( .A1(n7766), .A2(n8169), .ZN(n7767) );
  NAND2_X1 U9422 ( .A1(n7778), .A2(n7767), .ZN(n8396) );
  INV_X1 U9423 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U9424 ( .A1(n4407), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U9425 ( .A1(n4401), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n7769) );
  OAI211_X1 U9426 ( .C1(n8395), .C2(n7771), .A(n7770), .B(n7769), .ZN(n7772)
         );
  INV_X1 U9427 ( .A(n7772), .ZN(n7773) );
  XNOR2_X1 U9428 ( .A(n8599), .B(n8200), .ZN(n8032) );
  NAND2_X1 U9429 ( .A1(n7775), .A2(n7787), .ZN(n7777) );
  NAND2_X1 U9430 ( .A1(n7703), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7776) );
  NAND2_X1 U9431 ( .A1(n7778), .A2(n10185), .ZN(n7779) );
  NAND2_X1 U9432 ( .A1(n8384), .A2(n7780), .ZN(n7786) );
  INV_X1 U9433 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n10085) );
  NAND2_X1 U9434 ( .A1(n4407), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n7782) );
  NAND2_X1 U9435 ( .A1(n7798), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n7781) );
  OAI211_X1 U9436 ( .C1(n7783), .C2(n10085), .A(n7782), .B(n7781), .ZN(n7784)
         );
  INV_X1 U9437 ( .A(n7784), .ZN(n7785) );
  NAND2_X1 U9438 ( .A1(n8593), .A2(n8367), .ZN(n8364) );
  OR2_X1 U9439 ( .A1(n8599), .A2(n8200), .ZN(n8375) );
  NAND2_X1 U9440 ( .A1(n7788), .A2(n7787), .ZN(n7790) );
  NAND2_X1 U9441 ( .A1(n7703), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7789) );
  NAND2_X1 U9442 ( .A1(n8587), .A2(n8240), .ZN(n7939) );
  INV_X1 U9443 ( .A(n7791), .ZN(n7942) );
  NAND2_X1 U9444 ( .A1(n7792), .A2(n7787), .ZN(n7794) );
  NAND2_X1 U9445 ( .A1(n7703), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7793) );
  INV_X1 U9446 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8138) );
  INV_X1 U9447 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8127) );
  OAI21_X1 U9448 ( .B1(n7795), .B2(n8138), .A(n8127), .ZN(n7796) );
  NAND2_X1 U9449 ( .A1(n7797), .A2(n7796), .ZN(n8347) );
  INV_X1 U9450 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10066) );
  NAND2_X1 U9451 ( .A1(n7798), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n7801) );
  NAND2_X1 U9452 ( .A1(n4401), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7800) );
  OAI211_X1 U9453 ( .C1(n7802), .C2(n10066), .A(n7801), .B(n7800), .ZN(n7803)
         );
  INV_X1 U9454 ( .A(n7803), .ZN(n7804) );
  NAND2_X1 U9455 ( .A1(n8681), .A2(n7787), .ZN(n7808) );
  NAND2_X1 U9456 ( .A1(n7703), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7807) );
  NAND2_X1 U9457 ( .A1(n8579), .A2(n8124), .ZN(n7946) );
  INV_X1 U9458 ( .A(n7946), .ZN(n7809) );
  NAND2_X1 U9459 ( .A1(n9363), .A2(n7787), .ZN(n7812) );
  OR2_X1 U9460 ( .A1(n7810), .A2(n6119), .ZN(n7811) );
  INV_X1 U9461 ( .A(n8335), .ZN(n7814) );
  INV_X1 U9462 ( .A(n8577), .ZN(n8340) );
  INV_X1 U9463 ( .A(n8265), .ZN(n7813) );
  NAND2_X1 U9464 ( .A1(n8340), .A2(n7813), .ZN(n7948) );
  AND2_X1 U9465 ( .A1(n8570), .A2(n7814), .ZN(n7953) );
  INV_X1 U9466 ( .A(n7818), .ZN(n7957) );
  NOR2_X1 U9467 ( .A1(n8385), .A2(n7994), .ZN(n7820) );
  NAND2_X1 U9468 ( .A1(n7820), .A2(n7819), .ZN(n7821) );
  INV_X1 U9469 ( .A(n7821), .ZN(n7841) );
  INV_X1 U9470 ( .A(n7841), .ZN(n7956) );
  INV_X1 U9471 ( .A(n7940), .ZN(n7944) );
  INV_X1 U9472 ( .A(n7931), .ZN(n7938) );
  INV_X1 U9473 ( .A(n7823), .ZN(n7822) );
  AOI21_X1 U9474 ( .B1(n9796), .B2(n8284), .A(n7822), .ZN(n7827) );
  NAND2_X1 U9475 ( .A1(n7830), .A2(n7829), .ZN(n7825) );
  NAND2_X1 U9476 ( .A1(n7823), .A2(n7826), .ZN(n7824) );
  MUX2_X1 U9477 ( .A(n7825), .B(n7824), .S(n7821), .Z(n7839) );
  OAI211_X1 U9478 ( .C1(n7827), .C2(n7839), .A(n7826), .B(n7848), .ZN(n7850)
         );
  INV_X1 U9479 ( .A(n7830), .ZN(n7832) );
  INV_X1 U9480 ( .A(n7851), .ZN(n7831) );
  NAND3_X1 U9481 ( .A1(n7959), .A2(n7962), .A3(n7833), .ZN(n7844) );
  INV_X1 U9482 ( .A(n7845), .ZN(n7834) );
  AOI21_X1 U9483 ( .B1(n7835), .B2(n7844), .A(n7834), .ZN(n7838) );
  NAND2_X1 U9484 ( .A1(n7842), .A2(n7956), .ZN(n7837) );
  OAI21_X1 U9485 ( .B1(n7838), .B2(n7837), .A(n7836), .ZN(n7840) );
  NAND3_X1 U9486 ( .A1(n7844), .A2(n7843), .A3(n7842), .ZN(n7846) );
  NAND3_X1 U9487 ( .A1(n7846), .A2(n7841), .A3(n7845), .ZN(n7847) );
  AOI21_X1 U9488 ( .B1(n7841), .B2(n7850), .A(n7849), .ZN(n7856) );
  OAI21_X1 U9489 ( .B1(n7956), .B2(n7851), .A(n7971), .ZN(n7855) );
  MUX2_X1 U9490 ( .A(n7853), .B(n7852), .S(n7821), .Z(n7854) );
  OAI211_X1 U9491 ( .C1(n7856), .C2(n7855), .A(n7970), .B(n7854), .ZN(n7860)
         );
  MUX2_X1 U9492 ( .A(n7858), .B(n7857), .S(n7956), .Z(n7859) );
  NAND3_X1 U9493 ( .A1(n7860), .A2(n7861), .A3(n7859), .ZN(n7871) );
  INV_X1 U9494 ( .A(n7866), .ZN(n7870) );
  NAND2_X1 U9495 ( .A1(n7874), .A2(n7862), .ZN(n7868) );
  OAI211_X1 U9496 ( .C1(n7866), .C2(n7865), .A(n7864), .B(n7863), .ZN(n7867)
         );
  MUX2_X1 U9497 ( .A(n7868), .B(n7867), .S(n7821), .Z(n7869) );
  INV_X1 U9498 ( .A(n7872), .ZN(n7873) );
  OAI21_X1 U9499 ( .B1(n7878), .B2(n7873), .A(n7875), .ZN(n7880) );
  NAND2_X1 U9500 ( .A1(n7875), .A2(n7874), .ZN(n7877) );
  OAI21_X1 U9501 ( .B1(n7878), .B2(n7877), .A(n7876), .ZN(n7879) );
  INV_X1 U9502 ( .A(n7881), .ZN(n7882) );
  MUX2_X1 U9503 ( .A(n7883), .B(n7882), .S(n7821), .Z(n7885) );
  INV_X1 U9504 ( .A(n7982), .ZN(n7889) );
  MUX2_X1 U9505 ( .A(n7887), .B(n7886), .S(n7821), .Z(n7888) );
  MUX2_X1 U9506 ( .A(n7892), .B(n7891), .S(n7956), .Z(n7893) );
  INV_X1 U9507 ( .A(n7894), .ZN(n7895) );
  MUX2_X1 U9508 ( .A(n7896), .B(n7895), .S(n7956), .Z(n7897) );
  NOR2_X1 U9509 ( .A1(n7897), .A2(n8526), .ZN(n7903) );
  NAND2_X1 U9510 ( .A1(n7906), .A2(n7898), .ZN(n7901) );
  INV_X1 U9511 ( .A(n7899), .ZN(n7900) );
  MUX2_X1 U9512 ( .A(n7901), .B(n7900), .S(n7821), .Z(n7902) );
  NAND2_X1 U9513 ( .A1(n7904), .A2(n8498), .ZN(n7909) );
  OAI21_X1 U9514 ( .B1(n7908), .B2(n7909), .A(n8479), .ZN(n7905) );
  NAND2_X1 U9515 ( .A1(n7905), .A2(n7917), .ZN(n7912) );
  INV_X1 U9516 ( .A(n7906), .ZN(n7907) );
  OAI211_X1 U9517 ( .C1(n7910), .C2(n7909), .A(n8479), .B(n7913), .ZN(n7911)
         );
  MUX2_X1 U9518 ( .A(n7912), .B(n7911), .S(n7956), .Z(n7918) );
  NAND3_X1 U9519 ( .A1(n7918), .A2(n7913), .A3(n7919), .ZN(n7914) );
  NAND2_X1 U9520 ( .A1(n7914), .A2(n7916), .ZN(n7915) );
  NAND3_X1 U9521 ( .A1(n7918), .A2(n7917), .A3(n7916), .ZN(n7920) );
  NAND2_X1 U9522 ( .A1(n7920), .A2(n7919), .ZN(n7924) );
  INV_X1 U9523 ( .A(n7921), .ZN(n7922) );
  NAND2_X1 U9524 ( .A1(n7925), .A2(n7956), .ZN(n7927) );
  OAI21_X1 U9525 ( .B1(n8199), .B2(n8608), .A(n7929), .ZN(n7928) );
  NAND3_X1 U9526 ( .A1(n8602), .A2(n8426), .A3(n7841), .ZN(n7930) );
  NAND2_X1 U9527 ( .A1(n4947), .A2(n7930), .ZN(n7933) );
  NAND3_X1 U9528 ( .A1(n8394), .A2(n7841), .A3(n8416), .ZN(n7932) );
  OAI211_X1 U9529 ( .C1(n7934), .C2(n7933), .A(n7932), .B(n7931), .ZN(n7936)
         );
  OAI21_X1 U9530 ( .B1(n8394), .B2(n8416), .A(n8364), .ZN(n7935) );
  AOI22_X1 U9531 ( .A1(n7936), .A2(n8364), .B1(n7956), .B2(n7935), .ZN(n7937)
         );
  NAND2_X1 U9532 ( .A1(n7940), .A2(n7939), .ZN(n7941) );
  MUX2_X1 U9533 ( .A(n7942), .B(n7941), .S(n7821), .Z(n7943) );
  MUX2_X1 U9534 ( .A(n7946), .B(n7945), .S(n7956), .Z(n7947) );
  NAND3_X1 U9535 ( .A1(n7949), .A2(n7954), .A3(n7948), .ZN(n7952) );
  INV_X1 U9536 ( .A(n7953), .ZN(n7955) );
  NAND2_X1 U9537 ( .A1(n7955), .A2(n7954), .ZN(n7958) );
  INV_X1 U9538 ( .A(n7958), .ZN(n7989) );
  INV_X1 U9539 ( .A(n8447), .ZN(n8438) );
  INV_X1 U9540 ( .A(n8542), .ZN(n8546) );
  INV_X1 U9541 ( .A(n7959), .ZN(n7960) );
  NOR2_X1 U9542 ( .A1(n7961), .A2(n7960), .ZN(n9754) );
  NAND4_X1 U9543 ( .A1(n9754), .A2(n7964), .A3(n7963), .A4(n7962), .ZN(n7968)
         );
  NOR4_X1 U9544 ( .A1(n7968), .A2(n7967), .A3(n7966), .A4(n7965), .ZN(n7972)
         );
  NAND4_X1 U9545 ( .A1(n7972), .A2(n7971), .A3(n7970), .A4(n7969), .ZN(n7975)
         );
  NOR4_X1 U9546 ( .A1(n7976), .A2(n7975), .A3(n7974), .A4(n7973), .ZN(n7977)
         );
  NAND4_X1 U9547 ( .A1(n7980), .A2(n7979), .A3(n7978), .A4(n7977), .ZN(n7981)
         );
  NOR4_X1 U9548 ( .A1(n8526), .A2(n8546), .A3(n7982), .A4(n7981), .ZN(n7983)
         );
  NAND4_X1 U9549 ( .A1(n8478), .A2(n8512), .A3(n8497), .A4(n7983), .ZN(n7984)
         );
  NOR4_X1 U9550 ( .A1(n4966), .A2(n8438), .A3(n8458), .A4(n7984), .ZN(n7985)
         );
  NAND4_X1 U9551 ( .A1(n4938), .A2(n8414), .A3(n8377), .A4(n7985), .ZN(n7986)
         );
  NOR4_X1 U9552 ( .A1(n8036), .A2(n8352), .A3(n8032), .A4(n7986), .ZN(n7987)
         );
  NAND3_X1 U9553 ( .A1(n7989), .A2(n7988), .A3(n7987), .ZN(n7990) );
  XNOR2_X1 U9554 ( .A(n7990), .B(n8393), .ZN(n7995) );
  INV_X1 U9555 ( .A(n7991), .ZN(n7993) );
  AOI22_X1 U9556 ( .A1(n7995), .A2(n7994), .B1(n7993), .B2(n7992), .ZN(n7996)
         );
  INV_X1 U9557 ( .A(n7996), .ZN(n7997) );
  NAND2_X1 U9558 ( .A1(n7998), .A2(n7997), .ZN(n8001) );
  NAND3_X1 U9559 ( .A1(n7999), .A2(n7991), .A3(n5864), .ZN(n8000) );
  INV_X1 U9560 ( .A(n8037), .ZN(n8004) );
  NAND4_X1 U9561 ( .A1(n9771), .A2(n8004), .A3(n8003), .A4(n9751), .ZN(n8005)
         );
  OAI211_X1 U9562 ( .C1(n8007), .C2(n8006), .A(n8005), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8008) );
  INV_X1 U9563 ( .A(n8009), .ZN(n8010) );
  NAND2_X1 U9564 ( .A1(n8245), .A2(n8010), .ZN(n8013) );
  AND2_X1 U9565 ( .A1(P2_U3152), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9389) );
  AOI21_X1 U9566 ( .B1(n8011), .B2(P2_REG3_REG_2__SCAN_IN), .A(n9389), .ZN(
        n8012) );
  NAND2_X1 U9567 ( .A1(n8013), .A2(n8012), .ZN(n8019) );
  AOI22_X1 U9568 ( .A1(n8194), .A2(n6505), .B1(n8207), .B2(n8014), .ZN(n8017)
         );
  INV_X1 U9569 ( .A(n6379), .ZN(n8016) );
  NOR3_X1 U9570 ( .A1(n8017), .A2(n8016), .A3(n8015), .ZN(n8018) );
  AOI211_X1 U9571 ( .C1(n8020), .C2(n8259), .A(n8019), .B(n8018), .ZN(n8021)
         );
  OAI21_X1 U9572 ( .B1(n8022), .B2(n8263), .A(n8021), .ZN(P2_U3239) );
  INV_X1 U9573 ( .A(n8426), .ZN(n8268) );
  INV_X1 U9574 ( .A(n8047), .ZN(n8273) );
  NAND2_X1 U9575 ( .A1(n8645), .A2(n8549), .ZN(n8023) );
  INV_X1 U9576 ( .A(n8551), .ZN(n8514) );
  NAND2_X1 U9577 ( .A1(n8634), .A2(n8272), .ZN(n8026) );
  NAND2_X1 U9578 ( .A1(n8505), .A2(n8026), .ZN(n8029) );
  INV_X1 U9579 ( .A(n8634), .ZN(n8510) );
  NAND2_X1 U9580 ( .A1(n8510), .A2(n8027), .ZN(n8028) );
  INV_X1 U9581 ( .A(n8631), .ZN(n8492) );
  INV_X1 U9582 ( .A(n8461), .ZN(n8270) );
  AOI22_X2 U9583 ( .A1(n8470), .A2(n8469), .B1(n8624), .B2(n8270), .ZN(n8456)
         );
  NAND2_X1 U9584 ( .A1(n8619), .A2(n8449), .ZN(n8031) );
  INV_X1 U9585 ( .A(n8462), .ZN(n8269) );
  INV_X1 U9586 ( .A(n8367), .ZN(n8267) );
  INV_X1 U9587 ( .A(n8587), .ZN(n8363) );
  OAI22_X1 U9588 ( .A1(n8344), .A2(n8034), .B1(n8582), .B2(n8266), .ZN(n8035)
         );
  XOR2_X1 U9589 ( .A(n8036), .B(n4435), .Z(n8042) );
  NAND2_X1 U9590 ( .A1(n8266), .A2(n9751), .ZN(n8040) );
  INV_X1 U9591 ( .A(P2_B_REG_SCAN_IN), .ZN(n10173) );
  NOR2_X1 U9592 ( .A1(n8037), .A2(n10173), .ZN(n8038) );
  NOR2_X1 U9593 ( .A1(n8550), .A2(n8038), .ZN(n8334) );
  INV_X1 U9594 ( .A(n8602), .ZN(n8411) );
  INV_X1 U9595 ( .A(n8565), .ZN(n9442) );
  INV_X1 U9596 ( .A(n8624), .ZN(n8476) );
  NOR2_X1 U9597 ( .A1(n8599), .A2(n8392), .ZN(n8391) );
  AOI21_X1 U9598 ( .B1(n8579), .B2(n8345), .A(n8338), .ZN(n8580) );
  NAND2_X1 U9599 ( .A1(n8580), .A2(n8521), .ZN(n8045) );
  AOI22_X1 U9600 ( .A1(n8043), .A2(n9756), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n8535), .ZN(n8044) );
  OAI211_X1 U9601 ( .C1(n4612), .C2(n8538), .A(n8045), .B(n8044), .ZN(n8046)
         );
  XNOR2_X1 U9602 ( .A(n8565), .B(n8114), .ZN(n8050) );
  INV_X1 U9603 ( .A(n8050), .ZN(n8057) );
  NOR2_X1 U9604 ( .A1(n8047), .A2(n5905), .ZN(n8049) );
  INV_X1 U9605 ( .A(n8049), .ZN(n8056) );
  XNOR2_X1 U9606 ( .A(n8260), .B(n5934), .ZN(n8175) );
  OR2_X1 U9607 ( .A1(n8549), .A2(n5905), .ZN(n8177) );
  NAND2_X1 U9608 ( .A1(n8175), .A2(n8177), .ZN(n8054) );
  XNOR2_X1 U9609 ( .A(n8050), .B(n8049), .ZN(n8179) );
  INV_X1 U9610 ( .A(n8175), .ZN(n8052) );
  INV_X1 U9611 ( .A(n8177), .ZN(n8051) );
  XNOR2_X1 U9612 ( .A(n8641), .B(n8114), .ZN(n8060) );
  NAND2_X1 U9613 ( .A1(n8514), .A2(n8092), .ZN(n8058) );
  XNOR2_X1 U9614 ( .A(n8060), .B(n8058), .ZN(n8187) );
  INV_X1 U9615 ( .A(n8058), .ZN(n8059) );
  XNOR2_X1 U9616 ( .A(n8634), .B(n5934), .ZN(n8063) );
  NAND2_X1 U9617 ( .A1(n8272), .A2(n8092), .ZN(n8062) );
  XNOR2_X1 U9618 ( .A(n8063), .B(n8062), .ZN(n8227) );
  XNOR2_X1 U9619 ( .A(n8631), .B(n5934), .ZN(n8065) );
  NAND2_X1 U9620 ( .A1(n8515), .A2(n8092), .ZN(n8064) );
  NAND2_X1 U9621 ( .A1(n8065), .A2(n8064), .ZN(n8066) );
  OAI21_X1 U9622 ( .B1(n8065), .B2(n8064), .A(n8066), .ZN(n8151) );
  XNOR2_X1 U9623 ( .A(n8624), .B(n8114), .ZN(n8069) );
  NAND2_X1 U9624 ( .A1(n8270), .A2(n8092), .ZN(n8067) );
  XNOR2_X1 U9625 ( .A(n8069), .B(n8067), .ZN(n8220) );
  INV_X1 U9626 ( .A(n8067), .ZN(n8068) );
  AOI21_X2 U9627 ( .B1(n8221), .B2(n8220), .A(n8070), .ZN(n8158) );
  XNOR2_X1 U9628 ( .A(n8466), .B(n8114), .ZN(n8071) );
  NAND2_X1 U9629 ( .A1(n8449), .A2(n8092), .ZN(n8072) );
  XNOR2_X1 U9630 ( .A(n8071), .B(n8072), .ZN(n8157) );
  INV_X1 U9631 ( .A(n8071), .ZN(n8074) );
  INV_X1 U9632 ( .A(n8072), .ZN(n8073) );
  OAI21_X2 U9633 ( .B1(n8158), .B2(n8157), .A(n8075), .ZN(n8089) );
  XNOR2_X1 U9634 ( .A(n8613), .B(n8114), .ZN(n8088) );
  NAND2_X1 U9635 ( .A1(n8081), .A2(n5003), .ZN(n8091) );
  INV_X1 U9636 ( .A(n8443), .ZN(n8078) );
  OAI22_X1 U9637 ( .A1(n8078), .A2(n8253), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8077), .ZN(n8080) );
  OAI22_X1 U9638 ( .A1(n8199), .A2(n8230), .B1(n8482), .B2(n8231), .ZN(n8079)
         );
  AOI211_X1 U9639 ( .C1(n8613), .C2(n8259), .A(n8080), .B(n8079), .ZN(n8083)
         );
  OR3_X1 U9640 ( .A1(n8081), .A2(n8462), .A3(n8255), .ZN(n8082) );
  OAI211_X1 U9641 ( .C1(n8091), .C2(n8263), .A(n8083), .B(n8082), .ZN(P2_U3237) );
  OAI222_X1 U9642 ( .A1(n5773), .A2(P1_U3084), .B1(n9369), .B2(n8085), .C1(
        n8084), .C2(n9371), .ZN(P1_U3325) );
  INV_X1 U9643 ( .A(n8086), .ZN(n8130) );
  OAI222_X1 U9644 ( .A1(n9371), .A2(n10143), .B1(n9369), .B2(n8130), .C1(
        P1_U3084), .C2(n8087), .ZN(P1_U3323) );
  OR2_X1 U9645 ( .A1(n8089), .A2(n8088), .ZN(n8090) );
  NAND2_X2 U9646 ( .A1(n8091), .A2(n8090), .ZN(n8093) );
  XNOR2_X1 U9647 ( .A(n8608), .B(n5934), .ZN(n8094) );
  XNOR2_X2 U9648 ( .A(n8093), .B(n8094), .ZN(n8144) );
  NAND2_X1 U9649 ( .A1(n8450), .A2(n8092), .ZN(n8143) );
  OAI21_X2 U9650 ( .B1(n8144), .B2(n8143), .A(n8097), .ZN(n8100) );
  XNOR2_X1 U9651 ( .A(n8602), .B(n5934), .ZN(n8098) );
  NOR2_X1 U9652 ( .A1(n8426), .A2(n5905), .ZN(n8195) );
  NAND2_X1 U9653 ( .A1(n8196), .A2(n8195), .ZN(n8102) );
  INV_X1 U9654 ( .A(n8098), .ZN(n8099) );
  NAND2_X1 U9655 ( .A1(n8100), .A2(n8099), .ZN(n8101) );
  NAND2_X1 U9656 ( .A1(n8102), .A2(n8101), .ZN(n8168) );
  XNOR2_X1 U9657 ( .A(n8599), .B(n8114), .ZN(n8165) );
  NOR2_X1 U9658 ( .A1(n8200), .A2(n5905), .ZN(n8166) );
  XNOR2_X1 U9659 ( .A(n8593), .B(n8114), .ZN(n8133) );
  NOR2_X1 U9660 ( .A1(n8367), .A2(n5905), .ZN(n8103) );
  NAND2_X1 U9661 ( .A1(n8133), .A2(n8103), .ZN(n8106) );
  OAI21_X1 U9662 ( .B1(n8133), .B2(n8103), .A(n8106), .ZN(n8236) );
  XNOR2_X1 U9663 ( .A(n8587), .B(n8114), .ZN(n8107) );
  NOR2_X1 U9664 ( .A1(n8240), .A2(n5905), .ZN(n8108) );
  NAND2_X1 U9665 ( .A1(n8107), .A2(n8108), .ZN(n8113) );
  INV_X1 U9666 ( .A(n8107), .ZN(n8110) );
  INV_X1 U9667 ( .A(n8108), .ZN(n8109) );
  NAND2_X1 U9668 ( .A1(n8110), .A2(n8109), .ZN(n8111) );
  NOR2_X1 U9669 ( .A1(n8368), .A2(n5905), .ZN(n8115) );
  XNOR2_X1 U9670 ( .A(n8115), .B(n8114), .ZN(n8117) );
  INV_X1 U9671 ( .A(n8117), .ZN(n8118) );
  NOR3_X1 U9672 ( .A1(n8350), .A2(n8118), .A3(n8259), .ZN(n8116) );
  AOI21_X1 U9673 ( .B1(n8350), .B2(n8118), .A(n8116), .ZN(n8123) );
  OAI21_X1 U9674 ( .B1(n8350), .B2(n8248), .A(n8263), .ZN(n8122) );
  NOR3_X1 U9675 ( .A1(n8350), .A2(n8117), .A3(n8259), .ZN(n8120) );
  NOR2_X1 U9676 ( .A1(n8582), .A2(n8118), .ZN(n8119) );
  OR2_X1 U9677 ( .A1(n8240), .A2(n8548), .ZN(n8126) );
  OR2_X1 U9678 ( .A1(n8124), .A2(n8550), .ZN(n8125) );
  NAND2_X1 U9679 ( .A1(n8126), .A2(n8125), .ZN(n8354) );
  OAI22_X1 U9680 ( .A1(n8347), .A2(n8253), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8127), .ZN(n8128) );
  AOI21_X1 U9681 ( .B1(n8354), .B2(n8245), .A(n8128), .ZN(n8129) );
  OAI222_X1 U9682 ( .A1(n7404), .A2(n9992), .B1(n8131), .B2(n8130), .C1(n5888), 
        .C2(P2_U3152), .ZN(P2_U3328) );
  AOI21_X1 U9683 ( .B1(n8238), .B2(n4728), .A(n8263), .ZN(n8137) );
  INV_X1 U9684 ( .A(n8133), .ZN(n8134) );
  NOR3_X1 U9685 ( .A1(n8134), .A2(n8367), .A3(n8255), .ZN(n8136) );
  OAI21_X1 U9686 ( .B1(n8137), .B2(n8136), .A(n8135), .ZN(n8142) );
  OAI22_X1 U9687 ( .A1(n8367), .A2(n8231), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8138), .ZN(n8140) );
  NOR2_X1 U9688 ( .A1(n8368), .A2(n8230), .ZN(n8139) );
  AOI211_X1 U9689 ( .C1(n8211), .C2(n8361), .A(n8140), .B(n8139), .ZN(n8141)
         );
  OAI211_X1 U9690 ( .C1(n8363), .C2(n8248), .A(n8142), .B(n8141), .ZN(P2_U3216) );
  INV_X1 U9691 ( .A(n8608), .ZN(n8428) );
  NAND2_X1 U9692 ( .A1(n8143), .A2(n8207), .ZN(n8146) );
  NAND2_X1 U9693 ( .A1(n8450), .A2(n8194), .ZN(n8145) );
  MUX2_X1 U9694 ( .A(n8146), .B(n8145), .S(n8144), .Z(n8150) );
  NOR2_X1 U9695 ( .A1(n8430), .A2(n8253), .ZN(n8148) );
  OAI22_X1 U9696 ( .A1(n8426), .A2(n8230), .B1(n8462), .B2(n8231), .ZN(n8147)
         );
  AOI211_X1 U9697 ( .C1(P2_REG3_REG_23__SCAN_IN), .C2(P2_U3152), .A(n8148), 
        .B(n8147), .ZN(n8149) );
  OAI211_X1 U9698 ( .C1(n8428), .C2(n8248), .A(n8150), .B(n8149), .ZN(P2_U3218) );
  AOI21_X1 U9699 ( .B1(n8152), .B2(n8151), .A(n4484), .ZN(n8156) );
  NOR2_X1 U9700 ( .A1(n8253), .A2(n8493), .ZN(n8154) );
  AOI22_X1 U9701 ( .A1(n8270), .A2(n9752), .B1(n9751), .B2(n8272), .ZN(n8501)
         );
  INV_X1 U9702 ( .A(n8245), .ZN(n8189) );
  NAND2_X1 U9703 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8331) );
  OAI21_X1 U9704 ( .B1(n8501), .B2(n8189), .A(n8331), .ZN(n8153) );
  AOI211_X1 U9705 ( .C1(n8631), .C2(n8259), .A(n8154), .B(n8153), .ZN(n8155)
         );
  OAI21_X1 U9706 ( .B1(n8156), .B2(n8263), .A(n8155), .ZN(P2_U3221) );
  XNOR2_X1 U9707 ( .A(n8158), .B(n8157), .ZN(n8164) );
  INV_X1 U9708 ( .A(n8463), .ZN(n8160) );
  OAI22_X1 U9709 ( .A1(n8160), .A2(n8253), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8159), .ZN(n8162) );
  OAI22_X1 U9710 ( .A1(n8462), .A2(n8230), .B1(n8461), .B2(n8231), .ZN(n8161)
         );
  AOI211_X1 U9711 ( .C1(n8619), .C2(n8259), .A(n8162), .B(n8161), .ZN(n8163)
         );
  OAI21_X1 U9712 ( .B1(n8164), .B2(n8263), .A(n8163), .ZN(P2_U3225) );
  XOR2_X1 U9713 ( .A(n8166), .B(n8165), .Z(n8167) );
  XNOR2_X1 U9714 ( .A(n8168), .B(n8167), .ZN(n8173) );
  OAI22_X1 U9715 ( .A1(n8367), .A2(n8550), .B1(n8426), .B2(n8548), .ZN(n8401)
         );
  OAI22_X1 U9716 ( .A1(n8396), .A2(n8253), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8169), .ZN(n8171) );
  NOR2_X1 U9717 ( .A1(n8394), .A2(n8248), .ZN(n8170) );
  AOI211_X1 U9718 ( .C1(n8245), .C2(n8401), .A(n8171), .B(n8170), .ZN(n8172)
         );
  OAI21_X1 U9719 ( .B1(n8173), .B2(n8263), .A(n8172), .ZN(P2_U3227) );
  NAND2_X1 U9720 ( .A1(n8174), .A2(n8175), .ZN(n8178) );
  OR2_X1 U9721 ( .A1(n8174), .A2(n8175), .ZN(n8176) );
  AND2_X1 U9722 ( .A1(n8178), .A2(n8176), .ZN(n8256) );
  NAND2_X1 U9723 ( .A1(n8256), .A2(n8177), .ZN(n8262) );
  AND3_X1 U9724 ( .A1(n8262), .A2(n8179), .A3(n8178), .ZN(n8180) );
  OAI21_X1 U9725 ( .B1(n8181), .B2(n8180), .A(n8207), .ZN(n8186) );
  INV_X1 U9726 ( .A(n8557), .ZN(n8184) );
  OAI22_X1 U9727 ( .A1(n8549), .A2(n8231), .B1(n8230), .B2(n8551), .ZN(n8182)
         );
  AOI211_X1 U9728 ( .C1(n8184), .C2(n8211), .A(n8183), .B(n8182), .ZN(n8185)
         );
  OAI211_X1 U9729 ( .C1(n9442), .C2(n8248), .A(n8186), .B(n8185), .ZN(P2_U3228) );
  XNOR2_X1 U9730 ( .A(n8188), .B(n8187), .ZN(n8193) );
  AND2_X1 U9731 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8287) );
  AOI22_X1 U9732 ( .A1(n8273), .A2(n9751), .B1(n8272), .B2(n9752), .ZN(n8528)
         );
  NOR2_X1 U9733 ( .A1(n8189), .A2(n8528), .ZN(n8190) );
  AOI211_X1 U9734 ( .C1(n8211), .C2(n8534), .A(n8287), .B(n8190), .ZN(n8192)
         );
  NAND2_X1 U9735 ( .A1(n8641), .A2(n8259), .ZN(n8191) );
  OAI211_X1 U9736 ( .C1(n8193), .C2(n8263), .A(n8192), .B(n8191), .ZN(P2_U3230) );
  NAND2_X1 U9737 ( .A1(n8268), .A2(n8194), .ZN(n8198) );
  OR2_X1 U9738 ( .A1(n8195), .A2(n8263), .ZN(n8197) );
  MUX2_X1 U9739 ( .A(n8198), .B(n8197), .S(n8196), .Z(n8204) );
  NOR2_X1 U9740 ( .A1(n8419), .A2(n8253), .ZN(n8202) );
  OAI22_X1 U9741 ( .A1(n8200), .A2(n8230), .B1(n8199), .B2(n8231), .ZN(n8201)
         );
  AOI211_X1 U9742 ( .C1(P2_REG3_REG_24__SCAN_IN), .C2(P2_U3152), .A(n8202), 
        .B(n8201), .ZN(n8203) );
  OAI211_X1 U9743 ( .C1(n8411), .C2(n8248), .A(n8204), .B(n8203), .ZN(P2_U3231) );
  OAI21_X1 U9744 ( .B1(n8214), .B2(n8206), .A(n8205), .ZN(n8208) );
  NAND2_X1 U9745 ( .A1(n8208), .A2(n8207), .ZN(n8219) );
  AOI22_X1 U9746 ( .A1(n8259), .A2(n8209), .B1(P2_REG3_REG_4__SCAN_IN), .B2(
        P2_U3152), .ZN(n8218) );
  INV_X1 U9747 ( .A(n8210), .ZN(n8212) );
  AOI22_X1 U9748 ( .A1(n8250), .A2(n8282), .B1(n8212), .B2(n8211), .ZN(n8217)
         );
  NOR3_X1 U9749 ( .A1(n8255), .A2(n8214), .A3(n8213), .ZN(n8215) );
  OAI21_X1 U9750 ( .B1(n8215), .B2(n8249), .A(n8284), .ZN(n8216) );
  NAND4_X1 U9751 ( .A1(n8219), .A2(n8218), .A3(n8217), .A4(n8216), .ZN(
        P2_U3232) );
  XNOR2_X1 U9752 ( .A(n8221), .B(n8220), .ZN(n8226) );
  OAI22_X1 U9753 ( .A1(n8253), .A2(n8473), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8222), .ZN(n8224) );
  OAI22_X1 U9754 ( .A1(n8482), .A2(n8230), .B1(n8481), .B2(n8231), .ZN(n8223)
         );
  AOI211_X1 U9755 ( .C1(n8624), .C2(n8259), .A(n8224), .B(n8223), .ZN(n8225)
         );
  OAI21_X1 U9756 ( .B1(n8226), .B2(n8263), .A(n8225), .ZN(P2_U3235) );
  XNOR2_X1 U9757 ( .A(n8228), .B(n8227), .ZN(n8235) );
  NAND2_X1 U9758 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8311) );
  OAI21_X1 U9759 ( .B1(n8253), .B2(n8507), .A(n8311), .ZN(n8233) );
  OAI22_X1 U9760 ( .A1(n8551), .A2(n8231), .B1(n8230), .B2(n8481), .ZN(n8232)
         );
  AOI211_X1 U9761 ( .C1(n8634), .C2(n8259), .A(n8233), .B(n8232), .ZN(n8234)
         );
  OAI21_X1 U9762 ( .B1(n8235), .B2(n8263), .A(n8234), .ZN(P2_U3240) );
  AOI21_X1 U9763 ( .B1(n8237), .B2(n8236), .A(n8263), .ZN(n8239) );
  NAND2_X1 U9764 ( .A1(n8239), .A2(n8238), .ZN(n8247) );
  OR2_X1 U9765 ( .A1(n8240), .A2(n8550), .ZN(n8242) );
  NAND2_X1 U9766 ( .A1(n8416), .A2(n9751), .ZN(n8241) );
  NAND2_X1 U9767 ( .A1(n8242), .A2(n8241), .ZN(n8379) );
  INV_X1 U9768 ( .A(n8384), .ZN(n8243) );
  OAI22_X1 U9769 ( .A1(n8243), .A2(n8253), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10185), .ZN(n8244) );
  AOI21_X1 U9770 ( .B1(n8379), .B2(n8245), .A(n8244), .ZN(n8246) );
  OAI211_X1 U9771 ( .C1(n4950), .C2(n8248), .A(n8247), .B(n8246), .ZN(P2_U3242) );
  AOI22_X1 U9772 ( .A1(n8250), .A2(n8273), .B1(n8249), .B2(n8274), .ZN(n8252)
         );
  OAI211_X1 U9773 ( .C1(n8254), .C2(n8253), .A(n8252), .B(n8251), .ZN(n8258)
         );
  NOR3_X1 U9774 ( .A1(n8256), .A2(n8549), .A3(n8255), .ZN(n8257) );
  AOI211_X1 U9775 ( .C1(n8260), .C2(n8259), .A(n8258), .B(n8257), .ZN(n8261)
         );
  OAI21_X1 U9776 ( .B1(n8263), .B2(n8262), .A(n8261), .ZN(P2_U3243) );
  MUX2_X1 U9777 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8265), .S(n8264), .Z(
        P2_U3582) );
  MUX2_X1 U9778 ( .A(n8266), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8271), .Z(
        P2_U3580) );
  MUX2_X1 U9779 ( .A(n8267), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8271), .Z(
        P2_U3578) );
  MUX2_X1 U9780 ( .A(n8416), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8271), .Z(
        P2_U3577) );
  MUX2_X1 U9781 ( .A(n8268), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8271), .Z(
        P2_U3576) );
  MUX2_X1 U9782 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8450), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U9783 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8269), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9784 ( .A(n8270), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8271), .Z(
        P2_U3572) );
  MUX2_X1 U9785 ( .A(n8515), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8271), .Z(
        P2_U3571) );
  MUX2_X1 U9786 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8272), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9787 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8514), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9788 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8273), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9789 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8274), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9790 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8275), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9791 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8276), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9792 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8277), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9793 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8278), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9794 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8279), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9795 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8280), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9796 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n4535), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9797 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8281), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9798 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8282), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9799 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8283), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9800 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8284), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U9801 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n6506), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U9802 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6505), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U9803 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6484), .S(P2_U3966), .Z(
        P2_U3552) );
  INV_X1 U9804 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8304) );
  MUX2_X1 U9805 ( .A(n8304), .B(P2_REG1_REG_17__SCAN_IN), .S(n8308), .Z(n8299)
         );
  AOI21_X1 U9806 ( .B1(n10074), .B2(n8286), .A(n8285), .ZN(n8301) );
  XOR2_X1 U9807 ( .A(n8299), .B(n8301), .Z(n8298) );
  INV_X1 U9808 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8289) );
  INV_X1 U9809 ( .A(n8287), .ZN(n8288) );
  OAI21_X1 U9810 ( .B1(n9888), .B2(n8289), .A(n8288), .ZN(n8296) );
  AOI21_X1 U9811 ( .B1(n8291), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8290), .ZN(
        n8294) );
  NAND2_X1 U9812 ( .A1(n8308), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8292) );
  OAI21_X1 U9813 ( .B1(n8308), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8292), .ZN(
        n8293) );
  AOI211_X1 U9814 ( .C1(n8294), .C2(n8293), .A(n9740), .B(n8307), .ZN(n8295)
         );
  AOI211_X1 U9815 ( .C1(n9395), .C2(n8308), .A(n8296), .B(n8295), .ZN(n8297)
         );
  OAI21_X1 U9816 ( .B1(n9741), .B2(n8298), .A(n8297), .ZN(P2_U3262) );
  INV_X1 U9817 ( .A(n8299), .ZN(n8300) );
  NAND2_X1 U9818 ( .A1(n8301), .A2(n8300), .ZN(n8302) );
  OAI21_X1 U9819 ( .B1(n8304), .B2(n8303), .A(n8302), .ZN(n8306) );
  AOI22_X1 U9820 ( .A1(n8314), .A2(n10036), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8323), .ZN(n8305) );
  NOR2_X1 U9821 ( .A1(n8306), .A2(n8305), .ZN(n8322) );
  AOI21_X1 U9822 ( .B1(n8306), .B2(n8305), .A(n8322), .ZN(n8317) );
  OAI21_X1 U9823 ( .B1(n8309), .B2(n7708), .A(n8320), .ZN(n8310) );
  NAND2_X1 U9824 ( .A1(n8310), .A2(n9896), .ZN(n8316) );
  INV_X1 U9825 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8312) );
  OAI21_X1 U9826 ( .B1(n9888), .B2(n8312), .A(n8311), .ZN(n8313) );
  AOI21_X1 U9827 ( .B1(n9395), .B2(n8314), .A(n8313), .ZN(n8315) );
  OAI211_X1 U9828 ( .C1(n8317), .C2(n9741), .A(n8316), .B(n8315), .ZN(P2_U3263) );
  NAND2_X1 U9829 ( .A1(n8318), .A2(n8323), .ZN(n8319) );
  NAND2_X1 U9830 ( .A1(n8320), .A2(n8319), .ZN(n8321) );
  XNOR2_X1 U9831 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8321), .ZN(n8328) );
  INV_X1 U9832 ( .A(n8328), .ZN(n8326) );
  INV_X1 U9833 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n10042) );
  AOI21_X1 U9834 ( .B1(n8323), .B2(n10036), .A(n8322), .ZN(n8324) );
  XNOR2_X1 U9835 ( .A(n10042), .B(n8324), .ZN(n8327) );
  OAI21_X1 U9836 ( .B1(n8327), .B2(n9741), .A(n9900), .ZN(n8325) );
  AOI21_X1 U9837 ( .B1(n8326), .B2(n9896), .A(n8325), .ZN(n8330) );
  AOI22_X1 U9838 ( .A1(n8328), .A2(n9896), .B1(n9891), .B2(n8327), .ZN(n8329)
         );
  MUX2_X1 U9839 ( .A(n8330), .B(n8329), .S(n8385), .Z(n8332) );
  OAI211_X1 U9840 ( .C1(n4920), .C2(n9888), .A(n8332), .B(n8331), .ZN(P2_U3264) );
  NAND2_X1 U9841 ( .A1(n8577), .A2(n8338), .ZN(n8573) );
  XNOR2_X1 U9842 ( .A(n8573), .B(n8570), .ZN(n8572) );
  NOR2_X1 U9843 ( .A1(n9768), .A2(n8333), .ZN(n8336) );
  NAND2_X1 U9844 ( .A1(n8335), .A2(n8334), .ZN(n8575) );
  NOR2_X1 U9845 ( .A1(n8535), .A2(n8575), .ZN(n8341) );
  AOI211_X1 U9846 ( .C1(n8570), .C2(n8566), .A(n8336), .B(n8341), .ZN(n8337)
         );
  OAI21_X1 U9847 ( .B1(n8572), .B2(n8562), .A(n8337), .ZN(P2_U3265) );
  INV_X1 U9848 ( .A(n8338), .ZN(n8339) );
  NAND2_X1 U9849 ( .A1(n8340), .A2(n8339), .ZN(n8574) );
  NAND3_X1 U9850 ( .A1(n8574), .A2(n8521), .A3(n8573), .ZN(n8343) );
  AOI21_X1 U9851 ( .B1(n8518), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8341), .ZN(
        n8342) );
  OAI211_X1 U9852 ( .C1(n8577), .C2(n8538), .A(n8343), .B(n8342), .ZN(P2_U3266) );
  XNOR2_X1 U9853 ( .A(n8344), .B(n8352), .ZN(n8586) );
  INV_X1 U9854 ( .A(n8345), .ZN(n8346) );
  AOI21_X1 U9855 ( .B1(n8582), .B2(n4616), .A(n8346), .ZN(n8583) );
  INV_X1 U9856 ( .A(n8347), .ZN(n8348) );
  AOI22_X1 U9857 ( .A1(n8348), .A2(n9756), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n8535), .ZN(n8349) );
  OAI21_X1 U9858 ( .B1(n8350), .B2(n8538), .A(n8349), .ZN(n8357) );
  AOI211_X1 U9859 ( .C1(n8353), .C2(n8352), .A(n8529), .B(n8351), .ZN(n8355)
         );
  NOR2_X1 U9860 ( .A1(n8355), .A2(n8354), .ZN(n8585) );
  NOR2_X1 U9861 ( .A1(n8585), .A2(n8535), .ZN(n8356) );
  AOI211_X1 U9862 ( .C1(n8521), .C2(n8583), .A(n8357), .B(n8356), .ZN(n8358)
         );
  OAI21_X1 U9863 ( .B1(n8586), .B2(n8541), .A(n8358), .ZN(P2_U3268) );
  XNOR2_X1 U9864 ( .A(n8359), .B(n4938), .ZN(n8591) );
  AOI21_X1 U9865 ( .B1(n8587), .B2(n8381), .A(n8360), .ZN(n8588) );
  AOI22_X1 U9866 ( .A1(n8361), .A2(n9756), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n8535), .ZN(n8362) );
  OAI21_X1 U9867 ( .B1(n8363), .B2(n8538), .A(n8362), .ZN(n8372) );
  AOI21_X1 U9868 ( .B1(n8376), .B2(n8364), .A(n4938), .ZN(n8365) );
  NOR3_X1 U9869 ( .A1(n8366), .A2(n8365), .A3(n8529), .ZN(n8370) );
  OAI22_X1 U9870 ( .A1(n8368), .A2(n8550), .B1(n8367), .B2(n8548), .ZN(n8369)
         );
  NOR2_X1 U9871 ( .A1(n8370), .A2(n8369), .ZN(n8590) );
  NOR2_X1 U9872 ( .A1(n8590), .A2(n8518), .ZN(n8371) );
  AOI211_X1 U9873 ( .C1(n8521), .C2(n8588), .A(n8372), .B(n8371), .ZN(n8373)
         );
  OAI21_X1 U9874 ( .B1(n8591), .B2(n8541), .A(n8373), .ZN(P2_U3269) );
  XOR2_X1 U9875 ( .A(n8377), .B(n8374), .Z(n8596) );
  NOR2_X1 U9876 ( .A1(n4950), .A2(n8538), .ZN(n8388) );
  AND2_X1 U9877 ( .A1(n8399), .A2(n8375), .ZN(n8378) );
  OAI21_X1 U9878 ( .B1(n8378), .B2(n8377), .A(n8376), .ZN(n8380) );
  AOI21_X1 U9879 ( .B1(n8380), .B2(n9748), .A(n8379), .ZN(n8595) );
  INV_X1 U9880 ( .A(n8391), .ZN(n8383) );
  INV_X1 U9881 ( .A(n8381), .ZN(n8382) );
  AOI211_X1 U9882 ( .C1(n8593), .C2(n8383), .A(n9833), .B(n8382), .ZN(n8592)
         );
  AOI22_X1 U9883 ( .A1(n8592), .A2(n8385), .B1(n9756), .B2(n8384), .ZN(n8386)
         );
  AOI21_X1 U9884 ( .B1(n8595), .B2(n8386), .A(n8535), .ZN(n8387) );
  AOI211_X1 U9885 ( .C1(n8518), .C2(P2_REG2_REG_26__SCAN_IN), .A(n8388), .B(
        n8387), .ZN(n8389) );
  OAI21_X1 U9886 ( .B1(n8596), .B2(n8541), .A(n8389), .ZN(P2_U3270) );
  XNOR2_X1 U9887 ( .A(n8390), .B(n4947), .ZN(n8601) );
  AOI211_X1 U9888 ( .C1(n8599), .C2(n8392), .A(n9833), .B(n8391), .ZN(n8598)
         );
  NOR2_X1 U9889 ( .A1(n8535), .A2(n8393), .ZN(n8533) );
  NOR2_X1 U9890 ( .A1(n8394), .A2(n8538), .ZN(n8398) );
  OAI22_X1 U9891 ( .A1(n8396), .A2(n8556), .B1(n8395), .B2(n8555), .ZN(n8397)
         );
  AOI211_X1 U9892 ( .C1(n8598), .C2(n8533), .A(n8398), .B(n8397), .ZN(n8405)
         );
  OAI211_X1 U9893 ( .C1(n8400), .C2(n4947), .A(n8399), .B(n9748), .ZN(n8403)
         );
  INV_X1 U9894 ( .A(n8401), .ZN(n8402) );
  NAND2_X1 U9895 ( .A1(n8403), .A2(n8402), .ZN(n8597) );
  NAND2_X1 U9896 ( .A1(n8597), .A2(n8555), .ZN(n8404) );
  OAI211_X1 U9897 ( .C1(n8601), .C2(n8541), .A(n8405), .B(n8404), .ZN(P2_U3271) );
  OAI21_X1 U9898 ( .B1(n8408), .B2(n8407), .A(n8406), .ZN(n8409) );
  INV_X1 U9899 ( .A(n8409), .ZN(n8606) );
  XNOR2_X1 U9900 ( .A(n4476), .B(n8602), .ZN(n8603) );
  INV_X1 U9901 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8410) );
  OAI22_X1 U9902 ( .A1(n8411), .A2(n8538), .B1(n9768), .B2(n8410), .ZN(n8412)
         );
  AOI21_X1 U9903 ( .B1(n8521), .B2(n8603), .A(n8412), .ZN(n8422) );
  OAI211_X1 U9904 ( .C1(n8415), .C2(n8414), .A(n8413), .B(n9748), .ZN(n8418)
         );
  AOI22_X1 U9905 ( .A1(n8416), .A2(n9752), .B1(n9751), .B2(n8450), .ZN(n8417)
         );
  OAI21_X1 U9906 ( .B1(n8419), .B2(n8556), .A(n8605), .ZN(n8420) );
  NAND2_X1 U9907 ( .A1(n8420), .A2(n8555), .ZN(n8421) );
  OAI211_X1 U9908 ( .C1(n8606), .C2(n8541), .A(n8422), .B(n8421), .ZN(P2_U3272) );
  AOI21_X1 U9909 ( .B1(n4966), .B2(n8424), .A(n8423), .ZN(n8425) );
  OAI222_X1 U9910 ( .A1(n8548), .A2(n8462), .B1(n8550), .B2(n8426), .C1(n8529), 
        .C2(n8425), .ZN(n8427) );
  INV_X1 U9911 ( .A(n8427), .ZN(n8611) );
  AOI21_X1 U9912 ( .B1(n8608), .B2(n8440), .A(n4476), .ZN(n8609) );
  NOR2_X1 U9913 ( .A1(n8428), .A2(n8538), .ZN(n8432) );
  OAI22_X1 U9914 ( .A1(n8430), .A2(n8556), .B1(n8429), .B2(n8555), .ZN(n8431)
         );
  AOI211_X1 U9915 ( .C1(n8609), .C2(n8521), .A(n8432), .B(n8431), .ZN(n8437)
         );
  NAND2_X1 U9916 ( .A1(n8435), .A2(n8434), .ZN(n8607) );
  NAND3_X1 U9917 ( .A1(n4971), .A2(n9764), .A3(n8607), .ZN(n8436) );
  OAI211_X1 U9918 ( .C1(n8611), .C2(n8518), .A(n8437), .B(n8436), .ZN(P2_U3273) );
  XNOR2_X1 U9919 ( .A(n8439), .B(n8438), .ZN(n8617) );
  INV_X1 U9920 ( .A(n8440), .ZN(n8441) );
  AOI21_X1 U9921 ( .B1(n8613), .B2(n8442), .A(n8441), .ZN(n8614) );
  INV_X1 U9922 ( .A(n8613), .ZN(n8445) );
  AOI22_X1 U9923 ( .A1(n8535), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8443), .B2(
        n9756), .ZN(n8444) );
  OAI21_X1 U9924 ( .B1(n8445), .B2(n8538), .A(n8444), .ZN(n8454) );
  OAI211_X1 U9925 ( .C1(n8448), .C2(n8447), .A(n8446), .B(n9748), .ZN(n8452)
         );
  AOI22_X1 U9926 ( .A1(n8450), .A2(n9752), .B1(n9751), .B2(n8449), .ZN(n8451)
         );
  NOR2_X1 U9927 ( .A1(n8616), .A2(n8535), .ZN(n8453) );
  AOI211_X1 U9928 ( .C1(n8614), .C2(n8521), .A(n8454), .B(n8453), .ZN(n8455)
         );
  OAI21_X1 U9929 ( .B1(n8617), .B2(n8541), .A(n8455), .ZN(P2_U3274) );
  XOR2_X1 U9930 ( .A(n8458), .B(n8456), .Z(n8623) );
  AOI21_X1 U9931 ( .B1(n8459), .B2(n8458), .A(n8457), .ZN(n8460) );
  OAI222_X1 U9932 ( .A1(n8550), .A2(n8462), .B1(n8548), .B2(n8461), .C1(n8529), 
        .C2(n8460), .ZN(n8618) );
  XNOR2_X1 U9933 ( .A(n8471), .B(n8619), .ZN(n8620) );
  NAND2_X1 U9934 ( .A1(n8620), .A2(n8521), .ZN(n8465) );
  AOI22_X1 U9935 ( .A1(n8535), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8463), .B2(
        n9756), .ZN(n8464) );
  OAI211_X1 U9936 ( .C1(n8466), .C2(n8538), .A(n8465), .B(n8464), .ZN(n8467)
         );
  AOI21_X1 U9937 ( .B1(n8618), .B2(n9768), .A(n8467), .ZN(n8468) );
  OAI21_X1 U9938 ( .B1(n8623), .B2(n8541), .A(n8468), .ZN(P2_U3275) );
  XNOR2_X1 U9939 ( .A(n8470), .B(n8469), .ZN(n8628) );
  INV_X1 U9940 ( .A(n8491), .ZN(n8472) );
  AOI21_X1 U9941 ( .B1(n8624), .B2(n8472), .A(n8471), .ZN(n8625) );
  INV_X1 U9942 ( .A(n8473), .ZN(n8474) );
  AOI22_X1 U9943 ( .A1(n8535), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8474), .B2(
        n9756), .ZN(n8475) );
  OAI21_X1 U9944 ( .B1(n8476), .B2(n8538), .A(n8475), .ZN(n8487) );
  AOI21_X1 U9945 ( .B1(n8477), .B2(n8479), .A(n8478), .ZN(n8480) );
  NOR2_X1 U9946 ( .A1(n8480), .A2(n8529), .ZN(n8485) );
  OAI22_X1 U9947 ( .A1(n8482), .A2(n8550), .B1(n8481), .B2(n8548), .ZN(n8483)
         );
  AOI21_X1 U9948 ( .B1(n8485), .B2(n8484), .A(n8483), .ZN(n8627) );
  NOR2_X1 U9949 ( .A1(n8627), .A2(n8535), .ZN(n8486) );
  AOI211_X1 U9950 ( .C1(n8625), .C2(n8521), .A(n8487), .B(n8486), .ZN(n8488)
         );
  OAI21_X1 U9951 ( .B1(n8541), .B2(n8628), .A(n8488), .ZN(P2_U3276) );
  XOR2_X1 U9952 ( .A(n8497), .B(n8490), .Z(n8633) );
  AOI211_X1 U9953 ( .C1(n8631), .C2(n8506), .A(n9833), .B(n8491), .ZN(n8630)
         );
  NOR2_X1 U9954 ( .A1(n8492), .A2(n8538), .ZN(n8496) );
  OAI22_X1 U9955 ( .A1(n8555), .A2(n8494), .B1(n8493), .B2(n8556), .ZN(n8495)
         );
  AOI211_X1 U9956 ( .C1(n8630), .C2(n8533), .A(n8496), .B(n8495), .ZN(n8504)
         );
  INV_X1 U9957 ( .A(n8477), .ZN(n8500) );
  AOI21_X1 U9958 ( .B1(n8511), .B2(n8498), .A(n8497), .ZN(n8499) );
  OAI21_X1 U9959 ( .B1(n8500), .B2(n8499), .A(n9748), .ZN(n8502) );
  NAND2_X1 U9960 ( .A1(n8502), .A2(n8501), .ZN(n8629) );
  NAND2_X1 U9961 ( .A1(n8629), .A2(n8555), .ZN(n8503) );
  OAI211_X1 U9962 ( .C1(n8633), .C2(n8541), .A(n8504), .B(n8503), .ZN(P2_U3277) );
  XNOR2_X1 U9963 ( .A(n8505), .B(n8512), .ZN(n8638) );
  AOI21_X1 U9964 ( .B1(n8634), .B2(n8531), .A(n4622), .ZN(n8635) );
  INV_X1 U9965 ( .A(n8507), .ZN(n8508) );
  AOI22_X1 U9966 ( .A1(n8535), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8508), .B2(
        n9756), .ZN(n8509) );
  OAI21_X1 U9967 ( .B1(n8510), .B2(n8538), .A(n8509), .ZN(n8520) );
  OAI211_X1 U9968 ( .C1(n8513), .C2(n8512), .A(n8511), .B(n9748), .ZN(n8517)
         );
  AOI22_X1 U9969 ( .A1(n8515), .A2(n9752), .B1(n8514), .B2(n9751), .ZN(n8516)
         );
  AND2_X1 U9970 ( .A1(n8517), .A2(n8516), .ZN(n8637) );
  NOR2_X1 U9971 ( .A1(n8637), .A2(n8518), .ZN(n8519) );
  AOI211_X1 U9972 ( .C1(n8635), .C2(n8521), .A(n8520), .B(n8519), .ZN(n8522)
         );
  OAI21_X1 U9973 ( .B1(n8638), .B2(n8541), .A(n8522), .ZN(P2_U3278) );
  OAI21_X1 U9974 ( .B1(n8524), .B2(n8526), .A(n8523), .ZN(n8525) );
  INV_X1 U9975 ( .A(n8525), .ZN(n8643) );
  XNOR2_X1 U9976 ( .A(n8527), .B(n8526), .ZN(n8530) );
  OAI21_X1 U9977 ( .B1(n8530), .B2(n8529), .A(n8528), .ZN(n8639) );
  INV_X1 U9978 ( .A(n8561), .ZN(n8532) );
  AOI211_X1 U9979 ( .C1(n8641), .C2(n8532), .A(n9833), .B(n4618), .ZN(n8640)
         );
  NAND2_X1 U9980 ( .A1(n8640), .A2(n8533), .ZN(n8537) );
  AOI22_X1 U9981 ( .A1(n8535), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8534), .B2(
        n9756), .ZN(n8536) );
  OAI211_X1 U9982 ( .C1(n8025), .C2(n8538), .A(n8537), .B(n8536), .ZN(n8539)
         );
  AOI21_X1 U9983 ( .B1(n8639), .B2(n9768), .A(n8539), .ZN(n8540) );
  OAI21_X1 U9984 ( .B1(n8643), .B2(n8541), .A(n8540), .ZN(P2_U3279) );
  AND2_X1 U9985 ( .A1(n8543), .A2(n8542), .ZN(n8544) );
  XNOR2_X1 U9986 ( .A(n8547), .B(n8546), .ZN(n8553) );
  OAI22_X1 U9987 ( .A1(n8551), .A2(n8550), .B1(n8549), .B2(n8548), .ZN(n8552)
         );
  AOI21_X1 U9988 ( .B1(n8553), .B2(n9748), .A(n8552), .ZN(n8554) );
  OAI21_X1 U9989 ( .B1(n9441), .B2(n9797), .A(n8554), .ZN(n9444) );
  NAND2_X1 U9990 ( .A1(n9444), .A2(n8555), .ZN(n8568) );
  OAI22_X1 U9991 ( .A1(n8555), .A2(n8558), .B1(n8557), .B2(n8556), .ZN(n8564)
         );
  NOR2_X1 U9992 ( .A1(n8559), .A2(n9442), .ZN(n8560) );
  OR2_X1 U9993 ( .A1(n8561), .A2(n8560), .ZN(n9443) );
  NOR2_X1 U9994 ( .A1(n9443), .A2(n8562), .ZN(n8563) );
  AOI211_X1 U9995 ( .C1(n8566), .C2(n8565), .A(n8564), .B(n8563), .ZN(n8567)
         );
  OAI211_X1 U9996 ( .C1(n9441), .C2(n8569), .A(n8568), .B(n8567), .ZN(P2_U3280) );
  NAND2_X1 U9997 ( .A1(n8570), .A2(n9815), .ZN(n8571) );
  OAI211_X1 U9998 ( .C1(n8572), .C2(n9833), .A(n8571), .B(n8575), .ZN(n8657)
         );
  MUX2_X1 U9999 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8657), .S(n9853), .Z(
        P2_U3551) );
  NAND3_X1 U10000 ( .A1(n8574), .A2(n9816), .A3(n8573), .ZN(n8576) );
  OAI211_X1 U10001 ( .C1(n8577), .C2(n9831), .A(n8576), .B(n8575), .ZN(n8658)
         );
  MUX2_X1 U10002 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8658), .S(n9853), .Z(
        P2_U3550) );
  AOI22_X1 U10003 ( .A1(n8583), .A2(n9816), .B1(n9815), .B2(n8582), .ZN(n8584)
         );
  OAI211_X1 U10004 ( .C1(n8586), .C2(n8644), .A(n8585), .B(n8584), .ZN(n8660)
         );
  MUX2_X1 U10005 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8660), .S(n9853), .Z(
        P2_U3548) );
  AOI22_X1 U10006 ( .A1(n8588), .A2(n9816), .B1(n9815), .B2(n8587), .ZN(n8589)
         );
  OAI211_X1 U10007 ( .C1(n8591), .C2(n8644), .A(n8590), .B(n8589), .ZN(n8661)
         );
  MUX2_X1 U10008 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8661), .S(n9853), .Z(
        P2_U3547) );
  AOI21_X1 U10009 ( .B1(n9815), .B2(n8593), .A(n8592), .ZN(n8594) );
  OAI211_X1 U10010 ( .C1(n8596), .C2(n8644), .A(n8595), .B(n8594), .ZN(n8662)
         );
  MUX2_X1 U10011 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8662), .S(n9853), .Z(
        P2_U3546) );
  AOI211_X1 U10012 ( .C1(n9815), .C2(n8599), .A(n8598), .B(n8597), .ZN(n8600)
         );
  OAI21_X1 U10013 ( .B1(n8601), .B2(n8644), .A(n8600), .ZN(n8663) );
  MUX2_X1 U10014 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8663), .S(n9853), .Z(
        P2_U3545) );
  AOI22_X1 U10015 ( .A1(n8603), .A2(n9816), .B1(n9815), .B2(n8602), .ZN(n8604)
         );
  OAI211_X1 U10016 ( .C1(n8606), .C2(n8644), .A(n8605), .B(n8604), .ZN(n8664)
         );
  MUX2_X1 U10017 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8664), .S(n9853), .Z(
        P2_U3544) );
  NAND2_X1 U10018 ( .A1(n8607), .A2(n9837), .ZN(n8612) );
  AOI22_X1 U10019 ( .A1(n8609), .A2(n9816), .B1(n9815), .B2(n8608), .ZN(n8610)
         );
  OAI211_X1 U10020 ( .C1(n8433), .C2(n8612), .A(n8611), .B(n8610), .ZN(n8665)
         );
  MUX2_X1 U10021 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8665), .S(n9853), .Z(
        P2_U3543) );
  AOI22_X1 U10022 ( .A1(n8614), .A2(n9816), .B1(n9815), .B2(n8613), .ZN(n8615)
         );
  OAI211_X1 U10023 ( .C1(n8617), .C2(n8644), .A(n8616), .B(n8615), .ZN(n8666)
         );
  MUX2_X1 U10024 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8666), .S(n9853), .Z(
        P2_U3542) );
  INV_X1 U10025 ( .A(n8618), .ZN(n8622) );
  AOI22_X1 U10026 ( .A1(n8620), .A2(n9816), .B1(n9815), .B2(n8619), .ZN(n8621)
         );
  OAI211_X1 U10027 ( .C1(n8623), .C2(n8644), .A(n8622), .B(n8621), .ZN(n8667)
         );
  MUX2_X1 U10028 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8667), .S(n9853), .Z(
        P2_U3541) );
  AOI22_X1 U10029 ( .A1(n8625), .A2(n9816), .B1(n9815), .B2(n8624), .ZN(n8626)
         );
  OAI211_X1 U10030 ( .C1(n8628), .C2(n8644), .A(n8627), .B(n8626), .ZN(n8668)
         );
  MUX2_X1 U10031 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8668), .S(n9853), .Z(
        P2_U3540) );
  AOI211_X1 U10032 ( .C1(n9815), .C2(n8631), .A(n8630), .B(n8629), .ZN(n8632)
         );
  OAI21_X1 U10033 ( .B1(n8633), .B2(n8644), .A(n8632), .ZN(n8669) );
  MUX2_X1 U10034 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8669), .S(n9853), .Z(
        P2_U3539) );
  AOI22_X1 U10035 ( .A1(n8635), .A2(n9816), .B1(n9815), .B2(n8634), .ZN(n8636)
         );
  OAI211_X1 U10036 ( .C1(n8638), .C2(n8644), .A(n8637), .B(n8636), .ZN(n8670)
         );
  MUX2_X1 U10037 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8670), .S(n9853), .Z(
        P2_U3538) );
  AOI211_X1 U10038 ( .C1(n9815), .C2(n8641), .A(n8640), .B(n8639), .ZN(n8642)
         );
  OAI21_X1 U10039 ( .B1(n8644), .B2(n8643), .A(n8642), .ZN(n8671) );
  MUX2_X1 U10040 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8671), .S(n9853), .Z(
        P2_U3537) );
  OAI22_X1 U10041 ( .A1(n8646), .A2(n9833), .B1(n8645), .B2(n9831), .ZN(n8648)
         );
  AOI211_X1 U10042 ( .C1(n9837), .C2(n8649), .A(n8648), .B(n8647), .ZN(n8672)
         );
  MUX2_X1 U10043 ( .A(n6107), .B(n8672), .S(n9853), .Z(n8650) );
  INV_X1 U10044 ( .A(n8650), .ZN(P2_U3535) );
  OAI22_X1 U10045 ( .A1(n8652), .A2(n9833), .B1(n8651), .B2(n9831), .ZN(n8653)
         );
  AOI21_X1 U10046 ( .B1(n8654), .B2(n9829), .A(n8653), .ZN(n8655) );
  NAND2_X1 U10047 ( .A1(n8656), .A2(n8655), .ZN(n8674) );
  INV_X1 U10048 ( .A(n9853), .ZN(n9850) );
  MUX2_X1 U10049 ( .A(n8674), .B(P2_REG1_REG_13__SCAN_IN), .S(n9850), .Z(
        P2_U3533) );
  MUX2_X1 U10050 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8657), .S(n4405), .Z(
        P2_U3519) );
  MUX2_X1 U10051 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8658), .S(n4405), .Z(
        P2_U3518) );
  MUX2_X1 U10052 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8660), .S(n4405), .Z(
        P2_U3516) );
  MUX2_X1 U10053 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8661), .S(n4405), .Z(
        P2_U3515) );
  MUX2_X1 U10054 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8662), .S(n4405), .Z(
        P2_U3514) );
  MUX2_X1 U10055 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8663), .S(n4405), .Z(
        P2_U3513) );
  MUX2_X1 U10056 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8664), .S(n4405), .Z(
        P2_U3512) );
  MUX2_X1 U10057 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8665), .S(n4405), .Z(
        P2_U3511) );
  MUX2_X1 U10058 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8666), .S(n4405), .Z(
        P2_U3510) );
  MUX2_X1 U10059 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8667), .S(n4405), .Z(
        P2_U3509) );
  MUX2_X1 U10060 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8668), .S(n4405), .Z(
        P2_U3508) );
  MUX2_X1 U10061 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8669), .S(n4405), .Z(
        P2_U3507) );
  MUX2_X1 U10062 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8670), .S(n4405), .Z(
        P2_U3505) );
  MUX2_X1 U10063 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8671), .S(n4405), .Z(
        P2_U3502) );
  INV_X1 U10064 ( .A(n8672), .ZN(n8673) );
  MUX2_X1 U10065 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8673), .S(n4405), .Z(
        P2_U3496) );
  MUX2_X1 U10066 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8674), .S(n4405), .Z(
        P2_U3490) );
  NAND3_X1 U10067 ( .A1(n8676), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8677) );
  OAI22_X1 U10068 ( .A1(n8675), .A2(n8677), .B1(n6119), .B2(n7404), .ZN(n8678)
         );
  AOI21_X1 U10069 ( .B1(n9363), .B2(n8679), .A(n8678), .ZN(n8680) );
  INV_X1 U10070 ( .A(n8680), .ZN(P2_U3327) );
  INV_X1 U10071 ( .A(n8681), .ZN(n9374) );
  OAI222_X1 U10072 ( .A1(n8131), .A2(n9374), .B1(P2_U3152), .B2(n8683), .C1(
        n8682), .C2(n7404), .ZN(P2_U3329) );
  MUX2_X1 U10073 ( .A(n8684), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NOR2_X1 U10074 ( .A1(n4472), .A2(n4421), .ZN(n8686) );
  XNOR2_X1 U10075 ( .A(n8686), .B(n8685), .ZN(n8691) );
  INV_X1 U10076 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8687) );
  OAI22_X1 U10077 ( .A1(n8816), .A2(n9130), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8687), .ZN(n8689) );
  OAI22_X1 U10078 ( .A1(n8831), .A2(n9097), .B1(n9074), .B2(n8830), .ZN(n8688)
         );
  AOI211_X1 U10079 ( .C1(n9310), .C2(n8819), .A(n8689), .B(n8688), .ZN(n8690)
         );
  OAI21_X1 U10080 ( .B1(n8691), .B2(n8825), .A(n8690), .ZN(P1_U3214) );
  XNOR2_X1 U10081 ( .A(n8693), .B(n8692), .ZN(n8694) );
  XNOR2_X1 U10082 ( .A(n8775), .B(n8694), .ZN(n8695) );
  NAND2_X1 U10083 ( .A1(n8695), .A2(n8812), .ZN(n8704) );
  INV_X1 U10084 ( .A(n8696), .ZN(n8697) );
  AOI21_X1 U10085 ( .B1(n8833), .B2(n8841), .A(n8697), .ZN(n8703) );
  INV_X1 U10086 ( .A(n8698), .ZN(n8699) );
  AOI22_X1 U10087 ( .A1(n8807), .A2(n8839), .B1(n8806), .B2(n8699), .ZN(n8702)
         );
  NAND2_X1 U10088 ( .A1(n8819), .A2(n8700), .ZN(n8701) );
  NAND4_X1 U10089 ( .A1(n8704), .A2(n8703), .A3(n8702), .A4(n8701), .ZN(
        P1_U3215) );
  NAND2_X1 U10090 ( .A1(n4486), .A2(n8705), .ZN(n8706) );
  XNOR2_X1 U10091 ( .A(n8707), .B(n8706), .ZN(n8711) );
  NAND2_X1 U10092 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8932) );
  OAI21_X1 U10093 ( .B1(n9129), .B2(n8830), .A(n8932), .ZN(n8709) );
  OAI22_X1 U10094 ( .A1(n8831), .A2(n9155), .B1(n9200), .B2(n8816), .ZN(n8708)
         );
  AOI211_X1 U10095 ( .C1(n9330), .C2(n8819), .A(n8709), .B(n8708), .ZN(n8710)
         );
  OAI21_X1 U10096 ( .B1(n8711), .B2(n8825), .A(n8710), .ZN(P1_U3217) );
  NAND2_X1 U10097 ( .A1(n5008), .A2(n8712), .ZN(n8713) );
  XOR2_X1 U10098 ( .A(n8714), .B(n8713), .Z(n8715) );
  NAND2_X1 U10099 ( .A1(n8715), .A2(n8812), .ZN(n8721) );
  AND2_X1 U10100 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9594) );
  AOI21_X1 U10101 ( .B1(n8833), .B2(n8843), .A(n9594), .ZN(n8720) );
  INV_X1 U10102 ( .A(n8716), .ZN(n8717) );
  AOI22_X1 U10103 ( .A1(n8807), .A2(n8841), .B1(n8806), .B2(n8717), .ZN(n8719)
         );
  NAND2_X1 U10104 ( .A1(n8819), .A2(n4403), .ZN(n8718) );
  NAND4_X1 U10105 ( .A1(n8721), .A2(n8720), .A3(n8719), .A4(n8718), .ZN(
        P1_U3219) );
  XOR2_X1 U10106 ( .A(n8723), .B(n8722), .Z(n8728) );
  OAI22_X1 U10107 ( .A1(n8830), .A2(n9130), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8724), .ZN(n8726) );
  OAI22_X1 U10108 ( .A1(n8831), .A2(n9132), .B1(n9129), .B2(n8816), .ZN(n8725)
         );
  AOI211_X1 U10109 ( .C1(n9322), .C2(n8819), .A(n8726), .B(n8725), .ZN(n8727)
         );
  OAI21_X1 U10110 ( .B1(n8728), .B2(n8825), .A(n8727), .ZN(P1_U3221) );
  XOR2_X1 U10111 ( .A(n8730), .B(n8729), .Z(n8735) );
  OAI22_X1 U10112 ( .A1(n8830), .A2(n9076), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8731), .ZN(n8733) );
  OAI22_X1 U10113 ( .A1(n8831), .A2(n9068), .B1(n9074), .B2(n8816), .ZN(n8732)
         );
  AOI211_X1 U10114 ( .C1(n9302), .C2(n8819), .A(n8733), .B(n8732), .ZN(n8734)
         );
  OAI21_X1 U10115 ( .B1(n8735), .B2(n8825), .A(n8734), .ZN(P1_U3223) );
  XOR2_X1 U10116 ( .A(n8737), .B(n8736), .Z(n8738) );
  XNOR2_X1 U10117 ( .A(n8739), .B(n8738), .ZN(n8743) );
  NAND2_X1 U10118 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9644) );
  OAI21_X1 U10119 ( .B1(n8816), .B2(n9208), .A(n9644), .ZN(n8741) );
  OAI22_X1 U10120 ( .A1(n8831), .A2(n9215), .B1(n8953), .B2(n8830), .ZN(n8740)
         );
  AOI211_X1 U10121 ( .C1(n9220), .C2(n8819), .A(n8741), .B(n8740), .ZN(n8742)
         );
  OAI21_X1 U10122 ( .B1(n8743), .B2(n8825), .A(n8742), .ZN(P1_U3224) );
  XOR2_X1 U10123 ( .A(n8745), .B(n8744), .Z(n8749) );
  NAND2_X1 U10124 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9664) );
  OAI21_X1 U10125 ( .B1(n8816), .B2(n9198), .A(n9664), .ZN(n8747) );
  OAI22_X1 U10126 ( .A1(n8831), .A2(n9190), .B1(n9200), .B2(n8830), .ZN(n8746)
         );
  AOI211_X1 U10127 ( .C1(n9342), .C2(n8819), .A(n8747), .B(n8746), .ZN(n8748)
         );
  OAI21_X1 U10128 ( .B1(n8749), .B2(n8825), .A(n8748), .ZN(P1_U3226) );
  OAI21_X1 U10129 ( .B1(n8752), .B2(n8751), .A(n8750), .ZN(n8753) );
  NAND2_X1 U10130 ( .A1(n8753), .A2(n8812), .ZN(n8757) );
  INV_X1 U10131 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9997) );
  OAI22_X1 U10132 ( .A1(n8830), .A2(n9083), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9997), .ZN(n8755) );
  OAI22_X1 U10133 ( .A1(n8831), .A2(n9086), .B1(n9121), .B2(n8816), .ZN(n8754)
         );
  AOI211_X1 U10134 ( .C1(n9307), .C2(n8819), .A(n8755), .B(n8754), .ZN(n8756)
         );
  NAND2_X1 U10135 ( .A1(n8757), .A2(n8756), .ZN(P1_U3227) );
  AOI21_X1 U10136 ( .B1(n8759), .B2(n8758), .A(n4449), .ZN(n8764) );
  INV_X1 U10137 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8760) );
  OAI22_X1 U10138 ( .A1(n8830), .A2(n9119), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8760), .ZN(n8762) );
  OAI22_X1 U10139 ( .A1(n8831), .A2(n9143), .B1(n8955), .B2(n8816), .ZN(n8761)
         );
  AOI211_X1 U10140 ( .C1(n9325), .C2(n8819), .A(n8762), .B(n8761), .ZN(n8763)
         );
  OAI21_X1 U10141 ( .B1(n8764), .B2(n8825), .A(n8763), .ZN(P1_U3231) );
  NOR2_X1 U10142 ( .A1(n8766), .A2(n4775), .ZN(n8768) );
  XNOR2_X1 U10143 ( .A(n8768), .B(n8767), .ZN(n8773) );
  OAI22_X1 U10144 ( .A1(n8816), .A2(n9119), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8769), .ZN(n8771) );
  OAI22_X1 U10145 ( .A1(n8831), .A2(n9113), .B1(n9121), .B2(n8830), .ZN(n8770)
         );
  AOI211_X1 U10146 ( .C1(n9317), .C2(n8819), .A(n8771), .B(n8770), .ZN(n8772)
         );
  OAI21_X1 U10147 ( .B1(n8773), .B2(n8825), .A(n8772), .ZN(P1_U3233) );
  OR2_X1 U10148 ( .A1(n8775), .A2(n8774), .ZN(n8777) );
  NAND2_X1 U10149 ( .A1(n8777), .A2(n8776), .ZN(n8778) );
  XOR2_X1 U10150 ( .A(n8779), .B(n8778), .Z(n8780) );
  NAND2_X1 U10151 ( .A1(n8780), .A2(n8812), .ZN(n8787) );
  AOI21_X1 U10152 ( .B1(n8807), .B2(n8838), .A(n8781), .ZN(n8786) );
  INV_X1 U10153 ( .A(n9477), .ZN(n8782) );
  AOI22_X1 U10154 ( .A1(n8833), .A2(n8840), .B1(n8806), .B2(n8782), .ZN(n8785)
         );
  NAND2_X1 U10155 ( .A1(n8819), .A2(n8783), .ZN(n8784) );
  NAND4_X1 U10156 ( .A1(n8787), .A2(n8786), .A3(n8785), .A4(n8784), .ZN(
        P1_U3234) );
  INV_X1 U10157 ( .A(n8788), .ZN(n8789) );
  NOR2_X1 U10158 ( .A1(n8790), .A2(n8789), .ZN(n8792) );
  XNOR2_X1 U10159 ( .A(n8792), .B(n8791), .ZN(n8796) );
  NAND2_X1 U10160 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8896) );
  OAI21_X1 U10161 ( .B1(n8830), .B2(n8955), .A(n8896), .ZN(n8794) );
  OAI22_X1 U10162 ( .A1(n8831), .A2(n9171), .B1(n8953), .B2(n8816), .ZN(n8793)
         );
  AOI211_X1 U10163 ( .C1(n9335), .C2(n8819), .A(n8794), .B(n8793), .ZN(n8795)
         );
  OAI21_X1 U10164 ( .B1(n8796), .B2(n8825), .A(n8795), .ZN(P1_U3236) );
  OAI21_X1 U10165 ( .B1(n8799), .B2(n8798), .A(n8797), .ZN(n8803) );
  XNOR2_X1 U10166 ( .A(n8801), .B(n8800), .ZN(n8802) );
  XNOR2_X1 U10167 ( .A(n8803), .B(n8802), .ZN(n8804) );
  NAND2_X1 U10168 ( .A1(n8804), .A2(n8812), .ZN(n8811) );
  AND2_X1 U10169 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9576) );
  AOI21_X1 U10170 ( .B1(n8833), .B2(n8845), .A(n9576), .ZN(n8810) );
  AOI22_X1 U10171 ( .A1(n8807), .A2(n8843), .B1(n8806), .B2(n8805), .ZN(n8809)
         );
  NAND2_X1 U10172 ( .A1(n8819), .A2(n9696), .ZN(n8808) );
  NAND4_X1 U10173 ( .A1(n8811), .A2(n8810), .A3(n8809), .A4(n8808), .ZN(
        P1_U3237) );
  OAI211_X1 U10174 ( .C1(n8815), .C2(n8814), .A(n8813), .B(n8812), .ZN(n8821)
         );
  OAI22_X1 U10175 ( .A1(n8830), .A2(n9053), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9965), .ZN(n8818) );
  OAI22_X1 U10176 ( .A1(n8831), .A2(n9056), .B1(n9083), .B2(n8816), .ZN(n8817)
         );
  AOI211_X1 U10177 ( .C1(n9297), .C2(n8819), .A(n8818), .B(n8817), .ZN(n8820)
         );
  NAND2_X1 U10178 ( .A1(n8821), .A2(n8820), .ZN(P1_U3238) );
  INV_X1 U10179 ( .A(n9242), .ZN(n9488) );
  INV_X1 U10180 ( .A(n8824), .ZN(n8829) );
  AOI21_X1 U10181 ( .B1(n8822), .B2(n8824), .A(n8823), .ZN(n8826) );
  NOR2_X1 U10182 ( .A1(n8826), .A2(n8825), .ZN(n8827) );
  OAI21_X1 U10183 ( .B1(n8829), .B2(n8828), .A(n8827), .ZN(n8835) );
  AND2_X1 U10184 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9637) );
  OAI22_X1 U10185 ( .A1(n8831), .A2(n9235), .B1(n9198), .B2(n8830), .ZN(n8832)
         );
  AOI211_X1 U10186 ( .C1(n8833), .C2(n9229), .A(n9637), .B(n8832), .ZN(n8834)
         );
  OAI211_X1 U10187 ( .C1(n9488), .C2(n8836), .A(n8835), .B(n8834), .ZN(
        P1_U3239) );
  MUX2_X1 U10188 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n8999), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10189 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n8966), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10190 ( .A(n9044), .B(P1_DATAO_REG_26__SCAN_IN), .S(n8846), .Z(
        P1_U3581) );
  MUX2_X1 U10191 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n8962), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10192 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9106), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10193 ( .A(n8837), .B(P1_DATAO_REG_23__SCAN_IN), .S(n8846), .Z(
        P1_U3578) );
  MUX2_X1 U10194 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9107), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10195 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9142), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10196 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9163), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10197 ( .A(n9181), .B(P1_DATAO_REG_19__SCAN_IN), .S(n8846), .Z(
        P1_U3574) );
  MUX2_X1 U10198 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9162), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10199 ( .A(n9206), .B(P1_DATAO_REG_17__SCAN_IN), .S(n8846), .Z(
        P1_U3572) );
  MUX2_X1 U10200 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9230), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10201 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9255), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10202 ( .A(n9229), .B(P1_DATAO_REG_14__SCAN_IN), .S(n8846), .Z(
        P1_U3569) );
  MUX2_X1 U10203 ( .A(n9252), .B(P1_DATAO_REG_13__SCAN_IN), .S(n8846), .Z(
        P1_U3568) );
  MUX2_X1 U10204 ( .A(n8838), .B(P1_DATAO_REG_12__SCAN_IN), .S(n8846), .Z(
        P1_U3567) );
  MUX2_X1 U10205 ( .A(n8839), .B(P1_DATAO_REG_11__SCAN_IN), .S(n8846), .Z(
        P1_U3566) );
  MUX2_X1 U10206 ( .A(n8840), .B(P1_DATAO_REG_10__SCAN_IN), .S(n8846), .Z(
        P1_U3565) );
  MUX2_X1 U10207 ( .A(n8841), .B(P1_DATAO_REG_9__SCAN_IN), .S(n8846), .Z(
        P1_U3564) );
  MUX2_X1 U10208 ( .A(n8842), .B(P1_DATAO_REG_8__SCAN_IN), .S(n8846), .Z(
        P1_U3563) );
  MUX2_X1 U10209 ( .A(n8843), .B(P1_DATAO_REG_7__SCAN_IN), .S(n8846), .Z(
        P1_U3562) );
  MUX2_X1 U10210 ( .A(n8844), .B(P1_DATAO_REG_6__SCAN_IN), .S(n8846), .Z(
        P1_U3561) );
  MUX2_X1 U10211 ( .A(n8845), .B(P1_DATAO_REG_5__SCAN_IN), .S(n8846), .Z(
        P1_U3560) );
  MUX2_X1 U10212 ( .A(n8847), .B(P1_DATAO_REG_4__SCAN_IN), .S(n8846), .Z(
        P1_U3559) );
  MUX2_X1 U10213 ( .A(n8848), .B(P1_DATAO_REG_3__SCAN_IN), .S(n8846), .Z(
        P1_U3558) );
  MUX2_X1 U10214 ( .A(n6679), .B(P1_DATAO_REG_2__SCAN_IN), .S(n8846), .Z(
        P1_U3557) );
  MUX2_X1 U10215 ( .A(n6625), .B(P1_DATAO_REG_1__SCAN_IN), .S(n8846), .Z(
        P1_U3556) );
  NAND2_X1 U10216 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n8853) );
  INV_X1 U10217 ( .A(n8849), .ZN(n8852) );
  INV_X1 U10218 ( .A(n8850), .ZN(n8851) );
  AOI211_X1 U10219 ( .C1(n8853), .C2(n8852), .A(n8851), .B(n9630), .ZN(n8854)
         );
  AOI21_X1 U10220 ( .B1(n9651), .B2(n8855), .A(n8854), .ZN(n8861) );
  AOI22_X1 U10221 ( .A1(n9581), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3084), .ZN(n8860) );
  OAI211_X1 U10222 ( .C1(n8858), .C2(n8857), .A(n9663), .B(n8856), .ZN(n8859)
         );
  NAND3_X1 U10223 ( .A1(n8861), .A2(n8860), .A3(n8859), .ZN(P1_U3242) );
  OAI211_X1 U10224 ( .C1(n8864), .C2(n8863), .A(n9670), .B(n8862), .ZN(n8873)
         );
  AOI21_X1 U10225 ( .B1(n9581), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n8865), .ZN(
        n8872) );
  NAND2_X1 U10226 ( .A1(n9651), .A2(n8866), .ZN(n8871) );
  OAI211_X1 U10227 ( .C1(n8869), .C2(n8868), .A(n9663), .B(n8867), .ZN(n8870)
         );
  NAND4_X1 U10228 ( .A1(n8873), .A2(n8872), .A3(n8871), .A4(n8870), .ZN(
        P1_U3244) );
  OAI21_X1 U10229 ( .B1(n8876), .B2(n8875), .A(n8874), .ZN(n8877) );
  AOI22_X1 U10230 ( .A1(n8878), .A2(n9651), .B1(n9670), .B2(n8877), .ZN(n8887)
         );
  INV_X1 U10231 ( .A(n8879), .ZN(n8880) );
  AOI21_X1 U10232 ( .B1(n9581), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n8880), .ZN(
        n8886) );
  OAI21_X1 U10233 ( .B1(n8883), .B2(n8882), .A(n8881), .ZN(n8884) );
  NAND2_X1 U10234 ( .A1(n9663), .A2(n8884), .ZN(n8885) );
  NAND3_X1 U10235 ( .A1(n8887), .A2(n8886), .A3(n8885), .ZN(P1_U3248) );
  AOI22_X1 U10236 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n8921), .B1(n8918), .B2(
        n8922), .ZN(n8895) );
  XNOR2_X1 U10237 ( .A(n9667), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9672) );
  INV_X1 U10238 ( .A(n9652), .ZN(n8892) );
  MUX2_X1 U10239 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n8888), .S(n9652), .Z(n9654) );
  AOI21_X1 U10240 ( .B1(n8900), .B2(n9498), .A(n8889), .ZN(n8890) );
  NAND2_X1 U10241 ( .A1(n9638), .A2(n8890), .ZN(n8891) );
  XNOR2_X1 U10242 ( .A(n8890), .B(n8904), .ZN(n9640) );
  NAND2_X1 U10243 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9640), .ZN(n9639) );
  NAND2_X1 U10244 ( .A1(n8891), .A2(n9639), .ZN(n9655) );
  NAND2_X1 U10245 ( .A1(n9654), .A2(n9655), .ZN(n9653) );
  OAI21_X1 U10246 ( .B1(n8892), .B2(n8888), .A(n9653), .ZN(n9671) );
  NAND2_X1 U10247 ( .A1(n9672), .A2(n9671), .ZN(n9669) );
  OAI21_X1 U10248 ( .B1(n9667), .B2(n8893), .A(n9669), .ZN(n8894) );
  NOR2_X1 U10249 ( .A1(n8895), .A2(n8894), .ZN(n8920) );
  AOI21_X1 U10250 ( .B1(n8895), .B2(n8894), .A(n8920), .ZN(n8916) );
  INV_X1 U10251 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n8897) );
  OAI21_X1 U10252 ( .B1(n9675), .B2(n8897), .A(n8896), .ZN(n8914) );
  NOR2_X1 U10253 ( .A1(n8918), .A2(n8898), .ZN(n8899) );
  AOI21_X1 U10254 ( .B1(n8918), .B2(n8898), .A(n8899), .ZN(n8912) );
  NAND2_X1 U10255 ( .A1(n8901), .A2(n8900), .ZN(n8903) );
  NAND2_X1 U10256 ( .A1(n8903), .A2(n8902), .ZN(n8905) );
  NOR2_X1 U10257 ( .A1(n8904), .A2(n8905), .ZN(n8906) );
  XNOR2_X1 U10258 ( .A(n8905), .B(n8904), .ZN(n9635) );
  NOR2_X1 U10259 ( .A1(n9236), .A2(n9635), .ZN(n9634) );
  INV_X1 U10260 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n10116) );
  NOR2_X1 U10261 ( .A1(n9652), .A2(n10116), .ZN(n8907) );
  AOI21_X1 U10262 ( .B1(n10116), .B2(n9652), .A(n8907), .ZN(n9647) );
  NOR2_X1 U10263 ( .A1(n9648), .A2(n9647), .ZN(n9646) );
  AOI21_X1 U10264 ( .B1(n9652), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9646), .ZN(
        n9660) );
  OR2_X1 U10265 ( .A1(n9667), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8909) );
  NAND2_X1 U10266 ( .A1(n9667), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8908) );
  AND2_X1 U10267 ( .A1(n8909), .A2(n8908), .ZN(n9661) );
  NOR2_X1 U10268 ( .A1(n9660), .A2(n9661), .ZN(n9659) );
  NOR2_X1 U10269 ( .A1(n8911), .A2(n8912), .ZN(n8917) );
  AOI211_X1 U10270 ( .C1(n8912), .C2(n8911), .A(n8917), .B(n9645), .ZN(n8913)
         );
  AOI211_X1 U10271 ( .C1(n9651), .C2(n8918), .A(n8914), .B(n8913), .ZN(n8915)
         );
  OAI21_X1 U10272 ( .B1(n8916), .B2(n9630), .A(n8915), .ZN(P1_U3259) );
  AOI21_X1 U10273 ( .B1(n8918), .B2(P1_REG2_REG_18__SCAN_IN), .A(n8917), .ZN(
        n8919) );
  XNOR2_X1 U10274 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n8919), .ZN(n8928) );
  INV_X1 U10275 ( .A(n8928), .ZN(n8926) );
  AOI21_X1 U10276 ( .B1(n8922), .B2(n8921), .A(n8920), .ZN(n8923) );
  XNOR2_X1 U10277 ( .A(n8924), .B(n8923), .ZN(n8927) );
  OAI21_X1 U10278 ( .B1(n8927), .B2(n9630), .A(n9666), .ZN(n8925) );
  AOI21_X1 U10279 ( .B1(n9663), .B2(n8926), .A(n8925), .ZN(n8931) );
  AOI22_X1 U10280 ( .A1(n8928), .A2(n9663), .B1(n8927), .B2(n9670), .ZN(n8930)
         );
  MUX2_X1 U10281 ( .A(n8931), .B(n8930), .S(n8929), .Z(n8933) );
  OAI211_X1 U10282 ( .C1(n8934), .C2(n9675), .A(n8933), .B(n8932), .ZN(
        P1_U3260) );
  INV_X1 U10283 ( .A(n9265), .ZN(n9494) );
  INV_X1 U10284 ( .A(n9330), .ZN(n9158) );
  NAND2_X1 U10285 ( .A1(n9111), .A2(n9100), .ZN(n9094) );
  NAND2_X1 U10286 ( .A1(n8942), .A2(n9001), .ZN(n8935) );
  XNOR2_X1 U10287 ( .A(n7485), .B(n8935), .ZN(n9274) );
  AND2_X1 U10288 ( .A1(n8936), .A2(P1_B_REG_SCAN_IN), .ZN(n8937) );
  NOR2_X1 U10289 ( .A1(n9467), .A2(n8937), .ZN(n8998) );
  NAND2_X1 U10290 ( .A1(n8938), .A2(n8998), .ZN(n9277) );
  NOR2_X1 U10291 ( .A1(n9223), .A2(n9277), .ZN(n8944) );
  NOR2_X1 U10292 ( .A1(n8939), .A2(n9475), .ZN(n8940) );
  AOI211_X1 U10293 ( .C1(n9223), .C2(P1_REG2_REG_31__SCAN_IN), .A(n8944), .B(
        n8940), .ZN(n8941) );
  OAI21_X1 U10294 ( .B1(n9274), .B2(n9239), .A(n8941), .ZN(P1_U3261) );
  XNOR2_X1 U10295 ( .A(n8942), .B(n9001), .ZN(n9278) );
  NOR2_X1 U10296 ( .A1(n8942), .A2(n9475), .ZN(n8943) );
  AOI211_X1 U10297 ( .C1(n9223), .C2(P1_REG2_REG_30__SCAN_IN), .A(n8944), .B(
        n8943), .ZN(n8945) );
  OAI21_X1 U10298 ( .B1(n9278), .B2(n9239), .A(n8945), .ZN(P1_U3262) );
  OR2_X1 U10299 ( .A1(n9499), .A2(n9252), .ZN(n8946) );
  NAND2_X1 U10300 ( .A1(n9499), .A2(n9252), .ZN(n8948) );
  NAND2_X1 U10301 ( .A1(n8949), .A2(n8948), .ZN(n9247) );
  INV_X1 U10302 ( .A(n9247), .ZN(n8950) );
  OR2_X1 U10303 ( .A1(n9265), .A2(n9229), .ZN(n8951) );
  NAND2_X1 U10304 ( .A1(n8952), .A2(n8951), .ZN(n9224) );
  NOR2_X1 U10305 ( .A1(n9224), .A2(n9227), .ZN(n9226) );
  NOR2_X1 U10306 ( .A1(n9342), .A2(n9206), .ZN(n8954) );
  INV_X1 U10307 ( .A(n9342), .ZN(n9189) );
  NAND2_X1 U10308 ( .A1(n9330), .A2(n9181), .ZN(n8956) );
  AOI22_X1 U10309 ( .A1(n9151), .A2(n8956), .B1(n9158), .B2(n8955), .ZN(n9138)
         );
  NOR2_X1 U10310 ( .A1(n9297), .A2(n9044), .ZN(n8964) );
  NAND2_X1 U10311 ( .A1(n9036), .A2(n9053), .ZN(n9016) );
  AND2_X1 U10312 ( .A1(n9016), .A2(n9011), .ZN(n8965) );
  NAND2_X1 U10313 ( .A1(n9017), .A2(n8965), .ZN(n9021) );
  INV_X1 U10314 ( .A(n9285), .ZN(n9026) );
  NAND2_X1 U10315 ( .A1(n9285), .A2(n8966), .ZN(n8967) );
  NAND2_X1 U10316 ( .A1(n9021), .A2(n8967), .ZN(n8968) );
  XNOR2_X1 U10317 ( .A(n8968), .B(n8995), .ZN(n9279) );
  INV_X1 U10318 ( .A(n9279), .ZN(n9009) );
  NAND2_X1 U10319 ( .A1(n8970), .A2(n8969), .ZN(n8972) );
  NAND2_X1 U10320 ( .A1(n8972), .A2(n8971), .ZN(n9249) );
  INV_X1 U10321 ( .A(n8974), .ZN(n8975) );
  NAND2_X1 U10322 ( .A1(n9160), .A2(n9161), .ZN(n9159) );
  NAND2_X1 U10323 ( .A1(n9159), .A2(n8980), .ZN(n9139) );
  OAI21_X1 U10324 ( .B1(n9080), .B2(n9081), .A(n8987), .ZN(n9073) );
  INV_X1 U10325 ( .A(n9072), .ZN(n8990) );
  INV_X1 U10326 ( .A(n8988), .ZN(n8989) );
  INV_X1 U10327 ( .A(n8993), .ZN(n8994) );
  NOR2_X1 U10328 ( .A1(n9010), .A2(n8994), .ZN(n8997) );
  INV_X1 U10329 ( .A(n8995), .ZN(n8996) );
  AOI22_X1 U10330 ( .A1(n9253), .A2(n8966), .B1(n8999), .B2(n8998), .ZN(n9000)
         );
  INV_X1 U10331 ( .A(n9282), .ZN(n9006) );
  NAND2_X1 U10332 ( .A1(n9281), .A2(n9193), .ZN(n9005) );
  INV_X1 U10333 ( .A(n9002), .ZN(n9003) );
  AOI22_X1 U10334 ( .A1(n9223), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9003), .B2(
        n9172), .ZN(n9004) );
  OAI211_X1 U10335 ( .C1(n9006), .C2(n9475), .A(n9005), .B(n9004), .ZN(n9007)
         );
  AOI21_X1 U10336 ( .B1(n9280), .B2(n9269), .A(n9007), .ZN(n9008) );
  OAI21_X1 U10337 ( .B1(n9009), .B2(n9271), .A(n9008), .ZN(P1_U3355) );
  AOI211_X1 U10338 ( .C1(n9012), .C2(n9011), .A(n9234), .B(n9010), .ZN(n9015)
         );
  OAI22_X1 U10339 ( .A1(n9013), .A2(n9467), .B1(n9053), .B2(n9465), .ZN(n9014)
         );
  NOR2_X1 U10340 ( .A1(n9015), .A2(n9014), .ZN(n9288) );
  NAND2_X1 U10341 ( .A1(n9017), .A2(n9016), .ZN(n9019) );
  NAND2_X1 U10342 ( .A1(n9019), .A2(n9018), .ZN(n9020) );
  NAND2_X1 U10343 ( .A1(n9284), .A2(n9214), .ZN(n9029) );
  AOI21_X1 U10344 ( .B1(n9285), .B2(n9032), .A(n4648), .ZN(n9286) );
  INV_X1 U10345 ( .A(n9023), .ZN(n9024) );
  AOI22_X1 U10346 ( .A1(n9223), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9024), .B2(
        n9172), .ZN(n9025) );
  OAI21_X1 U10347 ( .B1(n9026), .B2(n9475), .A(n9025), .ZN(n9027) );
  AOI21_X1 U10348 ( .B1(n9286), .B2(n9461), .A(n9027), .ZN(n9028) );
  OAI211_X1 U10349 ( .C1(n9223), .C2(n9288), .A(n9029), .B(n9028), .ZN(
        P1_U3263) );
  XNOR2_X1 U10350 ( .A(n9031), .B(n9030), .ZN(n9294) );
  INV_X1 U10351 ( .A(n9054), .ZN(n9033) );
  AOI211_X1 U10352 ( .C1(n9291), .C2(n9033), .A(n9723), .B(n4649), .ZN(n9290)
         );
  AOI22_X1 U10353 ( .A1(n9223), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9034), .B2(
        n9172), .ZN(n9035) );
  OAI21_X1 U10354 ( .B1(n9036), .B2(n9475), .A(n9035), .ZN(n9046) );
  NOR2_X1 U10355 ( .A1(n9037), .A2(n9467), .ZN(n9043) );
  AOI21_X1 U10356 ( .B1(n4701), .B2(n9039), .A(n9038), .ZN(n9040) );
  NOR3_X1 U10357 ( .A1(n9041), .A2(n9040), .A3(n9234), .ZN(n9042) );
  AOI211_X1 U10358 ( .C1(n9253), .C2(n9044), .A(n9043), .B(n9042), .ZN(n9293)
         );
  NOR2_X1 U10359 ( .A1(n9293), .A2(n9223), .ZN(n9045) );
  AOI211_X1 U10360 ( .C1(n9193), .C2(n9290), .A(n9046), .B(n9045), .ZN(n9047)
         );
  OAI21_X1 U10361 ( .B1(n9294), .B2(n9271), .A(n9047), .ZN(P1_U3264) );
  XOR2_X1 U10362 ( .A(n9050), .B(n9048), .Z(n9299) );
  AOI21_X1 U10363 ( .B1(n9051), .B2(n9050), .A(n9049), .ZN(n9052) );
  OAI222_X1 U10364 ( .A1(n9467), .A2(n9053), .B1(n9465), .B2(n9083), .C1(n9234), .C2(n9052), .ZN(n9295) );
  INV_X1 U10365 ( .A(n9066), .ZN(n9055) );
  AOI211_X1 U10366 ( .C1(n9297), .C2(n9055), .A(n9723), .B(n9054), .ZN(n9296)
         );
  NAND2_X1 U10367 ( .A1(n9296), .A2(n9193), .ZN(n9059) );
  INV_X1 U10368 ( .A(n9056), .ZN(n9057) );
  AOI22_X1 U10369 ( .A1(n9223), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9057), .B2(
        n9172), .ZN(n9058) );
  OAI211_X1 U10370 ( .C1(n9060), .C2(n9475), .A(n9059), .B(n9058), .ZN(n9061)
         );
  AOI21_X1 U10371 ( .B1(n9295), .B2(n9269), .A(n9061), .ZN(n9062) );
  OAI21_X1 U10372 ( .B1(n9299), .B2(n9271), .A(n9062), .ZN(P1_U3265) );
  OAI21_X1 U10373 ( .B1(n9064), .B2(n9072), .A(n9063), .ZN(n9065) );
  INV_X1 U10374 ( .A(n9065), .ZN(n9304) );
  AOI211_X1 U10375 ( .C1(n9302), .C2(n9084), .A(n9723), .B(n9066), .ZN(n9301)
         );
  INV_X1 U10376 ( .A(n9302), .ZN(n9067) );
  NOR2_X1 U10377 ( .A1(n9067), .A2(n9475), .ZN(n9071) );
  OAI22_X1 U10378 ( .A1(n9479), .A2(n9069), .B1(n9068), .B2(n9476), .ZN(n9070)
         );
  AOI211_X1 U10379 ( .C1(n9301), .C2(n9193), .A(n9071), .B(n9070), .ZN(n9078)
         );
  XNOR2_X1 U10380 ( .A(n9073), .B(n9072), .ZN(n9075) );
  OAI222_X1 U10381 ( .A1(n9467), .A2(n9076), .B1(n9075), .B2(n9234), .C1(n9465), .C2(n9074), .ZN(n9300) );
  NAND2_X1 U10382 ( .A1(n9300), .A2(n9269), .ZN(n9077) );
  OAI211_X1 U10383 ( .C1(n9304), .C2(n9271), .A(n9078), .B(n9077), .ZN(
        P1_U3266) );
  XNOR2_X1 U10384 ( .A(n9079), .B(n9081), .ZN(n9309) );
  AOI22_X1 U10385 ( .A1(n9307), .A2(n9264), .B1(n9223), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n9091) );
  XOR2_X1 U10386 ( .A(n9081), .B(n9080), .Z(n9082) );
  OAI222_X1 U10387 ( .A1(n9467), .A2(n9083), .B1(n9082), .B2(n9234), .C1(n9465), .C2(n9121), .ZN(n9305) );
  INV_X1 U10388 ( .A(n9084), .ZN(n9085) );
  AOI211_X1 U10389 ( .C1(n9307), .C2(n9094), .A(n9723), .B(n9085), .ZN(n9306)
         );
  INV_X1 U10390 ( .A(n9306), .ZN(n9088) );
  OAI22_X1 U10391 ( .A1(n9088), .A2(n9087), .B1(n9476), .B2(n9086), .ZN(n9089)
         );
  OAI21_X1 U10392 ( .B1(n9305), .B2(n9089), .A(n9269), .ZN(n9090) );
  OAI211_X1 U10393 ( .C1(n9309), .C2(n9271), .A(n9091), .B(n9090), .ZN(
        P1_U3267) );
  XNOR2_X1 U10394 ( .A(n9093), .B(n9092), .ZN(n9314) );
  INV_X1 U10395 ( .A(n9111), .ZN(n9096) );
  INV_X1 U10396 ( .A(n9094), .ZN(n9095) );
  AOI21_X1 U10397 ( .B1(n9310), .B2(n9096), .A(n9095), .ZN(n9311) );
  INV_X1 U10398 ( .A(n9097), .ZN(n9098) );
  AOI22_X1 U10399 ( .A1(n9223), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9098), .B2(
        n9172), .ZN(n9099) );
  OAI21_X1 U10400 ( .B1(n9100), .B2(n9475), .A(n9099), .ZN(n9109) );
  NAND2_X1 U10401 ( .A1(n9102), .A2(n9101), .ZN(n9104) );
  XNOR2_X1 U10402 ( .A(n9104), .B(n9103), .ZN(n9105) );
  AOI222_X1 U10403 ( .A1(n9107), .A2(n9253), .B1(n9106), .B2(n9254), .C1(n9470), .C2(n9105), .ZN(n9313) );
  NOR2_X1 U10404 ( .A1(n9313), .A2(n9223), .ZN(n9108) );
  AOI211_X1 U10405 ( .C1(n9311), .C2(n9461), .A(n9109), .B(n9108), .ZN(n9110)
         );
  OAI21_X1 U10406 ( .B1(n9314), .B2(n9271), .A(n9110), .ZN(P1_U3268) );
  XNOR2_X1 U10407 ( .A(n4437), .B(n9117), .ZN(n9319) );
  AOI211_X1 U10408 ( .C1(n9317), .C2(n4639), .A(n9723), .B(n9111), .ZN(n9316)
         );
  NOR2_X1 U10409 ( .A1(n9112), .A2(n9475), .ZN(n9116) );
  OAI22_X1 U10410 ( .A1(n9479), .A2(n9114), .B1(n9113), .B2(n9476), .ZN(n9115)
         );
  AOI211_X1 U10411 ( .C1(n9316), .C2(n9193), .A(n9116), .B(n9115), .ZN(n9123)
         );
  XNOR2_X1 U10412 ( .A(n9118), .B(n9117), .ZN(n9120) );
  OAI222_X1 U10413 ( .A1(n9467), .A2(n9121), .B1(n9120), .B2(n9234), .C1(n9465), .C2(n9119), .ZN(n9315) );
  NAND2_X1 U10414 ( .A1(n9315), .A2(n9269), .ZN(n9122) );
  OAI211_X1 U10415 ( .C1(n9319), .C2(n9271), .A(n9123), .B(n9122), .ZN(
        P1_U3269) );
  XNOR2_X1 U10416 ( .A(n9124), .B(n9127), .ZN(n9324) );
  AOI21_X1 U10417 ( .B1(n9127), .B2(n9126), .A(n9125), .ZN(n9128) );
  OAI222_X1 U10418 ( .A1(n9467), .A2(n9130), .B1(n9465), .B2(n9129), .C1(n9234), .C2(n9128), .ZN(n9320) );
  AOI211_X1 U10419 ( .C1(n9322), .C2(n9145), .A(n9723), .B(n9131), .ZN(n9321)
         );
  NAND2_X1 U10420 ( .A1(n9321), .A2(n9193), .ZN(n9135) );
  INV_X1 U10421 ( .A(n9132), .ZN(n9133) );
  AOI22_X1 U10422 ( .A1(n9223), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9133), .B2(
        n9172), .ZN(n9134) );
  OAI211_X1 U10423 ( .C1(n4637), .C2(n9475), .A(n9135), .B(n9134), .ZN(n9136)
         );
  AOI21_X1 U10424 ( .B1(n9320), .B2(n9479), .A(n9136), .ZN(n9137) );
  OAI21_X1 U10425 ( .B1(n9324), .B2(n9271), .A(n9137), .ZN(P1_U3270) );
  XNOR2_X1 U10426 ( .A(n9138), .B(n9140), .ZN(n9329) );
  XOR2_X1 U10427 ( .A(n9140), .B(n9139), .Z(n9141) );
  AOI222_X1 U10428 ( .A1(n9181), .A2(n9253), .B1(n9142), .B2(n9254), .C1(n9470), .C2(n9141), .ZN(n9328) );
  OAI21_X1 U10429 ( .B1(n9143), .B2(n9476), .A(n9328), .ZN(n9149) );
  NAND2_X1 U10430 ( .A1(n9152), .A2(n9325), .ZN(n9144) );
  AND2_X1 U10431 ( .A1(n9145), .A2(n9144), .ZN(n9326) );
  INV_X1 U10432 ( .A(n9326), .ZN(n9147) );
  AOI22_X1 U10433 ( .A1(n9325), .A2(n9264), .B1(n9223), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9146) );
  OAI21_X1 U10434 ( .B1(n9147), .B2(n9239), .A(n9146), .ZN(n9148) );
  AOI21_X1 U10435 ( .B1(n9149), .B2(n9479), .A(n9148), .ZN(n9150) );
  OAI21_X1 U10436 ( .B1(n9329), .B2(n9271), .A(n9150), .ZN(P1_U3271) );
  XNOR2_X1 U10437 ( .A(n9151), .B(n9161), .ZN(n9334) );
  INV_X1 U10438 ( .A(n9170), .ZN(n9154) );
  INV_X1 U10439 ( .A(n9152), .ZN(n9153) );
  AOI21_X1 U10440 ( .B1(n9330), .B2(n9154), .A(n9153), .ZN(n9331) );
  INV_X1 U10441 ( .A(n9155), .ZN(n9156) );
  AOI22_X1 U10442 ( .A1(n9223), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9156), .B2(
        n9172), .ZN(n9157) );
  OAI21_X1 U10443 ( .B1(n9158), .B2(n9475), .A(n9157), .ZN(n9166) );
  OAI21_X1 U10444 ( .B1(n9161), .B2(n9160), .A(n9159), .ZN(n9164) );
  AOI222_X1 U10445 ( .A1(n9470), .A2(n9164), .B1(n9163), .B2(n9254), .C1(n9162), .C2(n9253), .ZN(n9333) );
  NOR2_X1 U10446 ( .A1(n9333), .A2(n9223), .ZN(n9165) );
  AOI211_X1 U10447 ( .C1(n9331), .C2(n9461), .A(n9166), .B(n9165), .ZN(n9167)
         );
  OAI21_X1 U10448 ( .B1(n9334), .B2(n9271), .A(n9167), .ZN(P1_U3272) );
  XNOR2_X1 U10449 ( .A(n9169), .B(n9168), .ZN(n9339) );
  AOI21_X1 U10450 ( .B1(n9335), .B2(n9187), .A(n9170), .ZN(n9336) );
  INV_X1 U10451 ( .A(n9335), .ZN(n9175) );
  INV_X1 U10452 ( .A(n9171), .ZN(n9173) );
  AOI22_X1 U10453 ( .A1(n9223), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9173), .B2(
        n9172), .ZN(n9174) );
  OAI21_X1 U10454 ( .B1(n9175), .B2(n9475), .A(n9174), .ZN(n9184) );
  INV_X1 U10455 ( .A(n9176), .ZN(n9177) );
  NOR2_X1 U10456 ( .A1(n9178), .A2(n9177), .ZN(n9180) );
  XNOR2_X1 U10457 ( .A(n9180), .B(n9179), .ZN(n9182) );
  AOI222_X1 U10458 ( .A1(n9470), .A2(n9182), .B1(n9181), .B2(n9254), .C1(n9206), .C2(n9253), .ZN(n9338) );
  NOR2_X1 U10459 ( .A1(n9338), .A2(n9223), .ZN(n9183) );
  AOI211_X1 U10460 ( .C1(n9336), .C2(n9461), .A(n9184), .B(n9183), .ZN(n9185)
         );
  OAI21_X1 U10461 ( .B1(n9339), .B2(n9271), .A(n9185), .ZN(P1_U3273) );
  XNOR2_X1 U10462 ( .A(n9186), .B(n9196), .ZN(n9344) );
  INV_X1 U10463 ( .A(n9187), .ZN(n9188) );
  AOI211_X1 U10464 ( .C1(n9342), .C2(n9216), .A(n9723), .B(n9188), .ZN(n9341)
         );
  NOR2_X1 U10465 ( .A1(n9189), .A2(n9475), .ZN(n9192) );
  INV_X1 U10466 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10089) );
  OAI22_X1 U10467 ( .A1(n9479), .A2(n10089), .B1(n9190), .B2(n9476), .ZN(n9191) );
  AOI211_X1 U10468 ( .C1(n9341), .C2(n9193), .A(n9192), .B(n9191), .ZN(n9202)
         );
  INV_X1 U10469 ( .A(n9194), .ZN(n9195) );
  NOR2_X1 U10470 ( .A1(n9205), .A2(n9195), .ZN(n9197) );
  XNOR2_X1 U10471 ( .A(n9197), .B(n9196), .ZN(n9199) );
  OAI222_X1 U10472 ( .A1(n9467), .A2(n9200), .B1(n9199), .B2(n9234), .C1(n9465), .C2(n9198), .ZN(n9340) );
  NAND2_X1 U10473 ( .A1(n9340), .A2(n9269), .ZN(n9201) );
  OAI211_X1 U10474 ( .C1(n9344), .C2(n9271), .A(n9202), .B(n9201), .ZN(
        P1_U3274) );
  NOR2_X1 U10475 ( .A1(n9203), .A2(n9212), .ZN(n9204) );
  OR2_X1 U10476 ( .A1(n9205), .A2(n9204), .ZN(n9210) );
  NAND2_X1 U10477 ( .A1(n9206), .A2(n9254), .ZN(n9207) );
  OAI21_X1 U10478 ( .B1(n9208), .B2(n9465), .A(n9207), .ZN(n9209) );
  AOI21_X1 U10479 ( .B1(n9210), .B2(n9470), .A(n9209), .ZN(n9485) );
  AOI21_X1 U10480 ( .B1(n9213), .B2(n9212), .A(n9211), .ZN(n9487) );
  NAND2_X1 U10481 ( .A1(n9487), .A2(n9214), .ZN(n9222) );
  OAI22_X1 U10482 ( .A1(n9479), .A2(n10116), .B1(n9215), .B2(n9476), .ZN(n9219) );
  INV_X1 U10483 ( .A(n9238), .ZN(n9217) );
  OAI211_X1 U10484 ( .C1(n9217), .C2(n4646), .A(n9711), .B(n9216), .ZN(n9484)
         );
  NOR2_X1 U10485 ( .A1(n9484), .A2(n9267), .ZN(n9218) );
  AOI211_X1 U10486 ( .C1(n9264), .C2(n9220), .A(n9219), .B(n9218), .ZN(n9221)
         );
  OAI211_X1 U10487 ( .C1(n9223), .C2(n9485), .A(n9222), .B(n9221), .ZN(
        P1_U3275) );
  AND2_X1 U10488 ( .A1(n9224), .A2(n9227), .ZN(n9225) );
  NOR2_X1 U10489 ( .A1(n9226), .A2(n9225), .ZN(n9492) );
  INV_X1 U10490 ( .A(n9492), .ZN(n9246) );
  XNOR2_X1 U10491 ( .A(n9228), .B(n9227), .ZN(n9233) );
  NAND2_X1 U10492 ( .A1(n9492), .A2(n9719), .ZN(n9232) );
  AOI22_X1 U10493 ( .A1(n9230), .A2(n9254), .B1(n9253), .B2(n9229), .ZN(n9231)
         );
  OAI211_X1 U10494 ( .C1(n9234), .C2(n9233), .A(n9232), .B(n9231), .ZN(n9490)
         );
  NAND2_X1 U10495 ( .A1(n9490), .A2(n9269), .ZN(n9244) );
  OAI22_X1 U10496 ( .A1(n9479), .A2(n9236), .B1(n9235), .B2(n9476), .ZN(n9241)
         );
  OR2_X1 U10497 ( .A1(n9258), .A2(n9488), .ZN(n9237) );
  NAND2_X1 U10498 ( .A1(n9238), .A2(n9237), .ZN(n9489) );
  NOR2_X1 U10499 ( .A1(n9489), .A2(n9239), .ZN(n9240) );
  AOI211_X1 U10500 ( .C1(n9264), .C2(n9242), .A(n9241), .B(n9240), .ZN(n9243)
         );
  OAI211_X1 U10501 ( .C1(n9246), .C2(n9245), .A(n9244), .B(n9243), .ZN(
        P1_U3276) );
  XOR2_X1 U10502 ( .A(n9247), .B(n9248), .Z(n9497) );
  INV_X1 U10503 ( .A(n9497), .ZN(n9272) );
  NAND2_X1 U10504 ( .A1(n9249), .A2(n9248), .ZN(n9250) );
  NAND3_X1 U10505 ( .A1(n9251), .A2(n9470), .A3(n9250), .ZN(n9257) );
  AOI22_X1 U10506 ( .A1(n9255), .A2(n9254), .B1(n9253), .B2(n9252), .ZN(n9256)
         );
  NAND2_X1 U10507 ( .A1(n9257), .A2(n9256), .ZN(n9496) );
  INV_X1 U10508 ( .A(n9258), .ZN(n9259) );
  OAI211_X1 U10509 ( .C1(n9494), .C2(n9260), .A(n9259), .B(n9711), .ZN(n9493)
         );
  OAI22_X1 U10510 ( .A1(n9479), .A2(n9262), .B1(n9261), .B2(n9476), .ZN(n9263)
         );
  AOI21_X1 U10511 ( .B1(n9265), .B2(n9264), .A(n9263), .ZN(n9266) );
  OAI21_X1 U10512 ( .B1(n9493), .B2(n9267), .A(n9266), .ZN(n9268) );
  AOI21_X1 U10513 ( .B1(n9496), .B2(n9269), .A(n9268), .ZN(n9270) );
  OAI21_X1 U10514 ( .B1(n9272), .B2(n9271), .A(n9270), .ZN(P1_U3277) );
  NAND2_X1 U10515 ( .A1(n7485), .A2(n9709), .ZN(n9273) );
  OAI211_X1 U10516 ( .C1(n9274), .C2(n9723), .A(n9273), .B(n9277), .ZN(n9346)
         );
  MUX2_X1 U10517 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9346), .S(n9737), .Z(
        P1_U3554) );
  NAND2_X1 U10518 ( .A1(n9275), .A2(n9709), .ZN(n9276) );
  OAI211_X1 U10519 ( .C1(n9278), .C2(n9723), .A(n9277), .B(n9276), .ZN(n9347)
         );
  MUX2_X1 U10520 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9347), .S(n9737), .Z(
        P1_U3553) );
  NAND2_X1 U10521 ( .A1(n9279), .A2(n9725), .ZN(n9283) );
  MUX2_X1 U10522 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9348), .S(n9737), .Z(
        P1_U3552) );
  NAND2_X1 U10523 ( .A1(n9284), .A2(n9725), .ZN(n9289) );
  AOI22_X1 U10524 ( .A1(n9286), .A2(n9711), .B1(n9285), .B2(n9709), .ZN(n9287)
         );
  NAND3_X1 U10525 ( .A1(n9289), .A2(n9288), .A3(n9287), .ZN(n9349) );
  MUX2_X1 U10526 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9349), .S(n9737), .Z(
        P1_U3551) );
  AOI21_X1 U10527 ( .B1(n9291), .B2(n9709), .A(n9290), .ZN(n9292) );
  OAI211_X1 U10528 ( .C1(n9294), .C2(n9687), .A(n9293), .B(n9292), .ZN(n9350)
         );
  MUX2_X1 U10529 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9350), .S(n9737), .Z(
        P1_U3550) );
  AOI211_X1 U10530 ( .C1(n9297), .C2(n9709), .A(n9296), .B(n9295), .ZN(n9298)
         );
  OAI21_X1 U10531 ( .B1(n9299), .B2(n9687), .A(n9298), .ZN(n9351) );
  MUX2_X1 U10532 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9351), .S(n9737), .Z(
        P1_U3549) );
  AOI211_X1 U10533 ( .C1(n9302), .C2(n9709), .A(n9301), .B(n9300), .ZN(n9303)
         );
  OAI21_X1 U10534 ( .B1(n9304), .B2(n9687), .A(n9303), .ZN(n9352) );
  MUX2_X1 U10535 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9352), .S(n9737), .Z(
        P1_U3548) );
  AOI211_X1 U10536 ( .C1(n9307), .C2(n9709), .A(n9306), .B(n9305), .ZN(n9308)
         );
  OAI21_X1 U10537 ( .B1(n9309), .B2(n9687), .A(n9308), .ZN(n9353) );
  MUX2_X1 U10538 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9353), .S(n9737), .Z(
        P1_U3547) );
  AOI22_X1 U10539 ( .A1(n9311), .A2(n9711), .B1(n9310), .B2(n9709), .ZN(n9312)
         );
  OAI211_X1 U10540 ( .C1(n9314), .C2(n9687), .A(n9313), .B(n9312), .ZN(n9354)
         );
  MUX2_X1 U10541 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9354), .S(n9737), .Z(
        P1_U3546) );
  AOI211_X1 U10542 ( .C1(n9317), .C2(n9709), .A(n9316), .B(n9315), .ZN(n9318)
         );
  OAI21_X1 U10543 ( .B1(n9319), .B2(n9687), .A(n9318), .ZN(n9355) );
  MUX2_X1 U10544 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9355), .S(n9737), .Z(
        P1_U3545) );
  AOI211_X1 U10545 ( .C1(n9322), .C2(n9709), .A(n9321), .B(n9320), .ZN(n9323)
         );
  OAI21_X1 U10546 ( .B1(n9324), .B2(n9687), .A(n9323), .ZN(n9356) );
  MUX2_X1 U10547 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9356), .S(n9737), .Z(
        P1_U3544) );
  AOI22_X1 U10548 ( .A1(n9326), .A2(n9711), .B1(n9325), .B2(n9709), .ZN(n9327)
         );
  OAI211_X1 U10549 ( .C1(n9329), .C2(n9687), .A(n9328), .B(n9327), .ZN(n9357)
         );
  MUX2_X1 U10550 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9357), .S(n9737), .Z(
        P1_U3543) );
  AOI22_X1 U10551 ( .A1(n9331), .A2(n9711), .B1(n9330), .B2(n9709), .ZN(n9332)
         );
  OAI211_X1 U10552 ( .C1(n9334), .C2(n9687), .A(n9333), .B(n9332), .ZN(n9358)
         );
  MUX2_X1 U10553 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9358), .S(n9737), .Z(
        P1_U3542) );
  AOI22_X1 U10554 ( .A1(n9336), .A2(n9711), .B1(n9335), .B2(n9709), .ZN(n9337)
         );
  OAI211_X1 U10555 ( .C1(n9339), .C2(n9687), .A(n9338), .B(n9337), .ZN(n9359)
         );
  MUX2_X1 U10556 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9359), .S(n9737), .Z(
        P1_U3541) );
  AOI211_X1 U10557 ( .C1(n9342), .C2(n9709), .A(n9341), .B(n9340), .ZN(n9343)
         );
  OAI21_X1 U10558 ( .B1(n9344), .B2(n9687), .A(n9343), .ZN(n9360) );
  MUX2_X1 U10559 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9360), .S(n9737), .Z(
        P1_U3540) );
  MUX2_X1 U10560 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9345), .S(n9737), .Z(
        P1_U3525) );
  MUX2_X1 U10561 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9346), .S(n9729), .Z(
        P1_U3522) );
  MUX2_X1 U10562 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9347), .S(n9729), .Z(
        P1_U3521) );
  MUX2_X1 U10563 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9348), .S(n9729), .Z(
        P1_U3520) );
  MUX2_X1 U10564 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9349), .S(n9729), .Z(
        P1_U3519) );
  MUX2_X1 U10565 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9350), .S(n9729), .Z(
        P1_U3518) );
  MUX2_X1 U10566 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9351), .S(n9729), .Z(
        P1_U3517) );
  MUX2_X1 U10567 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9352), .S(n9729), .Z(
        P1_U3516) );
  MUX2_X1 U10568 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9353), .S(n9729), .Z(
        P1_U3515) );
  MUX2_X1 U10569 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9354), .S(n9729), .Z(
        P1_U3514) );
  MUX2_X1 U10570 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9355), .S(n9729), .Z(
        P1_U3513) );
  MUX2_X1 U10571 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9356), .S(n9729), .Z(
        P1_U3512) );
  MUX2_X1 U10572 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9357), .S(n9729), .Z(
        P1_U3511) );
  MUX2_X1 U10573 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9358), .S(n9729), .Z(
        P1_U3510) );
  MUX2_X1 U10574 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9359), .S(n9729), .Z(
        P1_U3508) );
  MUX2_X1 U10575 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9360), .S(n9729), .Z(
        P1_U3505) );
  MUX2_X1 U10576 ( .A(P1_D_REG_1__SCAN_IN), .B(n9361), .S(n9678), .Z(P1_U3441)
         );
  MUX2_X1 U10577 ( .A(P1_D_REG_0__SCAN_IN), .B(n9362), .S(n9678), .Z(P1_U3440)
         );
  INV_X1 U10578 ( .A(n9363), .ZN(n9370) );
  NOR4_X1 U10579 ( .A1(n9365), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n5464), .ZN(n9366) );
  AOI21_X1 U10580 ( .B1(n9367), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9366), .ZN(
        n9368) );
  OAI21_X1 U10581 ( .B1(n9370), .B2(n9369), .A(n9368), .ZN(P1_U3322) );
  OAI222_X1 U10582 ( .A1(n9369), .A2(n9374), .B1(n9373), .B2(P1_U3084), .C1(
        n9372), .C2(n9371), .ZN(P1_U3324) );
  MUX2_X1 U10583 ( .A(n9375), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI21_X1 U10584 ( .B1(n9739), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n9376), .ZN(
        n9388) );
  AOI211_X1 U10585 ( .C1(n9379), .C2(n9378), .A(n9377), .B(n9740), .ZN(n9380)
         );
  AOI21_X1 U10586 ( .B1(n9395), .B2(n9381), .A(n9380), .ZN(n9387) );
  INV_X1 U10587 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9382) );
  NOR2_X1 U10588 ( .A1(n9382), .A2(n5897), .ZN(n9385) );
  OAI211_X1 U10589 ( .C1(n9385), .C2(n9384), .A(n9891), .B(n9383), .ZN(n9386)
         );
  NAND3_X1 U10590 ( .A1(n9388), .A2(n9387), .A3(n9386), .ZN(P2_U3246) );
  AOI21_X1 U10591 ( .B1(n9739), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n9389), .ZN(
        n9401) );
  AOI211_X1 U10592 ( .C1(n9392), .C2(n9391), .A(n9390), .B(n9740), .ZN(n9393)
         );
  AOI21_X1 U10593 ( .B1(n9395), .B2(n9394), .A(n9393), .ZN(n9400) );
  OAI211_X1 U10594 ( .C1(n9398), .C2(n9397), .A(n9891), .B(n9396), .ZN(n9399)
         );
  NAND3_X1 U10595 ( .A1(n9401), .A2(n9400), .A3(n9399), .ZN(P2_U3247) );
  INV_X1 U10596 ( .A(n9402), .ZN(n9407) );
  OAI21_X1 U10597 ( .B1(n9404), .B2(n9705), .A(n9403), .ZN(n9406) );
  AOI211_X1 U10598 ( .C1(n9686), .C2(n9407), .A(n9406), .B(n9405), .ZN(n9408)
         );
  INV_X1 U10599 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10105) );
  AOI22_X1 U10600 ( .A1(n9729), .A2(n9408), .B1(n10105), .B2(n9727), .ZN(
        P1_U3484) );
  AOI22_X1 U10601 ( .A1(n9737), .A2(n9408), .B1(n5400), .B2(n9735), .ZN(
        P1_U3533) );
  NOR2_X1 U10602 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9409) );
  AOI21_X1 U10603 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9409), .ZN(n9860) );
  NOR2_X1 U10604 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9410) );
  AOI21_X1 U10605 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9410), .ZN(n9863) );
  NOR2_X1 U10606 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9411) );
  AOI21_X1 U10607 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9411), .ZN(n9866) );
  NOR2_X1 U10608 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9412) );
  AOI21_X1 U10609 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9412), .ZN(n9869) );
  NOR2_X1 U10610 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9413) );
  AOI21_X1 U10611 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9413), .ZN(n9872) );
  NOR2_X1 U10612 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9421) );
  XNOR2_X1 U10613 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10227) );
  NAND2_X1 U10614 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9419) );
  INV_X1 U10615 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9414) );
  XOR2_X1 U10616 ( .A(n9414), .B(n9994), .Z(n10225) );
  NAND2_X1 U10617 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9417) );
  XOR2_X1 U10618 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10221) );
  AOI21_X1 U10619 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9854) );
  INV_X1 U10620 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9415) );
  NAND3_X1 U10621 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9856) );
  OAI21_X1 U10622 ( .B1(n9854), .B2(n9415), .A(n9856), .ZN(n10220) );
  NAND2_X1 U10623 ( .A1(n10221), .A2(n10220), .ZN(n9416) );
  NAND2_X1 U10624 ( .A1(n9417), .A2(n9416), .ZN(n10224) );
  NAND2_X1 U10625 ( .A1(n10225), .A2(n10224), .ZN(n9418) );
  NAND2_X1 U10626 ( .A1(n9419), .A2(n9418), .ZN(n10226) );
  NOR2_X1 U10627 ( .A1(n10227), .A2(n10226), .ZN(n9420) );
  NOR2_X1 U10628 ( .A1(n9421), .A2(n9420), .ZN(n9422) );
  NOR2_X1 U10629 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9422), .ZN(n10215) );
  AND2_X1 U10630 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9422), .ZN(n10214) );
  NOR2_X1 U10631 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10214), .ZN(n9423) );
  NOR2_X1 U10632 ( .A1(n10215), .A2(n9423), .ZN(n9424) );
  NAND2_X1 U10633 ( .A1(n9424), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9426) );
  XOR2_X1 U10634 ( .A(n9424), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10213) );
  NAND2_X1 U10635 ( .A1(n10213), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9425) );
  NAND2_X1 U10636 ( .A1(n9426), .A2(n9425), .ZN(n9427) );
  NAND2_X1 U10637 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9427), .ZN(n9429) );
  XOR2_X1 U10638 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9427), .Z(n10208) );
  NAND2_X1 U10639 ( .A1(n10208), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n9428) );
  NAND2_X1 U10640 ( .A1(n9429), .A2(n9428), .ZN(n9430) );
  NAND2_X1 U10641 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n9430), .ZN(n9432) );
  XOR2_X1 U10642 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n9430), .Z(n10223) );
  NAND2_X1 U10643 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n10223), .ZN(n9431) );
  NAND2_X1 U10644 ( .A1(n9432), .A2(n9431), .ZN(n9433) );
  AND2_X1 U10645 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9433), .ZN(n9434) );
  XNOR2_X1 U10646 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9433), .ZN(n10211) );
  INV_X1 U10647 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10210) );
  NAND2_X1 U10648 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9435) );
  OAI21_X1 U10649 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9435), .ZN(n9880) );
  NAND2_X1 U10650 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9436) );
  OAI21_X1 U10651 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9436), .ZN(n9877) );
  AOI21_X1 U10652 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9876), .ZN(n9875) );
  NOR2_X1 U10653 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9437) );
  AOI21_X1 U10654 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9437), .ZN(n9874) );
  NAND2_X1 U10655 ( .A1(n9875), .A2(n9874), .ZN(n9873) );
  OAI21_X1 U10656 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9873), .ZN(n9871) );
  NAND2_X1 U10657 ( .A1(n9872), .A2(n9871), .ZN(n9870) );
  OAI21_X1 U10658 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9870), .ZN(n9868) );
  NAND2_X1 U10659 ( .A1(n9869), .A2(n9868), .ZN(n9867) );
  OAI21_X1 U10660 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9867), .ZN(n9865) );
  NAND2_X1 U10661 ( .A1(n9866), .A2(n9865), .ZN(n9864) );
  OAI21_X1 U10662 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9864), .ZN(n9862) );
  NAND2_X1 U10663 ( .A1(n9863), .A2(n9862), .ZN(n9861) );
  OAI21_X1 U10664 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9861), .ZN(n9859) );
  NAND2_X1 U10665 ( .A1(n9860), .A2(n9859), .ZN(n9858) );
  OAI21_X1 U10666 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9858), .ZN(n10218) );
  NOR2_X1 U10667 ( .A1(n8312), .A2(n10218), .ZN(n9438) );
  NAND2_X1 U10668 ( .A1(n8312), .A2(n10218), .ZN(n10217) );
  OAI21_X1 U10669 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9438), .A(n10217), .ZN(
        n9440) );
  XOR2_X1 U10670 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .Z(n9439) );
  XNOR2_X1 U10671 ( .A(n9440), .B(n9439), .ZN(ADD_1071_U4) );
  INV_X1 U10672 ( .A(n9441), .ZN(n9446) );
  OAI22_X1 U10673 ( .A1(n9443), .A2(n9833), .B1(n9442), .B2(n9831), .ZN(n9445)
         );
  AOI211_X1 U10674 ( .C1(n9829), .C2(n9446), .A(n9445), .B(n9444), .ZN(n9454)
         );
  AOI22_X1 U10675 ( .A1(n9853), .A2(n9454), .B1(n10074), .B2(n9850), .ZN(
        P2_U3536) );
  OAI211_X1 U10676 ( .C1(n9449), .C2(n9831), .A(n9448), .B(n9447), .ZN(n9450)
         );
  AOI21_X1 U10677 ( .B1(n9451), .B2(n9837), .A(n9450), .ZN(n9456) );
  AOI22_X1 U10678 ( .A1(n9853), .A2(n9456), .B1(n9452), .B2(n9850), .ZN(
        P2_U3534) );
  INV_X1 U10679 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9453) );
  AOI22_X1 U10680 ( .A1(n4405), .A2(n9454), .B1(n9453), .B2(n9839), .ZN(
        P2_U3499) );
  INV_X1 U10681 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9455) );
  AOI22_X1 U10682 ( .A1(n4405), .A2(n9456), .B1(n9455), .B2(n9839), .ZN(
        P2_U3493) );
  XNOR2_X1 U10683 ( .A(n9457), .B(n9464), .ZN(n9474) );
  INV_X1 U10684 ( .A(n9474), .ZN(n9517) );
  OR2_X1 U10685 ( .A1(n9458), .A2(n9513), .ZN(n9459) );
  NAND2_X1 U10686 ( .A1(n4433), .A2(n9459), .ZN(n9514) );
  INV_X1 U10687 ( .A(n9514), .ZN(n9460) );
  AOI22_X1 U10688 ( .A1(n9517), .A2(n9462), .B1(n9461), .B2(n9460), .ZN(n9483)
         );
  XOR2_X1 U10689 ( .A(n9464), .B(n9463), .Z(n9471) );
  OAI22_X1 U10690 ( .A1(n9468), .A2(n9467), .B1(n9466), .B2(n9465), .ZN(n9469)
         );
  AOI21_X1 U10691 ( .B1(n9471), .B2(n9470), .A(n9469), .ZN(n9472) );
  OAI21_X1 U10692 ( .B1(n9474), .B2(n9473), .A(n9472), .ZN(n9515) );
  NOR2_X1 U10693 ( .A1(n9513), .A2(n9475), .ZN(n9481) );
  OAI22_X1 U10694 ( .A1(n9479), .A2(n9478), .B1(n9477), .B2(n9476), .ZN(n9480)
         );
  AOI211_X1 U10695 ( .C1(n9515), .C2(n9479), .A(n9481), .B(n9480), .ZN(n9482)
         );
  NAND2_X1 U10696 ( .A1(n9483), .A2(n9482), .ZN(P1_U3280) );
  OAI211_X1 U10697 ( .C1(n4646), .C2(n9705), .A(n9485), .B(n9484), .ZN(n9486)
         );
  AOI21_X1 U10698 ( .B1(n9487), .B2(n9725), .A(n9486), .ZN(n9519) );
  AOI22_X1 U10699 ( .A1(n9737), .A2(n9519), .B1(n8888), .B2(n9735), .ZN(
        P1_U3539) );
  OAI22_X1 U10700 ( .A1(n9489), .A2(n9723), .B1(n9488), .B2(n9705), .ZN(n9491)
         );
  AOI211_X1 U10701 ( .C1(n9686), .C2(n9492), .A(n9491), .B(n9490), .ZN(n9521)
         );
  AOI22_X1 U10702 ( .A1(n9737), .A2(n9521), .B1(n5513), .B2(n9735), .ZN(
        P1_U3538) );
  OAI21_X1 U10703 ( .B1(n9494), .B2(n9705), .A(n9493), .ZN(n9495) );
  AOI211_X1 U10704 ( .C1(n9497), .C2(n9725), .A(n9496), .B(n9495), .ZN(n9523)
         );
  AOI22_X1 U10705 ( .A1(n9737), .A2(n9523), .B1(n9498), .B2(n9735), .ZN(
        P1_U3537) );
  INV_X1 U10706 ( .A(n9499), .ZN(n9500) );
  OAI22_X1 U10707 ( .A1(n9501), .A2(n9723), .B1(n9500), .B2(n9705), .ZN(n9502)
         );
  AOI211_X1 U10708 ( .C1(n9504), .C2(n9725), .A(n9503), .B(n9502), .ZN(n9525)
         );
  AOI22_X1 U10709 ( .A1(n9737), .A2(n9525), .B1(n9505), .B2(n9735), .ZN(
        P1_U3536) );
  INV_X1 U10710 ( .A(n9510), .ZN(n9512) );
  AOI211_X1 U10711 ( .C1(n9508), .C2(n9709), .A(n9507), .B(n9506), .ZN(n9509)
         );
  OAI21_X1 U10712 ( .B1(n9715), .B2(n9510), .A(n9509), .ZN(n9511) );
  AOI21_X1 U10713 ( .B1(n9719), .B2(n9512), .A(n9511), .ZN(n9526) );
  AOI22_X1 U10714 ( .A1(n9737), .A2(n9526), .B1(n6389), .B2(n9735), .ZN(
        P1_U3535) );
  OAI22_X1 U10715 ( .A1(n9514), .A2(n9723), .B1(n9513), .B2(n9705), .ZN(n9516)
         );
  AOI211_X1 U10716 ( .C1(n9686), .C2(n9517), .A(n9516), .B(n9515), .ZN(n9527)
         );
  AOI22_X1 U10717 ( .A1(n9737), .A2(n9527), .B1(n6270), .B2(n9735), .ZN(
        P1_U3534) );
  INV_X1 U10718 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9518) );
  AOI22_X1 U10719 ( .A1(n9729), .A2(n9519), .B1(n9518), .B2(n9727), .ZN(
        P1_U3502) );
  INV_X1 U10720 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9520) );
  AOI22_X1 U10721 ( .A1(n9729), .A2(n9521), .B1(n9520), .B2(n9727), .ZN(
        P1_U3499) );
  INV_X1 U10722 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9522) );
  AOI22_X1 U10723 ( .A1(n9729), .A2(n9523), .B1(n9522), .B2(n9727), .ZN(
        P1_U3496) );
  INV_X1 U10724 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9524) );
  AOI22_X1 U10725 ( .A1(n9729), .A2(n9525), .B1(n9524), .B2(n9727), .ZN(
        P1_U3493) );
  AOI22_X1 U10726 ( .A1(n9729), .A2(n9526), .B1(n5448), .B2(n9727), .ZN(
        P1_U3490) );
  INV_X1 U10727 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U10728 ( .A1(n9729), .A2(n9527), .B1(n10176), .B2(n9727), .ZN(
        P1_U3487) );
  XNOR2_X1 U10729 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10730 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10731 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9538) );
  INV_X1 U10732 ( .A(n9528), .ZN(n9530) );
  AOI21_X1 U10733 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n9530), .A(n9529), .ZN(
        n9531) );
  AOI211_X1 U10734 ( .C1(n9533), .C2(P1_IR_REG_0__SCAN_IN), .A(n9532), .B(
        n9531), .ZN(n9536) );
  INV_X1 U10735 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9534) );
  NOR3_X1 U10736 ( .A1(n9630), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n9534), .ZN(
        n9535) );
  AOI211_X1 U10737 ( .C1(P1_ADDR_REG_0__SCAN_IN), .C2(n9581), .A(n9536), .B(
        n9535), .ZN(n9537) );
  OAI21_X1 U10738 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n9538), .A(n9537), .ZN(
        P1_U3241) );
  INV_X1 U10739 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9553) );
  AOI21_X1 U10740 ( .B1(n9541), .B2(n9540), .A(n9539), .ZN(n9543) );
  OAI21_X1 U10741 ( .B1(n9630), .B2(n9543), .A(n9542), .ZN(n9550) );
  AOI21_X1 U10742 ( .B1(n9546), .B2(n9545), .A(n9544), .ZN(n9548) );
  OAI22_X1 U10743 ( .A1(n9645), .A2(n9548), .B1(n9547), .B2(n9666), .ZN(n9549)
         );
  NOR3_X1 U10744 ( .A1(n9551), .A2(n9550), .A3(n9549), .ZN(n9552) );
  OAI21_X1 U10745 ( .B1(n9675), .B2(n9553), .A(n9552), .ZN(P1_U3245) );
  AND2_X1 U10746 ( .A1(n9555), .A2(n9554), .ZN(n9556) );
  NOR2_X1 U10747 ( .A1(n9557), .A2(n9556), .ZN(n9559) );
  AOI21_X1 U10748 ( .B1(n9670), .B2(n9559), .A(n9558), .ZN(n9565) );
  OAI21_X1 U10749 ( .B1(n9562), .B2(n9561), .A(n9560), .ZN(n9563) );
  NAND2_X1 U10750 ( .A1(n9663), .A2(n9563), .ZN(n9564) );
  AND2_X1 U10751 ( .A1(n9565), .A2(n9564), .ZN(n9568) );
  AOI22_X1 U10752 ( .A1(n9651), .A2(n9566), .B1(n9581), .B2(
        P1_ADDR_REG_5__SCAN_IN), .ZN(n9567) );
  NAND2_X1 U10753 ( .A1(n9568), .A2(n9567), .ZN(P1_U3246) );
  INV_X1 U10754 ( .A(n9569), .ZN(n9573) );
  INV_X1 U10755 ( .A(n9570), .ZN(n9572) );
  OAI211_X1 U10756 ( .C1(n9573), .C2(n9572), .A(n9663), .B(n9571), .ZN(n9579)
         );
  XNOR2_X1 U10757 ( .A(n9575), .B(n9574), .ZN(n9577) );
  AOI21_X1 U10758 ( .B1(n9670), .B2(n9577), .A(n9576), .ZN(n9578) );
  AND2_X1 U10759 ( .A1(n9579), .A2(n9578), .ZN(n9584) );
  INV_X1 U10760 ( .A(n9580), .ZN(n9582) );
  AOI22_X1 U10761 ( .A1(n9651), .A2(n9582), .B1(n9581), .B2(
        P1_ADDR_REG_6__SCAN_IN), .ZN(n9583) );
  NAND2_X1 U10762 ( .A1(n9584), .A2(n9583), .ZN(P1_U3247) );
  INV_X1 U10763 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10222) );
  INV_X1 U10764 ( .A(n9599), .ZN(n9586) );
  OAI21_X1 U10765 ( .B1(n9586), .B2(n9585), .A(n9613), .ZN(n9597) );
  MUX2_X1 U10766 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n6291), .S(n9587), .Z(n9590)
         );
  INV_X1 U10767 ( .A(n9588), .ZN(n9589) );
  NAND2_X1 U10768 ( .A1(n9590), .A2(n9589), .ZN(n9591) );
  NAND2_X1 U10769 ( .A1(n9592), .A2(n9591), .ZN(n9593) );
  NAND2_X1 U10770 ( .A1(n9663), .A2(n9593), .ZN(n9596) );
  INV_X1 U10771 ( .A(n9594), .ZN(n9595) );
  OAI211_X1 U10772 ( .C1(n9630), .C2(n9597), .A(n9596), .B(n9595), .ZN(n9598)
         );
  INV_X1 U10773 ( .A(n9598), .ZN(n9603) );
  NOR3_X1 U10774 ( .A1(n9630), .A2(n6266), .A3(n9599), .ZN(n9601) );
  OAI21_X1 U10775 ( .B1(n9601), .B2(n9651), .A(n9600), .ZN(n9602) );
  OAI211_X1 U10776 ( .C1(n10222), .C2(n9675), .A(n9603), .B(n9602), .ZN(
        P1_U3249) );
  INV_X1 U10777 ( .A(n9604), .ZN(n9608) );
  NAND2_X1 U10778 ( .A1(n9606), .A2(n9605), .ZN(n9607) );
  NAND3_X1 U10779 ( .A1(n9663), .A2(n9608), .A3(n9607), .ZN(n9610) );
  OAI211_X1 U10780 ( .C1(n9666), .C2(n9611), .A(n9610), .B(n9609), .ZN(n9612)
         );
  INV_X1 U10781 ( .A(n9612), .ZN(n9618) );
  NOR2_X1 U10782 ( .A1(n9614), .A2(n9613), .ZN(n9615) );
  OAI21_X1 U10783 ( .B1(n9616), .B2(n9615), .A(n9670), .ZN(n9617) );
  OAI211_X1 U10784 ( .C1(n10210), .C2(n9675), .A(n9618), .B(n9617), .ZN(
        P1_U3250) );
  INV_X1 U10785 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10175) );
  INV_X1 U10786 ( .A(n9619), .ZN(n9620) );
  OAI211_X1 U10787 ( .C1(n9622), .C2(n9621), .A(n9663), .B(n9620), .ZN(n9626)
         );
  AOI21_X1 U10788 ( .B1(n9651), .B2(n9624), .A(n9623), .ZN(n9625) );
  AND2_X1 U10789 ( .A1(n9626), .A2(n9625), .ZN(n9633) );
  AOI21_X1 U10790 ( .B1(n9629), .B2(n9628), .A(n9627), .ZN(n9631) );
  OR2_X1 U10791 ( .A1(n9631), .A2(n9630), .ZN(n9632) );
  OAI211_X1 U10792 ( .C1(n10175), .C2(n9675), .A(n9633), .B(n9632), .ZN(
        P1_U3253) );
  INV_X1 U10793 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9643) );
  AOI211_X1 U10794 ( .C1(n9635), .C2(n9236), .A(n9634), .B(n9645), .ZN(n9636)
         );
  AOI211_X1 U10795 ( .C1(n9651), .C2(n9638), .A(n9637), .B(n9636), .ZN(n9642)
         );
  OAI211_X1 U10796 ( .C1(n9640), .C2(P1_REG1_REG_15__SCAN_IN), .A(n9670), .B(
        n9639), .ZN(n9641) );
  OAI211_X1 U10797 ( .C1(n9643), .C2(n9675), .A(n9642), .B(n9641), .ZN(
        P1_U3256) );
  INV_X1 U10798 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9658) );
  INV_X1 U10799 ( .A(n9644), .ZN(n9650) );
  AOI211_X1 U10800 ( .C1(n9648), .C2(n9647), .A(n9646), .B(n9645), .ZN(n9649)
         );
  AOI211_X1 U10801 ( .C1(n9652), .C2(n9651), .A(n9650), .B(n9649), .ZN(n9657)
         );
  OAI211_X1 U10802 ( .C1(n9655), .C2(n9654), .A(n9670), .B(n9653), .ZN(n9656)
         );
  OAI211_X1 U10803 ( .C1(n9658), .C2(n9675), .A(n9657), .B(n9656), .ZN(
        P1_U3257) );
  INV_X1 U10804 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9676) );
  AOI21_X1 U10805 ( .B1(n9661), .B2(n9660), .A(n9659), .ZN(n9662) );
  NAND2_X1 U10806 ( .A1(n9663), .A2(n9662), .ZN(n9665) );
  OAI211_X1 U10807 ( .C1(n9667), .C2(n9666), .A(n9665), .B(n9664), .ZN(n9668)
         );
  INV_X1 U10808 ( .A(n9668), .ZN(n9674) );
  OAI211_X1 U10809 ( .C1(n9672), .C2(n9671), .A(n9670), .B(n9669), .ZN(n9673)
         );
  OAI211_X1 U10810 ( .C1(n9676), .C2(n9675), .A(n9674), .B(n9673), .ZN(
        P1_U3258) );
  INV_X1 U10811 ( .A(n9679), .ZN(n9680) );
  AND2_X1 U10812 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9680), .ZN(P1_U3292) );
  AND2_X1 U10813 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9680), .ZN(P1_U3293) );
  AND2_X1 U10814 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9680), .ZN(P1_U3294) );
  NOR2_X1 U10815 ( .A1(n9679), .A2(n9983), .ZN(P1_U3295) );
  AND2_X1 U10816 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9680), .ZN(P1_U3296) );
  AND2_X1 U10817 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9680), .ZN(P1_U3297) );
  NOR2_X1 U10818 ( .A1(n9679), .A2(n9967), .ZN(P1_U3298) );
  AND2_X1 U10819 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9680), .ZN(P1_U3299) );
  AND2_X1 U10820 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9680), .ZN(P1_U3300) );
  AND2_X1 U10821 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9680), .ZN(P1_U3301) );
  AND2_X1 U10822 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9680), .ZN(P1_U3302) );
  AND2_X1 U10823 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9680), .ZN(P1_U3303) );
  AND2_X1 U10824 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9680), .ZN(P1_U3304) );
  AND2_X1 U10825 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9680), .ZN(P1_U3305) );
  AND2_X1 U10826 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9680), .ZN(P1_U3306) );
  AND2_X1 U10827 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9680), .ZN(P1_U3307) );
  AND2_X1 U10828 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9680), .ZN(P1_U3308) );
  AND2_X1 U10829 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9680), .ZN(P1_U3309) );
  AND2_X1 U10830 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9680), .ZN(P1_U3310) );
  AND2_X1 U10831 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9680), .ZN(P1_U3311) );
  AND2_X1 U10832 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9680), .ZN(P1_U3312) );
  AND2_X1 U10833 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9680), .ZN(P1_U3313) );
  AND2_X1 U10834 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9680), .ZN(P1_U3314) );
  NOR2_X1 U10835 ( .A1(n9679), .A2(n10007), .ZN(P1_U3315) );
  AND2_X1 U10836 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9680), .ZN(P1_U3316) );
  AND2_X1 U10837 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9680), .ZN(P1_U3317) );
  AND2_X1 U10838 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9680), .ZN(P1_U3318) );
  NOR2_X1 U10839 ( .A1(n9679), .A2(n10054), .ZN(P1_U3319) );
  AND2_X1 U10840 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9680), .ZN(P1_U3320) );
  AND2_X1 U10841 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9680), .ZN(P1_U3321) );
  OAI22_X1 U10842 ( .A1(n9682), .A2(n9723), .B1(n9681), .B2(n9705), .ZN(n9684)
         );
  AOI211_X1 U10843 ( .C1(n9686), .C2(n9685), .A(n9684), .B(n9683), .ZN(n9730)
         );
  AOI22_X1 U10844 ( .A1(n9729), .A2(n9730), .B1(n5248), .B2(n9727), .ZN(
        P1_U3463) );
  OR2_X1 U10845 ( .A1(n9688), .A2(n9687), .ZN(n9694) );
  NAND2_X1 U10846 ( .A1(n9709), .A2(n9689), .ZN(n9690) );
  AND2_X1 U10847 ( .A1(n9691), .A2(n9690), .ZN(n9692) );
  INV_X1 U10848 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9695) );
  AOI22_X1 U10849 ( .A1(n9729), .A2(n9731), .B1(n9695), .B2(n9727), .ZN(
        P1_U3469) );
  INV_X1 U10850 ( .A(n9700), .ZN(n9702) );
  AOI22_X1 U10851 ( .A1(n9697), .A2(n9711), .B1(n9696), .B2(n9709), .ZN(n9698)
         );
  OAI211_X1 U10852 ( .C1(n9700), .C2(n9715), .A(n9699), .B(n9698), .ZN(n9701)
         );
  AOI21_X1 U10853 ( .B1(n9719), .B2(n9702), .A(n9701), .ZN(n9732) );
  AOI22_X1 U10854 ( .A1(n9729), .A2(n9732), .B1(n5308), .B2(n9727), .ZN(
        P1_U3472) );
  OAI211_X1 U10855 ( .C1(n9706), .C2(n9705), .A(n9704), .B(n9703), .ZN(n9707)
         );
  AOI21_X1 U10856 ( .B1(n9725), .B2(n9708), .A(n9707), .ZN(n9733) );
  INV_X1 U10857 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10130) );
  AOI22_X1 U10858 ( .A1(n9729), .A2(n9733), .B1(n10130), .B2(n9727), .ZN(
        P1_U3475) );
  AOI22_X1 U10859 ( .A1(n9712), .A2(n9711), .B1(n4403), .B2(n9709), .ZN(n9713)
         );
  OAI211_X1 U10860 ( .C1(n9716), .C2(n9715), .A(n9714), .B(n9713), .ZN(n9717)
         );
  AOI21_X1 U10861 ( .B1(n9719), .B2(n9718), .A(n9717), .ZN(n9734) );
  AOI22_X1 U10862 ( .A1(n9729), .A2(n9734), .B1(n5352), .B2(n9727), .ZN(
        P1_U3478) );
  OAI211_X1 U10863 ( .C1(n9723), .C2(n9722), .A(n9721), .B(n9720), .ZN(n9724)
         );
  AOI21_X1 U10864 ( .B1(n9726), .B2(n9725), .A(n9724), .ZN(n9736) );
  INV_X1 U10865 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9728) );
  AOI22_X1 U10866 ( .A1(n9729), .A2(n9736), .B1(n9728), .B2(n9727), .ZN(
        P1_U3481) );
  AOI22_X1 U10867 ( .A1(n9737), .A2(n9730), .B1(n6257), .B2(n9735), .ZN(
        P1_U3526) );
  AOI22_X1 U10868 ( .A1(n9737), .A2(n9731), .B1(n5291), .B2(n9735), .ZN(
        P1_U3528) );
  AOI22_X1 U10869 ( .A1(n9737), .A2(n9732), .B1(n6262), .B2(n9735), .ZN(
        P1_U3529) );
  AOI22_X1 U10870 ( .A1(n9737), .A2(n9733), .B1(n5333), .B2(n9735), .ZN(
        P1_U3530) );
  AOI22_X1 U10871 ( .A1(n9737), .A2(n9734), .B1(n6266), .B2(n9735), .ZN(
        P1_U3531) );
  AOI22_X1 U10872 ( .A1(n9737), .A2(n9736), .B1(n5373), .B2(n9735), .ZN(
        P1_U3532) );
  AOI22_X1 U10873 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n9896), .B1(n9891), .B2(
        P2_REG1_REG_0__SCAN_IN), .ZN(n9746) );
  AOI21_X1 U10874 ( .B1(n9739), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n9738), .ZN(
        n9745) );
  NOR2_X1 U10875 ( .A1(n9740), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9743) );
  OAI21_X1 U10876 ( .B1(n9741), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9900), .ZN(
        n9742) );
  OAI21_X1 U10877 ( .B1(n9743), .B2(n9742), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9744) );
  OAI211_X1 U10878 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9746), .A(n9745), .B(
        n9744), .ZN(P2_U3245) );
  INV_X1 U10879 ( .A(n9747), .ZN(n9750) );
  OAI21_X1 U10880 ( .B1(n9750), .B2(n9749), .A(n9748), .ZN(n9755) );
  AOI22_X1 U10881 ( .A1(n9752), .A2(n6506), .B1(n6484), .B2(n9751), .ZN(n9753)
         );
  OAI21_X1 U10882 ( .B1(n9755), .B2(n9754), .A(n9753), .ZN(n9785) );
  AOI22_X1 U10883 ( .A1(n9756), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n9768), .B2(
        n9785), .ZN(n9767) );
  OAI211_X1 U10884 ( .C1(n9759), .C2(n9758), .A(n9757), .B(n9816), .ZN(n9761)
         );
  NAND2_X1 U10885 ( .A1(n6504), .A2(n9815), .ZN(n9760) );
  NAND2_X1 U10886 ( .A1(n9761), .A2(n9760), .ZN(n9786) );
  OAI21_X1 U10887 ( .B1(n9747), .B2(n9763), .A(n9762), .ZN(n9787) );
  AOI22_X1 U10888 ( .A1(n9765), .A2(n9786), .B1(n9764), .B2(n9787), .ZN(n9766)
         );
  OAI211_X1 U10889 ( .C1(n6165), .C2(n9768), .A(n9767), .B(n9766), .ZN(
        P2_U3295) );
  INV_X1 U10890 ( .A(n9769), .ZN(n9770) );
  AND2_X1 U10891 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9775), .ZN(P2_U3297) );
  AND2_X1 U10892 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9775), .ZN(P2_U3298) );
  AND2_X1 U10893 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9775), .ZN(P2_U3299) );
  AND2_X1 U10894 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9775), .ZN(P2_U3300) );
  AND2_X1 U10895 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9775), .ZN(P2_U3301) );
  AND2_X1 U10896 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9775), .ZN(P2_U3302) );
  AND2_X1 U10897 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9775), .ZN(P2_U3303) );
  AND2_X1 U10898 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9775), .ZN(P2_U3304) );
  AND2_X1 U10899 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9775), .ZN(P2_U3305) );
  AND2_X1 U10900 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9775), .ZN(P2_U3306) );
  AND2_X1 U10901 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9775), .ZN(P2_U3307) );
  AND2_X1 U10902 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9775), .ZN(P2_U3308) );
  AND2_X1 U10903 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9775), .ZN(P2_U3309) );
  AND2_X1 U10904 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9775), .ZN(P2_U3310) );
  AND2_X1 U10905 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9775), .ZN(P2_U3311) );
  AND2_X1 U10906 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9775), .ZN(P2_U3312) );
  INV_X1 U10907 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10156) );
  NOR2_X1 U10908 ( .A1(n9772), .A2(n10156), .ZN(P2_U3313) );
  AND2_X1 U10909 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9775), .ZN(P2_U3314) );
  AND2_X1 U10910 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9775), .ZN(P2_U3315) );
  INV_X1 U10911 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10144) );
  NOR2_X1 U10912 ( .A1(n9772), .A2(n10144), .ZN(P2_U3316) );
  AND2_X1 U10913 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9775), .ZN(P2_U3317) );
  AND2_X1 U10914 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9775), .ZN(P2_U3318) );
  INV_X1 U10915 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10188) );
  NOR2_X1 U10916 ( .A1(n9772), .A2(n10188), .ZN(P2_U3319) );
  AND2_X1 U10917 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9775), .ZN(P2_U3320) );
  AND2_X1 U10918 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9775), .ZN(P2_U3321) );
  INV_X1 U10919 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n10099) );
  NOR2_X1 U10920 ( .A1(n9772), .A2(n10099), .ZN(P2_U3322) );
  AND2_X1 U10921 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9775), .ZN(P2_U3323) );
  INV_X1 U10922 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n10025) );
  NOR2_X1 U10923 ( .A1(n9772), .A2(n10025), .ZN(P2_U3324) );
  INV_X1 U10924 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10039) );
  NOR2_X1 U10925 ( .A1(n9772), .A2(n10039), .ZN(P2_U3325) );
  AND2_X1 U10926 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9775), .ZN(P2_U3326) );
  INV_X1 U10927 ( .A(n9773), .ZN(n9774) );
  AOI22_X1 U10928 ( .A1(n9774), .A2(n9777), .B1(n6013), .B2(n9775), .ZN(
        P2_U3437) );
  AOI22_X1 U10929 ( .A1(n9778), .A2(n9777), .B1(n9776), .B2(n9775), .ZN(
        P2_U3438) );
  AOI22_X1 U10930 ( .A1(n9781), .A2(n9837), .B1(n9780), .B2(n9779), .ZN(n9782)
         );
  AND2_X1 U10931 ( .A1(n9783), .A2(n9782), .ZN(n9841) );
  INV_X1 U10932 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9784) );
  AOI22_X1 U10933 ( .A1(n4405), .A2(n9841), .B1(n9784), .B2(n9839), .ZN(
        P2_U3451) );
  AOI211_X1 U10934 ( .C1(n9837), .C2(n9787), .A(n9786), .B(n9785), .ZN(n9842)
         );
  INV_X1 U10935 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10037) );
  AOI22_X1 U10936 ( .A1(n4405), .A2(n9842), .B1(n10037), .B2(n9839), .ZN(
        P2_U3454) );
  OAI21_X1 U10937 ( .B1(n9789), .B2(n9831), .A(n9788), .ZN(n9791) );
  AOI211_X1 U10938 ( .C1(n9837), .C2(n9792), .A(n9791), .B(n9790), .ZN(n9843)
         );
  INV_X1 U10939 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9793) );
  AOI22_X1 U10940 ( .A1(n4405), .A2(n9843), .B1(n9793), .B2(n9839), .ZN(
        P2_U3457) );
  INV_X1 U10941 ( .A(n9798), .ZN(n9801) );
  OAI211_X1 U10942 ( .C1(n9796), .C2(n9831), .A(n9795), .B(n9794), .ZN(n9800)
         );
  NOR2_X1 U10943 ( .A1(n9798), .A2(n9797), .ZN(n9799) );
  AOI211_X1 U10944 ( .C1(n9801), .C2(n9829), .A(n9800), .B(n9799), .ZN(n9844)
         );
  INV_X1 U10945 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9802) );
  AOI22_X1 U10946 ( .A1(n4405), .A2(n9844), .B1(n9802), .B2(n9839), .ZN(
        P2_U3460) );
  OAI22_X1 U10947 ( .A1(n9804), .A2(n9833), .B1(n9803), .B2(n9831), .ZN(n9806)
         );
  AOI211_X1 U10948 ( .C1(n9837), .C2(n9807), .A(n9806), .B(n9805), .ZN(n9845)
         );
  AOI22_X1 U10949 ( .A1(n4405), .A2(n9845), .B1(n5946), .B2(n9839), .ZN(
        P2_U3463) );
  OAI22_X1 U10950 ( .A1(n9809), .A2(n9833), .B1(n9808), .B2(n9831), .ZN(n9811)
         );
  AOI211_X1 U10951 ( .C1(n9812), .C2(n9837), .A(n9811), .B(n9810), .ZN(n9846)
         );
  INV_X1 U10952 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9813) );
  AOI22_X1 U10953 ( .A1(n4405), .A2(n9846), .B1(n9813), .B2(n9839), .ZN(
        P2_U3469) );
  AOI22_X1 U10954 ( .A1(n9817), .A2(n9816), .B1(n9815), .B2(n9814), .ZN(n9818)
         );
  OAI21_X1 U10955 ( .B1(n9820), .B2(n9819), .A(n9818), .ZN(n9821) );
  NOR2_X1 U10956 ( .A1(n9822), .A2(n9821), .ZN(n9848) );
  AOI22_X1 U10957 ( .A1(n4405), .A2(n9848), .B1(n6041), .B2(n9839), .ZN(
        P2_U3475) );
  INV_X1 U10958 ( .A(n9823), .ZN(n9828) );
  OAI22_X1 U10959 ( .A1(n9825), .A2(n9833), .B1(n9824), .B2(n9831), .ZN(n9827)
         );
  AOI211_X1 U10960 ( .C1(n9829), .C2(n9828), .A(n9827), .B(n9826), .ZN(n9849)
         );
  INV_X1 U10961 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9830) );
  AOI22_X1 U10962 ( .A1(n4405), .A2(n9849), .B1(n9830), .B2(n9839), .ZN(
        P2_U3481) );
  OAI22_X1 U10963 ( .A1(n9834), .A2(n9833), .B1(n9832), .B2(n9831), .ZN(n9836)
         );
  AOI211_X1 U10964 ( .C1(n9838), .C2(n9837), .A(n9836), .B(n9835), .ZN(n9852)
         );
  INV_X1 U10965 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9840) );
  AOI22_X1 U10966 ( .A1(n4405), .A2(n9852), .B1(n9840), .B2(n9839), .ZN(
        P2_U3487) );
  AOI22_X1 U10967 ( .A1(n9853), .A2(n9841), .B1(n5897), .B2(n9850), .ZN(
        P2_U3520) );
  AOI22_X1 U10968 ( .A1(n9853), .A2(n9842), .B1(n6147), .B2(n9850), .ZN(
        P2_U3521) );
  AOI22_X1 U10969 ( .A1(n9853), .A2(n9843), .B1(n6146), .B2(n9850), .ZN(
        P2_U3522) );
  AOI22_X1 U10970 ( .A1(n9853), .A2(n9844), .B1(n6145), .B2(n9850), .ZN(
        P2_U3523) );
  AOI22_X1 U10971 ( .A1(n9853), .A2(n9845), .B1(n6150), .B2(n9850), .ZN(
        P2_U3524) );
  AOI22_X1 U10972 ( .A1(n9853), .A2(n9846), .B1(n6208), .B2(n9850), .ZN(
        P2_U3526) );
  AOI22_X1 U10973 ( .A1(n9853), .A2(n9848), .B1(n9847), .B2(n9850), .ZN(
        P2_U3528) );
  AOI22_X1 U10974 ( .A1(n9853), .A2(n9849), .B1(n10098), .B2(n9850), .ZN(
        P2_U3530) );
  AOI22_X1 U10975 ( .A1(n9853), .A2(n9852), .B1(n9851), .B2(n9850), .ZN(
        P2_U3532) );
  INV_X1 U10976 ( .A(n9854), .ZN(n9855) );
  NAND2_X1 U10977 ( .A1(n9856), .A2(n9855), .ZN(n9857) );
  XNOR2_X1 U10978 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9857), .ZN(ADD_1071_U5) );
  XOR2_X1 U10979 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U10980 ( .B1(n9860), .B2(n9859), .A(n9858), .ZN(ADD_1071_U56) );
  OAI21_X1 U10981 ( .B1(n9863), .B2(n9862), .A(n9861), .ZN(ADD_1071_U57) );
  OAI21_X1 U10982 ( .B1(n9866), .B2(n9865), .A(n9864), .ZN(ADD_1071_U58) );
  OAI21_X1 U10983 ( .B1(n9869), .B2(n9868), .A(n9867), .ZN(ADD_1071_U59) );
  OAI21_X1 U10984 ( .B1(n9872), .B2(n9871), .A(n9870), .ZN(ADD_1071_U60) );
  OAI21_X1 U10985 ( .B1(n9875), .B2(n9874), .A(n9873), .ZN(ADD_1071_U61) );
  AOI21_X1 U10986 ( .B1(n9878), .B2(n9877), .A(n9876), .ZN(ADD_1071_U62) );
  AOI21_X1 U10987 ( .B1(n9881), .B2(n9880), .A(n9879), .ZN(ADD_1071_U63) );
  OAI21_X1 U10988 ( .B1(n9884), .B2(n9883), .A(n9882), .ZN(n9885) );
  INV_X1 U10989 ( .A(n9885), .ZN(n9890) );
  INV_X1 U10990 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n9887) );
  OAI21_X1 U10991 ( .B1(n9888), .B2(n9887), .A(n9886), .ZN(n9889) );
  AOI21_X1 U10992 ( .B1(n9891), .B2(n9890), .A(n9889), .ZN(n9898) );
  AOI21_X1 U10993 ( .B1(n9894), .B2(n9893), .A(n9892), .ZN(n9895) );
  NAND2_X1 U10994 ( .A1(n9896), .A2(n9895), .ZN(n9897) );
  OAI211_X1 U10995 ( .C1(n9900), .C2(n9899), .A(n9898), .B(n9897), .ZN(n9901)
         );
  INV_X1 U10996 ( .A(n9901), .ZN(n10207) );
  NOR4_X1 U10997 ( .A1(keyinput23), .A2(keyinput34), .A3(keyinput87), .A4(
        keyinput107), .ZN(n9902) );
  NAND4_X1 U10998 ( .A1(keyinput125), .A2(keyinput64), .A3(keyinput60), .A4(
        n9902), .ZN(n9916) );
  NOR2_X1 U10999 ( .A1(keyinput83), .A2(keyinput102), .ZN(n9903) );
  NAND3_X1 U11000 ( .A1(keyinput118), .A2(keyinput56), .A3(n9903), .ZN(n9915)
         );
  NOR2_X1 U11001 ( .A1(keyinput94), .A2(keyinput52), .ZN(n9904) );
  NAND3_X1 U11002 ( .A1(keyinput2), .A2(keyinput35), .A3(n9904), .ZN(n9914) );
  NAND2_X1 U11003 ( .A1(keyinput79), .A2(keyinput12), .ZN(n9905) );
  NOR3_X1 U11004 ( .A1(keyinput24), .A2(keyinput126), .A3(n9905), .ZN(n9912)
         );
  INV_X1 U11005 ( .A(keyinput63), .ZN(n9906) );
  NOR4_X1 U11006 ( .A1(keyinput25), .A2(keyinput114), .A3(keyinput10), .A4(
        n9906), .ZN(n9911) );
  NAND2_X1 U11007 ( .A1(keyinput106), .A2(keyinput57), .ZN(n9907) );
  NOR3_X1 U11008 ( .A1(keyinput95), .A2(keyinput30), .A3(n9907), .ZN(n9910) );
  INV_X1 U11009 ( .A(keyinput112), .ZN(n9908) );
  NOR4_X1 U11010 ( .A1(keyinput103), .A2(keyinput72), .A3(keyinput85), .A4(
        n9908), .ZN(n9909) );
  NAND4_X1 U11011 ( .A1(n9912), .A2(n9911), .A3(n9910), .A4(n9909), .ZN(n9913)
         );
  NOR4_X1 U11012 ( .A1(n9916), .A2(n9915), .A3(n9914), .A4(n9913), .ZN(n9963)
         );
  NAND4_X1 U11013 ( .A1(keyinput11), .A2(keyinput74), .A3(keyinput99), .A4(
        keyinput17), .ZN(n9917) );
  NOR3_X1 U11014 ( .A1(keyinput8), .A2(keyinput39), .A3(n9917), .ZN(n9931) );
  NAND2_X1 U11015 ( .A1(keyinput33), .A2(keyinput120), .ZN(n9918) );
  NOR3_X1 U11016 ( .A1(keyinput84), .A2(keyinput113), .A3(n9918), .ZN(n9919)
         );
  NAND3_X1 U11017 ( .A1(keyinput16), .A2(keyinput38), .A3(n9919), .ZN(n9929)
         );
  NAND2_X1 U11018 ( .A1(keyinput41), .A2(keyinput91), .ZN(n9920) );
  NOR3_X1 U11019 ( .A1(keyinput15), .A2(keyinput80), .A3(n9920), .ZN(n9927) );
  NAND2_X1 U11020 ( .A1(keyinput111), .A2(keyinput69), .ZN(n9921) );
  NOR3_X1 U11021 ( .A1(keyinput48), .A2(keyinput108), .A3(n9921), .ZN(n9926)
         );
  NAND2_X1 U11022 ( .A1(keyinput73), .A2(keyinput75), .ZN(n9922) );
  NOR3_X1 U11023 ( .A1(keyinput3), .A2(keyinput31), .A3(n9922), .ZN(n9925) );
  INV_X1 U11024 ( .A(keyinput123), .ZN(n9923) );
  NOR4_X1 U11025 ( .A1(keyinput104), .A2(keyinput21), .A3(keyinput27), .A4(
        n9923), .ZN(n9924) );
  NAND4_X1 U11026 ( .A1(n9927), .A2(n9926), .A3(n9925), .A4(n9924), .ZN(n9928)
         );
  NOR4_X1 U11027 ( .A1(keyinput62), .A2(keyinput96), .A3(n9929), .A4(n9928), 
        .ZN(n9930) );
  NAND4_X1 U11028 ( .A1(keyinput119), .A2(keyinput82), .A3(n9931), .A4(n9930), 
        .ZN(n9961) );
  NOR2_X1 U11029 ( .A1(keyinput77), .A2(keyinput90), .ZN(n9932) );
  NAND3_X1 U11030 ( .A1(keyinput50), .A2(keyinput47), .A3(n9932), .ZN(n9933)
         );
  NOR3_X1 U11031 ( .A1(keyinput6), .A2(keyinput117), .A3(n9933), .ZN(n9945) );
  NAND2_X1 U11032 ( .A1(keyinput61), .A2(keyinput65), .ZN(n9934) );
  NOR3_X1 U11033 ( .A1(keyinput122), .A2(keyinput110), .A3(n9934), .ZN(n9935)
         );
  NAND3_X1 U11034 ( .A1(keyinput36), .A2(keyinput46), .A3(n9935), .ZN(n9943)
         );
  NOR4_X1 U11035 ( .A1(keyinput116), .A2(keyinput5), .A3(keyinput40), .A4(
        keyinput121), .ZN(n9941) );
  NAND3_X1 U11036 ( .A1(keyinput66), .A2(keyinput93), .A3(keyinput43), .ZN(
        n9936) );
  NOR2_X1 U11037 ( .A1(keyinput71), .A2(n9936), .ZN(n9940) );
  NOR4_X1 U11038 ( .A1(keyinput59), .A2(keyinput22), .A3(keyinput20), .A4(
        keyinput45), .ZN(n9939) );
  NAND3_X1 U11039 ( .A1(keyinput49), .A2(keyinput28), .A3(keyinput13), .ZN(
        n9937) );
  NOR2_X1 U11040 ( .A1(keyinput92), .A2(n9937), .ZN(n9938) );
  NAND4_X1 U11041 ( .A1(n9941), .A2(n9940), .A3(n9939), .A4(n9938), .ZN(n9942)
         );
  NOR4_X1 U11042 ( .A1(keyinput55), .A2(keyinput37), .A3(n9943), .A4(n9942), 
        .ZN(n9944) );
  NAND4_X1 U11043 ( .A1(keyinput78), .A2(keyinput0), .A3(n9945), .A4(n9944), 
        .ZN(n9960) );
  AND4_X1 U11044 ( .A1(keyinput26), .A2(keyinput4), .A3(keyinput76), .A4(
        keyinput70), .ZN(n9951) );
  NAND2_X1 U11045 ( .A1(keyinput88), .A2(keyinput42), .ZN(n9946) );
  NOR3_X1 U11046 ( .A1(keyinput1), .A2(keyinput18), .A3(n9946), .ZN(n9950) );
  NAND2_X1 U11047 ( .A1(keyinput97), .A2(keyinput58), .ZN(n9947) );
  NOR3_X1 U11048 ( .A1(keyinput51), .A2(keyinput44), .A3(n9947), .ZN(n9949) );
  INV_X1 U11049 ( .A(keyinput100), .ZN(n10051) );
  NOR4_X1 U11050 ( .A1(keyinput9), .A2(keyinput53), .A3(keyinput109), .A4(
        n10051), .ZN(n9948) );
  NAND4_X1 U11051 ( .A1(n9951), .A2(n9950), .A3(n9949), .A4(n9948), .ZN(n9959)
         );
  NOR4_X1 U11052 ( .A1(keyinput54), .A2(keyinput105), .A3(keyinput32), .A4(
        keyinput68), .ZN(n9957) );
  INV_X1 U11053 ( .A(keyinput98), .ZN(n9952) );
  NOR4_X1 U11054 ( .A1(keyinput89), .A2(keyinput19), .A3(keyinput67), .A4(
        n9952), .ZN(n9956) );
  INV_X1 U11055 ( .A(keyinput81), .ZN(n9953) );
  NOR4_X1 U11056 ( .A1(keyinput101), .A2(keyinput7), .A3(keyinput86), .A4(
        n9953), .ZN(n9955) );
  AND4_X1 U11057 ( .A1(keyinput29), .A2(keyinput124), .A3(keyinput14), .A4(
        keyinput115), .ZN(n9954) );
  NAND4_X1 U11058 ( .A1(n9957), .A2(n9956), .A3(n9955), .A4(n9954), .ZN(n9958)
         );
  NOR4_X1 U11059 ( .A1(n9961), .A2(n9960), .A3(n9959), .A4(n9958), .ZN(n9962)
         );
  AOI21_X1 U11060 ( .B1(n9963), .B2(n9962), .A(keyinput127), .ZN(n10205) );
  AOI22_X1 U11061 ( .A1(n5151), .A2(keyinput43), .B1(keyinput116), .B2(n9965), 
        .ZN(n9964) );
  OAI221_X1 U11062 ( .B1(n5151), .B2(keyinput43), .C1(n9965), .C2(keyinput116), 
        .A(n9964), .ZN(n9977) );
  INV_X1 U11063 ( .A(SI_5_), .ZN(n9968) );
  AOI22_X1 U11064 ( .A1(n9968), .A2(keyinput5), .B1(n9967), .B2(keyinput40), 
        .ZN(n9966) );
  OAI221_X1 U11065 ( .B1(n9968), .B2(keyinput5), .C1(n9967), .C2(keyinput40), 
        .A(n9966), .ZN(n9976) );
  AOI22_X1 U11066 ( .A1(n9971), .A2(keyinput121), .B1(n9970), .B2(keyinput93), 
        .ZN(n9969) );
  OAI221_X1 U11067 ( .B1(n9971), .B2(keyinput121), .C1(n9970), .C2(keyinput93), 
        .A(n9969), .ZN(n9975) );
  AOI22_X1 U11068 ( .A1(n5850), .A2(keyinput66), .B1(n9973), .B2(keyinput77), 
        .ZN(n9972) );
  OAI221_X1 U11069 ( .B1(n5850), .B2(keyinput66), .C1(n9973), .C2(keyinput77), 
        .A(n9972), .ZN(n9974) );
  NOR4_X1 U11070 ( .A1(n9977), .A2(n9976), .A3(n9975), .A4(n9974), .ZN(n10023)
         );
  AOI22_X1 U11071 ( .A1(n9979), .A2(keyinput50), .B1(n4880), .B2(keyinput78), 
        .ZN(n9978) );
  OAI221_X1 U11072 ( .B1(n9979), .B2(keyinput50), .C1(n4880), .C2(keyinput78), 
        .A(n9978), .ZN(n9990) );
  AOI22_X1 U11073 ( .A1(n9981), .A2(keyinput0), .B1(keyinput47), .B2(n6827), 
        .ZN(n9980) );
  OAI221_X1 U11074 ( .B1(n9981), .B2(keyinput0), .C1(n6827), .C2(keyinput47), 
        .A(n9980), .ZN(n9989) );
  INV_X1 U11075 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n9984) );
  AOI22_X1 U11076 ( .A1(n9984), .A2(keyinput90), .B1(n9983), .B2(keyinput6), 
        .ZN(n9982) );
  OAI221_X1 U11077 ( .B1(n9984), .B2(keyinput90), .C1(n9983), .C2(keyinput6), 
        .A(n9982), .ZN(n9988) );
  INV_X1 U11078 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9986) );
  AOI22_X1 U11079 ( .A1(n9986), .A2(keyinput117), .B1(keyinput28), .B2(n5648), 
        .ZN(n9985) );
  OAI221_X1 U11080 ( .B1(n9986), .B2(keyinput117), .C1(n5648), .C2(keyinput28), 
        .A(n9985), .ZN(n9987) );
  NOR4_X1 U11081 ( .A1(n9990), .A2(n9989), .A3(n9988), .A4(n9987), .ZN(n10022)
         );
  AOI22_X1 U11082 ( .A1(n9992), .A2(keyinput13), .B1(n5567), .B2(keyinput92), 
        .ZN(n9991) );
  OAI221_X1 U11083 ( .B1(n9992), .B2(keyinput13), .C1(n5567), .C2(keyinput92), 
        .A(n9991), .ZN(n10004) );
  AOI22_X1 U11084 ( .A1(n6013), .A2(keyinput49), .B1(keyinput59), .B2(n9994), 
        .ZN(n9993) );
  OAI221_X1 U11085 ( .B1(n6013), .B2(keyinput49), .C1(n9994), .C2(keyinput59), 
        .A(n9993), .ZN(n10003) );
  AOI22_X1 U11086 ( .A1(n9997), .A2(keyinput22), .B1(keyinput20), .B2(n9996), 
        .ZN(n9995) );
  OAI221_X1 U11087 ( .B1(n9997), .B2(keyinput22), .C1(n9996), .C2(keyinput20), 
        .A(n9995), .ZN(n10002) );
  AOI22_X1 U11088 ( .A1(n10000), .A2(keyinput45), .B1(n9999), .B2(keyinput55), 
        .ZN(n9998) );
  OAI221_X1 U11089 ( .B1(n10000), .B2(keyinput45), .C1(n9999), .C2(keyinput55), 
        .A(n9998), .ZN(n10001) );
  NOR4_X1 U11090 ( .A1(n10004), .A2(n10003), .A3(n10002), .A4(n10001), .ZN(
        n10021) );
  AOI22_X1 U11091 ( .A1(n5448), .A2(keyinput65), .B1(n10006), .B2(keyinput61), 
        .ZN(n10005) );
  OAI221_X1 U11092 ( .B1(n5448), .B2(keyinput65), .C1(n10006), .C2(keyinput61), 
        .A(n10005), .ZN(n10011) );
  XNOR2_X1 U11093 ( .A(n10007), .B(keyinput37), .ZN(n10010) );
  XNOR2_X1 U11094 ( .A(n10008), .B(keyinput122), .ZN(n10009) );
  OR3_X1 U11095 ( .A1(n10011), .A2(n10010), .A3(n10009), .ZN(n10019) );
  INV_X1 U11096 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n10013) );
  AOI22_X1 U11097 ( .A1(n10013), .A2(keyinput110), .B1(n5897), .B2(keyinput36), 
        .ZN(n10012) );
  OAI221_X1 U11098 ( .B1(n10013), .B2(keyinput110), .C1(n5897), .C2(keyinput36), .A(n10012), .ZN(n10018) );
  INV_X1 U11099 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10015) );
  AOI22_X1 U11100 ( .A1(n10016), .A2(keyinput46), .B1(keyinput98), .B2(n10015), 
        .ZN(n10014) );
  OAI221_X1 U11101 ( .B1(n10016), .B2(keyinput46), .C1(n10015), .C2(keyinput98), .A(n10014), .ZN(n10017) );
  NOR3_X1 U11102 ( .A1(n10019), .A2(n10018), .A3(n10017), .ZN(n10020) );
  NAND4_X1 U11103 ( .A1(n10023), .A2(n10022), .A3(n10021), .A4(n10020), .ZN(
        n10203) );
  AOI22_X1 U11104 ( .A1(n10026), .A2(keyinput67), .B1(keyinput54), .B2(n10025), 
        .ZN(n10024) );
  OAI221_X1 U11105 ( .B1(n10026), .B2(keyinput67), .C1(n10025), .C2(keyinput54), .A(n10024), .ZN(n10034) );
  AOI22_X1 U11106 ( .A1(n6785), .A2(keyinput19), .B1(n5291), .B2(keyinput89), 
        .ZN(n10027) );
  OAI221_X1 U11107 ( .B1(n6785), .B2(keyinput19), .C1(n5291), .C2(keyinput89), 
        .A(n10027), .ZN(n10033) );
  AOI22_X1 U11108 ( .A1(n5248), .A2(keyinput68), .B1(n5308), .B2(keyinput42), 
        .ZN(n10028) );
  OAI221_X1 U11109 ( .B1(n5248), .B2(keyinput68), .C1(n5308), .C2(keyinput42), 
        .A(n10028), .ZN(n10032) );
  XOR2_X1 U11110 ( .A(n5122), .B(keyinput105), .Z(n10030) );
  XNOR2_X1 U11111 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput32), .ZN(n10029) );
  NAND2_X1 U11112 ( .A1(n10030), .A2(n10029), .ZN(n10031) );
  NOR4_X1 U11113 ( .A1(n10034), .A2(n10033), .A3(n10032), .A4(n10031), .ZN(
        n10082) );
  AOI22_X1 U11114 ( .A1(n10037), .A2(keyinput88), .B1(n10036), .B2(keyinput9), 
        .ZN(n10035) );
  OAI221_X1 U11115 ( .B1(n10037), .B2(keyinput88), .C1(n10036), .C2(keyinput9), 
        .A(n10035), .ZN(n10049) );
  AOI22_X1 U11116 ( .A1(n10040), .A2(keyinput4), .B1(n10039), .B2(keyinput76), 
        .ZN(n10038) );
  OAI221_X1 U11117 ( .B1(n10040), .B2(keyinput4), .C1(n10039), .C2(keyinput76), 
        .A(n10038), .ZN(n10048) );
  AOI22_X1 U11118 ( .A1(n10043), .A2(keyinput18), .B1(keyinput26), .B2(n10042), 
        .ZN(n10041) );
  OAI221_X1 U11119 ( .B1(n10043), .B2(keyinput18), .C1(n10042), .C2(keyinput26), .A(n10041), .ZN(n10047) );
  XNOR2_X1 U11120 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput1), .ZN(n10045) );
  XNOR2_X1 U11121 ( .A(SI_26_), .B(keyinput70), .ZN(n10044) );
  NAND2_X1 U11122 ( .A1(n10045), .A2(n10044), .ZN(n10046) );
  NOR4_X1 U11123 ( .A1(n10049), .A2(n10048), .A3(n10047), .A4(n10046), .ZN(
        n10081) );
  AOI22_X1 U11124 ( .A1(n10052), .A2(keyinput53), .B1(P2_WR_REG_SCAN_IN), .B2(
        n10051), .ZN(n10050) );
  OAI221_X1 U11125 ( .B1(n10052), .B2(keyinput53), .C1(n10051), .C2(
        P2_WR_REG_SCAN_IN), .A(n10050), .ZN(n10064) );
  AOI22_X1 U11126 ( .A1(n10055), .A2(keyinput109), .B1(n10054), .B2(keyinput58), .ZN(n10053) );
  OAI221_X1 U11127 ( .B1(n10055), .B2(keyinput109), .C1(n10054), .C2(
        keyinput58), .A(n10053), .ZN(n10063) );
  AOI22_X1 U11128 ( .A1(n10058), .A2(keyinput51), .B1(n10057), .B2(keyinput97), 
        .ZN(n10056) );
  OAI221_X1 U11129 ( .B1(n10058), .B2(keyinput51), .C1(n10057), .C2(keyinput97), .A(n10056), .ZN(n10062) );
  INV_X1 U11130 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10212) );
  AOI22_X1 U11131 ( .A1(n10212), .A2(keyinput44), .B1(n10060), .B2(keyinput29), 
        .ZN(n10059) );
  OAI221_X1 U11132 ( .B1(n10212), .B2(keyinput44), .C1(n10060), .C2(keyinput29), .A(n10059), .ZN(n10061) );
  NOR4_X1 U11133 ( .A1(n10064), .A2(n10063), .A3(n10062), .A4(n10061), .ZN(
        n10080) );
  AOI22_X1 U11134 ( .A1(n6266), .A2(keyinput124), .B1(keyinput14), .B2(n10066), 
        .ZN(n10065) );
  OAI221_X1 U11135 ( .B1(n6266), .B2(keyinput124), .C1(n10066), .C2(keyinput14), .A(n10065), .ZN(n10078) );
  AOI22_X1 U11136 ( .A1(n7708), .A2(keyinput115), .B1(keyinput101), .B2(n10068), .ZN(n10067) );
  OAI221_X1 U11137 ( .B1(n7708), .B2(keyinput115), .C1(n10068), .C2(
        keyinput101), .A(n10067), .ZN(n10077) );
  AOI22_X1 U11138 ( .A1(n10071), .A2(keyinput7), .B1(keyinput86), .B2(n10070), 
        .ZN(n10069) );
  OAI221_X1 U11139 ( .B1(n10071), .B2(keyinput7), .C1(n10070), .C2(keyinput86), 
        .A(n10069), .ZN(n10076) );
  INV_X1 U11140 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10073) );
  AOI22_X1 U11141 ( .A1(n10074), .A2(keyinput125), .B1(keyinput81), .B2(n10073), .ZN(n10072) );
  OAI221_X1 U11142 ( .B1(n10074), .B2(keyinput125), .C1(n10073), .C2(
        keyinput81), .A(n10072), .ZN(n10075) );
  NOR4_X1 U11143 ( .A1(n10078), .A2(n10077), .A3(n10076), .A4(n10075), .ZN(
        n10079) );
  NAND4_X1 U11144 ( .A1(n10082), .A2(n10081), .A3(n10080), .A4(n10079), .ZN(
        n10202) );
  AOI22_X1 U11145 ( .A1(n6208), .A2(keyinput111), .B1(keyinput15), .B2(n6586), 
        .ZN(n10083) );
  OAI221_X1 U11146 ( .B1(n6208), .B2(keyinput111), .C1(n6586), .C2(keyinput15), 
        .A(n10083), .ZN(n10096) );
  AOI22_X1 U11147 ( .A1(n10086), .A2(keyinput69), .B1(keyinput108), .B2(n10085), .ZN(n10084) );
  OAI221_X1 U11148 ( .B1(n10086), .B2(keyinput69), .C1(n10085), .C2(
        keyinput108), .A(n10084), .ZN(n10095) );
  INV_X1 U11149 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n10088) );
  AOI22_X1 U11150 ( .A1(n10089), .A2(keyinput80), .B1(keyinput62), .B2(n10088), 
        .ZN(n10087) );
  OAI221_X1 U11151 ( .B1(n10089), .B2(keyinput80), .C1(n10088), .C2(keyinput62), .A(n10087), .ZN(n10094) );
  AOI22_X1 U11152 ( .A1(n10092), .A2(keyinput91), .B1(keyinput41), .B2(n10091), 
        .ZN(n10090) );
  OAI221_X1 U11153 ( .B1(n10092), .B2(keyinput91), .C1(n10091), .C2(keyinput41), .A(n10090), .ZN(n10093) );
  NOR4_X1 U11154 ( .A1(n10096), .A2(n10095), .A3(n10094), .A4(n10093), .ZN(
        n10140) );
  AOI22_X1 U11155 ( .A1(n10099), .A2(keyinput39), .B1(keyinput48), .B2(n10098), 
        .ZN(n10097) );
  OAI221_X1 U11156 ( .B1(n10099), .B2(keyinput39), .C1(n10098), .C2(keyinput48), .A(n10097), .ZN(n10111) );
  INV_X1 U11157 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10101) );
  AOI22_X1 U11158 ( .A1(n8333), .A2(keyinput82), .B1(n10101), .B2(keyinput11), 
        .ZN(n10100) );
  OAI221_X1 U11159 ( .B1(n8333), .B2(keyinput82), .C1(n10101), .C2(keyinput11), 
        .A(n10100), .ZN(n10110) );
  AOI22_X1 U11160 ( .A1(n10104), .A2(keyinput74), .B1(keyinput99), .B2(n10103), 
        .ZN(n10102) );
  OAI221_X1 U11161 ( .B1(n10104), .B2(keyinput74), .C1(n10103), .C2(keyinput99), .A(n10102), .ZN(n10109) );
  XOR2_X1 U11162 ( .A(n10105), .B(keyinput8), .Z(n10107) );
  XNOR2_X1 U11163 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput17), .ZN(n10106) );
  NAND2_X1 U11164 ( .A1(n10107), .A2(n10106), .ZN(n10108) );
  NOR4_X1 U11165 ( .A1(n10111), .A2(n10110), .A3(n10109), .A4(n10108), .ZN(
        n10139) );
  AOI22_X1 U11166 ( .A1(n10222), .A2(keyinput27), .B1(n9478), .B2(keyinput75), 
        .ZN(n10112) );
  OAI221_X1 U11167 ( .B1(n10222), .B2(keyinput27), .C1(n9478), .C2(keyinput75), 
        .A(n10112), .ZN(n10123) );
  INV_X1 U11168 ( .A(P1_RD_REG_SCAN_IN), .ZN(n10114) );
  AOI22_X1 U11169 ( .A1(n6226), .A2(keyinput21), .B1(n10114), .B2(keyinput104), 
        .ZN(n10113) );
  OAI221_X1 U11170 ( .B1(n6226), .B2(keyinput21), .C1(n10114), .C2(keyinput104), .A(n10113), .ZN(n10122) );
  AOI22_X1 U11171 ( .A1(n10117), .A2(keyinput31), .B1(keyinput71), .B2(n10116), 
        .ZN(n10115) );
  OAI221_X1 U11172 ( .B1(n10117), .B2(keyinput31), .C1(n10116), .C2(keyinput71), .A(n10115), .ZN(n10121) );
  INV_X1 U11173 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n10119) );
  AOI22_X1 U11174 ( .A1(n10210), .A2(keyinput3), .B1(n10119), .B2(keyinput73), 
        .ZN(n10118) );
  OAI221_X1 U11175 ( .B1(n10210), .B2(keyinput3), .C1(n10119), .C2(keyinput73), 
        .A(n10118), .ZN(n10120) );
  NOR4_X1 U11176 ( .A1(n10123), .A2(n10122), .A3(n10121), .A4(n10120), .ZN(
        n10138) );
  AOI22_X1 U11177 ( .A1(n5722), .A2(keyinput120), .B1(keyinput16), .B2(n10125), 
        .ZN(n10124) );
  OAI221_X1 U11178 ( .B1(n5722), .B2(keyinput120), .C1(n10125), .C2(keyinput16), .A(n10124), .ZN(n10136) );
  INV_X1 U11179 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10128) );
  AOI22_X1 U11180 ( .A1(n10128), .A2(keyinput96), .B1(n10127), .B2(keyinput84), 
        .ZN(n10126) );
  OAI221_X1 U11181 ( .B1(n10128), .B2(keyinput96), .C1(n10127), .C2(keyinput84), .A(n10126), .ZN(n10135) );
  AOI22_X1 U11182 ( .A1(n10130), .A2(keyinput113), .B1(keyinput123), .B2(n4979), .ZN(n10129) );
  OAI221_X1 U11183 ( .B1(n10130), .B2(keyinput113), .C1(n4979), .C2(
        keyinput123), .A(n10129), .ZN(n10134) );
  AOI22_X1 U11184 ( .A1(n8897), .A2(keyinput38), .B1(n10132), .B2(keyinput33), 
        .ZN(n10131) );
  OAI221_X1 U11185 ( .B1(n8897), .B2(keyinput38), .C1(n10132), .C2(keyinput33), 
        .A(n10131), .ZN(n10133) );
  NOR4_X1 U11186 ( .A1(n10136), .A2(n10135), .A3(n10134), .A4(n10133), .ZN(
        n10137) );
  NAND4_X1 U11187 ( .A1(n10140), .A2(n10139), .A3(n10138), .A4(n10137), .ZN(
        n10201) );
  AOI22_X1 U11188 ( .A1(n10143), .A2(keyinput63), .B1(n10142), .B2(keyinput114), .ZN(n10141) );
  OAI221_X1 U11189 ( .B1(n10143), .B2(keyinput63), .C1(n10142), .C2(
        keyinput114), .A(n10141), .ZN(n10147) );
  XNOR2_X1 U11190 ( .A(n10144), .B(keyinput126), .ZN(n10146) );
  XOR2_X1 U11191 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput112), .Z(n10145) );
  OR3_X1 U11192 ( .A1(n10147), .A2(n10146), .A3(n10145), .ZN(n10154) );
  AOI22_X1 U11193 ( .A1(n8289), .A2(keyinput10), .B1(n7358), .B2(keyinput24), 
        .ZN(n10148) );
  OAI221_X1 U11194 ( .B1(n8289), .B2(keyinput10), .C1(n7358), .C2(keyinput24), 
        .A(n10148), .ZN(n10153) );
  INV_X1 U11195 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n10151) );
  AOI22_X1 U11196 ( .A1(n10151), .A2(keyinput12), .B1(n10150), .B2(keyinput79), 
        .ZN(n10149) );
  OAI221_X1 U11197 ( .B1(n10151), .B2(keyinput12), .C1(n10150), .C2(keyinput79), .A(n10149), .ZN(n10152) );
  NOR3_X1 U11198 ( .A1(n10154), .A2(n10153), .A3(n10152), .ZN(n10199) );
  NAND2_X1 U11199 ( .A1(n6172), .A2(keyinput23), .ZN(n10155) );
  OAI221_X1 U11200 ( .B1(n10156), .B2(keyinput127), .C1(n6172), .C2(keyinput23), .A(n10155), .ZN(n10167) );
  AOI22_X1 U11201 ( .A1(n10158), .A2(keyinput64), .B1(n5117), .B2(keyinput60), 
        .ZN(n10157) );
  OAI221_X1 U11202 ( .B1(n10158), .B2(keyinput64), .C1(n5117), .C2(keyinput60), 
        .A(n10157), .ZN(n10166) );
  AOI22_X1 U11203 ( .A1(n10161), .A2(keyinput107), .B1(keyinput25), .B2(n10160), .ZN(n10159) );
  OAI221_X1 U11204 ( .B1(n10161), .B2(keyinput107), .C1(n10160), .C2(
        keyinput25), .A(n10159), .ZN(n10165) );
  AOI22_X1 U11205 ( .A1(n10163), .A2(keyinput34), .B1(keyinput87), .B2(n8494), 
        .ZN(n10162) );
  OAI221_X1 U11206 ( .B1(n10163), .B2(keyinput34), .C1(n8494), .C2(keyinput87), 
        .A(n10162), .ZN(n10164) );
  NOR4_X1 U11207 ( .A1(n10167), .A2(n10166), .A3(n10165), .A4(n10164), .ZN(
        n10198) );
  INV_X1 U11208 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n10169) );
  AOI22_X1 U11209 ( .A1(n8888), .A2(keyinput35), .B1(n10169), .B2(keyinput118), 
        .ZN(n10168) );
  OAI221_X1 U11210 ( .B1(n8888), .B2(keyinput35), .C1(n10169), .C2(keyinput118), .A(n10168), .ZN(n10180) );
  AOI22_X1 U11211 ( .A1(n8312), .A2(keyinput52), .B1(n5840), .B2(keyinput94), 
        .ZN(n10170) );
  OAI221_X1 U11212 ( .B1(n8312), .B2(keyinput52), .C1(n5840), .C2(keyinput94), 
        .A(n10170), .ZN(n10179) );
  AOI22_X1 U11213 ( .A1(n10173), .A2(keyinput56), .B1(keyinput119), .B2(n10172), .ZN(n10171) );
  OAI221_X1 U11214 ( .B1(n10173), .B2(keyinput56), .C1(n10172), .C2(
        keyinput119), .A(n10171), .ZN(n10178) );
  AOI22_X1 U11215 ( .A1(n10176), .A2(keyinput102), .B1(keyinput83), .B2(n10175), .ZN(n10174) );
  OAI221_X1 U11216 ( .B1(n10176), .B2(keyinput102), .C1(n10175), .C2(
        keyinput83), .A(n10174), .ZN(n10177) );
  NOR4_X1 U11217 ( .A1(n10180), .A2(n10179), .A3(n10178), .A4(n10177), .ZN(
        n10197) );
  AOI22_X1 U11218 ( .A1(n10183), .A2(keyinput85), .B1(n10182), .B2(keyinput57), 
        .ZN(n10181) );
  OAI221_X1 U11219 ( .B1(n10183), .B2(keyinput85), .C1(n10182), .C2(keyinput57), .A(n10181), .ZN(n10195) );
  AOI22_X1 U11220 ( .A1(n8410), .A2(keyinput72), .B1(n10185), .B2(keyinput103), 
        .ZN(n10184) );
  OAI221_X1 U11221 ( .B1(n8410), .B2(keyinput72), .C1(n10185), .C2(keyinput103), .A(n10184), .ZN(n10194) );
  INV_X1 U11222 ( .A(SI_21_), .ZN(n10187) );
  AOI22_X1 U11223 ( .A1(n10188), .A2(keyinput30), .B1(n10187), .B2(keyinput2), 
        .ZN(n10186) );
  OAI221_X1 U11224 ( .B1(n10188), .B2(keyinput30), .C1(n10187), .C2(keyinput2), 
        .A(n10186), .ZN(n10193) );
  INV_X1 U11225 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n10191) );
  AOI22_X1 U11226 ( .A1(n10191), .A2(keyinput95), .B1(n10190), .B2(keyinput106), .ZN(n10189) );
  OAI221_X1 U11227 ( .B1(n10191), .B2(keyinput95), .C1(n10190), .C2(
        keyinput106), .A(n10189), .ZN(n10192) );
  NOR4_X1 U11228 ( .A1(n10195), .A2(n10194), .A3(n10193), .A4(n10192), .ZN(
        n10196) );
  NAND4_X1 U11229 ( .A1(n10199), .A2(n10198), .A3(n10197), .A4(n10196), .ZN(
        n10200) );
  NOR4_X1 U11230 ( .A1(n10203), .A2(n10202), .A3(n10201), .A4(n10200), .ZN(
        n10204) );
  OAI21_X1 U11231 ( .B1(P2_D_REG_15__SCAN_IN), .B2(n10205), .A(n10204), .ZN(
        n10206) );
  XOR2_X1 U11232 ( .A(n10207), .B(n10206), .Z(P2_U3255) );
  XOR2_X1 U11233 ( .A(n10208), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  AOI21_X1 U11234 ( .B1(n10211), .B2(n10210), .A(n10209), .ZN(ADD_1071_U47) );
  XNOR2_X1 U11235 ( .A(n10213), .B(n10212), .ZN(ADD_1071_U50) );
  NOR2_X1 U11236 ( .A1(n10215), .A2(n10214), .ZN(n10216) );
  XOR2_X1 U11237 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10216), .Z(ADD_1071_U51) );
  OAI21_X1 U11238 ( .B1(n8312), .B2(n10218), .A(n10217), .ZN(n10219) );
  XNOR2_X1 U11239 ( .A(n10219), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11240 ( .A(n10221), .B(n10220), .Z(ADD_1071_U54) );
  XNOR2_X1 U11241 ( .A(n10223), .B(n10222), .ZN(ADD_1071_U48) );
  XOR2_X1 U11242 ( .A(n10225), .B(n10224), .Z(ADD_1071_U53) );
  XNOR2_X1 U11243 ( .A(n10227), .B(n10226), .ZN(ADD_1071_U52) );
  NAND2_X1 U7391 ( .A1(n6143), .A2(n5880), .ZN(n6769) );
  AND2_X2 U4922 ( .A1(n5796), .A2(n5155), .ZN(n5801) );
  CLKBUF_X1 U4927 ( .A(n5178), .Z(n5670) );
  CLKBUF_X1 U4950 ( .A(n9710), .Z(n4403) );
endmodule

