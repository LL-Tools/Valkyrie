

module b20_C_SARLock_k_128_8 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4427, n4428, n4429, n4430, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436;

  INV_X4 U4934 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  AOI21_X1 U4935 ( .B1(n9765), .B2(n5443), .A(n4539), .ZN(n9716) );
  OR2_X1 U4936 ( .A1(n7882), .A2(n5525), .ZN(n4926) );
  OR2_X1 U4937 ( .A1(n9585), .A2(n7895), .ZN(n7893) );
  CLKBUF_X1 U4938 ( .A(n4438), .Z(n4446) );
  INV_X2 U4939 ( .A(n4430), .ZN(n4433) );
  INV_X1 U4941 ( .A(n9075), .ZN(n5483) );
  NAND2_X1 U4942 ( .A1(n5716), .A2(n5713), .ZN(n5765) );
  NAND4_X2 U4944 ( .A1(n5159), .A2(n5158), .A3(n5157), .A4(n5156), .ZN(n9829)
         );
  INV_X1 U4945 ( .A(n9848), .ZN(n9237) );
  OR2_X1 U4946 ( .A1(n6064), .A2(n6050), .ZN(n6091) );
  XNOR2_X1 U4947 ( .A(n6056), .B(n10268), .ZN(n6472) );
  NAND2_X1 U4948 ( .A1(n5098), .A2(n5097), .ZN(n7843) );
  INV_X1 U4950 ( .A(n6549), .ZN(n6550) );
  NAND2_X1 U4951 ( .A1(n5734), .A2(n5736), .ZN(n5728) );
  CLKBUF_X1 U4952 ( .A(n8047), .Z(n4427) );
  NOR2_X1 U4953 ( .A1(n6889), .A2(n6888), .ZN(n8047) );
  NAND2_X1 U4954 ( .A1(n5827), .A2(n5979), .ZN(n4643) );
  NOR2_X1 U4955 ( .A1(n5056), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n5055) );
  INV_X1 U4956 ( .A(n6077), .ZN(n4430) );
  INV_X1 U4957 ( .A(n6109), .ZN(n6183) );
  INV_X1 U4958 ( .A(n5979), .ZN(n5987) );
  INV_X1 U4959 ( .A(n6584), .ZN(n5482) );
  AND2_X1 U4960 ( .A1(n9804), .A2(n9937), .ZN(n7504) );
  OAI21_X1 U4962 ( .B1(n5126), .B2(n5100), .A(n5099), .ZN(n5124) );
  INV_X1 U4963 ( .A(n8353), .ZN(n6883) );
  NAND2_X1 U4964 ( .A1(n6064), .A2(n6048), .ZN(n6101) );
  INV_X1 U4965 ( .A(n4445), .ZN(n6365) );
  OR2_X1 U4966 ( .A1(n4445), .A2(n6713), .ZN(n6090) );
  OR2_X1 U4967 ( .A1(n6374), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6385) );
  INV_X1 U4968 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U4969 ( .A1(n4963), .A2(n5895), .ZN(n8971) );
  OAI21_X1 U4970 ( .B1(n7499), .B2(n4952), .A(n4949), .ZN(n5393) );
  NAND2_X1 U4971 ( .A1(n5330), .A2(n5329), .ZN(n7499) );
  NAND2_X1 U4972 ( .A1(n5098), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5096) );
  INV_X1 U4973 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U4974 ( .A1(n7819), .A2(n7818), .ZN(n7908) );
  NAND2_X1 U4975 ( .A1(n5800), .A2(n5799), .ZN(n6992) );
  MUX2_X1 U4976 ( .A(n9227), .B(n9226), .S(n5685), .Z(n9302) );
  AND4_X1 U4977 ( .A1(n5285), .A2(n5284), .A3(n5283), .A4(n5282), .ZN(n9927)
         );
  NAND2_X2 U4978 ( .A1(n4851), .A2(n5066), .ZN(n9848) );
  XNOR2_X1 U4979 ( .A(n5265), .B(n5264), .ZN(n6570) );
  OAI21_X1 U4980 ( .B1(n9302), .B2(n9301), .A(n9300), .ZN(n9309) );
  INV_X1 U4982 ( .A(n5685), .ZN(n5713) );
  XNOR2_X1 U4983 ( .A(n5096), .B(n5095), .ZN(n5717) );
  AND2_X1 U4984 ( .A1(n6064), .A2(n6050), .ZN(n6077) );
  AND2_X1 U4985 ( .A1(n5047), .A2(n5048), .ZN(n4428) );
  BUF_X2 U4986 ( .A(n8352), .Z(n4442) );
  NAND2_X2 U4987 ( .A1(n8025), .A2(n5068), .ZN(n8098) );
  OR2_X2 U4988 ( .A1(n9919), .A2(n9927), .ZN(n9156) );
  OAI21_X2 U4989 ( .B1(n5357), .B2(n4704), .A(n5356), .ZN(n5372) );
  OR2_X2 U4990 ( .A1(n7085), .A2(n4786), .ZN(n4782) );
  NOR2_X1 U4991 ( .A1(n9144), .A2(n5701), .ZN(n9087) );
  OAI22_X1 U4992 ( .A1(n7908), .A2(n7907), .B1(n8225), .B2(n7906), .ZN(n7975)
         );
  CLKBUF_X2 U4993 ( .A(n9828), .Z(n4429) );
  NAND4_X1 U4994 ( .A1(n5120), .A2(n5119), .A3(n5118), .A4(n5117), .ZN(n9828)
         );
  NAND3_X4 U4996 ( .A1(n6094), .A2(n6093), .A3(n6092), .ZN(n8351) );
  AND2_X2 U4997 ( .A1(n6090), .A2(n6089), .ZN(n6094) );
  NAND3_X2 U4998 ( .A1(n9478), .A2(n9475), .A3(n5724), .ZN(n5757) );
  NAND2_X2 U4999 ( .A1(n9762), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5085) );
  NOR3_X2 U5000 ( .A1(n8286), .A2(n8285), .A3(n8284), .ZN(n8293) );
  INV_X1 U5001 ( .A(n5137), .ZN(n4434) );
  NAND2_X1 U5002 ( .A1(n9225), .A2(n9298), .ZN(n7156) );
  XNOR2_X2 U5003 ( .A(n5686), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9225) );
  INV_X1 U5004 ( .A(n5691), .ZN(n5716) );
  NAND2_X2 U5005 ( .A1(n6883), .A2(n6913), .ZN(n8188) );
  NAND2_X2 U5006 ( .A1(n5091), .A2(n7868), .ZN(n5346) );
  NAND2_X2 U5007 ( .A1(n5251), .A2(n5250), .ZN(n7387) );
  NAND2_X1 U5008 ( .A1(n4759), .A2(n9133), .ZN(n7323) );
  AOI21_X2 U5009 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n7607), .A(n7606), .ZN(
        n9388) );
  XNOR2_X2 U5010 ( .A(n4795), .B(n6484), .ZN(n6490) );
  NOR4_X2 U5011 ( .A1(n9230), .A2(n9106), .A3(n9105), .A4(n9104), .ZN(n9224)
         );
  NOR2_X2 U5012 ( .A1(n7414), .A2(n7413), .ZN(n7417) );
  NAND3_X2 U5013 ( .A1(n4479), .A2(n5094), .A3(n5093), .ZN(n5762) );
  AND2_X1 U5014 ( .A1(n4471), .A2(n4768), .ZN(n9721) );
  NAND2_X1 U5015 ( .A1(n9554), .A2(n9196), .ZN(n9529) );
  AOI21_X2 U5016 ( .B1(n8083), .B2(n8082), .A(n8081), .ZN(n8004) );
  OAI21_X1 U5017 ( .B1(n8971), .B2(n4621), .A(n4619), .ZN(n9019) );
  NAND2_X1 U5018 ( .A1(n7705), .A2(n8151), .ZN(n6205) );
  NAND2_X1 U5019 ( .A1(n6127), .A2(n8217), .ZN(n7245) );
  OR2_X1 U5020 ( .A1(n6341), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6352) );
  OR2_X1 U5021 ( .A1(n6334), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6341) );
  BUF_X1 U5022 ( .A(n5307), .Z(n4558) );
  NAND2_X1 U5023 ( .A1(n8188), .A2(n8186), .ZN(n8192) );
  NAND2_X1 U5024 ( .A1(n8211), .A2(n8205), .ZN(n8306) );
  NAND2_X1 U5025 ( .A1(n4442), .A2(n10006), .ZN(n8198) );
  NAND2_X1 U5026 ( .A1(n9243), .A2(n9249), .ZN(n9083) );
  OR2_X1 U5027 ( .A1(n6266), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6280) );
  BUF_X1 U5028 ( .A(n6292), .Z(n4440) );
  INV_X1 U5029 ( .A(n6882), .ZN(n6913) );
  NAND2_X1 U5030 ( .A1(n6065), .A2(n6050), .ZN(n6292) );
  AND4_X1 U5031 ( .A1(n5233), .A2(n5232), .A3(n5231), .A4(n5230), .ZN(n7623)
         );
  CLKBUF_X1 U5032 ( .A(n5762), .Z(n9323) );
  CLKBUF_X2 U5033 ( .A(n5471), .Z(n6670) );
  INV_X1 U5035 ( .A(n5137), .ZN(n5434) );
  CLKBUF_X3 U5036 ( .A(n8525), .Z(n4438) );
  INV_X2 U5037 ( .A(n5585), .ZN(n4437) );
  XNOR2_X1 U5038 ( .A(n5087), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5092) );
  NAND3_X1 U5039 ( .A1(n6085), .A2(n4774), .A3(n4772), .ZN(n6737) );
  OR2_X1 U5040 ( .A1(n6532), .A2(n6533), .ZN(n6535) );
  OR2_X1 U5041 ( .A1(n6532), .A2(n10062), .ZN(n6519) );
  AND2_X1 U5042 ( .A1(n4726), .A2(n6480), .ZN(n5000) );
  OAI21_X1 U5043 ( .B1(n8096), .B2(n8095), .A(n8094), .ZN(n8097) );
  OR2_X1 U5044 ( .A1(n7964), .A2(n7685), .ZN(n4726) );
  AND2_X1 U5045 ( .A1(n4770), .A2(n4769), .ZN(n4768) );
  XNOR2_X1 U5046 ( .A(n8136), .B(n8279), .ZN(n7964) );
  AND2_X1 U5047 ( .A1(n9630), .A2(n9633), .ZN(n9713) );
  AOI21_X1 U5048 ( .B1(n8555), .B2(n8731), .A(n8554), .ZN(n8818) );
  AOI21_X1 U5049 ( .B1(n4428), .B2(n6469), .A(n6468), .ZN(n8551) );
  NAND2_X1 U5050 ( .A1(n4716), .A2(n4715), .ZN(n8562) );
  NAND2_X1 U5051 ( .A1(n4545), .A2(n4544), .ZN(n4833) );
  NAND2_X1 U5052 ( .A1(n8135), .A2(n8134), .ZN(n8756) );
  NAND2_X1 U5053 ( .A1(n4981), .A2(n4982), .ZN(n8920) );
  NAND2_X1 U5054 ( .A1(n9056), .A2(n9055), .ZN(n9719) );
  NAND2_X1 U5055 ( .A1(n8126), .A2(n8125), .ZN(n8758) );
  XNOR2_X1 U5056 ( .A(n8132), .B(n8131), .ZN(n9765) );
  OAI21_X1 U5057 ( .B1(n8129), .B2(n8128), .A(n8127), .ZN(n8132) );
  AOI21_X1 U5058 ( .B1(n5004), .B2(n5005), .A(n4513), .ZN(n5003) );
  OAI21_X2 U5059 ( .B1(n8004), .B2(n8006), .A(n8005), .ZN(n8063) );
  XNOR2_X1 U5060 ( .A(n8121), .B(SI_29_), .ZN(n7866) );
  AOI21_X1 U5061 ( .B1(n4452), .B2(n5049), .A(n4506), .ZN(n5048) );
  OAI21_X1 U5062 ( .B1(n6456), .B2(n6455), .A(n8629), .ZN(n8613) );
  NOR2_X1 U5063 ( .A1(n8476), .A2(n8693), .ZN(n8503) );
  AND2_X1 U5064 ( .A1(n5648), .A2(n5647), .ZN(n5663) );
  NAND2_X1 U5065 ( .A1(n4823), .A2(n4822), .ZN(n8032) );
  AOI21_X1 U5066 ( .B1(n8725), .B2(n6447), .A(n6446), .ZN(n8712) );
  NAND2_X1 U5067 ( .A1(n4792), .A2(n4791), .ZN(n4790) );
  NAND2_X1 U5068 ( .A1(n6349), .A2(n6348), .ZN(n8843) );
  OR2_X1 U5069 ( .A1(n8412), .A2(n8413), .ZN(n4565) );
  XNOR2_X1 U5070 ( .A(n4562), .B(n8414), .ZN(n8431) );
  OAI21_X1 U5071 ( .B1(n7707), .B2(n5025), .A(n5023), .ZN(n6442) );
  AOI21_X1 U5072 ( .B1(n5593), .B2(n5592), .A(n4559), .ZN(n5609) );
  NAND2_X1 U5073 ( .A1(n5560), .A2(n5559), .ZN(n5593) );
  NAND2_X1 U5074 ( .A1(n5552), .A2(n5551), .ZN(n5560) );
  NAND2_X1 U5075 ( .A1(n5467), .A2(n5466), .ZN(n9609) );
  INV_X1 U5076 ( .A(n9093), .ZN(n7732) );
  AOI21_X1 U5077 ( .B1(n9094), .B2(n5439), .A(n4459), .ZN(n4935) );
  NAND2_X1 U5078 ( .A1(n6155), .A2(n8153), .ZN(n7651) );
  NAND2_X1 U5079 ( .A1(n7501), .A2(n5351), .ZN(n7500) );
  NAND2_X1 U5080 ( .A1(n5447), .A2(n5446), .ZN(n9709) );
  NAND2_X1 U5081 ( .A1(n5404), .A2(n5403), .ZN(n9151) );
  OR2_X1 U5082 ( .A1(n5460), .A2(n4877), .ZN(n4872) );
  NAND2_X1 U5083 ( .A1(n7061), .A2(n7060), .ZN(n7200) );
  OAI21_X1 U5084 ( .B1(n5442), .B2(n5441), .A(n5440), .ZN(n5460) );
  NAND2_X1 U5085 ( .A1(n5383), .A2(n5382), .ZN(n9956) );
  AND2_X1 U5086 ( .A1(n9251), .A2(n9794), .ZN(n9086) );
  XNOR2_X1 U5087 ( .A(n10054), .B(n8344), .ZN(n8151) );
  NAND2_X1 U5088 ( .A1(n5319), .A2(n5318), .ZN(n9802) );
  AOI21_X1 U5089 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n7029), .A(n7025), .ZN(
        n7028) );
  NAND3_X1 U5090 ( .A1(n7992), .A2(n7991), .A3(n7009), .ZN(n7995) );
  OR2_X1 U5091 ( .A1(n7387), .A2(n9810), .ZN(n9136) );
  INV_X1 U5092 ( .A(n8306), .ZN(n6961) );
  NAND2_X1 U5093 ( .A1(n6088), .A2(n6887), .ZN(n8197) );
  NAND2_X1 U5094 ( .A1(n5225), .A2(n5224), .ZN(n9904) );
  XNOR2_X1 U5095 ( .A(n5288), .B(n5065), .ZN(n6574) );
  NAND2_X2 U5096 ( .A1(n6932), .A2(n8745), .ZN(n8748) );
  AND2_X1 U5097 ( .A1(n5202), .A2(n5201), .ZN(n9899) );
  NAND4_X2 U5098 ( .A1(n6108), .A2(n6107), .A3(n6106), .A4(n6105), .ZN(n7998)
         );
  NOR2_X2 U5099 ( .A1(n9857), .A2(n7132), .ZN(n7133) );
  NAND4_X2 U5100 ( .A1(n6055), .A2(n6054), .A3(n6053), .A4(n6052), .ZN(n8353)
         );
  OR2_X1 U5101 ( .A1(n9321), .A2(n5806), .ZN(n9243) );
  INV_X2 U5102 ( .A(n7938), .ZN(n7943) );
  XNOR2_X1 U5103 ( .A(n5766), .B(n5979), .ZN(n5777) );
  OAI21_X1 U5104 ( .B1(n6976), .B2(n6977), .A(n6975), .ZN(n7084) );
  NAND2_X1 U5105 ( .A1(n4871), .A2(n5217), .ZN(n5238) );
  CLKBUF_X2 U5106 ( .A(n6292), .Z(n4439) );
  INV_X1 U5107 ( .A(n7007), .ZN(n7938) );
  OR2_X1 U5108 ( .A1(n6091), .A2(n6997), .ZN(n6054) );
  AND3_X1 U5109 ( .A1(n6114), .A2(n6113), .A3(n6112), .ZN(n7003) );
  AND3_X1 U5110 ( .A1(n6100), .A2(n6099), .A3(n6098), .ZN(n7008) );
  CLKBUF_X3 U5111 ( .A(n6091), .Z(n4441) );
  OR2_X1 U5112 ( .A1(n6241), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6264) );
  NOR2_X1 U5113 ( .A1(n6855), .A2(n6845), .ZN(n6979) );
  NAND2_X2 U5114 ( .A1(n6879), .A2(n6878), .ZN(n7007) );
  AND4_X1 U5115 ( .A1(n5260), .A2(n5259), .A3(n5258), .A4(n5257), .ZN(n9810)
         );
  OR2_X1 U5116 ( .A1(n6492), .A2(P2_D_REG_0__SCAN_IN), .ZN(n4832) );
  NAND4_X1 U5117 ( .A1(n5141), .A2(n5140), .A3(n5139), .A4(n5138), .ZN(n9322)
         );
  INV_X2 U5118 ( .A(n6074), .ZN(n6646) );
  INV_X8 U5119 ( .A(n5966), .ZN(n5984) );
  NAND2_X1 U5120 ( .A1(n8893), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U5121 ( .A1(n6742), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6793) );
  AND2_X1 U5122 ( .A1(n6624), .A2(n6876), .ZN(n4831) );
  NAND2_X2 U5123 ( .A1(n4970), .A2(n5765), .ZN(n5979) );
  INV_X1 U5124 ( .A(n5116), .ZN(n5137) );
  INV_X2 U5125 ( .A(n5585), .ZN(n5135) );
  NAND2_X2 U5126 ( .A1(n5092), .A2(n9767), .ZN(n5471) );
  OR2_X1 U5127 ( .A1(n6199), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6218) );
  AOI21_X1 U5128 ( .B1(n4876), .B2(n4879), .A(n4875), .ZN(n4874) );
  NAND2_X1 U5129 ( .A1(n6045), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6047) );
  OR2_X2 U5130 ( .A1(n5091), .A2(n5092), .ZN(n5585) );
  INV_X1 U5131 ( .A(n6491), .ZN(n7828) );
  XNOR2_X1 U5132 ( .A(n4793), .B(P2_IR_REG_25__SCAN_IN), .ZN(n7758) );
  MUX2_X1 U5133 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6057), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n6059) );
  INV_X1 U5134 ( .A(n7359), .ZN(n8194) );
  AOI21_X1 U5135 ( .B1(n4661), .B2(n4659), .A(n4658), .ZN(n4657) );
  OR2_X1 U5136 ( .A1(n6188), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6199) );
  AND2_X1 U5137 ( .A1(n6488), .A2(n6487), .ZN(n6491) );
  XNOR2_X1 U5138 ( .A(n6415), .B(n6414), .ZN(n7359) );
  NAND2_X1 U5139 ( .A1(n4839), .A2(n4838), .ZN(n5097) );
  NAND2_X1 U5140 ( .A1(n6483), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4795) );
  NAND2_X1 U5141 ( .A1(n5690), .A2(n5689), .ZN(n9298) );
  NAND2_X1 U5142 ( .A1(n5689), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U5143 ( .A1(n6418), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6415) );
  OR2_X1 U5144 ( .A1(n5086), .A2(n5198), .ZN(n5087) );
  NAND2_X1 U5145 ( .A1(n5445), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5465) );
  INV_X2 U5146 ( .A(n9764), .ZN(n9769) );
  NOR2_X1 U5147 ( .A1(n5494), .A2(SI_19_), .ZN(n4875) );
  NAND2_X1 U5148 ( .A1(n6038), .A2(n6037), .ZN(n6482) );
  XNOR2_X1 U5149 ( .A(n5124), .B(SI_1_), .ZN(n5121) );
  AND2_X1 U5150 ( .A1(n4523), .A2(n6041), .ZN(n5051) );
  NAND2_X2 U5151 ( .A1(n6549), .A2(P1_U3086), .ZN(n9771) );
  AND2_X1 U5152 ( .A1(n4485), .A2(n6084), .ZN(n6163) );
  AND4_X1 U5153 ( .A1(n6035), .A2(n6034), .A3(n6033), .A4(n6032), .ZN(n4448)
         );
  AND3_X1 U5154 ( .A1(n6248), .A2(n6031), .A3(n6272), .ZN(n6035) );
  NAND2_X1 U5155 ( .A1(n5083), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4838) );
  NAND3_X1 U5156 ( .A1(n4894), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4893) );
  NAND2_X1 U5157 ( .A1(n6178), .A2(n5057), .ZN(n5056) );
  INV_X1 U5158 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5680) );
  NOR2_X1 U5159 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6033) );
  INV_X1 U5160 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5188) );
  INV_X1 U5161 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5293) );
  INV_X2 U5162 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9333) );
  INV_X1 U5163 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4573) );
  INV_X1 U5164 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6178) );
  NOR2_X1 U5165 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6032) );
  NOR2_X1 U5166 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4752) );
  NOR2_X1 U5167 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4754) );
  NOR2_X1 U5168 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4755) );
  NOR2_X1 U5169 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4753) );
  OR2_X2 U5170 ( .A1(n8351), .A2(n7008), .ZN(n8211) );
  AOI211_X2 U5171 ( .C1(n9652), .C2(n9887), .A(n9651), .B(n9650), .ZN(n9653)
         );
  OR2_X2 U5172 ( .A1(n7337), .A2(n7343), .ZN(n7335) );
  OAI21_X2 U5173 ( .B1(n6793), .B2(n4776), .A(n4775), .ZN(n6977) );
  AND2_X2 U5174 ( .A1(n5130), .A2(n4756), .ZN(n7300) );
  AOI21_X2 U5175 ( .B1(n4615), .B2(n4614), .A(n4613), .ZN(n4612) );
  OAI21_X2 U5176 ( .B1(n7245), .B2(n6141), .A(n8209), .ZN(n7445) );
  OAI21_X2 U5177 ( .B1(n7872), .B2(n5711), .A(n9113), .ZN(n9513) );
  OAI21_X2 U5178 ( .B1(n6205), .B2(n4750), .A(n4748), .ZN(n8735) );
  AOI21_X2 U5179 ( .B1(n5723), .B2(n9887), .A(n5722), .ZN(n9478) );
  OAI21_X2 U5180 ( .B1(n9529), .B2(n9100), .A(n9198), .ZN(n7872) );
  OAI21_X2 U5181 ( .B1(n9519), .B2(n9518), .A(n5627), .ZN(n9509) );
  OAI21_X2 U5182 ( .B1(n7651), .B2(n8154), .A(n8161), .ZN(n7674) );
  OR2_X1 U5183 ( .A1(n9080), .A2(n6945), .ZN(n7297) );
  OAI21_X2 U5184 ( .B1(n8697), .B2(n8227), .A(n8229), .ZN(n8690) );
  OAI21_X2 U5185 ( .B1(n5699), .B2(n4610), .A(n4612), .ZN(n9242) );
  CLKBUF_X1 U5186 ( .A(n6101), .Z(n4444) );
  BUF_X4 U5187 ( .A(n6101), .Z(n4445) );
  XNOR2_X2 U5188 ( .A(n6047), .B(n6046), .ZN(n6050) );
  NAND2_X1 U5189 ( .A1(n6059), .A2(n6058), .ZN(n8525) );
  NOR2_X1 U5190 ( .A1(n5264), .A2(n4662), .ZN(n4661) );
  INV_X1 U5191 ( .A(n5241), .ZN(n4662) );
  OAI21_X1 U5192 ( .B1(n6791), .B2(n6792), .A(n4564), .ZN(n4778) );
  OR2_X1 U5193 ( .A1(n8859), .A2(n8649), .ZN(n8254) );
  NAND2_X1 U5194 ( .A1(n4918), .A2(n4917), .ZN(n8411) );
  INV_X1 U5195 ( .A(n8384), .ZN(n4917) );
  NOR2_X1 U5196 ( .A1(n8431), .A2(n8432), .ZN(n8454) );
  AOI21_X1 U5197 ( .B1(n5020), .B2(n5018), .A(n4507), .ZN(n5017) );
  INV_X1 U5198 ( .A(n6469), .ZN(n5018) );
  INV_X1 U5199 ( .A(n6039), .ZN(n5053) );
  INV_X1 U5200 ( .A(n5527), .ZN(n5528) );
  NAND2_X1 U5201 ( .A1(n7925), .A2(n8061), .ZN(n4806) );
  OR2_X1 U5202 ( .A1(n6520), .A2(n8553), .ZN(n8291) );
  NAND2_X1 U5203 ( .A1(n8291), .A2(n8140), .ZN(n8284) );
  AOI21_X1 U5204 ( .B1(n4657), .B2(n4660), .A(n4655), .ZN(n4654) );
  NAND2_X1 U5205 ( .A1(n8197), .A2(n8198), .ZN(n6426) );
  NAND2_X1 U5206 ( .A1(n8298), .A2(n8265), .ZN(n4725) );
  OR2_X1 U5207 ( .A1(n8879), .A2(n8111), .ZN(n8232) );
  INV_X1 U5208 ( .A(n4447), .ZN(n4633) );
  OAI21_X1 U5209 ( .B1(n4633), .B2(n4631), .A(n4972), .ZN(n4630) );
  OR2_X1 U5210 ( .A1(n4476), .A2(n7693), .ZN(n4631) );
  AOI21_X1 U5211 ( .B1(n4447), .B2(n4975), .A(n4973), .ZN(n4972) );
  NAND2_X1 U5212 ( .A1(n4623), .A2(n4622), .ZN(n5890) );
  NAND2_X1 U5213 ( .A1(n5885), .A2(n8907), .ZN(n4622) );
  NAND2_X1 U5214 ( .A1(n7791), .A2(n4495), .ZN(n4623) );
  OR2_X1 U5215 ( .A1(n9956), .A2(n7829), .ZN(n9262) );
  INV_X1 U5216 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5082) );
  INV_X1 U5217 ( .A(n5081), .ZN(n4957) );
  NAND2_X1 U5218 ( .A1(n4890), .A2(n4888), .ZN(n5552) );
  NOR2_X1 U5219 ( .A1(n5536), .A2(n4889), .ZN(n4888) );
  INV_X1 U5220 ( .A(n5529), .ZN(n4889) );
  XNOR2_X1 U5221 ( .A(n5494), .B(SI_19_), .ZN(n5495) );
  NOR2_X1 U5222 ( .A1(n5462), .A2(n4882), .ZN(n4881) );
  INV_X1 U5223 ( .A(n4884), .ZN(n4882) );
  AND2_X1 U5224 ( .A1(n5444), .A2(n4618), .ZN(n5682) );
  INV_X1 U5225 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4618) );
  XNOR2_X1 U5226 ( .A(n5458), .B(SI_17_), .ZN(n5459) );
  INV_X1 U5227 ( .A(n5418), .ZN(n5419) );
  OAI21_X1 U5228 ( .B1(n7944), .B2(n4818), .A(n4815), .ZN(n4814) );
  NAND2_X1 U5229 ( .A1(n4816), .A2(n4818), .ZN(n4815) );
  OR2_X1 U5230 ( .A1(n7944), .A2(n7967), .ZN(n4816) );
  INV_X1 U5231 ( .A(n4441), .ZN(n6405) );
  NAND2_X1 U5232 ( .A1(n6852), .A2(n6790), .ZN(n4563) );
  NOR2_X1 U5233 ( .A1(n8375), .A2(n8365), .ZN(n8381) );
  AND2_X1 U5234 ( .A1(n8411), .A2(n8410), .ZN(n8438) );
  INV_X1 U5235 ( .A(n8457), .ZN(n4791) );
  NAND2_X1 U5236 ( .A1(n4908), .A2(n4907), .ZN(n4906) );
  INV_X1 U5237 ( .A(n8441), .ZN(n4907) );
  OR2_X1 U5238 ( .A1(n6394), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n7958) );
  AND2_X1 U5239 ( .A1(n8843), .A2(n8583), .ZN(n8298) );
  NAND2_X1 U5240 ( .A1(n6362), .A2(n6361), .ZN(n6374) );
  INV_X1 U5241 ( .A(n6363), .ZN(n6362) );
  INV_X1 U5242 ( .A(n8342), .ZN(n8594) );
  OR2_X1 U5243 ( .A1(n8872), .A2(n8659), .ZN(n8249) );
  AOI21_X1 U5244 ( .B1(n5024), .B2(n6440), .A(n4531), .ZN(n5023) );
  OR2_X1 U5245 ( .A1(n10060), .A2(n8741), .ZN(n8179) );
  AND2_X1 U5246 ( .A1(n4696), .A2(n4702), .ZN(n4695) );
  NAND2_X1 U5247 ( .A1(n4703), .A2(n5353), .ZN(n4702) );
  NAND2_X1 U5248 ( .A1(n4700), .A2(n4697), .ZN(n4696) );
  INV_X1 U5249 ( .A(n4705), .ZN(n4703) );
  AOI21_X1 U5250 ( .B1(n8315), .B2(n8156), .A(n4713), .ZN(n4712) );
  INV_X1 U5251 ( .A(n8163), .ZN(n4713) );
  INV_X1 U5252 ( .A(n8341), .ZN(n8574) );
  NAND2_X1 U5253 ( .A1(n6338), .A2(n8262), .ZN(n8602) );
  INV_X1 U5254 ( .A(n8133), .ZN(n6301) );
  NAND2_X1 U5255 ( .A1(n4438), .A2(n4737), .ZN(n4739) );
  AND2_X1 U5256 ( .A1(n6472), .A2(n9995), .ZN(n4737) );
  AOI21_X1 U5257 ( .B1(n4438), .B2(n6472), .A(n4741), .ZN(n4738) );
  OR2_X1 U5258 ( .A1(n6060), .A2(n4436), .ZN(n4741) );
  INV_X1 U5259 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4552) );
  INV_X1 U5260 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4551) );
  NAND2_X1 U5261 ( .A1(n7949), .A2(n7950), .ZN(n4992) );
  XNOR2_X1 U5262 ( .A(n5836), .B(n5837), .ZN(n7621) );
  NAND2_X1 U5263 ( .A1(n4648), .A2(n5962), .ZN(n4647) );
  AND2_X1 U5264 ( .A1(n5548), .A2(n5547), .ZN(n9058) );
  OAI21_X1 U5265 ( .B1(n9543), .B2(n4939), .A(n4937), .ZN(n9519) );
  NAND2_X1 U5266 ( .A1(n4940), .A2(n4472), .ZN(n4939) );
  AOI21_X1 U5267 ( .B1(n4519), .B2(n4940), .A(n4938), .ZN(n4937) );
  NOR2_X1 U5268 ( .A1(n7879), .A2(n8994), .ZN(n4938) );
  INV_X1 U5269 ( .A(n9543), .ZN(n4945) );
  OR2_X1 U5270 ( .A1(n7527), .A2(n9793), .ZN(n9163) );
  NAND2_X1 U5271 ( .A1(n7500), .A2(n4763), .ZN(n7662) );
  NOR2_X1 U5272 ( .A1(n9091), .A2(n4764), .ZN(n4763) );
  INV_X1 U5273 ( .A(n9163), .ZN(n4764) );
  NOR2_X1 U5274 ( .A1(n5338), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5377) );
  INV_X1 U5275 ( .A(n8535), .ZN(n10406) );
  AND2_X1 U5276 ( .A1(n8167), .A2(n8176), .ZN(n8218) );
  AOI21_X1 U5277 ( .B1(n4612), .B2(n4610), .A(n9219), .ZN(n4608) );
  NAND2_X1 U5278 ( .A1(n8223), .A2(n8224), .ZN(n4690) );
  NAND2_X1 U5279 ( .A1(n8736), .A2(n4503), .ZN(n4687) );
  NOR2_X1 U5280 ( .A1(n8727), .A2(n8317), .ZN(n4691) );
  INV_X1 U5281 ( .A(n9264), .ZN(n4605) );
  INV_X1 U5282 ( .A(n9257), .ZN(n4604) );
  NOR2_X1 U5283 ( .A1(n9259), .A2(n4601), .ZN(n4600) );
  NAND2_X1 U5284 ( .A1(n9261), .A2(n9251), .ZN(n4601) );
  NOR2_X1 U5285 ( .A1(n4602), .A2(n4599), .ZN(n4598) );
  INV_X1 U5286 ( .A(n9261), .ZN(n4599) );
  AOI21_X1 U5287 ( .B1(n4606), .B2(n9254), .A(n4603), .ZN(n4602) );
  INV_X1 U5288 ( .A(n9258), .ZN(n4603) );
  OAI21_X1 U5289 ( .B1(n9175), .B2(n4583), .A(n9174), .ZN(n9187) );
  OAI21_X1 U5290 ( .B1(n9154), .B2(n9217), .A(n4582), .ZN(n4583) );
  AOI21_X1 U5291 ( .B1(n8256), .B2(n8259), .A(n8255), .ZN(n4685) );
  INV_X1 U5292 ( .A(n4684), .ZN(n4683) );
  OAI21_X1 U5293 ( .B1(n8257), .B2(n8292), .A(n8615), .ZN(n4684) );
  NAND2_X1 U5294 ( .A1(n8300), .A2(n8262), .ZN(n4679) );
  NAND2_X1 U5295 ( .A1(n8267), .A2(n4863), .ZN(n4862) );
  INV_X1 U5296 ( .A(n4474), .ZN(n4863) );
  NAND2_X1 U5297 ( .A1(n8263), .A2(n8292), .ZN(n4681) );
  NOR2_X1 U5298 ( .A1(n8611), .A2(n4732), .ZN(n8322) );
  NAND2_X1 U5299 ( .A1(n4866), .A2(n8270), .ZN(n4865) );
  NAND2_X1 U5300 ( .A1(n4861), .A2(n4488), .ZN(n4866) );
  INV_X1 U5301 ( .A(n8273), .ZN(n4858) );
  INV_X1 U5302 ( .A(n4640), .ZN(n4639) );
  OAI21_X1 U5303 ( .B1(n5826), .B2(n4450), .A(n7349), .ZN(n4640) );
  AND2_X1 U5304 ( .A1(n5826), .A2(n4450), .ZN(n4638) );
  NAND2_X1 U5305 ( .A1(n4589), .A2(n9217), .ZN(n4588) );
  AND2_X1 U5306 ( .A1(n9676), .A2(n9681), .ZN(n9181) );
  NOR2_X2 U5307 ( .A1(n4765), .A2(n9246), .ZN(n4615) );
  NOR2_X1 U5308 ( .A1(n5332), .A2(n4709), .ZN(n4708) );
  INV_X1 U5309 ( .A(n5310), .ZN(n4709) );
  NAND2_X1 U5310 ( .A1(n5268), .A2(n5267), .ZN(n5289) );
  AOI21_X1 U5311 ( .B1(n4804), .B2(n4803), .A(n4802), .ZN(n4801) );
  INV_X1 U5312 ( .A(n4807), .ZN(n4803) );
  NOR2_X1 U5313 ( .A1(n8329), .A2(n8328), .ZN(n8330) );
  AND2_X1 U5314 ( .A1(n4896), .A2(n4543), .ZN(n4542) );
  OR2_X1 U5315 ( .A1(n8817), .A2(n8756), .ZN(n4543) );
  INV_X1 U5316 ( .A(n8333), .ZN(n4896) );
  NAND2_X1 U5317 ( .A1(n10415), .A2(n6726), .ZN(n6727) );
  AND2_X1 U5318 ( .A1(n8788), .A2(n8648), .ZN(n6453) );
  AOI21_X1 U5319 ( .B1(n4710), .B2(n4708), .A(n4706), .ZN(n4705) );
  INV_X1 U5320 ( .A(n5331), .ZN(n4706) );
  AND2_X1 U5321 ( .A1(n8826), .A2(n8574), .ZN(n8275) );
  NOR2_X1 U5322 ( .A1(n5050), .A2(n6467), .ZN(n5049) );
  INV_X1 U5323 ( .A(n6466), .ZN(n5050) );
  OR2_X1 U5324 ( .A1(n8826), .A2(n8574), .ZN(n8272) );
  OR2_X1 U5325 ( .A1(n8585), .A2(n8594), .ZN(n8269) );
  NAND2_X1 U5326 ( .A1(n5067), .A2(n5035), .ZN(n5034) );
  INV_X1 U5327 ( .A(n5036), .ZN(n5035) );
  INV_X1 U5328 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5057) );
  NOR2_X1 U5329 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n6030) );
  INV_X1 U5330 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6029) );
  INV_X1 U5331 ( .A(n5846), .ZN(n4976) );
  NAND2_X1 U5332 ( .A1(n4983), .A2(n4481), .ZN(n4982) );
  INV_X1 U5333 ( .A(n8940), .ZN(n4983) );
  AND2_X1 U5334 ( .A1(n4481), .A2(n5935), .ZN(n4984) );
  AND2_X1 U5335 ( .A1(n5769), .A2(n5770), .ZN(n5775) );
  AND2_X1 U5336 ( .A1(n6539), .A2(n7156), .ZN(n4970) );
  NAND2_X2 U5337 ( .A1(n5761), .A2(n6539), .ZN(n5966) );
  AOI21_X1 U5338 ( .B1(n9719), .B2(n9219), .A(n4466), .ZN(n4555) );
  NAND2_X1 U5339 ( .A1(n4586), .A2(n4585), .ZN(n9221) );
  OR2_X1 U5340 ( .A1(n9719), .A2(n9217), .ZN(n4585) );
  NAND2_X1 U5341 ( .A1(n9218), .A2(n9719), .ZN(n4586) );
  INV_X1 U5342 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5073) );
  INV_X1 U5343 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5074) );
  INV_X1 U5344 ( .A(n9210), .ZN(n9201) );
  OR2_X1 U5345 ( .A1(n5580), .A2(n5579), .ZN(n5601) );
  OR2_X1 U5346 ( .A1(n9540), .A2(n9648), .ZN(n9198) );
  INV_X1 U5347 ( .A(n9123), .ZN(n4762) );
  OR2_X1 U5348 ( .A1(n7813), .A2(n9622), .ZN(n9268) );
  NAND2_X1 U5349 ( .A1(n5351), .A2(n5352), .ZN(n4953) );
  INV_X1 U5350 ( .A(n5352), .ZN(n4950) );
  NAND2_X1 U5351 ( .A1(n5668), .A2(n5667), .ZN(n8118) );
  NAND2_X1 U5352 ( .A1(n5663), .A2(n5662), .ZN(n5668) );
  XNOR2_X1 U5353 ( .A(n8118), .B(n8117), .ZN(n8121) );
  NAND2_X1 U5354 ( .A1(n4524), .A2(n5083), .ZN(n4956) );
  INV_X1 U5355 ( .A(n5594), .ZN(n4559) );
  INV_X1 U5356 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5736) );
  INV_X1 U5357 ( .A(n5370), .ZN(n5371) );
  INV_X1 U5358 ( .A(n5263), .ZN(n4658) );
  INV_X1 U5359 ( .A(n5237), .ZN(n4659) );
  INV_X1 U5360 ( .A(n4661), .ZN(n4660) );
  AND3_X2 U5361 ( .A1(n4573), .A2(n9333), .A3(n5070), .ZN(n5072) );
  INV_X1 U5362 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5070) );
  NAND2_X2 U5363 ( .A1(n4895), .A2(n4893), .ZN(n5126) );
  NAND3_X1 U5364 ( .A1(n8531), .A2(n4652), .A3(n4651), .ZN(n4895) );
  INV_X1 U5365 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4651) );
  INV_X1 U5366 ( .A(n7931), .ZN(n4544) );
  INV_X1 U5367 ( .A(n7932), .ZN(n4545) );
  NAND2_X1 U5368 ( .A1(n7200), .A2(n4499), .ZN(n7286) );
  NOR2_X1 U5369 ( .A1(n8014), .A2(n4808), .ZN(n4807) );
  INV_X1 U5370 ( .A(n8062), .ZN(n4808) );
  AND2_X1 U5371 ( .A1(n8072), .A2(n7928), .ZN(n8013) );
  INV_X1 U5372 ( .A(n8729), .ZN(n8302) );
  INV_X1 U5373 ( .A(n4825), .ZN(n4824) );
  XNOR2_X1 U5374 ( .A(n8351), .B(n7010), .ZN(n7993) );
  NAND2_X1 U5375 ( .A1(n8106), .A2(n4826), .ZN(n4825) );
  INV_X1 U5376 ( .A(n4827), .ZN(n4826) );
  OR2_X1 U5377 ( .A1(n4439), .A2(n6934), .ZN(n6068) );
  OR2_X1 U5378 ( .A1(n4445), .A2(n6655), .ZN(n6069) );
  OAI21_X1 U5379 ( .B1(n6793), .B2(n6792), .A(n4517), .ZN(n4779) );
  INV_X1 U5380 ( .A(n6977), .ZN(n4780) );
  OR2_X1 U5381 ( .A1(n7178), .A2(n7070), .ZN(n4786) );
  NAND2_X1 U5382 ( .A1(n4785), .A2(n4784), .ZN(n4783) );
  INV_X1 U5383 ( .A(n7178), .ZN(n4784) );
  INV_X1 U5384 ( .A(n4787), .ZN(n4785) );
  OR2_X1 U5385 ( .A1(n7085), .A2(n7070), .ZN(n4788) );
  INV_X1 U5386 ( .A(n7416), .ZN(n4912) );
  AOI21_X1 U5387 ( .B1(n8363), .B2(n8362), .A(n8361), .ZN(n8368) );
  NOR2_X1 U5388 ( .A1(n8444), .A2(n8443), .ZN(n8468) );
  NOR2_X1 U5389 ( .A1(n8503), .A2(n8504), .ZN(n8507) );
  NAND2_X1 U5390 ( .A1(n8279), .A2(n5020), .ZN(n5016) );
  OAI21_X1 U5391 ( .B1(n8279), .B2(n4491), .A(n5013), .ZN(n5012) );
  INV_X1 U5392 ( .A(n8576), .ZN(n8571) );
  NAND2_X1 U5393 ( .A1(n4522), .A2(n4451), .ZN(n5004) );
  NAND2_X1 U5394 ( .A1(n8615), .A2(n6461), .ZN(n5006) );
  NAND2_X1 U5395 ( .A1(n4451), .A2(n6461), .ZN(n5005) );
  NAND2_X1 U5396 ( .A1(n6326), .A2(n6325), .ZN(n6334) );
  INV_X1 U5397 ( .A(n6327), .ZN(n6326) );
  OR2_X1 U5398 ( .A1(n6290), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6305) );
  AND4_X1 U5399 ( .A1(n6296), .A2(n6295), .A3(n6294), .A4(n6293), .ZN(n8659)
         );
  INV_X1 U5400 ( .A(n5046), .ZN(n5042) );
  NOR2_X1 U5401 ( .A1(n8703), .A2(n5044), .ZN(n5043) );
  INV_X1 U5402 ( .A(n6448), .ZN(n5044) );
  NAND2_X1 U5403 ( .A1(n6229), .A2(n6228), .ZN(n6241) );
  NAND2_X1 U5404 ( .A1(n5028), .A2(n5027), .ZN(n5030) );
  NAND2_X1 U5405 ( .A1(n6170), .A2(n6169), .ZN(n6188) );
  INV_X1 U5406 ( .A(n6171), .ZN(n6170) );
  OR2_X1 U5407 ( .A1(n6182), .A2(n7677), .ZN(n6434) );
  AND2_X1 U5408 ( .A1(n8215), .A2(n8209), .ZN(n8310) );
  OR2_X1 U5409 ( .A1(n4999), .A2(n8306), .ZN(n4997) );
  INV_X1 U5410 ( .A(n7120), .ZN(n4999) );
  AOI21_X1 U5411 ( .B1(n4717), .B2(n4723), .A(n4489), .ZN(n4715) );
  AND2_X1 U5412 ( .A1(n4720), .A2(n4718), .ZN(n4717) );
  AOI21_X1 U5413 ( .B1(n4475), .B2(n4722), .A(n4721), .ZN(n4720) );
  INV_X1 U5414 ( .A(n8269), .ZN(n4721) );
  INV_X1 U5415 ( .A(n4475), .ZN(n4723) );
  OR2_X1 U5416 ( .A1(n8271), .A2(n4489), .ZN(n8576) );
  OR2_X1 U5417 ( .A1(n4722), .A2(n8298), .ZN(n8597) );
  NAND2_X1 U5418 ( .A1(n6457), .A2(n8611), .ZN(n8617) );
  NOR2_X1 U5419 ( .A1(n4732), .A2(n4731), .ZN(n4730) );
  NAND2_X1 U5420 ( .A1(n6888), .A2(n8274), .ZN(n8744) );
  OR2_X1 U5421 ( .A1(n6888), .A2(n8292), .ZN(n8742) );
  INV_X1 U5422 ( .A(n8731), .ZN(n8740) );
  NAND2_X1 U5423 ( .A1(n4734), .A2(n8260), .ZN(n8641) );
  NAND2_X1 U5424 ( .A1(n8671), .A2(n4735), .ZN(n4734) );
  AND2_X1 U5425 ( .A1(n8232), .A2(n6449), .ZN(n8703) );
  NAND2_X1 U5426 ( .A1(n6263), .A2(n6262), .ZN(n8803) );
  INV_X1 U5427 ( .A(n8742), .ZN(n8726) );
  INV_X1 U5428 ( .A(n4749), .ZN(n4748) );
  OAI22_X1 U5429 ( .A1(n4751), .A2(n4750), .B1(n8727), .B2(n9774), .ZN(n4749)
         );
  NAND2_X1 U5430 ( .A1(n4516), .A2(n8179), .ZN(n4750) );
  NAND2_X1 U5431 ( .A1(n8137), .A2(n6509), .ZN(n8731) );
  NAND2_X1 U5432 ( .A1(n6487), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6057) );
  INV_X1 U5433 ( .A(n5056), .ZN(n5054) );
  CLKBUF_X1 U5434 ( .A(n6163), .Z(n6164) );
  OR2_X1 U5435 ( .A1(n7949), .A2(n7950), .ZN(n4993) );
  INV_X1 U5436 ( .A(n4982), .ZN(n4980) );
  AND2_X1 U5437 ( .A1(n4453), .A2(n4984), .ZN(n4979) );
  NAND2_X1 U5438 ( .A1(n6937), .A2(n4960), .ZN(n4958) );
  INV_X1 U5439 ( .A(n4630), .ZN(n4629) );
  NAND2_X1 U5440 ( .A1(n7692), .A2(n5846), .ZN(n7852) );
  NAND2_X1 U5441 ( .A1(n4645), .A2(n4644), .ZN(n9026) );
  AOI21_X1 U5442 ( .B1(n4454), .B2(n8989), .A(n4501), .ZN(n4644) );
  NAND2_X1 U5443 ( .A1(n5891), .A2(n5894), .ZN(n4963) );
  OR2_X1 U5444 ( .A1(n5890), .A2(n5889), .ZN(n5895) );
  NAND2_X1 U5445 ( .A1(n5764), .A2(n5765), .ZN(n4971) );
  NAND2_X1 U5446 ( .A1(n5135), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5110) );
  XOR2_X1 U5447 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6607), .Z(n9327) );
  NAND2_X1 U5448 ( .A1(n9520), .A2(n4842), .ZN(n9463) );
  NOR2_X1 U5449 ( .A1(n4843), .A2(n9719), .ZN(n4842) );
  INV_X1 U5450 ( .A(n4844), .ZN(n4843) );
  INV_X1 U5451 ( .A(n4932), .ZN(n4931) );
  OAI21_X1 U5452 ( .B1(n9508), .B2(n4933), .A(n5661), .ZN(n4932) );
  INV_X1 U5453 ( .A(n5642), .ZN(n4933) );
  AND2_X1 U5454 ( .A1(n9214), .A2(n9215), .ZN(n9111) );
  AND2_X1 U5455 ( .A1(n9201), .A2(n9110), .ZN(n9485) );
  NAND2_X1 U5456 ( .A1(n9520), .A2(n9505), .ZN(n9500) );
  AND2_X1 U5457 ( .A1(n5652), .A2(n5621), .ZN(n9523) );
  AND2_X1 U5458 ( .A1(n9116), .A2(n9114), .ZN(n9518) );
  AOI21_X1 U5459 ( .B1(n4943), .B2(n4941), .A(n4510), .ZN(n4940) );
  INV_X1 U5460 ( .A(n4473), .ZN(n4941) );
  AND2_X1 U5461 ( .A1(n9198), .A2(n9205), .ZN(n9532) );
  NAND2_X2 U5462 ( .A1(n5550), .A2(n5549), .ZN(n9543) );
  NOR2_X1 U5463 ( .A1(n4533), .A2(n4925), .ZN(n4924) );
  NAND2_X1 U5464 ( .A1(n9572), .A2(n9571), .ZN(n9570) );
  OR2_X1 U5465 ( .A1(n5517), .A2(n5516), .ZN(n5541) );
  OR2_X1 U5466 ( .A1(n7901), .A2(n4762), .ZN(n7885) );
  AND2_X1 U5467 ( .A1(n9174), .A2(n9273), .ZN(n4771) );
  NAND2_X1 U5468 ( .A1(n7803), .A2(n9094), .ZN(n5705) );
  AND2_X1 U5469 ( .A1(n9262), .A2(n9264), .ZN(n9166) );
  NAND2_X1 U5470 ( .A1(n5360), .A2(n5359), .ZN(n7668) );
  OR2_X1 U5471 ( .A1(n5299), .A2(n10141), .ZN(n5322) );
  AND4_X1 U5472 ( .A1(n5350), .A2(n5349), .A3(n5348), .A4(n5347), .ZN(n9793)
         );
  NAND2_X1 U5473 ( .A1(n4836), .A2(n9899), .ZN(n9823) );
  NAND2_X1 U5474 ( .A1(n5498), .A2(n5497), .ZN(n7895) );
  INV_X1 U5475 ( .A(n9887), .ZN(n9933) );
  INV_X1 U5476 ( .A(n9952), .ZN(n9918) );
  INV_X1 U5477 ( .A(n9950), .ZN(n9891) );
  XNOR2_X1 U5478 ( .A(n5634), .B(n5633), .ZN(n7841) );
  INV_X1 U5479 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5079) );
  XNOR2_X1 U5480 ( .A(n5629), .B(n5628), .ZN(n7800) );
  XNOR2_X1 U5481 ( .A(n5576), .B(n5575), .ZN(n7703) );
  NAND2_X1 U5482 ( .A1(n4890), .A2(n5529), .ZN(n5537) );
  NAND2_X1 U5483 ( .A1(n5682), .A2(n5681), .ZN(n5687) );
  OR2_X1 U5484 ( .A1(n5687), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U5485 ( .A1(n4873), .A2(n4879), .ZN(n5496) );
  NAND2_X1 U5486 ( .A1(n5460), .A2(n4881), .ZN(n4873) );
  NAND2_X1 U5487 ( .A1(n4883), .A2(n4881), .ZN(n5479) );
  NAND2_X1 U5488 ( .A1(n4883), .A2(n4884), .ZN(n5463) );
  NAND2_X1 U5489 ( .A1(n4966), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U5490 ( .A1(n5465), .A2(n5679), .ZN(n4966) );
  AND2_X1 U5491 ( .A1(n9333), .A2(n4573), .ZN(n5104) );
  NOR2_X1 U5492 ( .A1(n4456), .A2(n8039), .ZN(n4810) );
  INV_X1 U5493 ( .A(n4818), .ZN(n4813) );
  NAND2_X1 U5494 ( .A1(n4814), .A2(n4817), .ZN(n4812) );
  NAND2_X1 U5495 ( .A1(n7944), .A2(n7967), .ZN(n4817) );
  INV_X1 U5496 ( .A(n8346), .ZN(n7292) );
  AND4_X1 U5497 ( .A1(n6322), .A2(n6321), .A3(n6320), .A4(n6319), .ZN(n8660)
         );
  AND2_X1 U5498 ( .A1(n6358), .A2(n6357), .ZN(n8583) );
  OR2_X1 U5499 ( .A1(n7753), .A2(n8345), .ZN(n4829) );
  AND2_X1 U5500 ( .A1(n7753), .A2(n8345), .ZN(n4828) );
  INV_X1 U5501 ( .A(n8343), .ZN(n8741) );
  AND2_X1 U5502 ( .A1(n6773), .A2(n6772), .ZN(n8037) );
  INV_X1 U5503 ( .A(n8713), .ZN(n8111) );
  OR2_X1 U5504 ( .A1(n4674), .A2(n8533), .ZN(n4671) );
  NAND2_X1 U5505 ( .A1(n4674), .A2(n4669), .ZN(n4668) );
  NOR2_X1 U5506 ( .A1(n8339), .A2(n8519), .ZN(n4669) );
  AND2_X1 U5507 ( .A1(n7217), .A2(n6412), .ZN(n8553) );
  NAND2_X1 U5508 ( .A1(n6400), .A2(n6399), .ZN(n8564) );
  NAND2_X1 U5509 ( .A1(n6391), .A2(n6390), .ZN(n8341) );
  NAND2_X1 U5510 ( .A1(n6371), .A2(n6370), .ZN(n8342) );
  INV_X1 U5511 ( .A(n8583), .ZN(n8605) );
  INV_X1 U5512 ( .A(n6123), .ZN(n6110) );
  INV_X1 U5513 ( .A(n4567), .ZN(n7412) );
  OR2_X1 U5514 ( .A1(n8381), .A2(n8382), .ZN(n4918) );
  NAND2_X1 U5515 ( .A1(n4565), .A2(n4477), .ZN(n4908) );
  INV_X1 U5516 ( .A(n4792), .ZN(n8458) );
  INV_X1 U5517 ( .A(n4790), .ZN(n8465) );
  INV_X1 U5518 ( .A(n4906), .ZN(n8474) );
  NOR2_X1 U5519 ( .A1(n8507), .A2(n8506), .ZN(n8518) );
  INV_X1 U5520 ( .A(n4561), .ZN(n8486) );
  NOR2_X1 U5521 ( .A1(n4920), .A2(n8508), .ZN(n4919) );
  AND2_X1 U5522 ( .A1(n8509), .A2(n8522), .ZN(n4920) );
  NAND2_X1 U5523 ( .A1(n6393), .A2(n6392), .ZN(n8558) );
  NAND2_X1 U5524 ( .A1(n6316), .A2(n6315), .ZN(n8653) );
  NAND2_X1 U5525 ( .A1(n6197), .A2(n6196), .ZN(n10054) );
  AND3_X1 U5526 ( .A1(n6154), .A2(n6153), .A3(n6152), .ZN(n7515) );
  NAND2_X1 U5527 ( .A1(n5733), .A2(n5754), .ZN(n6539) );
  NOR2_X1 U5528 ( .A1(n7802), .A2(n7704), .ZN(n5733) );
  OR2_X1 U5529 ( .A1(n4993), .A2(n9052), .ZN(n4991) );
  INV_X1 U5530 ( .A(n4992), .ZN(n4990) );
  NAND2_X1 U5531 ( .A1(n4647), .A2(n4646), .ZN(n8960) );
  AOI21_X1 U5532 ( .B1(n4460), .B2(n4992), .A(n9052), .ZN(n4989) );
  INV_X1 U5533 ( .A(n4988), .ZN(n4987) );
  OAI21_X1 U5534 ( .B1(n4991), .B2(n5973), .A(n4994), .ZN(n4988) );
  INV_X1 U5535 ( .A(n4995), .ZN(n4994) );
  OAI21_X1 U5536 ( .B1(n9505), .B2(n9039), .A(n7956), .ZN(n4995) );
  NAND2_X1 U5537 ( .A1(n5563), .A2(n5562), .ZN(n9665) );
  AND4_X1 U5538 ( .A1(n5369), .A2(n5368), .A3(n5367), .A4(n5366), .ZN(n9953)
         );
  OAI21_X1 U5539 ( .B1(n7692), .B2(n4975), .A(n4447), .ZN(n7788) );
  AND4_X1 U5540 ( .A1(n5390), .A2(n5389), .A3(n5388), .A4(n5387), .ZN(n7829)
         );
  INV_X1 U5541 ( .A(n9058), .ZN(n9555) );
  INV_X1 U5542 ( .A(n9691), .ZN(n9583) );
  INV_X1 U5543 ( .A(n9603), .ZN(n9781) );
  INV_X1 U5544 ( .A(n9951), .ZN(n9780) );
  NAND2_X1 U5545 ( .A1(n4965), .A2(n4964), .ZN(n5481) );
  AOI21_X1 U5546 ( .B1(n4967), .B2(n5198), .A(n5198), .ZN(n4964) );
  AND2_X1 U5547 ( .A1(n5571), .A2(n5570), .ZN(n9659) );
  NAND2_X1 U5548 ( .A1(n7384), .A2(n7158), .ZN(n9841) );
  INV_X1 U5549 ( .A(n7133), .ZN(n9618) );
  INV_X2 U5550 ( .A(n9598), .ZN(n9857) );
  NAND2_X1 U5551 ( .A1(n6584), .A2(n4849), .ZN(n4851) );
  OR2_X1 U5552 ( .A1(n4850), .A2(n4462), .ZN(n4849) );
  OR2_X1 U5553 ( .A1(n6002), .A2(n9304), .ZN(n9846) );
  NAND2_X1 U5554 ( .A1(n5341), .A2(n5340), .ZN(n7527) );
  AND2_X1 U5555 ( .A1(n9473), .A2(n9741), .ZN(n5756) );
  OAI21_X1 U5556 ( .B1(n5699), .B2(n4610), .A(n4609), .ZN(n4617) );
  OAI21_X1 U5557 ( .B1(n4688), .B2(n4689), .A(n4686), .ZN(n8231) );
  NAND2_X1 U5558 ( .A1(n4480), .A2(n4687), .ZN(n4686) );
  NAND2_X1 U5559 ( .A1(n8222), .A2(n4690), .ZN(n4689) );
  NOR2_X1 U5560 ( .A1(n4511), .A2(n4598), .ZN(n4597) );
  AOI21_X1 U5561 ( .B1(n9219), .B2(n4584), .A(n4520), .ZN(n4582) );
  NAND2_X1 U5562 ( .A1(n9169), .A2(n9273), .ZN(n4584) );
  NAND2_X1 U5563 ( .A1(n9187), .A2(n9270), .ZN(n9189) );
  AND3_X1 U5564 ( .A1(n8179), .A2(n8178), .A3(n8151), .ZN(n8176) );
  INV_X1 U5565 ( .A(n8176), .ZN(n8316) );
  INV_X1 U5566 ( .A(n7306), .ZN(n5696) );
  AND2_X1 U5567 ( .A1(n4575), .A2(n4482), .ZN(n9207) );
  AOI21_X1 U5568 ( .B1(n4581), .B2(n9184), .A(n9183), .ZN(n4580) );
  NAND2_X1 U5569 ( .A1(n4869), .A2(n4868), .ZN(n4859) );
  NAND2_X1 U5570 ( .A1(n8265), .A2(n8300), .ZN(n4869) );
  NAND2_X1 U5571 ( .A1(n4474), .A2(n4870), .ZN(n4860) );
  OR2_X1 U5572 ( .A1(n8298), .A2(n8264), .ZN(n4870) );
  INV_X1 U5573 ( .A(n8587), .ZN(n4867) );
  AND2_X1 U5574 ( .A1(n4862), .A2(n4681), .ZN(n4680) );
  OAI21_X1 U5575 ( .B1(n4500), .B2(n4679), .A(n8274), .ZN(n4678) );
  OAI21_X1 U5576 ( .B1(n4685), .B2(n8274), .A(n4683), .ZN(n4682) );
  OAI21_X1 U5577 ( .B1(n9203), .B2(n9208), .A(n9201), .ZN(n4591) );
  AOI21_X1 U5578 ( .B1(n8493), .B2(n8502), .A(n8492), .ZN(n8495) );
  INV_X1 U5579 ( .A(n5065), .ZN(n4655) );
  INV_X1 U5580 ( .A(n7620), .ZN(n4634) );
  NOR2_X1 U5581 ( .A1(n5885), .A2(n8907), .ZN(n4626) );
  INV_X1 U5582 ( .A(n5878), .ZN(n4624) );
  NAND2_X1 U5583 ( .A1(n4595), .A2(n4593), .ZN(n4592) );
  NOR2_X1 U5584 ( .A1(n9210), .A2(n4594), .ZN(n4593) );
  NAND2_X1 U5585 ( .A1(n9212), .A2(n9213), .ZN(n4595) );
  NAND2_X1 U5586 ( .A1(n9283), .A2(n9219), .ZN(n4594) );
  AND2_X1 U5587 ( .A1(n9723), .A2(n9497), .ZN(n9210) );
  INV_X1 U5588 ( .A(n9148), .ZN(n4546) );
  NOR2_X1 U5589 ( .A1(n9151), .A2(n9956), .ZN(n4854) );
  NAND2_X1 U5590 ( .A1(n4879), .A2(n4878), .ZN(n4877) );
  INV_X1 U5591 ( .A(n5495), .ZN(n4878) );
  NOR2_X1 U5592 ( .A1(n4881), .A2(n5495), .ZN(n4876) );
  NAND2_X1 U5593 ( .A1(n5313), .A2(n5312), .ZN(n5331) );
  AOI21_X1 U5594 ( .B1(n4865), .B2(n8571), .A(n4857), .ZN(n8278) );
  INV_X1 U5595 ( .A(n8272), .ZN(n8276) );
  NAND2_X1 U5596 ( .A1(n9987), .A2(n6736), .ZN(n10401) );
  INV_X1 U5597 ( .A(SI_15_), .ZN(n10232) );
  INV_X1 U5598 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6096) );
  INV_X1 U5599 ( .A(n4778), .ZN(n4777) );
  NAND2_X1 U5600 ( .A1(n4916), .A2(n4915), .ZN(n4914) );
  INV_X1 U5601 ( .A(n7185), .ZN(n4915) );
  NAND2_X1 U5602 ( .A1(n7542), .A2(n7541), .ZN(n7579) );
  INV_X1 U5603 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6248) );
  AND2_X1 U5604 ( .A1(n4906), .A2(n4905), .ZN(n8501) );
  NAND2_X1 U5605 ( .A1(n8475), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4905) );
  NAND2_X1 U5606 ( .A1(n8279), .A2(n5017), .ZN(n5013) );
  NOR2_X1 U5607 ( .A1(n8279), .A2(n5015), .ZN(n5014) );
  INV_X1 U5608 ( .A(n5017), .ZN(n5015) );
  INV_X1 U5609 ( .A(n4708), .ZN(n4697) );
  NAND2_X1 U5610 ( .A1(n8151), .A2(n5029), .ZN(n5026) );
  OR2_X1 U5611 ( .A1(n6433), .A2(n6432), .ZN(n7677) );
  OR2_X1 U5612 ( .A1(n6157), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U5613 ( .A1(n6143), .A2(n6142), .ZN(n6157) );
  INV_X1 U5614 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6142) );
  INV_X1 U5615 ( .A(n6144), .ZN(n6143) );
  INV_X1 U5616 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6115) );
  INV_X1 U5617 ( .A(n8271), .ZN(n4718) );
  INV_X1 U5618 ( .A(n8275), .ZN(n4864) );
  AND2_X1 U5619 ( .A1(n4735), .A2(n8246), .ZN(n4729) );
  NOR2_X1 U5620 ( .A1(n4733), .A2(n8260), .ZN(n4731) );
  NAND2_X1 U5621 ( .A1(n6460), .A2(n8633), .ZN(n8262) );
  NAND2_X1 U5622 ( .A1(n5067), .A2(n5033), .ZN(n5032) );
  AND2_X1 U5623 ( .A1(n8249), .A2(n4736), .ZN(n4735) );
  NAND2_X1 U5624 ( .A1(n5040), .A2(n5045), .ZN(n5036) );
  NOR2_X1 U5625 ( .A1(n5038), .A2(n6451), .ZN(n5033) );
  AOI21_X1 U5626 ( .B1(n5040), .B2(n5039), .A(n8685), .ZN(n5038) );
  INV_X1 U5627 ( .A(n5043), .ZN(n5039) );
  AND2_X1 U5628 ( .A1(n8152), .A2(n8177), .ZN(n4751) );
  INV_X1 U5629 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n10268) );
  INV_X1 U5630 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U5631 ( .A1(n5052), .A2(n4523), .ZN(n6487) );
  INV_X1 U5632 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6508) );
  NOR2_X1 U5633 ( .A1(n5227), .A2(n5226), .ZN(n5253) );
  NAND2_X1 U5634 ( .A1(n4636), .A2(n4635), .ZN(n5836) );
  NAND2_X1 U5635 ( .A1(n4639), .A2(n4450), .ZN(n4635) );
  OR2_X1 U5636 ( .A1(n4639), .A2(n4638), .ZN(n4637) );
  NOR2_X1 U5637 ( .A1(n4633), .A2(n4476), .ZN(n4632) );
  NOR2_X1 U5638 ( .A1(n5469), .A2(n5468), .ZN(n5486) );
  NAND2_X1 U5639 ( .A1(n5764), .A2(n4502), .ZN(n4969) );
  AND2_X1 U5640 ( .A1(n5405), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5430) );
  NOR2_X1 U5641 ( .A1(n5384), .A2(n10279), .ZN(n5405) );
  AND2_X1 U5642 ( .A1(n5618), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5654) );
  NOR2_X1 U5643 ( .A1(n9473), .A2(n4845), .ZN(n4844) );
  INV_X1 U5644 ( .A(n4846), .ZN(n4845) );
  NOR2_X1 U5645 ( .A1(n9488), .A2(n4847), .ZN(n4846) );
  INV_X1 U5646 ( .A(n5526), .ZN(n4925) );
  NOR2_X1 U5647 ( .A1(n5541), .A2(n9012), .ZN(n5564) );
  OR2_X1 U5648 ( .A1(n5499), .A2(n9003), .ZN(n5517) );
  NAND2_X1 U5649 ( .A1(n4854), .A2(n9784), .ZN(n4853) );
  NAND2_X1 U5650 ( .A1(n5430), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5449) );
  INV_X1 U5651 ( .A(n9153), .ZN(n9265) );
  AND2_X1 U5652 ( .A1(n9267), .A2(n9265), .ZN(n9093) );
  NOR2_X1 U5653 ( .A1(n5322), .A2(n5321), .ZN(n5343) );
  NAND2_X1 U5654 ( .A1(n9088), .A2(n4758), .ZN(n9255) );
  INV_X1 U5655 ( .A(n9087), .ZN(n4758) );
  INV_X1 U5656 ( .A(n9127), .ZN(n4613) );
  NAND2_X1 U5657 ( .A1(n7300), .A2(n4560), .ZN(n7301) );
  INV_X1 U5658 ( .A(n7302), .ZN(n4560) );
  NOR2_X1 U5659 ( .A1(n7718), .A2(n4852), .ZN(n7810) );
  INV_X1 U5660 ( .A(n4854), .ZN(n4852) );
  OR2_X1 U5661 ( .A1(n5685), .A2(n9233), .ZN(n5763) );
  AND2_X1 U5662 ( .A1(n5644), .A2(n5615), .ZN(n5628) );
  NOR2_X1 U5663 ( .A1(n5530), .A2(n4892), .ZN(n4891) );
  INV_X1 U5664 ( .A(n5511), .ZN(n4892) );
  AOI21_X1 U5665 ( .B1(n4881), .B2(n5459), .A(n4880), .ZN(n4879) );
  INV_X1 U5666 ( .A(n5478), .ZN(n4880) );
  OR2_X1 U5667 ( .A1(n5460), .A2(n5459), .ZN(n4883) );
  NAND2_X1 U5668 ( .A1(n4886), .A2(n4885), .ZN(n4884) );
  INV_X1 U5669 ( .A(SI_17_), .ZN(n4885) );
  XNOR2_X1 U5670 ( .A(n5373), .B(SI_13_), .ZN(n5370) );
  INV_X1 U5671 ( .A(n5306), .ZN(n4710) );
  AND2_X1 U5672 ( .A1(n5219), .A2(n5218), .ZN(n5221) );
  NAND2_X1 U5673 ( .A1(n5126), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5099) );
  AND2_X1 U5674 ( .A1(n4819), .A2(n4487), .ZN(n4818) );
  NAND2_X1 U5675 ( .A1(n7967), .A2(n4820), .ZN(n4819) );
  AND2_X1 U5676 ( .A1(n8022), .A2(n7935), .ZN(n8051) );
  XNOR2_X1 U5677 ( .A(n7008), .B(n7007), .ZN(n7010) );
  NAND2_X1 U5678 ( .A1(n7555), .A2(n7554), .ZN(n4821) );
  AOI21_X1 U5679 ( .B1(n4801), .B2(n4805), .A(n4798), .ZN(n4797) );
  INV_X1 U5680 ( .A(n8073), .ZN(n4798) );
  NAND2_X1 U5681 ( .A1(n4897), .A2(n8756), .ZN(n4673) );
  AOI21_X1 U5682 ( .B1(n8139), .B2(n4542), .A(n8330), .ZN(n4677) );
  NAND2_X1 U5683 ( .A1(n8331), .A2(n4675), .ZN(n4897) );
  NAND2_X1 U5684 ( .A1(n4676), .A2(n4675), .ZN(n4674) );
  NOR2_X1 U5685 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n6036) );
  OR2_X1 U5686 ( .A1(n9984), .A2(n6715), .ZN(n9987) );
  XNOR2_X1 U5687 ( .A(n6717), .B(n9995), .ZN(n9992) );
  INV_X1 U5688 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10221) );
  NAND2_X1 U5689 ( .A1(n6084), .A2(n6096), .ZN(n6123) );
  AND2_X1 U5690 ( .A1(n4901), .A2(n6786), .ZN(n4902) );
  AND2_X1 U5691 ( .A1(n6785), .A2(n6728), .ZN(n6729) );
  NAND2_X1 U5692 ( .A1(n6729), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6788) );
  OR2_X1 U5693 ( .A1(n6854), .A2(n6861), .ZN(n4550) );
  OAI21_X1 U5694 ( .B1(n6979), .B2(n4904), .A(n6980), .ZN(n7077) );
  INV_X1 U5695 ( .A(n6982), .ZN(n4904) );
  NAND2_X1 U5696 ( .A1(n6861), .A2(n4781), .ZN(n4776) );
  NAND2_X1 U5697 ( .A1(n4778), .A2(n6861), .ZN(n4775) );
  INV_X1 U5698 ( .A(n4914), .ZN(n7401) );
  INV_X1 U5699 ( .A(n4916), .ZN(n7186) );
  AND3_X1 U5700 ( .A1(n4782), .A2(n7392), .A3(n4783), .ZN(n7426) );
  XNOR2_X1 U5701 ( .A(n4567), .B(n4566), .ZN(n7403) );
  INV_X1 U5702 ( .A(n7427), .ZN(n4566) );
  NAND2_X1 U5703 ( .A1(n7398), .A2(n7399), .ZN(n7420) );
  NAND2_X1 U5704 ( .A1(n4914), .A2(n4913), .ZN(n4567) );
  NAND2_X1 U5705 ( .A1(n7402), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4913) );
  OR2_X1 U5706 ( .A1(n7434), .A2(n7433), .ZN(n7542) );
  XNOR2_X1 U5707 ( .A(n7579), .B(n7571), .ZN(n7543) );
  NOR2_X1 U5708 ( .A1(n7543), .A2(n6198), .ZN(n7582) );
  OR2_X1 U5709 ( .A1(n8357), .A2(n8356), .ZN(n8395) );
  NOR2_X1 U5710 ( .A1(n7587), .A2(n6220), .ZN(n4570) );
  NOR2_X1 U5711 ( .A1(n8389), .A2(n8388), .ZN(n8390) );
  OR2_X1 U5712 ( .A1(n8454), .A2(n8455), .ZN(n4792) );
  INV_X1 U5713 ( .A(n4562), .ZN(n8452) );
  XNOR2_X1 U5714 ( .A(n8501), .B(n8502), .ZN(n8476) );
  NAND2_X1 U5715 ( .A1(n4790), .A2(n4789), .ZN(n4561) );
  NAND2_X1 U5716 ( .A1(n8475), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4789) );
  INV_X1 U5717 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8531) );
  NAND2_X1 U5718 ( .A1(n6384), .A2(n6383), .ZN(n6394) );
  INV_X1 U5719 ( .A(n6385), .ZN(n6384) );
  NAND2_X1 U5720 ( .A1(n6351), .A2(n6350), .ZN(n6363) );
  OR2_X1 U5721 ( .A1(n6317), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6327) );
  NAND2_X1 U5722 ( .A1(n6304), .A2(n10285), .ZN(n6317) );
  INV_X1 U5723 ( .A(n6305), .ZN(n6304) );
  NAND2_X1 U5724 ( .A1(n6279), .A2(n6278), .ZN(n6290) );
  INV_X1 U5725 ( .A(n6280), .ZN(n6279) );
  NAND2_X1 U5726 ( .A1(n6255), .A2(n6254), .ZN(n6266) );
  INV_X1 U5727 ( .A(n6264), .ZN(n6255) );
  INV_X1 U5728 ( .A(n8714), .ZN(n8743) );
  NAND2_X1 U5729 ( .A1(n6217), .A2(n6216), .ZN(n6230) );
  INV_X1 U5730 ( .A(n6218), .ZN(n6217) );
  NAND2_X1 U5731 ( .A1(n6205), .A2(n4751), .ZN(n7780) );
  NAND2_X1 U5732 ( .A1(n5030), .A2(n5029), .ZN(n7781) );
  OR2_X1 U5733 ( .A1(n5028), .A2(n6440), .ZN(n5022) );
  OR2_X1 U5734 ( .A1(n7292), .A2(n7688), .ZN(n8147) );
  AND2_X1 U5735 ( .A1(n8160), .A2(n8153), .ZN(n8311) );
  OR2_X1 U5736 ( .A1(n6128), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U5737 ( .A1(n5008), .A2(n6430), .ZN(n7248) );
  NAND2_X1 U5738 ( .A1(n7999), .A2(n6103), .ZN(n6117) );
  INV_X1 U5739 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U5740 ( .A1(n6116), .A2(n6115), .ZN(n6128) );
  INV_X1 U5741 ( .A(n6117), .ZN(n6116) );
  INV_X1 U5742 ( .A(n8197), .ZN(n4747) );
  NAND2_X1 U5743 ( .A1(n6954), .A2(n6955), .ZN(n4998) );
  NAND2_X1 U5744 ( .A1(n6425), .A2(n8192), .ZN(n6908) );
  NAND2_X1 U5745 ( .A1(n6757), .A2(n6625), .ZN(n6928) );
  AND2_X1 U5746 ( .A1(n6480), .A2(n6481), .ZN(n4727) );
  NAND2_X1 U5747 ( .A1(n6404), .A2(n6403), .ZN(n6520) );
  XNOR2_X1 U5748 ( .A(n8558), .B(n8564), .ZN(n8552) );
  NAND2_X1 U5749 ( .A1(n4864), .A2(n8272), .ZN(n8563) );
  INV_X1 U5750 ( .A(n8565), .ZN(n8584) );
  AND3_X1 U5751 ( .A1(n6331), .A2(n6330), .A3(n6329), .ZN(n8649) );
  NAND2_X1 U5752 ( .A1(n6303), .A2(n6302), .ZN(n8788) );
  OAI21_X1 U5753 ( .B1(n8712), .B2(n5036), .A(n5031), .ZN(n8677) );
  INV_X1 U5754 ( .A(n5033), .ZN(n5031) );
  NAND2_X1 U5755 ( .A1(n6277), .A2(n6276), .ZN(n8795) );
  AND2_X1 U5756 ( .A1(n8226), .A2(n8228), .ZN(n8736) );
  INV_X1 U5757 ( .A(n10039), .ZN(n10061) );
  INV_X1 U5758 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6046) );
  INV_X1 U5759 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6484) );
  AND2_X1 U5760 ( .A1(n6419), .A2(n6418), .ZN(n8280) );
  OR2_X1 U5761 ( .A1(n6123), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n6134) );
  INV_X1 U5762 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6135) );
  NOR2_X1 U5763 ( .A1(n9027), .A2(n9028), .ZN(n5973) );
  NAND2_X1 U5764 ( .A1(n8998), .A2(n4984), .ZN(n4981) );
  AND2_X1 U5765 ( .A1(n6690), .A2(n5776), .ZN(n6541) );
  INV_X1 U5766 ( .A(n5861), .ZN(n4975) );
  NAND2_X1 U5767 ( .A1(n5861), .A2(n4497), .ZN(n4974) );
  INV_X1 U5768 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5278) );
  OR2_X1 U5769 ( .A1(n5279), .A2(n5278), .ZN(n5299) );
  NAND2_X1 U5770 ( .A1(n5775), .A2(n4496), .ZN(n6692) );
  NAND2_X1 U5771 ( .A1(n4642), .A2(n4641), .ZN(n5766) );
  NAND2_X1 U5772 ( .A1(n4643), .A2(n9848), .ZN(n4642) );
  OR2_X1 U5773 ( .A1(n5449), .A2(n5448), .ZN(n5469) );
  OAI21_X1 U5774 ( .B1(n9218), .B2(n9719), .A(n4505), .ZN(n9223) );
  NAND2_X1 U5775 ( .A1(n4437), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5119) );
  AOI21_X1 U5776 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7237), .A(n7236), .ZN(
        n7240) );
  NOR2_X1 U5777 ( .A1(n7366), .A2(n7365), .ZN(n7369) );
  OR2_X1 U5778 ( .A1(n9394), .A2(n9393), .ZN(n9407) );
  NAND2_X1 U5779 ( .A1(n4571), .A2(n4478), .ZN(n4834) );
  AND2_X1 U5780 ( .A1(n9407), .A2(n9406), .ZN(n9410) );
  INV_X1 U5781 ( .A(n4968), .ZN(n4967) );
  OAI21_X1 U5782 ( .B1(n5679), .B2(n5198), .A(n5680), .ZN(n4968) );
  AND2_X1 U5783 ( .A1(n5660), .A2(n5659), .ZN(n7953) );
  NAND2_X1 U5784 ( .A1(n9520), .A2(n4844), .ZN(n9462) );
  AND2_X1 U5785 ( .A1(n9283), .A2(n9213), .ZN(n9496) );
  AND2_X1 U5786 ( .A1(n9060), .A2(n9196), .ZN(n9550) );
  AOI21_X1 U5787 ( .B1(n4951), .B2(n4950), .A(n4518), .ZN(n4949) );
  NOR2_X1 U5788 ( .A1(n7718), .A2(n9956), .ZN(n7737) );
  NAND2_X1 U5789 ( .A1(n4948), .A2(n4951), .ZN(n7716) );
  NAND2_X1 U5790 ( .A1(n7499), .A2(n5352), .ZN(n4948) );
  AND4_X1 U5791 ( .A1(n5304), .A2(n5303), .A3(n5302), .A4(n5301), .ZN(n9792)
         );
  OAI21_X1 U5792 ( .B1(n7323), .B2(n9247), .A(n9255), .ZN(n7337) );
  INV_X1 U5793 ( .A(n9086), .ZN(n7343) );
  INV_X1 U5794 ( .A(n7311), .ZN(n4837) );
  NAND2_X1 U5795 ( .A1(n9239), .A2(n5058), .ZN(n9834) );
  AND2_X1 U5796 ( .A1(n6584), .A2(n4461), .ZN(n4757) );
  NAND2_X1 U5797 ( .A1(n6801), .A2(n9080), .ZN(n4574) );
  NOR2_X1 U5798 ( .A1(n6549), .A2(n6558), .ZN(n4850) );
  NAND2_X1 U5799 ( .A1(n5617), .A2(n5616), .ZN(n9522) );
  AND2_X1 U5800 ( .A1(n5588), .A2(n5587), .ZN(n9648) );
  AND2_X1 U5801 ( .A1(n5626), .A2(n5625), .ZN(n9649) );
  NAND2_X1 U5802 ( .A1(n9217), .A2(n9298), .ZN(n9960) );
  INV_X1 U5803 ( .A(n9949), .ZN(n9894) );
  INV_X1 U5804 ( .A(n9304), .ZN(n6004) );
  OAI21_X1 U5805 ( .B1(n8121), .B2(n8120), .A(n8119), .ZN(n8129) );
  OR2_X1 U5806 ( .A1(n8118), .A2(n8117), .ZN(n8119) );
  NAND2_X1 U5807 ( .A1(n4955), .A2(n5095), .ZN(n4954) );
  INV_X1 U5808 ( .A(n4956), .ZN(n4955) );
  XNOR2_X1 U5809 ( .A(n8129), .B(n8128), .ZN(n9054) );
  XNOR2_X1 U5810 ( .A(n5732), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5754) );
  OAI211_X1 U5811 ( .C1(n4558), .C2(n4701), .A(n4692), .B(n4695), .ZN(n6696)
         );
  NAND2_X1 U5812 ( .A1(n4558), .A2(n4698), .ZN(n4692) );
  OR2_X1 U5813 ( .A1(n5238), .A2(n4660), .ZN(n4653) );
  NAND2_X1 U5814 ( .A1(n5072), .A2(n5071), .ZN(n5187) );
  NOR2_X1 U5815 ( .A1(n7975), .A2(n7977), .ZN(n7976) );
  XNOR2_X1 U5816 ( .A(n7752), .B(n8345), .ZN(n7598) );
  INV_X1 U5817 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U5818 ( .A1(n8063), .A2(n4807), .ZN(n4800) );
  AOI21_X1 U5819 ( .B1(n4824), .B2(n7977), .A(n4508), .ZN(n4822) );
  AND4_X1 U5820 ( .A1(n6313), .A2(n6312), .A3(n6311), .A4(n6310), .ZN(n8648)
         );
  AOI21_X1 U5821 ( .B1(n8063), .B2(n8062), .A(n8061), .ZN(n8065) );
  OR2_X1 U5822 ( .A1(n7976), .A2(n4825), .ZN(n8105) );
  NOR2_X1 U5823 ( .A1(n7976), .A2(n4827), .ZN(n8107) );
  OR2_X1 U5824 ( .A1(n7017), .A2(n7646), .ZN(n8113) );
  NAND4_X1 U5825 ( .A1(n6177), .A2(n6176), .A3(n6175), .A4(n6174), .ZN(n8346)
         );
  OR2_X1 U5826 ( .A1(n4441), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6093) );
  OR2_X1 U5827 ( .A1(n4439), .A2(n7115), .ZN(n6082) );
  OR2_X1 U5828 ( .A1(n6051), .A2(n6064), .ZN(n6053) );
  NAND2_X1 U5829 ( .A1(n6077), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6052) );
  NOR2_X1 U5830 ( .A1(n6780), .A2(n4498), .ZN(n6784) );
  AOI21_X1 U5831 ( .B1(n6793), .B2(n6791), .A(n6792), .ZN(n6848) );
  AOI21_X1 U5832 ( .B1(n7083), .B2(n7074), .A(n7073), .ZN(n7173) );
  NAND2_X1 U5833 ( .A1(n4782), .A2(n4783), .ZN(n7393) );
  NOR2_X1 U5834 ( .A1(n6168), .A2(n7394), .ZN(n7428) );
  NAND2_X1 U5835 ( .A1(n7571), .A2(n4912), .ZN(n4911) );
  AOI21_X1 U5836 ( .B1(n4465), .B2(n7416), .A(n4534), .ZN(n4910) );
  XNOR2_X1 U5837 ( .A(n8395), .B(n8374), .ZN(n8358) );
  NOR2_X1 U5838 ( .A1(n8358), .A2(n8364), .ZN(n8398) );
  XNOR2_X1 U5839 ( .A(n4561), .B(n8471), .ZN(n8466) );
  NAND2_X1 U5840 ( .A1(n5000), .A2(n6481), .ZN(n7957) );
  OAI21_X1 U5841 ( .B1(n8581), .B2(n4452), .A(n6466), .ZN(n8572) );
  NAND2_X1 U5842 ( .A1(n6360), .A2(n6359), .ZN(n8585) );
  NAND2_X1 U5843 ( .A1(n4724), .A2(n8265), .ZN(n8588) );
  OR2_X1 U5844 ( .A1(n8598), .A2(n8298), .ZN(n4724) );
  NAND2_X1 U5845 ( .A1(n5002), .A2(n5004), .ZN(n8592) );
  OR2_X1 U5846 ( .A1(n6457), .A2(n5005), .ZN(n5002) );
  NAND2_X1 U5847 ( .A1(n8671), .A2(n8249), .ZN(n8665) );
  INV_X1 U5848 ( .A(n5037), .ZN(n8686) );
  AOI21_X1 U5849 ( .B1(n8712), .B2(n5043), .A(n5041), .ZN(n5037) );
  NAND2_X1 U5850 ( .A1(n6215), .A2(n6214), .ZN(n10060) );
  OAI211_X1 U5851 ( .C1(n4558), .C2(n4694), .A(n4693), .B(n6183), .ZN(n6215)
         );
  NAND2_X1 U5852 ( .A1(n4695), .A2(n4701), .ZN(n4694) );
  INV_X1 U5853 ( .A(n5030), .ZN(n7706) );
  NAND2_X1 U5854 ( .A1(n6187), .A2(n6186), .ZN(n10049) );
  INV_X1 U5855 ( .A(n8720), .ZN(n8708) );
  NAND2_X1 U5856 ( .A1(n7104), .A2(n8197), .ZN(n6962) );
  INV_X1 U5857 ( .A(n8785), .ZN(n8808) );
  INV_X1 U5858 ( .A(n6520), .ZN(n7959) );
  XOR2_X1 U5859 ( .A(n8552), .B(n8550), .Z(n8820) );
  NAND2_X1 U5860 ( .A1(n6382), .A2(n6381), .ZN(n8826) );
  NAND2_X1 U5861 ( .A1(n6373), .A2(n6372), .ZN(n8832) );
  NAND2_X1 U5862 ( .A1(n4719), .A2(n4720), .ZN(n8577) );
  OR2_X1 U5863 ( .A1(n8598), .A2(n4723), .ZN(n4719) );
  NAND2_X1 U5864 ( .A1(n8617), .A2(n6461), .ZN(n8604) );
  NAND2_X1 U5865 ( .A1(n7451), .A2(n6183), .ZN(n4887) );
  NAND2_X1 U5866 ( .A1(n6324), .A2(n6323), .ZN(n8859) );
  NAND2_X1 U5867 ( .A1(n8641), .A2(n8246), .ZN(n8626) );
  NAND2_X1 U5868 ( .A1(n6289), .A2(n6288), .ZN(n8872) );
  NAND2_X1 U5869 ( .A1(n6253), .A2(n6252), .ZN(n8879) );
  AOI21_X1 U5870 ( .B1(n8712), .B2(n6448), .A(n5046), .ZN(n8702) );
  NAND2_X1 U5871 ( .A1(n6240), .A2(n6239), .ZN(n8887) );
  INV_X1 U5872 ( .A(n8864), .ZN(n8888) );
  INV_X1 U5873 ( .A(n8882), .ZN(n8889) );
  NAND2_X1 U5874 ( .A1(n6074), .A2(n4455), .ZN(n4742) );
  OR2_X1 U5875 ( .A1(n10062), .A2(n10039), .ZN(n8864) );
  AND2_X1 U5876 ( .A1(n6644), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6625) );
  INV_X1 U5877 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8894) );
  INV_X1 U5878 ( .A(n8280), .ZN(n8144) );
  INV_X1 U5879 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6299) );
  INV_X1 U5880 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6751) );
  INV_X1 U5881 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6689) );
  INV_X1 U5882 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10249) );
  INV_X1 U5883 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6573) );
  INV_X1 U5884 ( .A(n7079), .ZN(n7180) );
  INV_X1 U5885 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6565) );
  INV_X1 U5886 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6562) );
  NAND2_X1 U5887 ( .A1(n6209), .A2(n4773), .ZN(n4772) );
  NAND2_X1 U5888 ( .A1(n4625), .A2(n5885), .ZN(n8905) );
  INV_X1 U5889 ( .A(n4627), .ZN(n4625) );
  NAND2_X1 U5890 ( .A1(n4961), .A2(n5787), .ZN(n6938) );
  NAND2_X1 U5891 ( .A1(n6833), .A2(n6834), .ZN(n4961) );
  NOR2_X1 U5892 ( .A1(n9026), .A2(n4993), .ZN(n7951) );
  NAND2_X1 U5893 ( .A1(n8998), .A2(n5935), .ZN(n8939) );
  INV_X1 U5894 ( .A(n4647), .ZN(n8962) );
  NAND2_X1 U5895 ( .A1(n8970), .A2(n5907), .ZN(n8980) );
  AND2_X1 U5896 ( .A1(n5607), .A2(n5606), .ZN(n8994) );
  NAND2_X1 U5897 ( .A1(n4521), .A2(n4453), .ZN(n4978) );
  INV_X1 U5898 ( .A(n4648), .ZN(n8988) );
  INV_X1 U5899 ( .A(n6990), .ZN(n5799) );
  NAND2_X1 U5900 ( .A1(n7619), .A2(n4529), .ZN(n7692) );
  AND2_X1 U5901 ( .A1(n5524), .A2(n5523), .ZN(n9681) );
  INV_X1 U5902 ( .A(n8983), .ZN(n9045) );
  AOI21_X1 U5903 ( .B1(n5907), .B2(n4620), .A(n4492), .ZN(n4619) );
  INV_X1 U5904 ( .A(n5907), .ZN(n4621) );
  INV_X1 U5905 ( .A(n8972), .ZN(n4620) );
  INV_X1 U5906 ( .A(n4963), .ZN(n4962) );
  NAND2_X1 U5907 ( .A1(n5895), .A2(n5891), .ZN(n9041) );
  INV_X1 U5908 ( .A(n9039), .ZN(n9050) );
  NAND2_X1 U5909 ( .A1(n9299), .A2(n9298), .ZN(n9300) );
  NAND2_X1 U5910 ( .A1(n5641), .A2(n5640), .ZN(n9515) );
  INV_X1 U5911 ( .A(n8994), .ZN(n9530) );
  INV_X1 U5912 ( .A(n9648), .ZN(n9556) );
  CLKBUF_X1 U5913 ( .A(n5768), .Z(n9325) );
  AOI21_X1 U5914 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n9332), .A(n9326), .ZN(
        n6825) );
  NAND2_X1 U5915 ( .A1(n9371), .A2(n9370), .ZN(n9369) );
  NAND2_X1 U5916 ( .A1(n9356), .A2(n4553), .ZN(n9371) );
  NAND2_X1 U5917 ( .A1(n4554), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4553) );
  INV_X1 U5918 ( .A(n9353), .ZN(n4554) );
  AOI21_X1 U5919 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6629), .A(n6628), .ZN(
        n6631) );
  AOI21_X1 U5920 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6703), .A(n6699), .ZN(
        n6700) );
  OR2_X1 U5921 ( .A1(n6604), .A2(n6815), .ZN(n9445) );
  OR2_X1 U5922 ( .A1(n9438), .A2(n9437), .ZN(n9439) );
  AOI21_X1 U5923 ( .B1(n4931), .B2(n4933), .A(n4509), .ZN(n4930) );
  NAND2_X1 U5924 ( .A1(n9507), .A2(n5642), .ZN(n9487) );
  NAND2_X1 U5925 ( .A1(n4936), .A2(n4940), .ZN(n7871) );
  NAND2_X1 U5926 ( .A1(n9543), .A2(n4943), .ZN(n4936) );
  INV_X1 U5927 ( .A(n9649), .ZN(n9498) );
  NAND2_X1 U5928 ( .A1(n4944), .A2(n4946), .ZN(n9533) );
  NAND2_X1 U5929 ( .A1(n4945), .A2(n4473), .ZN(n4944) );
  NAND2_X1 U5930 ( .A1(n5578), .A2(n5577), .ZN(n9540) );
  NAND2_X1 U5931 ( .A1(n4926), .A2(n5526), .ZN(n9562) );
  NAND2_X1 U5932 ( .A1(n7885), .A2(n5708), .ZN(n7886) );
  NAND2_X1 U5933 ( .A1(n5485), .A2(n5484), .ZN(n9588) );
  AND4_X1 U5934 ( .A1(n5455), .A2(n5454), .A3(n5453), .A4(n5452), .ZN(n9603)
         );
  NAND2_X1 U5935 ( .A1(n5705), .A2(n9273), .ZN(n9621) );
  NAND2_X1 U5936 ( .A1(n9786), .A2(n5439), .ZN(n9613) );
  OR2_X1 U5937 ( .A1(n7804), .A2(n9094), .ZN(n9786) );
  NAND2_X1 U5938 ( .A1(n5429), .A2(n5428), .ZN(n7813) );
  AND4_X1 U5939 ( .A1(n5413), .A2(n5412), .A3(n5411), .A4(n5410), .ZN(n9951)
         );
  AND2_X1 U5940 ( .A1(n7662), .A2(n9257), .ZN(n7724) );
  NAND2_X1 U5941 ( .A1(n7500), .A2(n9163), .ZN(n7664) );
  AND4_X1 U5942 ( .A1(n5328), .A2(n5327), .A3(n5326), .A4(n5325), .ZN(n9926)
         );
  NAND2_X1 U5943 ( .A1(n5699), .A2(n5058), .ZN(n4616) );
  INV_X1 U5944 ( .A(n9822), .ZN(n9837) );
  OR3_X1 U5945 ( .A1(n7130), .A2(n7129), .A3(n7128), .ZN(n7131) );
  INV_X1 U5946 ( .A(n9606), .ZN(n9851) );
  NAND2_X1 U5947 ( .A1(n5600), .A2(n5599), .ZN(n9731) );
  NAND2_X1 U5948 ( .A1(n5540), .A2(n5539), .ZN(n9740) );
  INV_X1 U5949 ( .A(n5092), .ZN(n7868) );
  XNOR2_X1 U5950 ( .A(n5663), .B(n5662), .ZN(n7849) );
  NAND2_X1 U5951 ( .A1(n5726), .A2(n5727), .ZN(n7802) );
  MUX2_X1 U5952 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5725), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n5727) );
  OR2_X1 U5953 ( .A1(n5729), .A2(n5080), .ZN(n5730) );
  INV_X1 U5954 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5683) );
  OAI21_X1 U5955 ( .B1(n5689), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5684) );
  NOR2_X1 U5956 ( .A1(n5339), .A2(n5377), .ZN(n7275) );
  AND2_X1 U5957 ( .A1(n5316), .A2(n5295), .ZN(n7029) );
  INV_X1 U5958 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U5959 ( .A1(n5106), .A2(n5105), .ZN(n6607) );
  NAND2_X1 U5960 ( .A1(n7200), .A2(n7199), .ZN(n7203) );
  NAND2_X1 U5961 ( .A1(n4812), .A2(n8104), .ZN(n4811) );
  INV_X1 U5962 ( .A(n4918), .ZN(n8385) );
  INV_X1 U5963 ( .A(n4565), .ZN(n8439) );
  INV_X1 U5964 ( .A(n4908), .ZN(n8442) );
  AND2_X1 U5965 ( .A1(n4921), .A2(n4919), .ZN(n8510) );
  OAI21_X1 U5966 ( .B1(n8518), .B2(n4458), .A(n10419), .ZN(n4921) );
  NAND2_X1 U5967 ( .A1(n4989), .A2(n4990), .ZN(n4986) );
  OAI21_X1 U5968 ( .B1(n9721), .B2(n9981), .A(n4766), .ZN(P1_U3550) );
  AOI21_X1 U5969 ( .B1(n9488), .B2(n9673), .A(n4767), .ZN(n4766) );
  NOR2_X1 U5970 ( .A1(n9983), .A2(n10143), .ZN(n4767) );
  NAND2_X1 U5971 ( .A1(n4923), .A2(n4922), .ZN(P1_U3519) );
  NOR2_X1 U5972 ( .A1(n5756), .A2(n4537), .ZN(n4922) );
  NAND2_X1 U5973 ( .A1(n5757), .A2(n9967), .ZN(n4923) );
  OAI21_X1 U5974 ( .B1(n9721), .B2(n9965), .A(n4556), .ZN(P1_U3518) );
  INV_X1 U5975 ( .A(n4557), .ZN(n4556) );
  OAI22_X1 U5976 ( .A1(n9723), .A2(n9754), .B1(n9967), .B2(n9722), .ZN(n4557)
         );
  XNOR2_X1 U5977 ( .A(n5481), .B(P1_IR_REG_19__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U5978 ( .A1(n4564), .A2(n4563), .ZN(n6792) );
  NAND2_X2 U5979 ( .A1(n6584), .A2(n4436), .ZN(n5247) );
  AND2_X1 U5980 ( .A1(n4974), .A2(n8948), .ZN(n4447) );
  NOR2_X1 U5981 ( .A1(n7417), .A2(n7416), .ZN(n4449) );
  NAND4_X1 U5982 ( .A1(n6235), .A2(n6234), .A3(n6233), .A4(n6232), .ZN(n8727)
         );
  NAND2_X1 U5983 ( .A1(n5829), .A2(n5828), .ZN(n4450) );
  OR2_X1 U5984 ( .A1(n6462), .A2(n8618), .ZN(n4451) );
  NOR2_X1 U5985 ( .A1(n8837), .A2(n8594), .ZN(n4452) );
  INV_X1 U5986 ( .A(n8265), .ZN(n4722) );
  INV_X1 U5987 ( .A(n6440), .ZN(n5029) );
  NOR2_X1 U5988 ( .A1(n5955), .A2(n5954), .ZN(n4453) );
  AND2_X1 U5989 ( .A1(n5973), .A2(n5962), .ZN(n4454) );
  XNOR2_X1 U5990 ( .A(n5684), .B(n5683), .ZN(n5691) );
  OAI211_X1 U5991 ( .C1(n4445), .C2(n10129), .A(n6337), .B(n6336), .ZN(n8633)
         );
  AND2_X1 U5992 ( .A1(n4436), .A2(n5100), .ZN(n4455) );
  AND2_X1 U5993 ( .A1(n4814), .A2(n4483), .ZN(n4456) );
  INV_X1 U5994 ( .A(n8756), .ZN(n4676) );
  NAND2_X1 U5995 ( .A1(n9151), .A2(n9780), .ZN(n4457) );
  AND2_X1 U5996 ( .A1(n8507), .A2(n8506), .ZN(n4458) );
  NOR2_X1 U5997 ( .A1(n9709), .A2(n9781), .ZN(n4459) );
  NAND2_X1 U5998 ( .A1(n7949), .A2(n5973), .ZN(n4460) );
  AND2_X1 U5999 ( .A1(n6549), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4461) );
  AND2_X1 U6000 ( .A1(n6549), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4462) );
  INV_X1 U6001 ( .A(n6482), .ZN(n5052) );
  AND2_X1 U6002 ( .A1(n7560), .A2(n7558), .ZN(n4463) );
  AND2_X1 U6003 ( .A1(n5810), .A2(n5805), .ZN(n4464) );
  AND2_X1 U6004 ( .A1(n7581), .A2(n7530), .ZN(n4465) );
  NAND2_X1 U6005 ( .A1(n4821), .A2(n7558), .ZN(n7559) );
  INV_X1 U6006 ( .A(n9488), .ZN(n9723) );
  AND2_X1 U6007 ( .A1(n9459), .A2(n9310), .ZN(n4466) );
  NAND2_X1 U6008 ( .A1(n7995), .A2(n7011), .ZN(n7012) );
  NAND2_X1 U6009 ( .A1(n4969), .A2(n6539), .ZN(n5795) );
  OR2_X1 U6010 ( .A1(n7385), .A2(n9919), .ZN(n4467) );
  AND2_X1 U6011 ( .A1(n4677), .A2(n4673), .ZN(n4468) );
  OR3_X1 U6012 ( .A1(n7718), .A2(n9709), .A3(n4853), .ZN(n4469) );
  NAND2_X1 U6013 ( .A1(n6340), .A2(n6339), .ZN(n6462) );
  AND2_X1 U6014 ( .A1(n4800), .A2(n4804), .ZN(n4470) );
  AND2_X1 U6015 ( .A1(n9484), .A2(n9483), .ZN(n4471) );
  OR2_X1 U6016 ( .A1(n9731), .A2(n9530), .ZN(n4472) );
  INV_X2 U6017 ( .A(n5126), .ZN(n6549) );
  OR2_X1 U6018 ( .A1(n9665), .A2(n9311), .ZN(n4473) );
  AND2_X1 U6019 ( .A1(n8265), .A2(n8274), .ZN(n4474) );
  INV_X1 U6020 ( .A(n4701), .ZN(n4700) );
  NAND2_X1 U6021 ( .A1(n4705), .A2(n4704), .ZN(n4701) );
  AND2_X1 U6022 ( .A1(n8268), .A2(n4725), .ZN(n4475) );
  OAI22_X1 U6023 ( .A1(n8703), .A2(n5042), .B1(n6450), .B2(n8111), .ZN(n5041)
         );
  AND2_X1 U6024 ( .A1(n7693), .A2(n4634), .ZN(n4476) );
  NAND2_X1 U6025 ( .A1(n6074), .A2(n6549), .ZN(n6109) );
  OR2_X1 U6026 ( .A1(n8453), .A2(n8438), .ZN(n4477) );
  AND4_X1 U6027 ( .A1(n5293), .A2(n5073), .A3(n5074), .A4(n5188), .ZN(n4478)
         );
  AND2_X1 U6028 ( .A1(n5090), .A2(n5089), .ZN(n4479) );
  OR2_X1 U6029 ( .A1(n8226), .A2(n8292), .ZN(n4480) );
  INV_X1 U6030 ( .A(n8245), .ZN(n4736) );
  NAND2_X1 U6031 ( .A1(n4743), .A2(n4742), .ZN(n6882) );
  NAND2_X1 U6032 ( .A1(n5942), .A2(n5941), .ZN(n4481) );
  OR2_X1 U6033 ( .A1(n9198), .A2(n9219), .ZN(n4482) );
  NAND4_X1 U6034 ( .A1(n6082), .A2(n6081), .A3(n6080), .A4(n6079), .ZN(n8352)
         );
  INV_X1 U6035 ( .A(n8352), .ZN(n6088) );
  XNOR2_X1 U6036 ( .A(n5308), .B(SI_10_), .ZN(n5306) );
  OR2_X1 U6037 ( .A1(n7944), .A2(n4813), .ZN(n4483) );
  INV_X1 U6038 ( .A(n5058), .ZN(n4614) );
  OR2_X1 U6039 ( .A1(n5728), .A2(n5081), .ZN(n4484) );
  AND4_X1 U6040 ( .A1(n6030), .A2(n6029), .A3(n6096), .A4(n6135), .ZN(n4485)
         );
  NOR2_X1 U6041 ( .A1(n6584), .A2(n6822), .ZN(n4486) );
  NAND2_X1 U6042 ( .A1(n8258), .A2(n8262), .ZN(n8611) );
  NAND2_X1 U6043 ( .A1(n7942), .A2(n8341), .ZN(n4487) );
  INV_X1 U6044 ( .A(n8151), .ZN(n5027) );
  INV_X1 U6045 ( .A(n5353), .ZN(n4704) );
  XNOR2_X1 U6046 ( .A(n5354), .B(SI_12_), .ZN(n5353) );
  AND3_X1 U6047 ( .A1(n4867), .A2(n4860), .A3(n4859), .ZN(n4488) );
  AND2_X1 U6048 ( .A1(n8832), .A2(n8584), .ZN(n4489) );
  OR2_X1 U6049 ( .A1(n9802), .A2(n9317), .ZN(n4490) );
  AND2_X1 U6050 ( .A1(n5017), .A2(n5019), .ZN(n4491) );
  AND2_X1 U6051 ( .A1(n5910), .A2(n5909), .ZN(n4492) );
  NAND2_X1 U6052 ( .A1(n6227), .A2(n6226), .ZN(n8317) );
  AND2_X1 U6053 ( .A1(n9166), .A2(n9257), .ZN(n4493) );
  INV_X1 U6054 ( .A(n8259), .ZN(n4732) );
  OR2_X1 U6055 ( .A1(n8915), .A2(n5069), .ZN(n4494) );
  NOR2_X1 U6056 ( .A1(n4626), .A2(n4624), .ZN(n4495) );
  OR2_X1 U6057 ( .A1(n6539), .A2(n5771), .ZN(n4496) );
  INV_X1 U6058 ( .A(n4943), .ZN(n4942) );
  NOR2_X1 U6059 ( .A1(n5589), .A2(n4947), .ZN(n4943) );
  OR2_X1 U6060 ( .A1(n5862), .A2(n4976), .ZN(n4497) );
  AND2_X1 U6061 ( .A1(n6781), .A2(n6782), .ZN(n4498) );
  NAND2_X1 U6062 ( .A1(n9520), .A2(n4846), .ZN(n4848) );
  INV_X1 U6063 ( .A(n5806), .ZN(n9889) );
  AND3_X1 U6064 ( .A1(n5191), .A2(n5190), .A3(n5189), .ZN(n5806) );
  INV_X1 U6065 ( .A(n8152), .ZN(n6441) );
  AND2_X1 U6066 ( .A1(n8179), .A2(n8178), .ZN(n8152) );
  INV_X1 U6067 ( .A(n4805), .ZN(n4804) );
  NAND2_X1 U6068 ( .A1(n8013), .A2(n4806), .ZN(n4805) );
  AND2_X1 U6069 ( .A1(n7201), .A2(n7199), .ZN(n4499) );
  AND3_X1 U6070 ( .A1(n8261), .A2(n8322), .A3(n8260), .ZN(n4500) );
  AND2_X1 U6071 ( .A1(n5973), .A2(n8961), .ZN(n4501) );
  AND2_X1 U6072 ( .A1(n5765), .A2(n5761), .ZN(n4502) );
  OR2_X1 U6073 ( .A1(n4691), .A2(n8223), .ZN(n4503) );
  AND2_X1 U6074 ( .A1(n4468), .A2(n4671), .ZN(n4504) );
  INV_X1 U6075 ( .A(n6451), .ZN(n5045) );
  AND2_X1 U6076 ( .A1(n9295), .A2(n4555), .ZN(n4505) );
  AND2_X1 U6077 ( .A1(n8832), .A2(n8565), .ZN(n4506) );
  INV_X1 U6078 ( .A(n6792), .ZN(n4781) );
  INV_X1 U6079 ( .A(n9259), .ZN(n4606) );
  AND2_X1 U6080 ( .A1(n8558), .A2(n8564), .ZN(n4507) );
  INV_X1 U6081 ( .A(n5020), .ZN(n5019) );
  AND2_X1 U6082 ( .A1(n6470), .A2(n5021), .ZN(n5020) );
  NOR2_X1 U6083 ( .A1(n7910), .A2(n8302), .ZN(n4508) );
  NOR2_X1 U6084 ( .A1(n9488), .A2(n9497), .ZN(n4509) );
  NOR2_X1 U6085 ( .A1(n9540), .A2(n9556), .ZN(n4510) );
  INV_X1 U6086 ( .A(n4699), .ZN(n4698) );
  NAND2_X1 U6087 ( .A1(n4708), .A2(n5353), .ZN(n4699) );
  INV_X1 U6088 ( .A(n4947), .ZN(n4946) );
  NOR2_X1 U6089 ( .A1(n9549), .A2(n9659), .ZN(n4947) );
  OR2_X1 U6090 ( .A1(n4605), .A2(n4604), .ZN(n4511) );
  NAND2_X1 U6091 ( .A1(n8147), .A2(n8162), .ZN(n8315) );
  NAND2_X1 U6092 ( .A1(n5052), .A2(n5051), .ZN(n6058) );
  NAND3_X1 U6093 ( .A1(n6164), .A2(n5055), .A3(n4448), .ZN(n4512) );
  AND2_X1 U6094 ( .A1(n8060), .A2(n8583), .ZN(n4513) );
  OR2_X1 U6095 ( .A1(n6482), .A2(n6039), .ZN(n4514) );
  NAND3_X1 U6096 ( .A1(n6164), .A2(n4448), .A3(n5054), .ZN(n4515) );
  INV_X1 U6097 ( .A(n6468), .ZN(n5021) );
  OR2_X1 U6098 ( .A1(n8317), .A2(n8225), .ZN(n4516) );
  INV_X1 U6099 ( .A(n9174), .ZN(n9620) );
  AND2_X1 U6100 ( .A1(n9185), .A2(n9176), .ZN(n9174) );
  INV_X1 U6101 ( .A(n5025), .ZN(n5024) );
  NAND2_X1 U6102 ( .A1(n6441), .A2(n5026), .ZN(n5025) );
  AND2_X1 U6103 ( .A1(n4777), .A2(n6972), .ZN(n4517) );
  NAND2_X1 U6104 ( .A1(n5391), .A2(n7715), .ZN(n4518) );
  AND2_X1 U6105 ( .A1(n4942), .A2(n4472), .ZN(n4519) );
  OR2_X1 U6106 ( .A1(n6852), .A2(n6790), .ZN(n4564) );
  AND2_X1 U6107 ( .A1(n9155), .A2(n9217), .ZN(n4520) );
  NAND2_X1 U6108 ( .A1(n4887), .A2(n6333), .ZN(n6458) );
  AND2_X1 U6109 ( .A1(n9505), .A2(n9515), .ZN(n9211) );
  INV_X1 U6110 ( .A(n9211), .ZN(n9283) );
  INV_X1 U6111 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5083) );
  INV_X1 U6112 ( .A(n8267), .ZN(n4868) );
  INV_X1 U6113 ( .A(n5041), .ZN(n5040) );
  OR2_X1 U6114 ( .A1(n4494), .A2(n4980), .ZN(n4521) );
  NAND2_X1 U6115 ( .A1(n6463), .A2(n5006), .ZN(n4522) );
  AND2_X1 U6116 ( .A1(n5636), .A2(n5635), .ZN(n9505) );
  INV_X1 U6117 ( .A(n9505), .ZN(n4847) );
  AND2_X1 U6118 ( .A1(n9268), .A2(n9273), .ZN(n9094) );
  INV_X1 U6119 ( .A(n8246), .ZN(n4733) );
  OR2_X1 U6120 ( .A1(n8653), .A2(n8660), .ZN(n8246) );
  AND2_X1 U6121 ( .A1(n5053), .A2(n6040), .ZN(n4523) );
  AND2_X1 U6122 ( .A1(n4957), .A2(n5082), .ZN(n4524) );
  AND2_X1 U6123 ( .A1(n4695), .A2(n4699), .ZN(n4525) );
  NOR2_X1 U6124 ( .A1(n5419), .A2(n10232), .ZN(n4526) );
  AND2_X1 U6125 ( .A1(n4987), .A2(n4986), .ZN(n4527) );
  INV_X1 U6126 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4773) );
  AND2_X1 U6127 ( .A1(n7631), .A2(n8147), .ZN(n8156) );
  INV_X1 U6128 ( .A(n4952), .ZN(n4951) );
  NAND2_X1 U6129 ( .A1(n9091), .A2(n4953), .ZN(n4952) );
  OR2_X1 U6130 ( .A1(n6852), .A2(n7123), .ZN(n4528) );
  BUF_X1 U6131 ( .A(n5434), .Z(n5671) );
  NAND2_X1 U6132 ( .A1(n7791), .A2(n5878), .ZN(n4627) );
  INV_X1 U6133 ( .A(n7707), .ZN(n5028) );
  NAND2_X1 U6134 ( .A1(n7662), .A2(n4493), .ZN(n7723) );
  INV_X1 U6135 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U6136 ( .A1(n4714), .A2(n6182), .ZN(n7630) );
  NAND2_X1 U6137 ( .A1(n7621), .A2(n7620), .ZN(n7619) );
  NAND2_X1 U6138 ( .A1(n8971), .A2(n8972), .ZN(n8970) );
  INV_X1 U6139 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6140 ( .A1(n4928), .A2(n5305), .ZN(n9791) );
  NAND2_X1 U6141 ( .A1(n7780), .A2(n8179), .ZN(n8750) );
  INV_X1 U6142 ( .A(n8091), .ZN(n4820) );
  INV_X1 U6143 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6485) );
  INV_X1 U6144 ( .A(n8072), .ZN(n4802) );
  NAND2_X1 U6145 ( .A1(n4627), .A2(n5884), .ZN(n8904) );
  AND2_X1 U6146 ( .A1(n7691), .A2(n7693), .ZN(n4529) );
  INV_X1 U6147 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5376) );
  OR2_X1 U6148 ( .A1(n7718), .A2(n4853), .ZN(n4530) );
  NAND2_X1 U6149 ( .A1(n6347), .A2(n6346), .ZN(n8618) );
  INV_X1 U6150 ( .A(n8618), .ZN(n8595) );
  INV_X1 U6151 ( .A(n7530), .ZN(n4549) );
  AND2_X1 U6152 ( .A1(n7217), .A2(n7216), .ZN(n8543) );
  INV_X1 U6153 ( .A(n8543), .ZN(n4675) );
  INV_X1 U6154 ( .A(n8211), .ZN(n4746) );
  AND2_X1 U6155 ( .A1(n10060), .A2(n8343), .ZN(n4531) );
  AND2_X1 U6156 ( .A1(n4962), .A2(n5895), .ZN(n4532) );
  INV_X1 U6157 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5100) );
  AND2_X1 U6158 ( .A1(n9740), .A2(n9555), .ZN(n4533) );
  AND2_X1 U6159 ( .A1(n4549), .A2(n7571), .ZN(n4534) );
  NOR2_X1 U6160 ( .A1(n4834), .A2(n4835), .ZN(n5444) );
  AND2_X1 U6161 ( .A1(n5022), .A2(n5024), .ZN(n4535) );
  AND2_X1 U6162 ( .A1(n6205), .A2(n8177), .ZN(n4536) );
  NAND2_X1 U6163 ( .A1(n4832), .A2(n6624), .ZN(n6875) );
  INV_X1 U6164 ( .A(n9031), .ZN(n9052) );
  INV_X2 U6165 ( .A(n9965), .ZN(n9967) );
  INV_X1 U6166 ( .A(n8292), .ZN(n8274) );
  NAND2_X1 U6167 ( .A1(n8194), .A2(n8337), .ZN(n8292) );
  NAND2_X1 U6168 ( .A1(n7256), .A2(n5826), .ZN(n7348) );
  INV_X1 U6169 ( .A(n7789), .ZN(n4973) );
  NOR2_X1 U6170 ( .A1(n9967), .A2(n5755), .ZN(n4537) );
  NAND2_X1 U6171 ( .A1(n4837), .A2(n5806), .ZN(n7224) );
  INV_X1 U6172 ( .A(n7224), .ZN(n4836) );
  AND4_X1 U6173 ( .A1(n4572), .A2(n4571), .A3(n5078), .A4(n4478), .ZN(n5734)
         );
  NAND2_X1 U6174 ( .A1(n6482), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6507) );
  AND2_X1 U6175 ( .A1(n4788), .A2(n4787), .ZN(n4538) );
  INV_X1 U6176 ( .A(n8039), .ZN(n8104) );
  NOR2_X1 U6177 ( .A1(n9075), .A2(n9760), .ZN(n4539) );
  AND2_X1 U6178 ( .A1(n5691), .A2(n5685), .ZN(n9217) );
  INV_X1 U6179 ( .A(n9239), .ZN(n4765) );
  CLKBUF_X1 U6180 ( .A(n6424), .Z(n8354) );
  AND2_X1 U6181 ( .A1(n4616), .A2(n9239), .ZN(n4540) );
  XNOR2_X1 U6182 ( .A(n6300), .B(n6299), .ZN(n8519) );
  NAND2_X1 U6183 ( .A1(n6727), .A2(n6739), .ZN(n6785) );
  INV_X1 U6184 ( .A(n5091), .ZN(n9767) );
  INV_X1 U6185 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4652) );
  NAND2_X1 U6186 ( .A1(n6402), .A2(n6401), .ZN(n8136) );
  OAI21_X1 U6187 ( .B1(n8562), .B2(n8275), .A(n8272), .ZN(n8550) );
  NAND2_X1 U6188 ( .A1(n4468), .A2(n8519), .ZN(n4672) );
  AOI21_X1 U6189 ( .B1(n4541), .B2(n8519), .A(n4504), .ZN(n4665) );
  INV_X1 U6190 ( .A(n4468), .ZN(n4541) );
  OAI21_X2 U6191 ( .B1(n8690), .B2(n8689), .A(n8238), .ZN(n8673) );
  NOR2_X1 U6192 ( .A1(n4672), .A2(n8339), .ZN(n4670) );
  NAND2_X1 U6193 ( .A1(n4799), .A2(n4797), .ZN(n8074) );
  NAND2_X1 U6194 ( .A1(n7043), .A2(n7042), .ZN(n7059) );
  AOI21_X1 U6195 ( .B1(n7752), .B2(n4829), .A(n4828), .ZN(n7754) );
  NAND2_X4 U6196 ( .A1(n5717), .A2(n7843), .ZN(n6584) );
  INV_X1 U6197 ( .A(n4835), .ZN(n4572) );
  NAND2_X1 U6198 ( .A1(n9512), .A2(n9114), .ZN(n9495) );
  NAND2_X1 U6199 ( .A1(n9494), .A2(n9213), .ZN(n9480) );
  NAND2_X1 U6200 ( .A1(n9513), .A2(n9518), .ZN(n9512) );
  AND2_X2 U6201 ( .A1(n5697), .A2(n9240), .ZN(n7306) );
  NAND2_X1 U6202 ( .A1(n9592), .A2(n9594), .ZN(n9591) );
  NAND2_X1 U6203 ( .A1(n5703), .A2(n9159), .ZN(n7501) );
  NAND2_X1 U6204 ( .A1(n4653), .A2(n4657), .ZN(n5288) );
  INV_X1 U6205 ( .A(n9144), .ZN(n4547) );
  AOI21_X2 U6206 ( .B1(n4547), .B2(n9140), .A(n4546), .ZN(n9088) );
  NAND2_X1 U6207 ( .A1(n5126), .A2(n5101), .ZN(n5113) );
  INV_X1 U6208 ( .A(n9088), .ZN(n9247) );
  NAND4_X2 U6209 ( .A1(n5181), .A2(n5180), .A3(n5179), .A4(n5178), .ZN(n9321)
         );
  NAND2_X1 U6210 ( .A1(n4872), .A2(n4874), .ZN(n5508) );
  INV_X2 U6211 ( .A(n5346), .ZN(n6667) );
  OAI21_X1 U6212 ( .B1(n5417), .B2(n4526), .A(n5420), .ZN(n5442) );
  NAND2_X1 U6213 ( .A1(n4898), .A2(n5289), .ZN(n5307) );
  NAND2_X1 U6214 ( .A1(n5512), .A2(n5511), .ZN(n5531) );
  NAND2_X1 U6215 ( .A1(n4548), .A2(n6782), .ZN(n6728) );
  INV_X1 U6216 ( .A(n6727), .ZN(n4548) );
  NOR2_X1 U6217 ( .A1(n8372), .A2(n4570), .ZN(n8380) );
  NOR2_X1 U6218 ( .A1(n7568), .A2(n7567), .ZN(n7570) );
  NAND2_X1 U6219 ( .A1(n6982), .A2(n4550), .ZN(n6855) );
  NOR2_X1 U6220 ( .A1(n6173), .A2(n7403), .ZN(n7413) );
  NOR2_X1 U6221 ( .A1(n4449), .A2(n4549), .ZN(n7566) );
  NAND2_X1 U6222 ( .A1(n7183), .A2(n7182), .ZN(n4916) );
  NAND2_X1 U6223 ( .A1(n4902), .A2(n4903), .ZN(n4899) );
  AND2_X2 U6224 ( .A1(n4552), .A2(n4551), .ZN(n6734) );
  NAND2_X1 U6225 ( .A1(n10417), .A2(n10416), .ZN(n10415) );
  NOR2_X1 U6226 ( .A1(n8487), .A2(n8488), .ZN(n8490) );
  NOR2_X1 U6227 ( .A1(n7428), .A2(n7429), .ZN(n7434) );
  NOR2_X2 U6228 ( .A1(n7582), .A2(n7583), .ZN(n7585) );
  NOR2_X2 U6229 ( .A1(n6097), .A2(n6110), .ZN(n6782) );
  INV_X1 U6230 ( .A(n9827), .ZN(n5699) );
  NAND2_X1 U6231 ( .A1(n7307), .A2(n7306), .ZN(n5698) );
  AOI21_X1 U6232 ( .B1(n4762), .B2(n5708), .A(n9065), .ZN(n4761) );
  NOR2_X1 U6233 ( .A1(n4486), .A2(n4757), .ZN(n4756) );
  NAND2_X1 U6234 ( .A1(n7735), .A2(n9265), .ZN(n7803) );
  NOR2_X1 U6235 ( .A1(n9389), .A2(n9390), .ZN(n9394) );
  NAND2_X1 U6236 ( .A1(n5629), .A2(n5628), .ZN(n5646) );
  NAND2_X1 U6237 ( .A1(n4856), .A2(n5125), .ZN(n5143) );
  NAND2_X1 U6238 ( .A1(n5165), .A2(n5164), .ZN(n5183) );
  NAND2_X1 U6239 ( .A1(n4649), .A2(n5197), .ZN(n5214) );
  NAND4_X1 U6240 ( .A1(n4588), .A2(n9111), .A3(n4592), .A4(n9112), .ZN(n4587)
         );
  NAND2_X1 U6241 ( .A1(n7344), .A2(n7343), .ZN(n4928) );
  OR2_X1 U6242 ( .A1(n4429), .A2(n9865), .ZN(n5132) );
  NAND2_X1 U6243 ( .A1(n9638), .A2(n9949), .ZN(n4770) );
  OAI22_X2 U6244 ( .A1(n7892), .A2(n5506), .B1(n9583), .B2(n7895), .ZN(n7882)
         );
  NAND2_X1 U6245 ( .A1(n9495), .A2(n9496), .ZN(n9494) );
  INV_X1 U6246 ( .A(n7220), .ZN(n4759) );
  NAND2_X1 U6247 ( .A1(n5700), .A2(n9243), .ZN(n7220) );
  NAND2_X1 U6248 ( .A1(n9591), .A2(n9188), .ZN(n9577) );
  NAND2_X1 U6249 ( .A1(n5705), .A2(n4771), .ZN(n9624) );
  NAND2_X1 U6250 ( .A1(n4760), .A2(n4761), .ZN(n9572) );
  NAND2_X1 U6251 ( .A1(n5611), .A2(n5610), .ZN(n5629) );
  INV_X1 U6252 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6272) );
  INV_X2 U6253 ( .A(n5247), .ZN(n5443) );
  NAND2_X1 U6254 ( .A1(n5512), .A2(n4891), .ZN(n4890) );
  NAND2_X1 U6255 ( .A1(n4665), .A2(n7646), .ZN(n4664) );
  NAND2_X1 U6256 ( .A1(n4587), .A2(n9216), .ZN(n9218) );
  NAND2_X1 U6257 ( .A1(n4707), .A2(n4705), .ZN(n5357) );
  INV_X1 U6258 ( .A(n4591), .ZN(n4590) );
  NAND2_X1 U6259 ( .A1(n9202), .A2(n4590), .ZN(n4589) );
  NAND2_X1 U6260 ( .A1(n9544), .A2(n9549), .ZN(n9536) );
  NAND2_X1 U6261 ( .A1(n9604), .A2(n9751), .ZN(n9585) );
  NAND2_X1 U6262 ( .A1(n9821), .A2(n9911), .ZN(n7385) );
  INV_X1 U6263 ( .A(n9637), .ZN(n4769) );
  NOR2_X2 U6264 ( .A1(n7301), .A2(n9833), .ZN(n9836) );
  NOR2_X4 U6265 ( .A1(n9522), .A2(n9521), .ZN(n9520) );
  NAND2_X2 U6266 ( .A1(n8430), .A2(n8429), .ZN(n4562) );
  NAND2_X1 U6267 ( .A1(n6784), .A2(n6783), .ZN(n6842) );
  INV_X1 U6268 ( .A(n4446), .ZN(n6650) );
  NOR2_X1 U6269 ( .A1(n7531), .A2(n7711), .ZN(n7567) );
  XNOR2_X1 U6270 ( .A(n8380), .B(n8397), .ZN(n8375) );
  NAND2_X1 U6271 ( .A1(n5238), .A2(n5237), .ZN(n4663) );
  NAND2_X1 U6272 ( .A1(n4663), .A2(n5241), .ZN(n5265) );
  NAND2_X1 U6273 ( .A1(n6247), .A2(n8228), .ZN(n8697) );
  NAND2_X1 U6274 ( .A1(n7445), .A2(n8311), .ZN(n6155) );
  NAND3_X1 U6275 ( .A1(n4664), .A2(n4666), .A3(n8338), .ZN(P2_U3296) );
  NAND2_X1 U6276 ( .A1(n6083), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n4774) );
  MUX2_X1 U6277 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n7115), .S(n6737), .Z(n10417)
         );
  NAND2_X1 U6278 ( .A1(n5399), .A2(n5398), .ZN(n5417) );
  NAND2_X1 U6279 ( .A1(n5609), .A2(n5608), .ZN(n5611) );
  NAND2_X1 U6280 ( .A1(n4650), .A2(n5185), .ZN(n5195) );
  AOI21_X1 U6281 ( .B1(n4569), .B2(n9225), .A(n4568), .ZN(n9226) );
  AND2_X1 U6282 ( .A1(n9224), .A2(n9229), .ZN(n4568) );
  NAND2_X1 U6283 ( .A1(n9228), .A2(n5716), .ZN(n4569) );
  NAND2_X1 U6284 ( .A1(n4656), .A2(n4654), .ZN(n4898) );
  AND2_X2 U6285 ( .A1(n5072), .A2(n5071), .ZN(n4571) );
  NAND4_X1 U6286 ( .A1(n4752), .A2(n4754), .A3(n4755), .A4(n4753), .ZN(n4835)
         );
  NAND2_X1 U6287 ( .A1(n4574), .A2(n5695), .ZN(n7307) );
  XNOR2_X2 U6288 ( .A(n5762), .B(n9848), .ZN(n9080) );
  NOR2_X1 U6289 ( .A1(n5768), .A2(n7141), .ZN(n6801) );
  OAI211_X1 U6290 ( .C1(n4580), .C2(n9217), .A(n4576), .B(n9532), .ZN(n4575)
         );
  NAND2_X1 U6291 ( .A1(n4577), .A2(n9217), .ZN(n4576) );
  NAND2_X1 U6292 ( .A1(n4578), .A2(n9196), .ZN(n4577) );
  NAND2_X1 U6293 ( .A1(n4579), .A2(n9197), .ZN(n4578) );
  OAI21_X1 U6294 ( .B1(n9195), .B2(n9194), .A(n9571), .ZN(n4579) );
  OAI21_X1 U6295 ( .B1(n9182), .B2(n9181), .A(n9571), .ZN(n4581) );
  NAND2_X1 U6296 ( .A1(n9149), .A2(n4600), .ZN(n4596) );
  NAND2_X1 U6297 ( .A1(n4596), .A2(n4597), .ZN(n9150) );
  NAND2_X1 U6298 ( .A1(n5699), .A2(n4612), .ZN(n4611) );
  NAND2_X1 U6299 ( .A1(n4617), .A2(n4607), .ZN(n9131) );
  NAND2_X1 U6300 ( .A1(n4611), .A2(n4608), .ZN(n4607) );
  AOI21_X1 U6301 ( .B1(n4615), .B2(n4614), .A(n9217), .ZN(n4609) );
  INV_X1 U6302 ( .A(n4615), .ZN(n4610) );
  NAND2_X1 U6303 ( .A1(n7621), .A2(n4632), .ZN(n4628) );
  OAI211_X1 U6304 ( .C1(n7691), .C2(n4633), .A(n4628), .B(n4629), .ZN(n5877)
         );
  NAND2_X1 U6305 ( .A1(n7256), .A2(n4637), .ZN(n4636) );
  NAND2_X1 U6306 ( .A1(n9323), .A2(n5984), .ZN(n4641) );
  OR2_X1 U6307 ( .A1(n8990), .A2(n8989), .ZN(n4648) );
  NAND2_X1 U6308 ( .A1(n8990), .A2(n4454), .ZN(n4645) );
  INV_X1 U6309 ( .A(n8961), .ZN(n4646) );
  NAND2_X1 U6310 ( .A1(n5195), .A2(n5194), .ZN(n4649) );
  NAND2_X1 U6311 ( .A1(n5183), .A2(n5182), .ZN(n4650) );
  MUX2_X1 U6312 ( .A(n6552), .B(n6557), .S(n6549), .Z(n5162) );
  MUX2_X1 U6313 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n6549), .Z(n5184) );
  NAND2_X1 U6314 ( .A1(n5238), .A2(n4657), .ZN(n4656) );
  OAI21_X1 U6315 ( .B1(n8332), .B2(n4670), .A(n4667), .ZN(n4666) );
  NAND2_X1 U6316 ( .A1(n8332), .A2(n4668), .ZN(n4667) );
  NAND3_X1 U6317 ( .A1(n4682), .A2(n4680), .A3(n4678), .ZN(n4861) );
  NAND4_X1 U6318 ( .A1(n8219), .A2(n4480), .A3(n8220), .A4(n8221), .ZN(n4688)
         );
  NAND2_X1 U6319 ( .A1(n4558), .A2(n4525), .ZN(n4693) );
  NAND2_X1 U6320 ( .A1(n5307), .A2(n4708), .ZN(n4707) );
  OAI21_X1 U6321 ( .B1(n4558), .B2(n4710), .A(n5310), .ZN(n5333) );
  INV_X1 U6322 ( .A(n7674), .ZN(n4714) );
  NAND2_X1 U6323 ( .A1(n4711), .A2(n4712), .ZN(n7705) );
  NAND2_X1 U6324 ( .A1(n7674), .A2(n8156), .ZN(n4711) );
  NAND2_X1 U6325 ( .A1(n8598), .A2(n4717), .ZN(n4716) );
  NAND3_X1 U6326 ( .A1(n5062), .A2(n4727), .A3(n4726), .ZN(n6532) );
  NAND2_X1 U6327 ( .A1(n4728), .A2(n4730), .ZN(n6332) );
  NAND2_X1 U6328 ( .A1(n8671), .A2(n4729), .ZN(n4728) );
  INV_X1 U6329 ( .A(n4738), .ZN(n4740) );
  AND2_X1 U6330 ( .A1(n4740), .A2(n4739), .ZN(n4743) );
  NAND2_X2 U6331 ( .A1(n4438), .A2(n6472), .ZN(n6074) );
  NAND2_X2 U6332 ( .A1(n6074), .A2(n4436), .ZN(n8133) );
  NAND2_X1 U6333 ( .A1(n4745), .A2(n4744), .ZN(n7117) );
  AOI21_X1 U6334 ( .B1(n6961), .B2(n4747), .A(n4746), .ZN(n4744) );
  NAND3_X1 U6335 ( .A1(n7105), .A2(n7103), .A3(n6961), .ZN(n4745) );
  NAND2_X1 U6336 ( .A1(n7105), .A2(n7103), .ZN(n7104) );
  NAND2_X2 U6337 ( .A1(n6584), .A2(n6549), .ZN(n9075) );
  NAND2_X1 U6338 ( .A1(n7901), .A2(n5708), .ZN(n4760) );
  AND2_X2 U6339 ( .A1(n9624), .A2(n9185), .ZN(n9592) );
  OR2_X2 U6340 ( .A1(n5728), .A2(n4956), .ZN(n5098) );
  OR2_X2 U6341 ( .A1(n8402), .A2(n8401), .ZN(n8430) );
  NOR2_X1 U6342 ( .A1(n8398), .A2(n8399), .ZN(n8402) );
  MUX2_X1 U6343 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6078), .S(n6737), .Z(n10402)
         );
  NAND2_X1 U6344 ( .A1(n4780), .A2(n4779), .ZN(n6850) );
  INV_X1 U6345 ( .A(n4788), .ZN(n7176) );
  NAND2_X1 U6346 ( .A1(n7177), .A2(n7180), .ZN(n4787) );
  NAND2_X1 U6347 ( .A1(n4794), .A2(n7758), .ZN(n6489) );
  AOI21_X1 U6348 ( .B1(n4795), .B2(n6484), .A(n6209), .ZN(n4793) );
  XNOR2_X1 U6349 ( .A(n6490), .B(P2_B_REG_SCAN_IN), .ZN(n4794) );
  AND2_X1 U6350 ( .A1(n5055), .A2(n6036), .ZN(n4796) );
  INV_X1 U6351 ( .A(n6420), .ZN(n6038) );
  NAND3_X1 U6352 ( .A1(n4448), .A2(n6163), .A3(n4796), .ZN(n6420) );
  NAND2_X1 U6353 ( .A1(n8063), .A2(n4801), .ZN(n4799) );
  NAND2_X1 U6354 ( .A1(n8098), .A2(n4810), .ZN(n4809) );
  OAI211_X1 U6355 ( .C1(n8098), .C2(n4811), .A(n7948), .B(n4809), .ZN(P2_U3160) );
  NAND2_X1 U6356 ( .A1(n8098), .A2(n8091), .ZN(n7968) );
  NAND2_X1 U6357 ( .A1(n4821), .A2(n4463), .ZN(n7597) );
  NAND2_X1 U6358 ( .A1(n7975), .A2(n4824), .ZN(n4823) );
  AND2_X1 U6359 ( .A1(n7909), .A2(n8743), .ZN(n4827) );
  NAND3_X1 U6360 ( .A1(n7995), .A2(n4830), .A3(n7011), .ZN(n7043) );
  INV_X1 U6361 ( .A(n7014), .ZN(n4830) );
  XNOR2_X1 U6362 ( .A(n7039), .B(n7998), .ZN(n7014) );
  NAND2_X1 U6363 ( .A1(n4832), .A2(n4831), .ZN(n6879) );
  NAND3_X1 U6364 ( .A1(n4833), .A2(n8595), .A3(n8050), .ZN(n7984) );
  NAND2_X1 U6365 ( .A1(n7932), .A2(n7931), .ZN(n8050) );
  NAND2_X1 U6366 ( .A1(n4833), .A2(n8050), .ZN(n7985) );
  NAND2_X2 U6367 ( .A1(n5277), .A2(n5276), .ZN(n9919) );
  NAND2_X1 U6368 ( .A1(n4855), .A2(n5146), .ZN(n5161) );
  AND2_X2 U6369 ( .A1(n9566), .A2(n9567), .ZN(n9544) );
  NOR2_X2 U6370 ( .A1(n7893), .A2(n9676), .ZN(n9566) );
  INV_X1 U6371 ( .A(n5072), .ZN(n5147) );
  NOR2_X2 U6372 ( .A1(n9823), .A2(n9904), .ZN(n9821) );
  NAND2_X1 U6373 ( .A1(n4840), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4839) );
  NAND2_X1 U6374 ( .A1(n5726), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4840) );
  NAND2_X1 U6375 ( .A1(n4841), .A2(n4524), .ZN(n5726) );
  INV_X1 U6376 ( .A(n5728), .ZN(n4841) );
  INV_X1 U6377 ( .A(n4848), .ZN(n5693) );
  NAND2_X1 U6378 ( .A1(n5143), .A2(n5142), .ZN(n4855) );
  NAND2_X1 U6379 ( .A1(n5123), .A2(n5122), .ZN(n4856) );
  NAND3_X1 U6380 ( .A1(n4864), .A2(n4858), .A3(n8272), .ZN(n4857) );
  NAND2_X1 U6381 ( .A1(n5214), .A2(n5213), .ZN(n4871) );
  INV_X1 U6382 ( .A(n5458), .ZN(n4886) );
  INV_X2 U6383 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4894) );
  NAND3_X1 U6384 ( .A1(n4900), .A2(n4899), .A3(n4528), .ZN(n6854) );
  NAND2_X1 U6385 ( .A1(n6729), .A2(n4902), .ZN(n4900) );
  NAND2_X1 U6386 ( .A1(n6785), .A2(n6714), .ZN(n4901) );
  INV_X1 U6387 ( .A(n6785), .ZN(n4903) );
  OAI21_X1 U6388 ( .B1(n6729), .B2(n4903), .A(n4902), .ZN(n6853) );
  NAND2_X1 U6389 ( .A1(n7417), .A2(n4465), .ZN(n4909) );
  OAI211_X1 U6390 ( .C1(n7417), .C2(n4911), .A(n4910), .B(n4909), .ZN(n7531)
         );
  NAND2_X1 U6391 ( .A1(n4926), .A2(n4924), .ZN(n5550) );
  NAND2_X1 U6392 ( .A1(n4928), .A2(n4927), .ZN(n5330) );
  AND2_X1 U6393 ( .A1(n4490), .A2(n5305), .ZN(n4927) );
  NAND2_X1 U6394 ( .A1(n4929), .A2(n4930), .ZN(n5677) );
  NAND2_X1 U6395 ( .A1(n9509), .A2(n4931), .ZN(n4929) );
  NAND2_X1 U6396 ( .A1(n9509), .A2(n9508), .ZN(n9507) );
  NAND2_X1 U6397 ( .A1(n4934), .A2(n4935), .ZN(n5457) );
  NAND2_X1 U6398 ( .A1(n7804), .A2(n5439), .ZN(n4934) );
  OAI21_X1 U6399 ( .B1(n7499), .B2(n5351), .A(n5352), .ZN(n7661) );
  NOR2_X2 U6400 ( .A1(n5728), .A2(n4954), .ZN(n5086) );
  NAND3_X1 U6401 ( .A1(n4959), .A2(n5794), .A3(n4958), .ZN(n6991) );
  NAND3_X1 U6402 ( .A1(n6833), .A2(n6937), .A3(n6834), .ZN(n4959) );
  INV_X1 U6403 ( .A(n5787), .ZN(n4960) );
  NAND2_X1 U6404 ( .A1(n6992), .A2(n5805), .ZN(n5814) );
  NAND2_X1 U6405 ( .A1(n6992), .A2(n4464), .ZN(n7147) );
  NAND2_X1 U6406 ( .A1(n5465), .A2(n4967), .ZN(n4965) );
  NAND2_X2 U6407 ( .A1(n4971), .A2(n6539), .ZN(n5827) );
  NAND2_X1 U6408 ( .A1(n8998), .A2(n4979), .ZN(n4977) );
  NAND2_X1 U6409 ( .A1(n4977), .A2(n4978), .ZN(n8990) );
  OAI211_X1 U6410 ( .C1(n8960), .C2(n4991), .A(n4985), .B(n4527), .ZN(P1_U3214) );
  NAND2_X1 U6411 ( .A1(n8960), .A2(n4989), .ZN(n4985) );
  NAND2_X1 U6412 ( .A1(n6908), .A2(n7108), .ZN(n6427) );
  NAND2_X1 U6413 ( .A1(n8353), .A2(n6882), .ZN(n8186) );
  NAND3_X1 U6414 ( .A1(n6954), .A2(n6955), .A3(n7120), .ZN(n4996) );
  NAND3_X1 U6415 ( .A1(n6428), .A2(n4997), .A3(n4996), .ZN(n7119) );
  NAND2_X1 U6416 ( .A1(n4998), .A2(n8306), .ZN(n6953) );
  NAND2_X1 U6417 ( .A1(n5001), .A2(n5003), .ZN(n6465) );
  NAND2_X1 U6418 ( .A1(n6457), .A2(n5004), .ZN(n5001) );
  INV_X1 U6419 ( .A(n7246), .ZN(n5008) );
  NAND2_X1 U6420 ( .A1(n5007), .A2(n5009), .ZN(n7246) );
  NAND2_X1 U6421 ( .A1(n7092), .A2(n5010), .ZN(n5007) );
  NAND2_X1 U6422 ( .A1(n7056), .A2(n7099), .ZN(n5009) );
  OR2_X1 U6423 ( .A1(n7056), .A2(n7099), .ZN(n5010) );
  NAND2_X1 U6424 ( .A1(n4428), .A2(n5014), .ZN(n5011) );
  OAI211_X1 U6425 ( .C1(n4428), .C2(n5016), .A(n5011), .B(n5012), .ZN(n6471)
         );
  OAI21_X1 U6426 ( .B1(n8712), .B2(n5034), .A(n5032), .ZN(n6456) );
  AND2_X1 U6427 ( .A1(n8803), .A2(n8729), .ZN(n5046) );
  NAND2_X1 U6428 ( .A1(n8581), .A2(n5049), .ZN(n5047) );
  NAND3_X1 U6429 ( .A1(n6164), .A2(n4448), .A3(n6178), .ZN(n6286) );
  NAND2_X1 U6430 ( .A1(n5416), .A2(n5415), .ZN(n7804) );
  AOI21_X2 U6431 ( .B1(n7059), .B2(n7058), .A(n7057), .ZN(n7061) );
  NAND2_X1 U6433 ( .A1(n6539), .A2(n6537), .ZN(n9304) );
  NAND4_X1 U6434 ( .A1(n5110), .A2(n5109), .A3(n5108), .A4(n5107), .ZN(n5768)
         );
  OR2_X1 U6435 ( .A1(n7141), .A2(n5795), .ZN(n5769) );
  NAND2_X1 U6436 ( .A1(n6058), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6056) );
  INV_X1 U6437 ( .A(n6050), .ZN(n6048) );
  OAI22_X2 U6438 ( .A1(n9595), .A2(n5477), .B1(n9609), .B2(n9313), .ZN(n9579)
         );
  AND2_X1 U6439 ( .A1(n6516), .A2(n6515), .ZN(n10062) );
  OR2_X1 U6440 ( .A1(n9322), .A2(n9872), .ZN(n5058) );
  OR2_X1 U6441 ( .A1(n7083), .A2(n7082), .ZN(n5059) );
  INV_X1 U6442 ( .A(n10075), .ZN(n6533) );
  AND3_X1 U6443 ( .A1(n6023), .A2(n9031), .A3(n6022), .ZN(n5060) );
  OR2_X1 U6444 ( .A1(n7959), .A2(n8864), .ZN(n5061) );
  OR2_X1 U6445 ( .A1(n7964), .A2(n10045), .ZN(n5062) );
  OR2_X1 U6446 ( .A1(n7959), .A2(n8785), .ZN(n5063) );
  OR2_X1 U6447 ( .A1(n9983), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5064) );
  NAND2_X1 U6448 ( .A1(n7286), .A2(n7285), .ZN(n7555) );
  INV_X1 U6449 ( .A(n8315), .ZN(n6182) );
  AND2_X1 U6450 ( .A1(n5289), .A2(n5270), .ZN(n5065) );
  INV_X1 U6451 ( .A(n8284), .ZN(n8279) );
  INV_X1 U6452 ( .A(n6936), .ZN(n6075) );
  OR2_X1 U6453 ( .A1(n6584), .A2(n6607), .ZN(n5066) );
  INV_X1 U6454 ( .A(n7587), .ZN(n8373) );
  AND2_X1 U6455 ( .A1(n6213), .A2(n6225), .ZN(n7587) );
  INV_X1 U6456 ( .A(n8345), .ZN(n7708) );
  AND2_X1 U6457 ( .A1(n8643), .A2(n6452), .ZN(n5067) );
  AND2_X1 U6458 ( .A1(n7940), .A2(n8092), .ZN(n5068) );
  CLKBUF_X2 U6459 ( .A(P1_U3973), .Z(n9324) );
  INV_X1 U6460 ( .A(n6458), .ZN(n6460) );
  AND2_X1 U6461 ( .A1(n8919), .A2(n8918), .ZN(n5069) );
  OR2_X1 U6462 ( .A1(n8298), .A2(n8274), .ZN(n8267) );
  INV_X1 U6463 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6031) );
  AND2_X1 U6464 ( .A1(n8676), .A2(n8644), .ZN(n6452) );
  NOR2_X1 U6465 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6034) );
  INV_X1 U6466 ( .A(n7562), .ZN(n7560) );
  AND4_X1 U6467 ( .A1(n5077), .A2(n5076), .A3(n5075), .A4(n5680), .ZN(n5078)
         );
  INV_X1 U6468 ( .A(n8633), .ZN(n6459) );
  INV_X1 U6469 ( .A(n10049), .ZN(n6437) );
  INV_X1 U6470 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6037) );
  INV_X1 U6471 ( .A(n5802), .ZN(n5803) );
  NAND2_X1 U6472 ( .A1(n7929), .A2(n6459), .ZN(n7930) );
  INV_X1 U6473 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8355) );
  INV_X1 U6474 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6169) );
  INV_X1 U6475 ( .A(n8310), .ZN(n6430) );
  OR2_X1 U6476 ( .A1(n6492), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6493) );
  INV_X1 U6477 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6040) );
  NOR2_X1 U6478 ( .A1(n5601), .A2(n8964), .ZN(n5618) );
  AND2_X1 U6479 ( .A1(n9848), .A2(n5984), .ZN(n5767) );
  AND3_X1 U6480 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5204) );
  INV_X1 U6481 ( .A(n9111), .ZN(n9105) );
  INV_X1 U6482 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5321) );
  INV_X1 U6483 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U6484 ( .A1(n5080), .A2(n5079), .ZN(n5081) );
  NOR2_X1 U6485 ( .A1(n5528), .A2(SI_21_), .ZN(n5530) );
  INV_X1 U6486 ( .A(n5394), .ZN(n5395) );
  INV_X1 U6487 ( .A(n7204), .ZN(n7201) );
  INV_X1 U6488 ( .A(n8727), .ZN(n8225) );
  XNOR2_X1 U6489 ( .A(n7177), .B(n7180), .ZN(n7085) );
  NOR2_X1 U6490 ( .A1(n7587), .A2(n8355), .ZN(n8356) );
  INV_X1 U6491 ( .A(n6352), .ZN(n6351) );
  OR2_X1 U6492 ( .A1(n8350), .A2(n7099), .ZN(n8217) );
  AND2_X1 U6493 ( .A1(n8144), .A2(n8533), .ZN(n6770) );
  OR2_X1 U6494 ( .A1(n6184), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n6194) );
  INV_X1 U6495 ( .A(n5884), .ZN(n5885) );
  AND2_X1 U6496 ( .A1(n5952), .A2(n8917), .ZN(n5955) );
  OR2_X1 U6497 ( .A1(n5363), .A2(n5362), .ZN(n5384) );
  INV_X1 U6498 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10141) );
  INV_X1 U6499 ( .A(n9604), .ZN(n9605) );
  INV_X1 U6500 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5755) );
  AND2_X1 U6501 ( .A1(n5716), .A2(n9225), .ZN(n9076) );
  NAND2_X1 U6502 ( .A1(n5421), .A2(SI_16_), .ZN(n5440) );
  OR3_X1 U6503 ( .A1(n5335), .A2(P1_IR_REG_10__SCAN_IN), .A3(
        P1_IR_REG_11__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U6504 ( .A1(n5244), .A2(n5243), .ZN(n5263) );
  INV_X1 U6505 ( .A(n4439), .ZN(n6407) );
  OR2_X1 U6507 ( .A1(n6654), .A2(n7844), .ZN(n6731) );
  OR2_X1 U6508 ( .A1(n6875), .A2(n6921), .ZN(n6525) );
  INV_X1 U6509 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6517) );
  NAND2_X1 U6510 ( .A1(n6423), .A2(n6929), .ZN(n7685) );
  INV_X1 U6511 ( .A(n5654), .ZN(n5652) );
  AND2_X1 U6512 ( .A1(n5977), .A2(n5976), .ZN(n7950) );
  INV_X1 U6513 ( .A(n9298), .ZN(n9233) );
  AND2_X1 U6514 ( .A1(n5505), .A2(n5504), .ZN(n9691) );
  AND4_X1 U6515 ( .A1(n5438), .A2(n5437), .A3(n5436), .A4(n5435), .ZN(n9622)
         );
  OR2_X1 U6516 ( .A1(n6869), .A2(n6868), .ZN(n7032) );
  INV_X1 U6517 ( .A(n9096), .ZN(n9594) );
  AND2_X1 U6518 ( .A1(n7323), .A2(n9126), .ZN(n9809) );
  OR2_X1 U6519 ( .A1(n6803), .A2(n9233), .ZN(n9822) );
  OR2_X1 U6520 ( .A1(n5996), .A2(n4443), .ZN(n9952) );
  OR2_X1 U6521 ( .A1(n9960), .A2(n9225), .ZN(n6002) );
  AND2_X1 U6522 ( .A1(n5610), .A2(n5598), .ZN(n5608) );
  XNOR2_X1 U6523 ( .A(n5397), .B(SI_14_), .ZN(n5394) );
  INV_X1 U6524 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5071) );
  AND2_X1 U6525 ( .A1(n6653), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10411) );
  OR3_X1 U6526 ( .A1(n6928), .A2(n10039), .A3(n6927), .ZN(n8745) );
  INV_X1 U6527 ( .A(n8744), .ZN(n8728) );
  INV_X1 U6528 ( .A(n8745), .ZN(n8718) );
  INV_X1 U6529 ( .A(n8711), .ZN(n8753) );
  AND2_X1 U6530 ( .A1(n10075), .A2(n10020), .ZN(n8809) );
  AND2_X1 U6531 ( .A1(n6530), .A2(n6529), .ZN(n6531) );
  NAND2_X1 U6532 ( .A1(n7359), .A2(n7453), .ZN(n10039) );
  OR2_X1 U6533 ( .A1(n6775), .A2(n6514), .ZN(n6515) );
  AND2_X1 U6534 ( .A1(n6585), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6537) );
  INV_X1 U6535 ( .A(n8960), .ZN(n9029) );
  AND3_X1 U6536 ( .A1(n5476), .A2(n5475), .A3(n5474), .ZN(n9690) );
  OR2_X1 U6537 ( .A1(n6604), .A2(n9305), .ZN(n9428) );
  INV_X1 U6538 ( .A(n9446), .ZN(n9443) );
  AND2_X1 U6539 ( .A1(n9193), .A2(n5709), .ZN(n9099) );
  INV_X1 U6540 ( .A(n9872), .ZN(n9833) );
  NAND2_X1 U6541 ( .A1(n7131), .A2(n9846), .ZN(n9598) );
  NAND2_X1 U6542 ( .A1(n9814), .A2(n9960), .ZN(n9949) );
  NAND2_X1 U6543 ( .A1(n5715), .A2(n5714), .ZN(n9887) );
  NAND2_X1 U6544 ( .A1(n5741), .A2(n5740), .ZN(n5993) );
  AND2_X1 U6545 ( .A1(n5401), .A2(n5381), .ZN(n7607) );
  AND2_X1 U6546 ( .A1(n5248), .A2(n5223), .ZN(n6676) );
  INV_X1 U6547 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10391) );
  INV_X1 U6548 ( .A(n8585), .ZN(n8837) );
  NAND2_X1 U6549 ( .A1(n6769), .A2(n6768), .ZN(n8039) );
  INV_X1 U6550 ( .A(n8037), .ZN(n8116) );
  OR2_X1 U6551 ( .A1(n8497), .A2(n8334), .ZN(n8535) );
  INV_X1 U6552 ( .A(n10419), .ZN(n10002) );
  NAND2_X1 U6553 ( .A1(n8748), .A2(n6965), .ZN(n8711) );
  INV_X1 U6554 ( .A(n8748), .ZN(n8752) );
  AND2_X2 U6555 ( .A1(n6925), .A2(n6531), .ZN(n10075) );
  XNOR2_X1 U6556 ( .A(n8562), .B(n8563), .ZN(n8829) );
  AND3_X1 U6557 ( .A1(n10031), .A2(n10030), .A3(n10029), .ZN(n10069) );
  INV_X2 U6558 ( .A(n10062), .ZN(n10064) );
  AND2_X1 U6559 ( .A1(n6766), .A2(n6492), .ZN(n6620) );
  INV_X1 U6560 ( .A(n6620), .ZN(n6580) );
  INV_X1 U6561 ( .A(n8337), .ZN(n7453) );
  INV_X1 U6562 ( .A(n7813), .ZN(n9784) );
  INV_X1 U6563 ( .A(n8991), .ZN(n9048) );
  AND2_X1 U6564 ( .A1(n6003), .A2(n9846), .ZN(n9039) );
  INV_X1 U6565 ( .A(n7953), .ZN(n9497) );
  INV_X1 U6566 ( .A(n9681), .ZN(n9312) );
  INV_X1 U6567 ( .A(n9810), .ZN(n9917) );
  OR2_X1 U6568 ( .A1(n6604), .A2(n6812), .ZN(n9446) );
  INV_X1 U6569 ( .A(n9841), .ZN(n9629) );
  INV_X1 U6570 ( .A(n9673), .ZN(n9707) );
  OR3_X1 U6571 ( .A1(n7130), .A2(n5758), .A3(n5995), .ZN(n9981) );
  INV_X2 U6572 ( .A(n9981), .ZN(n9983) );
  INV_X1 U6573 ( .A(n9588), .ZN(n9751) );
  INV_X1 U6574 ( .A(n9741), .ZN(n9754) );
  OR3_X1 U6575 ( .A1(n7130), .A2(n5758), .A3(n7129), .ZN(n9965) );
  NAND2_X1 U6576 ( .A1(n6004), .A2(n5993), .ZN(n9859) );
  NAND2_X1 U6577 ( .A1(n5731), .A2(n5730), .ZN(n7704) );
  INV_X1 U6578 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10178) );
  INV_X1 U6579 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10251) );
  INV_X1 U6580 ( .A(n8497), .ZN(P2_U3893) );
  NOR2_X1 U6581 ( .A1(n6539), .A2(n6538), .ZN(P1_U3973) );
  NOR2_X1 U6582 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5077) );
  NOR2_X1 U6583 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5076) );
  NOR2_X1 U6584 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5075) );
  INV_X1 U6585 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5084) );
  NAND2_X1 U6586 ( .A1(n5086), .A2(n5084), .ZN(n9762) );
  XNOR2_X2 U6587 ( .A(n5085), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5091) );
  INV_X1 U6588 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5088) );
  OR2_X1 U6589 ( .A1(n5346), .A2(n5088), .ZN(n5090) );
  NAND2_X1 U6590 ( .A1(n5091), .A2(n5092), .ZN(n5116) );
  INV_X1 U6591 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9845) );
  OR2_X1 U6592 ( .A1(n5116), .A2(n9845), .ZN(n5089) );
  INV_X1 U6593 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6608) );
  OR2_X1 U6594 ( .A1(n5471), .A2(n6608), .ZN(n5094) );
  NAND2_X1 U6595 ( .A1(n4437), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5093) );
  INV_X1 U6596 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5095) );
  INV_X1 U6597 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6551) );
  AND2_X1 U6598 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5101) );
  AND2_X1 U6599 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5102) );
  NAND2_X1 U6600 ( .A1(n6549), .A2(n5102), .ZN(n6072) );
  NAND2_X1 U6601 ( .A1(n5113), .A2(n6072), .ZN(n5122) );
  XNOR2_X1 U6602 ( .A(n5121), .B(n5122), .ZN(n6060) );
  INV_X1 U6603 ( .A(n6060), .ZN(n6558) );
  NAND2_X1 U6604 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5103) );
  MUX2_X1 U6605 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5103), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5106) );
  INV_X1 U6606 ( .A(n5104), .ZN(n5105) );
  INV_X1 U6607 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7134) );
  OR2_X1 U6608 ( .A1(n4434), .A2(n7134), .ZN(n5109) );
  INV_X1 U6609 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6581) );
  OR2_X1 U6610 ( .A1(n5346), .A2(n6581), .ZN(n5108) );
  INV_X1 U6611 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5771) );
  OR2_X1 U6612 ( .A1(n5471), .A2(n5771), .ZN(n5107) );
  NAND2_X1 U6613 ( .A1(n4436), .A2(SI_0_), .ZN(n5112) );
  INV_X1 U6614 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5111) );
  NAND2_X1 U6615 ( .A1(n5112), .A2(n5111), .ZN(n5114) );
  NAND2_X1 U6616 ( .A1(n5114), .A2(n5113), .ZN(n9772) );
  MUX2_X1 U6617 ( .A(n9333), .B(n9772), .S(n6584), .Z(n7141) );
  INV_X1 U6618 ( .A(n7141), .ZN(n6693) );
  AND2_X1 U6619 ( .A1(n5768), .A2(n6693), .ZN(n6945) );
  INV_X1 U6620 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6606) );
  OR2_X1 U6621 ( .A1(n5471), .A2(n6606), .ZN(n5120) );
  INV_X1 U6622 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6597) );
  OR2_X1 U6623 ( .A1(n5346), .A2(n6597), .ZN(n5118) );
  INV_X1 U6624 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n5115) );
  OR2_X1 U6625 ( .A1(n5116), .A2(n5115), .ZN(n5117) );
  INV_X1 U6626 ( .A(n5121), .ZN(n5123) );
  NAND2_X1 U6627 ( .A1(n5124), .A2(SI_1_), .ZN(n5125) );
  INV_X1 U6628 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6555) );
  INV_X1 U6629 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6553) );
  MUX2_X1 U6630 ( .A(n6555), .B(n6553), .S(n5126), .Z(n5144) );
  XNOR2_X1 U6631 ( .A(n5144), .B(SI_2_), .ZN(n5142) );
  XNOR2_X1 U6632 ( .A(n5143), .B(n5142), .ZN(n6554) );
  OR2_X1 U6633 ( .A1(n5247), .A2(n6554), .ZN(n5130) );
  NOR2_X1 U6634 ( .A1(n5104), .A2(n5198), .ZN(n5127) );
  MUX2_X1 U6635 ( .A(n5198), .B(n5127), .S(P1_IR_REG_2__SCAN_IN), .Z(n5128) );
  INV_X1 U6636 ( .A(n5128), .ZN(n5129) );
  NAND2_X1 U6637 ( .A1(n5129), .A2(n5147), .ZN(n6822) );
  INV_X1 U6638 ( .A(n7300), .ZN(n9865) );
  OR2_X1 U6639 ( .A1(n5762), .A2(n9848), .ZN(n7296) );
  AND2_X1 U6640 ( .A1(n5132), .A2(n7296), .ZN(n5131) );
  NAND2_X1 U6641 ( .A1(n7297), .A2(n5131), .ZN(n5134) );
  OR2_X1 U6642 ( .A1(n9828), .A2(n7300), .ZN(n5697) );
  NAND2_X1 U6643 ( .A1(n4429), .A2(n7300), .ZN(n9240) );
  NAND2_X1 U6644 ( .A1(n7306), .A2(n5132), .ZN(n5133) );
  AND2_X1 U6645 ( .A1(n5134), .A2(n5133), .ZN(n9835) );
  NAND2_X1 U6646 ( .A1(n5135), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5141) );
  INV_X1 U6647 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6598) );
  OR2_X1 U6648 ( .A1(n5346), .A2(n6598), .ZN(n5140) );
  INV_X1 U6649 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5136) );
  OR2_X1 U6650 ( .A1(n5471), .A2(n5136), .ZN(n5139) );
  OR2_X1 U6651 ( .A1(n5116), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5138) );
  INV_X1 U6652 ( .A(n5144), .ZN(n5145) );
  NAND2_X1 U6653 ( .A1(n5145), .A2(SI_2_), .ZN(n5146) );
  INV_X1 U6654 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6557) );
  INV_X1 U6655 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6552) );
  XNOR2_X1 U6656 ( .A(n5162), .B(SI_3_), .ZN(n5160) );
  XNOR2_X1 U6657 ( .A(n5161), .B(n5160), .ZN(n6556) );
  OR2_X1 U6658 ( .A1(n5247), .A2(n6556), .ZN(n5152) );
  OR2_X1 U6659 ( .A1(n9075), .A2(n6552), .ZN(n5151) );
  NAND2_X1 U6660 ( .A1(n5147), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5148) );
  MUX2_X1 U6661 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5148), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n5149) );
  NAND2_X1 U6662 ( .A1(n5149), .A2(n5187), .ZN(n9340) );
  OR2_X1 U6663 ( .A1(n6584), .A2(n9340), .ZN(n5150) );
  AND3_X2 U6664 ( .A1(n5152), .A2(n5151), .A3(n5150), .ZN(n9872) );
  NAND2_X1 U6665 ( .A1(n9322), .A2(n9872), .ZN(n9239) );
  NAND2_X1 U6666 ( .A1(n9835), .A2(n9834), .ZN(n5154) );
  OR2_X1 U6667 ( .A1(n9322), .A2(n9833), .ZN(n5153) );
  NAND2_X1 U6668 ( .A1(n5154), .A2(n5153), .ZN(n7310) );
  NAND2_X1 U6669 ( .A1(n5135), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5159) );
  INV_X1 U6670 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5155) );
  OR2_X1 U6671 ( .A1(n5471), .A2(n5155), .ZN(n5158) );
  XNOR2_X1 U6672 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7312) );
  OR2_X1 U6673 ( .A1(n4434), .A2(n7312), .ZN(n5157) );
  INV_X1 U6674 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6599) );
  OR2_X1 U6675 ( .A1(n5346), .A2(n6599), .ZN(n5156) );
  NAND2_X1 U6676 ( .A1(n5161), .A2(n5160), .ZN(n5165) );
  INV_X1 U6677 ( .A(n5162), .ZN(n5163) );
  NAND2_X1 U6678 ( .A1(n5163), .A2(SI_3_), .ZN(n5164) );
  INV_X1 U6679 ( .A(SI_4_), .ZN(n5166) );
  XNOR2_X1 U6680 ( .A(n5184), .B(n5166), .ZN(n5182) );
  XNOR2_X1 U6681 ( .A(n5183), .B(n5182), .ZN(n6568) );
  OR2_X1 U6682 ( .A1(n5247), .A2(n6568), .ZN(n5172) );
  INV_X1 U6683 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5167) );
  OR2_X1 U6684 ( .A1(n9075), .A2(n5167), .ZN(n5171) );
  NAND2_X1 U6685 ( .A1(n5187), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5169) );
  INV_X1 U6686 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5168) );
  XNOR2_X1 U6687 ( .A(n5169), .B(n5168), .ZN(n9353) );
  OR2_X1 U6688 ( .A1(n6584), .A2(n9353), .ZN(n5170) );
  OR2_X1 U6690 ( .A1(n9829), .A2(n7316), .ZN(n9127) );
  NAND2_X1 U6691 ( .A1(n9829), .A2(n7316), .ZN(n9235) );
  NAND2_X1 U6692 ( .A1(n9127), .A2(n9235), .ZN(n9082) );
  NAND2_X1 U6693 ( .A1(n7310), .A2(n9082), .ZN(n5174) );
  INV_X1 U6694 ( .A(n7316), .ZN(n9881) );
  OR2_X1 U6695 ( .A1(n9829), .A2(n9881), .ZN(n5173) );
  NAND2_X1 U6696 ( .A1(n5174), .A2(n5173), .ZN(n7159) );
  NAND2_X1 U6697 ( .A1(n5135), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5181) );
  INV_X1 U6698 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6600) );
  OR2_X1 U6699 ( .A1(n5545), .A2(n6600), .ZN(n5180) );
  INV_X1 U6700 ( .A(n5204), .ZN(n5205) );
  INV_X1 U6701 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U6702 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5175) );
  NAND2_X1 U6703 ( .A1(n5176), .A2(n5175), .ZN(n5177) );
  NAND2_X1 U6704 ( .A1(n5205), .A2(n5177), .ZN(n7152) );
  OR2_X1 U6705 ( .A1(n5434), .A2(n7152), .ZN(n5179) );
  INV_X1 U6706 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6611) );
  OR2_X1 U6707 ( .A1(n5471), .A2(n6611), .ZN(n5178) );
  NAND2_X1 U6708 ( .A1(n5184), .A2(SI_4_), .ZN(n5185) );
  MUX2_X1 U6709 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n4435), .Z(n5196) );
  INV_X1 U6710 ( .A(SI_5_), .ZN(n5186) );
  XNOR2_X1 U6711 ( .A(n5196), .B(n5186), .ZN(n5194) );
  XNOR2_X1 U6712 ( .A(n5195), .B(n5194), .ZN(n6560) );
  OR2_X1 U6713 ( .A1(n6560), .A2(n5247), .ZN(n5191) );
  NOR2_X1 U6714 ( .A1(n5187), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5274) );
  OR2_X1 U6715 ( .A1(n5274), .A2(n5198), .ZN(n5219) );
  NAND2_X1 U6716 ( .A1(n5219), .A2(n5188), .ZN(n5199) );
  OAI21_X1 U6717 ( .B1(n5219), .B2(n5188), .A(n5199), .ZN(n9366) );
  OR2_X1 U6718 ( .A1(n6584), .A2(n9366), .ZN(n5190) );
  INV_X1 U6719 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6559) );
  OR2_X1 U6720 ( .A1(n9075), .A2(n6559), .ZN(n5189) );
  NAND2_X1 U6721 ( .A1(n9321), .A2(n5806), .ZN(n9249) );
  NAND2_X1 U6722 ( .A1(n7159), .A2(n9083), .ZN(n5193) );
  OR2_X1 U6723 ( .A1(n9321), .A2(n9889), .ZN(n5192) );
  NAND2_X1 U6724 ( .A1(n5193), .A2(n5192), .ZN(n7222) );
  NAND2_X1 U6725 ( .A1(n5196), .A2(SI_5_), .ZN(n5197) );
  INV_X1 U6726 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6564) );
  MUX2_X1 U6727 ( .A(n6562), .B(n6564), .S(n4436), .Z(n5215) );
  XNOR2_X1 U6728 ( .A(n5215), .B(SI_6_), .ZN(n5213) );
  XNOR2_X1 U6729 ( .A(n5214), .B(n5213), .ZN(n6563) );
  OR2_X1 U6730 ( .A1(n6563), .A2(n5247), .ZN(n5202) );
  NAND2_X1 U6731 ( .A1(n5199), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5200) );
  XNOR2_X1 U6732 ( .A(n5200), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6629) );
  AOI22_X1 U6733 ( .A1(n5483), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5482), .B2(
        n6629), .ZN(n5201) );
  INV_X1 U6734 ( .A(n5471), .ZN(n5582) );
  NAND2_X1 U6735 ( .A1(n5582), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5210) );
  INV_X1 U6736 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5203) );
  OR2_X1 U6737 ( .A1(n5585), .A2(n5203), .ZN(n5209) );
  NAND2_X1 U6738 ( .A1(n5204), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5227) );
  INV_X1 U6739 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U6740 ( .A1(n5205), .A2(n6603), .ZN(n5206) );
  NAND2_X1 U6741 ( .A1(n5227), .A2(n5206), .ZN(n7263) );
  OR2_X1 U6742 ( .A1(n5671), .A2(n7263), .ZN(n5208) );
  INV_X1 U6743 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7225) );
  OR2_X1 U6744 ( .A1(n5545), .A2(n7225), .ZN(n5207) );
  NAND4_X1 U6745 ( .A1(n5210), .A2(n5209), .A3(n5208), .A4(n5207), .ZN(n9890)
         );
  OR2_X1 U6746 ( .A1(n9899), .A2(n9890), .ZN(n9133) );
  NAND2_X1 U6747 ( .A1(n9899), .A2(n9890), .ZN(n9126) );
  NAND2_X1 U6748 ( .A1(n9133), .A2(n9126), .ZN(n7223) );
  NAND2_X1 U6749 ( .A1(n7222), .A2(n7223), .ZN(n5212) );
  INV_X1 U6750 ( .A(n9890), .ZN(n9811) );
  NAND2_X1 U6751 ( .A1(n9811), .A2(n9899), .ZN(n5211) );
  NAND2_X1 U6752 ( .A1(n5212), .A2(n5211), .ZN(n9812) );
  INV_X1 U6753 ( .A(n5215), .ZN(n5216) );
  NAND2_X1 U6754 ( .A1(n5216), .A2(SI_6_), .ZN(n5217) );
  MUX2_X1 U6755 ( .A(n6565), .B(n6567), .S(n4435), .Z(n5239) );
  XNOR2_X1 U6756 ( .A(n5239), .B(SI_7_), .ZN(n5237) );
  XNOR2_X1 U6757 ( .A(n5238), .B(n5237), .ZN(n6566) );
  OR2_X1 U6758 ( .A1(n6566), .A2(n5247), .ZN(n5225) );
  NOR2_X1 U6759 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5272) );
  OR2_X1 U6760 ( .A1(n5272), .A2(n5198), .ZN(n5218) );
  INV_X1 U6761 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5220) );
  NAND2_X1 U6762 ( .A1(n5221), .A2(n5220), .ZN(n5248) );
  INV_X1 U6763 ( .A(n5221), .ZN(n5222) );
  NAND2_X1 U6764 ( .A1(n5222), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5223) );
  AOI22_X1 U6765 ( .A1(n5483), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5482), .B2(
        n6676), .ZN(n5224) );
  NAND2_X1 U6766 ( .A1(n5135), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5233) );
  INV_X1 U6767 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6633) );
  OR2_X1 U6768 ( .A1(n5471), .A2(n6633), .ZN(n5232) );
  INV_X1 U6769 ( .A(n5253), .ZN(n5254) );
  NAND2_X1 U6770 ( .A1(n5227), .A2(n5226), .ZN(n5228) );
  NAND2_X1 U6771 ( .A1(n5254), .A2(n5228), .ZN(n9818) );
  OR2_X1 U6772 ( .A1(n5671), .A2(n9818), .ZN(n5231) );
  INV_X1 U6773 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5229) );
  OR2_X1 U6774 ( .A1(n5545), .A2(n5229), .ZN(n5230) );
  OR2_X1 U6775 ( .A1(n9904), .A2(n7623), .ZN(n9135) );
  NAND2_X1 U6776 ( .A1(n9904), .A2(n7623), .ZN(n7379) );
  NAND2_X1 U6777 ( .A1(n9135), .A2(n7379), .ZN(n9138) );
  NAND2_X1 U6778 ( .A1(n9812), .A2(n9138), .ZN(n5236) );
  INV_X1 U6779 ( .A(n9904), .ZN(n5234) );
  NAND2_X1 U6780 ( .A1(n5234), .A2(n7623), .ZN(n5235) );
  NAND2_X1 U6781 ( .A1(n5236), .A2(n5235), .ZN(n7375) );
  INV_X1 U6782 ( .A(n5239), .ZN(n5240) );
  NAND2_X1 U6783 ( .A1(n5240), .A2(SI_7_), .ZN(n5241) );
  INV_X1 U6784 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5242) );
  MUX2_X1 U6785 ( .A(n6573), .B(n5242), .S(n4435), .Z(n5244) );
  INV_X1 U6786 ( .A(SI_8_), .ZN(n5243) );
  INV_X1 U6787 ( .A(n5244), .ZN(n5245) );
  NAND2_X1 U6788 ( .A1(n5245), .A2(SI_8_), .ZN(n5246) );
  NAND2_X1 U6789 ( .A1(n5263), .A2(n5246), .ZN(n5264) );
  NAND2_X1 U6790 ( .A1(n6570), .A2(n5443), .ZN(n5251) );
  NAND2_X1 U6791 ( .A1(n5248), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5249) );
  XNOR2_X1 U6792 ( .A(n5249), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6703) );
  AOI22_X1 U6793 ( .A1(n5483), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5482), .B2(
        n6703), .ZN(n5250) );
  NAND2_X1 U6794 ( .A1(n5135), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5260) );
  INV_X1 U6795 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5252) );
  OR2_X1 U6796 ( .A1(n5545), .A2(n5252), .ZN(n5259) );
  NAND2_X1 U6797 ( .A1(n5253), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5279) );
  INV_X1 U6798 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6681) );
  NAND2_X1 U6799 ( .A1(n5254), .A2(n6681), .ZN(n5255) );
  NAND2_X1 U6800 ( .A1(n5279), .A2(n5255), .ZN(n7386) );
  OR2_X1 U6801 ( .A1(n5434), .A2(n7386), .ZN(n5258) );
  INV_X1 U6802 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5256) );
  OR2_X1 U6803 ( .A1(n6670), .A2(n5256), .ZN(n5257) );
  NAND2_X1 U6804 ( .A1(n7387), .A2(n9810), .ZN(n9143) );
  NAND2_X1 U6805 ( .A1(n9136), .A2(n9143), .ZN(n7377) );
  NAND2_X1 U6806 ( .A1(n7375), .A2(n7377), .ZN(n5262) );
  OR2_X1 U6807 ( .A1(n7387), .A2(n9917), .ZN(n5261) );
  NAND2_X1 U6808 ( .A1(n5262), .A2(n5261), .ZN(n7331) );
  INV_X1 U6809 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5266) );
  MUX2_X1 U6810 ( .A(n5266), .B(n10178), .S(n4436), .Z(n5268) );
  INV_X1 U6811 ( .A(SI_9_), .ZN(n5267) );
  INV_X1 U6812 ( .A(n5268), .ZN(n5269) );
  NAND2_X1 U6813 ( .A1(n5269), .A2(SI_9_), .ZN(n5270) );
  NAND2_X1 U6814 ( .A1(n6574), .A2(n5443), .ZN(n5277) );
  NOR2_X1 U6815 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5271) );
  AND2_X1 U6816 ( .A1(n5272), .A2(n5271), .ZN(n5273) );
  AND2_X1 U6817 ( .A1(n5274), .A2(n5273), .ZN(n5292) );
  OR2_X1 U6818 ( .A1(n5292), .A2(n5198), .ZN(n5275) );
  XNOR2_X1 U6819 ( .A(n5275), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6866) );
  AOI22_X1 U6820 ( .A1(n5483), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5482), .B2(
        n6866), .ZN(n5276) );
  NAND2_X1 U6821 ( .A1(n5135), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5285) );
  INV_X1 U6822 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6698) );
  OR2_X1 U6823 ( .A1(n5545), .A2(n6698), .ZN(n5284) );
  NAND2_X1 U6824 ( .A1(n5279), .A2(n5278), .ZN(n5280) );
  NAND2_X1 U6825 ( .A1(n5299), .A2(n5280), .ZN(n7695) );
  OR2_X1 U6826 ( .A1(n5434), .A2(n7695), .ZN(n5283) );
  INV_X1 U6827 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5281) );
  OR2_X1 U6828 ( .A1(n6670), .A2(n5281), .ZN(n5282) );
  NAND2_X1 U6829 ( .A1(n9919), .A2(n9927), .ZN(n9148) );
  NAND2_X1 U6830 ( .A1(n9156), .A2(n9148), .ZN(n7332) );
  NAND2_X1 U6831 ( .A1(n7331), .A2(n7332), .ZN(n5287) );
  INV_X1 U6832 ( .A(n9927), .ZN(n9319) );
  OR2_X1 U6833 ( .A1(n9919), .A2(n9319), .ZN(n5286) );
  NAND2_X1 U6834 ( .A1(n5287), .A2(n5286), .ZN(n7344) );
  INV_X1 U6835 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5290) );
  MUX2_X1 U6836 ( .A(n10249), .B(n5290), .S(n4436), .Z(n5308) );
  XNOR2_X1 U6837 ( .A(n4558), .B(n5306), .ZN(n6578) );
  NAND2_X1 U6838 ( .A1(n6578), .A2(n5443), .ZN(n5297) );
  INV_X1 U6839 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6840 ( .A1(n5292), .A2(n5291), .ZN(n5335) );
  NAND2_X1 U6841 ( .A1(n5335), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U6842 ( .A1(n5294), .A2(n5293), .ZN(n5316) );
  OR2_X1 U6843 ( .A1(n5294), .A2(n5293), .ZN(n5295) );
  AOI22_X1 U6844 ( .A1(n5483), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5482), .B2(
        n7029), .ZN(n5296) );
  NAND2_X2 U6845 ( .A1(n5297), .A2(n5296), .ZN(n9930) );
  NAND2_X1 U6846 ( .A1(n5582), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5304) );
  INV_X1 U6847 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5298) );
  OR2_X1 U6848 ( .A1(n5585), .A2(n5298), .ZN(n5303) );
  NAND2_X1 U6849 ( .A1(n5299), .A2(n10141), .ZN(n5300) );
  NAND2_X1 U6850 ( .A1(n5322), .A2(n5300), .ZN(n7776) );
  OR2_X1 U6851 ( .A1(n5671), .A2(n7776), .ZN(n5302) );
  INV_X1 U6852 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7338) );
  OR2_X1 U6853 ( .A1(n5545), .A2(n7338), .ZN(n5301) );
  OR2_X1 U6854 ( .A1(n9930), .A2(n9792), .ZN(n9251) );
  NAND2_X1 U6855 ( .A1(n9930), .A2(n9792), .ZN(n9794) );
  INV_X1 U6856 ( .A(n9792), .ZN(n9318) );
  OR2_X1 U6857 ( .A1(n9930), .A2(n9318), .ZN(n5305) );
  INV_X1 U6858 ( .A(n5308), .ZN(n5309) );
  NAND2_X1 U6859 ( .A1(n5309), .A2(SI_10_), .ZN(n5310) );
  INV_X1 U6860 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5311) );
  MUX2_X1 U6861 ( .A(n6689), .B(n5311), .S(n4436), .Z(n5313) );
  INV_X1 U6862 ( .A(SI_11_), .ZN(n5312) );
  INV_X1 U6863 ( .A(n5313), .ZN(n5314) );
  NAND2_X1 U6864 ( .A1(n5314), .A2(SI_11_), .ZN(n5315) );
  NAND2_X1 U6865 ( .A1(n5331), .A2(n5315), .ZN(n5332) );
  XNOR2_X1 U6866 ( .A(n5333), .B(n5332), .ZN(n6662) );
  NAND2_X1 U6867 ( .A1(n6662), .A2(n5443), .ZN(n5319) );
  NAND2_X1 U6868 ( .A1(n5316), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5317) );
  XNOR2_X1 U6869 ( .A(n5317), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7237) );
  AOI22_X1 U6870 ( .A1(n5483), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5482), .B2(
        n7237), .ZN(n5318) );
  NAND2_X1 U6871 ( .A1(n5135), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5328) );
  INV_X1 U6872 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5320) );
  OR2_X1 U6873 ( .A1(n6670), .A2(n5320), .ZN(n5327) );
  INV_X1 U6874 ( .A(n5343), .ZN(n5344) );
  NAND2_X1 U6875 ( .A1(n5322), .A2(n5321), .ZN(n5323) );
  NAND2_X1 U6876 ( .A1(n5344), .A2(n5323), .ZN(n9800) );
  OR2_X1 U6877 ( .A1(n5671), .A2(n9800), .ZN(n5326) );
  INV_X1 U6878 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5324) );
  OR2_X1 U6879 ( .A1(n5545), .A2(n5324), .ZN(n5325) );
  INV_X1 U6880 ( .A(n9926), .ZN(n9317) );
  NAND2_X1 U6881 ( .A1(n9802), .A2(n9317), .ZN(n5329) );
  INV_X1 U6882 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5334) );
  MUX2_X1 U6883 ( .A(n6751), .B(n5334), .S(n4436), .Z(n5354) );
  NAND2_X1 U6884 ( .A1(n6696), .A2(n5443), .ZN(n5341) );
  NAND2_X1 U6885 ( .A1(n5338), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5336) );
  MUX2_X1 U6886 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5336), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5337) );
  INV_X1 U6887 ( .A(n5337), .ZN(n5339) );
  AOI22_X1 U6888 ( .A1(n5483), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5482), .B2(
        n7275), .ZN(n5340) );
  NAND2_X1 U6889 ( .A1(n4437), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5350) );
  INV_X1 U6890 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5342) );
  OR2_X1 U6891 ( .A1(n5471), .A2(n5342), .ZN(n5349) );
  NAND2_X1 U6892 ( .A1(n5343), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5363) );
  INV_X1 U6893 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7235) );
  NAND2_X1 U6894 ( .A1(n5344), .A2(n7235), .ZN(n5345) );
  NAND2_X1 U6895 ( .A1(n5363), .A2(n5345), .ZN(n7506) );
  OR2_X1 U6896 ( .A1(n5671), .A2(n7506), .ZN(n5348) );
  INV_X1 U6897 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7238) );
  OR2_X1 U6898 ( .A1(n5545), .A2(n7238), .ZN(n5347) );
  NAND2_X1 U6899 ( .A1(n7527), .A2(n9793), .ZN(n9258) );
  NAND2_X1 U6900 ( .A1(n9163), .A2(n9258), .ZN(n9090) );
  INV_X1 U6901 ( .A(n9090), .ZN(n5351) );
  INV_X1 U6902 ( .A(n9793), .ZN(n9316) );
  OR2_X1 U6903 ( .A1(n7527), .A2(n9316), .ZN(n5352) );
  INV_X1 U6904 ( .A(n5354), .ZN(n5355) );
  NAND2_X1 U6905 ( .A1(n5355), .A2(SI_12_), .ZN(n5356) );
  MUX2_X1 U6906 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4436), .Z(n5373) );
  XNOR2_X1 U6907 ( .A(n5372), .B(n5370), .ZN(n6752) );
  NAND2_X1 U6908 ( .A1(n6752), .A2(n5443), .ZN(n5360) );
  OR2_X1 U6909 ( .A1(n5377), .A2(n5198), .ZN(n5358) );
  XNOR2_X1 U6910 ( .A(n5358), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7363) );
  AOI22_X1 U6911 ( .A1(n5483), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5482), .B2(
        n7363), .ZN(n5359) );
  NAND2_X1 U6912 ( .A1(n5135), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5369) );
  INV_X1 U6913 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n5361) );
  OR2_X1 U6914 ( .A1(n5545), .A2(n5361), .ZN(n5368) );
  INV_X1 U6915 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6916 ( .A1(n5363), .A2(n5362), .ZN(n5364) );
  NAND2_X1 U6917 ( .A1(n5384), .A2(n5364), .ZN(n7667) );
  OR2_X1 U6918 ( .A1(n5671), .A2(n7667), .ZN(n5367) );
  INV_X1 U6919 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n5365) );
  OR2_X1 U6920 ( .A1(n5471), .A2(n5365), .ZN(n5366) );
  OR2_X1 U6921 ( .A1(n7668), .A2(n9953), .ZN(n9261) );
  NAND2_X1 U6922 ( .A1(n7668), .A2(n9953), .ZN(n9257) );
  NAND2_X1 U6923 ( .A1(n9261), .A2(n9257), .ZN(n9091) );
  NAND2_X1 U6924 ( .A1(n5372), .A2(n5371), .ZN(n5375) );
  NAND2_X1 U6925 ( .A1(n5373), .A2(SI_13_), .ZN(n5374) );
  NAND2_X1 U6926 ( .A1(n5375), .A2(n5374), .ZN(n5396) );
  MUX2_X1 U6927 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4436), .Z(n5397) );
  XNOR2_X1 U6928 ( .A(n5396), .B(n5394), .ZN(n6830) );
  NAND2_X1 U6929 ( .A1(n6830), .A2(n5443), .ZN(n5383) );
  NAND2_X1 U6930 ( .A1(n5377), .A2(n5376), .ZN(n5378) );
  NAND2_X1 U6931 ( .A1(n5378), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U6932 ( .A1(n5380), .A2(n5379), .ZN(n5401) );
  OR2_X1 U6933 ( .A1(n5380), .A2(n5379), .ZN(n5381) );
  AOI22_X1 U6934 ( .A1(n5483), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5482), .B2(
        n7607), .ZN(n5382) );
  NAND2_X1 U6935 ( .A1(n5135), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5390) );
  INV_X1 U6936 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7719) );
  OR2_X1 U6937 ( .A1(n5545), .A2(n7719), .ZN(n5389) );
  INV_X1 U6938 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n10279) );
  INV_X1 U6939 ( .A(n5405), .ZN(n5407) );
  NAND2_X1 U6940 ( .A1(n5384), .A2(n10279), .ZN(n5385) );
  NAND2_X1 U6941 ( .A1(n5407), .A2(n5385), .ZN(n8911) );
  OR2_X1 U6942 ( .A1(n5671), .A2(n8911), .ZN(n5388) );
  INV_X1 U6943 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n5386) );
  OR2_X1 U6944 ( .A1(n6670), .A2(n5386), .ZN(n5387) );
  INV_X1 U6945 ( .A(n7829), .ZN(n9314) );
  OR2_X1 U6946 ( .A1(n9956), .A2(n9314), .ZN(n5391) );
  INV_X1 U6947 ( .A(n9953), .ZN(n9315) );
  OR2_X1 U6948 ( .A1(n7668), .A2(n9315), .ZN(n7715) );
  NAND2_X1 U6949 ( .A1(n9956), .A2(n9314), .ZN(n5392) );
  NAND2_X1 U6950 ( .A1(n5393), .A2(n5392), .ZN(n7731) );
  INV_X1 U6951 ( .A(n7731), .ZN(n5414) );
  NAND2_X1 U6952 ( .A1(n5396), .A2(n5395), .ZN(n5399) );
  NAND2_X1 U6953 ( .A1(n5397), .A2(SI_14_), .ZN(n5398) );
  MUX2_X1 U6954 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4436), .Z(n5418) );
  XNOR2_X1 U6955 ( .A(n5418), .B(SI_15_), .ZN(n5400) );
  XNOR2_X1 U6956 ( .A(n5417), .B(n5400), .ZN(n6902) );
  NAND2_X1 U6957 ( .A1(n6902), .A2(n5443), .ZN(n5404) );
  NAND2_X1 U6958 ( .A1(n5401), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5402) );
  XNOR2_X1 U6959 ( .A(n5402), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9381) );
  AOI22_X1 U6960 ( .A1(n5483), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9381), .B2(
        n5482), .ZN(n5403) );
  NAND2_X1 U6961 ( .A1(n5135), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5413) );
  INV_X1 U6962 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7739) );
  OR2_X1 U6963 ( .A1(n5545), .A2(n7739), .ZN(n5412) );
  INV_X1 U6964 ( .A(n5430), .ZN(n5432) );
  INV_X1 U6965 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U6966 ( .A1(n5407), .A2(n5406), .ZN(n5408) );
  NAND2_X1 U6967 ( .A1(n5432), .A2(n5408), .ZN(n9047) );
  OR2_X1 U6968 ( .A1(n5671), .A2(n9047), .ZN(n5411) );
  INV_X1 U6969 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5409) );
  OR2_X1 U6970 ( .A1(n5471), .A2(n5409), .ZN(n5410) );
  NAND2_X1 U6971 ( .A1(n5414), .A2(n4457), .ZN(n5416) );
  OR2_X1 U6972 ( .A1(n9151), .A2(n9780), .ZN(n5415) );
  NAND2_X1 U6973 ( .A1(n5419), .A2(n10232), .ZN(n5420) );
  MUX2_X1 U6974 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n4436), .Z(n5421) );
  INV_X1 U6975 ( .A(n5421), .ZN(n5423) );
  INV_X1 U6976 ( .A(SI_16_), .ZN(n5422) );
  NAND2_X1 U6977 ( .A1(n5423), .A2(n5422), .ZN(n5424) );
  NAND2_X1 U6978 ( .A1(n5440), .A2(n5424), .ZN(n5441) );
  INV_X1 U6979 ( .A(n5441), .ZN(n5425) );
  XNOR2_X1 U6980 ( .A(n5442), .B(n5425), .ZN(n6944) );
  NAND2_X1 U6981 ( .A1(n6944), .A2(n5443), .ZN(n5429) );
  INV_X1 U6982 ( .A(n5444), .ZN(n5426) );
  NAND2_X1 U6983 ( .A1(n5426), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5427) );
  XNOR2_X1 U6984 ( .A(n5427), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9397) );
  AOI22_X1 U6985 ( .A1(n5483), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5482), .B2(
        n9397), .ZN(n5428) );
  NAND2_X1 U6986 ( .A1(n4437), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5438) );
  INV_X1 U6987 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6988 ( .A1(n5432), .A2(n5431), .ZN(n5433) );
  NAND2_X1 U6989 ( .A1(n5449), .A2(n5433), .ZN(n8974) );
  OR2_X1 U6990 ( .A1(n5671), .A2(n8974), .ZN(n5437) );
  INV_X1 U6991 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7805) );
  OR2_X1 U6992 ( .A1(n5545), .A2(n7805), .ZN(n5436) );
  INV_X1 U6993 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9378) );
  OR2_X1 U6994 ( .A1(n6670), .A2(n9378), .ZN(n5435) );
  NAND2_X1 U6995 ( .A1(n7813), .A2(n9622), .ZN(n9273) );
  INV_X1 U6996 ( .A(n9622), .ZN(n7742) );
  NAND2_X1 U6997 ( .A1(n7813), .A2(n7742), .ZN(n5439) );
  MUX2_X1 U6998 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n4436), .Z(n5458) );
  XNOR2_X1 U6999 ( .A(n5460), .B(n5459), .ZN(n7052) );
  NAND2_X1 U7000 ( .A1(n7052), .A2(n5443), .ZN(n5447) );
  INV_X1 U7001 ( .A(n5682), .ZN(n5445) );
  XNOR2_X1 U7002 ( .A(n5465), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9423) );
  AOI22_X1 U7003 ( .A1(n5483), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5482), .B2(
        n9423), .ZN(n5446) );
  INV_X1 U7004 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10267) );
  OR2_X1 U7005 ( .A1(n5585), .A2(n10267), .ZN(n5455) );
  INV_X1 U7006 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U7007 ( .A1(n5449), .A2(n5448), .ZN(n5450) );
  NAND2_X1 U7008 ( .A1(n5469), .A2(n5450), .ZN(n9615) );
  OR2_X1 U7009 ( .A1(n9615), .A2(n5671), .ZN(n5454) );
  INV_X1 U7010 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9408) );
  OR2_X1 U7011 ( .A1(n5545), .A2(n9408), .ZN(n5453) );
  INV_X1 U7012 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n5451) );
  OR2_X1 U7013 ( .A1(n6670), .A2(n5451), .ZN(n5452) );
  NAND2_X1 U7014 ( .A1(n9709), .A2(n9781), .ZN(n5456) );
  NAND2_X1 U7015 ( .A1(n5457), .A2(n5456), .ZN(n9595) );
  MUX2_X1 U7016 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4436), .Z(n5461) );
  NAND2_X1 U7017 ( .A1(n5461), .A2(SI_18_), .ZN(n5478) );
  OAI21_X1 U7018 ( .B1(n5461), .B2(SI_18_), .A(n5478), .ZN(n5462) );
  NAND2_X1 U7019 ( .A1(n5463), .A2(n5462), .ZN(n5464) );
  AND2_X1 U7020 ( .A1(n5464), .A2(n5479), .ZN(n7143) );
  NAND2_X1 U7021 ( .A1(n7143), .A2(n5443), .ZN(n5467) );
  INV_X1 U7022 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5679) );
  XNOR2_X1 U7023 ( .A(n5480), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9441) );
  AOI22_X1 U7024 ( .A1(n5483), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5482), .B2(
        n9441), .ZN(n5466) );
  INV_X1 U7025 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5468) );
  INV_X1 U7026 ( .A(n5486), .ZN(n5488) );
  NAND2_X1 U7027 ( .A1(n5469), .A2(n5468), .ZN(n5470) );
  NAND2_X1 U7028 ( .A1(n5488), .A2(n5470), .ZN(n9596) );
  OR2_X1 U7029 ( .A1(n9596), .A2(n5434), .ZN(n5476) );
  INV_X1 U7030 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9705) );
  OR2_X1 U7031 ( .A1(n5471), .A2(n9705), .ZN(n5473) );
  INV_X1 U7032 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10254) );
  OR2_X1 U7033 ( .A1(n5585), .A2(n10254), .ZN(n5472) );
  AND2_X1 U7034 ( .A1(n5473), .A2(n5472), .ZN(n5475) );
  NAND2_X1 U7035 ( .A1(n6667), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5474) );
  INV_X1 U7036 ( .A(n9690), .ZN(n9313) );
  AND2_X1 U7037 ( .A1(n9609), .A2(n9313), .ZN(n5477) );
  MUX2_X1 U7038 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n4436), .Z(n5494) );
  XNOR2_X1 U7039 ( .A(n5496), .B(n5495), .ZN(n7268) );
  NAND2_X1 U7040 ( .A1(n7268), .A2(n5443), .ZN(n5485) );
  AOI22_X1 U7041 ( .A1(n5483), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n5685), .B2(
        n5482), .ZN(n5484) );
  INV_X1 U7042 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9581) );
  NAND2_X1 U7043 ( .A1(n5486), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5499) );
  INV_X1 U7044 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U7045 ( .A1(n5488), .A2(n5487), .ZN(n5489) );
  NAND2_X1 U7046 ( .A1(n5499), .A2(n5489), .ZN(n9580) );
  OR2_X1 U7047 ( .A1(n9580), .A2(n5671), .ZN(n5491) );
  AOI22_X1 U7048 ( .A1(n5582), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n5135), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5490) );
  OAI211_X1 U7049 ( .C1(n5545), .C2(n9581), .A(n5491), .B(n5490), .ZN(n9699)
         );
  NOR2_X1 U7050 ( .A1(n9588), .A2(n9699), .ZN(n9118) );
  OR2_X1 U7051 ( .A1(n9579), .A2(n9118), .ZN(n5493) );
  NAND2_X1 U7052 ( .A1(n9588), .A2(n9699), .ZN(n5492) );
  NAND2_X1 U7053 ( .A1(n5493), .A2(n5492), .ZN(n7892) );
  INV_X1 U7054 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6314) );
  INV_X1 U7055 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7322) );
  MUX2_X1 U7056 ( .A(n6314), .B(n7322), .S(n4436), .Z(n5510) );
  XNOR2_X1 U7057 ( .A(n5510), .B(SI_20_), .ZN(n5507) );
  XNOR2_X1 U7058 ( .A(n5508), .B(n5507), .ZN(n7321) );
  NAND2_X1 U7059 ( .A1(n7321), .A2(n5443), .ZN(n5498) );
  OR2_X1 U7060 ( .A1(n9075), .A2(n7322), .ZN(n5497) );
  INV_X1 U7061 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9003) );
  NAND2_X1 U7062 ( .A1(n5499), .A2(n9003), .ZN(n5500) );
  NAND2_X1 U7063 ( .A1(n5517), .A2(n5500), .ZN(n9002) );
  OR2_X1 U7064 ( .A1(n9002), .A2(n5434), .ZN(n5505) );
  INV_X1 U7065 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9688) );
  NAND2_X1 U7066 ( .A1(n4437), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U7067 ( .A1(n6667), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5501) );
  OAI211_X1 U7068 ( .C1(n9688), .C2(n6670), .A(n5502), .B(n5501), .ZN(n5503)
         );
  INV_X1 U7069 ( .A(n5503), .ZN(n5504) );
  AND2_X1 U7070 ( .A1(n7895), .A2(n9583), .ZN(n5506) );
  NAND2_X1 U7071 ( .A1(n5508), .A2(n5507), .ZN(n5512) );
  INV_X1 U7072 ( .A(SI_20_), .ZN(n5509) );
  NAND2_X1 U7073 ( .A1(n5510), .A2(n5509), .ZN(n5511) );
  INV_X1 U7074 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7361) );
  INV_X1 U7075 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7358) );
  MUX2_X1 U7076 ( .A(n7361), .B(n7358), .S(n4436), .Z(n5527) );
  XNOR2_X1 U7077 ( .A(n5527), .B(SI_21_), .ZN(n5513) );
  XNOR2_X1 U7078 ( .A(n5531), .B(n5513), .ZN(n7357) );
  NAND2_X1 U7079 ( .A1(n7357), .A2(n5443), .ZN(n5515) );
  OR2_X1 U7080 ( .A1(n9075), .A2(n7358), .ZN(n5514) );
  NAND2_X2 U7081 ( .A1(n5515), .A2(n5514), .ZN(n9676) );
  INV_X1 U7082 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U7083 ( .A1(n5517), .A2(n5516), .ZN(n5518) );
  AND2_X1 U7084 ( .A1(n5541), .A2(n5518), .ZN(n8941) );
  NAND2_X1 U7085 ( .A1(n8941), .A2(n5137), .ZN(n5524) );
  INV_X1 U7086 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U7087 ( .A1(n4437), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7088 ( .A1(n6667), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5519) );
  OAI211_X1 U7089 ( .C1(n5521), .C2(n6670), .A(n5520), .B(n5519), .ZN(n5522)
         );
  INV_X1 U7090 ( .A(n5522), .ZN(n5523) );
  NOR2_X1 U7091 ( .A1(n9676), .A2(n9312), .ZN(n5525) );
  NAND2_X1 U7092 ( .A1(n9676), .A2(n9312), .ZN(n5526) );
  NAND2_X1 U7093 ( .A1(n5528), .A2(SI_21_), .ZN(n5529) );
  INV_X1 U7094 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n10269) );
  INV_X1 U7095 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7452) );
  MUX2_X1 U7096 ( .A(n10269), .B(n7452), .S(n4436), .Z(n5533) );
  INV_X1 U7097 ( .A(SI_22_), .ZN(n5532) );
  NAND2_X1 U7098 ( .A1(n5533), .A2(n5532), .ZN(n5551) );
  INV_X1 U7099 ( .A(n5533), .ZN(n5534) );
  NAND2_X1 U7100 ( .A1(n5534), .A2(SI_22_), .ZN(n5535) );
  NAND2_X1 U7101 ( .A1(n5551), .A2(n5535), .ZN(n5536) );
  NAND2_X1 U7102 ( .A1(n5537), .A2(n5536), .ZN(n5538) );
  NAND2_X1 U7103 ( .A1(n5552), .A2(n5538), .ZN(n7451) );
  NAND2_X1 U7104 ( .A1(n7451), .A2(n5443), .ZN(n5540) );
  OR2_X1 U7105 ( .A1(n9075), .A2(n7452), .ZN(n5539) );
  INV_X1 U7106 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9012) );
  INV_X1 U7107 ( .A(n5564), .ZN(n5565) );
  NAND2_X1 U7108 ( .A1(n5541), .A2(n9012), .ZN(n5542) );
  NAND2_X1 U7109 ( .A1(n5565), .A2(n5542), .ZN(n9564) );
  OR2_X1 U7110 ( .A1(n9564), .A2(n5434), .ZN(n5548) );
  INV_X1 U7111 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9563) );
  NAND2_X1 U7112 ( .A1(n5135), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7113 ( .A1(n5582), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5543) );
  OAI211_X1 U7114 ( .C1(n9563), .C2(n5545), .A(n5544), .B(n5543), .ZN(n5546)
         );
  INV_X1 U7115 ( .A(n5546), .ZN(n5547) );
  OR2_X1 U7116 ( .A1(n9740), .A2(n9555), .ZN(n5549) );
  INV_X1 U7117 ( .A(n5560), .ZN(n5557) );
  INV_X1 U7118 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7648) );
  INV_X1 U7119 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7644) );
  MUX2_X1 U7120 ( .A(n7648), .B(n7644), .S(n4436), .Z(n5554) );
  INV_X1 U7121 ( .A(SI_23_), .ZN(n5553) );
  NAND2_X1 U7122 ( .A1(n5554), .A2(n5553), .ZN(n5591) );
  INV_X1 U7123 ( .A(n5554), .ZN(n5555) );
  NAND2_X1 U7124 ( .A1(n5555), .A2(SI_23_), .ZN(n5556) );
  NAND2_X1 U7125 ( .A1(n5591), .A2(n5556), .ZN(n5558) );
  NAND2_X1 U7126 ( .A1(n5557), .A2(n5558), .ZN(n5561) );
  INV_X1 U7127 ( .A(n5558), .ZN(n5559) );
  NAND2_X1 U7128 ( .A1(n5561), .A2(n5593), .ZN(n7645) );
  NAND2_X1 U7129 ( .A1(n7645), .A2(n5443), .ZN(n5563) );
  OR2_X1 U7130 ( .A1(n9075), .A2(n7644), .ZN(n5562) );
  NAND2_X1 U7131 ( .A1(n5564), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5580) );
  INV_X1 U7132 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8923) );
  NAND2_X1 U7133 ( .A1(n5565), .A2(n8923), .ZN(n5566) );
  NAND2_X1 U7134 ( .A1(n5580), .A2(n5566), .ZN(n9546) );
  OR2_X1 U7135 ( .A1(n9546), .A2(n5434), .ZN(n5571) );
  INV_X1 U7136 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10159) );
  NAND2_X1 U7137 ( .A1(n6667), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U7138 ( .A1(n4437), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5567) );
  OAI211_X1 U7139 ( .C1(n6670), .C2(n10159), .A(n5568), .B(n5567), .ZN(n5569)
         );
  INV_X1 U7140 ( .A(n5569), .ZN(n5570) );
  INV_X1 U7141 ( .A(n9659), .ZN(n9311) );
  INV_X1 U7142 ( .A(n9665), .ZN(n9549) );
  NAND2_X1 U7143 ( .A1(n5593), .A2(n5591), .ZN(n5576) );
  INV_X1 U7144 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n10301) );
  INV_X1 U7145 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10162) );
  MUX2_X1 U7146 ( .A(n10301), .B(n10162), .S(n4436), .Z(n5573) );
  INV_X1 U7147 ( .A(SI_24_), .ZN(n5572) );
  NAND2_X1 U7148 ( .A1(n5573), .A2(n5572), .ZN(n5590) );
  INV_X1 U7149 ( .A(n5573), .ZN(n5574) );
  NAND2_X1 U7150 ( .A1(n5574), .A2(SI_24_), .ZN(n5594) );
  AND2_X1 U7151 ( .A1(n5590), .A2(n5594), .ZN(n5575) );
  NAND2_X1 U7152 ( .A1(n7703), .A2(n5443), .ZN(n5578) );
  OR2_X1 U7153 ( .A1(n9075), .A2(n10162), .ZN(n5577) );
  INV_X1 U7154 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U7155 ( .A1(n5580), .A2(n5579), .ZN(n5581) );
  AND2_X1 U7156 ( .A1(n5601), .A2(n5581), .ZN(n9534) );
  NAND2_X1 U7157 ( .A1(n9534), .A2(n5137), .ZN(n5588) );
  INV_X1 U7158 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9734) );
  NAND2_X1 U7159 ( .A1(n6667), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U7160 ( .A1(n5582), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5583) );
  OAI211_X1 U7161 ( .C1(n5585), .C2(n9734), .A(n5584), .B(n5583), .ZN(n5586)
         );
  INV_X1 U7162 ( .A(n5586), .ZN(n5587) );
  AND2_X1 U7163 ( .A1(n9540), .A2(n9556), .ZN(n5589) );
  AND2_X1 U7164 ( .A1(n5591), .A2(n5590), .ZN(n5592) );
  INV_X1 U7165 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n10115) );
  INV_X1 U7166 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7729) );
  MUX2_X1 U7167 ( .A(n10115), .B(n7729), .S(n4436), .Z(n5596) );
  INV_X1 U7168 ( .A(SI_25_), .ZN(n5595) );
  NAND2_X1 U7169 ( .A1(n5596), .A2(n5595), .ZN(n5610) );
  INV_X1 U7170 ( .A(n5596), .ZN(n5597) );
  NAND2_X1 U7171 ( .A1(n5597), .A2(SI_25_), .ZN(n5598) );
  XNOR2_X1 U7172 ( .A(n5609), .B(n5608), .ZN(n7728) );
  NAND2_X1 U7173 ( .A1(n7728), .A2(n5443), .ZN(n5600) );
  OR2_X1 U7174 ( .A1(n9075), .A2(n7729), .ZN(n5599) );
  INV_X1 U7175 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8964) );
  INV_X1 U7176 ( .A(n5618), .ZN(n5620) );
  NAND2_X1 U7177 ( .A1(n5601), .A2(n8964), .ZN(n5602) );
  NAND2_X1 U7178 ( .A1(n5620), .A2(n5602), .ZN(n8963) );
  OR2_X1 U7179 ( .A1(n8963), .A2(n5434), .ZN(n5607) );
  INV_X1 U7180 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10237) );
  NAND2_X1 U7181 ( .A1(n5135), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U7182 ( .A1(n6667), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5603) );
  OAI211_X1 U7183 ( .C1(n6670), .C2(n10237), .A(n5604), .B(n5603), .ZN(n5605)
         );
  INV_X1 U7184 ( .A(n5605), .ZN(n5606) );
  INV_X1 U7185 ( .A(n9731), .ZN(n7879) );
  INV_X1 U7186 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7826) );
  INV_X1 U7187 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7801) );
  MUX2_X1 U7188 ( .A(n7826), .B(n7801), .S(n4436), .Z(n5613) );
  INV_X1 U7189 ( .A(SI_26_), .ZN(n5612) );
  NAND2_X1 U7190 ( .A1(n5613), .A2(n5612), .ZN(n5644) );
  INV_X1 U7191 ( .A(n5613), .ZN(n5614) );
  NAND2_X1 U7192 ( .A1(n5614), .A2(SI_26_), .ZN(n5615) );
  NAND2_X1 U7193 ( .A1(n7800), .A2(n5443), .ZN(n5617) );
  OR2_X1 U7194 ( .A1(n9075), .A2(n7801), .ZN(n5616) );
  INV_X1 U7195 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U7196 ( .A1(n5620), .A2(n5619), .ZN(n5621) );
  NAND2_X1 U7197 ( .A1(n9523), .A2(n5137), .ZN(n5626) );
  INV_X1 U7198 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10194) );
  NAND2_X1 U7199 ( .A1(n6667), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U7200 ( .A1(n4437), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5622) );
  OAI211_X1 U7201 ( .C1(n6670), .C2(n10194), .A(n5623), .B(n5622), .ZN(n5624)
         );
  INV_X1 U7202 ( .A(n5624), .ZN(n5625) );
  OR2_X1 U7203 ( .A1(n9522), .A2(n9649), .ZN(n9116) );
  NAND2_X1 U7204 ( .A1(n9522), .A2(n9649), .ZN(n9114) );
  OR2_X1 U7205 ( .A1(n9522), .A2(n9498), .ZN(n5627) );
  NAND2_X1 U7206 ( .A1(n5646), .A2(n5644), .ZN(n5634) );
  INV_X1 U7207 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7848) );
  INV_X1 U7208 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7842) );
  MUX2_X1 U7209 ( .A(n7848), .B(n7842), .S(n4436), .Z(n5631) );
  INV_X1 U7210 ( .A(SI_27_), .ZN(n5630) );
  NAND2_X1 U7211 ( .A1(n5631), .A2(n5630), .ZN(n5643) );
  INV_X1 U7212 ( .A(n5631), .ZN(n5632) );
  NAND2_X1 U7213 ( .A1(n5632), .A2(SI_27_), .ZN(n5647) );
  AND2_X1 U7214 ( .A1(n5643), .A2(n5647), .ZN(n5633) );
  NAND2_X1 U7215 ( .A1(n7841), .A2(n5443), .ZN(n5636) );
  OR2_X1 U7216 ( .A1(n9075), .A2(n7842), .ZN(n5635) );
  XNOR2_X1 U7217 ( .A(n5652), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9503) );
  NAND2_X1 U7218 ( .A1(n9503), .A2(n5137), .ZN(n5641) );
  INV_X1 U7219 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10286) );
  NAND2_X1 U7220 ( .A1(n4437), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U7221 ( .A1(n6667), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5637) );
  OAI211_X1 U7222 ( .C1(n6670), .C2(n10286), .A(n5638), .B(n5637), .ZN(n5639)
         );
  INV_X1 U7223 ( .A(n5639), .ZN(n5640) );
  INV_X1 U7224 ( .A(n9515), .ZN(n6021) );
  NAND2_X1 U7225 ( .A1(n4847), .A2(n6021), .ZN(n9213) );
  INV_X1 U7226 ( .A(n9496), .ZN(n9508) );
  NAND2_X1 U7227 ( .A1(n9505), .A2(n6021), .ZN(n5642) );
  AND2_X1 U7228 ( .A1(n5644), .A2(n5643), .ZN(n5645) );
  NAND2_X1 U7229 ( .A1(n5646), .A2(n5645), .ZN(n5648) );
  MUX2_X1 U7230 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n4436), .Z(n5664) );
  INV_X1 U7231 ( .A(SI_28_), .ZN(n5665) );
  XNOR2_X1 U7232 ( .A(n5664), .B(n5665), .ZN(n5662) );
  NAND2_X1 U7233 ( .A1(n7849), .A2(n5443), .ZN(n5650) );
  INV_X1 U7234 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7850) );
  OR2_X1 U7235 ( .A1(n9075), .A2(n7850), .ZN(n5649) );
  NAND2_X2 U7236 ( .A1(n5650), .A2(n5649), .ZN(n9488) );
  INV_X1 U7237 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7952) );
  INV_X1 U7238 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5651) );
  OAI21_X1 U7239 ( .B1(n5652), .B2(n7952), .A(n5651), .ZN(n5655) );
  AND2_X1 U7240 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5653) );
  NAND2_X1 U7241 ( .A1(n5654), .A2(n5653), .ZN(n9471) );
  NAND2_X1 U7242 ( .A1(n5655), .A2(n9471), .ZN(n6005) );
  OR2_X1 U7243 ( .A1(n6005), .A2(n5434), .ZN(n5660) );
  INV_X1 U7244 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n10143) );
  NAND2_X1 U7245 ( .A1(n5135), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U7246 ( .A1(n6667), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5656) );
  OAI211_X1 U7247 ( .C1(n6670), .C2(n10143), .A(n5657), .B(n5656), .ZN(n5658)
         );
  INV_X1 U7248 ( .A(n5658), .ZN(n5659) );
  NAND2_X1 U7249 ( .A1(n9488), .A2(n9497), .ZN(n5661) );
  INV_X1 U7250 ( .A(n5664), .ZN(n5666) );
  NAND2_X1 U7251 ( .A1(n5666), .A2(n5665), .ZN(n5667) );
  INV_X1 U7252 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7965) );
  INV_X1 U7253 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7867) );
  MUX2_X1 U7254 ( .A(n7965), .B(n7867), .S(n4436), .Z(n8117) );
  NAND2_X1 U7255 ( .A1(n7866), .A2(n5443), .ZN(n5670) );
  OR2_X1 U7256 ( .A1(n9075), .A2(n7867), .ZN(n5669) );
  NAND2_X2 U7257 ( .A1(n5670), .A2(n5669), .ZN(n9473) );
  OR2_X1 U7258 ( .A1(n9471), .A2(n5434), .ZN(n5676) );
  INV_X1 U7259 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n10173) );
  NAND2_X1 U7260 ( .A1(n4437), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U7261 ( .A1(n6667), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5672) );
  OAI211_X1 U7262 ( .C1(n6670), .C2(n10173), .A(n5673), .B(n5672), .ZN(n5674)
         );
  INV_X1 U7263 ( .A(n5674), .ZN(n5675) );
  AND2_X1 U7264 ( .A1(n5676), .A2(n5675), .ZN(n6017) );
  OR2_X1 U7265 ( .A1(n9473), .A2(n6017), .ZN(n9214) );
  NAND2_X1 U7266 ( .A1(n9473), .A2(n6017), .ZN(n9215) );
  XNOR2_X1 U7267 ( .A(n5677), .B(n9105), .ZN(n9469) );
  INV_X1 U7268 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5678) );
  AND3_X1 U7269 ( .A1(n5680), .A2(n5679), .A3(n5678), .ZN(n5681) );
  NAND2_X1 U7270 ( .A1(n5687), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5688) );
  MUX2_X1 U7271 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5688), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5690) );
  OR2_X1 U7272 ( .A1(n5765), .A2(n7156), .ZN(n9303) );
  INV_X1 U7273 ( .A(n9225), .ZN(n9236) );
  NAND2_X1 U7274 ( .A1(n5691), .A2(n9236), .ZN(n6803) );
  NAND2_X1 U7275 ( .A1(n5765), .A2(n5763), .ZN(n5692) );
  NAND3_X1 U7276 ( .A1(n9303), .A2(n6803), .A3(n5692), .ZN(n9814) );
  NAND2_X1 U7277 ( .A1(n9469), .A2(n9949), .ZN(n5724) );
  INV_X1 U7278 ( .A(n9740), .ZN(n9567) );
  NAND2_X1 U7279 ( .A1(n9237), .A2(n7141), .ZN(n7302) );
  NAND2_X1 U7280 ( .A1(n9836), .A2(n7316), .ZN(n7311) );
  INV_X1 U7281 ( .A(n9899), .ZN(n7265) );
  INV_X1 U7282 ( .A(n7387), .ZN(n9911) );
  NOR2_X2 U7283 ( .A1(n4467), .A2(n9930), .ZN(n9804) );
  INV_X1 U7284 ( .A(n9802), .ZN(n9937) );
  INV_X1 U7285 ( .A(n7527), .ZN(n8959) );
  NAND2_X1 U7286 ( .A1(n7504), .A2(n8959), .ZN(n7505) );
  OR2_X2 U7287 ( .A1(n7505), .A2(n7668), .ZN(n7718) );
  INV_X1 U7288 ( .A(n9151), .ZN(n7840) );
  NOR2_X2 U7289 ( .A1(n4469), .A2(n9609), .ZN(n9604) );
  OR2_X2 U7290 ( .A1(n9536), .A2(n9540), .ZN(n9537) );
  OR2_X2 U7291 ( .A1(n9537), .A2(n9731), .ZN(n9521) );
  AOI21_X1 U7292 ( .B1(n9473), .B2(n4848), .A(n9822), .ZN(n5694) );
  NAND2_X1 U7293 ( .A1(n5694), .A2(n9462), .ZN(n9475) );
  OR2_X1 U7294 ( .A1(n5762), .A2(n9237), .ZN(n5695) );
  NAND2_X1 U7295 ( .A1(n5698), .A2(n5697), .ZN(n9827) );
  INV_X1 U7296 ( .A(n9083), .ZN(n7160) );
  NAND2_X1 U7297 ( .A1(n9242), .A2(n7160), .ZN(n5700) );
  INV_X1 U7298 ( .A(n9133), .ZN(n9248) );
  NAND2_X1 U7299 ( .A1(n9156), .A2(n9136), .ZN(n9144) );
  NAND2_X1 U7300 ( .A1(n9143), .A2(n7379), .ZN(n9140) );
  INV_X1 U7301 ( .A(n9140), .ZN(n7324) );
  NAND2_X1 U7302 ( .A1(n9135), .A2(n9126), .ZN(n5701) );
  NAND2_X1 U7303 ( .A1(n9802), .A2(n9926), .ZN(n9161) );
  NAND2_X1 U7304 ( .A1(n9161), .A2(n9794), .ZN(n9254) );
  INV_X1 U7305 ( .A(n9254), .ZN(n5702) );
  NAND2_X1 U7306 ( .A1(n7335), .A2(n5702), .ZN(n5703) );
  OR2_X1 U7307 ( .A1(n9802), .A2(n9926), .ZN(n9159) );
  NAND2_X1 U7308 ( .A1(n9956), .A2(n7829), .ZN(n9264) );
  OR2_X1 U7309 ( .A1(n9151), .A2(n9951), .ZN(n9267) );
  AND2_X1 U7310 ( .A1(n9151), .A2(n9951), .ZN(n9153) );
  INV_X1 U7311 ( .A(n9262), .ZN(n7733) );
  NOR2_X1 U7312 ( .A1(n7732), .A2(n7733), .ZN(n5704) );
  NAND2_X1 U7313 ( .A1(n7723), .A2(n5704), .ZN(n7735) );
  OR2_X1 U7314 ( .A1(n9709), .A2(n9603), .ZN(n9185) );
  NAND2_X1 U7315 ( .A1(n9709), .A2(n9603), .ZN(n9176) );
  OR2_X1 U7316 ( .A1(n9609), .A2(n9690), .ZN(n9186) );
  NAND2_X1 U7317 ( .A1(n9609), .A2(n9690), .ZN(n9188) );
  NAND2_X1 U7318 ( .A1(n9186), .A2(n9188), .ZN(n9096) );
  INV_X1 U7319 ( .A(n9699), .ZN(n9680) );
  NOR2_X1 U7320 ( .A1(n9588), .A2(n9680), .ZN(n9120) );
  INV_X1 U7321 ( .A(n9120), .ZN(n9177) );
  NAND2_X1 U7322 ( .A1(n9588), .A2(n9680), .ZN(n9282) );
  NAND2_X1 U7323 ( .A1(n9177), .A2(n9282), .ZN(n9578) );
  INV_X1 U7324 ( .A(n9578), .ZN(n5706) );
  NAND2_X1 U7325 ( .A1(n9577), .A2(n5706), .ZN(n5707) );
  NAND2_X1 U7326 ( .A1(n5707), .A2(n9282), .ZN(n7901) );
  NAND2_X1 U7327 ( .A1(n7895), .A2(n9691), .ZN(n9123) );
  OR2_X1 U7328 ( .A1(n9676), .A2(n9681), .ZN(n9193) );
  INV_X1 U7329 ( .A(n9181), .ZN(n5709) );
  OR2_X1 U7330 ( .A1(n7895), .A2(n9691), .ZN(n9121) );
  AND2_X1 U7331 ( .A1(n9099), .A2(n9121), .ZN(n5708) );
  NAND2_X1 U7332 ( .A1(n5709), .A2(n9123), .ZN(n9190) );
  AND2_X1 U7333 ( .A1(n9190), .A2(n9193), .ZN(n9065) );
  XNOR2_X1 U7334 ( .A(n9740), .B(n9555), .ZN(n9571) );
  NAND2_X1 U7335 ( .A1(n9740), .A2(n9058), .ZN(n9552) );
  NAND2_X1 U7336 ( .A1(n9570), .A2(n9552), .ZN(n5710) );
  NOR2_X1 U7337 ( .A1(n9665), .A2(n9659), .ZN(n9183) );
  INV_X1 U7338 ( .A(n9183), .ZN(n9060) );
  NAND2_X1 U7339 ( .A1(n9665), .A2(n9659), .ZN(n9196) );
  NAND2_X1 U7340 ( .A1(n5710), .A2(n9550), .ZN(n9554) );
  NAND2_X1 U7341 ( .A1(n9540), .A2(n9648), .ZN(n9205) );
  INV_X1 U7342 ( .A(n9532), .ZN(n9100) );
  OR2_X1 U7343 ( .A1(n9731), .A2(n8994), .ZN(n9115) );
  INV_X1 U7344 ( .A(n9115), .ZN(n5711) );
  NAND2_X1 U7345 ( .A1(n9731), .A2(n8994), .ZN(n9113) );
  NAND2_X1 U7346 ( .A1(n9488), .A2(n7953), .ZN(n9110) );
  NAND2_X1 U7347 ( .A1(n9480), .A2(n9485), .ZN(n9479) );
  NAND2_X1 U7348 ( .A1(n9479), .A2(n9110), .ZN(n5712) );
  XNOR2_X1 U7349 ( .A(n5712), .B(n9111), .ZN(n5723) );
  OR2_X1 U7350 ( .A1(n5713), .A2(n5691), .ZN(n5715) );
  NAND2_X1 U7351 ( .A1(n9225), .A2(n9233), .ZN(n5714) );
  INV_X1 U7352 ( .A(n9076), .ZN(n5996) );
  INV_X1 U7353 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10179) );
  NAND2_X1 U7354 ( .A1(n6667), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U7355 ( .A1(n5135), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5718) );
  OAI211_X1 U7356 ( .C1(n6670), .C2(n10179), .A(n5719), .B(n5718), .ZN(n9310)
         );
  INV_X1 U7357 ( .A(n9310), .ZN(n5721) );
  NAND2_X1 U7358 ( .A1(n4443), .A2(n9076), .ZN(n9950) );
  INV_X1 U7359 ( .A(P1_B_REG_SCAN_IN), .ZN(n5738) );
  NOR2_X1 U7360 ( .A1(n7843), .A2(n5738), .ZN(n5720) );
  OR2_X1 U7361 ( .A1(n9950), .A2(n5720), .ZN(n9457) );
  OAI22_X1 U7362 ( .A1(n7953), .A2(n9952), .B1(n5721), .B2(n9457), .ZN(n5722)
         );
  NAND2_X1 U7363 ( .A1(n4484), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U7364 ( .A1(n5728), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U7365 ( .A1(n5729), .A2(n5080), .ZN(n5731) );
  NAND2_X1 U7366 ( .A1(n5731), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5732) );
  INV_X1 U7367 ( .A(n5734), .ZN(n5735) );
  NAND2_X1 U7368 ( .A1(n5735), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5737) );
  XNOR2_X1 U7369 ( .A(n5737), .B(n5736), .ZN(n6585) );
  OR2_X1 U7370 ( .A1(n5754), .A2(n5738), .ZN(n5739) );
  MUX2_X1 U7371 ( .A(P1_B_REG_SCAN_IN), .B(n5739), .S(n7704), .Z(n5741) );
  INV_X1 U7372 ( .A(n7802), .ZN(n5740) );
  NOR2_X1 U7373 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .ZN(
        n5745) );
  NOR4_X1 U7374 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n5744) );
  NOR4_X1 U7375 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5743) );
  NOR4_X1 U7376 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5742) );
  NAND4_X1 U7377 ( .A1(n5745), .A2(n5744), .A3(n5743), .A4(n5742), .ZN(n5751)
         );
  NOR4_X1 U7378 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n5749) );
  NOR4_X1 U7379 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5748) );
  NOR4_X1 U7380 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5747) );
  NOR4_X1 U7381 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5746) );
  NAND4_X1 U7382 ( .A1(n5749), .A2(n5748), .A3(n5747), .A4(n5746), .ZN(n5750)
         );
  NOR2_X1 U7383 ( .A1(n5751), .A2(n5750), .ZN(n5992) );
  NAND2_X1 U7384 ( .A1(n6004), .A2(n5992), .ZN(n5752) );
  NAND2_X1 U7385 ( .A1(n9859), .A2(n5752), .ZN(n5753) );
  NAND2_X1 U7386 ( .A1(n9076), .A2(n5763), .ZN(n6008) );
  NAND2_X1 U7387 ( .A1(n5753), .A2(n6008), .ZN(n7130) );
  INV_X1 U7388 ( .A(n5754), .ZN(n7730) );
  NAND2_X1 U7389 ( .A1(n7730), .A2(n7802), .ZN(n9757) );
  OAI21_X1 U7390 ( .B1(n5993), .B2(P1_D_REG_1__SCAN_IN), .A(n9757), .ZN(n7128)
         );
  NAND2_X1 U7391 ( .A1(n7128), .A2(n6002), .ZN(n5758) );
  NAND2_X1 U7392 ( .A1(n7802), .A2(n7704), .ZN(n9758) );
  OAI21_X1 U7393 ( .B1(n5993), .B2(P1_D_REG_0__SCAN_IN), .A(n9758), .ZN(n5995)
         );
  INV_X1 U7394 ( .A(n5995), .ZN(n7129) );
  INV_X1 U7395 ( .A(n6803), .ZN(n7135) );
  NAND2_X1 U7396 ( .A1(n7135), .A2(n5763), .ZN(n9944) );
  NOR2_X1 U7397 ( .A1(n9965), .A2(n9944), .ZN(n9741) );
  OAI21_X1 U7398 ( .B1(n5757), .B2(n9981), .A(n5064), .ZN(n5760) );
  NOR2_X1 U7399 ( .A1(n9981), .A2(n9944), .ZN(n9673) );
  NAND2_X1 U7400 ( .A1(n9473), .A2(n9673), .ZN(n5759) );
  NAND2_X1 U7401 ( .A1(n5760), .A2(n5759), .ZN(P1_U3551) );
  INV_X2 U7402 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7403 ( .A(n7156), .ZN(n5761) );
  NAND2_X1 U7404 ( .A1(n5763), .A2(n7156), .ZN(n5764) );
  AOI21_X1 U7405 ( .B1(n9323), .B2(n5981), .A(n5767), .ZN(n5778) );
  XNOR2_X1 U7406 ( .A(n5777), .B(n5778), .ZN(n6542) );
  NAND2_X1 U7407 ( .A1(n9325), .A2(n5984), .ZN(n5770) );
  NAND2_X1 U7408 ( .A1(n9325), .A2(n5981), .ZN(n5774) );
  OAI22_X1 U7409 ( .A1(n7141), .A2(n5966), .B1(n6539), .B2(n9333), .ZN(n5772)
         );
  INV_X1 U7410 ( .A(n5772), .ZN(n5773) );
  NAND2_X1 U7411 ( .A1(n5774), .A2(n5773), .ZN(n6691) );
  NAND2_X1 U7412 ( .A1(n6692), .A2(n6691), .ZN(n6690) );
  NAND2_X1 U7413 ( .A1(n5775), .A2(n5987), .ZN(n5776) );
  NAND2_X1 U7414 ( .A1(n6542), .A2(n6541), .ZN(n6540) );
  INV_X1 U7415 ( .A(n5777), .ZN(n5779) );
  NAND2_X1 U7416 ( .A1(n5779), .A2(n5778), .ZN(n5780) );
  NAND2_X1 U7417 ( .A1(n6540), .A2(n5780), .ZN(n6833) );
  NAND2_X1 U7418 ( .A1(n4429), .A2(n5984), .ZN(n5782) );
  OR2_X1 U7419 ( .A1(n7300), .A2(n5795), .ZN(n5781) );
  NAND2_X1 U7420 ( .A1(n5782), .A2(n5781), .ZN(n5783) );
  XNOR2_X1 U7421 ( .A(n5783), .B(n5979), .ZN(n5784) );
  AOI22_X1 U7422 ( .A1(n4429), .A2(n5981), .B1(n9865), .B2(n5984), .ZN(n5785)
         );
  XNOR2_X1 U7423 ( .A(n5784), .B(n5785), .ZN(n6834) );
  INV_X1 U7424 ( .A(n5784), .ZN(n5786) );
  NAND2_X1 U7425 ( .A1(n5786), .A2(n5785), .ZN(n5787) );
  NAND2_X1 U7426 ( .A1(n9322), .A2(n5984), .ZN(n5789) );
  OR2_X1 U7427 ( .A1(n9872), .A2(n5795), .ZN(n5788) );
  NAND2_X1 U7428 ( .A1(n5789), .A2(n5788), .ZN(n5790) );
  XNOR2_X1 U7429 ( .A(n5790), .B(n5979), .ZN(n5791) );
  AOI22_X1 U7430 ( .A1(n9322), .A2(n5981), .B1(n9833), .B2(n5984), .ZN(n5792)
         );
  XNOR2_X1 U7431 ( .A(n5791), .B(n5792), .ZN(n6937) );
  INV_X1 U7432 ( .A(n5791), .ZN(n5793) );
  NAND2_X1 U7433 ( .A1(n5793), .A2(n5792), .ZN(n5794) );
  INV_X1 U7434 ( .A(n6991), .ZN(n5800) );
  NAND2_X1 U7435 ( .A1(n9829), .A2(n5984), .ZN(n5797) );
  OR2_X1 U7436 ( .A1(n7316), .A2(n5795), .ZN(n5796) );
  NAND2_X1 U7437 ( .A1(n5797), .A2(n5796), .ZN(n5798) );
  XNOR2_X1 U7438 ( .A(n5798), .B(n5987), .ZN(n5801) );
  AOI22_X1 U7439 ( .A1(n9829), .A2(n5981), .B1(n9881), .B2(n5984), .ZN(n5802)
         );
  XNOR2_X1 U7440 ( .A(n5801), .B(n5802), .ZN(n6990) );
  INV_X1 U7441 ( .A(n5801), .ZN(n5804) );
  NAND2_X1 U7442 ( .A1(n5804), .A2(n5803), .ZN(n5805) );
  NAND2_X1 U7443 ( .A1(n9321), .A2(n5984), .ZN(n5808) );
  OR2_X1 U7444 ( .A1(n5806), .A2(n5795), .ZN(n5807) );
  NAND2_X1 U7445 ( .A1(n5808), .A2(n5807), .ZN(n5809) );
  XNOR2_X1 U7446 ( .A(n5809), .B(n5979), .ZN(n5813) );
  INV_X1 U7447 ( .A(n5813), .ZN(n5810) );
  NAND2_X1 U7448 ( .A1(n9321), .A2(n5981), .ZN(n5812) );
  NAND2_X1 U7449 ( .A1(n9889), .A2(n5984), .ZN(n5811) );
  NAND2_X1 U7450 ( .A1(n5812), .A2(n5811), .ZN(n7150) );
  NAND2_X1 U7451 ( .A1(n7147), .A2(n7150), .ZN(n5815) );
  NAND2_X1 U7452 ( .A1(n5814), .A2(n5813), .ZN(n7148) );
  NAND2_X1 U7453 ( .A1(n5815), .A2(n7148), .ZN(n7258) );
  INV_X1 U7454 ( .A(n7258), .ZN(n5821) );
  NAND2_X1 U7455 ( .A1(n9890), .A2(n5984), .ZN(n5816) );
  OAI21_X1 U7456 ( .B1(n9899), .B2(n5795), .A(n5816), .ZN(n5817) );
  XNOR2_X1 U7457 ( .A(n5817), .B(n5979), .ZN(n5822) );
  OR2_X1 U7458 ( .A1(n9899), .A2(n5966), .ZN(n5819) );
  NAND2_X1 U7459 ( .A1(n9890), .A2(n5981), .ZN(n5818) );
  NAND2_X1 U7460 ( .A1(n5819), .A2(n5818), .ZN(n5823) );
  XNOR2_X1 U7461 ( .A(n5822), .B(n5823), .ZN(n7259) );
  INV_X1 U7462 ( .A(n7259), .ZN(n5820) );
  NAND2_X1 U7463 ( .A1(n5821), .A2(n5820), .ZN(n7256) );
  INV_X1 U7464 ( .A(n5822), .ZN(n5825) );
  INV_X1 U7465 ( .A(n5823), .ZN(n5824) );
  NAND2_X1 U7466 ( .A1(n5825), .A2(n5824), .ZN(n5826) );
  NAND2_X1 U7467 ( .A1(n9904), .A2(n5984), .ZN(n5829) );
  OR2_X1 U7468 ( .A1(n7623), .A2(n5827), .ZN(n5828) );
  NAND2_X1 U7469 ( .A1(n9904), .A2(n5978), .ZN(n5831) );
  OR2_X1 U7470 ( .A1(n7623), .A2(n5966), .ZN(n5830) );
  NAND2_X1 U7471 ( .A1(n5831), .A2(n5830), .ZN(n5832) );
  XNOR2_X1 U7472 ( .A(n5832), .B(n5979), .ZN(n7349) );
  NAND2_X1 U7473 ( .A1(n7387), .A2(n5978), .ZN(n5834) );
  OR2_X1 U7474 ( .A1(n9810), .A2(n5966), .ZN(n5833) );
  NAND2_X1 U7475 ( .A1(n5834), .A2(n5833), .ZN(n5835) );
  XNOR2_X1 U7476 ( .A(n5835), .B(n5987), .ZN(n5837) );
  AOI22_X1 U7477 ( .A1(n7387), .A2(n5984), .B1(n5981), .B2(n9917), .ZN(n7620)
         );
  INV_X1 U7478 ( .A(n5836), .ZN(n5838) );
  NAND2_X1 U7479 ( .A1(n5838), .A2(n5837), .ZN(n7691) );
  NAND2_X1 U7480 ( .A1(n9919), .A2(n5978), .ZN(n5840) );
  OR2_X1 U7481 ( .A1(n9927), .A2(n5966), .ZN(n5839) );
  NAND2_X1 U7482 ( .A1(n5840), .A2(n5839), .ZN(n5841) );
  XNOR2_X1 U7483 ( .A(n5841), .B(n5979), .ZN(n5843) );
  NOR2_X1 U7484 ( .A1(n9927), .A2(n5827), .ZN(n5842) );
  AOI21_X1 U7485 ( .B1(n9919), .B2(n5984), .A(n5842), .ZN(n5844) );
  XNOR2_X1 U7486 ( .A(n5843), .B(n5844), .ZN(n7693) );
  INV_X1 U7487 ( .A(n5843), .ZN(n5845) );
  OR2_X1 U7488 ( .A1(n5845), .A2(n5844), .ZN(n5846) );
  NAND2_X1 U7489 ( .A1(n9930), .A2(n5978), .ZN(n5848) );
  OR2_X1 U7490 ( .A1(n9792), .A2(n5966), .ZN(n5847) );
  NAND2_X1 U7491 ( .A1(n5848), .A2(n5847), .ZN(n5849) );
  XNOR2_X1 U7492 ( .A(n5849), .B(n5987), .ZN(n7853) );
  NOR2_X1 U7493 ( .A1(n9792), .A2(n5827), .ZN(n5850) );
  AOI21_X1 U7494 ( .B1(n9930), .B2(n5984), .A(n5850), .ZN(n7855) );
  NAND2_X1 U7495 ( .A1(n9802), .A2(n5978), .ZN(n5852) );
  OR2_X1 U7496 ( .A1(n9926), .A2(n5966), .ZN(n5851) );
  NAND2_X1 U7497 ( .A1(n5852), .A2(n5851), .ZN(n5853) );
  XNOR2_X1 U7498 ( .A(n5853), .B(n5979), .ZN(n5856) );
  NAND2_X1 U7499 ( .A1(n9802), .A2(n5984), .ZN(n5855) );
  OR2_X1 U7500 ( .A1(n9926), .A2(n5827), .ZN(n5854) );
  NAND2_X1 U7501 ( .A1(n5855), .A2(n5854), .ZN(n5857) );
  NAND2_X1 U7502 ( .A1(n5856), .A2(n5857), .ZN(n7857) );
  OAI21_X1 U7503 ( .B1(n7853), .B2(n7855), .A(n7857), .ZN(n5862) );
  NAND3_X1 U7504 ( .A1(n7857), .A2(n7853), .A3(n7855), .ZN(n5860) );
  INV_X1 U7505 ( .A(n5856), .ZN(n5859) );
  INV_X1 U7506 ( .A(n5857), .ZN(n5858) );
  NAND2_X1 U7507 ( .A1(n5859), .A2(n5858), .ZN(n8947) );
  AND2_X1 U7508 ( .A1(n5860), .A2(n8947), .ZN(n5861) );
  NAND2_X1 U7509 ( .A1(n7527), .A2(n5978), .ZN(n5864) );
  OR2_X1 U7510 ( .A1(n9793), .A2(n5966), .ZN(n5863) );
  NAND2_X1 U7511 ( .A1(n5864), .A2(n5863), .ZN(n5865) );
  XNOR2_X1 U7512 ( .A(n5865), .B(n5987), .ZN(n5868) );
  NOR2_X1 U7513 ( .A1(n9793), .A2(n5827), .ZN(n5866) );
  AOI21_X1 U7514 ( .B1(n7527), .B2(n5984), .A(n5866), .ZN(n5867) );
  NAND2_X1 U7515 ( .A1(n5868), .A2(n5867), .ZN(n7789) );
  OR2_X1 U7516 ( .A1(n5868), .A2(n5867), .ZN(n5869) );
  AND2_X1 U7517 ( .A1(n7789), .A2(n5869), .ZN(n8948) );
  NAND2_X1 U7518 ( .A1(n7668), .A2(n5978), .ZN(n5871) );
  OR2_X1 U7519 ( .A1(n9953), .A2(n5966), .ZN(n5870) );
  NAND2_X1 U7520 ( .A1(n5871), .A2(n5870), .ZN(n5872) );
  XNOR2_X1 U7521 ( .A(n5872), .B(n5987), .ZN(n5875) );
  NOR2_X1 U7522 ( .A1(n9953), .A2(n5827), .ZN(n5873) );
  AOI21_X1 U7523 ( .B1(n7668), .B2(n5984), .A(n5873), .ZN(n5874) );
  NAND2_X1 U7524 ( .A1(n5875), .A2(n5874), .ZN(n5878) );
  OR2_X1 U7525 ( .A1(n5875), .A2(n5874), .ZN(n5876) );
  AND2_X1 U7526 ( .A1(n5878), .A2(n5876), .ZN(n7790) );
  NAND2_X1 U7527 ( .A1(n5877), .A2(n7790), .ZN(n7791) );
  INV_X1 U7528 ( .A(n5795), .ZN(n5978) );
  NAND2_X1 U7529 ( .A1(n9956), .A2(n5978), .ZN(n5880) );
  OR2_X1 U7530 ( .A1(n7829), .A2(n5966), .ZN(n5879) );
  NAND2_X1 U7531 ( .A1(n5880), .A2(n5879), .ZN(n5881) );
  XNOR2_X1 U7532 ( .A(n5881), .B(n5987), .ZN(n5884) );
  NAND2_X1 U7533 ( .A1(n9956), .A2(n5984), .ZN(n5883) );
  OR2_X1 U7534 ( .A1(n7829), .A2(n5827), .ZN(n5882) );
  NAND2_X1 U7535 ( .A1(n5883), .A2(n5882), .ZN(n8907) );
  NAND2_X1 U7536 ( .A1(n9151), .A2(n5978), .ZN(n5887) );
  OR2_X1 U7537 ( .A1(n9951), .A2(n5966), .ZN(n5886) );
  NAND2_X1 U7538 ( .A1(n5887), .A2(n5886), .ZN(n5888) );
  XNOR2_X1 U7539 ( .A(n5888), .B(n5979), .ZN(n5889) );
  NAND2_X1 U7540 ( .A1(n5890), .A2(n5889), .ZN(n5891) );
  NAND2_X1 U7541 ( .A1(n9151), .A2(n5984), .ZN(n5893) );
  OR2_X1 U7542 ( .A1(n9951), .A2(n5827), .ZN(n5892) );
  NAND2_X1 U7543 ( .A1(n5893), .A2(n5892), .ZN(n9040) );
  INV_X1 U7544 ( .A(n9040), .ZN(n5894) );
  NAND2_X1 U7545 ( .A1(n7813), .A2(n5978), .ZN(n5897) );
  OR2_X1 U7546 ( .A1(n9622), .A2(n5966), .ZN(n5896) );
  NAND2_X1 U7547 ( .A1(n5897), .A2(n5896), .ZN(n5898) );
  XNOR2_X1 U7548 ( .A(n5898), .B(n5979), .ZN(n5904) );
  NOR2_X1 U7549 ( .A1(n9622), .A2(n5827), .ZN(n5899) );
  AOI21_X1 U7550 ( .B1(n7813), .B2(n5984), .A(n5899), .ZN(n5905) );
  XNOR2_X1 U7551 ( .A(n5904), .B(n5905), .ZN(n8972) );
  NAND2_X1 U7552 ( .A1(n9709), .A2(n5978), .ZN(n5901) );
  NAND2_X1 U7553 ( .A1(n9781), .A2(n5984), .ZN(n5900) );
  NAND2_X1 U7554 ( .A1(n5901), .A2(n5900), .ZN(n5902) );
  XNOR2_X1 U7555 ( .A(n5902), .B(n5979), .ZN(n5910) );
  NOR2_X1 U7556 ( .A1(n9603), .A2(n5827), .ZN(n5903) );
  AOI21_X1 U7557 ( .B1(n9709), .B2(n5984), .A(n5903), .ZN(n5908) );
  XNOR2_X1 U7558 ( .A(n5910), .B(n5908), .ZN(n8981) );
  INV_X1 U7559 ( .A(n5904), .ZN(n5906) );
  NAND2_X1 U7560 ( .A1(n5906), .A2(n5905), .ZN(n8979) );
  AND2_X1 U7561 ( .A1(n8981), .A2(n8979), .ZN(n5907) );
  INV_X1 U7562 ( .A(n5908), .ZN(n5909) );
  NAND2_X1 U7563 ( .A1(n9609), .A2(n5978), .ZN(n5912) );
  OR2_X1 U7564 ( .A1(n9690), .A2(n5966), .ZN(n5911) );
  NAND2_X1 U7565 ( .A1(n5912), .A2(n5911), .ZN(n5913) );
  XNOR2_X1 U7566 ( .A(n5913), .B(n5987), .ZN(n5915) );
  NOR2_X1 U7567 ( .A1(n9690), .A2(n5827), .ZN(n5914) );
  AOI21_X1 U7568 ( .B1(n9609), .B2(n5984), .A(n5914), .ZN(n5916) );
  NAND2_X1 U7569 ( .A1(n5915), .A2(n5916), .ZN(n9018) );
  NAND2_X1 U7570 ( .A1(n9019), .A2(n9018), .ZN(n8929) );
  INV_X1 U7571 ( .A(n5915), .ZN(n5918) );
  INV_X1 U7572 ( .A(n5916), .ZN(n5917) );
  NAND2_X1 U7573 ( .A1(n5918), .A2(n5917), .ZN(n9017) );
  NAND2_X1 U7574 ( .A1(n9588), .A2(n5978), .ZN(n5920) );
  NAND2_X1 U7575 ( .A1(n9699), .A2(n5984), .ZN(n5919) );
  NAND2_X1 U7576 ( .A1(n5920), .A2(n5919), .ZN(n5921) );
  XNOR2_X1 U7577 ( .A(n5921), .B(n5987), .ZN(n5926) );
  AND2_X1 U7578 ( .A1(n9699), .A2(n5981), .ZN(n5922) );
  AOI21_X1 U7579 ( .B1(n9588), .B2(n5984), .A(n5922), .ZN(n5925) );
  XNOR2_X1 U7580 ( .A(n5926), .B(n5925), .ZN(n8933) );
  INV_X1 U7581 ( .A(n8933), .ZN(n5923) );
  AND2_X1 U7582 ( .A1(n9017), .A2(n5923), .ZN(n5924) );
  NAND2_X1 U7583 ( .A1(n8929), .A2(n5924), .ZN(n8930) );
  NAND2_X1 U7584 ( .A1(n5926), .A2(n5925), .ZN(n5927) );
  NAND2_X1 U7585 ( .A1(n8930), .A2(n5927), .ZN(n8999) );
  NAND2_X1 U7586 ( .A1(n7895), .A2(n5978), .ZN(n5929) );
  NAND2_X1 U7587 ( .A1(n9583), .A2(n5984), .ZN(n5928) );
  NAND2_X1 U7588 ( .A1(n5929), .A2(n5928), .ZN(n5930) );
  XNOR2_X1 U7589 ( .A(n5930), .B(n5979), .ZN(n5932) );
  NOR2_X1 U7590 ( .A1(n9691), .A2(n5827), .ZN(n5931) );
  AOI21_X1 U7591 ( .B1(n7895), .B2(n5984), .A(n5931), .ZN(n5933) );
  XNOR2_X1 U7592 ( .A(n5932), .B(n5933), .ZN(n9000) );
  NAND2_X1 U7593 ( .A1(n8999), .A2(n9000), .ZN(n8998) );
  INV_X1 U7594 ( .A(n5932), .ZN(n5934) );
  NAND2_X1 U7595 ( .A1(n5934), .A2(n5933), .ZN(n5935) );
  NAND2_X1 U7596 ( .A1(n9676), .A2(n5978), .ZN(n5937) );
  NAND2_X1 U7597 ( .A1(n9312), .A2(n5984), .ZN(n5936) );
  NAND2_X1 U7598 ( .A1(n5937), .A2(n5936), .ZN(n5938) );
  XNOR2_X1 U7599 ( .A(n5938), .B(n5979), .ZN(n5940) );
  NOR2_X1 U7600 ( .A1(n9681), .A2(n5827), .ZN(n5939) );
  AOI21_X1 U7601 ( .B1(n9676), .B2(n5984), .A(n5939), .ZN(n5941) );
  XNOR2_X1 U7602 ( .A(n5940), .B(n5941), .ZN(n8940) );
  INV_X1 U7603 ( .A(n5940), .ZN(n5942) );
  NAND2_X1 U7604 ( .A1(n9665), .A2(n5978), .ZN(n5944) );
  NAND2_X1 U7605 ( .A1(n9311), .A2(n5984), .ZN(n5943) );
  NAND2_X1 U7606 ( .A1(n5944), .A2(n5943), .ZN(n5945) );
  XNOR2_X1 U7607 ( .A(n5945), .B(n5987), .ZN(n8917) );
  NOR2_X1 U7608 ( .A1(n9659), .A2(n5827), .ZN(n5946) );
  AOI21_X1 U7609 ( .B1(n9665), .B2(n5984), .A(n5946), .ZN(n8916) );
  NOR2_X1 U7610 ( .A1(n8917), .A2(n8916), .ZN(n8915) );
  NAND2_X1 U7611 ( .A1(n9740), .A2(n5978), .ZN(n5948) );
  NAND2_X1 U7612 ( .A1(n9555), .A2(n5984), .ZN(n5947) );
  NAND2_X1 U7613 ( .A1(n5948), .A2(n5947), .ZN(n5949) );
  XNOR2_X1 U7614 ( .A(n5949), .B(n5979), .ZN(n8919) );
  NAND2_X1 U7615 ( .A1(n9740), .A2(n5984), .ZN(n5951) );
  NAND2_X1 U7616 ( .A1(n9555), .A2(n5981), .ZN(n5950) );
  NAND2_X1 U7617 ( .A1(n5951), .A2(n5950), .ZN(n8918) );
  INV_X1 U7618 ( .A(n8916), .ZN(n5953) );
  OAI21_X1 U7619 ( .B1(n8919), .B2(n8918), .A(n5953), .ZN(n5952) );
  NOR3_X1 U7620 ( .A1(n8919), .A2(n5953), .A3(n8918), .ZN(n5954) );
  NAND2_X1 U7621 ( .A1(n9540), .A2(n5978), .ZN(n5957) );
  NAND2_X1 U7622 ( .A1(n9556), .A2(n5984), .ZN(n5956) );
  NAND2_X1 U7623 ( .A1(n5957), .A2(n5956), .ZN(n5958) );
  XNOR2_X1 U7624 ( .A(n5958), .B(n5987), .ZN(n5961) );
  NOR2_X1 U7625 ( .A1(n9648), .A2(n5827), .ZN(n5959) );
  AOI21_X1 U7626 ( .B1(n9540), .B2(n5984), .A(n5959), .ZN(n5960) );
  NAND2_X1 U7627 ( .A1(n5961), .A2(n5960), .ZN(n5962) );
  OAI21_X1 U7628 ( .B1(n5961), .B2(n5960), .A(n5962), .ZN(n8989) );
  NAND2_X1 U7629 ( .A1(n9731), .A2(n5978), .ZN(n5964) );
  NAND2_X1 U7630 ( .A1(n9530), .A2(n5984), .ZN(n5963) );
  NAND2_X1 U7631 ( .A1(n5964), .A2(n5963), .ZN(n5965) );
  XNOR2_X1 U7632 ( .A(n5965), .B(n5979), .ZN(n5972) );
  OAI22_X1 U7633 ( .A1(n7879), .A2(n5966), .B1(n8994), .B2(n5827), .ZN(n5971)
         );
  XNOR2_X1 U7634 ( .A(n5972), .B(n5971), .ZN(n8961) );
  NAND2_X1 U7635 ( .A1(n9522), .A2(n5978), .ZN(n5968) );
  NAND2_X1 U7636 ( .A1(n9498), .A2(n5984), .ZN(n5967) );
  NAND2_X1 U7637 ( .A1(n5968), .A2(n5967), .ZN(n5969) );
  XNOR2_X1 U7638 ( .A(n5969), .B(n5987), .ZN(n5974) );
  NOR2_X1 U7639 ( .A1(n9649), .A2(n5827), .ZN(n5970) );
  AOI21_X1 U7640 ( .B1(n9522), .B2(n5984), .A(n5970), .ZN(n5975) );
  XNOR2_X1 U7641 ( .A(n5974), .B(n5975), .ZN(n9027) );
  NOR2_X1 U7642 ( .A1(n5972), .A2(n5971), .ZN(n9028) );
  INV_X1 U7643 ( .A(n5974), .ZN(n5977) );
  INV_X1 U7644 ( .A(n5975), .ZN(n5976) );
  AOI22_X1 U7645 ( .A1(n4847), .A2(n5978), .B1(n5984), .B2(n9515), .ZN(n5980)
         );
  XNOR2_X1 U7646 ( .A(n5980), .B(n5979), .ZN(n5983) );
  AOI22_X1 U7647 ( .A1(n4847), .A2(n5984), .B1(n5981), .B2(n9515), .ZN(n5982)
         );
  NAND2_X1 U7648 ( .A1(n5983), .A2(n5982), .ZN(n6022) );
  OAI21_X1 U7649 ( .B1(n5983), .B2(n5982), .A(n6022), .ZN(n7949) );
  INV_X1 U7650 ( .A(n7951), .ZN(n5998) );
  NAND2_X1 U7651 ( .A1(n9488), .A2(n5978), .ZN(n5986) );
  NAND2_X1 U7652 ( .A1(n9497), .A2(n5984), .ZN(n5985) );
  NAND2_X1 U7653 ( .A1(n5986), .A2(n5985), .ZN(n5988) );
  XNOR2_X1 U7654 ( .A(n5988), .B(n5987), .ZN(n5991) );
  NAND2_X1 U7655 ( .A1(n9488), .A2(n5984), .ZN(n5989) );
  OAI21_X1 U7656 ( .B1(n7953), .B2(n5827), .A(n5989), .ZN(n5990) );
  XNOR2_X1 U7657 ( .A(n5991), .B(n5990), .ZN(n5999) );
  INV_X1 U7658 ( .A(n5999), .ZN(n6023) );
  NOR2_X1 U7659 ( .A1(n5993), .A2(n5992), .ZN(n5994) );
  OR3_X1 U7660 ( .A1(n5995), .A2(n7128), .A3(n5994), .ZN(n6014) );
  NAND2_X1 U7661 ( .A1(n9944), .A2(n5996), .ZN(n6006) );
  OR2_X1 U7662 ( .A1(n9304), .A2(n6006), .ZN(n5997) );
  NOR2_X2 U7663 ( .A1(n6014), .A2(n5997), .ZN(n9031) );
  NAND2_X1 U7664 ( .A1(n5998), .A2(n5060), .ZN(n6028) );
  NAND3_X1 U7665 ( .A1(n7951), .A2(n5999), .A3(n9031), .ZN(n6027) );
  INV_X1 U7666 ( .A(n6014), .ZN(n6001) );
  OR2_X1 U7667 ( .A1(n6803), .A2(n9298), .ZN(n7132) );
  NOR2_X1 U7668 ( .A1(n9304), .A2(n7132), .ZN(n6000) );
  NAND2_X1 U7669 ( .A1(n6001), .A2(n6000), .ZN(n6003) );
  INV_X1 U7670 ( .A(n9303), .ZN(n7136) );
  NAND2_X1 U7671 ( .A1(n6004), .A2(n7136), .ZN(n6012) );
  NOR2_X1 U7672 ( .A1(n6014), .A2(n6012), .ZN(n6018) );
  INV_X1 U7673 ( .A(n4443), .ZN(n6815) );
  NAND2_X1 U7674 ( .A1(n6018), .A2(n6815), .ZN(n8983) );
  INV_X1 U7675 ( .A(n6005), .ZN(n9489) );
  INV_X1 U7676 ( .A(n6006), .ZN(n6007) );
  NAND2_X1 U7677 ( .A1(n6014), .A2(n6007), .ZN(n6010) );
  AND3_X1 U7678 ( .A1(n6008), .A2(n6539), .A3(n6585), .ZN(n6009) );
  NAND2_X1 U7679 ( .A1(n6010), .A2(n6009), .ZN(n6011) );
  NAND2_X1 U7680 ( .A1(n6011), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6016) );
  OAI21_X1 U7681 ( .B1(n7132), .B2(P1_U3086), .A(n6012), .ZN(n6013) );
  NAND2_X1 U7682 ( .A1(n6014), .A2(n6013), .ZN(n6015) );
  NAND2_X1 U7683 ( .A1(n6016), .A2(n6015), .ZN(n8991) );
  AOI22_X1 U7684 ( .A1(n9489), .A2(n8991), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6020) );
  INV_X1 U7685 ( .A(n6017), .ZN(n9482) );
  NAND2_X1 U7686 ( .A1(n6018), .A2(n4443), .ZN(n9043) );
  INV_X1 U7687 ( .A(n9043), .ZN(n9036) );
  NAND2_X1 U7688 ( .A1(n9482), .A2(n9036), .ZN(n6019) );
  OAI211_X1 U7689 ( .C1(n6021), .C2(n8983), .A(n6020), .B(n6019), .ZN(n6025)
         );
  NOR3_X1 U7690 ( .A1(n6023), .A2(n6022), .A3(n9052), .ZN(n6024) );
  AOI211_X1 U7691 ( .C1(n9488), .C2(n9050), .A(n6025), .B(n6024), .ZN(n6026)
         );
  NAND3_X1 U7692 ( .A1(n6028), .A2(n6027), .A3(n6026), .ZN(P1_U3220) );
  AND2_X2 U7693 ( .A1(n6734), .A2(n4773), .ZN(n6084) );
  NAND3_X1 U7694 ( .A1(n6508), .A2(n6484), .A3(n6485), .ZN(n6039) );
  INV_X1 U7695 ( .A(n6058), .ZN(n6042) );
  NAND2_X1 U7696 ( .A1(n6042), .A2(n10268), .ZN(n6045) );
  INV_X1 U7697 ( .A(n6045), .ZN(n6043) );
  NAND2_X1 U7698 ( .A1(n6043), .A2(n6046), .ZN(n8893) );
  XNOR2_X2 U7699 ( .A(n6044), .B(n8894), .ZN(n6064) );
  INV_X1 U7700 ( .A(n4444), .ZN(n6049) );
  NAND2_X1 U7701 ( .A1(n6049), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6055) );
  INV_X1 U7702 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6997) );
  NAND2_X1 U7703 ( .A1(P2_REG2_REG_1__SCAN_IN), .A2(n6050), .ZN(n6051) );
  NAND2_X1 U7704 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6061) );
  MUX2_X1 U7705 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6061), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n6063) );
  INV_X1 U7706 ( .A(n6734), .ZN(n6062) );
  NAND2_X1 U7707 ( .A1(n6063), .A2(n6062), .ZN(n9995) );
  INV_X1 U7708 ( .A(n8192), .ZN(n8304) );
  INV_X1 U7709 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6655) );
  INV_X1 U7710 ( .A(n6064), .ZN(n6065) );
  INV_X1 U7711 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6934) );
  INV_X1 U7712 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6779) );
  OR2_X1 U7713 ( .A1(n4441), .A2(n6779), .ZN(n6067) );
  NAND2_X1 U7714 ( .A1(n6077), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6066) );
  NAND4_X1 U7715 ( .A1(n6069), .A2(n6068), .A3(n6067), .A4(n6066), .ZN(n6424)
         );
  INV_X1 U7716 ( .A(n6424), .ZN(n6076) );
  INV_X1 U7717 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6733) );
  NAND2_X1 U7718 ( .A1(n6549), .A2(SI_0_), .ZN(n6071) );
  INV_X1 U7719 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7720 ( .A1(n6071), .A2(n6070), .ZN(n6073) );
  NAND2_X1 U7721 ( .A1(n6073), .A2(n6072), .ZN(n8902) );
  MUX2_X1 U7722 ( .A(n6733), .B(n8902), .S(n6074), .Z(n6936) );
  NAND2_X1 U7723 ( .A1(n6076), .A2(n6075), .ZN(n6881) );
  INV_X1 U7724 ( .A(n6881), .ZN(n6907) );
  NAND2_X1 U7725 ( .A1(n8304), .A2(n6907), .ZN(n6906) );
  NAND2_X1 U7726 ( .A1(n6906), .A2(n8188), .ZN(n7105) );
  INV_X1 U7727 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7115) );
  NAND2_X1 U7728 ( .A1(n6077), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6081) );
  INV_X1 U7729 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6078) );
  OR2_X1 U7730 ( .A1(n4444), .A2(n6078), .ZN(n6080) );
  INV_X1 U7731 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6890) );
  OR2_X1 U7732 ( .A1(n4441), .A2(n6890), .ZN(n6079) );
  NOR2_X1 U7733 ( .A1(n6734), .A2(n6209), .ZN(n6083) );
  INV_X1 U7734 ( .A(n6084), .ZN(n6085) );
  OR2_X1 U7735 ( .A1(n8133), .A2(n6555), .ZN(n6087) );
  OR2_X1 U7736 ( .A1(n6109), .A2(n6554), .ZN(n6086) );
  OAI211_X1 U7737 ( .C1(n6074), .C2(n6737), .A(n6087), .B(n6086), .ZN(n6887)
         );
  INV_X1 U7738 ( .A(n6887), .ZN(n10006) );
  INV_X1 U7739 ( .A(n6426), .ZN(n7103) );
  INV_X1 U7740 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6713) );
  INV_X1 U7741 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6714) );
  OR2_X1 U7742 ( .A1(n6292), .A2(n6714), .ZN(n6089) );
  NAND2_X1 U7743 ( .A1(n6077), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6092) );
  OR2_X1 U7744 ( .A1(n6109), .A2(n6556), .ZN(n6100) );
  OR2_X1 U7745 ( .A1(n8133), .A2(n6557), .ZN(n6099) );
  NOR2_X1 U7746 ( .A1(n6084), .A2(n6209), .ZN(n6095) );
  MUX2_X1 U7747 ( .A(n6209), .B(n6095), .S(P2_IR_REG_3__SCAN_IN), .Z(n6097) );
  NAND2_X1 U7748 ( .A1(n6646), .A2(n6782), .ZN(n6098) );
  NAND2_X1 U7749 ( .A1(n8351), .A2(n7008), .ZN(n8205) );
  NAND2_X1 U7750 ( .A1(n6365), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6108) );
  INV_X1 U7751 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6102) );
  OR2_X1 U7752 ( .A1(n4430), .A2(n6102), .ZN(n6107) );
  NAND2_X1 U7753 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6104) );
  AND2_X1 U7754 ( .A1(n6117), .A2(n6104), .ZN(n7015) );
  OR2_X1 U7755 ( .A1(n4441), .A2(n7015), .ZN(n6106) );
  INV_X1 U7756 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7123) );
  OR2_X1 U7757 ( .A1(n4440), .A2(n7123), .ZN(n6105) );
  OR2_X1 U7758 ( .A1(n6109), .A2(n6568), .ZN(n6114) );
  INV_X1 U7759 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6569) );
  OR2_X1 U7760 ( .A1(n8133), .A2(n6569), .ZN(n6113) );
  NAND2_X1 U7761 ( .A1(n6123), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6111) );
  XNOR2_X2 U7762 ( .A(n6111), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6852) );
  NAND2_X1 U7763 ( .A1(n6646), .A2(n6852), .ZN(n6112) );
  OR2_X1 U7764 ( .A1(n7998), .A2(n7003), .ZN(n8206) );
  NAND2_X1 U7765 ( .A1(n7998), .A2(n7003), .ZN(n8213) );
  NAND2_X1 U7766 ( .A1(n8206), .A2(n8213), .ZN(n6428) );
  INV_X1 U7767 ( .A(n6428), .ZN(n8303) );
  NAND2_X1 U7768 ( .A1(n7117), .A2(n8303), .ZN(n7118) );
  NAND2_X1 U7769 ( .A1(n7118), .A2(n8206), .ZN(n7097) );
  NAND2_X1 U7770 ( .A1(n4433), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6122) );
  INV_X1 U7771 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6844) );
  OR2_X1 U7772 ( .A1(n4445), .A2(n6844), .ZN(n6121) );
  NAND2_X1 U7773 ( .A1(n6117), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6118) );
  AND2_X1 U7774 ( .A1(n6128), .A2(n6118), .ZN(n7098) );
  OR2_X1 U7775 ( .A1(n4441), .A2(n7098), .ZN(n6120) );
  INV_X1 U7776 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6845) );
  OR2_X1 U7777 ( .A1(n4440), .A2(n6845), .ZN(n6119) );
  NAND4_X1 U7778 ( .A1(n6122), .A2(n6121), .A3(n6120), .A4(n6119), .ZN(n8350)
         );
  NAND2_X1 U7779 ( .A1(n6134), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6124) );
  XNOR2_X1 U7780 ( .A(n6124), .B(n6135), .ZN(n6861) );
  OR2_X1 U7781 ( .A1(n6109), .A2(n6560), .ZN(n6126) );
  INV_X1 U7782 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6561) );
  OR2_X1 U7783 ( .A1(n8133), .A2(n6561), .ZN(n6125) );
  OAI211_X1 U7784 ( .C1(n6074), .C2(n6861), .A(n6126), .B(n6125), .ZN(n10022)
         );
  INV_X1 U7785 ( .A(n10022), .ZN(n7099) );
  NAND2_X1 U7786 ( .A1(n8350), .A2(n7099), .ZN(n8212) );
  AND2_X1 U7787 ( .A1(n8217), .A2(n8212), .ZN(n7096) );
  NAND2_X1 U7788 ( .A1(n7097), .A2(n7096), .ZN(n6127) );
  NAND2_X1 U7789 ( .A1(n4433), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6133) );
  INV_X1 U7790 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7251) );
  OR2_X1 U7791 ( .A1(n4440), .A2(n7251), .ZN(n6132) );
  NAND2_X1 U7792 ( .A1(n6128), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6129) );
  AND2_X1 U7793 ( .A1(n6144), .A2(n6129), .ZN(n7252) );
  OR2_X1 U7794 ( .A1(n4441), .A2(n7252), .ZN(n6131) );
  INV_X1 U7795 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7082) );
  OR2_X1 U7796 ( .A1(n4445), .A2(n7082), .ZN(n6130) );
  NAND4_X1 U7797 ( .A1(n6133), .A2(n6132), .A3(n6131), .A4(n6130), .ZN(n8349)
         );
  INV_X1 U7798 ( .A(n6134), .ZN(n6136) );
  NAND2_X1 U7799 ( .A1(n6136), .A2(n6135), .ZN(n6150) );
  NAND2_X1 U7800 ( .A1(n6150), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6138) );
  INV_X1 U7801 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6137) );
  XNOR2_X1 U7802 ( .A(n6138), .B(n6137), .ZN(n7075) );
  OR2_X1 U7803 ( .A1(n6109), .A2(n6563), .ZN(n6140) );
  OR2_X1 U7804 ( .A1(n8133), .A2(n6562), .ZN(n6139) );
  OAI211_X1 U7805 ( .C1(n6074), .C2(n7075), .A(n6140), .B(n6139), .ZN(n10028)
         );
  INV_X1 U7806 ( .A(n10028), .ZN(n7063) );
  OR2_X1 U7807 ( .A1(n8349), .A2(n7063), .ZN(n8215) );
  INV_X1 U7808 ( .A(n8215), .ZN(n6141) );
  NAND2_X1 U7809 ( .A1(n8349), .A2(n7063), .ZN(n8209) );
  NAND2_X1 U7810 ( .A1(n4433), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6149) );
  INV_X1 U7811 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7071) );
  OR2_X1 U7812 ( .A1(n4440), .A2(n7071), .ZN(n6148) );
  NAND2_X1 U7813 ( .A1(n6144), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6145) );
  AND2_X1 U7814 ( .A1(n6157), .A2(n6145), .ZN(n7446) );
  OR2_X1 U7815 ( .A1(n4441), .A2(n7446), .ZN(n6147) );
  INV_X1 U7816 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7070) );
  OR2_X1 U7817 ( .A1(n4445), .A2(n7070), .ZN(n6146) );
  NAND4_X1 U7818 ( .A1(n6149), .A2(n6148), .A3(n6147), .A4(n6146), .ZN(n8348)
         );
  OR2_X1 U7819 ( .A1(n6109), .A2(n6566), .ZN(n6154) );
  OR2_X1 U7820 ( .A1(n8133), .A2(n6565), .ZN(n6153) );
  OAI21_X1 U7821 ( .B1(n6150), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6151) );
  XNOR2_X1 U7822 ( .A(n6151), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7079) );
  NAND2_X1 U7823 ( .A1(n6646), .A2(n7079), .ZN(n6152) );
  OR2_X1 U7824 ( .A1(n8348), .A2(n7515), .ZN(n8160) );
  NAND2_X1 U7825 ( .A1(n8348), .A2(n7515), .ZN(n8153) );
  NAND2_X1 U7826 ( .A1(n4433), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6162) );
  INV_X1 U7827 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6156) );
  OR2_X1 U7828 ( .A1(n4445), .A2(n6156), .ZN(n6161) );
  NAND2_X1 U7829 ( .A1(n6157), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6158) );
  AND2_X1 U7830 ( .A1(n6171), .A2(n6158), .ZN(n7287) );
  OR2_X1 U7831 ( .A1(n4441), .A2(n7287), .ZN(n6160) );
  INV_X1 U7832 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7656) );
  OR2_X1 U7833 ( .A1(n4440), .A2(n7656), .ZN(n6159) );
  NAND4_X1 U7834 ( .A1(n6162), .A2(n6161), .A3(n6160), .A4(n6159), .ZN(n8347)
         );
  OR2_X1 U7835 ( .A1(n6164), .A2(n6209), .ZN(n6165) );
  XNOR2_X1 U7836 ( .A(n6165), .B(n6178), .ZN(n7402) );
  INV_X1 U7837 ( .A(n7402), .ZN(n7189) );
  AOI22_X1 U7838 ( .A1(n6301), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6646), .B2(
        n7189), .ZN(n6167) );
  NAND2_X1 U7839 ( .A1(n6570), .A2(n6183), .ZN(n6166) );
  NAND2_X1 U7840 ( .A1(n6167), .A2(n6166), .ZN(n7658) );
  INV_X1 U7841 ( .A(n7658), .ZN(n10034) );
  AND2_X1 U7842 ( .A1(n8347), .A2(n10034), .ZN(n8154) );
  OR2_X1 U7843 ( .A1(n8347), .A2(n10034), .ZN(n8161) );
  NAND2_X1 U7844 ( .A1(n4433), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6177) );
  INV_X1 U7845 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6168) );
  OR2_X1 U7846 ( .A1(n4445), .A2(n6168), .ZN(n6176) );
  NAND2_X1 U7847 ( .A1(n6171), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6172) );
  AND2_X1 U7848 ( .A1(n6188), .A2(n6172), .ZN(n7550) );
  OR2_X1 U7849 ( .A1(n4441), .A2(n7550), .ZN(n6175) );
  INV_X1 U7850 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6173) );
  OR2_X1 U7851 ( .A1(n4439), .A2(n6173), .ZN(n6174) );
  NAND2_X1 U7852 ( .A1(n6574), .A2(n6183), .ZN(n6181) );
  NAND2_X1 U7853 ( .A1(n6164), .A2(n6178), .ZN(n6184) );
  NAND2_X1 U7854 ( .A1(n6184), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6179) );
  XNOR2_X1 U7855 ( .A(n6179), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7427) );
  AOI22_X1 U7856 ( .A1(n6301), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6646), .B2(
        n7427), .ZN(n6180) );
  NAND2_X1 U7857 ( .A1(n6181), .A2(n6180), .ZN(n7688) );
  NAND2_X1 U7858 ( .A1(n7292), .A2(n7688), .ZN(n8162) );
  NAND2_X1 U7859 ( .A1(n6578), .A2(n6183), .ZN(n6187) );
  NAND2_X1 U7860 ( .A1(n6194), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6185) );
  XNOR2_X1 U7861 ( .A(n6185), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7431) );
  AOI22_X1 U7862 ( .A1(n6301), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6646), .B2(
        n7431), .ZN(n6186) );
  NAND2_X1 U7863 ( .A1(n4433), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6193) );
  INV_X1 U7864 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7430) );
  OR2_X1 U7865 ( .A1(n4445), .A2(n7430), .ZN(n6192) );
  NAND2_X1 U7866 ( .A1(n6188), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6189) );
  AND2_X1 U7867 ( .A1(n6199), .A2(n6189), .ZN(n7638) );
  OR2_X1 U7868 ( .A1(n4441), .A2(n7638), .ZN(n6191) );
  INV_X1 U7869 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7639) );
  OR2_X1 U7870 ( .A1(n4440), .A2(n7639), .ZN(n6190) );
  NAND4_X1 U7871 ( .A1(n6193), .A2(n6192), .A3(n6191), .A4(n6190), .ZN(n8345)
         );
  OR2_X1 U7872 ( .A1(n10049), .A2(n7708), .ZN(n7631) );
  NAND2_X1 U7873 ( .A1(n10049), .A2(n7708), .ZN(n8163) );
  NAND2_X1 U7874 ( .A1(n6662), .A2(n6183), .ZN(n6197) );
  NOR2_X1 U7875 ( .A1(n6194), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n6207) );
  OR2_X1 U7876 ( .A1(n6207), .A2(n6209), .ZN(n6195) );
  XNOR2_X1 U7877 ( .A(n6195), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7581) );
  AOI22_X1 U7878 ( .A1(n6301), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6646), .B2(
        n7581), .ZN(n6196) );
  NAND2_X1 U7879 ( .A1(n4433), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6204) );
  INV_X1 U7880 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6198) );
  OR2_X1 U7881 ( .A1(n4445), .A2(n6198), .ZN(n6203) );
  NAND2_X1 U7882 ( .A1(n6199), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6200) );
  AND2_X1 U7883 ( .A1(n6218), .A2(n6200), .ZN(n7747) );
  OR2_X1 U7884 ( .A1(n4441), .A2(n7747), .ZN(n6202) );
  INV_X1 U7885 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7711) );
  OR2_X1 U7886 ( .A1(n4439), .A2(n7711), .ZN(n6201) );
  NAND4_X1 U7887 ( .A1(n6204), .A2(n6203), .A3(n6202), .A4(n6201), .ZN(n8344)
         );
  INV_X1 U7888 ( .A(n8344), .ZN(n7767) );
  NAND2_X1 U7889 ( .A1(n10054), .A2(n7767), .ZN(n8177) );
  INV_X1 U7890 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6206) );
  AND2_X1 U7891 ( .A1(n6207), .A2(n6206), .ZN(n6212) );
  NOR2_X1 U7892 ( .A1(n6212), .A2(n6209), .ZN(n6208) );
  MUX2_X1 U7893 ( .A(n6209), .B(n6208), .S(P2_IR_REG_12__SCAN_IN), .Z(n6210)
         );
  INV_X1 U7894 ( .A(n6210), .ZN(n6213) );
  INV_X1 U7895 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7896 ( .A1(n6212), .A2(n6211), .ZN(n6225) );
  AOI22_X1 U7897 ( .A1(n6301), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6646), .B2(
        n7587), .ZN(n6214) );
  NAND2_X1 U7898 ( .A1(n4433), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6224) );
  INV_X1 U7899 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7900 ( .A1(n6218), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6219) );
  AND2_X1 U7901 ( .A1(n6230), .A2(n6219), .ZN(n7784) );
  OR2_X1 U7902 ( .A1(n4441), .A2(n7784), .ZN(n6223) );
  INV_X1 U7903 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6220) );
  OR2_X1 U7904 ( .A1(n4439), .A2(n6220), .ZN(n6222) );
  OR2_X1 U7905 ( .A1(n4445), .A2(n8355), .ZN(n6221) );
  NAND4_X1 U7906 ( .A1(n6224), .A2(n6223), .A3(n6222), .A4(n6221), .ZN(n8343)
         );
  NAND2_X1 U7907 ( .A1(n10060), .A2(n8741), .ZN(n8178) );
  NAND2_X1 U7908 ( .A1(n6752), .A2(n6183), .ZN(n6227) );
  NAND2_X1 U7909 ( .A1(n6225), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6237) );
  XNOR2_X1 U7910 ( .A(n6237), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8397) );
  AOI22_X1 U7911 ( .A1(n6301), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6646), .B2(
        n8397), .ZN(n6226) );
  NAND2_X1 U7912 ( .A1(n4433), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6235) );
  INV_X1 U7913 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8364) );
  OR2_X1 U7914 ( .A1(n4445), .A2(n8364), .ZN(n6234) );
  INV_X1 U7915 ( .A(n6230), .ZN(n6229) );
  INV_X1 U7916 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6228) );
  NAND2_X1 U7917 ( .A1(n6230), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6231) );
  AND2_X1 U7918 ( .A1(n6241), .A2(n6231), .ZN(n8746) );
  OR2_X1 U7919 ( .A1(n4441), .A2(n8746), .ZN(n6233) );
  INV_X1 U7920 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8365) );
  OR2_X1 U7921 ( .A1(n4440), .A2(n8365), .ZN(n6232) );
  INV_X1 U7922 ( .A(n8317), .ZN(n9774) );
  NAND2_X1 U7923 ( .A1(n6830), .A2(n6183), .ZN(n6240) );
  INV_X1 U7924 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7925 ( .A1(n6237), .A2(n6236), .ZN(n6238) );
  NAND2_X1 U7926 ( .A1(n6238), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6249) );
  XNOR2_X1 U7927 ( .A(n6249), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8409) );
  AOI22_X1 U7928 ( .A1(n6301), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6646), .B2(
        n8409), .ZN(n6239) );
  NAND2_X1 U7929 ( .A1(n6365), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6246) );
  INV_X1 U7930 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8886) );
  OR2_X1 U7931 ( .A1(n4430), .A2(n8886), .ZN(n6245) );
  NAND2_X1 U7932 ( .A1(n6241), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6242) );
  AND2_X1 U7933 ( .A1(n6264), .A2(n6242), .ZN(n8724) );
  OR2_X1 U7934 ( .A1(n4441), .A2(n8724), .ZN(n6244) );
  INV_X1 U7935 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8408) );
  OR2_X1 U7936 ( .A1(n4439), .A2(n8408), .ZN(n6243) );
  NAND4_X1 U7937 ( .A1(n6246), .A2(n6245), .A3(n6244), .A4(n6243), .ZN(n8714)
         );
  OR2_X1 U7938 ( .A1(n8887), .A2(n8743), .ZN(n8226) );
  NAND2_X1 U7939 ( .A1(n8735), .A2(n8226), .ZN(n6247) );
  NAND2_X1 U7940 ( .A1(n8887), .A2(n8743), .ZN(n8228) );
  NAND2_X1 U7941 ( .A1(n6944), .A2(n6183), .ZN(n6253) );
  NAND2_X1 U7942 ( .A1(n6249), .A2(n6248), .ZN(n6250) );
  NAND2_X1 U7943 ( .A1(n6250), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6261) );
  INV_X1 U7944 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n10266) );
  NAND2_X1 U7945 ( .A1(n6261), .A2(n10266), .ZN(n6251) );
  NAND2_X1 U7946 ( .A1(n6251), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6273) );
  XNOR2_X1 U7947 ( .A(n6273), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8456) );
  AOI22_X1 U7948 ( .A1(n6301), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6646), .B2(
        n8456), .ZN(n6252) );
  NAND2_X1 U7949 ( .A1(n4433), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6260) );
  INV_X1 U7950 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8799) );
  OR2_X1 U7951 ( .A1(n4445), .A2(n8799), .ZN(n6259) );
  INV_X1 U7952 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U7953 ( .A1(n6266), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6256) );
  AND2_X1 U7954 ( .A1(n6280), .A2(n6256), .ZN(n8706) );
  OR2_X1 U7955 ( .A1(n4441), .A2(n8706), .ZN(n6258) );
  INV_X1 U7956 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8445) );
  OR2_X1 U7957 ( .A1(n4439), .A2(n8445), .ZN(n6257) );
  NAND4_X1 U7958 ( .A1(n6260), .A2(n6259), .A3(n6258), .A4(n6257), .ZN(n8713)
         );
  NAND2_X1 U7959 ( .A1(n8879), .A2(n8111), .ZN(n6449) );
  NAND2_X1 U7960 ( .A1(n6902), .A2(n6183), .ZN(n6263) );
  XNOR2_X1 U7961 ( .A(n6261), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8453) );
  AOI22_X1 U7962 ( .A1(n6301), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6646), .B2(
        n8453), .ZN(n6262) );
  NAND2_X1 U7963 ( .A1(n4433), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6270) );
  INV_X1 U7964 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8432) );
  OR2_X1 U7965 ( .A1(n4445), .A2(n8432), .ZN(n6269) );
  NAND2_X1 U7966 ( .A1(n6264), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6265) );
  AND2_X1 U7967 ( .A1(n6266), .A2(n6265), .ZN(n8108) );
  OR2_X1 U7968 ( .A1(n4441), .A2(n8108), .ZN(n6268) );
  INV_X1 U7969 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8413) );
  OR2_X1 U7970 ( .A1(n4440), .A2(n8413), .ZN(n6267) );
  NAND4_X1 U7971 ( .A1(n6270), .A2(n6269), .A3(n6268), .A4(n6267), .ZN(n8729)
         );
  NAND2_X1 U7972 ( .A1(n8803), .A2(n8302), .ZN(n8698) );
  NAND2_X1 U7973 ( .A1(n6449), .A2(n8698), .ZN(n8227) );
  OR2_X1 U7974 ( .A1(n8803), .A2(n8302), .ZN(n8699) );
  NAND2_X1 U7975 ( .A1(n8232), .A2(n8699), .ZN(n6271) );
  NAND2_X1 U7976 ( .A1(n6271), .A2(n6449), .ZN(n8229) );
  NAND2_X1 U7977 ( .A1(n7052), .A2(n6183), .ZN(n6277) );
  NAND2_X1 U7978 ( .A1(n6273), .A2(n6272), .ZN(n6274) );
  NAND2_X1 U7979 ( .A1(n6274), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6275) );
  XNOR2_X1 U7980 ( .A(n6275), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8502) );
  AOI22_X1 U7981 ( .A1(n6301), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6646), .B2(
        n8502), .ZN(n6276) );
  NAND2_X1 U7982 ( .A1(n4433), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6285) );
  INV_X1 U7983 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8470) );
  OR2_X1 U7984 ( .A1(n4445), .A2(n8470), .ZN(n6284) );
  INV_X1 U7985 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U7986 ( .A1(n6280), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6281) );
  AND2_X1 U7987 ( .A1(n6290), .A2(n6281), .ZN(n8692) );
  OR2_X1 U7988 ( .A1(n4441), .A2(n8692), .ZN(n6283) );
  INV_X1 U7989 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8693) );
  OR2_X1 U7990 ( .A1(n4440), .A2(n8693), .ZN(n6282) );
  NAND4_X1 U7991 ( .A1(n6285), .A2(n6284), .A3(n6283), .A4(n6282), .ZN(n8704)
         );
  INV_X1 U7992 ( .A(n8704), .ZN(n8033) );
  OR2_X1 U7993 ( .A1(n8795), .A2(n8033), .ZN(n8242) );
  NAND2_X1 U7994 ( .A1(n8795), .A2(n8033), .ZN(n8238) );
  NAND2_X1 U7995 ( .A1(n8242), .A2(n8238), .ZN(n8689) );
  INV_X1 U7996 ( .A(n8673), .ZN(n6298) );
  NAND2_X1 U7997 ( .A1(n7143), .A2(n6183), .ZN(n6289) );
  NAND2_X1 U7998 ( .A1(n6286), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6287) );
  XNOR2_X1 U7999 ( .A(n6287), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8522) );
  AOI22_X1 U8000 ( .A1(n6301), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6646), .B2(
        n8522), .ZN(n6288) );
  NAND2_X1 U8001 ( .A1(n6365), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6296) );
  INV_X1 U8002 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8871) );
  OR2_X1 U8003 ( .A1(n4430), .A2(n8871), .ZN(n6295) );
  NAND2_X1 U8004 ( .A1(n6290), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6291) );
  AND2_X1 U8005 ( .A1(n6305), .A2(n6291), .ZN(n8085) );
  OR2_X1 U8006 ( .A1(n4441), .A2(n8085), .ZN(n6294) );
  INV_X1 U8007 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8680) );
  OR2_X1 U8008 ( .A1(n4440), .A2(n8680), .ZN(n6293) );
  NAND2_X1 U8009 ( .A1(n8872), .A2(n8659), .ZN(n8239) );
  NAND2_X1 U8010 ( .A1(n8249), .A2(n8239), .ZN(n8676) );
  INV_X1 U8011 ( .A(n8676), .ZN(n6297) );
  NAND2_X1 U8012 ( .A1(n6298), .A2(n6297), .ZN(n8671) );
  NAND2_X1 U8013 ( .A1(n7268), .A2(n6183), .ZN(n6303) );
  NAND2_X1 U8014 ( .A1(n4515), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6300) );
  INV_X1 U8015 ( .A(n8519), .ZN(n8533) );
  AOI22_X1 U8016 ( .A1(n6301), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6646), .B2(
        n8533), .ZN(n6302) );
  INV_X1 U8017 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10285) );
  NAND2_X1 U8018 ( .A1(n6305), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U8019 ( .A1(n6317), .A2(n6306), .ZN(n8666) );
  NAND2_X1 U8020 ( .A1(n6405), .A2(n8666), .ZN(n6313) );
  INV_X1 U8021 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n6307) );
  OR2_X1 U8022 ( .A1(n4430), .A2(n6307), .ZN(n6312) );
  INV_X1 U8023 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n10236) );
  OR2_X1 U8024 ( .A1(n4445), .A2(n10236), .ZN(n6311) );
  INV_X1 U8025 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6309) );
  OR2_X1 U8026 ( .A1(n4440), .A2(n6309), .ZN(n6310) );
  NOR2_X1 U8027 ( .A1(n8788), .A2(n8648), .ZN(n8245) );
  INV_X1 U8028 ( .A(n6453), .ZN(n8260) );
  NAND2_X1 U8029 ( .A1(n7321), .A2(n6183), .ZN(n6316) );
  OR2_X1 U8030 ( .A1(n8133), .A2(n6314), .ZN(n6315) );
  NAND2_X1 U8031 ( .A1(n6317), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6318) );
  NAND2_X1 U8032 ( .A1(n6327), .A2(n6318), .ZN(n8652) );
  NAND2_X1 U8033 ( .A1(n8652), .A2(n6405), .ZN(n6322) );
  INV_X1 U8034 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n10299) );
  OR2_X1 U8035 ( .A1(n4445), .A2(n10299), .ZN(n6321) );
  NAND2_X1 U8036 ( .A1(n4433), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U8037 ( .A1(n6407), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U8038 ( .A1(n7357), .A2(n6183), .ZN(n6324) );
  OR2_X1 U8039 ( .A1(n8133), .A2(n7361), .ZN(n6323) );
  INV_X1 U8040 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U8041 ( .A1(n6327), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6328) );
  NAND2_X1 U8042 ( .A1(n6334), .A2(n6328), .ZN(n8637) );
  NAND2_X1 U8043 ( .A1(n8637), .A2(n6405), .ZN(n6331) );
  AOI22_X1 U8044 ( .A1(n6365), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n4433), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U8045 ( .A1(n6407), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6329) );
  NAND2_X1 U8046 ( .A1(n8859), .A2(n8649), .ZN(n8146) );
  NAND2_X1 U8047 ( .A1(n8653), .A2(n8660), .ZN(n8625) );
  AND2_X1 U8048 ( .A1(n8146), .A2(n8625), .ZN(n8259) );
  NAND2_X1 U8049 ( .A1(n6332), .A2(n8254), .ZN(n8612) );
  OR2_X1 U8050 ( .A1(n8133), .A2(n10269), .ZN(n6333) );
  INV_X1 U8051 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n10129) );
  NAND2_X1 U8052 ( .A1(n6334), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U8053 ( .A1(n6341), .A2(n6335), .ZN(n8621) );
  NAND2_X1 U8054 ( .A1(n8621), .A2(n6405), .ZN(n6337) );
  AOI22_X1 U8055 ( .A1(n4433), .A2(P2_REG0_REG_22__SCAN_IN), .B1(n6407), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U8056 ( .A1(n6458), .A2(n6459), .ZN(n8258) );
  NAND2_X1 U8057 ( .A1(n8612), .A2(n8258), .ZN(n6338) );
  NAND2_X1 U8058 ( .A1(n7645), .A2(n6183), .ZN(n6340) );
  OR2_X1 U8059 ( .A1(n8133), .A2(n7648), .ZN(n6339) );
  NAND2_X1 U8060 ( .A1(n6341), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6342) );
  NAND2_X1 U8061 ( .A1(n6352), .A2(n6342), .ZN(n8608) );
  NAND2_X1 U8062 ( .A1(n8608), .A2(n6405), .ZN(n6347) );
  INV_X1 U8063 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8778) );
  NAND2_X1 U8064 ( .A1(n6407), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6344) );
  NAND2_X1 U8065 ( .A1(n4433), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6343) );
  OAI211_X1 U8066 ( .C1(n4445), .C2(n8778), .A(n6344), .B(n6343), .ZN(n6345)
         );
  INV_X1 U8067 ( .A(n6345), .ZN(n6346) );
  NOR2_X1 U8068 ( .A1(n6462), .A2(n8595), .ZN(n8266) );
  NAND2_X1 U8069 ( .A1(n6462), .A2(n8595), .ZN(n8299) );
  OAI21_X2 U8070 ( .B1(n8602), .B2(n8266), .A(n8299), .ZN(n8598) );
  NAND2_X1 U8071 ( .A1(n7703), .A2(n6183), .ZN(n6349) );
  OR2_X1 U8072 ( .A1(n8133), .A2(n10301), .ZN(n6348) );
  INV_X1 U8073 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6350) );
  NAND2_X1 U8074 ( .A1(n6352), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6353) );
  NAND2_X1 U8075 ( .A1(n6363), .A2(n6353), .ZN(n8596) );
  NAND2_X1 U8076 ( .A1(n8596), .A2(n6405), .ZN(n6358) );
  INV_X1 U8077 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8775) );
  NAND2_X1 U8078 ( .A1(n6407), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U8079 ( .A1(n4433), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6354) );
  OAI211_X1 U8080 ( .C1(n4445), .C2(n8775), .A(n6355), .B(n6354), .ZN(n6356)
         );
  INV_X1 U8081 ( .A(n6356), .ZN(n6357) );
  OR2_X1 U8082 ( .A1(n8843), .A2(n8583), .ZN(n8265) );
  NAND2_X1 U8083 ( .A1(n7728), .A2(n6183), .ZN(n6360) );
  OR2_X1 U8084 ( .A1(n8133), .A2(n10115), .ZN(n6359) );
  INV_X1 U8085 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6361) );
  NAND2_X1 U8086 ( .A1(n6363), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6364) );
  NAND2_X1 U8087 ( .A1(n6374), .A2(n6364), .ZN(n8586) );
  NAND2_X1 U8088 ( .A1(n8586), .A2(n6405), .ZN(n6371) );
  INV_X1 U8089 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6368) );
  NAND2_X1 U8090 ( .A1(n6365), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6367) );
  NAND2_X1 U8091 ( .A1(n4433), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6366) );
  OAI211_X1 U8092 ( .C1(n6368), .C2(n4439), .A(n6367), .B(n6366), .ZN(n6369)
         );
  INV_X1 U8093 ( .A(n6369), .ZN(n6370) );
  NAND2_X1 U8094 ( .A1(n8585), .A2(n8594), .ZN(n8268) );
  NAND2_X1 U8095 ( .A1(n7800), .A2(n6183), .ZN(n6373) );
  OR2_X1 U8096 ( .A1(n8133), .A2(n7826), .ZN(n6372) );
  NAND2_X1 U8097 ( .A1(n6374), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6375) );
  NAND2_X1 U8098 ( .A1(n6385), .A2(n6375), .ZN(n8575) );
  NAND2_X1 U8099 ( .A1(n8575), .A2(n6405), .ZN(n6380) );
  INV_X1 U8100 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8768) );
  NAND2_X1 U8101 ( .A1(n4433), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6377) );
  NAND2_X1 U8102 ( .A1(n6407), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6376) );
  OAI211_X1 U8103 ( .C1(n8768), .C2(n4445), .A(n6377), .B(n6376), .ZN(n6378)
         );
  INV_X1 U8104 ( .A(n6378), .ZN(n6379) );
  NAND2_X2 U8105 ( .A1(n6380), .A2(n6379), .ZN(n8565) );
  NOR2_X1 U8106 ( .A1(n8832), .A2(n8584), .ZN(n8271) );
  NAND2_X1 U8107 ( .A1(n7841), .A2(n6183), .ZN(n6382) );
  OR2_X1 U8108 ( .A1(n8133), .A2(n7848), .ZN(n6381) );
  INV_X1 U8109 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6383) );
  NAND2_X1 U8110 ( .A1(n6385), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U8111 ( .A1(n6394), .A2(n6386), .ZN(n8568) );
  NAND2_X1 U8112 ( .A1(n8568), .A2(n6405), .ZN(n6391) );
  INV_X1 U8113 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U8114 ( .A1(n6407), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U8115 ( .A1(n4433), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6387) );
  OAI211_X1 U8116 ( .C1(n4445), .C2(n8764), .A(n6388), .B(n6387), .ZN(n6389)
         );
  INV_X1 U8117 ( .A(n6389), .ZN(n6390) );
  NAND2_X1 U8118 ( .A1(n7849), .A2(n6183), .ZN(n6393) );
  INV_X1 U8119 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7846) );
  OR2_X1 U8120 ( .A1(n8133), .A2(n7846), .ZN(n6392) );
  NAND2_X1 U8121 ( .A1(n6394), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6395) );
  NAND2_X1 U8122 ( .A1(n7958), .A2(n6395), .ZN(n8557) );
  NAND2_X1 U8123 ( .A1(n8557), .A2(n6405), .ZN(n6400) );
  INV_X1 U8124 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8761) );
  NAND2_X1 U8125 ( .A1(n6407), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6397) );
  NAND2_X1 U8126 ( .A1(n4433), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6396) );
  OAI211_X1 U8127 ( .C1(n4445), .C2(n8761), .A(n6397), .B(n6396), .ZN(n6398)
         );
  INV_X1 U8128 ( .A(n6398), .ZN(n6399) );
  NAND2_X1 U8129 ( .A1(n8550), .A2(n8552), .ZN(n6402) );
  INV_X1 U8130 ( .A(n8564), .ZN(n7971) );
  OR2_X1 U8131 ( .A1(n8558), .A2(n7971), .ZN(n6401) );
  NAND2_X1 U8132 ( .A1(n7866), .A2(n6183), .ZN(n6404) );
  OR2_X1 U8133 ( .A1(n8133), .A2(n7965), .ZN(n6403) );
  INV_X1 U8134 ( .A(n7958), .ZN(n6406) );
  NAND2_X1 U8135 ( .A1(n6406), .A2(n6405), .ZN(n7217) );
  INV_X1 U8136 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6410) );
  NAND2_X1 U8137 ( .A1(n4433), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6409) );
  NAND2_X1 U8138 ( .A1(n6407), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6408) );
  OAI211_X1 U8139 ( .C1(n6410), .C2(n4445), .A(n6409), .B(n6408), .ZN(n6411)
         );
  INV_X1 U8140 ( .A(n6411), .ZN(n6412) );
  NAND2_X1 U8141 ( .A1(n6520), .A2(n8553), .ZN(n8140) );
  NAND2_X1 U8142 ( .A1(n4512), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6416) );
  INV_X1 U8143 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U8144 ( .A1(n6416), .A2(n6413), .ZN(n6418) );
  INV_X1 U8145 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6414) );
  INV_X1 U8146 ( .A(n6416), .ZN(n6417) );
  NAND2_X1 U8147 ( .A1(n6417), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n6419) );
  NAND2_X1 U8148 ( .A1(n8194), .A2(n8144), .ZN(n6963) );
  NAND2_X1 U8149 ( .A1(n6420), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6421) );
  XNOR2_X1 U8150 ( .A(n6421), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8337) );
  NAND2_X1 U8151 ( .A1(n6963), .A2(n7453), .ZN(n6422) );
  NAND2_X1 U8152 ( .A1(n6422), .A2(n8519), .ZN(n6526) );
  INV_X1 U8153 ( .A(n6526), .ZN(n6423) );
  NAND2_X1 U8154 ( .A1(n8144), .A2(n8519), .ZN(n6877) );
  OR2_X1 U8155 ( .A1(n8292), .A2(n6877), .ZN(n6929) );
  INV_X1 U8156 ( .A(n7688), .ZN(n10040) );
  NAND2_X1 U8157 ( .A1(n8354), .A2(n6075), .ZN(n6425) );
  OR2_X1 U8158 ( .A1(n8353), .A2(n6913), .ZN(n7108) );
  NAND2_X1 U8159 ( .A1(n6427), .A2(n6426), .ZN(n6954) );
  OR2_X1 U8160 ( .A1(n4442), .A2(n6887), .ZN(n6955) );
  INV_X1 U8161 ( .A(n7008), .ZN(n10011) );
  OR2_X1 U8162 ( .A1(n10011), .A2(n8351), .ZN(n7120) );
  INV_X1 U8163 ( .A(n7003), .ZN(n10016) );
  OR2_X1 U8164 ( .A1(n10016), .A2(n7998), .ZN(n6429) );
  NAND2_X1 U8165 ( .A1(n7119), .A2(n6429), .ZN(n7092) );
  INV_X1 U8166 ( .A(n8350), .ZN(n7056) );
  NAND2_X1 U8167 ( .A1(n8349), .A2(n10028), .ZN(n6431) );
  NAND2_X1 U8168 ( .A1(n7248), .A2(n6431), .ZN(n7441) );
  NAND2_X1 U8169 ( .A1(n8347), .A2(n7658), .ZN(n7649) );
  INV_X1 U8170 ( .A(n7649), .ZN(n6433) );
  OR2_X1 U8171 ( .A1(n8311), .A2(n6433), .ZN(n7676) );
  OR2_X1 U8172 ( .A1(n7676), .A2(n6182), .ZN(n6435) );
  INV_X1 U8173 ( .A(n7515), .ZN(n7518) );
  OR2_X1 U8174 ( .A1(n7518), .A2(n8348), .ZN(n7652) );
  OR2_X1 U8175 ( .A1(n8347), .A2(n7658), .ZN(n7650) );
  AND2_X1 U8176 ( .A1(n7652), .A2(n7650), .ZN(n6432) );
  OAI21_X1 U8177 ( .B1(n7441), .B2(n6435), .A(n6434), .ZN(n7681) );
  AOI21_X1 U8178 ( .B1(n10040), .B2(n7292), .A(n7681), .ZN(n6436) );
  INV_X1 U8179 ( .A(n6436), .ZN(n7634) );
  OAI21_X1 U8180 ( .B1(n7634), .B2(n7708), .A(n6437), .ZN(n6439) );
  NAND2_X1 U8181 ( .A1(n7634), .A2(n7708), .ZN(n6438) );
  NAND2_X1 U8182 ( .A1(n6439), .A2(n6438), .ZN(n7707) );
  AND2_X1 U8183 ( .A1(n10054), .A2(n8344), .ZN(n6440) );
  NAND2_X1 U8184 ( .A1(n6443), .A2(n8225), .ZN(n6445) );
  INV_X1 U8185 ( .A(n6442), .ZN(n6443) );
  NOR2_X1 U8186 ( .A1(n6443), .A2(n8225), .ZN(n6444) );
  AOI21_X1 U8187 ( .B1(n6445), .B2(n8317), .A(n6444), .ZN(n8725) );
  NAND2_X1 U8188 ( .A1(n8887), .A2(n8714), .ZN(n6447) );
  NOR2_X1 U8189 ( .A1(n8887), .A2(n8714), .ZN(n6446) );
  INV_X1 U8190 ( .A(n8803), .ZN(n8721) );
  NAND2_X1 U8191 ( .A1(n8721), .A2(n8302), .ZN(n6448) );
  INV_X1 U8192 ( .A(n8879), .ZN(n6450) );
  INV_X1 U8193 ( .A(n8795), .ZN(n8691) );
  NOR2_X1 U8194 ( .A1(n8691), .A2(n8033), .ZN(n6451) );
  NAND2_X1 U8195 ( .A1(n8246), .A2(n8625), .ZN(n8643) );
  INV_X1 U8196 ( .A(n8648), .ZN(n8678) );
  NAND2_X1 U8197 ( .A1(n8788), .A2(n8678), .ZN(n8644) );
  NOR2_X1 U8198 ( .A1(n8245), .A2(n6453), .ZN(n8657) );
  INV_X1 U8199 ( .A(n8659), .ZN(n8687) );
  NOR2_X1 U8200 ( .A1(n8872), .A2(n8687), .ZN(n8628) );
  OAI211_X1 U8201 ( .C1(n8657), .C2(n8628), .A(n8644), .B(n8643), .ZN(n6454)
         );
  INV_X1 U8202 ( .A(n8653), .ZN(n8865) );
  NAND2_X1 U8203 ( .A1(n8865), .A2(n8660), .ZN(n8630) );
  NAND2_X1 U8204 ( .A1(n6454), .A2(n8630), .ZN(n6455) );
  NAND2_X1 U8205 ( .A1(n8254), .A2(n8146), .ZN(n8629) );
  INV_X1 U8206 ( .A(n8859), .ZN(n8020) );
  NAND2_X1 U8207 ( .A1(n8020), .A2(n8649), .ZN(n8614) );
  NAND2_X1 U8208 ( .A1(n8613), .A2(n8614), .ZN(n6457) );
  NAND2_X1 U8209 ( .A1(n6460), .A2(n6459), .ZN(n6461) );
  NAND2_X1 U8210 ( .A1(n6462), .A2(n8618), .ZN(n6463) );
  INV_X1 U8211 ( .A(n8843), .ZN(n8060) );
  NAND2_X1 U8212 ( .A1(n8843), .A2(n8605), .ZN(n6464) );
  NAND2_X1 U8213 ( .A1(n6465), .A2(n6464), .ZN(n8581) );
  NAND2_X1 U8214 ( .A1(n8837), .A2(n8594), .ZN(n6466) );
  NOR2_X1 U8215 ( .A1(n8832), .A2(n8565), .ZN(n6467) );
  NAND2_X1 U8216 ( .A1(n8826), .A2(n8341), .ZN(n6469) );
  NOR2_X1 U8217 ( .A1(n8826), .A2(n8341), .ZN(n6468) );
  INV_X1 U8218 ( .A(n8558), .ZN(n8823) );
  NAND2_X1 U8219 ( .A1(n8823), .A2(n7971), .ZN(n6470) );
  OR2_X1 U8220 ( .A1(n8144), .A2(n7359), .ZN(n8137) );
  NAND2_X1 U8221 ( .A1(n8337), .A2(n8533), .ZN(n6509) );
  NAND2_X1 U8222 ( .A1(n6471), .A2(n8731), .ZN(n6481) );
  INV_X1 U8223 ( .A(n6472), .ZN(n8334) );
  NAND2_X1 U8224 ( .A1(n8334), .A2(n6650), .ZN(n6473) );
  NAND2_X1 U8225 ( .A1(n6074), .A2(n6473), .ZN(n6888) );
  INV_X1 U8226 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6476) );
  NAND2_X1 U8227 ( .A1(n4433), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6475) );
  INV_X1 U8228 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8549) );
  OR2_X1 U8229 ( .A1(n4440), .A2(n8549), .ZN(n6474) );
  OAI211_X1 U8230 ( .C1(n4445), .C2(n6476), .A(n6475), .B(n6474), .ZN(n6477)
         );
  INV_X1 U8231 ( .A(n6477), .ZN(n6478) );
  NAND2_X1 U8232 ( .A1(n7217), .A2(n6478), .ZN(n8340) );
  AND2_X1 U8233 ( .A1(n6074), .A2(P2_B_REG_SCAN_IN), .ZN(n6479) );
  NOR2_X1 U8234 ( .A1(n8744), .A2(n6479), .ZN(n8541) );
  AOI22_X1 U8235 ( .A1(n8726), .A2(n8564), .B1(n8340), .B2(n8541), .ZN(n6480)
         );
  NAND2_X1 U8236 ( .A1(n7453), .A2(n6770), .ZN(n10045) );
  NAND2_X1 U8237 ( .A1(n6507), .A2(n6508), .ZN(n6483) );
  NAND2_X1 U8238 ( .A1(n4514), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6486) );
  MUX2_X1 U8239 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6486), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6488) );
  NAND2_X1 U8240 ( .A1(n6489), .A2(n6491), .ZN(n6492) );
  NAND2_X1 U8241 ( .A1(n6490), .A2(n7828), .ZN(n6624) );
  NAND2_X1 U8242 ( .A1(n7758), .A2(n7828), .ZN(n6621) );
  NAND2_X1 U8243 ( .A1(n6493), .A2(n6621), .ZN(n6921) );
  INV_X1 U8244 ( .A(n6525), .ZN(n6504) );
  NOR4_X1 U8245 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6502) );
  INV_X1 U8246 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10295) );
  INV_X1 U8247 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10245) );
  INV_X1 U8248 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10114) );
  INV_X1 U8249 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10202) );
  NAND4_X1 U8250 ( .A1(n10295), .A2(n10245), .A3(n10114), .A4(n10202), .ZN(
        n6499) );
  NOR4_X1 U8251 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6497) );
  NOR4_X1 U8252 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6496) );
  NOR4_X1 U8253 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6495) );
  NOR4_X1 U8254 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6494) );
  NAND4_X1 U8255 ( .A1(n6497), .A2(n6496), .A3(n6495), .A4(n6494), .ZN(n6498)
         );
  NOR4_X1 U8256 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        n6499), .A4(n6498), .ZN(n6501) );
  NOR4_X1 U8257 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6500) );
  AND3_X1 U8258 ( .A1(n6502), .A2(n6501), .A3(n6500), .ZN(n6503) );
  OR2_X1 U8259 ( .A1(n6492), .A2(n6503), .ZN(n6523) );
  NAND2_X1 U8260 ( .A1(n6504), .A2(n6523), .ZN(n6771) );
  INV_X1 U8261 ( .A(n6771), .ZN(n6511) );
  NOR2_X1 U8262 ( .A1(n6490), .A2(n7828), .ZN(n6506) );
  INV_X1 U8263 ( .A(n7758), .ZN(n6505) );
  NAND2_X1 U8264 ( .A1(n6506), .A2(n6505), .ZN(n6757) );
  XNOR2_X1 U8265 ( .A(n6507), .B(n6508), .ZN(n6644) );
  NAND2_X1 U8266 ( .A1(n7359), .A2(n8280), .ZN(n8328) );
  OR2_X1 U8267 ( .A1(n8328), .A2(n6509), .ZN(n6764) );
  OR2_X1 U8268 ( .A1(n6928), .A2(n6929), .ZN(n6774) );
  OAI21_X1 U8269 ( .B1(n6928), .B2(n6764), .A(n6774), .ZN(n6510) );
  NAND2_X1 U8270 ( .A1(n6511), .A2(n6510), .ZN(n6516) );
  NAND3_X1 U8271 ( .A1(n6875), .A2(n6921), .A3(n6523), .ZN(n6775) );
  AND2_X1 U8272 ( .A1(n8292), .A2(n10039), .ZN(n6763) );
  NAND2_X1 U8273 ( .A1(n6763), .A2(n6764), .ZN(n6512) );
  OR2_X1 U8274 ( .A1(n10039), .A2(n6770), .ZN(n8747) );
  NAND2_X1 U8275 ( .A1(n6512), .A2(n8747), .ZN(n6754) );
  INV_X1 U8276 ( .A(n6754), .ZN(n6513) );
  OR2_X1 U8277 ( .A1(n6928), .A2(n6513), .ZN(n6514) );
  NAND2_X1 U8278 ( .A1(n10062), .A2(n6517), .ZN(n6518) );
  NAND2_X1 U8279 ( .A1(n6519), .A2(n6518), .ZN(n6521) );
  NAND2_X1 U8280 ( .A1(n6521), .A2(n5061), .ZN(P2_U3456) );
  INV_X1 U8281 ( .A(n6928), .ZN(n6766) );
  INV_X1 U8282 ( .A(n6877), .ZN(n6522) );
  OR2_X1 U8283 ( .A1(n8292), .A2(n6522), .ZN(n6756) );
  AND3_X1 U8284 ( .A1(n6523), .A2(n6766), .A3(n6756), .ZN(n6524) );
  AND2_X1 U8285 ( .A1(n6525), .A2(n6524), .ZN(n6925) );
  NOR2_X1 U8286 ( .A1(n10045), .A2(n8194), .ZN(n6528) );
  OR2_X1 U8287 ( .A1(n6526), .A2(n8144), .ZN(n6527) );
  AND2_X1 U8288 ( .A1(n6527), .A2(n8292), .ZN(n6920) );
  OAI21_X1 U8289 ( .B1(n6875), .B2(n6528), .A(n6920), .ZN(n6530) );
  INV_X1 U8290 ( .A(n6920), .ZN(n6919) );
  NAND2_X1 U8291 ( .A1(n6921), .A2(n6919), .ZN(n6529) );
  NAND2_X1 U8292 ( .A1(n6533), .A2(n6410), .ZN(n6534) );
  NAND2_X1 U8293 ( .A1(n6535), .A2(n6534), .ZN(n6536) );
  NAND2_X1 U8294 ( .A1(n10075), .A2(n10061), .ZN(n8785) );
  NAND2_X1 U8295 ( .A1(n6536), .A2(n5063), .ZN(P2_U3488) );
  INV_X1 U8296 ( .A(n6537), .ZN(n6538) );
  INV_X1 U8297 ( .A(n6625), .ZN(n6762) );
  OR2_X2 U8298 ( .A1(n6757), .A2(n6762), .ZN(n8497) );
  OAI21_X1 U8299 ( .B1(n6542), .B2(n6541), .A(n6540), .ZN(n6543) );
  AND2_X1 U8300 ( .A1(n6543), .A2(n9031), .ZN(n6548) );
  NAND2_X1 U8301 ( .A1(n9048), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6838) );
  AND2_X1 U8302 ( .A1(n6838), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6547) );
  INV_X1 U8303 ( .A(n4429), .ZN(n6940) );
  NOR2_X1 U8304 ( .A1(n9043), .A2(n6940), .ZN(n6546) );
  INV_X1 U8305 ( .A(n9325), .ZN(n6544) );
  OAI22_X1 U8306 ( .A1(n6544), .A2(n8983), .B1(n9039), .B2(n9237), .ZN(n6545)
         );
  OR4_X1 U8307 ( .A1(n6548), .A2(n6547), .A3(n6546), .A4(n6545), .ZN(P1_U3222)
         );
  AND2_X1 U8308 ( .A1(n4436), .A2(P1_U3086), .ZN(n9764) );
  OAI222_X1 U8309 ( .A1(n9771), .A2(n6551), .B1(n9769), .B2(n6558), .C1(
        P1_U3086), .C2(n6607), .ZN(P1_U3354) );
  OAI222_X1 U8310 ( .A1(n9353), .A2(P1_U3086), .B1(n9769), .B2(n6568), .C1(
        n9771), .C2(n5167), .ZN(P1_U3351) );
  OAI222_X1 U8311 ( .A1(n9771), .A2(n6552), .B1(n9769), .B2(n6556), .C1(
        P1_U3086), .C2(n9340), .ZN(P1_U3352) );
  OAI222_X1 U8312 ( .A1(n9771), .A2(n6553), .B1(n9769), .B2(n6554), .C1(
        P1_U3086), .C2(n6822), .ZN(P1_U3353) );
  AND2_X1 U8313 ( .A1(n4436), .A2(P2_U3151), .ZN(n6575) );
  INV_X2 U8314 ( .A(n6575), .ZN(n8899) );
  NOR2_X1 U8315 ( .A1(n4436), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8897) );
  INV_X2 U8316 ( .A(n8897), .ZN(n8900) );
  OAI222_X1 U8317 ( .A1(n8899), .A2(n6555), .B1(n8900), .B2(n6554), .C1(
        P2_U3151), .C2(n6737), .ZN(P2_U3293) );
  INV_X1 U8318 ( .A(n6782), .ZN(n6739) );
  OAI222_X1 U8319 ( .A1(n8899), .A2(n6557), .B1(n8900), .B2(n6556), .C1(
        P2_U3151), .C2(n6739), .ZN(P2_U3292) );
  OAI222_X1 U8320 ( .A1(n9995), .A2(P2_U3151), .B1(n8900), .B2(n6558), .C1(
        n5100), .C2(n8899), .ZN(P2_U3294) );
  OAI222_X1 U8321 ( .A1(n9771), .A2(n6559), .B1(n9769), .B2(n6560), .C1(
        P1_U3086), .C2(n9366), .ZN(P1_U3350) );
  OAI222_X1 U8322 ( .A1(n8899), .A2(n6561), .B1(n8900), .B2(n6560), .C1(
        P2_U3151), .C2(n6861), .ZN(P2_U3290) );
  OAI222_X1 U8323 ( .A1(n8899), .A2(n6562), .B1(n8900), .B2(n6563), .C1(
        P2_U3151), .C2(n7075), .ZN(P2_U3289) );
  INV_X1 U8324 ( .A(n6629), .ZN(n6632) );
  OAI222_X1 U8325 ( .A1(n9771), .A2(n6564), .B1(n9769), .B2(n6563), .C1(
        P1_U3086), .C2(n6632), .ZN(P1_U3349) );
  OAI222_X1 U8326 ( .A1(n8899), .A2(n6565), .B1(n8900), .B2(n6566), .C1(
        P2_U3151), .C2(n7180), .ZN(P2_U3288) );
  INV_X1 U8327 ( .A(n6676), .ZN(n6640) );
  OAI222_X1 U8328 ( .A1(n9771), .A2(n6567), .B1(n9769), .B2(n6566), .C1(
        P1_U3086), .C2(n6640), .ZN(P1_U3348) );
  INV_X1 U8329 ( .A(n6852), .ZN(n6849) );
  OAI222_X1 U8330 ( .A1(n8899), .A2(n6569), .B1(n8900), .B2(n6568), .C1(
        P2_U3151), .C2(n6849), .ZN(P2_U3291) );
  INV_X1 U8331 ( .A(n6570), .ZN(n6572) );
  INV_X1 U8332 ( .A(n9771), .ZN(n7053) );
  AOI22_X1 U8333 ( .A1(n6703), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n7053), .ZN(n6571) );
  OAI21_X1 U8334 ( .B1(n6572), .B2(n9769), .A(n6571), .ZN(P1_U3347) );
  NOR2_X1 U8335 ( .A1(n6620), .A2(n10295), .ZN(P2_U3242) );
  NOR2_X1 U8336 ( .A1(n6620), .A2(n10114), .ZN(P2_U3255) );
  NOR2_X1 U8337 ( .A1(n6620), .A2(n10202), .ZN(P2_U3252) );
  NOR2_X1 U8338 ( .A1(n6620), .A2(n10245), .ZN(P2_U3260) );
  OAI222_X1 U8339 ( .A1(n8899), .A2(n6573), .B1(n8900), .B2(n6572), .C1(
        P2_U3151), .C2(n7402), .ZN(P2_U3287) );
  INV_X1 U8340 ( .A(n6574), .ZN(n6577) );
  AOI22_X1 U8341 ( .A1(n7427), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n6575), .ZN(n6576) );
  OAI21_X1 U8342 ( .B1(n6577), .B2(n8900), .A(n6576), .ZN(P2_U3286) );
  INV_X1 U8343 ( .A(n6866), .ZN(n6709) );
  OAI222_X1 U8344 ( .A1(n9769), .A2(n6577), .B1(n6709), .B2(P1_U3086), .C1(
        n10178), .C2(n9771), .ZN(P1_U3346) );
  INV_X1 U8345 ( .A(n6578), .ZN(n6595) );
  AOI22_X1 U8346 ( .A1(n7029), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n7053), .ZN(n6579) );
  OAI21_X1 U8347 ( .B1(n6595), .B2(n9769), .A(n6579), .ZN(P1_U3345) );
  AND2_X1 U8348 ( .A1(n6580), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8349 ( .A1(n6580), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8350 ( .A1(n6580), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8351 ( .A1(n6580), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8352 ( .A1(n6580), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8353 ( .A1(n6580), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8354 ( .A1(n6580), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8355 ( .A1(n6580), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8356 ( .A1(n6580), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8357 ( .A1(n6580), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8358 ( .A1(n6580), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  INV_X1 U8359 ( .A(n7843), .ZN(n6812) );
  AOI21_X1 U8360 ( .B1(n6812), .B2(n6581), .A(n4443), .ZN(n6818) );
  OAI21_X1 U8361 ( .B1(n6812), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6818), .ZN(
        n6582) );
  MUX2_X1 U8362 ( .A(n6818), .B(n6582), .S(n9333), .Z(n6594) );
  NAND2_X1 U8363 ( .A1(n9076), .A2(n6585), .ZN(n6583) );
  AND2_X1 U8364 ( .A1(n6584), .A2(n6583), .ZN(n6588) );
  INV_X1 U8365 ( .A(n6585), .ZN(n6586) );
  NAND2_X1 U8366 ( .A1(n6586), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9308) );
  NAND2_X1 U8367 ( .A1(n9304), .A2(n9308), .ZN(n6587) );
  NAND2_X1 U8368 ( .A1(n6588), .A2(n6587), .ZN(n6604) );
  NAND3_X1 U8369 ( .A1(n9443), .A2(P1_IR_REG_0__SCAN_IN), .A3(n5771), .ZN(
        n6593) );
  INV_X1 U8370 ( .A(n6587), .ZN(n6589) );
  OR2_X1 U8371 ( .A1(n6589), .A2(n6588), .ZN(n9455) );
  INV_X1 U8372 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6590) );
  OAI22_X1 U8373 ( .A1(n9455), .A2(n6590), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7134), .ZN(n6591) );
  INV_X1 U8374 ( .A(n6591), .ZN(n6592) );
  OAI211_X1 U8375 ( .C1(n6594), .C2(n6604), .A(n6593), .B(n6592), .ZN(P1_U3243) );
  INV_X1 U8376 ( .A(n7431), .ZN(n7532) );
  OAI222_X1 U8377 ( .A1(n8899), .A2(n10249), .B1(n8900), .B2(n6595), .C1(n7532), .C2(P2_U3151), .ZN(P2_U3285) );
  INV_X1 U8378 ( .A(n6607), .ZN(n9332) );
  NAND2_X1 U8379 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9328) );
  NOR2_X1 U8380 ( .A1(n9327), .A2(n9328), .ZN(n9326) );
  INV_X1 U8381 ( .A(n6822), .ZN(n6609) );
  XNOR2_X1 U8382 ( .A(n6609), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6824) );
  NOR2_X1 U8383 ( .A1(n6825), .A2(n6824), .ZN(n6823) );
  INV_X1 U8384 ( .A(n6823), .ZN(n6596) );
  OAI21_X1 U8385 ( .B1(n6597), .B2(n6822), .A(n6596), .ZN(n9344) );
  XNOR2_X1 U8386 ( .A(n9340), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9345) );
  NAND2_X1 U8387 ( .A1(n9344), .A2(n9345), .ZN(n9343) );
  OAI21_X1 U8388 ( .B1(n6598), .B2(n9340), .A(n9343), .ZN(n9357) );
  MUX2_X1 U8389 ( .A(n6599), .B(P1_REG2_REG_4__SCAN_IN), .S(n9353), .Z(n9358)
         );
  NAND2_X1 U8390 ( .A1(n9357), .A2(n9358), .ZN(n9356) );
  XNOR2_X1 U8391 ( .A(n9366), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n9370) );
  OAI21_X1 U8392 ( .B1(n6600), .B2(n9366), .A(n9369), .ZN(n6602) );
  MUX2_X1 U8393 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7225), .S(n6629), .Z(n6601)
         );
  NAND2_X1 U8394 ( .A1(n6815), .A2(n6812), .ZN(n9305) );
  INV_X1 U8395 ( .A(n9428), .ZN(n9450) );
  OAI21_X1 U8396 ( .B1(n6602), .B2(n6601), .A(n9450), .ZN(n6619) );
  AND2_X1 U8397 ( .A1(n6602), .A2(n6601), .ZN(n6628) );
  INV_X1 U8398 ( .A(n9455), .ZN(n9433) );
  NOR2_X1 U8399 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6603), .ZN(n7261) );
  NOR2_X1 U8400 ( .A1(n9445), .A2(n6632), .ZN(n6605) );
  AOI211_X1 U8401 ( .C1(n9433), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n7261), .B(
        n6605), .ZN(n6618) );
  INV_X1 U8402 ( .A(n9340), .ZN(n6610) );
  MUX2_X1 U8403 ( .A(n6606), .B(P1_REG1_REG_2__SCAN_IN), .S(n6822), .Z(n6819)
         );
  XNOR2_X1 U8404 ( .A(n6607), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9336) );
  NAND3_X1 U8405 ( .A1(n9336), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9334) );
  OAI21_X1 U8406 ( .B1(n6608), .B2(n6607), .A(n9334), .ZN(n6820) );
  AOI22_X1 U8407 ( .A1(n6819), .A2(n6820), .B1(n6609), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n9348) );
  MUX2_X1 U8408 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n5136), .S(n9340), .Z(n9347)
         );
  NOR2_X1 U8409 ( .A1(n9348), .A2(n9347), .ZN(n9346) );
  AOI21_X1 U8410 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n6610), .A(n9346), .ZN(
        n9359) );
  MUX2_X1 U8411 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n5155), .S(n9353), .Z(n9360)
         );
  OAI22_X1 U8412 ( .A1(n9359), .A2(n9360), .B1(n5155), .B2(n9353), .ZN(n9373)
         );
  MUX2_X1 U8413 ( .A(n6611), .B(P1_REG1_REG_5__SCAN_IN), .S(n9366), .Z(n9374)
         );
  NAND2_X1 U8414 ( .A1(n9373), .A2(n9374), .ZN(n9372) );
  INV_X1 U8415 ( .A(n9366), .ZN(n6612) );
  NAND2_X1 U8416 ( .A1(n6612), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6614) );
  INV_X1 U8417 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9972) );
  MUX2_X1 U8418 ( .A(n9972), .B(P1_REG1_REG_6__SCAN_IN), .S(n6629), .Z(n6613)
         );
  AOI21_X1 U8419 ( .B1(n9372), .B2(n6614), .A(n6613), .ZN(n6636) );
  INV_X1 U8420 ( .A(n6636), .ZN(n6616) );
  NAND3_X1 U8421 ( .A1(n9372), .A2(n6614), .A3(n6613), .ZN(n6615) );
  NAND3_X1 U8422 ( .A1(n6616), .A2(n9443), .A3(n6615), .ZN(n6617) );
  OAI211_X1 U8423 ( .C1(n6619), .C2(n6628), .A(n6618), .B(n6617), .ZN(P1_U3249) );
  INV_X1 U8424 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6623) );
  INV_X1 U8425 ( .A(n6621), .ZN(n6622) );
  AOI22_X1 U8426 ( .A1(n6580), .A2(n6623), .B1(n6622), .B2(n6625), .ZN(
        P2_U3377) );
  INV_X1 U8427 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6627) );
  INV_X1 U8428 ( .A(n6624), .ZN(n6626) );
  AOI22_X1 U8429 ( .A1(n6580), .A2(n6627), .B1(n6626), .B2(n6625), .ZN(
        P2_U3376) );
  NOR2_X1 U8430 ( .A1(n9433), .A2(n9324), .ZN(P1_U3085) );
  XNOR2_X1 U8431 ( .A(n6676), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n6630) );
  NOR2_X1 U8432 ( .A1(n6631), .A2(n6630), .ZN(n6673) );
  AOI211_X1 U8433 ( .C1(n6631), .C2(n6630), .A(n9428), .B(n6673), .ZN(n6643)
         );
  NOR2_X1 U8434 ( .A1(n6632), .A2(n9972), .ZN(n6635) );
  MUX2_X1 U8435 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6633), .S(n6676), .Z(n6634)
         );
  OAI21_X1 U8436 ( .B1(n6636), .B2(n6635), .A(n6634), .ZN(n6679) );
  INV_X1 U8437 ( .A(n6679), .ZN(n6638) );
  NOR3_X1 U8438 ( .A1(n6636), .A2(n6635), .A3(n6634), .ZN(n6637) );
  NOR3_X1 U8439 ( .A1(n6638), .A2(n6637), .A3(n9446), .ZN(n6642) );
  NOR2_X1 U8440 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5226), .ZN(n7352) );
  AOI21_X1 U8441 ( .B1(n9433), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n7352), .ZN(
        n6639) );
  OAI21_X1 U8442 ( .B1(n6640), .B2(n9445), .A(n6639), .ZN(n6641) );
  OR3_X1 U8443 ( .A1(n6643), .A2(n6642), .A3(n6641), .ZN(P1_U3250) );
  AND2_X1 U8444 ( .A1(n6580), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8445 ( .A1(n6580), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8446 ( .A1(n6580), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8447 ( .A1(n6580), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8448 ( .A1(n6580), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8449 ( .A1(n6580), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8450 ( .A1(n6580), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8451 ( .A1(n6580), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8452 ( .A1(n6580), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8453 ( .A1(n6580), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8454 ( .A1(n6580), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8455 ( .A1(n6580), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8456 ( .A1(n6580), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8457 ( .A1(n6580), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8458 ( .A1(n6580), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  INV_X1 U8459 ( .A(n6644), .ZN(n7016) );
  OR2_X1 U8460 ( .A1(n6757), .A2(n7016), .ZN(n6649) );
  NAND2_X1 U8461 ( .A1(n8274), .A2(n6644), .ZN(n6645) );
  NAND2_X1 U8462 ( .A1(n6649), .A2(n6645), .ZN(n6654) );
  OR2_X1 U8463 ( .A1(n6654), .A2(n6646), .ZN(n6647) );
  NAND2_X1 U8464 ( .A1(n6647), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8465 ( .A(P2_U3150), .ZN(n6648) );
  NAND2_X1 U8466 ( .A1(n6648), .A2(n6649), .ZN(n10005) );
  INV_X1 U8467 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6661) );
  INV_X1 U8468 ( .A(n6649), .ZN(n6652) );
  NOR2_X1 U8469 ( .A1(n6654), .A2(n4446), .ZN(n6651) );
  MUX2_X1 U8470 ( .A(n6652), .B(n6651), .S(n6472), .Z(n6653) );
  NAND2_X1 U8472 ( .A1(n10411), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6660) );
  OR2_X1 U8473 ( .A1(n6472), .A2(P2_U3151), .ZN(n7844) );
  NAND2_X1 U8474 ( .A1(n6731), .A2(n8535), .ZN(n6658) );
  MUX2_X1 U8475 ( .A(n6934), .B(n6655), .S(n4438), .Z(n6656) );
  NAND2_X1 U8476 ( .A1(n6656), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9991) );
  OAI21_X1 U8477 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6656), .A(n9991), .ZN(n6657) );
  AOI22_X1 U8478 ( .A1(n6658), .A2(n6657), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n6659) );
  OAI211_X1 U8479 ( .C1(n10005), .C2(n6661), .A(n6660), .B(n6659), .ZN(
        P2_U3182) );
  INV_X1 U8480 ( .A(n6662), .ZN(n6688) );
  AOI22_X1 U8481 ( .A1(n7237), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n7053), .ZN(n6663) );
  OAI21_X1 U8482 ( .B1(n6688), .B2(n9769), .A(n6663), .ZN(P1_U3344) );
  INV_X1 U8483 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7269) );
  NAND2_X1 U8484 ( .A1(n9699), .A2(n9324), .ZN(n6664) );
  OAI21_X1 U8485 ( .B1(n7269), .B2(n9324), .A(n6664), .ZN(P1_U3573) );
  INV_X1 U8486 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6969) );
  NAND2_X1 U8487 ( .A1(n7742), .A2(n9324), .ZN(n6665) );
  OAI21_X1 U8488 ( .B1(n6969), .B2(n9324), .A(n6665), .ZN(P1_U3570) );
  NAND2_X1 U8489 ( .A1(n9583), .A2(n9324), .ZN(n6666) );
  OAI21_X1 U8490 ( .B1(n6314), .B2(n9324), .A(n6666), .ZN(P1_U3574) );
  INV_X1 U8491 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6672) );
  INV_X1 U8492 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9631) );
  NAND2_X1 U8493 ( .A1(n6667), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U8494 ( .A1(n4437), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6668) );
  OAI211_X1 U8495 ( .C1(n6670), .C2(n9631), .A(n6669), .B(n6668), .ZN(n9459)
         );
  NAND2_X1 U8496 ( .A1(n9459), .A2(n9324), .ZN(n6671) );
  OAI21_X1 U8497 ( .B1(n9324), .B2(n6672), .A(n6671), .ZN(P1_U3585) );
  AOI21_X1 U8498 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6676), .A(n6673), .ZN(
        n6675) );
  XNOR2_X1 U8499 ( .A(n6703), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6674) );
  NOR2_X1 U8500 ( .A1(n6675), .A2(n6674), .ZN(n6699) );
  AOI211_X1 U8501 ( .C1(n6675), .C2(n6674), .A(n9428), .B(n6699), .ZN(n6686)
         );
  NAND2_X1 U8502 ( .A1(n6676), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6678) );
  MUX2_X1 U8503 ( .A(n5256), .B(P1_REG1_REG_8__SCAN_IN), .S(n6703), .Z(n6677)
         );
  AOI21_X1 U8504 ( .B1(n6679), .B2(n6678), .A(n6677), .ZN(n6702) );
  AND3_X1 U8505 ( .A1(n6679), .A2(n6678), .A3(n6677), .ZN(n6680) );
  NOR3_X1 U8506 ( .A1(n6702), .A2(n6680), .A3(n9446), .ZN(n6685) );
  INV_X1 U8507 ( .A(n6703), .ZN(n6683) );
  NOR2_X1 U8508 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6681), .ZN(n7624) );
  AOI21_X1 U8509 ( .B1(n9433), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n7624), .ZN(
        n6682) );
  OAI21_X1 U8510 ( .B1(n6683), .B2(n9445), .A(n6682), .ZN(n6684) );
  OR3_X1 U8511 ( .A1(n6686), .A2(n6685), .A3(n6684), .ZN(P1_U3251) );
  NAND2_X1 U8512 ( .A1(n7998), .A2(P2_U3893), .ZN(n6687) );
  OAI21_X1 U8513 ( .B1(P2_U3893), .B2(n5167), .A(n6687), .ZN(P2_U3495) );
  INV_X1 U8514 ( .A(n7581), .ZN(n7571) );
  OAI222_X1 U8515 ( .A1(n8899), .A2(n6689), .B1(n8900), .B2(n6688), .C1(
        P2_U3151), .C2(n7571), .ZN(P2_U3284) );
  OAI21_X1 U8516 ( .B1(n6692), .B2(n6691), .A(n6690), .ZN(n6814) );
  AOI22_X1 U8517 ( .A1(n6693), .A2(n9050), .B1(n9036), .B2(n9323), .ZN(n6695)
         );
  NAND2_X1 U8518 ( .A1(n6838), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6694) );
  OAI211_X1 U8519 ( .C1(n6814), .C2(n9052), .A(n6695), .B(n6694), .ZN(P1_U3232) );
  INV_X1 U8520 ( .A(n6696), .ZN(n6750) );
  AOI22_X1 U8521 ( .A1(n7275), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n7053), .ZN(n6697) );
  OAI21_X1 U8522 ( .B1(n6750), .B2(n9769), .A(n6697), .ZN(P1_U3343) );
  XNOR2_X1 U8523 ( .A(n6866), .B(n6698), .ZN(n6701) );
  NAND2_X1 U8524 ( .A1(n6700), .A2(n6701), .ZN(n6862) );
  OAI21_X1 U8525 ( .B1(n6701), .B2(n6700), .A(n6862), .ZN(n6711) );
  MUX2_X1 U8526 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n5281), .S(n6866), .Z(n6705)
         );
  AOI21_X1 U8527 ( .B1(n6703), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6702), .ZN(
        n6704) );
  NAND2_X1 U8528 ( .A1(n6704), .A2(n6705), .ZN(n6865) );
  OAI21_X1 U8529 ( .B1(n6705), .B2(n6704), .A(n6865), .ZN(n6706) );
  NAND2_X1 U8530 ( .A1(n6706), .A2(n9443), .ZN(n6708) );
  AND2_X1 U8531 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7696) );
  AOI21_X1 U8532 ( .B1(n9433), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7696), .ZN(
        n6707) );
  OAI211_X1 U8533 ( .C1(n9445), .C2(n6709), .A(n6708), .B(n6707), .ZN(n6710)
         );
  AOI21_X1 U8534 ( .B1(n6711), .B2(n9450), .A(n6710), .ZN(n6712) );
  INV_X1 U8535 ( .A(n6712), .ZN(P1_U3252) );
  MUX2_X1 U8536 ( .A(n6714), .B(n6713), .S(n4438), .Z(n6781) );
  XNOR2_X1 U8537 ( .A(n6781), .B(n6782), .ZN(n6723) );
  INV_X1 U8538 ( .A(n6737), .ZN(n10410) );
  MUX2_X1 U8539 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n4438), .Z(n6720) );
  INV_X1 U8540 ( .A(n6720), .ZN(n6721) );
  INV_X1 U8541 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6716) );
  INV_X1 U8542 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6715) );
  MUX2_X1 U8543 ( .A(n6716), .B(n6715), .S(n4438), .Z(n6717) );
  NAND2_X1 U8544 ( .A1(n9992), .A2(n9991), .ZN(n9990) );
  INV_X1 U8545 ( .A(n6717), .ZN(n6718) );
  NAND2_X1 U8546 ( .A1(n6718), .A2(n9995), .ZN(n6719) );
  NAND2_X1 U8547 ( .A1(n9990), .A2(n6719), .ZN(n10409) );
  XNOR2_X1 U8548 ( .A(n6720), .B(n10410), .ZN(n10408) );
  NAND2_X1 U8549 ( .A1(n10409), .A2(n10408), .ZN(n10407) );
  OAI21_X1 U8550 ( .B1(n10410), .B2(n6721), .A(n10407), .ZN(n6722) );
  NOR2_X1 U8551 ( .A1(n6722), .A2(n6723), .ZN(n6780) );
  AOI21_X1 U8552 ( .B1(n6723), .B2(n6722), .A(n6780), .ZN(n6749) );
  INV_X1 U8553 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6746) );
  NOR2_X1 U8554 ( .A1(n6731), .A2(n4446), .ZN(n10419) );
  AND2_X1 U8555 ( .A1(n6733), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6724) );
  NAND2_X1 U8556 ( .A1(n6734), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6725) );
  OAI21_X1 U8557 ( .B1(n9995), .B2(n6724), .A(n6725), .ZN(n10000) );
  OR2_X1 U8558 ( .A1(n10000), .A2(n6716), .ZN(n9998) );
  NAND2_X1 U8559 ( .A1(n9998), .A2(n6725), .ZN(n10416) );
  NAND2_X1 U8560 ( .A1(n6737), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6726) );
  OAI21_X1 U8561 ( .B1(n6729), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6788), .ZN(
        n6730) );
  AND2_X1 U8562 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7997) );
  AOI21_X1 U8563 ( .B1(n10419), .B2(n6730), .A(n7997), .ZN(n6745) );
  INV_X1 U8564 ( .A(n6731), .ZN(n6732) );
  NAND2_X1 U8565 ( .A1(n6732), .A2(n4446), .ZN(n9985) );
  INV_X1 U8566 ( .A(n9985), .ZN(n10404) );
  AND2_X1 U8567 ( .A1(n6733), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6735) );
  NAND2_X1 U8568 ( .A1(n6734), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6736) );
  OAI21_X1 U8569 ( .B1(n9995), .B2(n6735), .A(n6736), .ZN(n9984) );
  NAND2_X1 U8570 ( .A1(n10402), .A2(n10401), .ZN(n10400) );
  NAND2_X1 U8571 ( .A1(n6737), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6738) );
  NAND2_X1 U8572 ( .A1(n10400), .A2(n6738), .ZN(n6740) );
  NAND2_X1 U8573 ( .A1(n6740), .A2(n6739), .ZN(n6791) );
  OR2_X1 U8574 ( .A1(n6740), .A2(n6739), .ZN(n6741) );
  AND2_X1 U8575 ( .A1(n6791), .A2(n6741), .ZN(n6742) );
  OAI21_X1 U8576 ( .B1(n6742), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6793), .ZN(
        n6743) );
  NAND2_X1 U8577 ( .A1(n10404), .A2(n6743), .ZN(n6744) );
  OAI211_X1 U8578 ( .C1(n6746), .C2(n10005), .A(n6745), .B(n6744), .ZN(n6747)
         );
  AOI21_X1 U8579 ( .B1(n6782), .B2(n10411), .A(n6747), .ZN(n6748) );
  OAI21_X1 U8580 ( .B1(n6749), .B2(n8535), .A(n6748), .ZN(P2_U3185) );
  OAI222_X1 U8581 ( .A1(n8899), .A2(n6751), .B1(n8900), .B2(n6750), .C1(n8373), 
        .C2(P2_U3151), .ZN(P2_U3283) );
  INV_X1 U8582 ( .A(n6752), .ZN(n6800) );
  AOI22_X1 U8583 ( .A1(n7363), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n7053), .ZN(n6753) );
  OAI21_X1 U8584 ( .B1(n6800), .B2(n9769), .A(n6753), .ZN(P1_U3342) );
  NAND2_X1 U8585 ( .A1(n6771), .A2(n6754), .ZN(n6758) );
  INV_X1 U8586 ( .A(n6764), .ZN(n6755) );
  NAND2_X1 U8587 ( .A1(n6775), .A2(n6755), .ZN(n6767) );
  NAND4_X1 U8588 ( .A1(n6758), .A2(n6757), .A3(n6767), .A4(n6756), .ZN(n6759)
         );
  NAND2_X1 U8589 ( .A1(n6759), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6761) );
  INV_X1 U8590 ( .A(n6774), .ZN(n8335) );
  NAND2_X1 U8591 ( .A1(n6775), .A2(n8335), .ZN(n6760) );
  NAND2_X1 U8592 ( .A1(n6761), .A2(n6760), .ZN(n7017) );
  NOR2_X1 U8593 ( .A1(n7017), .A2(n6762), .ZN(n6897) );
  INV_X1 U8594 ( .A(n6763), .ZN(n6765) );
  OAI21_X1 U8595 ( .B1(n6771), .B2(n6765), .A(n6764), .ZN(n6769) );
  AND2_X1 U8596 ( .A1(n6767), .A2(n6766), .ZN(n6768) );
  NAND2_X1 U8597 ( .A1(n8354), .A2(n6936), .ZN(n8187) );
  NAND2_X1 U8598 ( .A1(n6881), .A2(n8187), .ZN(n8305) );
  INV_X1 U8599 ( .A(n6770), .ZN(n6927) );
  NAND2_X1 U8600 ( .A1(n6771), .A2(n6927), .ZN(n6773) );
  NOR2_X1 U8601 ( .A1(n6928), .A2(n10039), .ZN(n6772) );
  OR2_X1 U8602 ( .A1(n6775), .A2(n6774), .ZN(n6889) );
  INV_X1 U8603 ( .A(n6889), .ZN(n6776) );
  NAND2_X1 U8604 ( .A1(n6776), .A2(n6888), .ZN(n8110) );
  OAI22_X1 U8605 ( .A1(n8116), .A2(n6936), .B1(n6883), .B2(n8110), .ZN(n6777)
         );
  AOI21_X1 U8606 ( .B1(n8104), .B2(n8305), .A(n6777), .ZN(n6778) );
  OAI21_X1 U8607 ( .B1(n6897), .B2(n6779), .A(n6778), .ZN(P2_U3172) );
  INV_X1 U8608 ( .A(n10411), .ZN(n9996) );
  MUX2_X1 U8609 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n4438), .Z(n6841) );
  XNOR2_X1 U8610 ( .A(n6841), .B(n6852), .ZN(n6783) );
  OAI211_X1 U8611 ( .C1(n6784), .C2(n6783), .A(n6842), .B(n10406), .ZN(n6799)
         );
  INV_X1 U8612 ( .A(n10005), .ZN(n10405) );
  MUX2_X1 U8613 ( .A(n7123), .B(P2_REG2_REG_4__SCAN_IN), .S(n6852), .Z(n6786)
         );
  NOR2_X1 U8614 ( .A1(n4903), .A2(n6786), .ZN(n6789) );
  INV_X1 U8615 ( .A(n6853), .ZN(n6787) );
  AOI21_X1 U8616 ( .B1(n6789), .B2(n6788), .A(n6787), .ZN(n6796) );
  INV_X1 U8617 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6790) );
  AND3_X1 U8618 ( .A1(n6793), .A2(n6792), .A3(n6791), .ZN(n6794) );
  OAI21_X1 U8619 ( .B1(n6848), .B2(n6794), .A(n10404), .ZN(n6795) );
  NAND2_X1 U8620 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7018) );
  OAI211_X1 U8621 ( .C1(n10002), .C2(n6796), .A(n6795), .B(n7018), .ZN(n6797)
         );
  AOI21_X1 U8622 ( .B1(n10405), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n6797), .ZN(
        n6798) );
  OAI211_X1 U8623 ( .C1(n9996), .C2(n6849), .A(n6799), .B(n6798), .ZN(P2_U3186) );
  INV_X1 U8624 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10164) );
  INV_X1 U8625 ( .A(n8397), .ZN(n8374) );
  OAI222_X1 U8626 ( .A1(n8899), .A2(n10164), .B1(n8900), .B2(n6800), .C1(
        P2_U3151), .C2(n8374), .ZN(P2_U3282) );
  INV_X1 U8627 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6805) );
  INV_X1 U8628 ( .A(n6801), .ZN(n6946) );
  NAND2_X1 U8629 ( .A1(n9325), .A2(n7141), .ZN(n9238) );
  NAND2_X1 U8630 ( .A1(n6946), .A2(n9238), .ZN(n9079) );
  INV_X1 U8631 ( .A(n9079), .ZN(n7137) );
  NOR2_X1 U8632 ( .A1(n9949), .A2(n9887), .ZN(n6802) );
  INV_X1 U8633 ( .A(n9323), .ZN(n9862) );
  OAI222_X1 U8634 ( .A1(n7141), .A2(n6803), .B1(n7137), .B2(n6802), .C1(n9950), 
        .C2(n9862), .ZN(n6806) );
  NAND2_X1 U8635 ( .A1(n6806), .A2(n9967), .ZN(n6804) );
  OAI21_X1 U8636 ( .B1(n9967), .B2(n6805), .A(n6804), .ZN(P1_U3453) );
  NAND2_X1 U8637 ( .A1(n6806), .A2(n9983), .ZN(n6807) );
  OAI21_X1 U8638 ( .B1(n9983), .B2(n5771), .A(n6807), .ZN(P1_U3522) );
  INV_X1 U8639 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6811) );
  NOR2_X1 U8640 ( .A1(n6883), .A2(n8744), .ZN(n6931) );
  INV_X1 U8641 ( .A(n6931), .ZN(n6809) );
  NAND2_X1 U8642 ( .A1(n7685), .A2(n10045), .ZN(n10020) );
  OAI21_X1 U8643 ( .B1(n8731), .B2(n10020), .A(n8305), .ZN(n6808) );
  OAI211_X1 U8644 ( .C1(n10039), .C2(n6936), .A(n6809), .B(n6808), .ZN(n8812)
         );
  NAND2_X1 U8645 ( .A1(n8812), .A2(n10064), .ZN(n6810) );
  OAI21_X1 U8646 ( .B1(n6811), .B2(n10064), .A(n6810), .ZN(P2_U3390) );
  INV_X1 U8647 ( .A(n9328), .ZN(n6813) );
  MUX2_X1 U8648 ( .A(n6814), .B(n6813), .S(n6812), .Z(n6816) );
  NAND2_X1 U8649 ( .A1(n6816), .A2(n6815), .ZN(n6817) );
  OAI211_X1 U8650 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n6818), .A(n6817), .B(n9324), .ZN(n9365) );
  XOR2_X1 U8651 ( .A(n6820), .B(n6819), .Z(n6828) );
  AOI22_X1 U8652 ( .A1(n9433), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6821) );
  OAI21_X1 U8653 ( .B1(n6822), .B2(n9445), .A(n6821), .ZN(n6827) );
  AOI211_X1 U8654 ( .C1(n6825), .C2(n6824), .A(n6823), .B(n9428), .ZN(n6826)
         );
  AOI211_X1 U8655 ( .C1(n9443), .C2(n6828), .A(n6827), .B(n6826), .ZN(n6829)
         );
  NAND2_X1 U8656 ( .A1(n9365), .A2(n6829), .ZN(P1_U3245) );
  INV_X1 U8657 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10280) );
  INV_X1 U8658 ( .A(n6830), .ZN(n6832) );
  INV_X1 U8659 ( .A(n8409), .ZN(n6831) );
  OAI222_X1 U8660 ( .A1(n8899), .A2(n10280), .B1(n8900), .B2(n6832), .C1(
        P2_U3151), .C2(n6831), .ZN(P2_U3281) );
  INV_X1 U8661 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10234) );
  INV_X1 U8662 ( .A(n7607), .ZN(n7612) );
  OAI222_X1 U8663 ( .A1(n9771), .A2(n10234), .B1(n9769), .B2(n6832), .C1(
        P1_U3086), .C2(n7612), .ZN(P1_U3341) );
  XOR2_X1 U8664 ( .A(n6834), .B(n6833), .Z(n6840) );
  OR2_X1 U8665 ( .A1(n8983), .A2(n9862), .ZN(n6836) );
  INV_X1 U8666 ( .A(n9322), .ZN(n9879) );
  OR2_X1 U8667 ( .A1(n9043), .A2(n9879), .ZN(n6835) );
  OAI211_X1 U8668 ( .C1(n7300), .C2(n9039), .A(n6836), .B(n6835), .ZN(n6837)
         );
  AOI21_X1 U8669 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n6838), .A(n6837), .ZN(
        n6839) );
  OAI21_X1 U8670 ( .B1(n6840), .B2(n9052), .A(n6839), .ZN(P1_U3237) );
  INV_X1 U8671 ( .A(n6841), .ZN(n6843) );
  OAI21_X1 U8672 ( .B1(n6852), .B2(n6843), .A(n6842), .ZN(n6847) );
  MUX2_X1 U8673 ( .A(n6845), .B(n6844), .S(n4438), .Z(n6971) );
  XNOR2_X1 U8674 ( .A(n6971), .B(n6861), .ZN(n6846) );
  NAND2_X1 U8675 ( .A1(n6847), .A2(n6846), .ZN(n6970) );
  OAI211_X1 U8676 ( .C1(n6847), .C2(n6846), .A(n6970), .B(n10406), .ZN(n6860)
         );
  INV_X1 U8677 ( .A(n6861), .ZN(n6972) );
  NOR2_X1 U8678 ( .A1(n6844), .A2(n6850), .ZN(n6976) );
  AOI21_X1 U8679 ( .B1(n6850), .B2(n6844), .A(n6976), .ZN(n6851) );
  NOR2_X1 U8680 ( .A1(n6851), .A2(n9985), .ZN(n6858) );
  NAND2_X1 U8681 ( .A1(n6854), .A2(n6861), .ZN(n6982) );
  AOI21_X1 U8682 ( .B1(n6855), .B2(n6845), .A(n6979), .ZN(n6856) );
  NAND2_X1 U8683 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7044) );
  OAI21_X1 U8684 ( .B1(n10002), .B2(n6856), .A(n7044), .ZN(n6857) );
  AOI211_X1 U8685 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n10405), .A(n6858), .B(
        n6857), .ZN(n6859) );
  OAI211_X1 U8686 ( .C1(n9996), .C2(n6861), .A(n6860), .B(n6859), .ZN(P2_U3187) );
  XNOR2_X1 U8687 ( .A(n7029), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n6864) );
  OAI21_X1 U8688 ( .B1(n6866), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6862), .ZN(
        n6863) );
  NOR2_X1 U8689 ( .A1(n6863), .A2(n6864), .ZN(n7025) );
  AOI211_X1 U8690 ( .C1(n6864), .C2(n6863), .A(n9428), .B(n7025), .ZN(n6874)
         );
  OAI21_X1 U8691 ( .B1(n6866), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6865), .ZN(
        n6869) );
  INV_X1 U8692 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9977) );
  MUX2_X1 U8693 ( .A(n9977), .B(P1_REG1_REG_10__SCAN_IN), .S(n7029), .Z(n6868)
         );
  INV_X1 U8694 ( .A(n7032), .ZN(n6867) );
  AOI211_X1 U8695 ( .C1(n6869), .C2(n6868), .A(n9446), .B(n6867), .ZN(n6873)
         );
  INV_X1 U8696 ( .A(n7029), .ZN(n6871) );
  NOR2_X1 U8697 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10141), .ZN(n7774) );
  AOI21_X1 U8698 ( .B1(n9433), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7774), .ZN(
        n6870) );
  OAI21_X1 U8699 ( .B1(n6871), .B2(n9445), .A(n6870), .ZN(n6872) );
  OR3_X1 U8700 ( .A1(n6874), .A2(n6873), .A3(n6872), .ZN(P1_U3253) );
  INV_X1 U8701 ( .A(n8328), .ZN(n6876) );
  AND2_X1 U8702 ( .A1(n6963), .A2(n6877), .ZN(n6878) );
  NAND2_X1 U8703 ( .A1(n7938), .A2(n6936), .ZN(n6880) );
  NAND2_X1 U8704 ( .A1(n6881), .A2(n6880), .ZN(n6896) );
  XNOR2_X1 U8705 ( .A(n6913), .B(n7007), .ZN(n6884) );
  XNOR2_X1 U8706 ( .A(n6884), .B(n8353), .ZN(n6895) );
  NAND2_X1 U8707 ( .A1(n6896), .A2(n6895), .ZN(n6886) );
  NAND2_X1 U8708 ( .A1(n6884), .A2(n6883), .ZN(n6885) );
  NAND2_X1 U8709 ( .A1(n6886), .A2(n6885), .ZN(n7005) );
  XNOR2_X1 U8710 ( .A(n7007), .B(n6887), .ZN(n7006) );
  XNOR2_X1 U8711 ( .A(n4442), .B(n7006), .ZN(n7004) );
  XOR2_X1 U8712 ( .A(n7005), .B(n7004), .Z(n6894) );
  INV_X1 U8713 ( .A(n8110), .ZN(n8066) );
  INV_X1 U8714 ( .A(n4427), .ZN(n8068) );
  OAI22_X1 U8715 ( .A1(n8116), .A2(n10006), .B1(n8068), .B2(n6883), .ZN(n6892)
         );
  NOR2_X1 U8716 ( .A1(n6897), .A2(n6890), .ZN(n6891) );
  AOI211_X1 U8717 ( .C1(n8066), .C2(n8351), .A(n6892), .B(n6891), .ZN(n6893)
         );
  OAI21_X1 U8718 ( .B1(n6894), .B2(n8039), .A(n6893), .ZN(P2_U3177) );
  XOR2_X1 U8719 ( .A(n6896), .B(n6895), .Z(n6901) );
  OAI22_X1 U8720 ( .A1(n8116), .A2(n6882), .B1(n8068), .B2(n6076), .ZN(n6899)
         );
  NOR2_X1 U8721 ( .A1(n6897), .A2(n6997), .ZN(n6898) );
  AOI211_X1 U8722 ( .C1(n8066), .C2(n4442), .A(n6899), .B(n6898), .ZN(n6900)
         );
  OAI21_X1 U8723 ( .B1(n8039), .B2(n6901), .A(n6900), .ZN(P2_U3162) );
  INV_X1 U8724 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6903) );
  INV_X1 U8725 ( .A(n6902), .ZN(n6904) );
  INV_X1 U8726 ( .A(n9381), .ZN(n9387) );
  OAI222_X1 U8727 ( .A1(n9771), .A2(n6903), .B1(n9769), .B2(n6904), .C1(
        P1_U3086), .C2(n9387), .ZN(P1_U3340) );
  INV_X1 U8728 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6905) );
  INV_X1 U8729 ( .A(n8453), .ZN(n8414) );
  OAI222_X1 U8730 ( .A1(n8899), .A2(n6905), .B1(n8900), .B2(n6904), .C1(
        P2_U3151), .C2(n8414), .ZN(P2_U3280) );
  OAI21_X1 U8731 ( .B1(n8304), .B2(n6907), .A(n6906), .ZN(n7001) );
  NAND2_X1 U8732 ( .A1(n6075), .A2(n8731), .ZN(n6909) );
  OAI21_X1 U8733 ( .B1(n8192), .B2(n6909), .A(n8742), .ZN(n6910) );
  NAND2_X1 U8734 ( .A1(n6910), .A2(n8354), .ZN(n6912) );
  NAND2_X1 U8735 ( .A1(n4442), .A2(n8728), .ZN(n6911) );
  OAI211_X1 U8736 ( .C1(n6908), .C2(n8740), .A(n6912), .B(n6911), .ZN(n6998)
         );
  AOI21_X1 U8737 ( .B1(n10020), .B2(n7001), .A(n6998), .ZN(n6918) );
  AOI22_X1 U8738 ( .A1(n8808), .A2(n6913), .B1(n6533), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n6914) );
  OAI21_X1 U8739 ( .B1(n6918), .B2(n6533), .A(n6914), .ZN(P2_U3460) );
  INV_X1 U8740 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6915) );
  OAI22_X1 U8741 ( .A1(n6882), .A2(n8864), .B1(n10064), .B2(n6915), .ZN(n6916)
         );
  INV_X1 U8742 ( .A(n6916), .ZN(n6917) );
  OAI21_X1 U8743 ( .B1(n6918), .B2(n10062), .A(n6917), .ZN(P2_U3393) );
  NAND2_X1 U8744 ( .A1(n6875), .A2(n6919), .ZN(n6923) );
  NAND2_X1 U8745 ( .A1(n6921), .A2(n6920), .ZN(n6922) );
  AND2_X1 U8746 ( .A1(n6923), .A2(n6922), .ZN(n6924) );
  NAND2_X1 U8747 ( .A1(n6925), .A2(n6924), .ZN(n6932) );
  INV_X1 U8748 ( .A(n6932), .ZN(n6926) );
  INV_X1 U8749 ( .A(n8747), .ZN(n8734) );
  NAND2_X1 U8750 ( .A1(n6926), .A2(n8734), .ZN(n8720) );
  AND3_X1 U8751 ( .A1(n8305), .A2(n10039), .A3(n6929), .ZN(n6930) );
  AOI211_X1 U8752 ( .C1(n8718), .C2(P2_REG3_REG_0__SCAN_IN), .A(n6931), .B(
        n6930), .ZN(n6933) );
  MUX2_X1 U8753 ( .A(n6934), .B(n6933), .S(n8748), .Z(n6935) );
  OAI21_X1 U8754 ( .B1(n8720), .B2(n6936), .A(n6935), .ZN(P2_U3233) );
  XNOR2_X1 U8755 ( .A(n6938), .B(n6937), .ZN(n6939) );
  NAND2_X1 U8756 ( .A1(n6939), .A2(n9031), .ZN(n6943) );
  INV_X1 U8757 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10172) );
  NOR2_X1 U8758 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10172), .ZN(n9342) );
  INV_X1 U8759 ( .A(n9829), .ZN(n7161) );
  OAI22_X1 U8760 ( .A1(n6940), .A2(n8983), .B1(n9043), .B2(n7161), .ZN(n6941)
         );
  AOI211_X1 U8761 ( .C1(n9833), .C2(n9050), .A(n9342), .B(n6941), .ZN(n6942)
         );
  OAI211_X1 U8762 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9048), .A(n6943), .B(
        n6942), .ZN(P1_U3218) );
  INV_X1 U8763 ( .A(n6944), .ZN(n6968) );
  INV_X1 U8764 ( .A(n9397), .ZN(n9402) );
  INV_X1 U8765 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10283) );
  OAI222_X1 U8766 ( .A1(n9769), .A2(n6968), .B1(n9402), .B2(P1_U3086), .C1(
        n10283), .C2(n9771), .ZN(P1_U3339) );
  INV_X1 U8767 ( .A(n9960), .ZN(n9942) );
  XNOR2_X1 U8768 ( .A(n9080), .B(n6945), .ZN(n9853) );
  OAI211_X1 U8769 ( .C1(n9237), .C2(n7141), .A(n9837), .B(n7302), .ZN(n9849)
         );
  OAI21_X1 U8770 ( .B1(n9237), .B2(n9944), .A(n9849), .ZN(n6951) );
  INV_X1 U8771 ( .A(n9814), .ZN(n9964) );
  XNOR2_X1 U8772 ( .A(n6946), .B(n9080), .ZN(n6948) );
  AOI22_X1 U8773 ( .A1(n9918), .A2(n9325), .B1(n4429), .B2(n9891), .ZN(n6947)
         );
  OAI21_X1 U8774 ( .B1(n6948), .B2(n9933), .A(n6947), .ZN(n6949) );
  AOI21_X1 U8775 ( .B1(n9964), .B2(n9853), .A(n6949), .ZN(n9856) );
  INV_X1 U8776 ( .A(n9856), .ZN(n6950) );
  AOI211_X1 U8777 ( .C1(n9942), .C2(n9853), .A(n6951), .B(n6950), .ZN(n9861)
         );
  NAND2_X1 U8778 ( .A1(n9981), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6952) );
  OAI21_X1 U8779 ( .B1(n9861), .B2(n9981), .A(n6952), .ZN(P1_U3523) );
  NAND3_X1 U8780 ( .A1(n6954), .A2(n6961), .A3(n6955), .ZN(n6956) );
  NAND2_X1 U8781 ( .A1(n6953), .A2(n6956), .ZN(n6957) );
  NAND2_X1 U8782 ( .A1(n6957), .A2(n8731), .ZN(n6959) );
  AOI22_X1 U8783 ( .A1(n8726), .A2(n4442), .B1(n7998), .B2(n8728), .ZN(n6958)
         );
  AND2_X1 U8784 ( .A1(n6959), .A2(n6958), .ZN(n10013) );
  OAI22_X1 U8785 ( .A1(n8720), .A2(n7008), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8745), .ZN(n6960) );
  AOI21_X1 U8786 ( .B1(n8752), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6960), .ZN(
        n6967) );
  XNOR2_X1 U8787 ( .A(n6961), .B(n6962), .ZN(n10010) );
  NOR2_X1 U8788 ( .A1(n6963), .A2(n8519), .ZN(n7107) );
  INV_X1 U8789 ( .A(n7107), .ZN(n6964) );
  NAND2_X1 U8790 ( .A1(n7685), .A2(n6964), .ZN(n6965) );
  NAND2_X1 U8791 ( .A1(n10010), .A2(n8753), .ZN(n6966) );
  OAI211_X1 U8792 ( .C1(n10013), .C2(n8752), .A(n6967), .B(n6966), .ZN(
        P2_U3230) );
  INV_X1 U8793 ( .A(n8456), .ZN(n8475) );
  OAI222_X1 U8794 ( .A1(P2_U3151), .A2(n8475), .B1(n8899), .B2(n6969), .C1(
        n6968), .C2(n8900), .ZN(P2_U3279) );
  MUX2_X1 U8795 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n4446), .Z(n7072) );
  XNOR2_X1 U8796 ( .A(n7072), .B(n7075), .ZN(n6974) );
  OAI21_X1 U8797 ( .B1(n6972), .B2(n6971), .A(n6970), .ZN(n6973) );
  NOR2_X1 U8798 ( .A1(n6973), .A2(n6974), .ZN(n7073) );
  AOI21_X1 U8799 ( .B1(n6974), .B2(n6973), .A(n7073), .ZN(n6989) );
  INV_X1 U8800 ( .A(n7075), .ZN(n7083) );
  XNOR2_X1 U8801 ( .A(n7083), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n6975) );
  OR3_X1 U8802 ( .A1(n6977), .A2(n6976), .A3(n6975), .ZN(n6978) );
  AOI21_X1 U8803 ( .B1(n7084), .B2(n6978), .A(n9985), .ZN(n6986) );
  XNOR2_X1 U8804 ( .A(n7075), .B(n7251), .ZN(n6980) );
  NOR2_X1 U8805 ( .A1(n6980), .A2(n6979), .ZN(n6983) );
  INV_X1 U8806 ( .A(n7077), .ZN(n6981) );
  AOI21_X1 U8807 ( .B1(n6983), .B2(n6982), .A(n6981), .ZN(n6984) );
  NAND2_X1 U8808 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7062) );
  OAI21_X1 U8809 ( .B1(n10002), .B2(n6984), .A(n7062), .ZN(n6985) );
  AOI211_X1 U8810 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n10405), .A(n6986), .B(
        n6985), .ZN(n6988) );
  NAND2_X1 U8811 ( .A1(n10411), .A2(n7083), .ZN(n6987) );
  OAI211_X1 U8812 ( .C1(n6989), .C2(n8535), .A(n6988), .B(n6987), .ZN(P2_U3188) );
  AOI21_X1 U8813 ( .B1(n6991), .B2(n6990), .A(n9052), .ZN(n6993) );
  NAND2_X1 U8814 ( .A1(n6993), .A2(n6992), .ZN(n6996) );
  AND2_X1 U8815 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9355) );
  INV_X1 U8816 ( .A(n9321), .ZN(n9878) );
  OAI22_X1 U8817 ( .A1(n9879), .A2(n8983), .B1(n9043), .B2(n9878), .ZN(n6994)
         );
  AOI211_X1 U8818 ( .C1(n9881), .C2(n9050), .A(n9355), .B(n6994), .ZN(n6995)
         );
  OAI211_X1 U8819 ( .C1(n9048), .C2(n7312), .A(n6996), .B(n6995), .ZN(P1_U3230) );
  OAI22_X1 U8820 ( .A1(n8720), .A2(n6882), .B1(n6997), .B2(n8745), .ZN(n7000)
         );
  MUX2_X1 U8821 ( .A(n6998), .B(P2_REG2_REG_1__SCAN_IN), .S(n8752), .Z(n6999)
         );
  AOI211_X1 U8822 ( .C1(n8753), .C2(n7001), .A(n7000), .B(n6999), .ZN(n7002)
         );
  INV_X1 U8823 ( .A(n7002), .ZN(P2_U3232) );
  XNOR2_X1 U8824 ( .A(n7003), .B(n7007), .ZN(n7039) );
  NAND2_X1 U8825 ( .A1(n7005), .A2(n7004), .ZN(n7992) );
  NAND2_X1 U8826 ( .A1(n6088), .A2(n7006), .ZN(n7991) );
  INV_X1 U8827 ( .A(n7993), .ZN(n7009) );
  NAND2_X1 U8828 ( .A1(n7010), .A2(n8351), .ZN(n7011) );
  INV_X1 U8829 ( .A(n7043), .ZN(n7013) );
  AOI21_X1 U8830 ( .B1(n7014), .B2(n7012), .A(n7013), .ZN(n7024) );
  INV_X1 U8831 ( .A(n7015), .ZN(n7124) );
  AND2_X1 U8832 ( .A1(n7016), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7646) );
  INV_X1 U8833 ( .A(n7018), .ZN(n7019) );
  AOI21_X1 U8834 ( .B1(n4427), .B2(n8351), .A(n7019), .ZN(n7021) );
  NAND2_X1 U8835 ( .A1(n8037), .A2(n10016), .ZN(n7020) );
  OAI211_X1 U8836 ( .C1(n7056), .C2(n8110), .A(n7021), .B(n7020), .ZN(n7022)
         );
  AOI21_X1 U8837 ( .B1(n7124), .B2(n8113), .A(n7022), .ZN(n7023) );
  OAI21_X1 U8838 ( .B1(n7024), .B2(n8039), .A(n7023), .ZN(P2_U3170) );
  NAND2_X1 U8839 ( .A1(n7237), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7026) );
  OAI21_X1 U8840 ( .B1(n7237), .B2(P1_REG2_REG_11__SCAN_IN), .A(n7026), .ZN(
        n7027) );
  NOR2_X1 U8841 ( .A1(n7028), .A2(n7027), .ZN(n7236) );
  AOI211_X1 U8842 ( .C1(n7028), .C2(n7027), .A(n9428), .B(n7236), .ZN(n7038)
         );
  NAND2_X1 U8843 ( .A1(n7029), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7031) );
  MUX2_X1 U8844 ( .A(n5320), .B(P1_REG1_REG_11__SCAN_IN), .S(n7237), .Z(n7030)
         );
  AOI21_X1 U8845 ( .B1(n7032), .B2(n7031), .A(n7030), .ZN(n7231) );
  AND3_X1 U8846 ( .A1(n7032), .A2(n7031), .A3(n7030), .ZN(n7033) );
  NOR3_X1 U8847 ( .A1(n7231), .A2(n7033), .A3(n9446), .ZN(n7037) );
  INV_X1 U8848 ( .A(n7237), .ZN(n7035) );
  AND2_X1 U8849 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7861) );
  AOI21_X1 U8850 ( .B1(n9433), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n7861), .ZN(
        n7034) );
  OAI21_X1 U8851 ( .B1(n7035), .B2(n9445), .A(n7034), .ZN(n7036) );
  OR3_X1 U8852 ( .A1(n7038), .A2(n7037), .A3(n7036), .ZN(P1_U3254) );
  INV_X1 U8853 ( .A(n7998), .ZN(n7041) );
  INV_X1 U8854 ( .A(n7039), .ZN(n7040) );
  NAND2_X1 U8855 ( .A1(n7041), .A2(n7040), .ZN(n7042) );
  XNOR2_X1 U8856 ( .A(n7007), .B(n10022), .ZN(n7055) );
  XNOR2_X1 U8857 ( .A(n7055), .B(n8350), .ZN(n7058) );
  XOR2_X1 U8858 ( .A(n7059), .B(n7058), .Z(n7051) );
  INV_X1 U8859 ( .A(n7098), .ZN(n7049) );
  INV_X1 U8860 ( .A(n8349), .ZN(n7444) );
  INV_X1 U8861 ( .A(n7044), .ZN(n7045) );
  AOI21_X1 U8862 ( .B1(n4427), .B2(n7998), .A(n7045), .ZN(n7047) );
  NAND2_X1 U8863 ( .A1(n8037), .A2(n10022), .ZN(n7046) );
  OAI211_X1 U8864 ( .C1(n7444), .C2(n8110), .A(n7047), .B(n7046), .ZN(n7048)
         );
  AOI21_X1 U8865 ( .B1(n7049), .B2(n8113), .A(n7048), .ZN(n7050) );
  OAI21_X1 U8866 ( .B1(n7051), .B2(n8039), .A(n7050), .ZN(P2_U3167) );
  INV_X1 U8867 ( .A(n7052), .ZN(n7068) );
  AOI22_X1 U8868 ( .A1(n9423), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n7053), .ZN(n7054) );
  OAI21_X1 U8869 ( .B1(n7068), .B2(n9769), .A(n7054), .ZN(P1_U3338) );
  INV_X1 U8870 ( .A(n8113), .ZN(n8044) );
  AND2_X1 U8871 ( .A1(n7056), .A2(n7055), .ZN(n7057) );
  XNOR2_X1 U8872 ( .A(n7007), .B(n10028), .ZN(n7197) );
  XNOR2_X1 U8873 ( .A(n7197), .B(n8349), .ZN(n7060) );
  OAI211_X1 U8874 ( .C1(n7061), .C2(n7060), .A(n7200), .B(n8104), .ZN(n7067)
         );
  INV_X1 U8875 ( .A(n7062), .ZN(n7065) );
  INV_X1 U8876 ( .A(n8348), .ZN(n7284) );
  OAI22_X1 U8877 ( .A1(n8116), .A2(n7063), .B1(n7284), .B2(n8110), .ZN(n7064)
         );
  AOI211_X1 U8878 ( .C1(n4427), .C2(n8350), .A(n7065), .B(n7064), .ZN(n7066)
         );
  OAI211_X1 U8879 ( .C1(n7252), .C2(n8044), .A(n7067), .B(n7066), .ZN(P2_U3179) );
  INV_X1 U8880 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7069) );
  INV_X1 U8881 ( .A(n8502), .ZN(n8471) );
  OAI222_X1 U8882 ( .A1(n8899), .A2(n7069), .B1(n8900), .B2(n7068), .C1(
        P2_U3151), .C2(n8471), .ZN(P2_U3278) );
  MUX2_X1 U8883 ( .A(n7071), .B(n7070), .S(n4446), .Z(n7170) );
  XNOR2_X1 U8884 ( .A(n7170), .B(n7079), .ZN(n7172) );
  INV_X1 U8885 ( .A(n7072), .ZN(n7074) );
  XOR2_X1 U8886 ( .A(n7172), .B(n7173), .Z(n7091) );
  NAND2_X1 U8887 ( .A1(n7075), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7076) );
  NAND2_X1 U8888 ( .A1(n7077), .A2(n7076), .ZN(n7181) );
  XNOR2_X1 U8889 ( .A(n7181), .B(n7079), .ZN(n7078) );
  NAND2_X1 U8890 ( .A1(n7078), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7183) );
  OAI21_X1 U8891 ( .B1(n7078), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7183), .ZN(
        n7089) );
  INV_X1 U8892 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7081) );
  NAND2_X1 U8893 ( .A1(n10411), .A2(n7079), .ZN(n7080) );
  NAND2_X1 U8894 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7205) );
  OAI211_X1 U8895 ( .C1(n10005), .C2(n7081), .A(n7080), .B(n7205), .ZN(n7088)
         );
  NAND2_X1 U8896 ( .A1(n7084), .A2(n5059), .ZN(n7177) );
  AOI21_X1 U8897 ( .B1(n7070), .B2(n7085), .A(n7176), .ZN(n7086) );
  NOR2_X1 U8898 ( .A1(n7086), .A2(n9985), .ZN(n7087) );
  AOI211_X1 U8899 ( .C1(n10419), .C2(n7089), .A(n7088), .B(n7087), .ZN(n7090)
         );
  OAI21_X1 U8900 ( .B1(n7091), .B2(n8535), .A(n7090), .ZN(P2_U3189) );
  INV_X1 U8901 ( .A(n7096), .ZN(n8307) );
  XNOR2_X1 U8902 ( .A(n7092), .B(n8307), .ZN(n7093) );
  NAND2_X1 U8903 ( .A1(n7093), .A2(n8731), .ZN(n7095) );
  AOI22_X1 U8904 ( .A1(n8726), .A2(n7998), .B1(n8349), .B2(n8728), .ZN(n7094)
         );
  AND2_X1 U8905 ( .A1(n7095), .A2(n7094), .ZN(n10025) );
  XNOR2_X1 U8906 ( .A(n7097), .B(n7096), .ZN(n10021) );
  NOR2_X1 U8907 ( .A1(n8748), .A2(n6845), .ZN(n7101) );
  OAI22_X1 U8908 ( .A1(n8720), .A2(n7099), .B1(n7098), .B2(n8745), .ZN(n7100)
         );
  AOI211_X1 U8909 ( .C1(n10021), .C2(n8753), .A(n7101), .B(n7100), .ZN(n7102)
         );
  OAI21_X1 U8910 ( .B1(n8752), .B2(n10025), .A(n7102), .ZN(P2_U3228) );
  OAI21_X1 U8911 ( .B1(n7105), .B2(n7103), .A(n7104), .ZN(n7106) );
  INV_X1 U8912 ( .A(n7106), .ZN(n10007) );
  NAND2_X1 U8913 ( .A1(n8748), .A2(n7107), .ZN(n7963) );
  AOI22_X1 U8914 ( .A1(n8726), .A2(n8353), .B1(n8351), .B2(n8728), .ZN(n7112)
         );
  INV_X1 U8915 ( .A(n6954), .ZN(n7110) );
  AND3_X1 U8916 ( .A1(n6908), .A2(n7103), .A3(n7108), .ZN(n7109) );
  OAI21_X1 U8917 ( .B1(n7110), .B2(n7109), .A(n8731), .ZN(n7111) );
  OAI211_X1 U8918 ( .C1(n10007), .C2(n7685), .A(n7112), .B(n7111), .ZN(n10009)
         );
  OAI22_X1 U8919 ( .A1(n10006), .A2(n8747), .B1(n6890), .B2(n8745), .ZN(n7113)
         );
  NOR2_X1 U8920 ( .A1(n10009), .A2(n7113), .ZN(n7114) );
  MUX2_X1 U8921 ( .A(n7115), .B(n7114), .S(n8748), .Z(n7116) );
  OAI21_X1 U8922 ( .B1(n10007), .B2(n7963), .A(n7116), .ZN(P2_U3231) );
  OAI21_X1 U8923 ( .B1(n7117), .B2(n8303), .A(n7118), .ZN(n10017) );
  INV_X1 U8924 ( .A(n10017), .ZN(n7127) );
  NAND3_X1 U8925 ( .A1(n6953), .A2(n8303), .A3(n7120), .ZN(n7121) );
  NAND2_X1 U8926 ( .A1(n7119), .A2(n7121), .ZN(n7122) );
  AOI222_X1 U8927 ( .A1(n8731), .A2(n7122), .B1(n8351), .B2(n8726), .C1(n8350), 
        .C2(n8728), .ZN(n10019) );
  MUX2_X1 U8928 ( .A(n7123), .B(n10019), .S(n8748), .Z(n7126) );
  AOI22_X1 U8929 ( .A1(n8708), .A2(n10016), .B1(n8718), .B2(n7124), .ZN(n7125)
         );
  OAI211_X1 U8930 ( .C1(n7127), .C2(n8711), .A(n7126), .B(n7125), .ZN(P2_U3229) );
  NAND2_X1 U8931 ( .A1(n9598), .A2(n5713), .ZN(n9606) );
  AOI21_X1 U8932 ( .B1(n9851), .B2(n9837), .A(n7133), .ZN(n7142) );
  NOR2_X1 U8933 ( .A1(n9857), .A2(n9950), .ZN(n9600) );
  OAI22_X1 U8934 ( .A1(n9598), .A2(n6581), .B1(n7134), .B2(n9846), .ZN(n7139)
         );
  NOR4_X1 U8935 ( .A1(n7137), .A2(n7136), .A3(n7135), .A4(n9857), .ZN(n7138)
         );
  AOI211_X1 U8936 ( .C1(n9600), .C2(n9323), .A(n7139), .B(n7138), .ZN(n7140)
         );
  OAI21_X1 U8937 ( .B1(n7142), .B2(n7141), .A(n7140), .ZN(P1_U3293) );
  INV_X1 U8938 ( .A(n8522), .ZN(n8505) );
  INV_X1 U8939 ( .A(n7143), .ZN(n7145) );
  INV_X1 U8940 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7144) );
  OAI222_X1 U8941 ( .A1(P2_U3151), .A2(n8505), .B1(n8900), .B2(n7145), .C1(
        n7144), .C2(n8899), .ZN(P2_U3277) );
  INV_X1 U8942 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7146) );
  INV_X1 U8943 ( .A(n9441), .ZN(n9436) );
  OAI222_X1 U8944 ( .A1(n9771), .A2(n7146), .B1(n9436), .B2(P1_U3086), .C1(
        n9769), .C2(n7145), .ZN(P1_U3337) );
  NAND2_X1 U8945 ( .A1(n7147), .A2(n7148), .ZN(n7149) );
  XOR2_X1 U8946 ( .A(n7150), .B(n7149), .Z(n7155) );
  NOR2_X1 U8947 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5176), .ZN(n9368) );
  NOR2_X1 U8948 ( .A1(n9043), .A2(n9811), .ZN(n7151) );
  AOI211_X1 U8949 ( .C1(n9045), .C2(n9829), .A(n9368), .B(n7151), .ZN(n7154)
         );
  INV_X1 U8950 ( .A(n7152), .ZN(n7163) );
  AOI22_X1 U8951 ( .A1(n9050), .A2(n9889), .B1(n7163), .B2(n8991), .ZN(n7153)
         );
  OAI211_X1 U8952 ( .C1(n7155), .C2(n9052), .A(n7154), .B(n7153), .ZN(P1_U3227) );
  NOR2_X1 U8953 ( .A1(n5713), .A2(n7156), .ZN(n7157) );
  NAND2_X1 U8954 ( .A1(n9598), .A2(n7157), .ZN(n7384) );
  NAND2_X1 U8955 ( .A1(n9598), .A2(n9964), .ZN(n7158) );
  XNOR2_X1 U8956 ( .A(n7160), .B(n7159), .ZN(n9895) );
  XNOR2_X1 U8957 ( .A(n9242), .B(n9083), .ZN(n7162) );
  OAI22_X1 U8958 ( .A1(n7162), .A2(n9933), .B1(n7161), .B2(n9952), .ZN(n9897)
         );
  NAND2_X1 U8959 ( .A1(n9897), .A2(n9598), .ZN(n7169) );
  INV_X1 U8960 ( .A(n9600), .ZN(n7809) );
  INV_X1 U8961 ( .A(n9846), .ZN(n9820) );
  AOI22_X1 U8962 ( .A1(n9857), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7163), .B2(
        n9820), .ZN(n7164) );
  OAI21_X1 U8963 ( .B1(n7809), .B2(n9811), .A(n7164), .ZN(n7167) );
  AOI21_X1 U8964 ( .B1(n7311), .B2(n9889), .A(n9822), .ZN(n7165) );
  NAND2_X1 U8965 ( .A1(n7165), .A2(n7224), .ZN(n9892) );
  NOR2_X1 U8966 ( .A1(n9892), .A2(n9606), .ZN(n7166) );
  AOI211_X1 U8967 ( .C1(n7133), .C2(n9889), .A(n7167), .B(n7166), .ZN(n7168)
         );
  OAI211_X1 U8968 ( .C1(n9629), .C2(n9895), .A(n7169), .B(n7168), .ZN(P1_U3288) );
  INV_X1 U8969 ( .A(n7170), .ZN(n7171) );
  OAI22_X1 U8970 ( .A1(n7173), .A2(n7172), .B1(n7171), .B2(n7180), .ZN(n7175)
         );
  MUX2_X1 U8971 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n4446), .Z(n7395) );
  XNOR2_X1 U8972 ( .A(n7395), .B(n7189), .ZN(n7174) );
  NAND2_X1 U8973 ( .A1(n7175), .A2(n7174), .ZN(n7396) );
  OAI21_X1 U8974 ( .B1(n7175), .B2(n7174), .A(n7396), .ZN(n7195) );
  NAND2_X1 U8975 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7402), .ZN(n7392) );
  OAI21_X1 U8976 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7402), .A(n7392), .ZN(
        n7178) );
  AOI21_X1 U8977 ( .B1(n4538), .B2(n7178), .A(n7393), .ZN(n7179) );
  NOR2_X1 U8978 ( .A1(n7179), .A2(n9985), .ZN(n7194) );
  NAND2_X1 U8979 ( .A1(n7181), .A2(n7180), .ZN(n7182) );
  NAND2_X1 U8980 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7402), .ZN(n7184) );
  OAI21_X1 U8981 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7402), .A(n7184), .ZN(
        n7185) );
  AOI21_X1 U8982 ( .B1(n7186), .B2(n7185), .A(n7401), .ZN(n7192) );
  INV_X1 U8983 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7187) );
  NAND2_X1 U8984 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7288) );
  OAI21_X1 U8985 ( .B1(n10005), .B2(n7187), .A(n7288), .ZN(n7188) );
  INV_X1 U8986 ( .A(n7188), .ZN(n7191) );
  NAND2_X1 U8987 ( .A1(n10411), .A2(n7189), .ZN(n7190) );
  OAI211_X1 U8988 ( .C1(n7192), .C2(n10002), .A(n7191), .B(n7190), .ZN(n7193)
         );
  AOI211_X1 U8989 ( .C1(n7195), .C2(n10406), .A(n7194), .B(n7193), .ZN(n7196)
         );
  INV_X1 U8990 ( .A(n7196), .ZN(P2_U3190) );
  XNOR2_X1 U8991 ( .A(n7515), .B(n7943), .ZN(n7282) );
  XNOR2_X1 U8992 ( .A(n7282), .B(n8348), .ZN(n7204) );
  INV_X1 U8993 ( .A(n7197), .ZN(n7198) );
  NAND2_X1 U8994 ( .A1(n7198), .A2(n8349), .ZN(n7199) );
  INV_X1 U8995 ( .A(n7286), .ZN(n7202) );
  AOI21_X1 U8996 ( .B1(n7204), .B2(n7203), .A(n7202), .ZN(n7211) );
  INV_X1 U8997 ( .A(n8347), .ZN(n7556) );
  INV_X1 U8998 ( .A(n7205), .ZN(n7206) );
  AOI21_X1 U8999 ( .B1(n4427), .B2(n8349), .A(n7206), .ZN(n7207) );
  OAI21_X1 U9000 ( .B1(n7556), .B2(n8110), .A(n7207), .ZN(n7209) );
  NOR2_X1 U9001 ( .A1(n8044), .A2(n7446), .ZN(n7208) );
  AOI211_X1 U9002 ( .C1(n8037), .C2(n7518), .A(n7209), .B(n7208), .ZN(n7210)
         );
  OAI21_X1 U9003 ( .B1(n7211), .B2(n8039), .A(n7210), .ZN(P2_U3153) );
  INV_X1 U9004 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7214) );
  NAND2_X1 U9005 ( .A1(n4433), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7213) );
  INV_X1 U9006 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8546) );
  OR2_X1 U9007 ( .A1(n4439), .A2(n8546), .ZN(n7212) );
  OAI211_X1 U9008 ( .C1(n4445), .C2(n7214), .A(n7213), .B(n7212), .ZN(n7215)
         );
  INV_X1 U9009 ( .A(n7215), .ZN(n7216) );
  NAND2_X1 U9010 ( .A1(n8497), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7218) );
  OAI21_X1 U9011 ( .B1(n8543), .B2(n8497), .A(n7218), .ZN(P2_U3522) );
  NAND2_X1 U9012 ( .A1(n8497), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7219) );
  OAI21_X1 U9013 ( .B1(n8553), .B2(n8497), .A(n7219), .ZN(P2_U3520) );
  XNOR2_X1 U9014 ( .A(n7220), .B(n7223), .ZN(n7221) );
  OAI222_X1 U9015 ( .A1(n9950), .A2(n7623), .B1(n9952), .B2(n9878), .C1(n7221), 
        .C2(n9933), .ZN(n9900) );
  INV_X1 U9016 ( .A(n9900), .ZN(n7230) );
  XNOR2_X1 U9017 ( .A(n7222), .B(n7223), .ZN(n9902) );
  OAI211_X1 U9018 ( .C1(n4836), .C2(n9899), .A(n9837), .B(n9823), .ZN(n9898)
         );
  OAI22_X1 U9019 ( .A1(n9598), .A2(n7225), .B1(n7263), .B2(n9846), .ZN(n7226)
         );
  AOI21_X1 U9020 ( .B1(n7133), .B2(n7265), .A(n7226), .ZN(n7227) );
  OAI21_X1 U9021 ( .B1(n9898), .B2(n9606), .A(n7227), .ZN(n7228) );
  AOI21_X1 U9022 ( .B1(n9902), .B2(n9841), .A(n7228), .ZN(n7229) );
  OAI21_X1 U9023 ( .B1(n7230), .B2(n9857), .A(n7229), .ZN(P1_U3287) );
  INV_X1 U9024 ( .A(n7275), .ZN(n7244) );
  MUX2_X1 U9025 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n5342), .S(n7275), .Z(n7233)
         );
  AOI21_X1 U9026 ( .B1(n7237), .B2(P1_REG1_REG_11__SCAN_IN), .A(n7231), .ZN(
        n7232) );
  NAND2_X1 U9027 ( .A1(n7232), .A2(n7233), .ZN(n7270) );
  OAI21_X1 U9028 ( .B1(n7233), .B2(n7232), .A(n7270), .ZN(n7234) );
  NAND2_X1 U9029 ( .A1(n7234), .A2(n9443), .ZN(n7243) );
  NOR2_X1 U9030 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7235), .ZN(n8953) );
  XNOR2_X1 U9031 ( .A(n7275), .B(n7238), .ZN(n7239) );
  NAND2_X1 U9032 ( .A1(n7239), .A2(n7240), .ZN(n7274) );
  AOI221_X1 U9033 ( .B1(n7240), .B2(n7274), .C1(n7239), .C2(n7274), .A(n9428), 
        .ZN(n7241) );
  AOI211_X1 U9034 ( .C1(n9433), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n8953), .B(
        n7241), .ZN(n7242) );
  OAI211_X1 U9035 ( .C1(n9445), .C2(n7244), .A(n7243), .B(n7242), .ZN(P1_U3255) );
  XNOR2_X1 U9036 ( .A(n7245), .B(n6430), .ZN(n10027) );
  NAND2_X1 U9037 ( .A1(n7246), .A2(n8310), .ZN(n7247) );
  NAND3_X1 U9038 ( .A1(n7248), .A2(n8731), .A3(n7247), .ZN(n7250) );
  AOI22_X1 U9039 ( .A1(n8726), .A2(n8350), .B1(n8348), .B2(n8728), .ZN(n7249)
         );
  AND2_X1 U9040 ( .A1(n7250), .A2(n7249), .ZN(n10031) );
  MUX2_X1 U9041 ( .A(n10031), .B(n7251), .S(n8752), .Z(n7255) );
  INV_X1 U9042 ( .A(n7252), .ZN(n7253) );
  AOI22_X1 U9043 ( .A1(n8708), .A2(n10028), .B1(n8718), .B2(n7253), .ZN(n7254)
         );
  OAI211_X1 U9044 ( .C1(n8711), .C2(n10027), .A(n7255), .B(n7254), .ZN(
        P2_U3227) );
  INV_X1 U9045 ( .A(n7256), .ZN(n7257) );
  AOI21_X1 U9046 ( .B1(n7259), .B2(n7258), .A(n7257), .ZN(n7267) );
  NOR2_X1 U9047 ( .A1(n9043), .A2(n7623), .ZN(n7260) );
  AOI211_X1 U9048 ( .C1(n9045), .C2(n9321), .A(n7261), .B(n7260), .ZN(n7262)
         );
  OAI21_X1 U9049 ( .B1(n9048), .B2(n7263), .A(n7262), .ZN(n7264) );
  AOI21_X1 U9050 ( .B1(n7265), .B2(n9050), .A(n7264), .ZN(n7266) );
  OAI21_X1 U9051 ( .B1(n7267), .B2(n9052), .A(n7266), .ZN(P1_U3239) );
  INV_X1 U9052 ( .A(n7268), .ZN(n7870) );
  OAI222_X1 U9053 ( .A1(P2_U3151), .A2(n8519), .B1(n8900), .B2(n7870), .C1(
        n8899), .C2(n7269), .ZN(P2_U3276) );
  INV_X1 U9054 ( .A(n7363), .ZN(n7281) );
  OAI21_X1 U9055 ( .B1(n7275), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7270), .ZN(
        n7272) );
  MUX2_X1 U9056 ( .A(n5365), .B(P1_REG1_REG_13__SCAN_IN), .S(n7363), .Z(n7271)
         );
  NOR2_X1 U9057 ( .A1(n7272), .A2(n7271), .ZN(n7362) );
  AOI211_X1 U9058 ( .C1(n7272), .C2(n7271), .A(n9446), .B(n7362), .ZN(n7273)
         );
  INV_X1 U9059 ( .A(n7273), .ZN(n7280) );
  AND2_X1 U9060 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7794) );
  NAND2_X1 U9061 ( .A1(n7363), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7364) );
  OAI21_X1 U9062 ( .B1(n7363), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7364), .ZN(
        n7277) );
  OAI21_X1 U9063 ( .B1(n7275), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7274), .ZN(
        n7276) );
  NOR2_X1 U9064 ( .A1(n7276), .A2(n7277), .ZN(n7366) );
  AOI211_X1 U9065 ( .C1(n7277), .C2(n7276), .A(n7366), .B(n9428), .ZN(n7278)
         );
  AOI211_X1 U9066 ( .C1(n9433), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n7794), .B(
        n7278), .ZN(n7279) );
  OAI211_X1 U9067 ( .C1(n9445), .C2(n7281), .A(n7280), .B(n7279), .ZN(P1_U3256) );
  INV_X1 U9068 ( .A(n7282), .ZN(n7283) );
  NAND2_X1 U9069 ( .A1(n7284), .A2(n7283), .ZN(n7285) );
  XNOR2_X1 U9070 ( .A(n7658), .B(n7943), .ZN(n7557) );
  XNOR2_X1 U9071 ( .A(n7557), .B(n8347), .ZN(n7554) );
  XOR2_X1 U9072 ( .A(n7555), .B(n7554), .Z(n7295) );
  INV_X1 U9073 ( .A(n7287), .ZN(n7657) );
  NAND2_X1 U9074 ( .A1(n8113), .A2(n7657), .ZN(n7291) );
  INV_X1 U9075 ( .A(n7288), .ZN(n7289) );
  AOI21_X1 U9076 ( .B1(n4427), .B2(n8348), .A(n7289), .ZN(n7290) );
  OAI211_X1 U9077 ( .C1(n7292), .C2(n8110), .A(n7291), .B(n7290), .ZN(n7293)
         );
  AOI21_X1 U9078 ( .B1(n8037), .B2(n7658), .A(n7293), .ZN(n7294) );
  OAI21_X1 U9079 ( .B1(n7295), .B2(n8039), .A(n7294), .ZN(P2_U3161) );
  NAND2_X1 U9080 ( .A1(n7297), .A2(n7296), .ZN(n7298) );
  XNOR2_X1 U9081 ( .A(n7298), .B(n7306), .ZN(n9867) );
  NAND2_X1 U9082 ( .A1(n9598), .A2(n9918), .ZN(n9602) );
  INV_X1 U9083 ( .A(n9602), .ZN(n7807) );
  AOI22_X1 U9084 ( .A1(n9857), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9820), .ZN(n7299) );
  OAI21_X1 U9085 ( .B1(n9618), .B2(n7300), .A(n7299), .ZN(n7305) );
  INV_X1 U9086 ( .A(n7301), .ZN(n9839) );
  AOI211_X1 U9087 ( .C1(n9865), .C2(n7302), .A(n9822), .B(n9839), .ZN(n9863)
         );
  INV_X1 U9088 ( .A(n9863), .ZN(n7303) );
  OAI22_X1 U9089 ( .A1(n7303), .A2(n9606), .B1(n9879), .B2(n7809), .ZN(n7304)
         );
  AOI211_X1 U9090 ( .C1(n7807), .C2(n9323), .A(n7305), .B(n7304), .ZN(n7309)
         );
  XNOR2_X1 U9091 ( .A(n7307), .B(n7306), .ZN(n9869) );
  NOR2_X1 U9092 ( .A1(n9857), .A2(n9933), .ZN(n7902) );
  NAND2_X1 U9093 ( .A1(n9869), .A2(n7902), .ZN(n7308) );
  OAI211_X1 U9094 ( .C1(n9629), .C2(n9867), .A(n7309), .B(n7308), .ZN(P1_U3291) );
  XOR2_X1 U9095 ( .A(n7310), .B(n9082), .Z(n9884) );
  XOR2_X1 U9096 ( .A(n9082), .B(n4540), .Z(n9886) );
  NAND2_X1 U9097 ( .A1(n9886), .A2(n7902), .ZN(n7320) );
  OAI211_X1 U9098 ( .C1(n9836), .C2(n7316), .A(n7311), .B(n9837), .ZN(n9882)
         );
  INV_X1 U9099 ( .A(n9882), .ZN(n7318) );
  AOI22_X1 U9100 ( .A1(n7807), .A2(n9322), .B1(n9600), .B2(n9321), .ZN(n7315)
         );
  INV_X1 U9101 ( .A(n7312), .ZN(n7313) );
  AOI22_X1 U9102 ( .A1(n9857), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7313), .B2(
        n9820), .ZN(n7314) );
  OAI211_X1 U9103 ( .C1(n7316), .C2(n9618), .A(n7315), .B(n7314), .ZN(n7317)
         );
  AOI21_X1 U9104 ( .B1(n9851), .B2(n7318), .A(n7317), .ZN(n7319) );
  OAI211_X1 U9105 ( .C1(n9629), .C2(n9884), .A(n7320), .B(n7319), .ZN(P1_U3289) );
  INV_X1 U9106 ( .A(n7321), .ZN(n7347) );
  OAI222_X1 U9107 ( .A1(n9769), .A2(n7347), .B1(P1_U3086), .B2(n9298), .C1(
        n7322), .C2(n9771), .ZN(P1_U3335) );
  INV_X1 U9108 ( .A(n9138), .ZN(n9813) );
  NAND2_X1 U9109 ( .A1(n9809), .A2(n9813), .ZN(n9808) );
  NAND2_X1 U9110 ( .A1(n9808), .A2(n7324), .ZN(n7376) );
  NAND2_X1 U9111 ( .A1(n7376), .A2(n9136), .ZN(n7325) );
  XOR2_X1 U9112 ( .A(n7332), .B(n7325), .Z(n9922) );
  INV_X1 U9113 ( .A(n7902), .ZN(n9612) );
  AOI21_X1 U9114 ( .B1(n7385), .B2(n9919), .A(n9822), .ZN(n7326) );
  AOI22_X1 U9115 ( .A1(n7326), .A2(n4467), .B1(n9891), .B2(n9318), .ZN(n9921)
         );
  INV_X1 U9116 ( .A(n9921), .ZN(n7330) );
  INV_X1 U9117 ( .A(n9919), .ZN(n7702) );
  OAI22_X1 U9118 ( .A1(n9598), .A2(n6698), .B1(n7695), .B2(n9846), .ZN(n7327)
         );
  AOI21_X1 U9119 ( .B1(n7807), .B2(n9917), .A(n7327), .ZN(n7328) );
  OAI21_X1 U9120 ( .B1(n7702), .B2(n9618), .A(n7328), .ZN(n7329) );
  AOI21_X1 U9121 ( .B1(n7330), .B2(n9851), .A(n7329), .ZN(n7334) );
  XNOR2_X1 U9122 ( .A(n7331), .B(n7332), .ZN(n9924) );
  NAND2_X1 U9123 ( .A1(n9924), .A2(n9841), .ZN(n7333) );
  OAI211_X1 U9124 ( .C1(n9922), .C2(n9612), .A(n7334), .B(n7333), .ZN(P1_U3284) );
  INV_X1 U9125 ( .A(n7335), .ZN(n7336) );
  AOI21_X1 U9126 ( .B1(n7343), .B2(n7337), .A(n7336), .ZN(n9932) );
  AOI211_X1 U9127 ( .C1(n9930), .C2(n4467), .A(n9822), .B(n9804), .ZN(n9928)
         );
  NAND2_X1 U9128 ( .A1(n9930), .A2(n7133), .ZN(n7341) );
  OAI22_X1 U9129 ( .A1(n9598), .A2(n7338), .B1(n7776), .B2(n9846), .ZN(n7339)
         );
  AOI21_X1 U9130 ( .B1(n7807), .B2(n9319), .A(n7339), .ZN(n7340) );
  OAI211_X1 U9131 ( .C1(n9926), .C2(n7809), .A(n7341), .B(n7340), .ZN(n7342)
         );
  AOI21_X1 U9132 ( .B1(n9928), .B2(n9851), .A(n7342), .ZN(n7346) );
  XNOR2_X1 U9133 ( .A(n7344), .B(n7343), .ZN(n9935) );
  NAND2_X1 U9134 ( .A1(n9935), .A2(n9841), .ZN(n7345) );
  OAI211_X1 U9135 ( .C1(n9932), .C2(n9612), .A(n7346), .B(n7345), .ZN(P1_U3283) );
  OAI222_X1 U9136 ( .A1(P2_U3151), .A2(n8144), .B1(n8899), .B2(n6314), .C1(
        n7347), .C2(n8900), .ZN(P2_U3275) );
  XNOR2_X1 U9137 ( .A(n7349), .B(n4450), .ZN(n7350) );
  XNOR2_X1 U9138 ( .A(n7348), .B(n7350), .ZN(n7356) );
  NOR2_X1 U9139 ( .A1(n9043), .A2(n9810), .ZN(n7351) );
  AOI211_X1 U9140 ( .C1(n9045), .C2(n9890), .A(n7352), .B(n7351), .ZN(n7353)
         );
  OAI21_X1 U9141 ( .B1(n9048), .B2(n9818), .A(n7353), .ZN(n7354) );
  AOI21_X1 U9142 ( .B1(n9904), .B2(n9050), .A(n7354), .ZN(n7355) );
  OAI21_X1 U9143 ( .B1(n7356), .B2(n9052), .A(n7355), .ZN(P1_U3213) );
  INV_X1 U9144 ( .A(n7357), .ZN(n7360) );
  OAI222_X1 U9145 ( .A1(n9769), .A2(n7360), .B1(P1_U3086), .B2(n9236), .C1(
        n7358), .C2(n9771), .ZN(P1_U3334) );
  OAI222_X1 U9146 ( .A1(n8899), .A2(n7361), .B1(n8900), .B2(n7360), .C1(n7359), 
        .C2(P2_U3151), .ZN(P2_U3274) );
  MUX2_X1 U9147 ( .A(n5386), .B(P1_REG1_REG_14__SCAN_IN), .S(n7607), .Z(n7610)
         );
  AOI21_X1 U9148 ( .B1(n7363), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7362), .ZN(
        n7609) );
  XOR2_X1 U9149 ( .A(n7610), .B(n7609), .Z(n7373) );
  INV_X1 U9150 ( .A(n7364), .ZN(n7365) );
  NAND2_X1 U9151 ( .A1(n7607), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7367) );
  OAI21_X1 U9152 ( .B1(n7607), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7367), .ZN(
        n7368) );
  NOR2_X1 U9153 ( .A1(n7369), .A2(n7368), .ZN(n7606) );
  AOI211_X1 U9154 ( .C1(n7369), .C2(n7368), .A(n7606), .B(n9428), .ZN(n7372)
         );
  NOR2_X1 U9155 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10279), .ZN(n8909) );
  AOI21_X1 U9156 ( .B1(n9433), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n8909), .ZN(
        n7370) );
  OAI21_X1 U9157 ( .B1(n7612), .B2(n9445), .A(n7370), .ZN(n7371) );
  AOI211_X1 U9158 ( .C1(n7373), .C2(n9443), .A(n7372), .B(n7371), .ZN(n7374)
         );
  INV_X1 U9159 ( .A(n7374), .ZN(P1_U3257) );
  XNOR2_X1 U9160 ( .A(n7375), .B(n7377), .ZN(n9915) );
  OAI22_X1 U9161 ( .A1(n7623), .A2(n9952), .B1(n9927), .B2(n9950), .ZN(n7383)
         );
  INV_X1 U9162 ( .A(n7376), .ZN(n7381) );
  INV_X1 U9163 ( .A(n7377), .ZN(n7378) );
  AOI21_X1 U9164 ( .B1(n9808), .B2(n7379), .A(n7378), .ZN(n7380) );
  AOI211_X1 U9165 ( .C1(n7381), .C2(n9136), .A(n9933), .B(n7380), .ZN(n7382)
         );
  AOI211_X1 U9166 ( .C1(n9964), .C2(n9915), .A(n7383), .B(n7382), .ZN(n9912)
         );
  INV_X1 U9167 ( .A(n7384), .ZN(n9852) );
  OAI211_X1 U9168 ( .C1(n9821), .C2(n9911), .A(n7385), .B(n9837), .ZN(n9910)
         );
  INV_X1 U9169 ( .A(n7386), .ZN(n7627) );
  AOI22_X1 U9170 ( .A1(n9857), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7627), .B2(
        n9820), .ZN(n7389) );
  NAND2_X1 U9171 ( .A1(n7387), .A2(n7133), .ZN(n7388) );
  OAI211_X1 U9172 ( .C1(n9910), .C2(n9606), .A(n7389), .B(n7388), .ZN(n7390)
         );
  AOI21_X1 U9173 ( .B1(n9915), .B2(n9852), .A(n7390), .ZN(n7391) );
  OAI21_X1 U9174 ( .B1(n9912), .B2(n9857), .A(n7391), .ZN(P1_U3285) );
  XNOR2_X1 U9175 ( .A(n7426), .B(n7427), .ZN(n7394) );
  AOI21_X1 U9176 ( .B1(n6168), .B2(n7394), .A(n7428), .ZN(n7411) );
  MUX2_X1 U9177 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n4446), .Z(n7418) );
  XNOR2_X1 U9178 ( .A(n7418), .B(n7427), .ZN(n7399) );
  OR2_X1 U9179 ( .A1(n7395), .A2(n7402), .ZN(n7397) );
  NAND2_X1 U9180 ( .A1(n7397), .A2(n7396), .ZN(n7398) );
  OAI21_X1 U9181 ( .B1(n7399), .B2(n7398), .A(n7420), .ZN(n7400) );
  AND2_X1 U9182 ( .A1(n7400), .A2(n10406), .ZN(n7409) );
  INV_X1 U9183 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7407) );
  AND2_X1 U9184 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7551) );
  INV_X1 U9185 ( .A(n7551), .ZN(n7406) );
  AND2_X1 U9186 ( .A1(n7403), .A2(n6173), .ZN(n7404) );
  OAI21_X1 U9187 ( .B1(n7413), .B2(n7404), .A(n10419), .ZN(n7405) );
  OAI211_X1 U9188 ( .C1(n10005), .C2(n7407), .A(n7406), .B(n7405), .ZN(n7408)
         );
  AOI211_X1 U9189 ( .C1(n10411), .C2(n7427), .A(n7409), .B(n7408), .ZN(n7410)
         );
  OAI21_X1 U9190 ( .B1(n7411), .B2(n9985), .A(n7410), .ZN(P2_U3191) );
  NOR2_X1 U9191 ( .A1(n7427), .A2(n7412), .ZN(n7414) );
  OR2_X1 U9192 ( .A1(n7431), .A2(n7639), .ZN(n7530) );
  NAND2_X1 U9193 ( .A1(n7431), .A2(n7639), .ZN(n7415) );
  NAND2_X1 U9194 ( .A1(n7530), .A2(n7415), .ZN(n7416) );
  AOI21_X1 U9195 ( .B1(n7417), .B2(n7416), .A(n4449), .ZN(n7440) );
  MUX2_X1 U9196 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n4446), .Z(n7533) );
  XNOR2_X1 U9197 ( .A(n7533), .B(n7431), .ZN(n7423) );
  INV_X1 U9198 ( .A(n7418), .ZN(n7419) );
  NAND2_X1 U9199 ( .A1(n7427), .A2(n7419), .ZN(n7421) );
  NAND2_X1 U9200 ( .A1(n7421), .A2(n7420), .ZN(n7422) );
  NAND2_X1 U9201 ( .A1(n7423), .A2(n7422), .ZN(n7534) );
  OAI21_X1 U9202 ( .B1(n7423), .B2(n7422), .A(n7534), .ZN(n7438) );
  INV_X1 U9203 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10248) );
  NAND2_X1 U9204 ( .A1(n10411), .A2(n7431), .ZN(n7425) );
  AND2_X1 U9205 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7600) );
  INV_X1 U9206 ( .A(n7600), .ZN(n7424) );
  OAI211_X1 U9207 ( .C1(n10248), .C2(n10005), .A(n7425), .B(n7424), .ZN(n7437)
         );
  NOR2_X1 U9208 ( .A1(n7427), .A2(n7426), .ZN(n7429) );
  OR2_X1 U9209 ( .A1(n7431), .A2(n7430), .ZN(n7541) );
  NAND2_X1 U9210 ( .A1(n7431), .A2(n7430), .ZN(n7432) );
  NAND2_X1 U9211 ( .A1(n7541), .A2(n7432), .ZN(n7433) );
  NAND2_X1 U9212 ( .A1(n7434), .A2(n7433), .ZN(n7435) );
  AOI21_X1 U9213 ( .B1(n7542), .B2(n7435), .A(n9985), .ZN(n7436) );
  AOI211_X1 U9214 ( .C1(n10406), .C2(n7438), .A(n7437), .B(n7436), .ZN(n7439)
         );
  OAI21_X1 U9215 ( .B1(n7440), .B2(n10002), .A(n7439), .ZN(P2_U3192) );
  OR2_X1 U9216 ( .A1(n7441), .A2(n8311), .ZN(n7653) );
  INV_X1 U9217 ( .A(n7653), .ZN(n7442) );
  AOI21_X1 U9218 ( .B1(n8311), .B2(n7441), .A(n7442), .ZN(n7443) );
  OAI222_X1 U9219 ( .A1(n8742), .A2(n7444), .B1(n8744), .B2(n7556), .C1(n8740), 
        .C2(n7443), .ZN(n7512) );
  INV_X1 U9220 ( .A(n7512), .ZN(n7450) );
  XOR2_X1 U9221 ( .A(n7445), .B(n8311), .Z(n7513) );
  NOR2_X1 U9222 ( .A1(n8720), .A2(n7515), .ZN(n7448) );
  OAI22_X1 U9223 ( .A1(n8748), .A2(n7071), .B1(n7446), .B2(n8745), .ZN(n7447)
         );
  AOI211_X1 U9224 ( .C1(n7513), .C2(n8753), .A(n7448), .B(n7447), .ZN(n7449)
         );
  OAI21_X1 U9225 ( .B1(n7450), .B2(n8752), .A(n7449), .ZN(P2_U3226) );
  INV_X1 U9226 ( .A(n7451), .ZN(n7454) );
  OAI222_X1 U9227 ( .A1(n9771), .A2(n7452), .B1(n9769), .B2(n7454), .C1(n5691), 
        .C2(P1_U3086), .ZN(P1_U3333) );
  OAI222_X1 U9228 ( .A1(n8899), .A2(n10269), .B1(n8900), .B2(n7454), .C1(
        P2_U3151), .C2(n7453), .ZN(P2_U3273) );
  INV_X1 U9229 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10082) );
  NOR2_X1 U9230 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7495) );
  NOR2_X1 U9231 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7492) );
  NOR2_X1 U9232 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7489) );
  NOR2_X1 U9233 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7486) );
  NOR2_X1 U9234 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7482) );
  NOR2_X1 U9235 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7480) );
  XNOR2_X1 U9236 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10095) );
  NAND2_X1 U9237 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7478) );
  INV_X1 U9238 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7540) );
  XNOR2_X1 U9239 ( .A(P1_ADDR_REG_11__SCAN_IN), .B(n7540), .ZN(n10097) );
  NAND2_X1 U9240 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7476) );
  XNOR2_X1 U9241 ( .A(n10248), .B(P1_ADDR_REG_10__SCAN_IN), .ZN(n10099) );
  NOR2_X1 U9242 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7460) );
  XOR2_X1 U9243 ( .A(n10391), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10436) );
  NAND2_X1 U9244 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7458) );
  XOR2_X1 U9245 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10434) );
  NAND2_X1 U9246 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7456) );
  XOR2_X1 U9247 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10432) );
  AOI21_X1 U9248 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10076) );
  NAND3_X1 U9249 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10078) );
  OAI21_X1 U9250 ( .B1(n10076), .B2(n10251), .A(n10078), .ZN(n10431) );
  NAND2_X1 U9251 ( .A1(n10432), .A2(n10431), .ZN(n7455) );
  NAND2_X1 U9252 ( .A1(n7456), .A2(n7455), .ZN(n10433) );
  NAND2_X1 U9253 ( .A1(n10434), .A2(n10433), .ZN(n7457) );
  NAND2_X1 U9254 ( .A1(n7458), .A2(n7457), .ZN(n10435) );
  NOR2_X1 U9255 ( .A1(n10436), .A2(n10435), .ZN(n7459) );
  NOR2_X1 U9256 ( .A1(n7460), .A2(n7459), .ZN(n7461) );
  NOR2_X1 U9257 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7461), .ZN(n10426) );
  AND2_X1 U9258 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7461), .ZN(n10425) );
  NOR2_X1 U9259 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10425), .ZN(n7462) );
  NOR2_X1 U9260 ( .A1(n10426), .A2(n7462), .ZN(n7463) );
  NAND2_X1 U9261 ( .A1(n7463), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7465) );
  INV_X1 U9262 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10101) );
  XNOR2_X1 U9263 ( .A(n7463), .B(n10101), .ZN(n10424) );
  NAND2_X1 U9264 ( .A1(n10424), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7464) );
  NAND2_X1 U9265 ( .A1(n7465), .A2(n7464), .ZN(n7466) );
  NAND2_X1 U9266 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7466), .ZN(n7468) );
  INV_X1 U9267 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10176) );
  XNOR2_X1 U9268 ( .A(n10176), .B(n7466), .ZN(n10429) );
  NAND2_X1 U9269 ( .A1(n10429), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7467) );
  NAND2_X1 U9270 ( .A1(n7468), .A2(n7467), .ZN(n7469) );
  NAND2_X1 U9271 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7469), .ZN(n7471) );
  INV_X1 U9272 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10161) );
  XNOR2_X1 U9273 ( .A(n10161), .B(n7469), .ZN(n10430) );
  NAND2_X1 U9274 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10430), .ZN(n7470) );
  NAND2_X1 U9275 ( .A1(n7471), .A2(n7470), .ZN(n7472) );
  NAND2_X1 U9276 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n7472), .ZN(n7474) );
  XOR2_X1 U9277 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n7472), .Z(n10428) );
  NAND2_X1 U9278 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10428), .ZN(n7473) );
  NAND2_X1 U9279 ( .A1(n7474), .A2(n7473), .ZN(n10098) );
  NAND2_X1 U9280 ( .A1(n10099), .A2(n10098), .ZN(n7475) );
  NAND2_X1 U9281 ( .A1(n7476), .A2(n7475), .ZN(n10096) );
  NAND2_X1 U9282 ( .A1(n10097), .A2(n10096), .ZN(n7477) );
  NAND2_X1 U9283 ( .A1(n7478), .A2(n7477), .ZN(n10094) );
  NOR2_X1 U9284 ( .A1(n10095), .A2(n10094), .ZN(n7479) );
  NOR2_X1 U9285 ( .A1(n7480), .A2(n7479), .ZN(n10093) );
  INV_X1 U9286 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10206) );
  INV_X1 U9287 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10294) );
  AOI22_X1 U9288 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n10206), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n10294), .ZN(n10092) );
  NOR2_X1 U9289 ( .A1(n10093), .A2(n10092), .ZN(n7481) );
  NOR2_X1 U9290 ( .A1(n7482), .A2(n7481), .ZN(n10091) );
  INV_X1 U9291 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7484) );
  INV_X1 U9292 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7483) );
  AOI22_X1 U9293 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n7484), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(n7483), .ZN(n10090) );
  NOR2_X1 U9294 ( .A1(n10091), .A2(n10090), .ZN(n7485) );
  NOR2_X1 U9295 ( .A1(n7486), .A2(n7485), .ZN(n10089) );
  INV_X1 U9296 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7487) );
  INV_X1 U9297 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8425) );
  AOI22_X1 U9298 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n7487), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n8425), .ZN(n10088) );
  NOR2_X1 U9299 ( .A1(n10089), .A2(n10088), .ZN(n7488) );
  NOR2_X1 U9300 ( .A1(n7489), .A2(n7488), .ZN(n10087) );
  INV_X1 U9301 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7490) );
  INV_X1 U9302 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8451) );
  AOI22_X1 U9303 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n7490), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n8451), .ZN(n10086) );
  NOR2_X1 U9304 ( .A1(n10087), .A2(n10086), .ZN(n7491) );
  NOR2_X1 U9305 ( .A1(n7492), .A2(n7491), .ZN(n10085) );
  INV_X1 U9306 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7493) );
  INV_X1 U9307 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8478) );
  AOI22_X1 U9308 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n7493), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n8478), .ZN(n10084) );
  NOR2_X1 U9309 ( .A1(n10085), .A2(n10084), .ZN(n7494) );
  NOR2_X1 U9310 ( .A1(n7495), .A2(n7494), .ZN(n10081) );
  NOR2_X1 U9311 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10081), .ZN(n7496) );
  NAND2_X1 U9312 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10081), .ZN(n10080) );
  OAI21_X1 U9313 ( .B1(n10082), .B2(n7496), .A(n10080), .ZN(n7498) );
  XNOR2_X1 U9314 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7497) );
  XNOR2_X1 U9315 ( .A(n7498), .B(n7497), .ZN(ADD_1068_U4) );
  XNOR2_X1 U9316 ( .A(n7499), .B(n5351), .ZN(n7523) );
  INV_X1 U9317 ( .A(n7523), .ZN(n7511) );
  OAI211_X1 U9318 ( .C1(n7501), .C2(n5351), .A(n7500), .B(n9887), .ZN(n7503)
         );
  OR2_X1 U9319 ( .A1(n9926), .A2(n9952), .ZN(n7502) );
  OAI211_X1 U9320 ( .C1(n9953), .C2(n9950), .A(n7503), .B(n7502), .ZN(n7521)
         );
  INV_X1 U9321 ( .A(n7504), .ZN(n9803) );
  INV_X1 U9322 ( .A(n7505), .ZN(n7666) );
  AOI211_X1 U9323 ( .C1(n7527), .C2(n9803), .A(n9822), .B(n7666), .ZN(n7522)
         );
  NAND2_X1 U9324 ( .A1(n7522), .A2(n9851), .ZN(n7508) );
  INV_X1 U9325 ( .A(n7506), .ZN(n8956) );
  AOI22_X1 U9326 ( .A1(n9857), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8956), .B2(
        n9820), .ZN(n7507) );
  OAI211_X1 U9327 ( .C1(n8959), .C2(n9618), .A(n7508), .B(n7507), .ZN(n7509)
         );
  AOI21_X1 U9328 ( .B1(n9598), .B2(n7521), .A(n7509), .ZN(n7510) );
  OAI21_X1 U9329 ( .B1(n7511), .B2(n9629), .A(n7510), .ZN(P1_U3281) );
  AOI21_X1 U9330 ( .B1(n10020), .B2(n7513), .A(n7512), .ZN(n7520) );
  INV_X1 U9331 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7514) );
  OAI22_X1 U9332 ( .A1(n7515), .A2(n8864), .B1(n10064), .B2(n7514), .ZN(n7516)
         );
  INV_X1 U9333 ( .A(n7516), .ZN(n7517) );
  OAI21_X1 U9334 ( .B1(n7520), .B2(n10062), .A(n7517), .ZN(P2_U3411) );
  AOI22_X1 U9335 ( .A1(n8808), .A2(n7518), .B1(n6533), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n7519) );
  OAI21_X1 U9336 ( .B1(n7520), .B2(n6533), .A(n7519), .ZN(P2_U3466) );
  AOI211_X1 U9337 ( .C1(n7523), .C2(n9949), .A(n7522), .B(n7521), .ZN(n7529)
         );
  INV_X1 U9338 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7524) );
  OAI22_X1 U9339 ( .A1(n8959), .A2(n9754), .B1(n9967), .B2(n7524), .ZN(n7525)
         );
  INV_X1 U9340 ( .A(n7525), .ZN(n7526) );
  OAI21_X1 U9341 ( .B1(n7529), .B2(n9965), .A(n7526), .ZN(P1_U3489) );
  AOI22_X1 U9342 ( .A1(n7527), .A2(n9673), .B1(n9981), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7528) );
  OAI21_X1 U9343 ( .B1(n7529), .B2(n9981), .A(n7528), .ZN(P1_U3534) );
  AOI21_X1 U9344 ( .B1(n7531), .B2(n7711), .A(n7567), .ZN(n7549) );
  MUX2_X1 U9345 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n4446), .Z(n7572) );
  XNOR2_X1 U9346 ( .A(n7572), .B(n7581), .ZN(n7537) );
  OR2_X1 U9347 ( .A1(n7533), .A2(n7532), .ZN(n7535) );
  NAND2_X1 U9348 ( .A1(n7535), .A2(n7534), .ZN(n7536) );
  NAND2_X1 U9349 ( .A1(n7537), .A2(n7536), .ZN(n7573) );
  OAI21_X1 U9350 ( .B1(n7537), .B2(n7536), .A(n7573), .ZN(n7547) );
  NAND2_X1 U9351 ( .A1(n10411), .A2(n7581), .ZN(n7539) );
  AND2_X1 U9352 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7749) );
  INV_X1 U9353 ( .A(n7749), .ZN(n7538) );
  OAI211_X1 U9354 ( .C1(n7540), .C2(n10005), .A(n7539), .B(n7538), .ZN(n7546)
         );
  AOI21_X1 U9355 ( .B1(n6198), .B2(n7543), .A(n7582), .ZN(n7544) );
  NOR2_X1 U9356 ( .A1(n7544), .A2(n9985), .ZN(n7545) );
  AOI211_X1 U9357 ( .C1(n10406), .C2(n7547), .A(n7546), .B(n7545), .ZN(n7548)
         );
  OAI21_X1 U9358 ( .B1(n7549), .B2(n10002), .A(n7548), .ZN(P2_U3193) );
  INV_X1 U9359 ( .A(n7550), .ZN(n7687) );
  NAND2_X1 U9360 ( .A1(n8113), .A2(n7687), .ZN(n7553) );
  AOI21_X1 U9361 ( .B1(n4427), .B2(n8347), .A(n7551), .ZN(n7552) );
  OAI211_X1 U9362 ( .C1(n7708), .C2(n8110), .A(n7553), .B(n7552), .ZN(n7564)
         );
  XNOR2_X1 U9363 ( .A(n7688), .B(n7938), .ZN(n7595) );
  XNOR2_X1 U9364 ( .A(n7595), .B(n8346), .ZN(n7562) );
  NAND2_X1 U9365 ( .A1(n7557), .A2(n7556), .ZN(n7558) );
  INV_X1 U9366 ( .A(n7597), .ZN(n7561) );
  AOI211_X1 U9367 ( .C1(n7562), .C2(n7559), .A(n8039), .B(n7561), .ZN(n7563)
         );
  AOI211_X1 U9368 ( .C1(n8037), .C2(n7688), .A(n7564), .B(n7563), .ZN(n7565)
         );
  INV_X1 U9369 ( .A(n7565), .ZN(P2_U3171) );
  NOR2_X1 U9370 ( .A1(n7581), .A2(n7566), .ZN(n7568) );
  AOI22_X1 U9371 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n7587), .B1(n8373), .B2(
        n6220), .ZN(n7569) );
  NOR2_X1 U9372 ( .A1(n7570), .A2(n7569), .ZN(n8372) );
  AOI21_X1 U9373 ( .B1(n7570), .B2(n7569), .A(n8372), .ZN(n7594) );
  OR2_X1 U9374 ( .A1(n7572), .A2(n7571), .ZN(n7574) );
  NAND2_X1 U9375 ( .A1(n7574), .A2(n7573), .ZN(n8362) );
  MUX2_X1 U9376 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n4446), .Z(n7575) );
  NOR2_X1 U9377 ( .A1(n7575), .A2(n8373), .ZN(n8361) );
  NAND2_X1 U9378 ( .A1(n7575), .A2(n8373), .ZN(n8363) );
  INV_X1 U9379 ( .A(n8363), .ZN(n7576) );
  NOR2_X1 U9380 ( .A1(n8361), .A2(n7576), .ZN(n7577) );
  XNOR2_X1 U9381 ( .A(n8362), .B(n7577), .ZN(n7578) );
  NAND2_X1 U9382 ( .A1(n7578), .A2(n10406), .ZN(n7593) );
  INV_X1 U9383 ( .A(n7579), .ZN(n7580) );
  NOR2_X1 U9384 ( .A1(n7581), .A2(n7580), .ZN(n7583) );
  AOI22_X1 U9385 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n7587), .B1(n8373), .B2(
        n8355), .ZN(n7584) );
  NOR2_X1 U9386 ( .A1(n7585), .A2(n7584), .ZN(n8357) );
  AOI21_X1 U9387 ( .B1(n7585), .B2(n7584), .A(n8357), .ZN(n7586) );
  INV_X1 U9388 ( .A(n7586), .ZN(n7591) );
  INV_X1 U9389 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7589) );
  NAND2_X1 U9390 ( .A1(n10411), .A2(n7587), .ZN(n7588) );
  NAND2_X1 U9391 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7766) );
  OAI211_X1 U9392 ( .C1(n10005), .C2(n7589), .A(n7588), .B(n7766), .ZN(n7590)
         );
  AOI21_X1 U9393 ( .B1(n7591), .B2(n10404), .A(n7590), .ZN(n7592) );
  OAI211_X1 U9394 ( .C1(n7594), .C2(n10002), .A(n7593), .B(n7592), .ZN(
        P2_U3194) );
  NAND2_X1 U9395 ( .A1(n7595), .A2(n8346), .ZN(n7596) );
  NAND2_X1 U9396 ( .A1(n7597), .A2(n7596), .ZN(n7752) );
  XOR2_X1 U9397 ( .A(n7943), .B(n10049), .Z(n7753) );
  XOR2_X1 U9398 ( .A(n7598), .B(n7753), .Z(n7605) );
  INV_X1 U9399 ( .A(n7638), .ZN(n7599) );
  NAND2_X1 U9400 ( .A1(n8113), .A2(n7599), .ZN(n7602) );
  AOI21_X1 U9401 ( .B1(n4427), .B2(n8346), .A(n7600), .ZN(n7601) );
  OAI211_X1 U9402 ( .C1(n7767), .C2(n8110), .A(n7602), .B(n7601), .ZN(n7603)
         );
  AOI21_X1 U9403 ( .B1(n8037), .B2(n10049), .A(n7603), .ZN(n7604) );
  OAI21_X1 U9404 ( .B1(n7605), .B2(n8039), .A(n7604), .ZN(P2_U3157) );
  XNOR2_X1 U9405 ( .A(n9387), .B(n9388), .ZN(n7608) );
  NOR2_X1 U9406 ( .A1(n7739), .A2(n7608), .ZN(n9389) );
  AOI211_X1 U9407 ( .C1(n7739), .C2(n7608), .A(n9389), .B(n9428), .ZN(n7618)
         );
  OR2_X1 U9408 ( .A1(n7610), .A2(n7609), .ZN(n7611) );
  OAI21_X1 U9409 ( .B1(n5386), .B2(n7612), .A(n7611), .ZN(n9380) );
  XNOR2_X1 U9410 ( .A(n9387), .B(n9380), .ZN(n7613) );
  NAND2_X1 U9411 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n7613), .ZN(n9382) );
  OAI211_X1 U9412 ( .C1(n7613), .C2(P1_REG1_REG_15__SCAN_IN), .A(n9443), .B(
        n9382), .ZN(n7616) );
  NAND2_X1 U9413 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9042) );
  INV_X1 U9414 ( .A(n9042), .ZN(n7614) );
  AOI21_X1 U9415 ( .B1(n9433), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n7614), .ZN(
        n7615) );
  OAI211_X1 U9416 ( .C1(n9445), .C2(n9387), .A(n7616), .B(n7615), .ZN(n7617)
         );
  OR2_X1 U9417 ( .A1(n7618), .A2(n7617), .ZN(P1_U3258) );
  OAI21_X1 U9418 ( .B1(n7621), .B2(n7620), .A(n7619), .ZN(n7622) );
  NAND2_X1 U9419 ( .A1(n7622), .A2(n9031), .ZN(n7629) );
  INV_X1 U9420 ( .A(n7623), .ZN(n9320) );
  AOI21_X1 U9421 ( .B1(n9045), .B2(n9320), .A(n7624), .ZN(n7625) );
  OAI21_X1 U9422 ( .B1(n9927), .B2(n9043), .A(n7625), .ZN(n7626) );
  AOI21_X1 U9423 ( .B1(n7627), .B2(n8991), .A(n7626), .ZN(n7628) );
  OAI211_X1 U9424 ( .C1(n9911), .C2(n9039), .A(n7629), .B(n7628), .ZN(P1_U3221) );
  NAND2_X1 U9425 ( .A1(n7630), .A2(n8147), .ZN(n7633) );
  NAND2_X1 U9426 ( .A1(n7631), .A2(n8163), .ZN(n8314) );
  INV_X1 U9427 ( .A(n8314), .ZN(n7632) );
  XNOR2_X1 U9428 ( .A(n7633), .B(n7632), .ZN(n10046) );
  XNOR2_X1 U9429 ( .A(n7634), .B(n8314), .ZN(n7635) );
  NAND2_X1 U9430 ( .A1(n7635), .A2(n8731), .ZN(n7637) );
  AOI22_X1 U9431 ( .A1(n8726), .A2(n8346), .B1(n8344), .B2(n8728), .ZN(n7636)
         );
  OAI211_X1 U9432 ( .C1(n10046), .C2(n7685), .A(n7637), .B(n7636), .ZN(n10047)
         );
  NAND2_X1 U9433 ( .A1(n10047), .A2(n8748), .ZN(n7642) );
  OAI22_X1 U9434 ( .A1(n8748), .A2(n7639), .B1(n7638), .B2(n8745), .ZN(n7640)
         );
  AOI21_X1 U9435 ( .B1(n8708), .B2(n10049), .A(n7640), .ZN(n7641) );
  OAI211_X1 U9436 ( .C1(n10046), .C2(n7963), .A(n7642), .B(n7641), .ZN(
        P2_U3223) );
  NAND2_X1 U9437 ( .A1(n7645), .A2(n9764), .ZN(n7643) );
  OAI211_X1 U9438 ( .C1(n7644), .C2(n9771), .A(n7643), .B(n9308), .ZN(P1_U3332) );
  NAND2_X1 U9439 ( .A1(n7645), .A2(n8897), .ZN(n7647) );
  INV_X1 U9440 ( .A(n7646), .ZN(n8339) );
  OAI211_X1 U9441 ( .C1(n7648), .C2(n8899), .A(n7647), .B(n8339), .ZN(P2_U3272) );
  NAND2_X1 U9442 ( .A1(n7650), .A2(n7649), .ZN(n8309) );
  XNOR2_X1 U9443 ( .A(n7651), .B(n8309), .ZN(n10035) );
  NAND2_X1 U9444 ( .A1(n7653), .A2(n7652), .ZN(n7654) );
  XOR2_X1 U9445 ( .A(n8309), .B(n7654), .Z(n7655) );
  AOI222_X1 U9446 ( .A1(n8731), .A2(n7655), .B1(n8346), .B2(n8728), .C1(n8348), 
        .C2(n8726), .ZN(n10033) );
  MUX2_X1 U9447 ( .A(n7656), .B(n10033), .S(n8748), .Z(n7660) );
  AOI22_X1 U9448 ( .A1(n8708), .A2(n7658), .B1(n8718), .B2(n7657), .ZN(n7659)
         );
  OAI211_X1 U9449 ( .C1(n8711), .C2(n10035), .A(n7660), .B(n7659), .ZN(
        P2_U3225) );
  OAI21_X1 U9450 ( .B1(n7661), .B2(n9091), .A(n7716), .ZN(n9948) );
  INV_X1 U9451 ( .A(n9948), .ZN(n7673) );
  INV_X1 U9452 ( .A(n7662), .ZN(n7663) );
  AOI21_X1 U9453 ( .B1(n9091), .B2(n7664), .A(n7663), .ZN(n7665) );
  OAI222_X1 U9454 ( .A1(n9950), .A2(n7829), .B1(n9952), .B2(n9793), .C1(n9933), 
        .C2(n7665), .ZN(n9946) );
  INV_X1 U9455 ( .A(n7668), .ZN(n9945) );
  OAI211_X1 U9456 ( .C1(n7666), .C2(n9945), .A(n9837), .B(n7718), .ZN(n9943)
         );
  INV_X1 U9457 ( .A(n7667), .ZN(n7797) );
  AOI22_X1 U9458 ( .A1(n9857), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7797), .B2(
        n9820), .ZN(n7670) );
  NAND2_X1 U9459 ( .A1(n7668), .A2(n7133), .ZN(n7669) );
  OAI211_X1 U9460 ( .C1(n9943), .C2(n9606), .A(n7670), .B(n7669), .ZN(n7671)
         );
  AOI21_X1 U9461 ( .B1(n9946), .B2(n9598), .A(n7671), .ZN(n7672) );
  OAI21_X1 U9462 ( .B1(n9629), .B2(n7673), .A(n7672), .ZN(P1_U3280) );
  NAND2_X1 U9463 ( .A1(n7674), .A2(n8315), .ZN(n7675) );
  NAND2_X1 U9464 ( .A1(n7630), .A2(n7675), .ZN(n10041) );
  OR2_X1 U9465 ( .A1(n7441), .A2(n7676), .ZN(n7678) );
  NAND2_X1 U9466 ( .A1(n7678), .A2(n7677), .ZN(n7679) );
  NOR2_X1 U9467 ( .A1(n7679), .A2(n8315), .ZN(n7680) );
  OR2_X1 U9468 ( .A1(n7681), .A2(n7680), .ZN(n7682) );
  NAND2_X1 U9469 ( .A1(n7682), .A2(n8731), .ZN(n7684) );
  AOI22_X1 U9470 ( .A1(n8726), .A2(n8347), .B1(n8345), .B2(n8728), .ZN(n7683)
         );
  OAI211_X1 U9471 ( .C1(n7685), .C2(n10041), .A(n7684), .B(n7683), .ZN(n10043)
         );
  MUX2_X1 U9472 ( .A(n10043), .B(P2_REG2_REG_9__SCAN_IN), .S(n8752), .Z(n7686)
         );
  INV_X1 U9473 ( .A(n7686), .ZN(n7690) );
  AOI22_X1 U9474 ( .A1(n8708), .A2(n7688), .B1(n8718), .B2(n7687), .ZN(n7689)
         );
  OAI211_X1 U9475 ( .C1(n10041), .C2(n7963), .A(n7690), .B(n7689), .ZN(
        P2_U3224) );
  AND2_X1 U9476 ( .A1(n7619), .A2(n7691), .ZN(n7694) );
  OAI211_X1 U9477 ( .C1(n7694), .C2(n7693), .A(n9031), .B(n7692), .ZN(n7701)
         );
  INV_X1 U9478 ( .A(n7695), .ZN(n7699) );
  AOI21_X1 U9479 ( .B1(n9045), .B2(n9917), .A(n7696), .ZN(n7697) );
  OAI21_X1 U9480 ( .B1(n9792), .B2(n9043), .A(n7697), .ZN(n7698) );
  AOI21_X1 U9481 ( .B1(n7699), .B2(n8991), .A(n7698), .ZN(n7700) );
  OAI211_X1 U9482 ( .C1(n7702), .C2(n9039), .A(n7701), .B(n7700), .ZN(P1_U3231) );
  INV_X1 U9483 ( .A(n7703), .ZN(n7869) );
  OAI222_X1 U9484 ( .A1(n9769), .A2(n7869), .B1(P1_U3086), .B2(n7704), .C1(
        n10162), .C2(n9771), .ZN(P1_U3331) );
  XOR2_X1 U9485 ( .A(n7705), .B(n8151), .Z(n10051) );
  AOI211_X1 U9486 ( .C1(n8151), .C2(n7707), .A(n8740), .B(n7706), .ZN(n7710)
         );
  OAI22_X1 U9487 ( .A1(n7708), .A2(n8742), .B1(n8741), .B2(n8744), .ZN(n7709)
         );
  OR2_X1 U9488 ( .A1(n7710), .A2(n7709), .ZN(n10052) );
  NAND2_X1 U9489 ( .A1(n10052), .A2(n8748), .ZN(n7714) );
  OAI22_X1 U9490 ( .A1(n8748), .A2(n7711), .B1(n7747), .B2(n8745), .ZN(n7712)
         );
  AOI21_X1 U9491 ( .B1(n10054), .B2(n8708), .A(n7712), .ZN(n7713) );
  OAI211_X1 U9492 ( .C1(n10051), .C2(n8711), .A(n7714), .B(n7713), .ZN(
        P2_U3222) );
  NAND2_X1 U9493 ( .A1(n7716), .A2(n7715), .ZN(n7717) );
  XOR2_X1 U9494 ( .A(n9166), .B(n7717), .Z(n9963) );
  INV_X1 U9495 ( .A(n9963), .ZN(n9961) );
  AOI211_X1 U9496 ( .C1(n9956), .C2(n7718), .A(n9822), .B(n7737), .ZN(n9954)
         );
  NAND2_X1 U9497 ( .A1(n9956), .A2(n7133), .ZN(n7722) );
  OAI22_X1 U9498 ( .A1(n9598), .A2(n7719), .B1(n8911), .B2(n9846), .ZN(n7720)
         );
  AOI21_X1 U9499 ( .B1(n7807), .B2(n9315), .A(n7720), .ZN(n7721) );
  OAI211_X1 U9500 ( .C1(n9951), .C2(n7809), .A(n7722), .B(n7721), .ZN(n7726)
         );
  OAI211_X1 U9501 ( .C1(n7724), .C2(n9166), .A(n9887), .B(n7723), .ZN(n9958)
         );
  NOR2_X1 U9502 ( .A1(n9958), .A2(n9857), .ZN(n7725) );
  AOI211_X1 U9503 ( .C1(n9954), .C2(n9851), .A(n7726), .B(n7725), .ZN(n7727)
         );
  OAI21_X1 U9504 ( .B1(n9961), .B2(n9629), .A(n7727), .ZN(P1_U3279) );
  INV_X1 U9505 ( .A(n7728), .ZN(n7759) );
  OAI222_X1 U9506 ( .A1(n9769), .A2(n7759), .B1(P1_U3086), .B2(n7730), .C1(
        n7729), .C2(n9771), .ZN(P1_U3330) );
  XNOR2_X1 U9507 ( .A(n7731), .B(n7732), .ZN(n7834) );
  INV_X1 U9508 ( .A(n7723), .ZN(n7734) );
  OAI21_X1 U9509 ( .B1(n7734), .B2(n7733), .A(n7732), .ZN(n7736) );
  NAND2_X1 U9510 ( .A1(n7736), .A2(n7735), .ZN(n7832) );
  INV_X1 U9511 ( .A(n7737), .ZN(n7738) );
  AOI211_X1 U9512 ( .C1(n9151), .C2(n7738), .A(n9822), .B(n7810), .ZN(n7831)
         );
  NAND2_X1 U9513 ( .A1(n7831), .A2(n9851), .ZN(n7744) );
  OAI22_X1 U9514 ( .A1(n9598), .A2(n7739), .B1(n9047), .B2(n9846), .ZN(n7741)
         );
  NOR2_X1 U9515 ( .A1(n9602), .A2(n7829), .ZN(n7740) );
  AOI211_X1 U9516 ( .C1(n9600), .C2(n7742), .A(n7741), .B(n7740), .ZN(n7743)
         );
  OAI211_X1 U9517 ( .C1(n7840), .C2(n9618), .A(n7744), .B(n7743), .ZN(n7745)
         );
  AOI21_X1 U9518 ( .B1(n7832), .B2(n7902), .A(n7745), .ZN(n7746) );
  OAI21_X1 U9519 ( .B1(n7834), .B2(n9629), .A(n7746), .ZN(P1_U3278) );
  INV_X1 U9520 ( .A(n7747), .ZN(n7748) );
  NAND2_X1 U9521 ( .A1(n8113), .A2(n7748), .ZN(n7751) );
  AOI21_X1 U9522 ( .B1(n4427), .B2(n8345), .A(n7749), .ZN(n7750) );
  OAI211_X1 U9523 ( .C1(n8741), .C2(n8110), .A(n7751), .B(n7750), .ZN(n7756)
         );
  XOR2_X1 U9524 ( .A(n7943), .B(n8151), .Z(n7760) );
  NOR2_X1 U9525 ( .A1(n7754), .A2(n7760), .ZN(n7762) );
  AOI211_X1 U9526 ( .C1(n7760), .C2(n7754), .A(n8039), .B(n7762), .ZN(n7755)
         );
  AOI211_X1 U9527 ( .C1(n8037), .C2(n10054), .A(n7756), .B(n7755), .ZN(n7757)
         );
  INV_X1 U9528 ( .A(n7757), .ZN(P2_U3176) );
  OAI222_X1 U9529 ( .A1(n8899), .A2(n10115), .B1(n8900), .B2(n7759), .C1(n7758), .C2(P2_U3151), .ZN(P2_U3270) );
  INV_X1 U9530 ( .A(n10060), .ZN(n7772) );
  AND2_X1 U9531 ( .A1(n7760), .A2(n8344), .ZN(n7761) );
  NOR2_X1 U9532 ( .A1(n7762), .A2(n7761), .ZN(n7764) );
  XNOR2_X1 U9533 ( .A(n10060), .B(n7943), .ZN(n7817) );
  XNOR2_X1 U9534 ( .A(n7817), .B(n8343), .ZN(n7763) );
  NAND2_X1 U9535 ( .A1(n7764), .A2(n7763), .ZN(n7819) );
  OAI21_X1 U9536 ( .B1(n7764), .B2(n7763), .A(n7819), .ZN(n7765) );
  NAND2_X1 U9537 ( .A1(n7765), .A2(n8104), .ZN(n7771) );
  OAI21_X1 U9538 ( .B1(n8068), .B2(n7767), .A(n7766), .ZN(n7769) );
  NOR2_X1 U9539 ( .A1(n8044), .A2(n7784), .ZN(n7768) );
  AOI211_X1 U9540 ( .C1(n8066), .C2(n8727), .A(n7769), .B(n7768), .ZN(n7770)
         );
  OAI211_X1 U9541 ( .C1(n7772), .C2(n8116), .A(n7771), .B(n7770), .ZN(P2_U3164) );
  XOR2_X1 U9542 ( .A(n7852), .B(n7853), .Z(n7856) );
  XNOR2_X1 U9543 ( .A(n7856), .B(n7855), .ZN(n7779) );
  NOR2_X1 U9544 ( .A1(n8983), .A2(n9927), .ZN(n7773) );
  AOI211_X1 U9545 ( .C1(n9036), .C2(n9317), .A(n7774), .B(n7773), .ZN(n7775)
         );
  OAI21_X1 U9546 ( .B1(n9048), .B2(n7776), .A(n7775), .ZN(n7777) );
  AOI21_X1 U9547 ( .B1(n9930), .B2(n9050), .A(n7777), .ZN(n7778) );
  OAI21_X1 U9548 ( .B1(n7779), .B2(n9052), .A(n7778), .ZN(P1_U3217) );
  OAI21_X1 U9549 ( .B1(n4536), .B2(n8152), .A(n7780), .ZN(n10057) );
  OAI21_X1 U9550 ( .B1(n7781), .B2(n6441), .A(n8731), .ZN(n7783) );
  AOI22_X1 U9551 ( .A1(n8726), .A2(n8344), .B1(n8727), .B2(n8728), .ZN(n7782)
         );
  OAI21_X1 U9552 ( .B1(n7783), .B2(n4535), .A(n7782), .ZN(n10058) );
  NAND2_X1 U9553 ( .A1(n10058), .A2(n8748), .ZN(n7787) );
  OAI22_X1 U9554 ( .A1(n8748), .A2(n6220), .B1(n7784), .B2(n8745), .ZN(n7785)
         );
  AOI21_X1 U9555 ( .B1(n10060), .B2(n8708), .A(n7785), .ZN(n7786) );
  OAI211_X1 U9556 ( .C1(n8711), .C2(n10057), .A(n7787), .B(n7786), .ZN(
        P2_U3221) );
  INV_X1 U9557 ( .A(n7788), .ZN(n8951) );
  NOR3_X1 U9558 ( .A1(n8951), .A2(n4973), .A3(n7790), .ZN(n7793) );
  INV_X1 U9559 ( .A(n7791), .ZN(n7792) );
  OAI21_X1 U9560 ( .B1(n7793), .B2(n7792), .A(n9031), .ZN(n7799) );
  AOI21_X1 U9561 ( .B1(n9045), .B2(n9316), .A(n7794), .ZN(n7795) );
  OAI21_X1 U9562 ( .B1(n7829), .B2(n9043), .A(n7795), .ZN(n7796) );
  AOI21_X1 U9563 ( .B1(n7797), .B2(n8991), .A(n7796), .ZN(n7798) );
  OAI211_X1 U9564 ( .C1(n9945), .C2(n9039), .A(n7799), .B(n7798), .ZN(P1_U3234) );
  INV_X1 U9565 ( .A(n7800), .ZN(n7827) );
  OAI222_X1 U9566 ( .A1(n9769), .A2(n7827), .B1(P1_U3086), .B2(n7802), .C1(
        n7801), .C2(n9771), .ZN(P1_U3329) );
  XNOR2_X1 U9567 ( .A(n7803), .B(n9094), .ZN(n9789) );
  INV_X1 U9568 ( .A(n9789), .ZN(n7816) );
  NAND2_X1 U9569 ( .A1(n7804), .A2(n9094), .ZN(n9785) );
  NAND3_X1 U9570 ( .A1(n9786), .A2(n9785), .A3(n9841), .ZN(n7815) );
  OAI22_X1 U9571 ( .A1(n9598), .A2(n7805), .B1(n8974), .B2(n9846), .ZN(n7806)
         );
  AOI21_X1 U9572 ( .B1(n7807), .B2(n9780), .A(n7806), .ZN(n7808) );
  OAI21_X1 U9573 ( .B1(n9603), .B2(n7809), .A(n7808), .ZN(n7812) );
  OAI211_X1 U9574 ( .C1(n7810), .C2(n9784), .A(n9837), .B(n4530), .ZN(n9783)
         );
  NOR2_X1 U9575 ( .A1(n9783), .A2(n9606), .ZN(n7811) );
  AOI211_X1 U9576 ( .C1(n7133), .C2(n7813), .A(n7812), .B(n7811), .ZN(n7814)
         );
  OAI211_X1 U9577 ( .C1(n7816), .C2(n9612), .A(n7815), .B(n7814), .ZN(P1_U3277) );
  NAND2_X1 U9578 ( .A1(n7817), .A2(n8741), .ZN(n7818) );
  XOR2_X1 U9579 ( .A(n7943), .B(n8317), .Z(n7905) );
  XNOR2_X1 U9580 ( .A(n7905), .B(n8727), .ZN(n7820) );
  XNOR2_X1 U9581 ( .A(n7908), .B(n7820), .ZN(n7825) );
  AND2_X1 U9582 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8359) );
  NOR2_X1 U9583 ( .A1(n8110), .A2(n8743), .ZN(n7821) );
  AOI211_X1 U9584 ( .C1(n4427), .C2(n8343), .A(n8359), .B(n7821), .ZN(n7822)
         );
  OAI21_X1 U9585 ( .B1(n8746), .B2(n8044), .A(n7822), .ZN(n7823) );
  AOI21_X1 U9586 ( .B1(n8037), .B2(n8317), .A(n7823), .ZN(n7824) );
  OAI21_X1 U9587 ( .B1(n7825), .B2(n8039), .A(n7824), .ZN(P2_U3174) );
  OAI222_X1 U9588 ( .A1(P2_U3151), .A2(n7828), .B1(n8900), .B2(n7827), .C1(
        n7826), .C2(n8899), .ZN(P2_U3269) );
  INV_X1 U9589 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7836) );
  OAI22_X1 U9590 ( .A1(n7829), .A2(n9952), .B1(n9622), .B2(n9950), .ZN(n7830)
         );
  AOI211_X1 U9591 ( .C1(n7832), .C2(n9887), .A(n7831), .B(n7830), .ZN(n7833)
         );
  OAI21_X1 U9592 ( .B1(n7834), .B2(n9894), .A(n7833), .ZN(n7835) );
  INV_X1 U9593 ( .A(n7835), .ZN(n7838) );
  MUX2_X1 U9594 ( .A(n7836), .B(n7838), .S(n9967), .Z(n7837) );
  OAI21_X1 U9595 ( .B1(n7840), .B2(n9754), .A(n7837), .ZN(P1_U3498) );
  MUX2_X1 U9596 ( .A(n5409), .B(n7838), .S(n9983), .Z(n7839) );
  OAI21_X1 U9597 ( .B1(n7840), .B2(n9707), .A(n7839), .ZN(P1_U3537) );
  INV_X1 U9598 ( .A(n7841), .ZN(n7847) );
  OAI222_X1 U9599 ( .A1(n9769), .A2(n7847), .B1(n7843), .B2(P1_U3086), .C1(
        n7842), .C2(n9771), .ZN(P1_U3328) );
  NAND2_X1 U9600 ( .A1(n7849), .A2(n8897), .ZN(n7845) );
  OAI211_X1 U9601 ( .C1(n8899), .C2(n7846), .A(n7845), .B(n7844), .ZN(P2_U3267) );
  OAI222_X1 U9602 ( .A1(n8899), .A2(n7848), .B1(n8900), .B2(n7847), .C1(n4446), 
        .C2(P2_U3151), .ZN(P2_U3268) );
  INV_X1 U9603 ( .A(n7849), .ZN(n7851) );
  OAI222_X1 U9604 ( .A1(n9769), .A2(n7851), .B1(n4443), .B2(P1_U3086), .C1(
        n7850), .C2(n9771), .ZN(P1_U3327) );
  INV_X1 U9605 ( .A(n7852), .ZN(n7854) );
  OAI22_X1 U9606 ( .A1(n7856), .A2(n7855), .B1(n7854), .B2(n7853), .ZN(n7859)
         );
  NAND2_X1 U9607 ( .A1(n7857), .A2(n8947), .ZN(n7858) );
  NOR2_X1 U9608 ( .A1(n7859), .A2(n7858), .ZN(n8950) );
  AOI21_X1 U9609 ( .B1(n7859), .B2(n7858), .A(n8950), .ZN(n7865) );
  NOR2_X1 U9610 ( .A1(n9043), .A2(n9793), .ZN(n7860) );
  AOI211_X1 U9611 ( .C1(n9045), .C2(n9318), .A(n7861), .B(n7860), .ZN(n7862)
         );
  OAI21_X1 U9612 ( .B1(n9048), .B2(n9800), .A(n7862), .ZN(n7863) );
  AOI21_X1 U9613 ( .B1(n9802), .B2(n9050), .A(n7863), .ZN(n7864) );
  OAI21_X1 U9614 ( .B1(n7865), .B2(n9052), .A(n7864), .ZN(P1_U3236) );
  INV_X1 U9615 ( .A(n7866), .ZN(n7966) );
  OAI222_X1 U9616 ( .A1(n9769), .A2(n7966), .B1(n7868), .B2(P1_U3086), .C1(
        n7867), .C2(n9771), .ZN(P1_U3326) );
  OAI222_X1 U9617 ( .A1(n8899), .A2(n10301), .B1(n8900), .B2(n7869), .C1(n6490), .C2(P2_U3151), .ZN(P2_U3271) );
  INV_X1 U9618 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10189) );
  OAI222_X1 U9619 ( .A1(n9771), .A2(n10189), .B1(n9769), .B2(n7870), .C1(n5713), .C2(P1_U3086), .ZN(P1_U3336) );
  NAND2_X1 U9620 ( .A1(n9115), .A2(n9113), .ZN(n9102) );
  XOR2_X1 U9621 ( .A(n9102), .B(n7871), .Z(n9654) );
  XNOR2_X1 U9622 ( .A(n7872), .B(n9102), .ZN(n9652) );
  INV_X1 U9623 ( .A(n9521), .ZN(n7873) );
  AOI211_X1 U9624 ( .C1(n9731), .C2(n9537), .A(n9822), .B(n7873), .ZN(n9650)
         );
  NAND2_X1 U9625 ( .A1(n9650), .A2(n9851), .ZN(n7878) );
  INV_X1 U9626 ( .A(n8963), .ZN(n7874) );
  AOI22_X1 U9627 ( .A1(n7874), .A2(n9820), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9857), .ZN(n7875) );
  OAI21_X1 U9628 ( .B1(n9648), .B2(n9602), .A(n7875), .ZN(n7876) );
  AOI21_X1 U9629 ( .B1(n9498), .B2(n9600), .A(n7876), .ZN(n7877) );
  OAI211_X1 U9630 ( .C1(n7879), .C2(n9618), .A(n7878), .B(n7877), .ZN(n7880)
         );
  AOI21_X1 U9631 ( .B1(n7902), .B2(n9652), .A(n7880), .ZN(n7881) );
  OAI21_X1 U9632 ( .B1(n9654), .B2(n9629), .A(n7881), .ZN(P1_U3268) );
  XNOR2_X1 U9633 ( .A(n7882), .B(n9099), .ZN(n9679) );
  AOI211_X1 U9634 ( .C1(n9676), .C2(n7893), .A(n9822), .B(n9566), .ZN(n9675)
         );
  INV_X1 U9635 ( .A(n9676), .ZN(n7884) );
  AOI22_X1 U9636 ( .A1(n8941), .A2(n9820), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9857), .ZN(n7883) );
  OAI21_X1 U9637 ( .B1(n7884), .B2(n9618), .A(n7883), .ZN(n7890) );
  AND2_X1 U9638 ( .A1(n7885), .A2(n9121), .ZN(n7887) );
  OAI21_X1 U9639 ( .B1(n7887), .B2(n9099), .A(n7886), .ZN(n7888) );
  AOI222_X1 U9640 ( .A1(n9887), .A2(n7888), .B1(n9583), .B2(n9918), .C1(n9555), 
        .C2(n9891), .ZN(n9678) );
  NOR2_X1 U9641 ( .A1(n9678), .A2(n9857), .ZN(n7889) );
  AOI211_X1 U9642 ( .C1(n9675), .C2(n9851), .A(n7890), .B(n7889), .ZN(n7891)
         );
  OAI21_X1 U9643 ( .B1(n9629), .B2(n9679), .A(n7891), .ZN(P1_U3272) );
  XNOR2_X1 U9644 ( .A(n7895), .B(n9583), .ZN(n9097) );
  XOR2_X1 U9645 ( .A(n9097), .B(n7892), .Z(n9686) );
  INV_X1 U9646 ( .A(n7893), .ZN(n7894) );
  AOI211_X1 U9647 ( .C1(n7895), .C2(n9585), .A(n9822), .B(n7894), .ZN(n9683)
         );
  INV_X1 U9648 ( .A(n7895), .ZN(n9747) );
  NOR2_X1 U9649 ( .A1(n9747), .A2(n9618), .ZN(n7900) );
  NAND2_X1 U9650 ( .A1(n9312), .A2(n9600), .ZN(n7898) );
  INV_X1 U9651 ( .A(n9002), .ZN(n7896) );
  AOI22_X1 U9652 ( .A1(n7896), .A2(n9820), .B1(P1_REG2_REG_20__SCAN_IN), .B2(
        n9857), .ZN(n7897) );
  OAI211_X1 U9653 ( .C1(n9680), .C2(n9602), .A(n7898), .B(n7897), .ZN(n7899)
         );
  AOI211_X1 U9654 ( .C1(n9683), .C2(n9851), .A(n7900), .B(n7899), .ZN(n7904)
         );
  XNOR2_X1 U9655 ( .A(n7901), .B(n9097), .ZN(n9684) );
  NAND2_X1 U9656 ( .A1(n9684), .A2(n7902), .ZN(n7903) );
  OAI211_X1 U9657 ( .C1(n9686), .C2(n9629), .A(n7904), .B(n7903), .ZN(P1_U3273) );
  XNOR2_X1 U9658 ( .A(n8887), .B(n7943), .ZN(n7909) );
  NOR2_X1 U9659 ( .A1(n7905), .A2(n8727), .ZN(n7907) );
  INV_X1 U9660 ( .A(n7905), .ZN(n7906) );
  XOR2_X1 U9661 ( .A(n8714), .B(n7909), .Z(n7977) );
  XNOR2_X1 U9662 ( .A(n8803), .B(n7943), .ZN(n7910) );
  XNOR2_X1 U9663 ( .A(n7910), .B(n8729), .ZN(n8106) );
  XNOR2_X1 U9664 ( .A(n8879), .B(n7943), .ZN(n7911) );
  XNOR2_X1 U9665 ( .A(n7911), .B(n8713), .ZN(n8031) );
  INV_X1 U9666 ( .A(n7911), .ZN(n7912) );
  AOI22_X2 U9667 ( .A1(n8032), .A2(n8031), .B1(n7912), .B2(n8713), .ZN(n8041)
         );
  XNOR2_X1 U9668 ( .A(n8795), .B(n7938), .ZN(n7913) );
  NOR2_X1 U9669 ( .A1(n7913), .A2(n8704), .ZN(n7914) );
  AOI21_X1 U9670 ( .B1(n7913), .B2(n8704), .A(n7914), .ZN(n8042) );
  INV_X1 U9671 ( .A(n7914), .ZN(n8082) );
  XNOR2_X1 U9672 ( .A(n8872), .B(n7943), .ZN(n7915) );
  NAND2_X1 U9673 ( .A1(n7915), .A2(n8659), .ZN(n7918) );
  INV_X1 U9674 ( .A(n7915), .ZN(n7916) );
  NAND2_X1 U9675 ( .A1(n7916), .A2(n8687), .ZN(n7917) );
  NAND2_X1 U9676 ( .A1(n7918), .A2(n7917), .ZN(n8081) );
  INV_X1 U9677 ( .A(n7918), .ZN(n8006) );
  XNOR2_X1 U9678 ( .A(n8788), .B(n7943), .ZN(n7919) );
  NAND2_X1 U9679 ( .A1(n7919), .A2(n8648), .ZN(n8062) );
  INV_X1 U9680 ( .A(n7919), .ZN(n7920) );
  NAND2_X1 U9681 ( .A1(n7920), .A2(n8678), .ZN(n7921) );
  AND2_X1 U9682 ( .A1(n8062), .A2(n7921), .ZN(n8005) );
  XNOR2_X1 U9683 ( .A(n8653), .B(n7943), .ZN(n7922) );
  NAND2_X1 U9684 ( .A1(n7922), .A2(n8660), .ZN(n7925) );
  INV_X1 U9685 ( .A(n7922), .ZN(n7923) );
  INV_X1 U9686 ( .A(n8660), .ZN(n8634) );
  NAND2_X1 U9687 ( .A1(n7923), .A2(n8634), .ZN(n7924) );
  NAND2_X1 U9688 ( .A1(n7925), .A2(n7924), .ZN(n8061) );
  INV_X1 U9689 ( .A(n7925), .ZN(n8014) );
  XNOR2_X1 U9690 ( .A(n8859), .B(n7943), .ZN(n7926) );
  NAND2_X1 U9691 ( .A1(n7926), .A2(n8649), .ZN(n8072) );
  INV_X1 U9692 ( .A(n7926), .ZN(n7927) );
  INV_X1 U9693 ( .A(n8649), .ZN(n8619) );
  NAND2_X1 U9694 ( .A1(n7927), .A2(n8619), .ZN(n7928) );
  XNOR2_X1 U9695 ( .A(n6458), .B(n7943), .ZN(n7929) );
  XNOR2_X1 U9696 ( .A(n7929), .B(n8633), .ZN(n8073) );
  NAND2_X1 U9697 ( .A1(n8074), .A2(n7930), .ZN(n7932) );
  XNOR2_X1 U9698 ( .A(n6462), .B(n7943), .ZN(n7931) );
  NAND2_X1 U9699 ( .A1(n7984), .A2(n8050), .ZN(n7936) );
  XNOR2_X1 U9700 ( .A(n8843), .B(n7943), .ZN(n7933) );
  NAND2_X1 U9701 ( .A1(n7933), .A2(n8583), .ZN(n8022) );
  INV_X1 U9702 ( .A(n7933), .ZN(n7934) );
  NAND2_X1 U9703 ( .A1(n7934), .A2(n8605), .ZN(n7935) );
  NAND2_X1 U9704 ( .A1(n7936), .A2(n8051), .ZN(n8021) );
  NAND2_X1 U9705 ( .A1(n8021), .A2(n8022), .ZN(n7937) );
  XNOR2_X1 U9706 ( .A(n8585), .B(n7943), .ZN(n7939) );
  XNOR2_X1 U9707 ( .A(n7939), .B(n8342), .ZN(n8023) );
  NAND2_X1 U9708 ( .A1(n7937), .A2(n8023), .ZN(n8025) );
  XNOR2_X1 U9709 ( .A(n8832), .B(n7938), .ZN(n8093) );
  OR2_X1 U9710 ( .A1(n8093), .A2(n8565), .ZN(n7940) );
  NAND2_X1 U9711 ( .A1(n7939), .A2(n8594), .ZN(n8092) );
  NAND2_X1 U9712 ( .A1(n8093), .A2(n8565), .ZN(n8091) );
  XNOR2_X1 U9713 ( .A(n8826), .B(n7943), .ZN(n7941) );
  XNOR2_X1 U9714 ( .A(n7941), .B(n8341), .ZN(n7967) );
  INV_X1 U9715 ( .A(n7941), .ZN(n7942) );
  XOR2_X1 U9716 ( .A(n7943), .B(n8552), .Z(n7944) );
  AOI22_X1 U9717 ( .A1(n8341), .A2(n4427), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7946) );
  NAND2_X1 U9718 ( .A1(n8557), .A2(n8113), .ZN(n7945) );
  OAI211_X1 U9719 ( .C1(n8553), .C2(n8110), .A(n7946), .B(n7945), .ZN(n7947)
         );
  AOI21_X1 U9720 ( .B1(n8558), .B2(n8037), .A(n7947), .ZN(n7948) );
  OAI22_X1 U9721 ( .A1(n9649), .A2(n8983), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7952), .ZN(n7955) );
  NOR2_X1 U9722 ( .A1(n7953), .A2(n9043), .ZN(n7954) );
  AOI211_X1 U9723 ( .C1(n9503), .C2(n8991), .A(n7955), .B(n7954), .ZN(n7956)
         );
  NAND2_X1 U9724 ( .A1(n7957), .A2(n8748), .ZN(n7962) );
  NOR2_X1 U9725 ( .A1(n7958), .A2(n8745), .ZN(n8544) );
  NOR2_X1 U9726 ( .A1(n7959), .A2(n8720), .ZN(n7960) );
  AOI211_X1 U9727 ( .C1(n8752), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8544), .B(
        n7960), .ZN(n7961) );
  OAI211_X1 U9728 ( .C1(n7964), .C2(n7963), .A(n7962), .B(n7961), .ZN(P2_U3204) );
  OAI222_X1 U9729 ( .A1(n6050), .A2(P2_U3151), .B1(n8900), .B2(n7966), .C1(
        n7965), .C2(n8899), .ZN(P2_U3266) );
  XNOR2_X1 U9730 ( .A(n7968), .B(n7967), .ZN(n7974) );
  AOI22_X1 U9731 ( .A1(n8565), .A2(n4427), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7970) );
  NAND2_X1 U9732 ( .A1(n8568), .A2(n8113), .ZN(n7969) );
  OAI211_X1 U9733 ( .C1(n7971), .C2(n8110), .A(n7970), .B(n7969), .ZN(n7972)
         );
  AOI21_X1 U9734 ( .B1(n8826), .B2(n8037), .A(n7972), .ZN(n7973) );
  OAI21_X1 U9735 ( .B1(n7974), .B2(n8039), .A(n7973), .ZN(P2_U3154) );
  AOI21_X1 U9736 ( .B1(n7977), .B2(n7975), .A(n7976), .ZN(n7983) );
  INV_X1 U9737 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7978) );
  NOR2_X1 U9738 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7978), .ZN(n8392) );
  NOR2_X1 U9739 ( .A1(n8110), .A2(n8302), .ZN(n7979) );
  AOI211_X1 U9740 ( .C1(n4427), .C2(n8727), .A(n8392), .B(n7979), .ZN(n7980)
         );
  OAI21_X1 U9741 ( .B1(n8724), .B2(n8044), .A(n7980), .ZN(n7981) );
  AOI21_X1 U9742 ( .B1(n8887), .B2(n8037), .A(n7981), .ZN(n7982) );
  OAI21_X1 U9743 ( .B1(n7983), .B2(n8039), .A(n7982), .ZN(P2_U3155) );
  INV_X1 U9744 ( .A(n7984), .ZN(n8053) );
  AOI21_X1 U9745 ( .B1(n8618), .B2(n7985), .A(n8053), .ZN(n7990) );
  AOI22_X1 U9746 ( .A1(n8633), .A2(n4427), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n7987) );
  NAND2_X1 U9747 ( .A1(n8113), .A2(n8608), .ZN(n7986) );
  OAI211_X1 U9748 ( .C1(n8583), .C2(n8110), .A(n7987), .B(n7986), .ZN(n7988)
         );
  AOI21_X1 U9749 ( .B1(n6462), .B2(n8037), .A(n7988), .ZN(n7989) );
  OAI21_X1 U9750 ( .B1(n7990), .B2(n8039), .A(n7989), .ZN(P2_U3156) );
  NAND2_X1 U9751 ( .A1(n7992), .A2(n7991), .ZN(n7994) );
  AOI21_X1 U9752 ( .B1(n7994), .B2(n7993), .A(n8039), .ZN(n7996) );
  NAND2_X1 U9753 ( .A1(n7996), .A2(n7995), .ZN(n8003) );
  AOI21_X1 U9754 ( .B1(n4427), .B2(n4442), .A(n7997), .ZN(n8002) );
  AOI22_X1 U9755 ( .A1(n8066), .A2(n7998), .B1(n8037), .B2(n10011), .ZN(n8001)
         );
  NAND2_X1 U9756 ( .A1(n8113), .A2(n7999), .ZN(n8000) );
  NAND4_X1 U9757 ( .A1(n8003), .A2(n8002), .A3(n8001), .A4(n8000), .ZN(
        P2_U3158) );
  INV_X1 U9758 ( .A(n8788), .ZN(n8668) );
  INV_X1 U9759 ( .A(n8063), .ZN(n8008) );
  NOR3_X1 U9760 ( .A1(n8004), .A2(n8006), .A3(n8005), .ZN(n8007) );
  OAI21_X1 U9761 ( .B1(n8008), .B2(n8007), .A(n8104), .ZN(n8012) );
  NAND2_X1 U9762 ( .A1(n8687), .A2(n4427), .ZN(n8009) );
  NAND2_X1 U9763 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8530) );
  OAI211_X1 U9764 ( .C1(n8660), .C2(n8110), .A(n8009), .B(n8530), .ZN(n8010)
         );
  AOI21_X1 U9765 ( .B1(n8666), .B2(n8113), .A(n8010), .ZN(n8011) );
  OAI211_X1 U9766 ( .C1(n8668), .C2(n8116), .A(n8012), .B(n8011), .ZN(P2_U3159) );
  NOR3_X1 U9767 ( .A1(n8065), .A2(n8014), .A3(n8013), .ZN(n8015) );
  OAI21_X1 U9768 ( .B1(n4470), .B2(n8015), .A(n8104), .ZN(n8019) );
  AOI22_X1 U9769 ( .A1(n8633), .A2(n8066), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8016) );
  OAI21_X1 U9770 ( .B1(n8660), .B2(n8068), .A(n8016), .ZN(n8017) );
  AOI21_X1 U9771 ( .B1(n8637), .B2(n8113), .A(n8017), .ZN(n8018) );
  OAI211_X1 U9772 ( .C1(n8020), .C2(n8116), .A(n8019), .B(n8018), .ZN(P2_U3163) );
  INV_X1 U9773 ( .A(n8021), .ZN(n8054) );
  INV_X1 U9774 ( .A(n8022), .ZN(n8024) );
  NOR3_X1 U9775 ( .A1(n8054), .A2(n8024), .A3(n8023), .ZN(n8026) );
  INV_X1 U9776 ( .A(n8025), .ZN(n8096) );
  OAI21_X1 U9777 ( .B1(n8026), .B2(n8096), .A(n8104), .ZN(n8030) );
  AOI22_X1 U9778 ( .A1(n8565), .A2(n8066), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8027) );
  OAI21_X1 U9779 ( .B1(n8583), .B2(n8068), .A(n8027), .ZN(n8028) );
  AOI21_X1 U9780 ( .B1(n8586), .B2(n8113), .A(n8028), .ZN(n8029) );
  OAI211_X1 U9781 ( .C1(n8837), .C2(n8116), .A(n8030), .B(n8029), .ZN(P2_U3165) );
  XNOR2_X1 U9782 ( .A(n8032), .B(n8031), .ZN(n8040) );
  INV_X1 U9783 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10288) );
  OR2_X1 U9784 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10288), .ZN(n8449) );
  OAI21_X1 U9785 ( .B1(n8110), .B2(n8033), .A(n8449), .ZN(n8034) );
  AOI21_X1 U9786 ( .B1(n4427), .B2(n8729), .A(n8034), .ZN(n8035) );
  OAI21_X1 U9787 ( .B1(n8044), .B2(n8706), .A(n8035), .ZN(n8036) );
  AOI21_X1 U9788 ( .B1(n8879), .B2(n8037), .A(n8036), .ZN(n8038) );
  OAI21_X1 U9789 ( .B1(n8040), .B2(n8039), .A(n8038), .ZN(P2_U3166) );
  OAI21_X1 U9790 ( .B1(n8042), .B2(n8041), .A(n8083), .ZN(n8043) );
  NAND2_X1 U9791 ( .A1(n8043), .A2(n8104), .ZN(n8049) );
  NAND2_X1 U9792 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8477) );
  OAI21_X1 U9793 ( .B1(n8110), .B2(n8659), .A(n8477), .ZN(n8046) );
  NOR2_X1 U9794 ( .A1(n8044), .A2(n8692), .ZN(n8045) );
  AOI211_X1 U9795 ( .C1(n4427), .C2(n8713), .A(n8046), .B(n8045), .ZN(n8048)
         );
  OAI211_X1 U9796 ( .C1(n8691), .C2(n8116), .A(n8049), .B(n8048), .ZN(P2_U3168) );
  INV_X1 U9797 ( .A(n8050), .ZN(n8052) );
  NOR3_X1 U9798 ( .A1(n8053), .A2(n8052), .A3(n8051), .ZN(n8055) );
  OAI21_X1 U9799 ( .B1(n8055), .B2(n8054), .A(n8104), .ZN(n8059) );
  AOI22_X1 U9800 ( .A1(n8342), .A2(n8066), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8056) );
  OAI21_X1 U9801 ( .B1(n8595), .B2(n8068), .A(n8056), .ZN(n8057) );
  AOI21_X1 U9802 ( .B1(n8596), .B2(n8113), .A(n8057), .ZN(n8058) );
  OAI211_X1 U9803 ( .C1(n8060), .C2(n8116), .A(n8059), .B(n8058), .ZN(P2_U3169) );
  AND3_X1 U9804 ( .A1(n8063), .A2(n8062), .A3(n8061), .ZN(n8064) );
  OAI21_X1 U9805 ( .B1(n8065), .B2(n8064), .A(n8104), .ZN(n8071) );
  AOI22_X1 U9806 ( .A1(n8619), .A2(n8066), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8067) );
  OAI21_X1 U9807 ( .B1(n8648), .B2(n8068), .A(n8067), .ZN(n8069) );
  AOI21_X1 U9808 ( .B1(n8652), .B2(n8113), .A(n8069), .ZN(n8070) );
  OAI211_X1 U9809 ( .C1(n8865), .C2(n8116), .A(n8071), .B(n8070), .ZN(P2_U3173) );
  NOR3_X1 U9810 ( .A1(n4470), .A2(n4802), .A3(n8073), .ZN(n8076) );
  INV_X1 U9811 ( .A(n8074), .ZN(n8075) );
  OAI21_X1 U9812 ( .B1(n8076), .B2(n8075), .A(n8104), .ZN(n8080) );
  AOI22_X1 U9813 ( .A1(n8619), .A2(n4427), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8077) );
  OAI21_X1 U9814 ( .B1(n8595), .B2(n8110), .A(n8077), .ZN(n8078) );
  AOI21_X1 U9815 ( .B1(n8621), .B2(n8113), .A(n8078), .ZN(n8079) );
  OAI211_X1 U9816 ( .C1(n6460), .C2(n8116), .A(n8080), .B(n8079), .ZN(P2_U3175) );
  INV_X1 U9817 ( .A(n8872), .ZN(n8090) );
  AND3_X1 U9818 ( .A1(n8083), .A2(n8082), .A3(n8081), .ZN(n8084) );
  OAI21_X1 U9819 ( .B1(n8004), .B2(n8084), .A(n8104), .ZN(n8089) );
  INV_X1 U9820 ( .A(n8085), .ZN(n8681) );
  NAND2_X1 U9821 ( .A1(n4427), .A2(n8704), .ZN(n8086) );
  NAND2_X1 U9822 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8499) );
  OAI211_X1 U9823 ( .C1(n8110), .C2(n8648), .A(n8086), .B(n8499), .ZN(n8087)
         );
  AOI21_X1 U9824 ( .B1(n8113), .B2(n8681), .A(n8087), .ZN(n8088) );
  OAI211_X1 U9825 ( .C1(n8090), .C2(n8116), .A(n8089), .B(n8088), .ZN(P2_U3178) );
  INV_X1 U9826 ( .A(n8832), .ZN(n8103) );
  INV_X1 U9827 ( .A(n8092), .ZN(n8095) );
  XNOR2_X1 U9828 ( .A(n8093), .B(n8565), .ZN(n8094) );
  OAI211_X1 U9829 ( .C1(n4820), .C2(n8098), .A(n8097), .B(n8104), .ZN(n8102)
         );
  AOI22_X1 U9830 ( .A1(n8342), .A2(n4427), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8099) );
  OAI21_X1 U9831 ( .B1(n8574), .B2(n8110), .A(n8099), .ZN(n8100) );
  AOI21_X1 U9832 ( .B1(n8575), .B2(n8113), .A(n8100), .ZN(n8101) );
  OAI211_X1 U9833 ( .C1(n8103), .C2(n8116), .A(n8102), .B(n8101), .ZN(P2_U3180) );
  OAI211_X1 U9834 ( .C1(n8107), .C2(n8106), .A(n8105), .B(n8104), .ZN(n8115)
         );
  INV_X1 U9835 ( .A(n8108), .ZN(n8717) );
  NOR2_X1 U9836 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6254), .ZN(n8423) );
  AOI21_X1 U9837 ( .B1(n4427), .B2(n8714), .A(n8423), .ZN(n8109) );
  OAI21_X1 U9838 ( .B1(n8111), .B2(n8110), .A(n8109), .ZN(n8112) );
  AOI21_X1 U9839 ( .B1(n8717), .B2(n8113), .A(n8112), .ZN(n8114) );
  OAI211_X1 U9840 ( .C1(n8721), .C2(n8116), .A(n8115), .B(n8114), .ZN(P2_U3181) );
  INV_X1 U9841 ( .A(SI_29_), .ZN(n8120) );
  INV_X1 U9842 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n10317) );
  INV_X1 U9843 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9770) );
  MUX2_X1 U9844 ( .A(n10317), .B(n9770), .S(n4436), .Z(n8122) );
  NAND2_X1 U9845 ( .A1(n8122), .A2(n10126), .ZN(n8127) );
  INV_X1 U9846 ( .A(n8122), .ZN(n8123) );
  NAND2_X1 U9847 ( .A1(n8123), .A2(SI_30_), .ZN(n8124) );
  NAND2_X1 U9848 ( .A1(n8127), .A2(n8124), .ZN(n8128) );
  NAND2_X1 U9849 ( .A1(n9054), .A2(n6183), .ZN(n8126) );
  OR2_X1 U9850 ( .A1(n8133), .A2(n10317), .ZN(n8125) );
  INV_X1 U9851 ( .A(n8758), .ZN(n8817) );
  INV_X1 U9852 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9760) );
  MUX2_X1 U9853 ( .A(n6672), .B(n9760), .S(n4436), .Z(n8130) );
  XNOR2_X1 U9854 ( .A(n8130), .B(SI_31_), .ZN(n8131) );
  NAND2_X1 U9855 ( .A1(n9765), .A2(n6183), .ZN(n8135) );
  OR2_X1 U9856 ( .A1(n8133), .A2(n6672), .ZN(n8134) );
  INV_X1 U9857 ( .A(n8136), .ZN(n8138) );
  AOI21_X1 U9858 ( .B1(n8138), .B2(n8291), .A(n8137), .ZN(n8139) );
  OR2_X1 U9859 ( .A1(n8756), .A2(n8543), .ZN(n8143) );
  INV_X1 U9860 ( .A(n8340), .ZN(n8290) );
  NAND2_X1 U9861 ( .A1(n8758), .A2(n8290), .ZN(n8141) );
  NAND2_X1 U9862 ( .A1(n8141), .A2(n8140), .ZN(n8281) );
  INV_X1 U9863 ( .A(n8281), .ZN(n8142) );
  NAND2_X1 U9864 ( .A1(n8143), .A2(n8142), .ZN(n8333) );
  OAI21_X1 U9865 ( .B1(n8290), .B2(n8292), .A(n8758), .ZN(n8145) );
  OAI211_X1 U9866 ( .C1(n8274), .C2(n8340), .A(n8145), .B(n8144), .ZN(n8297)
         );
  INV_X1 U9867 ( .A(n8611), .ZN(n8615) );
  NAND2_X1 U9868 ( .A1(n8254), .A2(n8246), .ZN(n8301) );
  AND2_X1 U9869 ( .A1(n8301), .A2(n8146), .ZN(n8257) );
  INV_X1 U9870 ( .A(n8154), .ZN(n8148) );
  NAND2_X1 U9871 ( .A1(n8148), .A2(n8147), .ZN(n8150) );
  NAND2_X1 U9872 ( .A1(n8162), .A2(n8161), .ZN(n8149) );
  MUX2_X1 U9873 ( .A(n8150), .B(n8149), .S(n8292), .Z(n8158) );
  INV_X1 U9874 ( .A(n8158), .ZN(n8166) );
  NAND2_X1 U9875 ( .A1(n8166), .A2(n8311), .ZN(n8168) );
  INV_X1 U9876 ( .A(n8153), .ZN(n8155) );
  NOR2_X1 U9877 ( .A1(n8155), .A2(n8154), .ZN(n8157) );
  OAI211_X1 U9878 ( .C1(n8158), .C2(n8157), .A(n8156), .B(n8292), .ZN(n8159)
         );
  NOR2_X1 U9879 ( .A1(n8316), .A2(n8159), .ZN(n8210) );
  OAI21_X1 U9880 ( .B1(n6141), .B2(n8168), .A(n8210), .ZN(n8172) );
  NAND2_X1 U9881 ( .A1(n8161), .A2(n8160), .ZN(n8165) );
  NAND3_X1 U9882 ( .A1(n8163), .A2(n8274), .A3(n8162), .ZN(n8164) );
  AOI21_X1 U9883 ( .B1(n8166), .B2(n8165), .A(n8164), .ZN(n8167) );
  INV_X1 U9884 ( .A(n8168), .ZN(n8169) );
  NAND2_X1 U9885 ( .A1(n8169), .A2(n8209), .ZN(n8170) );
  NAND2_X1 U9886 ( .A1(n8218), .A2(n8170), .ZN(n8171) );
  AND2_X1 U9887 ( .A1(n8172), .A2(n8171), .ZN(n8222) );
  AND2_X1 U9888 ( .A1(n8345), .A2(n8274), .ZN(n8174) );
  OAI21_X1 U9889 ( .B1(n8274), .B2(n8345), .A(n10049), .ZN(n8173) );
  OAI21_X1 U9890 ( .B1(n8174), .B2(n10049), .A(n8173), .ZN(n8175) );
  NAND2_X1 U9891 ( .A1(n8176), .A2(n8175), .ZN(n8185) );
  NAND2_X1 U9892 ( .A1(n8178), .A2(n8177), .ZN(n8180) );
  NAND2_X1 U9893 ( .A1(n8180), .A2(n8179), .ZN(n8182) );
  NAND2_X1 U9894 ( .A1(n8182), .A2(n8274), .ZN(n8181) );
  NAND2_X1 U9895 ( .A1(n8316), .A2(n8181), .ZN(n8184) );
  NOR2_X1 U9896 ( .A1(n8182), .A2(n8274), .ZN(n8183) );
  AOI21_X1 U9897 ( .B1(n8185), .B2(n8184), .A(n8183), .ZN(n8221) );
  MUX2_X1 U9898 ( .A(n8188), .B(n8186), .S(n8292), .Z(n8196) );
  NAND2_X1 U9899 ( .A1(n8187), .A2(n8337), .ZN(n8191) );
  NAND2_X1 U9900 ( .A1(n8187), .A2(n8194), .ZN(n8189) );
  NAND3_X1 U9901 ( .A1(n8189), .A2(n8292), .A3(n8188), .ZN(n8190) );
  OAI21_X1 U9902 ( .B1(n8192), .B2(n8191), .A(n8190), .ZN(n8193) );
  OAI21_X1 U9903 ( .B1(n8194), .B2(n6881), .A(n8193), .ZN(n8195) );
  NAND3_X1 U9904 ( .A1(n8196), .A2(n8195), .A3(n7103), .ZN(n8203) );
  NAND2_X1 U9905 ( .A1(n8211), .A2(n8197), .ZN(n8200) );
  NAND2_X1 U9906 ( .A1(n8205), .A2(n8198), .ZN(n8199) );
  MUX2_X1 U9907 ( .A(n8200), .B(n8199), .S(n8274), .Z(n8201) );
  INV_X1 U9908 ( .A(n8201), .ZN(n8202) );
  NAND2_X1 U9909 ( .A1(n8203), .A2(n8202), .ZN(n8204) );
  NAND2_X1 U9910 ( .A1(n8204), .A2(n8303), .ZN(n8214) );
  INV_X1 U9911 ( .A(n8205), .ZN(n8207) );
  OAI211_X1 U9912 ( .C1(n8214), .C2(n8207), .A(n8217), .B(n8206), .ZN(n8208)
         );
  NAND4_X1 U9913 ( .A1(n8210), .A2(n8209), .A3(n8208), .A4(n8212), .ZN(n8220)
         );
  OAI211_X1 U9914 ( .C1(n8214), .C2(n4746), .A(n8213), .B(n8212), .ZN(n8216)
         );
  NAND4_X1 U9915 ( .A1(n8218), .A2(n8217), .A3(n8216), .A4(n8215), .ZN(n8219)
         );
  NAND2_X1 U9916 ( .A1(n8317), .A2(n8727), .ZN(n8224) );
  MUX2_X1 U9917 ( .A(n8727), .B(n8317), .S(n8292), .Z(n8223) );
  INV_X1 U9918 ( .A(n8227), .ZN(n8234) );
  NAND3_X1 U9919 ( .A1(n8231), .A2(n8234), .A3(n8228), .ZN(n8230) );
  NAND2_X1 U9920 ( .A1(n8230), .A2(n8229), .ZN(n8237) );
  NAND2_X1 U9921 ( .A1(n8231), .A2(n8699), .ZN(n8235) );
  INV_X1 U9922 ( .A(n8232), .ZN(n8233) );
  AOI21_X1 U9923 ( .B1(n8235), .B2(n8234), .A(n8233), .ZN(n8236) );
  MUX2_X1 U9924 ( .A(n8237), .B(n8236), .S(n8274), .Z(n8241) );
  INV_X1 U9925 ( .A(n8689), .ZN(n8685) );
  AOI21_X1 U9926 ( .B1(n8239), .B2(n8238), .A(n8292), .ZN(n8240) );
  AOI21_X1 U9927 ( .B1(n8241), .B2(n8685), .A(n8240), .ZN(n8248) );
  NAND3_X1 U9928 ( .A1(n8248), .A2(n8242), .A3(n8249), .ZN(n8244) );
  NAND3_X1 U9929 ( .A1(n8872), .A2(n8659), .A3(n8292), .ZN(n8243) );
  NAND3_X1 U9930 ( .A1(n8244), .A2(n8260), .A3(n8243), .ZN(n8247) );
  NAND3_X1 U9931 ( .A1(n8247), .A2(n4736), .A3(n8246), .ZN(n8253) );
  INV_X1 U9932 ( .A(n8248), .ZN(n8250) );
  NAND3_X1 U9933 ( .A1(n8250), .A2(n8249), .A3(n4736), .ZN(n8251) );
  NAND2_X1 U9934 ( .A1(n8251), .A2(n8274), .ZN(n8252) );
  NAND2_X1 U9935 ( .A1(n8253), .A2(n8252), .ZN(n8261) );
  INV_X1 U9936 ( .A(n8261), .ZN(n8256) );
  INV_X1 U9937 ( .A(n8254), .ZN(n8255) );
  NAND2_X1 U9938 ( .A1(n8299), .A2(n8258), .ZN(n8263) );
  INV_X1 U9939 ( .A(n8266), .ZN(n8300) );
  INV_X1 U9940 ( .A(n8299), .ZN(n8264) );
  NAND2_X1 U9941 ( .A1(n8269), .A2(n8268), .ZN(n8587) );
  MUX2_X1 U9942 ( .A(n8269), .B(n8268), .S(n8292), .Z(n8270) );
  MUX2_X1 U9943 ( .A(n8271), .B(n4489), .S(n8292), .Z(n8273) );
  MUX2_X1 U9944 ( .A(n8276), .B(n8275), .S(n8274), .Z(n8277) );
  NOR2_X1 U9945 ( .A1(n8278), .A2(n8277), .ZN(n8282) );
  MUX2_X1 U9946 ( .A(n8564), .B(n8558), .S(n8292), .Z(n8283) );
  OAI21_X1 U9947 ( .B1(n8282), .B2(n8283), .A(n8279), .ZN(n8289) );
  NOR2_X1 U9948 ( .A1(n8281), .A2(n8280), .ZN(n8288) );
  INV_X1 U9949 ( .A(n8282), .ZN(n8286) );
  INV_X1 U9950 ( .A(n8283), .ZN(n8285) );
  INV_X1 U9951 ( .A(n8293), .ZN(n8287) );
  OAI211_X1 U9952 ( .C1(n8289), .C2(n8564), .A(n8288), .B(n8287), .ZN(n8296)
         );
  NOR2_X1 U9953 ( .A1(n8289), .A2(n8558), .ZN(n8294) );
  OR2_X1 U9954 ( .A1(n8758), .A2(n8290), .ZN(n8331) );
  NAND2_X1 U9955 ( .A1(n8331), .A2(n8291), .ZN(n8327) );
  NOR4_X1 U9956 ( .A1(n8294), .A2(n8293), .A3(n8292), .A4(n8327), .ZN(n8295)
         );
  AOI21_X1 U9957 ( .B1(n8297), .B2(n8296), .A(n8295), .ZN(n8332) );
  INV_X1 U9958 ( .A(n8563), .ZN(n8325) );
  NAND2_X1 U9959 ( .A1(n8300), .A2(n8299), .ZN(n8603) );
  INV_X1 U9960 ( .A(n8301), .ZN(n8321) );
  XNOR2_X1 U9961 ( .A(n8803), .B(n8302), .ZN(n8716) );
  NAND3_X1 U9962 ( .A1(n8304), .A2(n8303), .A3(n7103), .ZN(n8308) );
  NOR4_X1 U9963 ( .A1(n8308), .A2(n8307), .A3(n8306), .A4(n8305), .ZN(n8312)
         );
  NAND4_X1 U9964 ( .A1(n8312), .A2(n8311), .A3(n8310), .A4(n8309), .ZN(n8313)
         );
  NOR4_X1 U9965 ( .A1(n8316), .A2(n8315), .A3(n8314), .A4(n8313), .ZN(n8318)
         );
  XNOR2_X1 U9966 ( .A(n8317), .B(n8727), .ZN(n8751) );
  NAND4_X1 U9967 ( .A1(n8703), .A2(n8736), .A3(n8318), .A4(n8751), .ZN(n8319)
         );
  NOR4_X1 U9968 ( .A1(n8676), .A2(n8716), .A3(n8689), .A4(n8319), .ZN(n8320)
         );
  NAND4_X1 U9969 ( .A1(n8322), .A2(n8321), .A3(n8657), .A4(n8320), .ZN(n8323)
         );
  NOR4_X1 U9970 ( .A1(n8597), .A2(n8587), .A3(n8603), .A4(n8323), .ZN(n8324)
         );
  NAND4_X1 U9971 ( .A1(n8325), .A2(n8571), .A3(n8324), .A4(n8552), .ZN(n8326)
         );
  NOR3_X1 U9972 ( .A1(n8333), .A2(n8327), .A3(n8326), .ZN(n8329) );
  NAND3_X1 U9973 ( .A1(n8335), .A2(n8334), .A3(n4446), .ZN(n8336) );
  OAI211_X1 U9974 ( .C1(n8337), .C2(n8339), .A(n8336), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8338) );
  MUX2_X1 U9975 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8340), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9976 ( .A(n8564), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8497), .Z(
        P2_U3519) );
  MUX2_X1 U9977 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8341), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9978 ( .A(n8565), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8497), .Z(
        P2_U3517) );
  MUX2_X1 U9979 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8342), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9980 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8605), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9981 ( .A(n8618), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8497), .Z(
        P2_U3514) );
  MUX2_X1 U9982 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8633), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9983 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8619), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9984 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8634), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9985 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8678), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9986 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8687), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9987 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8704), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9988 ( .A(n8713), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8497), .Z(
        P2_U3507) );
  MUX2_X1 U9989 ( .A(n8729), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8497), .Z(
        P2_U3506) );
  MUX2_X1 U9990 ( .A(n8714), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8497), .Z(
        P2_U3505) );
  MUX2_X1 U9991 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8727), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9992 ( .A(n8343), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8497), .Z(
        P2_U3503) );
  MUX2_X1 U9993 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8344), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U9994 ( .A(n8345), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8497), .Z(
        P2_U3501) );
  MUX2_X1 U9995 ( .A(n8346), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8497), .Z(
        P2_U3500) );
  MUX2_X1 U9996 ( .A(n8347), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8497), .Z(
        P2_U3499) );
  MUX2_X1 U9997 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8348), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U9998 ( .A(n8349), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8497), .Z(
        P2_U3497) );
  MUX2_X1 U9999 ( .A(n8350), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8497), .Z(
        P2_U3496) );
  MUX2_X1 U10000 ( .A(n8351), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8497), .Z(
        P2_U3494) );
  MUX2_X1 U10001 ( .A(n4442), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8497), .Z(
        P2_U3493) );
  MUX2_X1 U10002 ( .A(n8353), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8497), .Z(
        P2_U3492) );
  MUX2_X1 U10003 ( .A(n8354), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8497), .Z(
        P2_U3491) );
  AOI21_X1 U10004 ( .B1(n8364), .B2(n8358), .A(n8398), .ZN(n8379) );
  INV_X1 U10005 ( .A(n8359), .ZN(n8360) );
  OAI21_X1 U10006 ( .B1(n10005), .B2(n10294), .A(n8360), .ZN(n8371) );
  MUX2_X1 U10007 ( .A(n8365), .B(n8364), .S(n4446), .Z(n8366) );
  NAND2_X1 U10008 ( .A1(n8366), .A2(n8397), .ZN(n8387) );
  OAI21_X1 U10009 ( .B1(n8366), .B2(n8397), .A(n8387), .ZN(n8367) );
  NOR2_X1 U10010 ( .A1(n8368), .A2(n8367), .ZN(n8388) );
  AOI21_X1 U10011 ( .B1(n8368), .B2(n8367), .A(n8388), .ZN(n8369) );
  NOR2_X1 U10012 ( .A1(n8369), .A2(n8535), .ZN(n8370) );
  AOI211_X1 U10013 ( .C1(n10411), .C2(n8397), .A(n8371), .B(n8370), .ZN(n8378)
         );
  AOI21_X1 U10014 ( .B1(n8365), .B2(n8375), .A(n8381), .ZN(n8376) );
  OR2_X1 U10015 ( .A1(n8376), .A2(n10002), .ZN(n8377) );
  OAI211_X1 U10016 ( .C1(n8379), .C2(n9985), .A(n8378), .B(n8377), .ZN(
        P2_U3195) );
  NOR2_X1 U10017 ( .A1(n8397), .A2(n8380), .ZN(n8382) );
  MUX2_X1 U10018 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n8408), .S(n8409), .Z(n8384) );
  INV_X1 U10019 ( .A(n8411), .ZN(n8383) );
  AOI21_X1 U10020 ( .B1(n8385), .B2(n8384), .A(n8383), .ZN(n8407) );
  INV_X1 U10021 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8807) );
  MUX2_X1 U10022 ( .A(n8408), .B(n8807), .S(n4446), .Z(n8386) );
  NAND2_X1 U10023 ( .A1(n8386), .A2(n8409), .ZN(n8418) );
  OAI21_X1 U10024 ( .B1(n8386), .B2(n8409), .A(n8418), .ZN(n8391) );
  INV_X1 U10025 ( .A(n8387), .ZN(n8389) );
  NOR2_X1 U10026 ( .A1(n8390), .A2(n8391), .ZN(n8419) );
  AOI21_X1 U10027 ( .B1(n8391), .B2(n8390), .A(n8419), .ZN(n8394) );
  AOI21_X1 U10028 ( .B1(n10405), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n8392), .ZN(
        n8393) );
  OAI21_X1 U10029 ( .B1(n8394), .B2(n8535), .A(n8393), .ZN(n8405) );
  INV_X1 U10030 ( .A(n8395), .ZN(n8396) );
  NOR2_X1 U10031 ( .A1(n8397), .A2(n8396), .ZN(n8399) );
  OR2_X1 U10032 ( .A1(n8409), .A2(n8807), .ZN(n8429) );
  NAND2_X1 U10033 ( .A1(n8409), .A2(n8807), .ZN(n8400) );
  NAND2_X1 U10034 ( .A1(n8429), .A2(n8400), .ZN(n8401) );
  NAND2_X1 U10035 ( .A1(n8402), .A2(n8401), .ZN(n8403) );
  AOI21_X1 U10036 ( .B1(n8430), .B2(n8403), .A(n9985), .ZN(n8404) );
  AOI211_X1 U10037 ( .C1(n10411), .C2(n8409), .A(n8405), .B(n8404), .ZN(n8406)
         );
  OAI21_X1 U10038 ( .B1(n8407), .B2(n10002), .A(n8406), .ZN(P2_U3196) );
  OR2_X1 U10039 ( .A1(n8409), .A2(n8408), .ZN(n8410) );
  XNOR2_X1 U10040 ( .A(n8438), .B(n8453), .ZN(n8412) );
  AOI21_X1 U10041 ( .B1(n8413), .B2(n8412), .A(n8439), .ZN(n8437) );
  MUX2_X1 U10042 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n4446), .Z(n8415) );
  INV_X1 U10043 ( .A(n8415), .ZN(n8417) );
  NOR2_X1 U10044 ( .A1(n8415), .A2(n8414), .ZN(n8444) );
  INV_X1 U10045 ( .A(n8444), .ZN(n8416) );
  OAI21_X1 U10046 ( .B1(n8453), .B2(n8417), .A(n8416), .ZN(n8422) );
  INV_X1 U10047 ( .A(n8418), .ZN(n8420) );
  NOR2_X1 U10048 ( .A1(n8420), .A2(n8419), .ZN(n8421) );
  NOR2_X1 U10049 ( .A1(n8421), .A2(n8422), .ZN(n8443) );
  AOI21_X1 U10050 ( .B1(n8422), .B2(n8421), .A(n8443), .ZN(n8428) );
  INV_X1 U10051 ( .A(n8423), .ZN(n8424) );
  OAI21_X1 U10052 ( .B1(n10005), .B2(n8425), .A(n8424), .ZN(n8426) );
  INV_X1 U10053 ( .A(n8426), .ZN(n8427) );
  OAI21_X1 U10054 ( .B1(n8428), .B2(n8535), .A(n8427), .ZN(n8435) );
  AOI21_X1 U10055 ( .B1(n8432), .B2(n8431), .A(n8454), .ZN(n8433) );
  NOR2_X1 U10056 ( .A1(n8433), .A2(n9985), .ZN(n8434) );
  AOI211_X1 U10057 ( .C1(n10411), .C2(n8453), .A(n8435), .B(n8434), .ZN(n8436)
         );
  OAI21_X1 U10058 ( .B1(n8437), .B2(n10002), .A(n8436), .ZN(P2_U3197) );
  NAND2_X1 U10059 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8475), .ZN(n8440) );
  OAI21_X1 U10060 ( .B1(n8475), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8440), .ZN(
        n8441) );
  AOI21_X1 U10061 ( .B1(n8442), .B2(n8441), .A(n8474), .ZN(n8464) );
  MUX2_X1 U10062 ( .A(n8445), .B(n8799), .S(n4446), .Z(n8446) );
  NAND2_X1 U10063 ( .A1(n8446), .A2(n8456), .ZN(n8467) );
  NOR2_X1 U10064 ( .A1(n8446), .A2(n8456), .ZN(n8469) );
  INV_X1 U10065 ( .A(n8469), .ZN(n8447) );
  NAND2_X1 U10066 ( .A1(n8467), .A2(n8447), .ZN(n8448) );
  XNOR2_X1 U10067 ( .A(n8468), .B(n8448), .ZN(n8462) );
  NAND2_X1 U10068 ( .A1(n10411), .A2(n8456), .ZN(n8450) );
  OAI211_X1 U10069 ( .C1(n8451), .C2(n10005), .A(n8450), .B(n8449), .ZN(n8461)
         );
  NOR2_X1 U10070 ( .A1(n8453), .A2(n8452), .ZN(n8455) );
  AOI22_X1 U10071 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8456), .B1(n8475), .B2(
        n8799), .ZN(n8457) );
  AOI21_X1 U10072 ( .B1(n8458), .B2(n8457), .A(n8465), .ZN(n8459) );
  NOR2_X1 U10073 ( .A1(n8459), .A2(n9985), .ZN(n8460) );
  AOI211_X1 U10074 ( .C1(n10406), .C2(n8462), .A(n8461), .B(n8460), .ZN(n8463)
         );
  OAI21_X1 U10075 ( .B1(n8464), .B2(n10002), .A(n8463), .ZN(P2_U3198) );
  NOR2_X1 U10076 ( .A1(n8470), .A2(n8466), .ZN(n8487) );
  AOI21_X1 U10077 ( .B1(n8470), .B2(n8466), .A(n8487), .ZN(n8485) );
  OAI21_X1 U10078 ( .B1(n8469), .B2(n8468), .A(n8467), .ZN(n8473) );
  MUX2_X1 U10079 ( .A(n8693), .B(n8470), .S(n4446), .Z(n8493) );
  XNOR2_X1 U10080 ( .A(n8471), .B(n8493), .ZN(n8472) );
  NAND2_X1 U10081 ( .A1(n8472), .A2(n8473), .ZN(n8491) );
  OAI21_X1 U10082 ( .B1(n8473), .B2(n8472), .A(n8491), .ZN(n8483) );
  AOI21_X1 U10083 ( .B1(n8476), .B2(n8693), .A(n8503), .ZN(n8481) );
  OAI21_X1 U10084 ( .B1(n10005), .B2(n8478), .A(n8477), .ZN(n8479) );
  AOI21_X1 U10085 ( .B1(n8502), .B2(n10411), .A(n8479), .ZN(n8480) );
  OAI21_X1 U10086 ( .B1(n8481), .B2(n10002), .A(n8480), .ZN(n8482) );
  AOI21_X1 U10087 ( .B1(n8483), .B2(n10406), .A(n8482), .ZN(n8484) );
  OAI21_X1 U10088 ( .B1(n8485), .B2(n9985), .A(n8484), .ZN(P2_U3199) );
  NOR2_X1 U10089 ( .A1(n8502), .A2(n8486), .ZN(n8488) );
  NAND2_X1 U10090 ( .A1(n8505), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8512) );
  OAI21_X1 U10091 ( .B1(n8505), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8512), .ZN(
        n8489) );
  NOR2_X1 U10092 ( .A1(n8490), .A2(n8489), .ZN(n8514) );
  AOI21_X1 U10093 ( .B1(n8490), .B2(n8489), .A(n8514), .ZN(n8511) );
  INV_X1 U10094 ( .A(n8491), .ZN(n8492) );
  MUX2_X1 U10095 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n4446), .Z(n8494) );
  NOR2_X1 U10096 ( .A1(n8495), .A2(n8494), .ZN(n8523) );
  INV_X1 U10097 ( .A(n8523), .ZN(n8496) );
  NAND2_X1 U10098 ( .A1(n8495), .A2(n8494), .ZN(n8521) );
  NAND2_X1 U10099 ( .A1(n8496), .A2(n8521), .ZN(n8498) );
  OAI21_X1 U10100 ( .B1(n8498), .B2(n8497), .A(n9996), .ZN(n8509) );
  NAND3_X1 U10101 ( .A1(n8498), .A2(n10406), .A3(n8505), .ZN(n8500) );
  OAI211_X1 U10102 ( .C1(n10082), .C2(n10005), .A(n8500), .B(n8499), .ZN(n8508) );
  NOR2_X1 U10103 ( .A1(n8502), .A2(n8501), .ZN(n8504) );
  NAND2_X1 U10104 ( .A1(n8505), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8516) );
  OAI21_X1 U10105 ( .B1(n8505), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8516), .ZN(
        n8506) );
  OAI21_X1 U10106 ( .B1(n8511), .B2(n9985), .A(n8510), .ZN(P2_U3200) );
  INV_X1 U10107 ( .A(n8512), .ZN(n8513) );
  NOR2_X1 U10108 ( .A1(n8514), .A2(n8513), .ZN(n8515) );
  XNOR2_X1 U10109 ( .A(n8533), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8526) );
  XNOR2_X1 U10110 ( .A(n8515), .B(n8526), .ZN(n8540) );
  INV_X1 U10111 ( .A(n8516), .ZN(n8517) );
  NOR2_X1 U10112 ( .A1(n8518), .A2(n8517), .ZN(n8520) );
  XNOR2_X1 U10113 ( .A(n8519), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8524) );
  XNOR2_X1 U10114 ( .A(n8520), .B(n8524), .ZN(n8538) );
  OAI21_X1 U10115 ( .B1(n8523), .B2(n8522), .A(n8521), .ZN(n8529) );
  INV_X1 U10116 ( .A(n8524), .ZN(n8527) );
  MUX2_X1 U10117 ( .A(n8527), .B(n8526), .S(n4446), .Z(n8528) );
  XNOR2_X1 U10118 ( .A(n8529), .B(n8528), .ZN(n8536) );
  OAI21_X1 U10119 ( .B1(n10005), .B2(n8531), .A(n8530), .ZN(n8532) );
  AOI21_X1 U10120 ( .B1(n8533), .B2(n10411), .A(n8532), .ZN(n8534) );
  OAI21_X1 U10121 ( .B1(n8536), .B2(n8535), .A(n8534), .ZN(n8537) );
  AOI21_X1 U10122 ( .B1(n8538), .B2(n10419), .A(n8537), .ZN(n8539) );
  OAI21_X1 U10123 ( .B1(n8540), .B2(n9985), .A(n8539), .ZN(P2_U3201) );
  NAND2_X1 U10124 ( .A1(n8756), .A2(n8708), .ZN(n8545) );
  INV_X1 U10125 ( .A(n8541), .ZN(n8542) );
  NOR2_X1 U10126 ( .A1(n8543), .A2(n8542), .ZN(n8813) );
  AOI21_X1 U10127 ( .B1(n8813), .B2(n8748), .A(n8544), .ZN(n8547) );
  OAI211_X1 U10128 ( .C1(n8748), .C2(n8546), .A(n8545), .B(n8547), .ZN(
        P2_U3202) );
  NAND2_X1 U10129 ( .A1(n8758), .A2(n8708), .ZN(n8548) );
  OAI211_X1 U10130 ( .C1(n8748), .C2(n8549), .A(n8548), .B(n8547), .ZN(
        P2_U3203) );
  INV_X1 U10131 ( .A(n8820), .ZN(n8561) );
  INV_X1 U10132 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8556) );
  XNOR2_X1 U10133 ( .A(n8551), .B(n8552), .ZN(n8555) );
  OAI22_X1 U10134 ( .A1(n8553), .A2(n8744), .B1(n8574), .B2(n8742), .ZN(n8554)
         );
  MUX2_X1 U10135 ( .A(n8556), .B(n8818), .S(n8748), .Z(n8560) );
  AOI22_X1 U10136 ( .A1(n8558), .A2(n8708), .B1(n8718), .B2(n8557), .ZN(n8559)
         );
  OAI211_X1 U10137 ( .C1(n8561), .C2(n8711), .A(n8560), .B(n8559), .ZN(
        P2_U3205) );
  INV_X1 U10138 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8567) );
  XNOR2_X1 U10139 ( .A(n4428), .B(n8563), .ZN(n8566) );
  AOI222_X1 U10140 ( .A1(n8731), .A2(n8566), .B1(n8565), .B2(n8726), .C1(n8564), .C2(n8728), .ZN(n8824) );
  MUX2_X1 U10141 ( .A(n8567), .B(n8824), .S(n8748), .Z(n8570) );
  AOI22_X1 U10142 ( .A1(n8826), .A2(n8708), .B1(n8718), .B2(n8568), .ZN(n8569)
         );
  OAI211_X1 U10143 ( .C1(n8829), .C2(n8711), .A(n8570), .B(n8569), .ZN(
        P2_U3206) );
  XNOR2_X1 U10144 ( .A(n8572), .B(n8571), .ZN(n8573) );
  OAI222_X1 U10145 ( .A1(n8742), .A2(n8594), .B1(n8744), .B2(n8574), .C1(n8740), .C2(n8573), .ZN(n8767) );
  AOI21_X1 U10146 ( .B1(n8718), .B2(n8575), .A(n8767), .ZN(n8580) );
  AOI22_X1 U10147 ( .A1(n8832), .A2(n8708), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n8752), .ZN(n8579) );
  XNOR2_X1 U10148 ( .A(n8577), .B(n8576), .ZN(n8833) );
  NAND2_X1 U10149 ( .A1(n8833), .A2(n8753), .ZN(n8578) );
  OAI211_X1 U10150 ( .C1(n8580), .C2(n8752), .A(n8579), .B(n8578), .ZN(
        P2_U3207) );
  XNOR2_X1 U10151 ( .A(n8581), .B(n8587), .ZN(n8582) );
  OAI222_X1 U10152 ( .A1(n8744), .A2(n8584), .B1(n8742), .B2(n8583), .C1(n8582), .C2(n8740), .ZN(n8836) );
  AOI21_X1 U10153 ( .B1(n8734), .B2(n8585), .A(n8836), .ZN(n8591) );
  AOI22_X1 U10154 ( .A1(n8586), .A2(n8718), .B1(n8752), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8590) );
  XNOR2_X1 U10155 ( .A(n8588), .B(n8587), .ZN(n8771) );
  NAND2_X1 U10156 ( .A1(n8771), .A2(n8753), .ZN(n8589) );
  OAI211_X1 U10157 ( .C1(n8591), .C2(n8752), .A(n8590), .B(n8589), .ZN(
        P2_U3208) );
  XNOR2_X1 U10158 ( .A(n8592), .B(n8597), .ZN(n8593) );
  OAI222_X1 U10159 ( .A1(n8742), .A2(n8595), .B1(n8744), .B2(n8594), .C1(n8740), .C2(n8593), .ZN(n8774) );
  AOI21_X1 U10160 ( .B1(n8734), .B2(n8843), .A(n8774), .ZN(n8601) );
  AOI22_X1 U10161 ( .A1(n8596), .A2(n8718), .B1(n8752), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8600) );
  XOR2_X1 U10162 ( .A(n8598), .B(n8597), .Z(n8844) );
  NAND2_X1 U10163 ( .A1(n8844), .A2(n8753), .ZN(n8599) );
  OAI211_X1 U10164 ( .C1(n8601), .C2(n8752), .A(n8600), .B(n8599), .ZN(
        P2_U3209) );
  XOR2_X1 U10165 ( .A(n8603), .B(n8602), .Z(n8851) );
  INV_X1 U10166 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8607) );
  XNOR2_X1 U10167 ( .A(n8604), .B(n8603), .ZN(n8606) );
  AOI222_X1 U10168 ( .A1(n8731), .A2(n8606), .B1(n8605), .B2(n8728), .C1(n8633), .C2(n8726), .ZN(n8847) );
  MUX2_X1 U10169 ( .A(n8607), .B(n8847), .S(n8748), .Z(n8610) );
  AOI22_X1 U10170 ( .A1(n6462), .A2(n8708), .B1(n8718), .B2(n8608), .ZN(n8609)
         );
  OAI211_X1 U10171 ( .C1(n8851), .C2(n8711), .A(n8610), .B(n8609), .ZN(
        P2_U3210) );
  XNOR2_X1 U10172 ( .A(n8612), .B(n8611), .ZN(n8854) );
  INV_X1 U10173 ( .A(n8854), .ZN(n8624) );
  INV_X1 U10174 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n10127) );
  NAND3_X1 U10175 ( .A1(n8613), .A2(n8615), .A3(n8614), .ZN(n8616) );
  NAND2_X1 U10176 ( .A1(n8617), .A2(n8616), .ZN(n8620) );
  AOI222_X1 U10177 ( .A1(n8731), .A2(n8620), .B1(n8619), .B2(n8726), .C1(n8618), .C2(n8728), .ZN(n8852) );
  MUX2_X1 U10178 ( .A(n10127), .B(n8852), .S(n8748), .Z(n8623) );
  AOI22_X1 U10179 ( .A1(n6458), .A2(n8708), .B1(n8718), .B2(n8621), .ZN(n8622)
         );
  OAI211_X1 U10180 ( .C1(n8624), .C2(n8711), .A(n8623), .B(n8622), .ZN(
        P2_U3211) );
  NAND2_X1 U10181 ( .A1(n8626), .A2(n8625), .ZN(n8627) );
  XOR2_X1 U10182 ( .A(n8629), .B(n8627), .Z(n8860) );
  INV_X1 U10183 ( .A(n8860), .ZN(n8640) );
  INV_X1 U10184 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8636) );
  AND2_X1 U10185 ( .A1(n8677), .A2(n8676), .ZN(n8674) );
  NOR2_X1 U10186 ( .A1(n8674), .A2(n8628), .ZN(n8656) );
  INV_X1 U10187 ( .A(n8657), .ZN(n8664) );
  NAND2_X1 U10188 ( .A1(n8656), .A2(n8664), .ZN(n8662) );
  NAND3_X1 U10189 ( .A1(n8662), .A2(n8643), .A3(n8644), .ZN(n8642) );
  INV_X1 U10190 ( .A(n8629), .ZN(n8631) );
  NAND3_X1 U10191 ( .A1(n8642), .A2(n8631), .A3(n8630), .ZN(n8632) );
  NAND2_X1 U10192 ( .A1(n8632), .A2(n8613), .ZN(n8635) );
  AOI222_X1 U10193 ( .A1(n8731), .A2(n8635), .B1(n8634), .B2(n8726), .C1(n8633), .C2(n8728), .ZN(n8857) );
  MUX2_X1 U10194 ( .A(n8636), .B(n8857), .S(n8748), .Z(n8639) );
  AOI22_X1 U10195 ( .A1(n8859), .A2(n8708), .B1(n8718), .B2(n8637), .ZN(n8638)
         );
  OAI211_X1 U10196 ( .C1(n8640), .C2(n8711), .A(n8639), .B(n8638), .ZN(
        P2_U3212) );
  XNOR2_X1 U10197 ( .A(n8641), .B(n8643), .ZN(n8866) );
  INV_X1 U10198 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8651) );
  INV_X1 U10199 ( .A(n8642), .ZN(n8646) );
  AOI21_X1 U10200 ( .B1(n8662), .B2(n8644), .A(n8643), .ZN(n8645) );
  NOR2_X1 U10201 ( .A1(n8646), .A2(n8645), .ZN(n8647) );
  OAI222_X1 U10202 ( .A1(n8744), .A2(n8649), .B1(n8742), .B2(n8648), .C1(n8740), .C2(n8647), .ZN(n8863) );
  INV_X1 U10203 ( .A(n8863), .ZN(n8650) );
  MUX2_X1 U10204 ( .A(n8651), .B(n8650), .S(n8748), .Z(n8655) );
  AOI22_X1 U10205 ( .A1(n8653), .A2(n8708), .B1(n8718), .B2(n8652), .ZN(n8654)
         );
  OAI211_X1 U10206 ( .C1(n8866), .C2(n8711), .A(n8655), .B(n8654), .ZN(
        P2_U3213) );
  INV_X1 U10207 ( .A(n8656), .ZN(n8658) );
  AOI21_X1 U10208 ( .B1(n8658), .B2(n8657), .A(n8740), .ZN(n8663) );
  OAI22_X1 U10209 ( .A1(n8660), .A2(n8744), .B1(n8659), .B2(n8742), .ZN(n8661)
         );
  AOI21_X1 U10210 ( .B1(n8663), .B2(n8662), .A(n8661), .ZN(n8791) );
  XNOR2_X1 U10211 ( .A(n8665), .B(n8664), .ZN(n8789) );
  AOI22_X1 U10212 ( .A1(n8752), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8718), .B2(
        n8666), .ZN(n8667) );
  OAI21_X1 U10213 ( .B1(n8668), .B2(n8720), .A(n8667), .ZN(n8669) );
  AOI21_X1 U10214 ( .B1(n8789), .B2(n8753), .A(n8669), .ZN(n8670) );
  OAI21_X1 U10215 ( .B1(n8791), .B2(n8752), .A(n8670), .ZN(P2_U3214) );
  INV_X1 U10216 ( .A(n8671), .ZN(n8672) );
  AOI21_X1 U10217 ( .B1(n8673), .B2(n8676), .A(n8672), .ZN(n8873) );
  INV_X1 U10218 ( .A(n8873), .ZN(n8684) );
  INV_X1 U10219 ( .A(n8674), .ZN(n8675) );
  OAI21_X1 U10220 ( .B1(n8677), .B2(n8676), .A(n8675), .ZN(n8679) );
  AOI222_X1 U10221 ( .A1(n8731), .A2(n8679), .B1(n8678), .B2(n8728), .C1(n8704), .C2(n8726), .ZN(n8870) );
  MUX2_X1 U10222 ( .A(n8680), .B(n8870), .S(n8748), .Z(n8683) );
  AOI22_X1 U10223 ( .A1(n8872), .A2(n8708), .B1(n8718), .B2(n8681), .ZN(n8682)
         );
  OAI211_X1 U10224 ( .C1(n8684), .C2(n8711), .A(n8683), .B(n8682), .ZN(
        P2_U3215) );
  XNOR2_X1 U10225 ( .A(n8686), .B(n8685), .ZN(n8688) );
  AOI222_X1 U10226 ( .A1(n8731), .A2(n8688), .B1(n8687), .B2(n8728), .C1(n8713), .C2(n8726), .ZN(n8798) );
  XNOR2_X1 U10227 ( .A(n8690), .B(n8689), .ZN(n8796) );
  NOR2_X1 U10228 ( .A1(n8691), .A2(n8720), .ZN(n8695) );
  OAI22_X1 U10229 ( .A1(n8748), .A2(n8693), .B1(n8692), .B2(n8745), .ZN(n8694)
         );
  AOI211_X1 U10230 ( .C1(n8796), .C2(n8753), .A(n8695), .B(n8694), .ZN(n8696)
         );
  OAI21_X1 U10231 ( .B1(n8798), .B2(n8752), .A(n8696), .ZN(P2_U3216) );
  INV_X1 U10232 ( .A(n8698), .ZN(n8700) );
  OAI21_X1 U10233 ( .B1(n8697), .B2(n8700), .A(n8699), .ZN(n8701) );
  XNOR2_X1 U10234 ( .A(n8701), .B(n8703), .ZN(n8883) );
  XOR2_X1 U10235 ( .A(n8703), .B(n8702), .Z(n8705) );
  AOI222_X1 U10236 ( .A1(n8731), .A2(n8705), .B1(n8704), .B2(n8728), .C1(n8729), .C2(n8726), .ZN(n8877) );
  OAI21_X1 U10237 ( .B1(n8706), .B2(n8745), .A(n8877), .ZN(n8707) );
  NAND2_X1 U10238 ( .A1(n8707), .A2(n8748), .ZN(n8710) );
  AOI22_X1 U10239 ( .A1(n8879), .A2(n8708), .B1(P2_REG2_REG_16__SCAN_IN), .B2(
        n8752), .ZN(n8709) );
  OAI211_X1 U10240 ( .C1(n8883), .C2(n8711), .A(n8710), .B(n8709), .ZN(
        P2_U3217) );
  XOR2_X1 U10241 ( .A(n8716), .B(n8712), .Z(n8715) );
  AOI222_X1 U10242 ( .A1(n8731), .A2(n8715), .B1(n8714), .B2(n8726), .C1(n8713), .C2(n8728), .ZN(n8806) );
  XOR2_X1 U10243 ( .A(n8697), .B(n8716), .Z(n8804) );
  AOI22_X1 U10244 ( .A1(n8752), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8718), .B2(
        n8717), .ZN(n8719) );
  OAI21_X1 U10245 ( .B1(n8721), .B2(n8720), .A(n8719), .ZN(n8722) );
  AOI21_X1 U10246 ( .B1(n8804), .B2(n8753), .A(n8722), .ZN(n8723) );
  OAI21_X1 U10247 ( .B1(n8806), .B2(n8752), .A(n8723), .ZN(P2_U3218) );
  NOR2_X1 U10248 ( .A1(n8745), .A2(n8724), .ZN(n8733) );
  XOR2_X1 U10249 ( .A(n8725), .B(n8736), .Z(n8730) );
  AOI222_X1 U10250 ( .A1(n8731), .A2(n8730), .B1(n8729), .B2(n8728), .C1(n8727), .C2(n8726), .ZN(n8885) );
  INV_X1 U10251 ( .A(n8885), .ZN(n8732) );
  AOI211_X1 U10252 ( .C1(n8734), .C2(n8887), .A(n8733), .B(n8732), .ZN(n8738)
         );
  XNOR2_X1 U10253 ( .A(n8735), .B(n8736), .ZN(n8890) );
  AOI22_X1 U10254 ( .A1(n8890), .A2(n8753), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n8752), .ZN(n8737) );
  OAI21_X1 U10255 ( .B1(n8738), .B2(n8752), .A(n8737), .ZN(P2_U3219) );
  XNOR2_X1 U10256 ( .A(n6443), .B(n8751), .ZN(n8739) );
  OAI222_X1 U10257 ( .A1(n8744), .A2(n8743), .B1(n8742), .B2(n8741), .C1(n8740), .C2(n8739), .ZN(n9775) );
  OAI22_X1 U10258 ( .A1(n9774), .A2(n8747), .B1(n8746), .B2(n8745), .ZN(n8749)
         );
  OAI21_X1 U10259 ( .B1(n9775), .B2(n8749), .A(n8748), .ZN(n8755) );
  XOR2_X1 U10260 ( .A(n8750), .B(n8751), .Z(n9777) );
  AOI22_X1 U10261 ( .A1(n9777), .A2(n8753), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n8752), .ZN(n8754) );
  NAND2_X1 U10262 ( .A1(n8755), .A2(n8754), .ZN(P2_U3220) );
  NAND2_X1 U10263 ( .A1(n8756), .A2(n8808), .ZN(n8757) );
  NAND2_X1 U10264 ( .A1(n8813), .A2(n10075), .ZN(n8759) );
  OAI211_X1 U10265 ( .C1(n10075), .C2(n7214), .A(n8757), .B(n8759), .ZN(
        P2_U3490) );
  NAND2_X1 U10266 ( .A1(n8758), .A2(n8808), .ZN(n8760) );
  OAI211_X1 U10267 ( .C1(n10075), .C2(n6476), .A(n8760), .B(n8759), .ZN(
        P2_U3489) );
  MUX2_X1 U10268 ( .A(n8761), .B(n8818), .S(n10075), .Z(n8763) );
  NAND2_X1 U10269 ( .A1(n8820), .A2(n8809), .ZN(n8762) );
  OAI211_X1 U10270 ( .C1(n8823), .C2(n8785), .A(n8763), .B(n8762), .ZN(
        P2_U3487) );
  INV_X1 U10271 ( .A(n8809), .ZN(n8802) );
  MUX2_X1 U10272 ( .A(n8764), .B(n8824), .S(n10075), .Z(n8766) );
  NAND2_X1 U10273 ( .A1(n8826), .A2(n8808), .ZN(n8765) );
  OAI211_X1 U10274 ( .C1(n8802), .C2(n8829), .A(n8766), .B(n8765), .ZN(
        P2_U3486) );
  INV_X1 U10275 ( .A(n8767), .ZN(n8830) );
  MUX2_X1 U10276 ( .A(n8768), .B(n8830), .S(n10075), .Z(n8770) );
  AOI22_X1 U10277 ( .A1(n8833), .A2(n8809), .B1(n8808), .B2(n8832), .ZN(n8769)
         );
  NAND2_X1 U10278 ( .A1(n8770), .A2(n8769), .ZN(P2_U3485) );
  MUX2_X1 U10279 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8836), .S(n10075), .Z(
        n8773) );
  INV_X1 U10280 ( .A(n8771), .ZN(n8838) );
  OAI22_X1 U10281 ( .A1(n8838), .A2(n8802), .B1(n8837), .B2(n8785), .ZN(n8772)
         );
  OR2_X1 U10282 ( .A1(n8773), .A2(n8772), .ZN(P2_U3484) );
  INV_X1 U10283 ( .A(n8774), .ZN(n8841) );
  MUX2_X1 U10284 ( .A(n8775), .B(n8841), .S(n10075), .Z(n8777) );
  AOI22_X1 U10285 ( .A1(n8844), .A2(n8809), .B1(n8808), .B2(n8843), .ZN(n8776)
         );
  NAND2_X1 U10286 ( .A1(n8777), .A2(n8776), .ZN(P2_U3483) );
  MUX2_X1 U10287 ( .A(n8778), .B(n8847), .S(n10075), .Z(n8780) );
  NAND2_X1 U10288 ( .A1(n6462), .A2(n8808), .ZN(n8779) );
  OAI211_X1 U10289 ( .C1(n8851), .C2(n8802), .A(n8780), .B(n8779), .ZN(
        P2_U3482) );
  MUX2_X1 U10290 ( .A(n10129), .B(n8852), .S(n10075), .Z(n8782) );
  AOI22_X1 U10291 ( .A1(n8854), .A2(n8809), .B1(n8808), .B2(n6458), .ZN(n8781)
         );
  NAND2_X1 U10292 ( .A1(n8782), .A2(n8781), .ZN(P2_U3481) );
  INV_X1 U10293 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n10282) );
  MUX2_X1 U10294 ( .A(n10282), .B(n8857), .S(n10075), .Z(n8784) );
  AOI22_X1 U10295 ( .A1(n8860), .A2(n8809), .B1(n8808), .B2(n8859), .ZN(n8783)
         );
  NAND2_X1 U10296 ( .A1(n8784), .A2(n8783), .ZN(P2_U3480) );
  MUX2_X1 U10297 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8863), .S(n10075), .Z(
        n8787) );
  OAI22_X1 U10298 ( .A1(n8866), .A2(n8802), .B1(n8865), .B2(n8785), .ZN(n8786)
         );
  OR2_X1 U10299 ( .A1(n8787), .A2(n8786), .ZN(P2_U3479) );
  AOI22_X1 U10300 ( .A1(n8789), .A2(n10020), .B1(n10061), .B2(n8788), .ZN(
        n8790) );
  NAND2_X1 U10301 ( .A1(n8791), .A2(n8790), .ZN(n8869) );
  MUX2_X1 U10302 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8869), .S(n10075), .Z(
        P2_U3478) );
  INV_X1 U10303 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8792) );
  MUX2_X1 U10304 ( .A(n8792), .B(n8870), .S(n10075), .Z(n8794) );
  AOI22_X1 U10305 ( .A1(n8873), .A2(n8809), .B1(n8808), .B2(n8872), .ZN(n8793)
         );
  NAND2_X1 U10306 ( .A1(n8794), .A2(n8793), .ZN(P2_U3477) );
  AOI22_X1 U10307 ( .A1(n8796), .A2(n10020), .B1(n10061), .B2(n8795), .ZN(
        n8797) );
  NAND2_X1 U10308 ( .A1(n8798), .A2(n8797), .ZN(n8876) );
  MUX2_X1 U10309 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8876), .S(n10075), .Z(
        P2_U3476) );
  MUX2_X1 U10310 ( .A(n8799), .B(n8877), .S(n10075), .Z(n8801) );
  NAND2_X1 U10311 ( .A1(n8879), .A2(n8808), .ZN(n8800) );
  OAI211_X1 U10312 ( .C1(n8883), .C2(n8802), .A(n8801), .B(n8800), .ZN(
        P2_U3475) );
  AOI22_X1 U10313 ( .A1(n8804), .A2(n10020), .B1(n10061), .B2(n8803), .ZN(
        n8805) );
  NAND2_X1 U10314 ( .A1(n8806), .A2(n8805), .ZN(n8884) );
  MUX2_X1 U10315 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8884), .S(n10075), .Z(
        P2_U3474) );
  MUX2_X1 U10316 ( .A(n8807), .B(n8885), .S(n10075), .Z(n8811) );
  AOI22_X1 U10317 ( .A1(n8890), .A2(n8809), .B1(n8808), .B2(n8887), .ZN(n8810)
         );
  NAND2_X1 U10318 ( .A1(n8811), .A2(n8810), .ZN(P2_U3473) );
  MUX2_X1 U10319 ( .A(n8812), .B(P2_REG1_REG_0__SCAN_IN), .S(n6533), .Z(
        P2_U3459) );
  NAND2_X1 U10320 ( .A1(n8813), .A2(n10064), .ZN(n8815) );
  NAND2_X1 U10321 ( .A1(n10062), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8814) );
  OAI211_X1 U10322 ( .C1(n4676), .C2(n8864), .A(n8815), .B(n8814), .ZN(
        P2_U3458) );
  NAND2_X1 U10323 ( .A1(n10062), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8816) );
  OAI211_X1 U10324 ( .C1(n8817), .C2(n8864), .A(n8816), .B(n8815), .ZN(
        P2_U3457) );
  INV_X1 U10325 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8819) );
  MUX2_X1 U10326 ( .A(n8819), .B(n8818), .S(n10064), .Z(n8822) );
  INV_X1 U10327 ( .A(n10020), .ZN(n10056) );
  OR2_X1 U10328 ( .A1(n10062), .A2(n10056), .ZN(n8882) );
  NAND2_X1 U10329 ( .A1(n8820), .A2(n8889), .ZN(n8821) );
  OAI211_X1 U10330 ( .C1(n8823), .C2(n8864), .A(n8822), .B(n8821), .ZN(
        P2_U3455) );
  INV_X1 U10331 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8825) );
  MUX2_X1 U10332 ( .A(n8825), .B(n8824), .S(n10064), .Z(n8828) );
  NAND2_X1 U10333 ( .A1(n8826), .A2(n8888), .ZN(n8827) );
  OAI211_X1 U10334 ( .C1(n8829), .C2(n8882), .A(n8828), .B(n8827), .ZN(
        P2_U3454) );
  INV_X1 U10335 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8831) );
  MUX2_X1 U10336 ( .A(n8831), .B(n8830), .S(n10064), .Z(n8835) );
  AOI22_X1 U10337 ( .A1(n8833), .A2(n8889), .B1(n8888), .B2(n8832), .ZN(n8834)
         );
  NAND2_X1 U10338 ( .A1(n8835), .A2(n8834), .ZN(P2_U3453) );
  MUX2_X1 U10339 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8836), .S(n10064), .Z(
        n8840) );
  OAI22_X1 U10340 ( .A1(n8838), .A2(n8882), .B1(n8837), .B2(n8864), .ZN(n8839)
         );
  OR2_X1 U10341 ( .A1(n8840), .A2(n8839), .ZN(P2_U3452) );
  INV_X1 U10342 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8842) );
  MUX2_X1 U10343 ( .A(n8842), .B(n8841), .S(n10064), .Z(n8846) );
  AOI22_X1 U10344 ( .A1(n8844), .A2(n8889), .B1(n8888), .B2(n8843), .ZN(n8845)
         );
  NAND2_X1 U10345 ( .A1(n8846), .A2(n8845), .ZN(P2_U3451) );
  INV_X1 U10346 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8848) );
  MUX2_X1 U10347 ( .A(n8848), .B(n8847), .S(n10064), .Z(n8850) );
  NAND2_X1 U10348 ( .A1(n6462), .A2(n8888), .ZN(n8849) );
  OAI211_X1 U10349 ( .C1(n8851), .C2(n8882), .A(n8850), .B(n8849), .ZN(
        P2_U3450) );
  INV_X1 U10350 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8853) );
  MUX2_X1 U10351 ( .A(n8853), .B(n8852), .S(n10064), .Z(n8856) );
  AOI22_X1 U10352 ( .A1(n8854), .A2(n8889), .B1(n8888), .B2(n6458), .ZN(n8855)
         );
  NAND2_X1 U10353 ( .A1(n8856), .A2(n8855), .ZN(P2_U3449) );
  INV_X1 U10354 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8858) );
  MUX2_X1 U10355 ( .A(n8858), .B(n8857), .S(n10064), .Z(n8862) );
  AOI22_X1 U10356 ( .A1(n8860), .A2(n8889), .B1(n8888), .B2(n8859), .ZN(n8861)
         );
  NAND2_X1 U10357 ( .A1(n8862), .A2(n8861), .ZN(P2_U3448) );
  MUX2_X1 U10358 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8863), .S(n10064), .Z(
        n8868) );
  OAI22_X1 U10359 ( .A1(n8866), .A2(n8882), .B1(n8865), .B2(n8864), .ZN(n8867)
         );
  OR2_X1 U10360 ( .A1(n8868), .A2(n8867), .ZN(P2_U3447) );
  MUX2_X1 U10361 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8869), .S(n10064), .Z(
        P2_U3446) );
  MUX2_X1 U10362 ( .A(n8871), .B(n8870), .S(n10064), .Z(n8875) );
  AOI22_X1 U10363 ( .A1(n8873), .A2(n8889), .B1(n8888), .B2(n8872), .ZN(n8874)
         );
  NAND2_X1 U10364 ( .A1(n8875), .A2(n8874), .ZN(P2_U3444) );
  MUX2_X1 U10365 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8876), .S(n10064), .Z(
        P2_U3441) );
  INV_X1 U10366 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8878) );
  MUX2_X1 U10367 ( .A(n8878), .B(n8877), .S(n10064), .Z(n8881) );
  NAND2_X1 U10368 ( .A1(n8879), .A2(n8888), .ZN(n8880) );
  OAI211_X1 U10369 ( .C1(n8883), .C2(n8882), .A(n8881), .B(n8880), .ZN(
        P2_U3438) );
  MUX2_X1 U10370 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8884), .S(n10064), .Z(
        P2_U3435) );
  MUX2_X1 U10371 ( .A(n8886), .B(n8885), .S(n10064), .Z(n8892) );
  AOI22_X1 U10372 ( .A1(n8890), .A2(n8889), .B1(n8888), .B2(n8887), .ZN(n8891)
         );
  NAND2_X1 U10373 ( .A1(n8892), .A2(n8891), .ZN(P2_U3432) );
  NAND3_X1 U10374 ( .A1(n8894), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8895) );
  OAI22_X1 U10375 ( .A1(n8893), .A2(n8895), .B1(n6672), .B2(n8899), .ZN(n8896)
         );
  AOI21_X1 U10376 ( .B1(n9765), .B2(n8897), .A(n8896), .ZN(n8898) );
  INV_X1 U10377 ( .A(n8898), .ZN(P2_U3264) );
  INV_X1 U10378 ( .A(n9054), .ZN(n9768) );
  OAI222_X1 U10379 ( .A1(P2_U3151), .A2(n6064), .B1(n8900), .B2(n9768), .C1(
        n10317), .C2(n8899), .ZN(P2_U3265) );
  INV_X1 U10380 ( .A(n8902), .ZN(n8903) );
  MUX2_X1 U10381 ( .A(n8903), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10382 ( .A1(n8905), .A2(n8904), .ZN(n8906) );
  XOR2_X1 U10383 ( .A(n8907), .B(n8906), .Z(n8914) );
  NOR2_X1 U10384 ( .A1(n8983), .A2(n9953), .ZN(n8908) );
  AOI211_X1 U10385 ( .C1(n9036), .C2(n9780), .A(n8909), .B(n8908), .ZN(n8910)
         );
  OAI21_X1 U10386 ( .B1(n9048), .B2(n8911), .A(n8910), .ZN(n8912) );
  AOI21_X1 U10387 ( .B1(n9956), .B2(n9050), .A(n8912), .ZN(n8913) );
  OAI21_X1 U10388 ( .B1(n8914), .B2(n9052), .A(n8913), .ZN(P1_U3215) );
  AOI21_X1 U10389 ( .B1(n8917), .B2(n8916), .A(n8915), .ZN(n8922) );
  XOR2_X1 U10390 ( .A(n8919), .B(n8920), .Z(n9010) );
  INV_X1 U10391 ( .A(n8918), .ZN(n9009) );
  NAND2_X1 U10392 ( .A1(n9010), .A2(n9009), .ZN(n9008) );
  OAI21_X1 U10393 ( .B1(n8920), .B2(n8919), .A(n9008), .ZN(n8921) );
  XOR2_X1 U10394 ( .A(n8922), .B(n8921), .Z(n8928) );
  OAI22_X1 U10395 ( .A1(n9058), .A2(n8983), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8923), .ZN(n8924) );
  AOI21_X1 U10396 ( .B1(n9556), .B2(n9036), .A(n8924), .ZN(n8925) );
  OAI21_X1 U10397 ( .B1(n9048), .B2(n9546), .A(n8925), .ZN(n8926) );
  AOI21_X1 U10398 ( .B1(n9665), .B2(n9050), .A(n8926), .ZN(n8927) );
  OAI21_X1 U10399 ( .B1(n8928), .B2(n9052), .A(n8927), .ZN(P1_U3216) );
  NAND2_X1 U10400 ( .A1(n8929), .A2(n9017), .ZN(n8932) );
  INV_X1 U10401 ( .A(n8930), .ZN(n8931) );
  AOI21_X1 U10402 ( .B1(n8933), .B2(n8932), .A(n8931), .ZN(n8938) );
  AOI22_X1 U10403 ( .A1(n9583), .A2(n9036), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n8935) );
  NAND2_X1 U10404 ( .A1(n9313), .A2(n9045), .ZN(n8934) );
  OAI211_X1 U10405 ( .C1(n9048), .C2(n9580), .A(n8935), .B(n8934), .ZN(n8936)
         );
  AOI21_X1 U10406 ( .B1(n9588), .B2(n9050), .A(n8936), .ZN(n8937) );
  OAI21_X1 U10407 ( .B1(n8938), .B2(n9052), .A(n8937), .ZN(P1_U3219) );
  XOR2_X1 U10408 ( .A(n8940), .B(n8939), .Z(n8946) );
  AOI22_X1 U10409 ( .A1(n9555), .A2(n9036), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n8943) );
  NAND2_X1 U10410 ( .A1(n8941), .A2(n8991), .ZN(n8942) );
  OAI211_X1 U10411 ( .C1(n9691), .C2(n8983), .A(n8943), .B(n8942), .ZN(n8944)
         );
  AOI21_X1 U10412 ( .B1(n9676), .B2(n9050), .A(n8944), .ZN(n8945) );
  OAI21_X1 U10413 ( .B1(n8946), .B2(n9052), .A(n8945), .ZN(P1_U3223) );
  INV_X1 U10414 ( .A(n8947), .ZN(n8949) );
  NOR3_X1 U10415 ( .A1(n8950), .A2(n8949), .A3(n8948), .ZN(n8952) );
  OAI21_X1 U10416 ( .B1(n8952), .B2(n8951), .A(n9031), .ZN(n8958) );
  AOI21_X1 U10417 ( .B1(n9045), .B2(n9317), .A(n8953), .ZN(n8954) );
  OAI21_X1 U10418 ( .B1(n9953), .B2(n9043), .A(n8954), .ZN(n8955) );
  AOI21_X1 U10419 ( .B1(n8956), .B2(n8991), .A(n8955), .ZN(n8957) );
  OAI211_X1 U10420 ( .C1(n8959), .C2(n9039), .A(n8958), .B(n8957), .ZN(
        P1_U3224) );
  AOI21_X1 U10421 ( .B1(n8962), .B2(n8961), .A(n9029), .ZN(n8969) );
  NOR2_X1 U10422 ( .A1(n8963), .A2(n9048), .ZN(n8966) );
  OAI22_X1 U10423 ( .A1(n9648), .A2(n8983), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8964), .ZN(n8965) );
  AOI211_X1 U10424 ( .C1(n9498), .C2(n9036), .A(n8966), .B(n8965), .ZN(n8968)
         );
  NAND2_X1 U10425 ( .A1(n9731), .A2(n9050), .ZN(n8967) );
  OAI211_X1 U10426 ( .C1(n8969), .C2(n9052), .A(n8968), .B(n8967), .ZN(
        P1_U3225) );
  OAI21_X1 U10427 ( .B1(n8972), .B2(n8971), .A(n8970), .ZN(n8973) );
  NAND2_X1 U10428 ( .A1(n8973), .A2(n9031), .ZN(n8978) );
  NAND2_X1 U10429 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9386) );
  OAI21_X1 U10430 ( .B1(n9043), .B2(n9603), .A(n9386), .ZN(n8976) );
  NOR2_X1 U10431 ( .A1(n9048), .A2(n8974), .ZN(n8975) );
  AOI211_X1 U10432 ( .C1(n9045), .C2(n9780), .A(n8976), .B(n8975), .ZN(n8977)
         );
  OAI211_X1 U10433 ( .C1(n9784), .C2(n9039), .A(n8978), .B(n8977), .ZN(
        P1_U3226) );
  INV_X1 U10434 ( .A(n9709), .ZN(n9619) );
  AND2_X1 U10435 ( .A1(n8970), .A2(n8979), .ZN(n8982) );
  OAI211_X1 U10436 ( .C1(n8982), .C2(n8981), .A(n9031), .B(n8980), .ZN(n8987)
         );
  NAND2_X1 U10437 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9405) );
  OAI21_X1 U10438 ( .B1(n8983), .B2(n9622), .A(n9405), .ZN(n8985) );
  NOR2_X1 U10439 ( .A1(n9048), .A2(n9615), .ZN(n8984) );
  AOI211_X1 U10440 ( .C1(n9036), .C2(n9313), .A(n8985), .B(n8984), .ZN(n8986)
         );
  OAI211_X1 U10441 ( .C1(n9619), .C2(n9039), .A(n8987), .B(n8986), .ZN(
        P1_U3228) );
  AOI21_X1 U10442 ( .B1(n8990), .B2(n8989), .A(n8988), .ZN(n8997) );
  AOI22_X1 U10443 ( .A1(n9311), .A2(n9045), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8993) );
  NAND2_X1 U10444 ( .A1(n9534), .A2(n8991), .ZN(n8992) );
  OAI211_X1 U10445 ( .C1(n8994), .C2(n9043), .A(n8993), .B(n8992), .ZN(n8995)
         );
  AOI21_X1 U10446 ( .B1(n9540), .B2(n9050), .A(n8995), .ZN(n8996) );
  OAI21_X1 U10447 ( .B1(n8997), .B2(n9052), .A(n8996), .ZN(P1_U3229) );
  OAI21_X1 U10448 ( .B1(n9000), .B2(n8999), .A(n8998), .ZN(n9001) );
  NAND2_X1 U10449 ( .A1(n9001), .A2(n9031), .ZN(n9007) );
  NOR2_X1 U10450 ( .A1(n9048), .A2(n9002), .ZN(n9005) );
  OAI22_X1 U10451 ( .A1(n9681), .A2(n9043), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9003), .ZN(n9004) );
  AOI211_X1 U10452 ( .C1(n9045), .C2(n9699), .A(n9005), .B(n9004), .ZN(n9006)
         );
  OAI211_X1 U10453 ( .C1(n9747), .C2(n9039), .A(n9007), .B(n9006), .ZN(
        P1_U3233) );
  OAI21_X1 U10454 ( .B1(n9010), .B2(n9009), .A(n9008), .ZN(n9011) );
  NAND2_X1 U10455 ( .A1(n9011), .A2(n9031), .ZN(n9016) );
  NOR2_X1 U10456 ( .A1(n9564), .A2(n9048), .ZN(n9014) );
  OAI22_X1 U10457 ( .A1(n9659), .A2(n9043), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9012), .ZN(n9013) );
  AOI211_X1 U10458 ( .C1(n9045), .C2(n9312), .A(n9014), .B(n9013), .ZN(n9015)
         );
  OAI211_X1 U10459 ( .C1(n9567), .C2(n9039), .A(n9016), .B(n9015), .ZN(
        P1_U3235) );
  NAND2_X1 U10460 ( .A1(n9018), .A2(n9017), .ZN(n9020) );
  XOR2_X1 U10461 ( .A(n9020), .B(n9019), .Z(n9025) );
  NAND2_X1 U10462 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9422) );
  OAI21_X1 U10463 ( .B1(n9680), .B2(n9043), .A(n9422), .ZN(n9021) );
  AOI21_X1 U10464 ( .B1(n9045), .B2(n9781), .A(n9021), .ZN(n9022) );
  OAI21_X1 U10465 ( .B1(n9048), .B2(n9596), .A(n9022), .ZN(n9023) );
  AOI21_X1 U10466 ( .B1(n9609), .B2(n9050), .A(n9023), .ZN(n9024) );
  OAI21_X1 U10467 ( .B1(n9025), .B2(n9052), .A(n9024), .ZN(P1_U3238) );
  INV_X1 U10468 ( .A(n9522), .ZN(n9728) );
  INV_X1 U10469 ( .A(n9026), .ZN(n9032) );
  OAI21_X1 U10470 ( .B1(n9029), .B2(n9028), .A(n9027), .ZN(n9030) );
  NAND3_X1 U10471 ( .A1(n9032), .A2(n9031), .A3(n9030), .ZN(n9038) );
  INV_X1 U10472 ( .A(n9523), .ZN(n9034) );
  AOI22_X1 U10473 ( .A1(n9530), .A2(n9045), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9033) );
  OAI21_X1 U10474 ( .B1(n9048), .B2(n9034), .A(n9033), .ZN(n9035) );
  AOI21_X1 U10475 ( .B1(n9036), .B2(n9515), .A(n9035), .ZN(n9037) );
  OAI211_X1 U10476 ( .C1(n9728), .C2(n9039), .A(n9038), .B(n9037), .ZN(
        P1_U3240) );
  AOI21_X1 U10477 ( .B1(n9041), .B2(n9040), .A(n4532), .ZN(n9053) );
  OAI21_X1 U10478 ( .B1(n9043), .B2(n9622), .A(n9042), .ZN(n9044) );
  AOI21_X1 U10479 ( .B1(n9045), .B2(n9314), .A(n9044), .ZN(n9046) );
  OAI21_X1 U10480 ( .B1(n9048), .B2(n9047), .A(n9046), .ZN(n9049) );
  AOI21_X1 U10481 ( .B1(n9151), .B2(n9050), .A(n9049), .ZN(n9051) );
  OAI21_X1 U10482 ( .B1(n9053), .B2(n9052), .A(n9051), .ZN(P1_U3241) );
  NAND2_X1 U10483 ( .A1(n9054), .A2(n5443), .ZN(n9056) );
  OR2_X1 U10484 ( .A1(n9075), .A2(n9770), .ZN(n9055) );
  INV_X1 U10485 ( .A(n9719), .ZN(n9465) );
  AND2_X1 U10486 ( .A1(n9465), .A2(n9310), .ZN(n9290) );
  INV_X1 U10487 ( .A(n9214), .ZN(n9057) );
  NOR2_X1 U10488 ( .A1(n9057), .A2(n9210), .ZN(n9286) );
  OR2_X1 U10489 ( .A1(n9740), .A2(n9058), .ZN(n9059) );
  AND2_X1 U10490 ( .A1(n9060), .A2(n9059), .ZN(n9197) );
  INV_X1 U10491 ( .A(n9197), .ZN(n9061) );
  NAND3_X1 U10492 ( .A1(n9205), .A2(n9196), .A3(n9061), .ZN(n9062) );
  AND2_X1 U10493 ( .A1(n9062), .A2(n9198), .ZN(n9063) );
  NAND2_X1 U10494 ( .A1(n9063), .A2(n9115), .ZN(n9068) );
  NAND2_X1 U10495 ( .A1(n9193), .A2(n9121), .ZN(n9179) );
  NOR2_X1 U10496 ( .A1(n9068), .A2(n9179), .ZN(n9278) );
  INV_X1 U10497 ( .A(n9114), .ZN(n9284) );
  AOI21_X1 U10498 ( .B1(n9278), .B2(n7901), .A(n9284), .ZN(n9072) );
  INV_X1 U10499 ( .A(n9116), .ZN(n9279) );
  NOR2_X1 U10500 ( .A1(n9211), .A2(n9279), .ZN(n9070) );
  INV_X1 U10501 ( .A(n9070), .ZN(n9071) );
  INV_X1 U10502 ( .A(n9205), .ZN(n9066) );
  AND2_X1 U10503 ( .A1(n9196), .A2(n9552), .ZN(n9184) );
  INV_X1 U10504 ( .A(n9184), .ZN(n9064) );
  NOR3_X1 U10505 ( .A1(n9066), .A2(n9065), .A3(n9064), .ZN(n9067) );
  OAI21_X1 U10506 ( .B1(n9068), .B2(n9067), .A(n9113), .ZN(n9069) );
  AND2_X1 U10507 ( .A1(n9110), .A2(n9213), .ZN(n9200) );
  INV_X1 U10508 ( .A(n9200), .ZN(n9203) );
  AOI21_X1 U10509 ( .B1(n9070), .B2(n9069), .A(n9203), .ZN(n9289) );
  OAI21_X1 U10510 ( .B1(n9072), .B2(n9071), .A(n9289), .ZN(n9073) );
  OAI21_X1 U10511 ( .B1(n9465), .B2(n9310), .A(n9215), .ZN(n9292) );
  AOI21_X1 U10512 ( .B1(n9286), .B2(n9073), .A(n9292), .ZN(n9074) );
  AOI21_X1 U10513 ( .B1(n9290), .B2(n9459), .A(n9074), .ZN(n9078) );
  NAND2_X1 U10514 ( .A1(n9716), .A2(n9459), .ZN(n9295) );
  OAI21_X1 U10515 ( .B1(n9465), .B2(n9459), .A(n9295), .ZN(n9077) );
  OAI21_X1 U10516 ( .B1(n9078), .B2(n9077), .A(n9076), .ZN(n9109) );
  INV_X1 U10517 ( .A(n9295), .ZN(n9230) );
  XOR2_X1 U10518 ( .A(n9310), .B(n9719), .Z(n9106) );
  INV_X1 U10519 ( .A(n9571), .ZN(n9561) );
  NAND2_X1 U10520 ( .A1(n9159), .A2(n9161), .ZN(n9795) );
  NOR4_X1 U10521 ( .A1(n5696), .A2(n9834), .A3(n9079), .A4(n9225), .ZN(n9081)
         );
  NAND2_X1 U10522 ( .A1(n9081), .A2(n9080), .ZN(n9084) );
  NOR4_X1 U10523 ( .A1(n9084), .A2(n9248), .A3(n9083), .A4(n9082), .ZN(n9085)
         );
  NAND4_X1 U10524 ( .A1(n9088), .A2(n9087), .A3(n9086), .A4(n9085), .ZN(n9089)
         );
  NOR4_X1 U10525 ( .A1(n9091), .A2(n9090), .A3(n9795), .A4(n9089), .ZN(n9092)
         );
  NAND4_X1 U10526 ( .A1(n9094), .A2(n9166), .A3(n9093), .A4(n9092), .ZN(n9095)
         );
  NOR4_X1 U10527 ( .A1(n9578), .A2(n9620), .A3(n9096), .A4(n9095), .ZN(n9098)
         );
  NAND4_X1 U10528 ( .A1(n9550), .A2(n9099), .A3(n9098), .A4(n9097), .ZN(n9101)
         );
  NOR4_X1 U10529 ( .A1(n9102), .A2(n9561), .A3(n9101), .A4(n9100), .ZN(n9103)
         );
  NAND4_X1 U10530 ( .A1(n9485), .A2(n9496), .A3(n9518), .A4(n9103), .ZN(n9104)
         );
  INV_X1 U10531 ( .A(n9224), .ZN(n9108) );
  INV_X1 U10532 ( .A(n9716), .ZN(n9220) );
  INV_X1 U10533 ( .A(n9459), .ZN(n9107) );
  NAND2_X1 U10534 ( .A1(n9220), .A2(n9107), .ZN(n9229) );
  INV_X1 U10535 ( .A(n9229), .ZN(n9294) );
  AOI21_X1 U10536 ( .B1(n9109), .B2(n9108), .A(n9294), .ZN(n9227) );
  OR2_X1 U10537 ( .A1(n9217), .A2(n9110), .ZN(n9112) );
  NAND2_X1 U10538 ( .A1(n9114), .A2(n9113), .ZN(n9204) );
  OR2_X1 U10539 ( .A1(n9204), .A2(n9115), .ZN(n9117) );
  AND2_X1 U10540 ( .A1(n9117), .A2(n9116), .ZN(n9208) );
  INV_X1 U10541 ( .A(n9217), .ZN(n9219) );
  NAND2_X1 U10542 ( .A1(n9123), .A2(n9118), .ZN(n9119) );
  OAI21_X1 U10543 ( .B1(n9120), .B2(n9219), .A(n9119), .ZN(n9122) );
  NAND2_X1 U10544 ( .A1(n9122), .A2(n9121), .ZN(n9125) );
  NAND3_X1 U10545 ( .A1(n9123), .A2(n9699), .A3(n9219), .ZN(n9124) );
  NAND2_X1 U10546 ( .A1(n9125), .A2(n9124), .ZN(n9192) );
  INV_X1 U10547 ( .A(n9268), .ZN(n9155) );
  AND2_X1 U10548 ( .A1(n9126), .A2(n9249), .ZN(n9132) );
  NAND3_X1 U10549 ( .A1(n9132), .A2(n9133), .A3(n9243), .ZN(n9130) );
  NAND2_X1 U10550 ( .A1(n9243), .A2(n9127), .ZN(n9128) );
  AOI21_X1 U10551 ( .B1(n9132), .B2(n9128), .A(n9248), .ZN(n9129) );
  OAI22_X1 U10552 ( .A1(n9131), .A2(n9130), .B1(n9217), .B2(n9129), .ZN(n9142)
         );
  INV_X1 U10553 ( .A(n9132), .ZN(n9134) );
  NAND2_X1 U10554 ( .A1(n9134), .A2(n9133), .ZN(n9137) );
  OAI211_X1 U10555 ( .C1(n9138), .C2(n9137), .A(n9136), .B(n9135), .ZN(n9139)
         );
  MUX2_X1 U10556 ( .A(n9140), .B(n9139), .S(n9217), .Z(n9141) );
  AOI21_X1 U10557 ( .B1(n9142), .B2(n9813), .A(n9141), .ZN(n9147) );
  NAND2_X1 U10558 ( .A1(n9148), .A2(n9143), .ZN(n9145) );
  MUX2_X1 U10559 ( .A(n9145), .B(n9144), .S(n9219), .Z(n9146) );
  OR2_X1 U10560 ( .A1(n9147), .A2(n9146), .ZN(n9157) );
  NAND2_X1 U10561 ( .A1(n9157), .A2(n9148), .ZN(n9149) );
  NAND2_X1 U10562 ( .A1(n9163), .A2(n9159), .ZN(n9259) );
  NAND4_X1 U10563 ( .A1(n9150), .A2(n9268), .A3(n9267), .A4(n9262), .ZN(n9154)
         );
  NOR2_X1 U10564 ( .A1(n9151), .A2(n9219), .ZN(n9152) );
  AOI21_X1 U10565 ( .B1(n9268), .B2(n9153), .A(n9152), .ZN(n9169) );
  NAND2_X1 U10566 ( .A1(n9157), .A2(n9156), .ZN(n9158) );
  NAND2_X1 U10567 ( .A1(n9158), .A2(n9794), .ZN(n9160) );
  NAND3_X1 U10568 ( .A1(n9160), .A2(n9251), .A3(n9159), .ZN(n9162) );
  NAND3_X1 U10569 ( .A1(n9162), .A2(n9161), .A3(n9258), .ZN(n9164) );
  NAND2_X1 U10570 ( .A1(n9164), .A2(n9163), .ZN(n9165) );
  NAND2_X1 U10571 ( .A1(n9165), .A2(n9257), .ZN(n9167) );
  NAND3_X1 U10572 ( .A1(n9167), .A2(n9166), .A3(n9261), .ZN(n9168) );
  NAND4_X1 U10573 ( .A1(n9168), .A2(n9217), .A3(n9265), .A4(n9264), .ZN(n9173)
         );
  INV_X1 U10574 ( .A(n9169), .ZN(n9170) );
  NAND2_X1 U10575 ( .A1(n9170), .A2(n9780), .ZN(n9172) );
  INV_X1 U10576 ( .A(n9273), .ZN(n9171) );
  AOI21_X1 U10577 ( .B1(n9173), .B2(n9172), .A(n9171), .ZN(n9175) );
  AND2_X1 U10578 ( .A1(n9188), .A2(n9176), .ZN(n9274) );
  NAND2_X1 U10579 ( .A1(n9187), .A2(n9274), .ZN(n9178) );
  AND2_X1 U10580 ( .A1(n9177), .A2(n9186), .ZN(n9275) );
  NAND2_X1 U10581 ( .A1(n9178), .A2(n9275), .ZN(n9180) );
  AOI21_X1 U10582 ( .B1(n9192), .B2(n9180), .A(n9179), .ZN(n9182) );
  AND2_X1 U10583 ( .A1(n9186), .A2(n9185), .ZN(n9270) );
  NAND3_X1 U10584 ( .A1(n9189), .A2(n9282), .A3(n9188), .ZN(n9191) );
  AOI21_X1 U10585 ( .B1(n9192), .B2(n9191), .A(n9190), .ZN(n9195) );
  INV_X1 U10586 ( .A(n9193), .ZN(n9194) );
  OAI21_X1 U10587 ( .B1(n9207), .B2(n9204), .A(n9283), .ZN(n9199) );
  NAND2_X1 U10588 ( .A1(n9200), .A2(n9199), .ZN(n9202) );
  INV_X1 U10589 ( .A(n9204), .ZN(n9206) );
  NAND3_X1 U10590 ( .A1(n9207), .A2(n9206), .A3(n9205), .ZN(n9209) );
  NAND2_X1 U10591 ( .A1(n9209), .A2(n9208), .ZN(n9212) );
  MUX2_X1 U10592 ( .A(n9215), .B(n9214), .S(n9219), .Z(n9216) );
  NAND3_X1 U10593 ( .A1(n9221), .A2(n9220), .A3(n9310), .ZN(n9222) );
  NAND3_X1 U10594 ( .A1(n9223), .A2(n9222), .A3(n9229), .ZN(n9228) );
  OAI21_X1 U10595 ( .B1(n9229), .B2(n5713), .A(n9228), .ZN(n9232) );
  AOI211_X1 U10596 ( .C1(n9230), .C2(n5685), .A(n5716), .B(n9236), .ZN(n9231)
         );
  NAND2_X1 U10597 ( .A1(n9232), .A2(n9231), .ZN(n9234) );
  NAND2_X1 U10598 ( .A1(n9234), .A2(n9233), .ZN(n9301) );
  INV_X1 U10599 ( .A(n9235), .ZN(n9246) );
  AOI21_X1 U10600 ( .B1(n9323), .B2(n9237), .A(n9236), .ZN(n9241) );
  NAND4_X1 U10601 ( .A1(n9241), .A2(n9240), .A3(n9239), .A4(n9238), .ZN(n9245)
         );
  INV_X1 U10602 ( .A(n9242), .ZN(n9244) );
  OAI211_X1 U10603 ( .C1(n9246), .C2(n9245), .A(n9244), .B(n9243), .ZN(n9250)
         );
  AOI211_X1 U10604 ( .C1(n9250), .C2(n9249), .A(n9248), .B(n9247), .ZN(n9253)
         );
  INV_X1 U10605 ( .A(n9251), .ZN(n9252) );
  NOR2_X1 U10606 ( .A1(n9253), .A2(n9252), .ZN(n9256) );
  AOI21_X1 U10607 ( .B1(n9256), .B2(n9255), .A(n9254), .ZN(n9260) );
  OAI211_X1 U10608 ( .C1(n9260), .C2(n9259), .A(n9258), .B(n9257), .ZN(n9263)
         );
  NAND3_X1 U10609 ( .A1(n9263), .A2(n9262), .A3(n9261), .ZN(n9266) );
  NAND3_X1 U10610 ( .A1(n9266), .A2(n9265), .A3(n9264), .ZN(n9269) );
  NAND3_X1 U10611 ( .A1(n9269), .A2(n9268), .A3(n9267), .ZN(n9272) );
  INV_X1 U10612 ( .A(n9270), .ZN(n9271) );
  AOI21_X1 U10613 ( .B1(n9273), .B2(n9272), .A(n9271), .ZN(n9277) );
  INV_X1 U10614 ( .A(n9274), .ZN(n9276) );
  OAI21_X1 U10615 ( .B1(n9277), .B2(n9276), .A(n9275), .ZN(n9281) );
  INV_X1 U10616 ( .A(n9278), .ZN(n9280) );
  AOI211_X1 U10617 ( .C1(n9282), .C2(n9281), .A(n9280), .B(n9279), .ZN(n9285)
         );
  OAI21_X1 U10618 ( .B1(n9285), .B2(n9284), .A(n9283), .ZN(n9288) );
  INV_X1 U10619 ( .A(n9286), .ZN(n9287) );
  AOI21_X1 U10620 ( .B1(n9289), .B2(n9288), .A(n9287), .ZN(n9293) );
  INV_X1 U10621 ( .A(n9290), .ZN(n9291) );
  OAI21_X1 U10622 ( .B1(n9293), .B2(n9292), .A(n9291), .ZN(n9296) );
  AOI21_X1 U10623 ( .B1(n9296), .B2(n9295), .A(n9294), .ZN(n9297) );
  XNOR2_X1 U10624 ( .A(n9297), .B(n5685), .ZN(n9299) );
  NOR3_X1 U10625 ( .A1(n9305), .A2(n9304), .A3(n9303), .ZN(n9307) );
  OAI21_X1 U10626 ( .B1(n5716), .B2(n9308), .A(P1_B_REG_SCAN_IN), .ZN(n9306)
         );
  OAI22_X1 U10627 ( .A1(n9309), .A2(n9308), .B1(n9307), .B2(n9306), .ZN(
        P1_U3242) );
  MUX2_X1 U10628 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9310), .S(n9324), .Z(
        P1_U3584) );
  MUX2_X1 U10629 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9482), .S(n9324), .Z(
        P1_U3583) );
  MUX2_X1 U10630 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9497), .S(n9324), .Z(
        P1_U3582) );
  MUX2_X1 U10631 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9515), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10632 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9498), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10633 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9530), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10634 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9556), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10635 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9311), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10636 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9555), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10637 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9312), .S(n9324), .Z(
        P1_U3575) );
  MUX2_X1 U10638 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9313), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10639 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9781), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10640 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9780), .S(n9324), .Z(
        P1_U3569) );
  MUX2_X1 U10641 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9314), .S(n9324), .Z(
        P1_U3568) );
  MUX2_X1 U10642 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9315), .S(n9324), .Z(
        P1_U3567) );
  MUX2_X1 U10643 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9316), .S(n9324), .Z(
        P1_U3566) );
  MUX2_X1 U10644 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9317), .S(n9324), .Z(
        P1_U3565) );
  MUX2_X1 U10645 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9318), .S(n9324), .Z(
        P1_U3564) );
  MUX2_X1 U10646 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9319), .S(n9324), .Z(
        P1_U3563) );
  MUX2_X1 U10647 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9917), .S(n9324), .Z(
        P1_U3562) );
  MUX2_X1 U10648 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9320), .S(n9324), .Z(
        P1_U3561) );
  MUX2_X1 U10649 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9890), .S(n9324), .Z(
        P1_U3560) );
  MUX2_X1 U10650 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9321), .S(n9324), .Z(
        P1_U3559) );
  MUX2_X1 U10651 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9829), .S(n9324), .Z(
        P1_U3558) );
  MUX2_X1 U10652 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9322), .S(n9324), .Z(
        P1_U3557) );
  MUX2_X1 U10653 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n4429), .S(n9324), .Z(
        P1_U3556) );
  MUX2_X1 U10654 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9323), .S(n9324), .Z(
        P1_U3555) );
  MUX2_X1 U10655 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9325), .S(n9324), .Z(
        P1_U3554) );
  AOI211_X1 U10656 ( .C1(n9328), .C2(n9327), .A(n9326), .B(n9428), .ZN(n9329)
         );
  INV_X1 U10657 ( .A(n9329), .ZN(n9339) );
  INV_X1 U10658 ( .A(n9445), .ZN(n9413) );
  INV_X1 U10659 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9330) );
  OAI22_X1 U10660 ( .A1(n9455), .A2(n9330), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9845), .ZN(n9331) );
  AOI21_X1 U10661 ( .B1(n9332), .B2(n9413), .A(n9331), .ZN(n9338) );
  NOR2_X1 U10662 ( .A1(n9333), .A2(n5771), .ZN(n9335) );
  OAI211_X1 U10663 ( .C1(n9336), .C2(n9335), .A(n9443), .B(n9334), .ZN(n9337)
         );
  NAND3_X1 U10664 ( .A1(n9339), .A2(n9338), .A3(n9337), .ZN(P1_U3244) );
  NOR2_X1 U10665 ( .A1(n9445), .A2(n9340), .ZN(n9341) );
  AOI211_X1 U10666 ( .C1(n9433), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n9342), .B(
        n9341), .ZN(n9352) );
  OAI211_X1 U10667 ( .C1(n9345), .C2(n9344), .A(n9450), .B(n9343), .ZN(n9351)
         );
  AOI211_X1 U10668 ( .C1(n9348), .C2(n9347), .A(n9346), .B(n9446), .ZN(n9349)
         );
  INV_X1 U10669 ( .A(n9349), .ZN(n9350) );
  NAND3_X1 U10670 ( .A1(n9352), .A2(n9351), .A3(n9350), .ZN(P1_U3246) );
  NOR2_X1 U10671 ( .A1(n9445), .A2(n9353), .ZN(n9354) );
  AOI211_X1 U10672 ( .C1(n9433), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n9355), .B(
        n9354), .ZN(n9364) );
  OAI211_X1 U10673 ( .C1(n9358), .C2(n9357), .A(n9450), .B(n9356), .ZN(n9363)
         );
  XOR2_X1 U10674 ( .A(n9360), .B(n9359), .Z(n9361) );
  NAND2_X1 U10675 ( .A1(n9443), .A2(n9361), .ZN(n9362) );
  NAND4_X1 U10676 ( .A1(n9365), .A2(n9364), .A3(n9363), .A4(n9362), .ZN(
        P1_U3247) );
  NOR2_X1 U10677 ( .A1(n9445), .A2(n9366), .ZN(n9367) );
  AOI211_X1 U10678 ( .C1(n9433), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n9368), .B(
        n9367), .ZN(n9377) );
  OAI211_X1 U10679 ( .C1(n9371), .C2(n9370), .A(n9369), .B(n9450), .ZN(n9376)
         );
  OAI211_X1 U10680 ( .C1(n9374), .C2(n9373), .A(n9443), .B(n9372), .ZN(n9375)
         );
  NAND3_X1 U10681 ( .A1(n9377), .A2(n9376), .A3(n9375), .ZN(P1_U3248) );
  NOR2_X1 U10682 ( .A1(n9397), .A2(n9378), .ZN(n9379) );
  AOI21_X1 U10683 ( .B1(n9397), .B2(n9378), .A(n9379), .ZN(n9385) );
  NAND2_X1 U10684 ( .A1(n9381), .A2(n9380), .ZN(n9383) );
  NAND2_X1 U10685 ( .A1(n9383), .A2(n9382), .ZN(n9384) );
  NOR2_X1 U10686 ( .A1(n9384), .A2(n9385), .ZN(n9401) );
  AOI21_X1 U10687 ( .B1(n9385), .B2(n9384), .A(n9401), .ZN(n9400) );
  INV_X1 U10688 ( .A(n9386), .ZN(n9396) );
  NOR2_X1 U10689 ( .A1(n9388), .A2(n9387), .ZN(n9390) );
  NAND2_X1 U10690 ( .A1(n9397), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9406) );
  OR2_X1 U10691 ( .A1(n9397), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9391) );
  NAND2_X1 U10692 ( .A1(n9406), .A2(n9391), .ZN(n9393) );
  INV_X1 U10693 ( .A(n9407), .ZN(n9392) );
  AOI211_X1 U10694 ( .C1(n9394), .C2(n9393), .A(n9392), .B(n9428), .ZN(n9395)
         );
  AOI211_X1 U10695 ( .C1(n9433), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9396), .B(
        n9395), .ZN(n9399) );
  NAND2_X1 U10696 ( .A1(n9413), .A2(n9397), .ZN(n9398) );
  OAI211_X1 U10697 ( .C1(n9400), .C2(n9446), .A(n9399), .B(n9398), .ZN(
        P1_U3259) );
  AOI21_X1 U10698 ( .B1(n9378), .B2(n9402), .A(n9401), .ZN(n9404) );
  XNOR2_X1 U10699 ( .A(n9423), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9403) );
  NOR2_X1 U10700 ( .A1(n9404), .A2(n9403), .ZN(n9419) );
  AOI21_X1 U10701 ( .B1(n9404), .B2(n9403), .A(n9419), .ZN(n9416) );
  INV_X1 U10702 ( .A(n9405), .ZN(n9412) );
  XNOR2_X1 U10703 ( .A(n9423), .B(n9408), .ZN(n9409) );
  NAND2_X1 U10704 ( .A1(n9410), .A2(n9409), .ZN(n9425) );
  AOI221_X1 U10705 ( .B1(n9410), .B2(n9425), .C1(n9409), .C2(n9425), .A(n9428), 
        .ZN(n9411) );
  AOI211_X1 U10706 ( .C1(n9433), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n9412), .B(
        n9411), .ZN(n9415) );
  NAND2_X1 U10707 ( .A1(n9413), .A2(n9423), .ZN(n9414) );
  OAI211_X1 U10708 ( .C1(n9416), .C2(n9446), .A(n9415), .B(n9414), .ZN(
        P1_U3260) );
  NOR2_X1 U10709 ( .A1(n9423), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9418) );
  XNOR2_X1 U10710 ( .A(n9441), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9417) );
  NOR3_X1 U10711 ( .A1(n9419), .A2(n9418), .A3(n9417), .ZN(n9440) );
  INV_X1 U10712 ( .A(n9440), .ZN(n9421) );
  OAI21_X1 U10713 ( .B1(n9419), .B2(n9418), .A(n9417), .ZN(n9420) );
  NAND3_X1 U10714 ( .A1(n9421), .A2(n9443), .A3(n9420), .ZN(n9435) );
  INV_X1 U10715 ( .A(n9422), .ZN(n9432) );
  OR2_X1 U10716 ( .A1(n9423), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9424) );
  NAND2_X1 U10717 ( .A1(n9425), .A2(n9424), .ZN(n9430) );
  INV_X1 U10718 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9597) );
  OR2_X1 U10719 ( .A1(n9441), .A2(n9597), .ZN(n9427) );
  NAND2_X1 U10720 ( .A1(n9441), .A2(n9597), .ZN(n9426) );
  AND2_X1 U10721 ( .A1(n9427), .A2(n9426), .ZN(n9429) );
  NOR2_X1 U10722 ( .A1(n9430), .A2(n9429), .ZN(n9438) );
  AOI211_X1 U10723 ( .C1(n9430), .C2(n9429), .A(n9438), .B(n9428), .ZN(n9431)
         );
  AOI211_X1 U10724 ( .C1(n9433), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9432), .B(
        n9431), .ZN(n9434) );
  OAI211_X1 U10725 ( .C1(n9445), .C2(n9436), .A(n9435), .B(n9434), .ZN(
        P1_U3261) );
  AND2_X1 U10726 ( .A1(n9441), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9437) );
  XNOR2_X1 U10727 ( .A(n9439), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9449) );
  INV_X1 U10728 ( .A(n9449), .ZN(n9444) );
  AOI21_X1 U10729 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n9441), .A(n9440), .ZN(
        n9442) );
  XNOR2_X1 U10730 ( .A(n9442), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9447) );
  AOI22_X1 U10731 ( .A1(n9444), .A2(n9450), .B1(n9447), .B2(n9443), .ZN(n9452)
         );
  OAI21_X1 U10732 ( .B1(n9447), .B2(n9446), .A(n9445), .ZN(n9448) );
  AOI21_X1 U10733 ( .B1(n9450), .B2(n9449), .A(n9448), .ZN(n9451) );
  MUX2_X1 U10734 ( .A(n9452), .B(n9451), .S(n5685), .Z(n9454) );
  NAND2_X1 U10735 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9453) );
  OAI211_X1 U10736 ( .C1(n4652), .C2(n9455), .A(n9454), .B(n9453), .ZN(
        P1_U3262) );
  XNOR2_X1 U10737 ( .A(n9716), .B(n9463), .ZN(n9456) );
  NAND2_X1 U10738 ( .A1(n9456), .A2(n9837), .ZN(n9630) );
  INV_X1 U10739 ( .A(n9457), .ZN(n9458) );
  NAND2_X1 U10740 ( .A1(n9459), .A2(n9458), .ZN(n9633) );
  NOR2_X1 U10741 ( .A1(n9633), .A2(n9857), .ZN(n9467) );
  NOR2_X1 U10742 ( .A1(n9716), .A2(n9618), .ZN(n9460) );
  AOI211_X1 U10743 ( .C1(n9857), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9467), .B(
        n9460), .ZN(n9461) );
  OAI21_X1 U10744 ( .B1(n9630), .B2(n9606), .A(n9461), .ZN(P1_U3263) );
  AOI21_X1 U10745 ( .B1(n9719), .B2(n9462), .A(n9822), .ZN(n9464) );
  NAND2_X1 U10746 ( .A1(n9464), .A2(n9463), .ZN(n9634) );
  NOR2_X1 U10747 ( .A1(n9465), .A2(n9618), .ZN(n9466) );
  AOI211_X1 U10748 ( .C1(n9857), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9467), .B(
        n9466), .ZN(n9468) );
  OAI21_X1 U10749 ( .B1(n9634), .B2(n9606), .A(n9468), .ZN(P1_U3264) );
  INV_X1 U10750 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9470) );
  OAI22_X1 U10751 ( .A1(n9471), .A2(n9846), .B1(n9470), .B2(n9598), .ZN(n9472)
         );
  AOI21_X1 U10752 ( .B1(n9473), .B2(n7133), .A(n9472), .ZN(n9474) );
  OAI21_X1 U10753 ( .B1(n9475), .B2(n9606), .A(n9474), .ZN(n9476) );
  AOI21_X1 U10754 ( .B1(n9469), .B2(n9841), .A(n9476), .ZN(n9477) );
  OAI21_X1 U10755 ( .B1(n9478), .B2(n9857), .A(n9477), .ZN(P1_U3356) );
  OAI21_X1 U10756 ( .B1(n9485), .B2(n9480), .A(n9479), .ZN(n9481) );
  NAND2_X1 U10757 ( .A1(n9481), .A2(n9887), .ZN(n9484) );
  AOI22_X1 U10758 ( .A1(n9482), .A2(n9891), .B1(n9515), .B2(n9918), .ZN(n9483)
         );
  INV_X1 U10759 ( .A(n9485), .ZN(n9486) );
  XNOR2_X1 U10760 ( .A(n9487), .B(n9486), .ZN(n9638) );
  NAND2_X1 U10761 ( .A1(n9638), .A2(n9841), .ZN(n9493) );
  AOI211_X1 U10762 ( .C1(n9488), .C2(n9500), .A(n9822), .B(n5693), .ZN(n9637)
         );
  AOI22_X1 U10763 ( .A1(n9489), .A2(n9820), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9857), .ZN(n9490) );
  OAI21_X1 U10764 ( .B1(n9723), .B2(n9618), .A(n9490), .ZN(n9491) );
  AOI21_X1 U10765 ( .B1(n9637), .B2(n9851), .A(n9491), .ZN(n9492) );
  OAI211_X1 U10766 ( .C1(n4471), .C2(n9857), .A(n9493), .B(n9492), .ZN(
        P1_U3265) );
  OAI21_X1 U10767 ( .B1(n9496), .B2(n9495), .A(n9494), .ZN(n9499) );
  AOI222_X1 U10768 ( .A1(n9887), .A2(n9499), .B1(n9498), .B2(n9918), .C1(n9497), .C2(n9891), .ZN(n9642) );
  INV_X1 U10769 ( .A(n9520), .ZN(n9502) );
  INV_X1 U10770 ( .A(n9500), .ZN(n9501) );
  AOI211_X1 U10771 ( .C1(n4847), .C2(n9502), .A(n9822), .B(n9501), .ZN(n9640)
         );
  AOI22_X1 U10772 ( .A1(n9503), .A2(n9820), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9857), .ZN(n9504) );
  OAI21_X1 U10773 ( .B1(n9505), .B2(n9618), .A(n9504), .ZN(n9506) );
  AOI21_X1 U10774 ( .B1(n9640), .B2(n9851), .A(n9506), .ZN(n9511) );
  OAI21_X1 U10775 ( .B1(n9509), .B2(n9508), .A(n9507), .ZN(n9639) );
  NAND2_X1 U10776 ( .A1(n9639), .A2(n9841), .ZN(n9510) );
  OAI211_X1 U10777 ( .C1(n9642), .C2(n9857), .A(n9511), .B(n9510), .ZN(
        P1_U3266) );
  OAI21_X1 U10778 ( .B1(n9518), .B2(n9513), .A(n9512), .ZN(n9514) );
  NAND2_X1 U10779 ( .A1(n9514), .A2(n9887), .ZN(n9517) );
  AOI22_X1 U10780 ( .A1(n9515), .A2(n9891), .B1(n9918), .B2(n9530), .ZN(n9516)
         );
  NAND2_X1 U10781 ( .A1(n9517), .A2(n9516), .ZN(n9644) );
  INV_X1 U10782 ( .A(n9644), .ZN(n9528) );
  XNOR2_X1 U10783 ( .A(n9519), .B(n9518), .ZN(n9646) );
  NAND2_X1 U10784 ( .A1(n9646), .A2(n9841), .ZN(n9527) );
  AOI211_X1 U10785 ( .C1(n9522), .C2(n9521), .A(n9822), .B(n9520), .ZN(n9645)
         );
  AOI22_X1 U10786 ( .A1(n9523), .A2(n9820), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9857), .ZN(n9524) );
  OAI21_X1 U10787 ( .B1(n9728), .B2(n9618), .A(n9524), .ZN(n9525) );
  AOI21_X1 U10788 ( .B1(n9645), .B2(n9851), .A(n9525), .ZN(n9526) );
  OAI211_X1 U10789 ( .C1(n9857), .C2(n9528), .A(n9527), .B(n9526), .ZN(
        P1_U3267) );
  XNOR2_X1 U10790 ( .A(n9529), .B(n9532), .ZN(n9531) );
  AOI22_X1 U10791 ( .A1(n9531), .A2(n9887), .B1(n9891), .B2(n9530), .ZN(n9658)
         );
  XNOR2_X1 U10792 ( .A(n9533), .B(n9532), .ZN(n9661) );
  NAND2_X1 U10793 ( .A1(n9661), .A2(n9841), .ZN(n9542) );
  AOI22_X1 U10794 ( .A1(n9534), .A2(n9820), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9857), .ZN(n9535) );
  OAI21_X1 U10795 ( .B1(n9659), .B2(n9602), .A(n9535), .ZN(n9539) );
  INV_X1 U10796 ( .A(n9540), .ZN(n9736) );
  INV_X1 U10797 ( .A(n9536), .ZN(n9545) );
  OAI211_X1 U10798 ( .C1(n9736), .C2(n9545), .A(n9537), .B(n9837), .ZN(n9657)
         );
  NOR2_X1 U10799 ( .A1(n9657), .A2(n9606), .ZN(n9538) );
  AOI211_X1 U10800 ( .C1(n7133), .C2(n9540), .A(n9539), .B(n9538), .ZN(n9541)
         );
  OAI211_X1 U10801 ( .C1(n9857), .C2(n9658), .A(n9542), .B(n9541), .ZN(
        P1_U3269) );
  XNOR2_X1 U10802 ( .A(n9543), .B(n9550), .ZN(n9668) );
  INV_X1 U10803 ( .A(n9544), .ZN(n9565) );
  AOI211_X1 U10804 ( .C1(n9665), .C2(n9565), .A(n9822), .B(n9545), .ZN(n9664)
         );
  INV_X1 U10805 ( .A(n9546), .ZN(n9547) );
  AOI22_X1 U10806 ( .A1(n9547), .A2(n9820), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9857), .ZN(n9548) );
  OAI21_X1 U10807 ( .B1(n9549), .B2(n9618), .A(n9548), .ZN(n9559) );
  INV_X1 U10808 ( .A(n9550), .ZN(n9551) );
  NAND3_X1 U10809 ( .A1(n9570), .A2(n9552), .A3(n9551), .ZN(n9553) );
  NAND2_X1 U10810 ( .A1(n9554), .A2(n9553), .ZN(n9557) );
  AOI222_X1 U10811 ( .A1(n9887), .A2(n9557), .B1(n9556), .B2(n9891), .C1(n9555), .C2(n9918), .ZN(n9667) );
  NOR2_X1 U10812 ( .A1(n9667), .A2(n9857), .ZN(n9558) );
  AOI211_X1 U10813 ( .C1(n9664), .C2(n9851), .A(n9559), .B(n9558), .ZN(n9560)
         );
  OAI21_X1 U10814 ( .B1(n9629), .B2(n9668), .A(n9560), .ZN(P1_U3270) );
  XNOR2_X1 U10815 ( .A(n9562), .B(n9561), .ZN(n9671) );
  OAI22_X1 U10816 ( .A1(n9564), .A2(n9846), .B1(n9563), .B2(n9598), .ZN(n9569)
         );
  OAI211_X1 U10817 ( .C1(n9567), .C2(n9566), .A(n9565), .B(n9837), .ZN(n9669)
         );
  NOR2_X1 U10818 ( .A1(n9669), .A2(n9606), .ZN(n9568) );
  AOI211_X1 U10819 ( .C1(n7133), .C2(n9740), .A(n9569), .B(n9568), .ZN(n9576)
         );
  OAI21_X1 U10820 ( .B1(n9572), .B2(n9571), .A(n9570), .ZN(n9574) );
  OAI22_X1 U10821 ( .A1(n9659), .A2(n9950), .B1(n9681), .B2(n9952), .ZN(n9573)
         );
  AOI21_X1 U10822 ( .B1(n9574), .B2(n9887), .A(n9573), .ZN(n9670) );
  OR2_X1 U10823 ( .A1(n9670), .A2(n9857), .ZN(n9575) );
  OAI211_X1 U10824 ( .C1(n9671), .C2(n9629), .A(n9576), .B(n9575), .ZN(
        P1_U3271) );
  XNOR2_X1 U10825 ( .A(n9577), .B(n9578), .ZN(n9695) );
  XNOR2_X1 U10826 ( .A(n9579), .B(n9578), .ZN(n9697) );
  NAND2_X1 U10827 ( .A1(n9697), .A2(n9841), .ZN(n9590) );
  OAI22_X1 U10828 ( .A1(n9598), .A2(n9581), .B1(n9580), .B2(n9846), .ZN(n9582)
         );
  AOI21_X1 U10829 ( .B1(n9583), .B2(n9600), .A(n9582), .ZN(n9584) );
  OAI21_X1 U10830 ( .B1(n9690), .B2(n9602), .A(n9584), .ZN(n9587) );
  OAI211_X1 U10831 ( .C1(n9751), .C2(n9604), .A(n9837), .B(n9585), .ZN(n9693)
         );
  NOR2_X1 U10832 ( .A1(n9693), .A2(n9606), .ZN(n9586) );
  AOI211_X1 U10833 ( .C1(n7133), .C2(n9588), .A(n9587), .B(n9586), .ZN(n9589)
         );
  OAI211_X1 U10834 ( .C1(n9695), .C2(n9612), .A(n9590), .B(n9589), .ZN(
        P1_U3274) );
  OAI21_X1 U10835 ( .B1(n9592), .B2(n9594), .A(n9591), .ZN(n9593) );
  INV_X1 U10836 ( .A(n9593), .ZN(n9702) );
  XNOR2_X1 U10837 ( .A(n9595), .B(n9594), .ZN(n9704) );
  NAND2_X1 U10838 ( .A1(n9704), .A2(n9841), .ZN(n9611) );
  OAI22_X1 U10839 ( .A1(n9598), .A2(n9597), .B1(n9596), .B2(n9846), .ZN(n9599)
         );
  AOI21_X1 U10840 ( .B1(n9600), .B2(n9699), .A(n9599), .ZN(n9601) );
  OAI21_X1 U10841 ( .B1(n9603), .B2(n9602), .A(n9601), .ZN(n9608) );
  INV_X1 U10842 ( .A(n4469), .ZN(n9614) );
  INV_X1 U10843 ( .A(n9609), .ZN(n9755) );
  OAI211_X1 U10844 ( .C1(n9614), .C2(n9755), .A(n9837), .B(n9605), .ZN(n9700)
         );
  NOR2_X1 U10845 ( .A1(n9700), .A2(n9606), .ZN(n9607) );
  AOI211_X1 U10846 ( .C1(n7133), .C2(n9609), .A(n9608), .B(n9607), .ZN(n9610)
         );
  OAI211_X1 U10847 ( .C1(n9702), .C2(n9612), .A(n9611), .B(n9610), .ZN(
        P1_U3275) );
  XNOR2_X1 U10848 ( .A(n9613), .B(n9620), .ZN(n9712) );
  AOI211_X1 U10849 ( .C1(n9709), .C2(n4530), .A(n9822), .B(n9614), .ZN(n9708)
         );
  INV_X1 U10850 ( .A(n9615), .ZN(n9616) );
  AOI22_X1 U10851 ( .A1(n9857), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9616), .B2(
        n9820), .ZN(n9617) );
  OAI21_X1 U10852 ( .B1(n9619), .B2(n9618), .A(n9617), .ZN(n9627) );
  AOI21_X1 U10853 ( .B1(n9621), .B2(n9620), .A(n9933), .ZN(n9625) );
  OAI22_X1 U10854 ( .A1(n9690), .A2(n9950), .B1(n9622), .B2(n9952), .ZN(n9623)
         );
  AOI21_X1 U10855 ( .B1(n9625), .B2(n9624), .A(n9623), .ZN(n9711) );
  NOR2_X1 U10856 ( .A1(n9711), .A2(n9857), .ZN(n9626) );
  AOI211_X1 U10857 ( .C1(n9708), .C2(n9851), .A(n9627), .B(n9626), .ZN(n9628)
         );
  OAI21_X1 U10858 ( .B1(n9629), .B2(n9712), .A(n9628), .ZN(P1_U3276) );
  MUX2_X1 U10859 ( .A(n9631), .B(n9713), .S(n9983), .Z(n9632) );
  OAI21_X1 U10860 ( .B1(n9716), .B2(n9707), .A(n9632), .ZN(P1_U3553) );
  NAND2_X1 U10861 ( .A1(n9634), .A2(n9633), .ZN(n9717) );
  MUX2_X1 U10862 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9717), .S(n9983), .Z(n9635) );
  AOI21_X1 U10863 ( .B1(n9673), .B2(n9719), .A(n9635), .ZN(n9636) );
  INV_X1 U10864 ( .A(n9636), .ZN(P1_U3552) );
  INV_X1 U10865 ( .A(n9639), .ZN(n9643) );
  INV_X1 U10866 ( .A(n9944), .ZN(n9957) );
  AOI21_X1 U10867 ( .B1(n9957), .B2(n4847), .A(n9640), .ZN(n9641) );
  OAI211_X1 U10868 ( .C1(n9643), .C2(n9894), .A(n9642), .B(n9641), .ZN(n9724)
         );
  MUX2_X1 U10869 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9724), .S(n9983), .Z(
        P1_U3549) );
  AOI211_X1 U10870 ( .C1(n9646), .C2(n9949), .A(n9645), .B(n9644), .ZN(n9725)
         );
  MUX2_X1 U10871 ( .A(n10194), .B(n9725), .S(n9983), .Z(n9647) );
  OAI21_X1 U10872 ( .B1(n9728), .B2(n9707), .A(n9647), .ZN(P1_U3548) );
  OAI22_X1 U10873 ( .A1(n9649), .A2(n9950), .B1(n9648), .B2(n9952), .ZN(n9651)
         );
  OAI21_X1 U10874 ( .B1(n9654), .B2(n9894), .A(n9653), .ZN(n9729) );
  MUX2_X1 U10875 ( .A(n9729), .B(P1_REG1_REG_25__SCAN_IN), .S(n9981), .Z(n9655) );
  AOI21_X1 U10876 ( .B1(n9673), .B2(n9731), .A(n9655), .ZN(n9656) );
  INV_X1 U10877 ( .A(n9656), .ZN(P1_U3547) );
  INV_X1 U10878 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9662) );
  OAI211_X1 U10879 ( .C1(n9659), .C2(n9952), .A(n9658), .B(n9657), .ZN(n9660)
         );
  AOI21_X1 U10880 ( .B1(n9661), .B2(n9949), .A(n9660), .ZN(n9733) );
  MUX2_X1 U10881 ( .A(n9662), .B(n9733), .S(n9983), .Z(n9663) );
  OAI21_X1 U10882 ( .B1(n9736), .B2(n9707), .A(n9663), .ZN(P1_U3546) );
  AOI21_X1 U10883 ( .B1(n9957), .B2(n9665), .A(n9664), .ZN(n9666) );
  OAI211_X1 U10884 ( .C1(n9668), .C2(n9894), .A(n9667), .B(n9666), .ZN(n9737)
         );
  MUX2_X1 U10885 ( .A(n9737), .B(P1_REG1_REG_23__SCAN_IN), .S(n9981), .Z(
        P1_U3545) );
  OAI211_X1 U10886 ( .C1(n9671), .C2(n9894), .A(n9670), .B(n9669), .ZN(n9738)
         );
  MUX2_X1 U10887 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9738), .S(n9983), .Z(n9672) );
  AOI21_X1 U10888 ( .B1(n9673), .B2(n9740), .A(n9672), .ZN(n9674) );
  INV_X1 U10889 ( .A(n9674), .ZN(P1_U3544) );
  AOI21_X1 U10890 ( .B1(n9957), .B2(n9676), .A(n9675), .ZN(n9677) );
  OAI211_X1 U10891 ( .C1(n9894), .C2(n9679), .A(n9678), .B(n9677), .ZN(n9743)
         );
  MUX2_X1 U10892 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9743), .S(n9983), .Z(
        P1_U3543) );
  OAI22_X1 U10893 ( .A1(n9681), .A2(n9950), .B1(n9680), .B2(n9952), .ZN(n9682)
         );
  AOI211_X1 U10894 ( .C1(n9684), .C2(n9887), .A(n9683), .B(n9682), .ZN(n9685)
         );
  OAI21_X1 U10895 ( .B1(n9686), .B2(n9894), .A(n9685), .ZN(n9687) );
  INV_X1 U10896 ( .A(n9687), .ZN(n9744) );
  MUX2_X1 U10897 ( .A(n9688), .B(n9744), .S(n9983), .Z(n9689) );
  OAI21_X1 U10898 ( .B1(n9747), .B2(n9707), .A(n9689), .ZN(P1_U3542) );
  INV_X1 U10899 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10105) );
  OAI22_X1 U10900 ( .A1(n9691), .A2(n9950), .B1(n9690), .B2(n9952), .ZN(n9692)
         );
  INV_X1 U10901 ( .A(n9692), .ZN(n9694) );
  OAI211_X1 U10902 ( .C1(n9695), .C2(n9933), .A(n9694), .B(n9693), .ZN(n9696)
         );
  AOI21_X1 U10903 ( .B1(n9697), .B2(n9949), .A(n9696), .ZN(n9748) );
  MUX2_X1 U10904 ( .A(n10105), .B(n9748), .S(n9983), .Z(n9698) );
  OAI21_X1 U10905 ( .B1(n9751), .B2(n9707), .A(n9698), .ZN(P1_U3541) );
  AOI22_X1 U10906 ( .A1(n9891), .A2(n9699), .B1(n9781), .B2(n9918), .ZN(n9701)
         );
  OAI211_X1 U10907 ( .C1(n9702), .C2(n9933), .A(n9701), .B(n9700), .ZN(n9703)
         );
  AOI21_X1 U10908 ( .B1(n9704), .B2(n9949), .A(n9703), .ZN(n9752) );
  MUX2_X1 U10909 ( .A(n9705), .B(n9752), .S(n9983), .Z(n9706) );
  OAI21_X1 U10910 ( .B1(n9755), .B2(n9707), .A(n9706), .ZN(P1_U3540) );
  AOI21_X1 U10911 ( .B1(n9957), .B2(n9709), .A(n9708), .ZN(n9710) );
  OAI211_X1 U10912 ( .C1(n9712), .C2(n9894), .A(n9711), .B(n9710), .ZN(n9756)
         );
  MUX2_X1 U10913 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9756), .S(n9983), .Z(
        P1_U3539) );
  INV_X1 U10914 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9714) );
  MUX2_X1 U10915 ( .A(n9714), .B(n9713), .S(n9967), .Z(n9715) );
  OAI21_X1 U10916 ( .B1(n9716), .B2(n9754), .A(n9715), .ZN(P1_U3521) );
  MUX2_X1 U10917 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9717), .S(n9967), .Z(n9718) );
  AOI21_X1 U10918 ( .B1(n9741), .B2(n9719), .A(n9718), .ZN(n9720) );
  INV_X1 U10919 ( .A(n9720), .ZN(P1_U3520) );
  INV_X1 U10920 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9722) );
  MUX2_X1 U10921 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9724), .S(n9967), .Z(
        P1_U3517) );
  INV_X1 U10922 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9726) );
  MUX2_X1 U10923 ( .A(n9726), .B(n9725), .S(n9967), .Z(n9727) );
  OAI21_X1 U10924 ( .B1(n9728), .B2(n9754), .A(n9727), .ZN(P1_U3516) );
  MUX2_X1 U10925 ( .A(n9729), .B(P1_REG0_REG_25__SCAN_IN), .S(n9965), .Z(n9730) );
  AOI21_X1 U10926 ( .B1(n9741), .B2(n9731), .A(n9730), .ZN(n9732) );
  INV_X1 U10927 ( .A(n9732), .ZN(P1_U3515) );
  MUX2_X1 U10928 ( .A(n9734), .B(n9733), .S(n9967), .Z(n9735) );
  OAI21_X1 U10929 ( .B1(n9736), .B2(n9754), .A(n9735), .ZN(P1_U3514) );
  MUX2_X1 U10930 ( .A(n9737), .B(P1_REG0_REG_23__SCAN_IN), .S(n9965), .Z(
        P1_U3513) );
  MUX2_X1 U10931 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9738), .S(n9967), .Z(n9739) );
  AOI21_X1 U10932 ( .B1(n9741), .B2(n9740), .A(n9739), .ZN(n9742) );
  INV_X1 U10933 ( .A(n9742), .ZN(P1_U3512) );
  MUX2_X1 U10934 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9743), .S(n9967), .Z(
        P1_U3511) );
  INV_X1 U10935 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9745) );
  MUX2_X1 U10936 ( .A(n9745), .B(n9744), .S(n9967), .Z(n9746) );
  OAI21_X1 U10937 ( .B1(n9747), .B2(n9754), .A(n9746), .ZN(P1_U3510) );
  INV_X1 U10938 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9749) );
  MUX2_X1 U10939 ( .A(n9749), .B(n9748), .S(n9967), .Z(n9750) );
  OAI21_X1 U10940 ( .B1(n9751), .B2(n9754), .A(n9750), .ZN(P1_U3509) );
  MUX2_X1 U10941 ( .A(n10254), .B(n9752), .S(n9967), .Z(n9753) );
  OAI21_X1 U10942 ( .B1(n9755), .B2(n9754), .A(n9753), .ZN(P1_U3507) );
  MUX2_X1 U10943 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9756), .S(n9967), .Z(
        P1_U3504) );
  MUX2_X1 U10944 ( .A(n9757), .B(P1_D_REG_1__SCAN_IN), .S(n9859), .Z(P1_U3440)
         );
  MUX2_X1 U10945 ( .A(n9758), .B(P1_D_REG_0__SCAN_IN), .S(n9859), .Z(P1_U3439)
         );
  INV_X1 U10946 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9759) );
  NAND3_X1 U10947 ( .A1(n9759), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9761) );
  OAI22_X1 U10948 ( .A1(n9762), .A2(n9761), .B1(n9760), .B2(n9771), .ZN(n9763)
         );
  AOI21_X1 U10949 ( .B1(n9765), .B2(n9764), .A(n9763), .ZN(n9766) );
  INV_X1 U10950 ( .A(n9766), .ZN(P1_U3324) );
  OAI222_X1 U10951 ( .A1(n9771), .A2(n9770), .B1(n9769), .B2(n9768), .C1(
        P1_U3086), .C2(n9767), .ZN(P1_U3325) );
  INV_X1 U10952 ( .A(n9772), .ZN(n9773) );
  MUX2_X1 U10953 ( .A(n9773), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NOR2_X1 U10954 ( .A1(n9774), .A2(n10039), .ZN(n9776) );
  AOI211_X1 U10955 ( .C1(n9777), .C2(n10020), .A(n9776), .B(n9775), .ZN(n9779)
         );
  AOI22_X1 U10956 ( .A1(n10075), .A2(n9779), .B1(n8364), .B2(n6533), .ZN(
        P2_U3472) );
  INV_X1 U10957 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9778) );
  AOI22_X1 U10958 ( .A1(n10064), .A2(n9779), .B1(n9778), .B2(n10062), .ZN(
        P2_U3429) );
  AOI22_X1 U10959 ( .A1(n9891), .A2(n9781), .B1(n9780), .B2(n9918), .ZN(n9782)
         );
  OAI211_X1 U10960 ( .C1(n9784), .C2(n9944), .A(n9783), .B(n9782), .ZN(n9788)
         );
  AND3_X1 U10961 ( .A1(n9786), .A2(n9949), .A3(n9785), .ZN(n9787) );
  AOI211_X1 U10962 ( .C1(n9789), .C2(n9887), .A(n9788), .B(n9787), .ZN(n9790)
         );
  AOI22_X1 U10963 ( .A1(n9983), .A2(n9790), .B1(n9378), .B2(n9981), .ZN(
        P1_U3538) );
  INV_X1 U10964 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10252) );
  AOI22_X1 U10965 ( .A1(n9967), .A2(n9790), .B1(n10252), .B2(n9965), .ZN(
        P1_U3501) );
  XNOR2_X1 U10966 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XOR2_X1 U10967 ( .A(P1_RD_REG_SCAN_IN), .B(n4894), .Z(U126) );
  XNOR2_X1 U10968 ( .A(n9791), .B(n9795), .ZN(n9941) );
  OAI22_X1 U10969 ( .A1(n9793), .A2(n9950), .B1(n9792), .B2(n9952), .ZN(n9799)
         );
  NAND2_X1 U10970 ( .A1(n7335), .A2(n9794), .ZN(n9796) );
  XNOR2_X1 U10971 ( .A(n9796), .B(n9795), .ZN(n9797) );
  NOR2_X1 U10972 ( .A1(n9797), .A2(n9933), .ZN(n9798) );
  AOI211_X1 U10973 ( .C1(n9941), .C2(n9964), .A(n9799), .B(n9798), .ZN(n9938)
         );
  INV_X1 U10974 ( .A(n9800), .ZN(n9801) );
  AOI222_X1 U10975 ( .A1(n9802), .A2(n7133), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n9857), .C1(n9820), .C2(n9801), .ZN(n9807) );
  OAI211_X1 U10976 ( .C1(n9937), .C2(n9804), .A(n9803), .B(n9837), .ZN(n9936)
         );
  INV_X1 U10977 ( .A(n9936), .ZN(n9805) );
  AOI22_X1 U10978 ( .A1(n9941), .A2(n9852), .B1(n9851), .B2(n9805), .ZN(n9806)
         );
  OAI211_X1 U10979 ( .C1(n9857), .C2(n9938), .A(n9807), .B(n9806), .ZN(
        P1_U3282) );
  OAI21_X1 U10980 ( .B1(n9813), .B2(n9809), .A(n9808), .ZN(n9817) );
  OAI22_X1 U10981 ( .A1(n9811), .A2(n9952), .B1(n9810), .B2(n9950), .ZN(n9816)
         );
  XNOR2_X1 U10982 ( .A(n9812), .B(n9813), .ZN(n9907) );
  NOR2_X1 U10983 ( .A1(n9907), .A2(n9814), .ZN(n9815) );
  AOI211_X1 U10984 ( .C1(n9887), .C2(n9817), .A(n9816), .B(n9815), .ZN(n9906)
         );
  INV_X1 U10985 ( .A(n9818), .ZN(n9819) );
  AOI222_X1 U10986 ( .A1(n9904), .A2(n7133), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n9857), .C1(n9820), .C2(n9819), .ZN(n9826) );
  INV_X1 U10987 ( .A(n9907), .ZN(n9824) );
  AOI211_X1 U10988 ( .C1(n9904), .C2(n9823), .A(n9822), .B(n9821), .ZN(n9903)
         );
  AOI22_X1 U10989 ( .A1(n9824), .A2(n9852), .B1(n9851), .B2(n9903), .ZN(n9825)
         );
  OAI211_X1 U10990 ( .C1(n9857), .C2(n9906), .A(n9826), .B(n9825), .ZN(
        P1_U3286) );
  XOR2_X1 U10991 ( .A(n9827), .B(n9834), .Z(n9830) );
  AOI222_X1 U10992 ( .A1(n9887), .A2(n9830), .B1(n9829), .B2(n9891), .C1(n4429), .C2(n9918), .ZN(n9873) );
  NAND2_X1 U10993 ( .A1(n9857), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9831) );
  OAI21_X1 U10994 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(n9846), .A(n9831), .ZN(
        n9832) );
  AOI21_X1 U10995 ( .B1(n7133), .B2(n9833), .A(n9832), .ZN(n9843) );
  XNOR2_X1 U10996 ( .A(n9835), .B(n9834), .ZN(n9876) );
  INV_X1 U10997 ( .A(n9836), .ZN(n9838) );
  OAI211_X1 U10998 ( .C1(n9872), .C2(n9839), .A(n9838), .B(n9837), .ZN(n9871)
         );
  INV_X1 U10999 ( .A(n9871), .ZN(n9840) );
  AOI22_X1 U11000 ( .A1(n9876), .A2(n9841), .B1(n9851), .B2(n9840), .ZN(n9842)
         );
  OAI211_X1 U11001 ( .C1(n9857), .C2(n9873), .A(n9843), .B(n9842), .ZN(
        P1_U3290) );
  NAND2_X1 U11002 ( .A1(n9857), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9844) );
  OAI21_X1 U11003 ( .B1(n9846), .B2(n9845), .A(n9844), .ZN(n9847) );
  AOI21_X1 U11004 ( .B1(n7133), .B2(n9848), .A(n9847), .ZN(n9855) );
  INV_X1 U11005 ( .A(n9849), .ZN(n9850) );
  AOI22_X1 U11006 ( .A1(n9853), .A2(n9852), .B1(n9851), .B2(n9850), .ZN(n9854)
         );
  OAI211_X1 U11007 ( .C1(n9857), .C2(n9856), .A(n9855), .B(n9854), .ZN(
        P1_U3292) );
  AND2_X1 U11008 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9859), .ZN(P1_U3294) );
  INV_X1 U11009 ( .A(n9859), .ZN(n9858) );
  INV_X1 U11010 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10210) );
  NOR2_X1 U11011 ( .A1(n9858), .A2(n10210), .ZN(P1_U3295) );
  AND2_X1 U11012 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9859), .ZN(P1_U3296) );
  AND2_X1 U11013 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9859), .ZN(P1_U3297) );
  AND2_X1 U11014 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9859), .ZN(P1_U3298) );
  AND2_X1 U11015 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9859), .ZN(P1_U3299) );
  INV_X1 U11016 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10188) );
  NOR2_X1 U11017 ( .A1(n9858), .A2(n10188), .ZN(P1_U3300) );
  AND2_X1 U11018 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9859), .ZN(P1_U3301) );
  AND2_X1 U11019 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9859), .ZN(P1_U3302) );
  AND2_X1 U11020 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9859), .ZN(P1_U3303) );
  INV_X1 U11021 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10130) );
  NOR2_X1 U11022 ( .A1(n9858), .A2(n10130), .ZN(P1_U3304) );
  AND2_X1 U11023 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9859), .ZN(P1_U3305) );
  AND2_X1 U11024 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9859), .ZN(P1_U3306) );
  AND2_X1 U11025 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9859), .ZN(P1_U3307) );
  AND2_X1 U11026 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9859), .ZN(P1_U3308) );
  INV_X1 U11027 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10261) );
  NOR2_X1 U11028 ( .A1(n9858), .A2(n10261), .ZN(P1_U3309) );
  INV_X1 U11029 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10191) );
  NOR2_X1 U11030 ( .A1(n9858), .A2(n10191), .ZN(P1_U3310) );
  AND2_X1 U11031 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9859), .ZN(P1_U3311) );
  AND2_X1 U11032 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9859), .ZN(P1_U3312) );
  INV_X1 U11033 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10146) );
  NOR2_X1 U11034 ( .A1(n9858), .A2(n10146), .ZN(P1_U3313) );
  AND2_X1 U11035 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9859), .ZN(P1_U3314) );
  AND2_X1 U11036 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9859), .ZN(P1_U3315) );
  AND2_X1 U11037 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9859), .ZN(P1_U3316) );
  AND2_X1 U11038 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9859), .ZN(P1_U3317) );
  AND2_X1 U11039 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9859), .ZN(P1_U3318) );
  AND2_X1 U11040 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9859), .ZN(P1_U3319) );
  AND2_X1 U11041 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9859), .ZN(P1_U3320) );
  AND2_X1 U11042 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9859), .ZN(P1_U3321) );
  AND2_X1 U11043 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9859), .ZN(P1_U3322) );
  AND2_X1 U11044 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9859), .ZN(P1_U3323) );
  INV_X1 U11045 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9860) );
  AOI22_X1 U11046 ( .A1(n9967), .A2(n9861), .B1(n9860), .B2(n9965), .ZN(
        P1_U3456) );
  OAI22_X1 U11047 ( .A1(n9862), .A2(n9952), .B1(n9879), .B2(n9950), .ZN(n9864)
         );
  AOI211_X1 U11048 ( .C1(n9957), .C2(n9865), .A(n9864), .B(n9863), .ZN(n9866)
         );
  OAI21_X1 U11049 ( .B1(n9894), .B2(n9867), .A(n9866), .ZN(n9868) );
  AOI21_X1 U11050 ( .B1(n9869), .B2(n9887), .A(n9868), .ZN(n9968) );
  INV_X1 U11051 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9870) );
  AOI22_X1 U11052 ( .A1(n9967), .A2(n9968), .B1(n9870), .B2(n9965), .ZN(
        P1_U3459) );
  OAI21_X1 U11053 ( .B1(n9872), .B2(n9944), .A(n9871), .ZN(n9875) );
  INV_X1 U11054 ( .A(n9873), .ZN(n9874) );
  AOI211_X1 U11055 ( .C1(n9949), .C2(n9876), .A(n9875), .B(n9874), .ZN(n9969)
         );
  INV_X1 U11056 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9877) );
  AOI22_X1 U11057 ( .A1(n9967), .A2(n9969), .B1(n9877), .B2(n9965), .ZN(
        P1_U3462) );
  OAI22_X1 U11058 ( .A1(n9879), .A2(n9952), .B1(n9878), .B2(n9950), .ZN(n9880)
         );
  AOI21_X1 U11059 ( .B1(n9957), .B2(n9881), .A(n9880), .ZN(n9883) );
  OAI211_X1 U11060 ( .C1(n9884), .C2(n9894), .A(n9883), .B(n9882), .ZN(n9885)
         );
  AOI21_X1 U11061 ( .B1(n9887), .B2(n9886), .A(n9885), .ZN(n9970) );
  INV_X1 U11062 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9888) );
  AOI22_X1 U11063 ( .A1(n9967), .A2(n9970), .B1(n9888), .B2(n9965), .ZN(
        P1_U3465) );
  AOI22_X1 U11064 ( .A1(n9891), .A2(n9890), .B1(n9889), .B2(n9957), .ZN(n9893)
         );
  OAI211_X1 U11065 ( .C1(n9895), .C2(n9894), .A(n9893), .B(n9892), .ZN(n9896)
         );
  NOR2_X1 U11066 ( .A1(n9897), .A2(n9896), .ZN(n9971) );
  INV_X1 U11067 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10133) );
  AOI22_X1 U11068 ( .A1(n9967), .A2(n9971), .B1(n10133), .B2(n9965), .ZN(
        P1_U3468) );
  OAI21_X1 U11069 ( .B1(n9899), .B2(n9944), .A(n9898), .ZN(n9901) );
  AOI211_X1 U11070 ( .C1(n9949), .C2(n9902), .A(n9901), .B(n9900), .ZN(n9973)
         );
  AOI22_X1 U11071 ( .A1(n9967), .A2(n9973), .B1(n5203), .B2(n9965), .ZN(
        P1_U3471) );
  AOI21_X1 U11072 ( .B1(n9957), .B2(n9904), .A(n9903), .ZN(n9905) );
  OAI211_X1 U11073 ( .C1(n9907), .C2(n9960), .A(n9906), .B(n9905), .ZN(n9908)
         );
  INV_X1 U11074 ( .A(n9908), .ZN(n9974) );
  INV_X1 U11075 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9909) );
  AOI22_X1 U11076 ( .A1(n9967), .A2(n9974), .B1(n9909), .B2(n9965), .ZN(
        P1_U3474) );
  OAI21_X1 U11077 ( .B1(n9911), .B2(n9944), .A(n9910), .ZN(n9914) );
  INV_X1 U11078 ( .A(n9912), .ZN(n9913) );
  AOI211_X1 U11079 ( .C1(n9942), .C2(n9915), .A(n9914), .B(n9913), .ZN(n9975)
         );
  INV_X1 U11080 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9916) );
  AOI22_X1 U11081 ( .A1(n9967), .A2(n9975), .B1(n9916), .B2(n9965), .ZN(
        P1_U3477) );
  AOI22_X1 U11082 ( .A1(n9919), .A2(n9957), .B1(n9918), .B2(n9917), .ZN(n9920)
         );
  OAI211_X1 U11083 ( .C1(n9922), .C2(n9933), .A(n9921), .B(n9920), .ZN(n9923)
         );
  AOI21_X1 U11084 ( .B1(n9949), .B2(n9924), .A(n9923), .ZN(n9976) );
  INV_X1 U11085 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9925) );
  AOI22_X1 U11086 ( .A1(n9967), .A2(n9976), .B1(n9925), .B2(n9965), .ZN(
        P1_U3480) );
  OAI22_X1 U11087 ( .A1(n9927), .A2(n9952), .B1(n9926), .B2(n9950), .ZN(n9929)
         );
  AOI211_X1 U11088 ( .C1(n9957), .C2(n9930), .A(n9929), .B(n9928), .ZN(n9931)
         );
  OAI21_X1 U11089 ( .B1(n9933), .B2(n9932), .A(n9931), .ZN(n9934) );
  AOI21_X1 U11090 ( .B1(n9949), .B2(n9935), .A(n9934), .ZN(n9978) );
  AOI22_X1 U11091 ( .A1(n9967), .A2(n9978), .B1(n5298), .B2(n9965), .ZN(
        P1_U3483) );
  OAI21_X1 U11092 ( .B1(n9937), .B2(n9944), .A(n9936), .ZN(n9940) );
  INV_X1 U11093 ( .A(n9938), .ZN(n9939) );
  AOI211_X1 U11094 ( .C1(n9942), .C2(n9941), .A(n9940), .B(n9939), .ZN(n9979)
         );
  INV_X1 U11095 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10103) );
  AOI22_X1 U11096 ( .A1(n9967), .A2(n9979), .B1(n10103), .B2(n9965), .ZN(
        P1_U3486) );
  OAI21_X1 U11097 ( .B1(n9945), .B2(n9944), .A(n9943), .ZN(n9947) );
  AOI211_X1 U11098 ( .C1(n9949), .C2(n9948), .A(n9947), .B(n9946), .ZN(n9980)
         );
  INV_X1 U11099 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10262) );
  AOI22_X1 U11100 ( .A1(n9967), .A2(n9980), .B1(n10262), .B2(n9965), .ZN(
        P1_U3492) );
  OAI22_X1 U11101 ( .A1(n9953), .A2(n9952), .B1(n9951), .B2(n9950), .ZN(n9955)
         );
  AOI211_X1 U11102 ( .C1(n9957), .C2(n9956), .A(n9955), .B(n9954), .ZN(n9959)
         );
  OAI211_X1 U11103 ( .C1(n9961), .C2(n9960), .A(n9959), .B(n9958), .ZN(n9962)
         );
  AOI21_X1 U11104 ( .B1(n9964), .B2(n9963), .A(n9962), .ZN(n9982) );
  INV_X1 U11105 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9966) );
  AOI22_X1 U11106 ( .A1(n9967), .A2(n9982), .B1(n9966), .B2(n9965), .ZN(
        P1_U3495) );
  AOI22_X1 U11107 ( .A1(n9983), .A2(n9968), .B1(n6606), .B2(n9981), .ZN(
        P1_U3524) );
  AOI22_X1 U11108 ( .A1(n9983), .A2(n9969), .B1(n5136), .B2(n9981), .ZN(
        P1_U3525) );
  AOI22_X1 U11109 ( .A1(n9983), .A2(n9970), .B1(n5155), .B2(n9981), .ZN(
        P1_U3526) );
  AOI22_X1 U11110 ( .A1(n9983), .A2(n9971), .B1(n6611), .B2(n9981), .ZN(
        P1_U3527) );
  AOI22_X1 U11111 ( .A1(n9983), .A2(n9973), .B1(n9972), .B2(n9981), .ZN(
        P1_U3528) );
  AOI22_X1 U11112 ( .A1(n9983), .A2(n9974), .B1(n6633), .B2(n9981), .ZN(
        P1_U3529) );
  AOI22_X1 U11113 ( .A1(n9983), .A2(n9975), .B1(n5256), .B2(n9981), .ZN(
        P1_U3530) );
  AOI22_X1 U11114 ( .A1(n9983), .A2(n9976), .B1(n5281), .B2(n9981), .ZN(
        P1_U3531) );
  AOI22_X1 U11115 ( .A1(n9983), .A2(n9978), .B1(n9977), .B2(n9981), .ZN(
        P1_U3532) );
  AOI22_X1 U11116 ( .A1(n9983), .A2(n9979), .B1(n5320), .B2(n9981), .ZN(
        P1_U3533) );
  AOI22_X1 U11117 ( .A1(n9983), .A2(n9980), .B1(n5365), .B2(n9981), .ZN(
        P1_U3535) );
  AOI22_X1 U11118 ( .A1(n9983), .A2(n9982), .B1(n5386), .B2(n9981), .ZN(
        P1_U3536) );
  NAND2_X1 U11119 ( .A1(n9984), .A2(n6715), .ZN(n9986) );
  AOI21_X1 U11120 ( .B1(n9987), .B2(n9986), .A(n9985), .ZN(n9988) );
  AOI21_X1 U11121 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(P2_U3151), .A(n9988), 
        .ZN(n9994) );
  OAI211_X1 U11122 ( .C1(n9992), .C2(n9991), .A(n9990), .B(n10406), .ZN(n9993)
         );
  OAI211_X1 U11123 ( .C1(n9996), .C2(n9995), .A(n9994), .B(n9993), .ZN(n9997)
         );
  INV_X1 U11124 ( .A(n9997), .ZN(n10004) );
  INV_X1 U11125 ( .A(n9998), .ZN(n9999) );
  AOI21_X1 U11126 ( .B1(n6716), .B2(n10000), .A(n9999), .ZN(n10001) );
  OR2_X1 U11127 ( .A1(n10002), .A2(n10001), .ZN(n10003) );
  OAI211_X1 U11128 ( .C1(n10251), .C2(n10005), .A(n10004), .B(n10003), .ZN(
        P2_U3183) );
  OAI22_X1 U11129 ( .A1(n10007), .A2(n10045), .B1(n10006), .B2(n10039), .ZN(
        n10008) );
  NOR2_X1 U11130 ( .A1(n10009), .A2(n10008), .ZN(n10065) );
  INV_X1 U11131 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10117) );
  AOI22_X1 U11132 ( .A1(n10064), .A2(n10065), .B1(n10117), .B2(n10062), .ZN(
        P2_U3396) );
  NAND2_X1 U11133 ( .A1(n10010), .A2(n10020), .ZN(n10014) );
  NAND2_X1 U11134 ( .A1(n10011), .A2(n10061), .ZN(n10012) );
  AND3_X1 U11135 ( .A1(n10014), .A2(n10013), .A3(n10012), .ZN(n10066) );
  INV_X1 U11136 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10015) );
  AOI22_X1 U11137 ( .A1(n10064), .A2(n10066), .B1(n10015), .B2(n10062), .ZN(
        P2_U3399) );
  AOI22_X1 U11138 ( .A1(n10017), .A2(n10020), .B1(n10061), .B2(n10016), .ZN(
        n10018) );
  AND2_X1 U11139 ( .A1(n10019), .A2(n10018), .ZN(n10067) );
  AOI22_X1 U11140 ( .A1(n10064), .A2(n10067), .B1(n6102), .B2(n10062), .ZN(
        P2_U3402) );
  NAND2_X1 U11141 ( .A1(n10021), .A2(n10020), .ZN(n10024) );
  NAND2_X1 U11142 ( .A1(n10022), .A2(n10061), .ZN(n10023) );
  AND3_X1 U11143 ( .A1(n10025), .A2(n10024), .A3(n10023), .ZN(n10068) );
  INV_X1 U11144 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10026) );
  AOI22_X1 U11145 ( .A1(n10064), .A2(n10068), .B1(n10026), .B2(n10062), .ZN(
        P2_U3405) );
  OR2_X1 U11146 ( .A1(n10027), .A2(n10056), .ZN(n10030) );
  NAND2_X1 U11147 ( .A1(n10028), .A2(n10061), .ZN(n10029) );
  INV_X1 U11148 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10032) );
  AOI22_X1 U11149 ( .A1(n10064), .A2(n10069), .B1(n10032), .B2(n10062), .ZN(
        P2_U3408) );
  INV_X1 U11150 ( .A(n10033), .ZN(n10037) );
  OAI22_X1 U11151 ( .A1(n10035), .A2(n10056), .B1(n10034), .B2(n10039), .ZN(
        n10036) );
  NOR2_X1 U11152 ( .A1(n10037), .A2(n10036), .ZN(n10070) );
  INV_X1 U11153 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10038) );
  AOI22_X1 U11154 ( .A1(n10064), .A2(n10070), .B1(n10038), .B2(n10062), .ZN(
        P2_U3414) );
  OAI22_X1 U11155 ( .A1(n10041), .A2(n10045), .B1(n10040), .B2(n10039), .ZN(
        n10042) );
  NOR2_X1 U11156 ( .A1(n10043), .A2(n10042), .ZN(n10071) );
  INV_X1 U11157 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10044) );
  AOI22_X1 U11158 ( .A1(n10064), .A2(n10071), .B1(n10044), .B2(n10062), .ZN(
        P2_U3417) );
  NOR2_X1 U11159 ( .A1(n10046), .A2(n10045), .ZN(n10048) );
  AOI211_X1 U11160 ( .C1(n10061), .C2(n10049), .A(n10048), .B(n10047), .ZN(
        n10072) );
  INV_X1 U11161 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10050) );
  AOI22_X1 U11162 ( .A1(n10064), .A2(n10072), .B1(n10050), .B2(n10062), .ZN(
        P2_U3420) );
  NOR2_X1 U11163 ( .A1(n10051), .A2(n10056), .ZN(n10053) );
  AOI211_X1 U11164 ( .C1(n10061), .C2(n10054), .A(n10053), .B(n10052), .ZN(
        n10073) );
  INV_X1 U11165 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10055) );
  AOI22_X1 U11166 ( .A1(n10064), .A2(n10073), .B1(n10055), .B2(n10062), .ZN(
        P2_U3423) );
  NOR2_X1 U11167 ( .A1(n10057), .A2(n10056), .ZN(n10059) );
  AOI211_X1 U11168 ( .C1(n10061), .C2(n10060), .A(n10059), .B(n10058), .ZN(
        n10074) );
  INV_X1 U11169 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10063) );
  AOI22_X1 U11170 ( .A1(n10064), .A2(n10074), .B1(n10063), .B2(n10062), .ZN(
        P2_U3426) );
  AOI22_X1 U11171 ( .A1(n10075), .A2(n10065), .B1(n6078), .B2(n6533), .ZN(
        P2_U3461) );
  AOI22_X1 U11172 ( .A1(n10075), .A2(n10066), .B1(n6713), .B2(n6533), .ZN(
        P2_U3462) );
  AOI22_X1 U11173 ( .A1(n10075), .A2(n10067), .B1(n6790), .B2(n6533), .ZN(
        P2_U3463) );
  AOI22_X1 U11174 ( .A1(n10075), .A2(n10068), .B1(n6844), .B2(n6533), .ZN(
        P2_U3464) );
  AOI22_X1 U11175 ( .A1(n10075), .A2(n10069), .B1(n7082), .B2(n6533), .ZN(
        P2_U3465) );
  AOI22_X1 U11176 ( .A1(n10075), .A2(n10070), .B1(n6156), .B2(n6533), .ZN(
        P2_U3467) );
  AOI22_X1 U11177 ( .A1(n10075), .A2(n10071), .B1(n6168), .B2(n6533), .ZN(
        P2_U3468) );
  AOI22_X1 U11178 ( .A1(n10075), .A2(n10072), .B1(n7430), .B2(n6533), .ZN(
        P2_U3469) );
  AOI22_X1 U11179 ( .A1(n10075), .A2(n10073), .B1(n6198), .B2(n6533), .ZN(
        P2_U3470) );
  AOI22_X1 U11180 ( .A1(n10075), .A2(n10074), .B1(n8355), .B2(n6533), .ZN(
        P2_U3471) );
  INV_X1 U11181 ( .A(n10076), .ZN(n10077) );
  NAND2_X1 U11182 ( .A1(n10078), .A2(n10077), .ZN(n10079) );
  XOR2_X1 U11183 ( .A(n10251), .B(n10079), .Z(ADD_1068_U5) );
  XOR2_X1 U11184 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U11185 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10081), .A(n10080), 
        .ZN(n10083) );
  XOR2_X1 U11186 ( .A(n10083), .B(n10082), .Z(ADD_1068_U55) );
  XNOR2_X1 U11187 ( .A(n10085), .B(n10084), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11188 ( .A(n10087), .B(n10086), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11189 ( .A(n10089), .B(n10088), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11190 ( .A(n10091), .B(n10090), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11191 ( .A(n10093), .B(n10092), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11192 ( .A(n10095), .B(n10094), .ZN(ADD_1068_U61) );
  XOR2_X1 U11193 ( .A(n10097), .B(n10096), .Z(ADD_1068_U62) );
  XOR2_X1 U11194 ( .A(n10099), .B(n10098), .Z(ADD_1068_U63) );
  AOI22_X1 U11195 ( .A1(n8364), .A2(keyinput7), .B1(keyinput26), .B2(n10101), 
        .ZN(n10100) );
  OAI221_X1 U11196 ( .B1(n8364), .B2(keyinput7), .C1(n10101), .C2(keyinput26), 
        .A(n10100), .ZN(n10112) );
  AOI22_X1 U11197 ( .A1(n10103), .A2(keyinput119), .B1(keyinput9), .B2(n5252), 
        .ZN(n10102) );
  OAI221_X1 U11198 ( .B1(n10103), .B2(keyinput119), .C1(n5252), .C2(keyinput9), 
        .A(n10102), .ZN(n10111) );
  INV_X1 U11199 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n10106) );
  AOI22_X1 U11200 ( .A1(n10106), .A2(keyinput63), .B1(keyinput108), .B2(n10105), .ZN(n10104) );
  OAI221_X1 U11201 ( .B1(n10106), .B2(keyinput63), .C1(n10105), .C2(
        keyinput108), .A(n10104), .ZN(n10110) );
  XOR2_X1 U11202 ( .A(n5665), .B(keyinput8), .Z(n10108) );
  XNOR2_X1 U11203 ( .A(P1_REG2_REG_2__SCAN_IN), .B(keyinput109), .ZN(n10107)
         );
  NAND2_X1 U11204 ( .A1(n10108), .A2(n10107), .ZN(n10109) );
  NOR4_X1 U11205 ( .A1(n10112), .A2(n10111), .A3(n10110), .A4(n10109), .ZN(
        n10157) );
  AOI22_X1 U11206 ( .A1(n10115), .A2(keyinput85), .B1(keyinput104), .B2(n10114), .ZN(n10113) );
  OAI221_X1 U11207 ( .B1(n10115), .B2(keyinput85), .C1(n10114), .C2(
        keyinput104), .A(n10113), .ZN(n10124) );
  AOI22_X1 U11208 ( .A1(n5226), .A2(keyinput5), .B1(keyinput92), .B2(n5176), 
        .ZN(n10116) );
  OAI221_X1 U11209 ( .B1(n5226), .B2(keyinput5), .C1(n5176), .C2(keyinput92), 
        .A(n10116), .ZN(n10123) );
  XOR2_X1 U11210 ( .A(n9378), .B(keyinput13), .Z(n10121) );
  XOR2_X1 U11211 ( .A(n10117), .B(keyinput24), .Z(n10120) );
  XNOR2_X1 U11212 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput121), .ZN(n10119)
         );
  XNOR2_X1 U11213 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput122), .ZN(n10118) );
  NAND4_X1 U11214 ( .A1(n10121), .A2(n10120), .A3(n10119), .A4(n10118), .ZN(
        n10122) );
  NOR3_X1 U11215 ( .A1(n10124), .A2(n10123), .A3(n10122), .ZN(n10156) );
  INV_X1 U11216 ( .A(SI_30_), .ZN(n10126) );
  AOI22_X1 U11217 ( .A1(n10127), .A2(keyinput79), .B1(keyinput116), .B2(n10126), .ZN(n10125) );
  OAI221_X1 U11218 ( .B1(n10127), .B2(keyinput79), .C1(n10126), .C2(
        keyinput116), .A(n10125), .ZN(n10139) );
  AOI22_X1 U11219 ( .A1(n10130), .A2(keyinput35), .B1(keyinput82), .B2(n10129), 
        .ZN(n10128) );
  OAI221_X1 U11220 ( .B1(n10130), .B2(keyinput35), .C1(n10129), .C2(keyinput82), .A(n10128), .ZN(n10138) );
  INV_X1 U11221 ( .A(SI_13_), .ZN(n10132) );
  AOI22_X1 U11222 ( .A1(n10133), .A2(keyinput47), .B1(n10132), .B2(keyinput101), .ZN(n10131) );
  OAI221_X1 U11223 ( .B1(n10133), .B2(keyinput47), .C1(n10132), .C2(
        keyinput101), .A(n10131), .ZN(n10137) );
  XNOR2_X1 U11224 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput114), .ZN(n10135) );
  XNOR2_X1 U11225 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(keyinput33), .ZN(n10134)
         );
  NAND2_X1 U11226 ( .A1(n10135), .A2(n10134), .ZN(n10136) );
  NOR4_X1 U11227 ( .A1(n10139), .A2(n10138), .A3(n10137), .A4(n10136), .ZN(
        n10155) );
  AOI22_X1 U11228 ( .A1(n10141), .A2(keyinput75), .B1(keyinput124), .B2(n6115), 
        .ZN(n10140) );
  OAI221_X1 U11229 ( .B1(n10141), .B2(keyinput75), .C1(n6115), .C2(keyinput124), .A(n10140), .ZN(n10153) );
  AOI22_X1 U11230 ( .A1(n4894), .A2(keyinput113), .B1(keyinput65), .B2(n10143), 
        .ZN(n10142) );
  OAI221_X1 U11231 ( .B1(n4894), .B2(keyinput113), .C1(n10143), .C2(keyinput65), .A(n10142), .ZN(n10152) );
  INV_X1 U11232 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10145) );
  AOI22_X1 U11233 ( .A1(n10146), .A2(keyinput95), .B1(keyinput88), .B2(n10145), 
        .ZN(n10144) );
  OAI221_X1 U11234 ( .B1(n10146), .B2(keyinput95), .C1(n10145), .C2(keyinput88), .A(n10144), .ZN(n10151) );
  XOR2_X1 U11235 ( .A(n6698), .B(keyinput29), .Z(n10149) );
  XNOR2_X1 U11236 ( .A(P2_IR_REG_0__SCAN_IN), .B(keyinput94), .ZN(n10148) );
  NAND2_X1 U11237 ( .A1(n10149), .A2(n10148), .ZN(n10150) );
  NOR4_X1 U11238 ( .A1(n10153), .A2(n10152), .A3(n10151), .A4(n10150), .ZN(
        n10154) );
  NAND4_X1 U11239 ( .A1(n10157), .A2(n10156), .A3(n10155), .A4(n10154), .ZN(
        n10399) );
  AOI22_X1 U11240 ( .A1(n10159), .A2(keyinput39), .B1(keyinput106), .B2(n7187), 
        .ZN(n10158) );
  OAI221_X1 U11241 ( .B1(n10159), .B2(keyinput39), .C1(n7187), .C2(keyinput106), .A(n10158), .ZN(n10170) );
  AOI22_X1 U11242 ( .A1(n10162), .A2(keyinput111), .B1(keyinput22), .B2(n10161), .ZN(n10160) );
  OAI221_X1 U11243 ( .B1(n10162), .B2(keyinput111), .C1(n10161), .C2(
        keyinput22), .A(n10160), .ZN(n10169) );
  AOI22_X1 U11244 ( .A1(n5365), .A2(keyinput34), .B1(n10164), .B2(keyinput126), 
        .ZN(n10163) );
  OAI221_X1 U11245 ( .B1(n5365), .B2(keyinput34), .C1(n10164), .C2(keyinput126), .A(n10163), .ZN(n10168) );
  XOR2_X1 U11246 ( .A(n6102), .B(keyinput14), .Z(n10166) );
  XNOR2_X1 U11247 ( .A(SI_0_), .B(keyinput77), .ZN(n10165) );
  NAND2_X1 U11248 ( .A1(n10166), .A2(n10165), .ZN(n10167) );
  NOR4_X1 U11249 ( .A1(n10170), .A2(n10169), .A3(n10168), .A4(n10167), .ZN(
        n10218) );
  AOI22_X1 U11250 ( .A1(n10173), .A2(keyinput4), .B1(n10172), .B2(keyinput102), 
        .ZN(n10171) );
  OAI221_X1 U11251 ( .B1(n10173), .B2(keyinput4), .C1(n10172), .C2(keyinput102), .A(n10171), .ZN(n10186) );
  INV_X1 U11252 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U11253 ( .A1(n10176), .A2(keyinput36), .B1(n10175), .B2(keyinput72), 
        .ZN(n10174) );
  OAI221_X1 U11254 ( .B1(n10176), .B2(keyinput36), .C1(n10175), .C2(keyinput72), .A(n10174), .ZN(n10185) );
  AOI22_X1 U11255 ( .A1(n10179), .A2(keyinput27), .B1(n10178), .B2(keyinput20), 
        .ZN(n10177) );
  OAI221_X1 U11256 ( .B1(n10179), .B2(keyinput27), .C1(n10178), .C2(keyinput20), .A(n10177), .ZN(n10184) );
  INV_X1 U11257 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10180) );
  XOR2_X1 U11258 ( .A(n10180), .B(keyinput53), .Z(n10182) );
  XNOR2_X1 U11259 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput18), .ZN(n10181) );
  NAND2_X1 U11260 ( .A1(n10182), .A2(n10181), .ZN(n10183) );
  NOR4_X1 U11261 ( .A1(n10186), .A2(n10185), .A3(n10184), .A4(n10183), .ZN(
        n10217) );
  AOI22_X1 U11262 ( .A1(n10189), .A2(keyinput64), .B1(n10188), .B2(keyinput80), 
        .ZN(n10187) );
  OAI221_X1 U11263 ( .B1(n10189), .B2(keyinput64), .C1(n10188), .C2(keyinput80), .A(n10187), .ZN(n10200) );
  AOI22_X1 U11264 ( .A1(n10191), .A2(keyinput86), .B1(keyinput62), .B2(n6368), 
        .ZN(n10190) );
  OAI221_X1 U11265 ( .B1(n10191), .B2(keyinput86), .C1(n6368), .C2(keyinput62), 
        .A(n10190), .ZN(n10199) );
  INV_X1 U11266 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10193) );
  AOI22_X1 U11267 ( .A1(n10194), .A2(keyinput57), .B1(keyinput125), .B2(n10193), .ZN(n10192) );
  OAI221_X1 U11268 ( .B1(n10194), .B2(keyinput57), .C1(n10193), .C2(
        keyinput125), .A(n10192), .ZN(n10198) );
  XNOR2_X1 U11269 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(keyinput37), .ZN(n10196)
         );
  XNOR2_X1 U11270 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput115), .ZN(n10195) );
  NAND2_X1 U11271 ( .A1(n10196), .A2(n10195), .ZN(n10197) );
  NOR4_X1 U11272 ( .A1(n10200), .A2(n10199), .A3(n10198), .A4(n10197), .ZN(
        n10216) );
  INV_X1 U11273 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U11274 ( .A1(n10203), .A2(keyinput118), .B1(n10202), .B2(keyinput44), .ZN(n10201) );
  OAI221_X1 U11275 ( .B1(n10203), .B2(keyinput118), .C1(n10202), .C2(
        keyinput44), .A(n10201), .ZN(n10214) );
  INV_X1 U11276 ( .A(SI_21_), .ZN(n10205) );
  AOI22_X1 U11277 ( .A1(n10206), .A2(keyinput89), .B1(n10205), .B2(keyinput70), 
        .ZN(n10204) );
  OAI221_X1 U11278 ( .B1(n10206), .B2(keyinput89), .C1(n10205), .C2(keyinput70), .A(n10204), .ZN(n10213) );
  XNOR2_X1 U11279 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput74), .ZN(n10209) );
  XNOR2_X1 U11280 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput127), .ZN(n10208) );
  XNOR2_X1 U11281 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput19), .ZN(n10207)
         );
  NAND3_X1 U11282 ( .A1(n10209), .A2(n10208), .A3(n10207), .ZN(n10212) );
  XNOR2_X1 U11283 ( .A(n10210), .B(keyinput46), .ZN(n10211) );
  NOR4_X1 U11284 ( .A1(n10214), .A2(n10213), .A3(n10212), .A4(n10211), .ZN(
        n10215) );
  NAND4_X1 U11285 ( .A1(n10218), .A2(n10217), .A3(n10216), .A4(n10215), .ZN(
        n10398) );
  INV_X1 U11286 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n10220) );
  AOI22_X1 U11287 ( .A1(n5203), .A2(keyinput16), .B1(n10220), .B2(keyinput51), 
        .ZN(n10219) );
  OAI221_X1 U11288 ( .B1(n5203), .B2(keyinput16), .C1(n10220), .C2(keyinput51), 
        .A(n10219), .ZN(n10230) );
  XNOR2_X1 U11289 ( .A(n10221), .B(keyinput76), .ZN(n10229) );
  INV_X1 U11290 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10222) );
  XNOR2_X1 U11291 ( .A(keyinput107), .B(n10222), .ZN(n10228) );
  XNOR2_X1 U11292 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput52), .ZN(n10226) );
  XNOR2_X1 U11293 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput43), .ZN(n10225) );
  XNOR2_X1 U11294 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput71), .ZN(n10224)
         );
  XNOR2_X1 U11295 ( .A(SI_5_), .B(keyinput100), .ZN(n10223) );
  NAND4_X1 U11296 ( .A1(n10226), .A2(n10225), .A3(n10224), .A4(n10223), .ZN(
        n10227) );
  NOR4_X1 U11297 ( .A1(n10230), .A2(n10229), .A3(n10228), .A4(n10227), .ZN(
        n10396) );
  AOI22_X1 U11298 ( .A1(n10232), .A2(keyinput10), .B1(keyinput117), .B2(n5281), 
        .ZN(n10231) );
  OAI221_X1 U11299 ( .B1(n10232), .B2(keyinput10), .C1(n5281), .C2(keyinput117), .A(n10231), .ZN(n10243) );
  AOI22_X1 U11300 ( .A1(n6779), .A2(keyinput49), .B1(n10234), .B2(keyinput54), 
        .ZN(n10233) );
  OAI221_X1 U11301 ( .B1(n6779), .B2(keyinput49), .C1(n10234), .C2(keyinput54), 
        .A(n10233), .ZN(n10242) );
  AOI22_X1 U11302 ( .A1(n10237), .A2(keyinput32), .B1(keyinput23), .B2(n10236), 
        .ZN(n10235) );
  OAI221_X1 U11303 ( .B1(n10237), .B2(keyinput32), .C1(n10236), .C2(keyinput23), .A(n10235), .ZN(n10241) );
  XOR2_X1 U11304 ( .A(n7656), .B(keyinput60), .Z(n10239) );
  XNOR2_X1 U11305 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput90), .ZN(n10238) );
  NAND2_X1 U11306 ( .A1(n10239), .A2(n10238), .ZN(n10240) );
  NOR4_X1 U11307 ( .A1(n10243), .A2(n10242), .A3(n10241), .A4(n10240), .ZN(
        n10395) );
  INV_X1 U11308 ( .A(SI_18_), .ZN(n10246) );
  AOI22_X1 U11309 ( .A1(n10246), .A2(keyinput40), .B1(keyinput56), .B2(n10245), 
        .ZN(n10244) );
  OAI221_X1 U11310 ( .B1(n10246), .B2(keyinput40), .C1(n10245), .C2(keyinput56), .A(n10244), .ZN(n10258) );
  AOI22_X1 U11311 ( .A1(n10249), .A2(keyinput0), .B1(keyinput97), .B2(n10248), 
        .ZN(n10247) );
  OAI221_X1 U11312 ( .B1(n10249), .B2(keyinput0), .C1(n10248), .C2(keyinput97), 
        .A(n10247), .ZN(n10257) );
  AOI22_X1 U11313 ( .A1(n10252), .A2(keyinput11), .B1(keyinput93), .B2(n10251), 
        .ZN(n10250) );
  OAI221_X1 U11314 ( .B1(n10252), .B2(keyinput11), .C1(n10251), .C2(keyinput93), .A(n10250), .ZN(n10256) );
  AOI22_X1 U11315 ( .A1(n10254), .A2(keyinput98), .B1(keyinput30), .B2(n7430), 
        .ZN(n10253) );
  OAI221_X1 U11316 ( .B1(n10254), .B2(keyinput98), .C1(n7430), .C2(keyinput30), 
        .A(n10253), .ZN(n10255) );
  OR4_X1 U11317 ( .A1(n10258), .A2(n10257), .A3(n10256), .A4(n10255), .ZN(
        n10277) );
  AOI22_X1 U11318 ( .A1(n7081), .A2(keyinput59), .B1(n6254), .B2(keyinput2), 
        .ZN(n10259) );
  OAI221_X1 U11319 ( .B1(n7081), .B2(keyinput59), .C1(n6254), .C2(keyinput2), 
        .A(n10259), .ZN(n10276) );
  AOI22_X1 U11320 ( .A1(n10262), .A2(keyinput42), .B1(n10261), .B2(keyinput1), 
        .ZN(n10260) );
  OAI221_X1 U11321 ( .B1(n10262), .B2(keyinput42), .C1(n10261), .C2(keyinput1), 
        .A(n10260), .ZN(n10275) );
  INV_X1 U11322 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10264) );
  AOI22_X1 U11323 ( .A1(n10264), .A2(keyinput55), .B1(keyinput12), .B2(n9563), 
        .ZN(n10263) );
  OAI221_X1 U11324 ( .B1(n10264), .B2(keyinput55), .C1(n9563), .C2(keyinput12), 
        .A(n10263), .ZN(n10273) );
  AOI22_X1 U11325 ( .A1(n10267), .A2(keyinput6), .B1(keyinput15), .B2(n10266), 
        .ZN(n10265) );
  OAI221_X1 U11326 ( .B1(n10267), .B2(keyinput6), .C1(n10266), .C2(keyinput15), 
        .A(n10265), .ZN(n10272) );
  XNOR2_X1 U11327 ( .A(n10268), .B(keyinput120), .ZN(n10271) );
  XNOR2_X1 U11328 ( .A(n10269), .B(keyinput25), .ZN(n10270) );
  OR4_X1 U11329 ( .A1(n10273), .A2(n10272), .A3(n10271), .A4(n10270), .ZN(
        n10274) );
  NOR4_X1 U11330 ( .A1(n10277), .A2(n10276), .A3(n10275), .A4(n10274), .ZN(
        n10327) );
  AOI22_X1 U11331 ( .A1(n10280), .A2(keyinput96), .B1(keyinput17), .B2(n10279), 
        .ZN(n10278) );
  OAI221_X1 U11332 ( .B1(n10280), .B2(keyinput96), .C1(n10279), .C2(keyinput17), .A(n10278), .ZN(n10292) );
  AOI22_X1 U11333 ( .A1(n10283), .A2(keyinput67), .B1(keyinput58), .B2(n10282), 
        .ZN(n10281) );
  OAI221_X1 U11334 ( .B1(n10283), .B2(keyinput67), .C1(n10282), .C2(keyinput58), .A(n10281), .ZN(n10291) );
  AOI22_X1 U11335 ( .A1(n10286), .A2(keyinput73), .B1(keyinput123), .B2(n10285), .ZN(n10284) );
  OAI221_X1 U11336 ( .B1(n10286), .B2(keyinput73), .C1(n10285), .C2(
        keyinput123), .A(n10284), .ZN(n10290) );
  AOI22_X1 U11337 ( .A1(n6598), .A2(keyinput81), .B1(keyinput99), .B2(n10288), 
        .ZN(n10287) );
  OAI221_X1 U11338 ( .B1(n6598), .B2(keyinput81), .C1(n10288), .C2(keyinput99), 
        .A(n10287), .ZN(n10289) );
  NOR4_X1 U11339 ( .A1(n10292), .A2(n10291), .A3(n10290), .A4(n10289), .ZN(
        n10326) );
  INV_X1 U11340 ( .A(keyinput91), .ZN(n10297) );
  AOI22_X1 U11341 ( .A1(n10295), .A2(keyinput31), .B1(keyinput21), .B2(n10294), 
        .ZN(n10293) );
  OAI221_X1 U11342 ( .B1(n10295), .B2(keyinput31), .C1(n10294), .C2(keyinput21), .A(n10293), .ZN(n10296) );
  AOI221_X1 U11343 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n10297), .C1(n6845), 
        .C2(keyinput91), .A(n10296), .ZN(n10325) );
  AOI22_X1 U11344 ( .A1(n10299), .A2(keyinput87), .B1(keyinput48), .B2(n6714), 
        .ZN(n10298) );
  OAI221_X1 U11345 ( .B1(n10299), .B2(keyinput87), .C1(n6714), .C2(keyinput48), 
        .A(n10298), .ZN(n10323) );
  AOI22_X1 U11346 ( .A1(n7071), .A2(keyinput45), .B1(n10301), .B2(keyinput50), 
        .ZN(n10300) );
  OAI221_X1 U11347 ( .B1(n7071), .B2(keyinput45), .C1(n10301), .C2(keyinput50), 
        .A(n10300), .ZN(n10315) );
  XNOR2_X1 U11348 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput110), .ZN(n10305) );
  XNOR2_X1 U11349 ( .A(SI_4_), .B(keyinput112), .ZN(n10304) );
  XNOR2_X1 U11350 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput66), .ZN(n10303) );
  XNOR2_X1 U11351 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput68), .ZN(n10302) );
  NAND4_X1 U11352 ( .A1(n10305), .A2(n10304), .A3(n10303), .A4(n10302), .ZN(
        n10314) );
  XNOR2_X1 U11353 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput61), .ZN(n10309) );
  XNOR2_X1 U11354 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput105), .ZN(n10308) );
  XNOR2_X1 U11355 ( .A(P2_REG1_REG_0__SCAN_IN), .B(keyinput84), .ZN(n10307) );
  XNOR2_X1 U11356 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(keyinput41), .ZN(n10306)
         );
  NAND4_X1 U11357 ( .A1(n10309), .A2(n10308), .A3(n10307), .A4(n10306), .ZN(
        n10313) );
  XNOR2_X1 U11358 ( .A(P1_REG0_REG_24__SCAN_IN), .B(keyinput28), .ZN(n10311)
         );
  XNOR2_X1 U11359 ( .A(keyinput69), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n10310)
         );
  OAI211_X1 U11360 ( .C1(n10391), .C2(keyinput38), .A(n10311), .B(n10310), 
        .ZN(n10312) );
  OR4_X1 U11361 ( .A1(n10315), .A2(n10314), .A3(n10313), .A4(n10312), .ZN(
        n10322) );
  AOI22_X1 U11362 ( .A1(n6600), .A2(keyinput83), .B1(keyinput3), .B2(n10317), 
        .ZN(n10316) );
  OAI221_X1 U11363 ( .B1(n6600), .B2(keyinput83), .C1(n10317), .C2(keyinput3), 
        .A(n10316), .ZN(n10321) );
  INV_X1 U11364 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U11365 ( .A1(P1_U3086), .A2(keyinput103), .B1(keyinput78), .B2(
        n10319), .ZN(n10318) );
  OAI221_X1 U11366 ( .B1(P1_U3086), .B2(keyinput103), .C1(n10319), .C2(
        keyinput78), .A(n10318), .ZN(n10320) );
  NOR4_X1 U11367 ( .A1(n10323), .A2(n10322), .A3(n10321), .A4(n10320), .ZN(
        n10324) );
  AND4_X1 U11368 ( .A1(n10327), .A2(n10326), .A3(n10325), .A4(n10324), .ZN(
        n10394) );
  NAND4_X1 U11369 ( .A1(keyinput58), .A2(keyinput96), .A3(keyinput99), .A4(
        keyinput73), .ZN(n10390) );
  NOR2_X1 U11370 ( .A1(keyinput17), .A2(keyinput67), .ZN(n10328) );
  NAND3_X1 U11371 ( .A1(keyinput100), .A2(keyinput81), .A3(n10328), .ZN(n10389) );
  NOR2_X1 U11372 ( .A1(keyinput87), .A2(keyinput59), .ZN(n10329) );
  NAND3_X1 U11373 ( .A1(keyinput15), .A2(keyinput105), .A3(n10329), .ZN(n10330) );
  NOR3_X1 U11374 ( .A1(keyinput56), .A2(keyinput41), .A3(n10330), .ZN(n10338)
         );
  NAND4_X1 U11375 ( .A1(keyinput97), .A2(keyinput103), .A3(keyinput78), .A4(
        keyinput68), .ZN(n10336) );
  NOR3_X1 U11376 ( .A1(keyinput123), .A2(keyinput83), .A3(keyinput0), .ZN(
        n10331) );
  NAND2_X1 U11377 ( .A1(keyinput84), .A2(n10331), .ZN(n10335) );
  NAND4_X1 U11378 ( .A1(keyinput25), .A2(keyinput98), .A3(keyinput30), .A4(
        keyinput45), .ZN(n10334) );
  NOR3_X1 U11379 ( .A1(keyinput3), .A2(keyinput50), .A3(keyinput120), .ZN(
        n10332) );
  NAND2_X1 U11380 ( .A1(keyinput6), .A2(n10332), .ZN(n10333) );
  NOR4_X1 U11381 ( .A1(n10336), .A2(n10335), .A3(n10334), .A4(n10333), .ZN(
        n10337) );
  NAND4_X1 U11382 ( .A1(keyinput48), .A2(keyinput40), .A3(n10338), .A4(n10337), 
        .ZN(n10388) );
  NAND2_X1 U11383 ( .A1(keyinput21), .A2(keyinput31), .ZN(n10339) );
  NOR3_X1 U11384 ( .A1(keyinput91), .A2(keyinput61), .A3(n10339), .ZN(n10340)
         );
  NAND4_X1 U11385 ( .A1(keyinput74), .A2(keyinput112), .A3(keyinput69), .A4(
        n10340), .ZN(n10354) );
  NOR3_X1 U11386 ( .A1(keyinput12), .A2(keyinput11), .A3(keyinput55), .ZN(
        n10341) );
  NAND2_X1 U11387 ( .A1(keyinput1), .A2(n10341), .ZN(n10353) );
  INV_X1 U11388 ( .A(keyinput42), .ZN(n10342) );
  NAND4_X1 U11389 ( .A1(keyinput110), .A2(keyinput66), .A3(keyinput28), .A4(
        n10342), .ZN(n10352) );
  NAND2_X1 U11390 ( .A1(keyinput10), .A2(keyinput32), .ZN(n10343) );
  NOR3_X1 U11391 ( .A1(keyinput54), .A2(keyinput23), .A3(n10343), .ZN(n10350)
         );
  INV_X1 U11392 ( .A(keyinput90), .ZN(n10344) );
  NOR4_X1 U11393 ( .A1(keyinput93), .A2(keyinput60), .A3(keyinput49), .A4(
        n10344), .ZN(n10349) );
  NAND2_X1 U11394 ( .A1(keyinput76), .A2(keyinput51), .ZN(n10345) );
  NOR3_X1 U11395 ( .A1(keyinput71), .A2(keyinput107), .A3(n10345), .ZN(n10348)
         );
  INV_X1 U11396 ( .A(keyinput52), .ZN(n10346) );
  NOR4_X1 U11397 ( .A1(keyinput117), .A2(keyinput43), .A3(keyinput16), .A4(
        n10346), .ZN(n10347) );
  NAND4_X1 U11398 ( .A1(n10350), .A2(n10349), .A3(n10348), .A4(n10347), .ZN(
        n10351) );
  NOR4_X1 U11399 ( .A1(n10354), .A2(n10353), .A3(n10352), .A4(n10351), .ZN(
        n10386) );
  NOR2_X1 U11400 ( .A1(keyinput85), .A2(keyinput5), .ZN(n10355) );
  NAND3_X1 U11401 ( .A1(keyinput122), .A2(keyinput104), .A3(n10355), .ZN(
        n10362) );
  INV_X1 U11402 ( .A(keyinput108), .ZN(n10356) );
  NAND4_X1 U11403 ( .A1(keyinput13), .A2(keyinput121), .A3(keyinput24), .A4(
        n10356), .ZN(n10361) );
  NOR2_X1 U11404 ( .A1(keyinput75), .A2(keyinput95), .ZN(n10357) );
  NAND3_X1 U11405 ( .A1(keyinput29), .A2(keyinput124), .A3(n10357), .ZN(n10360) );
  INV_X1 U11406 ( .A(keyinput65), .ZN(n10358) );
  NAND4_X1 U11407 ( .A1(keyinput113), .A2(keyinput114), .A3(keyinput94), .A4(
        n10358), .ZN(n10359) );
  NOR4_X1 U11408 ( .A1(n10362), .A2(n10361), .A3(n10360), .A4(n10359), .ZN(
        n10385) );
  NOR4_X1 U11409 ( .A1(keyinput9), .A2(keyinput8), .A3(keyinput26), .A4(
        keyinput63), .ZN(n10368) );
  NAND2_X1 U11410 ( .A1(keyinput7), .A2(keyinput119), .ZN(n10363) );
  NOR3_X1 U11411 ( .A1(keyinput2), .A2(keyinput109), .A3(n10363), .ZN(n10367)
         );
  NOR4_X1 U11412 ( .A1(keyinput82), .A2(keyinput79), .A3(keyinput116), .A4(
        keyinput33), .ZN(n10366) );
  NAND2_X1 U11413 ( .A1(keyinput101), .A2(keyinput47), .ZN(n10364) );
  NOR3_X1 U11414 ( .A1(keyinput92), .A2(keyinput35), .A3(n10364), .ZN(n10365)
         );
  AND4_X1 U11415 ( .A1(n10368), .A2(n10367), .A3(n10366), .A4(n10365), .ZN(
        n10384) );
  NAND2_X1 U11416 ( .A1(keyinput126), .A2(keyinput34), .ZN(n10369) );
  NOR3_X1 U11417 ( .A1(keyinput88), .A2(keyinput111), .A3(n10369), .ZN(n10370)
         );
  NAND3_X1 U11418 ( .A1(keyinput22), .A2(keyinput77), .A3(n10370), .ZN(n10382)
         );
  NAND4_X1 U11419 ( .A1(keyinput62), .A2(keyinput57), .A3(keyinput125), .A4(
        keyinput115), .ZN(n10371) );
  NOR3_X1 U11420 ( .A1(keyinput37), .A2(keyinput64), .A3(n10371), .ZN(n10380)
         );
  NOR2_X1 U11421 ( .A1(keyinput20), .A2(keyinput27), .ZN(n10372) );
  NAND3_X1 U11422 ( .A1(keyinput53), .A2(keyinput4), .A3(n10372), .ZN(n10378)
         );
  NAND4_X1 U11423 ( .A1(keyinput106), .A2(keyinput36), .A3(keyinput72), .A4(
        keyinput18), .ZN(n10377) );
  INV_X1 U11424 ( .A(keyinput118), .ZN(n10373) );
  NAND4_X1 U11425 ( .A1(keyinput46), .A2(keyinput44), .A3(keyinput19), .A4(
        n10373), .ZN(n10376) );
  NOR3_X1 U11426 ( .A1(keyinput70), .A2(keyinput127), .A3(keyinput89), .ZN(
        n10374) );
  NAND2_X1 U11427 ( .A1(keyinput80), .A2(n10374), .ZN(n10375) );
  NOR4_X1 U11428 ( .A1(n10378), .A2(n10377), .A3(n10376), .A4(n10375), .ZN(
        n10379) );
  NAND4_X1 U11429 ( .A1(keyinput102), .A2(keyinput86), .A3(n10380), .A4(n10379), .ZN(n10381) );
  NOR4_X1 U11430 ( .A1(keyinput14), .A2(keyinput39), .A3(n10382), .A4(n10381), 
        .ZN(n10383) );
  NAND4_X1 U11431 ( .A1(n10386), .A2(n10385), .A3(n10384), .A4(n10383), .ZN(
        n10387) );
  NOR4_X1 U11432 ( .A1(n10390), .A2(n10389), .A3(n10388), .A4(n10387), .ZN(
        n10392) );
  OAI21_X1 U11433 ( .B1(keyinput38), .B2(n10392), .A(n10391), .ZN(n10393) );
  NAND4_X1 U11434 ( .A1(n10396), .A2(n10395), .A3(n10394), .A4(n10393), .ZN(
        n10397) );
  NOR3_X1 U11435 ( .A1(n10399), .A2(n10398), .A3(n10397), .ZN(n10423) );
  OAI21_X1 U11436 ( .B1(n10402), .B2(n10401), .A(n10400), .ZN(n10403) );
  AOI22_X1 U11437 ( .A1(n10405), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n10404), 
        .B2(n10403), .ZN(n10414) );
  OAI211_X1 U11438 ( .C1(n10409), .C2(n10408), .A(n10407), .B(n10406), .ZN(
        n10413) );
  NAND2_X1 U11439 ( .A1(n10411), .A2(n10410), .ZN(n10412) );
  AND3_X1 U11440 ( .A1(n10414), .A2(n10413), .A3(n10412), .ZN(n10421) );
  OAI21_X1 U11441 ( .B1(n10417), .B2(n10416), .A(n10415), .ZN(n10418) );
  NAND2_X1 U11442 ( .A1(n10419), .A2(n10418), .ZN(n10420) );
  OAI211_X1 U11443 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6890), .A(n10421), .B(
        n10420), .ZN(n10422) );
  XOR2_X1 U11444 ( .A(n10423), .B(n10422), .Z(P2_U3184) );
  XOR2_X1 U11445 ( .A(n10424), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1068_U50) );
  NOR2_X1 U11446 ( .A1(n10426), .A2(n10425), .ZN(n10427) );
  XOR2_X1 U11447 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10427), .Z(ADD_1068_U51) );
  XOR2_X1 U11448 ( .A(n10428), .B(P2_ADDR_REG_9__SCAN_IN), .Z(ADD_1068_U47) );
  XOR2_X1 U11449 ( .A(n10429), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1068_U49) );
  XOR2_X1 U11450 ( .A(n10430), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1068_U48) );
  XOR2_X1 U11451 ( .A(n10432), .B(n10431), .Z(ADD_1068_U54) );
  XOR2_X1 U11452 ( .A(n10434), .B(n10433), .Z(ADD_1068_U53) );
  XNOR2_X1 U11453 ( .A(n10436), .B(n10435), .ZN(ADD_1068_U52) );
  INV_X1 U4940 ( .A(n5827), .ZN(n5981) );
  CLKBUF_X1 U4943 ( .A(n6550), .Z(n4435) );
  NAND2_X1 U4949 ( .A1(n8041), .A2(n8042), .ZN(n8083) );
  INV_X2 U4961 ( .A(n6667), .ZN(n5545) );
  AND3_X1 U4981 ( .A1(n5172), .A2(n5171), .A3(n5170), .ZN(n7316) );
  CLKBUF_X3 U4995 ( .A(n6550), .Z(n4436) );
  CLKBUF_X1 U5034 ( .A(n5717), .Z(n4443) );
endmodule

